// Benchmark "testing" written by ABC on Thu Oct  8 22:16:59 2020

module testing ( 
    G5873, G5872, G5871, G5870, G5869, G5868, G5806, G5805, G5804, G5803,
    G5802, G5801, G5739, G5738, G5737, G5736, G5735, G5734, G5672, G5671,
    G5670, G5669, G5668, G5667, G5605, G5604, G5603, G5602, G5601, G5600,
    G5538, G5537, G5536, G5535, G5534, G5533, G5471, G5470, G5469, G5468,
    G5467, G5466, G5404, G5403, G5402, G5401, G5400, G5399, G5337, G5336,
    G5335, G5334, G5333, G5332, G5270, G5269, G5268, G5267, G5266, G5265,
    G5203, G5202, G5201, G5200, G5199, G5198, G5136, G5135, G5134, G5133,
    G5132, G5131, G5069, G5068, G5067, G5066, G5065, G5064, G5002, G5001,
    G5000, G4999, G4998, G4997, G4935, G4934, G4933, G4932, G4931, G4930,
    G4868, G4867, G4866, G4865, G4864, G4863, G4801, G4800, G4799, G4798,
    G4797, G4796, G4734, G4733, G4732, G4731, G4730, G4729, G4667, G4666,
    G4665, G4664, G4663, G4662, G4600, G4599, G4598, G4597, G4596, G4595,
    G4533, G4532, G4531, G4530, G4529, G4528, G4466, G4465, G4464, G4463,
    G4462, G4461, G4399, G4398, G4397, G4396, G4395, G4394, G4332, G4331,
    G4330, G4329, G4328, G4327, G4265, G4264, G4263, G4262, G4261, G4260,
    G4198, G4197, G4196, G4195, G4194, G4193, G4131, G4130, G4129, G4128,
    G4127, G4126, G4064, G4063, G4062, G4061, G4060, G4059, G3997, G3996,
    G3995, G3994, G3993, G3992, G3930, G3929, G3928, G3927, G3926, G3925,
    G3863, G3862, G3861, G3860, G3859, G3858, G3796, G3795, G3794, G3793,
    G3792, G3791, G3729, G3728, G3727, G3726, G3725, G3724, G3662, G3661,
    G3660, G3659, G3658, G3657, G3595, G3594, G3593, G3592, G3591, G3590,
    G3528, G3527, G3526, G3525, G3524, G3523, G3461, G3460, G3459, G3458,
    G3457, G3456, G3394, G3393, G3392, G3391, G3390, G3389, G3327, G3326,
    G3325, G3324, G3323, G3322, G3260, G3259, G3258, G3257, G3256, G3255,
    G3193, G3192, G3191, G3190, G3189, G3188, G3126, G3125, G3124, G3123,
    G3122, G3121, G3059, G3058, G3057, G3056, G3055, G3054, G2992, G2991,
    G2990, G2989, G2988, G2987, G2925, G2924, G2923, G2922, G2921, G2920,
    G2858, G2857, G2856, G2855, G2854, G2853, G2791, G2790, G2789, G2788,
    G2787, G2786, G2724, G2723, G2722, G2721, G2720, G2719, G2657, G2656,
    G2655, G2654, G2653, G2652, G2590, G2589, G2588, G2587, G2586, G2585,
    G2523, G2522, G2521, G2520, G2519, G2518, G2456, G2455, G2454, G2453,
    G2452, G2451, G2389, G2388, G2387, G2386, G2385, G2384, G2322, G2321,
    G2320, G2319, G2318, G2317, G2255, G2254, G2253, G2252, G2251, G2250,
    G2188, G2187, G2186, G2185, G2184, G2183, G2121, G2120, G2119, G2118,
    G2117, G2116, G2054, G2053, G2052, G2051, G2050, G2049, G1987, G1986,
    G1985, G1984, G1983, G1982, G1920, G1919, G1918, G1917, G1916, G1915,
    G1853, G1852, G1851, G1850, G1849, G1848, G1786, G1785, G1784, G1783,
    G1782, G1781, G1719, G1718, G1717, G1716, G1715, G1714, G1652, G1651,
    G1650, G1649, G1648, G1647, G1585, G1584, G1583, G1582, G1581, G1580,
    G1518, G1517, G1516, G1515, G1514, G1513, G1451, G1450, G1449, G1448,
    G1447, G1446, G1384, G1383, G1382, G1381, G1380, G1379, G1317, G1316,
    G1315, G1314, G1313, G1312, G1250, G1249, G1248, G1247, G1246, G1245,
    G1183, G1182, G1181, G1180, G1179, G1178, G1116, G1115, G1114, G1113,
    G1112, G1111, G1049, G1048, G1047, G1046, G1045, G1044, G982, G981,
    G980, G979, G978, G977, G915, G914, G913, G912, G911, G910, G848, G847,
    G846, G845, G844, G843, G781, G780, G779, G778, G777, G776, G714, G713,
    G712, G711, G710, G709, G647, G646, G645, G644, G643, G642, G580, G579,
    G578, G577, G576, G575, G513, G512, G511, G510, G509, G508, G446, G445,
    G444, G443, G442, G441, G379, G378, G377, G376, G375, G374, G312, G311,
    G310, G309, G308, G307, G245, G244, G243, G242, G241, G240, G178, G177,
    G176, G175, G174, G173, G111, G110, G109, G108, G107, G106, G44, G43,
    G42, G41, G40, G39, F9976, F9975, F9974, F9973, F9972, F9971, F9909,
    F9908, F9907, F9906, F9905, F9904, F9842, F9841, F9840, F9839, F9838,
    F9837, F9775, F9774, F9773, F9772, F9771, F9770, F9708, F9707, F9706,
    F9705, F9704, F9703, F9641, F9640, F9639, F9638, F9637, F9636, F9574,
    F9573, F9572, F9571, F9570, F9569, F9507, F9506, F9505, F9504, F9503,
    F9502, F9440, F9439, F9438, F9437, F9436, F9435, F9373, F9372, F9371,
    F9370, F9369, F9368, F9306, F9305, F9304, F9303, F9302, F9301, F9239,
    F9238, F9237, F9236, F9235, F9234, F9172, F9171, F9170, F9169, F9168,
    F9167, F9105, F9104, F9103, F9102, F9101, F9100, F9038, F9037, F9036,
    F9035, F9034, F9033, F8971, F8970, F8969, F8968, F8967, F8966, F8904,
    F8903, F8902, F8901, F8900, F8899, F8837, F8836, F8835, F8834, F8833,
    F8832, F8770, F8769, F8768, F8767, F8766, F8765, F8703, F8702, F8701,
    F8700, F8699, F8698, F8636, F8635, F8634, F8633, F8632, F8631, F8569,
    F8568, F8567, F8566, F8565, F8564, F8502, F8501, F8500, F8499, F8498,
    F8497, F8435, F8434, F8433, F8432, F8431, F8430, F8368, F8367, F8366,
    F8365, F8364, F8363, F8301, F8300, F8299, F8298, F8297, F8296, F8234,
    F8233, F8232, F8231, F8230, F8229, F8167, F8166, F8165, F8164, F8163,
    F8162, F8100, F8099, F8098, F8097, F8096, F8095, F8033, F8032, F8031,
    F8030, F8029, F8028, F7966, F7965, F7964, F7963, F7962, F7961, F7899,
    F7898, F7897, F7896, F7895, F7894, F7832, F7831, F7830, F7829, F7828,
    F7827, F7765, F7764, F7763, F7762, F7761, F7760, F7698, F7697, F7696,
    F7695, F7694, F7693, F7631, F7630, F7629, F7628, F7627, F7626, F7564,
    F7563, F7562, F7561, F7560, F7559, F7497, F7496, F7495, F7494, F7493,
    F7492, F7430, F7429, F7428, F7427, F7426, F7425, F7363, F7362, F7361,
    F7360, F7359, F7358, F7296, F7295, F7294, F7293, F7292, F7291, F7229,
    F7228, F7227, F7226, F7225, F7224, F7162, F7161, F7160, F7159, F7158,
    F7157, F7095, F7094, F7093, F7092, F7091, F7090, F7028, F7027, F7026,
    F7025, F7024, F7023, F6961, F6960, F6959, F6958, F6957, F6956, F6894,
    F6893, F6892, F6891, F6890, F6889, F6827, F6826, F6825, F6824, F6823,
    F6822, F6760, F6759, F6758, F6757, F6756, F6755, F6693, F6692, F6691,
    F6690, F6689, F6688, F6626, F6625, F6624, F6623, F6622, F6621, F6559,
    F6558, F6557, F6556, F6555, F6554, F6492, F6491, F6490, F6489, F6488,
    F6487, F6425, F6424, F6423, F6422, F6421, F6420, F6358, F6357, F6356,
    F6355, F6354, F6353, F6291, F6290, F6289, F6288, F6287, F6286, F6224,
    F6223, F6222, F6221, F6220, F6219, F6157, F6156, F6155, F6154, F6153,
    F6152, F6090, F6089, F6088, F6087, F6086, F6085, F6023, F6022, F6021,
    F6020, F6019, F6018, F5956, F5955, F5954, F5953, F5952, F5951, F5889,
    F5888, F5887, F5886, F5885, F5884, F5822, F5821, F5820, F5819, F5818,
    F5817, F5755, F5754, F5753, F5752, F5751, F5750, F5688, F5687, F5686,
    F5685, F5684, F5683, F5621, F5620, F5619, F5618, F5617, F5616, F5554,
    F5553, F5552, F5551, F5550, F5549, F5487, F5486, F5485, F5484, F5483,
    F5482, F5420, F5419, F5418, F5417, F5416, F5415, F5353, F5352, F5351,
    F5350, F5349, F5348, F5286, F5285, F5284, F5283, F5282, F5281, F5219,
    F5218, F5217, F5216, F5215, F5214, F5152, F5151, F5150, F5149, F5148,
    F5147, F5085, F5084, F5083, F5082, F5081, F5080, F5018, F5017, F5016,
    F5015, F5014, F5013, F4951, F4950, F4949, F4948, F4947, F4946, F4884,
    F4883, F4882, F4881, F4880, F4879, F4817, F4816, F4815, F4814, F4813,
    F4812, F4750, F4749, F4748, F4747, F4746, F4745, F4683, F4682, F4681,
    F4680, F4679, F4678, F4616, F4615, F4614, F4613, F4612, F4611, F4549,
    F4548, F4547, F4546, F4545, F4544, F4482, F4481, F4480, F4479, F4478,
    F4477, F4415, F4414, F4413, F4412, F4411, F4410, F4348, F4347, F4346,
    F4345, F4344, F4343, F4281, F4280, F4279, F4278, F4277, F4276, F4214,
    F4213, F4212, F4211, F4210, F4209, F4147, F4146, F4145, F4144, F4143,
    F4142, F4080, F4079, F4078, F4077, F4076, F4075, F4013, F4012, F4011,
    F4010, F4009, F4008, F3946, F3945, F3944, F3943, F3942, F3941, F3879,
    F3878, F3877, F3876, F3875, F3874, F3812, F3811, F3810, F3809, F3808,
    F3807, F3745, F3744, F3743, F3742, F3741, F3740, F3678, F3677, F3676,
    F3675, F3674, F3673, F3611, F3610, F3609, F3608, F3607, F3606, F3544,
    F3543, F3542, F3541, F3540, F3539, F3477, F3476, F3475, F3474, F3473,
    F3472, F3410, F3409, F3408, F3407, F3406, F3405, F3343, F3342, F3341,
    F3340, F3339, F3338, F3276, F3275, F3274, F3273, F3272, F3271, F3209,
    F3208, F3207, F3206, F3205, F3204, F3142, F3141, F3140, F3139, F3138,
    F3137, F3075, F3074, F3073, F3072, F3071, F3070, F3008, F3007, F3006,
    F3005, F3004, F3003, F2941, F2940, F2939, F2938, F2937, F2936, F2874,
    F2873, F2872, F2871, F2870, F2869, F2807, F2806, F2805, F2804, F2803,
    F2802, F2740, F2739, F2738, F2737, F2736, F2735, F2673, F2672, F2671,
    F2670, F2669, F2668, F2606, F2605, F2604, F2603, F2602, F2601, F2539,
    F2538, F2537, F2536, F2535, F2534, F2472, F2471, F2470, F2469, F2468,
    F2467, F2405, F2404, F2403, F2402, F2401, F2400, F2338, F2337, F2336,
    F2335, F2334, F2333, F2271, F2270, F2269, F2268, F2267, F2266, F2204,
    F2203, F2202, F2201, F2200, F2199, F2137, F2136, F2135, F2134, F2133,
    F2132, F2070, F2069, F2068, F2067, F2066, F2065, F2003, F2002, F2001,
    F2000, F1999, F1998, F1936, F1935, F1934, F1933, F1932, F1931, F1869,
    F1868, F1867, F1866, F1865, F1864, F1802, F1801, F1800, F1799, F1798,
    F1797, F1735, F1734, F1733, F1732, F1731, F1730, F1668, F1667, F1666,
    F1665, F1664, F1663, F1601, F1600, F1599, F1598, F1597, F1596, F1534,
    F1533, F1532, F1531, F1530, F1529, F1462, F1463, F1464, F1465, F1466,
    F1467,
    C2459, C2458, C2457, C2456, C2455, C2454, C2392, C2391, C2390, C2389,
    C2388, C2387, C2325, C2324, C2323, C2322, C2321, C2320, C2258, C2257,
    C2256, C2255, C2254, C2253, C2191, C2190, C2189, C2188, C2187, C2186,
    C2124, C2123, C2122, C2121, C2120, C2119, C2057, C2056, C2055, C2054,
    C2053, C2052, C1990, C1989, C1988, C1987, C1986, C1985, C1923, C1922,
    C1921, C1920, C1919, C1918, C1856, C1855, C1854, C1853, C1852, C1851,
    C1789, C1788, C1787, C1786, C1785, C1784, C1722, C1721, C1720, C1719,
    C1718, C1717, C1655, C1654, C1653, C1652, C1651, C1650, C1588, C1587,
    C1586, C1585, C1584, C1583, C1521, C1520, C1519, C1518, C1517, C1516,
    C1454, C1453, C1452, C1451, C1450, C1449, C1387, C1386, C1385, C1384,
    C1383, C1382, C1320, C1319, C1318, C1317, C1316, C1315, C1253, C1252,
    C1251, C1250, C1249, C1248, C1186, C1185, C1184, C1183, C1182, C1181,
    C1119, C1118, C1117, C1116, C1115, C1114, C1052, C1051, C1050, C1049,
    C1048, C1047, C985, C984, C983, C982, C981, C980, C918, C917, C916,
    C915, C914, C913, C851, C850, C849, C848, C847, C846, C784, C783, C782,
    C781, C780, C779, C717, C716, C715, C714, C713, C712, C650, C649, C648,
    C647, C646, C645, C583, C582, C581, C580, C579, C578, C516, C515, C514,
    C513, C512, C511, C449, C448, C447, C446, C445, C444, C382, C381, C380,
    C379, C378, C377, C315, C314, C313, C312, C311, C310, C248, C247, C246,
    C245, C244, C243, C181, C180, C179, C178, C177, C176, C114, C113, C112,
    C111, C110, C109, C47, C46, C45, C44, C43, C42, B9979, B9978, B9977,
    B9976, B9975, B9974, B9912, B9911, B9910, B9909, B9908, B9907, B9845,
    B9844, B9843, B9842, B9841, B9840, B9778, B9777, B9776, B9775, B9774,
    B9773, B9711, B9710, B9709, B9708, B9707, B9706, B9644, B9643, B9642,
    B9641, B9640, B9639, B9577, B9576, B9575, B9574, B9573, B9572, B9510,
    B9509, B9508, B9507, B9506, B9505, B9443, B9442, B9441, B9440, B9439,
    B9438, B9376, B9375, B9374, B9373, B9372, B9371, B9309, B9308, B9307,
    B9306, B9305, B9304, B9242, B9241, B9240, B9239, B9238, B9237, B9175,
    B9174, B9173, B9172, B9171, B9170, B9108, B9107, B9106, B9105, B9104,
    B9103, B9041, B9040, B9039, B9038, B9037, B9036, B8974, B8973, B8972,
    B8971, B8970, B8969, B8907, B8906, B8905, B8904, B8903, B8902, B8840,
    B8839, B8838, B8837, B8836, B8835, B8773, B8772, B8771, B8770, B8769,
    B8768, B8706, B8705, B8704, B8703, B8702, B8701, B8639, B8638, B8637,
    B8636, B8635, B8634, B8572, B8571, B8570, B8569, B8568, B8567, B8505,
    B8504, B8503, B8502, B8501, B8500, B8438, B8437, B8436, B8435, B8434,
    B8433, B8371, B8370, B8369, B8368, B8367, B8366, B8304, B8303, B8302,
    B8301, B8300, B8299, B8237, B8236, B8235, B8234, B8233, B8232, B8170,
    B8169, B8168, B8167, B8166, B8165, B8103, B8102, B8101, B8100, B8099,
    B8098, B8036, B8035, B8034, B8033, B8032, B8031, B7969, B7968, B7967,
    B7966, B7965, B7964, B7902, B7901, B7900, B7899, B7898, B7897, B7835,
    B7834, B7833, B7832, B7831, B7830, B7768, B7767, B7766, B7765, B7764,
    B7763, B7701, B7700, B7699, B7698, B7697, B7696, B7634, B7633, B7632,
    B7631, B7630, B7629, B7567, B7566, B7565, B7564, B7563, B7562, B7500,
    B7499, B7498, B7497, B7496, B7495, B7433, B7432, B7431, B7430, B7429,
    B7428, B7366, B7365, B7364, B7363, B7362, B7361, B7299, B7298, B7297,
    B7296, B7295, B7294, B7232, B7231, B7230, B7229, B7228, B7227, B7165,
    B7164, B7163, B7162, B7161, B7160, B7098, B7097, B7096, B7095, B7094,
    B7093, B7031, B7030, B7029, B7028, B7027, B7026, B6964, B6963, B6962,
    B6961, B6960, B6959, B6897, B6896, B6895, B6894, B6893, B6892, B6830,
    B6829, B6828, B6827, B6826, B6825, B6763, B6762, B6761, B6760, B6759,
    B6758, B6696, B6695, B6694, B6693, B6692, B6691, B6629, B6628, B6627,
    B6626, B6625, B6624, B6562, B6561, B6560, B6559, B6558, B6557, B6495,
    B6494, B6493, B6492, B6491, B6490, B6428, B6427, B6426, B6425, B6424,
    B6423, B6361, B6360, B6359, B6358, B6357, B6356, B6294, B6293, B6292,
    B6291, B6290, B6289, B6227, B6226, B6225, B6224, B6223, B6222, B6160,
    B6159, B6158, B6157, B6156, B6155, B6093, B6092, B6091, B6090, B6089,
    B6088, B6026, B6025, B6024, B6023, B6022, B6021, B5959, B5958, B5957,
    B5956, B5955, B5954, B5892, B5891, B5890, B5889, B5888, B5887, B5825,
    B5824, B5823, B5822, B5821, B5820, B5758, B5757, B5756, B5755, B5754,
    B5753, B5691, B5690, B5689, B5688, B5687, B5686, B5624, B5623, B5622,
    B5621, B5620, B5619, B5557, B5556, B5555, B5554, B5553, B5552, B5490,
    B5489, B5488, B5487, B5486, B5485, B5423, B5422, B5421, B5420, B5419,
    B5418, B5356, B5355, B5354, B5353, B5352, B5351, B5289, B5288, B5287,
    B5286, B5285, B5284, B5222, B5221, B5220, B5219, B5218, B5217, B5155,
    B5154, B5153, B5152, B5151, B5150, B5088, B5087, B5086, B5085, B5084,
    B5083, B5021, B5020, B5019, B5018, B5017, B5016, B4954, B4953, B4952,
    B4951, B4950, B4949, B4887, B4886, B4885, B4884, B4883, B4882, B4820,
    B4819, B4818, B4817, B4816, B4815, B4753, B4752, B4751, B4750, B4749,
    B4748, B4686, B4685, B4684, B4683, B4682, B4681, B4619, B4618, B4617,
    B4616, B4615, B4614, B4552, B4551, B4550, B4549, B4548, B4547, B4485,
    B4484, B4483, B4482, B4481, B4480, B4418, B4417, B4416, B4415, B4414,
    B4413, B4351, B4350, B4349, B4348, B4347, B4346, B4284, B4283, B4282,
    B4281, B4280, B4279, B4217, B4216, B4215, B4214, B4213, B4212, B4150,
    B4149, B4148, B4147, B4146, B4145, B4083, B4082, B4081, B4080, B4079,
    B4078, B4016, B4015, B4014, B4013, B4012, B4011, B3949, B3948, B3947,
    B3946, B3945, B3944, B3882, B3881, B3880, B3879, B3878, B3877, B3815,
    B3814, B3813, B3812, B3811, B3810, B3748, B3747, B3746, B3745, B3744,
    B3743, B3681, B3680, B3679, B3678, B3677, B3676, B3614, B3613, B3612,
    B3611, B3610, B3609, B3547, B3546, B3545, B3544, B3543, B3542, B3480,
    B3479, B3478, B3477, B3476, B3475, B3413, B3412, B3411, B3410, B3409,
    B3408, B3346, B3345, B3344, B3343, B3342, B3341, B3279, B3278, B3277,
    B3276, B3275, B3274, B3212, B3211, B3210, B3209, B3208, B3207, B3145,
    B3144, B3143, B3142, B3141, B3140, B3078, B3077, B3076, B3075, B3074,
    B3073, B3011, B3010, B3009, B3008, B3007, B3006, B2944, B2943, B2942,
    B2941, B2940, B2939, B2877, B2876, B2875, B2874, B2873, B2872, B2810,
    B2809, B2808, B2807, B2806, B2805, B2743, B2742, B2741, B2740, B2739,
    B2738, B2676, B2675, B2674, B2673, B2672, B2671, B2609, B2608, B2607,
    B2606, B2605, B2604, B2542, B2541, B2540, B2539, B2538, B2537, B2475,
    B2474, B2473, B2472, B2471, B2470, B2408, B2407, B2406, B2405, B2404,
    B2403, B2341, B2340, B2339, B2338, B2337, B2336, B2274, B2273, B2272,
    B2271, B2270, B2269, B2207, B2206, B2205, B2204, B2203, B2202, B2140,
    B2139, B2138, B2137, B2136, B2135, B2073, B2072, B2071, B2070, B2069,
    B2068, B2006, B2005, B2004, B2003, B2002, B2001, B1939, B1938, B1937,
    B1936, B1935, B1934, B1872, B1871, B1870, B1869, B1868, B1867, B1805,
    B1804, B1803, B1802, B1801, B1800, B1738, B1737, B1736, B1735, B1734,
    B1733, B1671, B1670, B1669, B1668, B1667, B1666, B1604, B1603, B1602,
    B1601, B1600, B1599, B1537, B1536, B1535, B1534, B1533, B1532, B1470,
    B1469, B1468, B1467, B1466, B1465, B1403, B1402, B1401, B1400, B1399,
    B1398, B1336, B1335, B1334, B1333, B1332, B1331, B1269, B1268, B1267,
    B1266, B1265, B1264, B1202, B1201, B1200, B1199, B1198, B1197, B1135,
    B1134, B1133, B1132, B1131, B1130, B1068, B1067, B1066, B1065, B1064,
    B1063, B1001, B1000, B999, B998, B997, B996, B934, B933, B932, B931,
    B930, B929, B867, B866, B865, B864, B863, B862, B800, B799, B798, B797,
    B796, B795, B733, B732, B731, B730, B729, B728, B666, B665, B664, B663,
    B662, B661, B599, B598, B597, B596, B595, B594, B532, B531, B530, B529,
    B528, B527, B465, B464, B463, B462, B461, B460, B398, B397, B396, B395,
    B394, B393, B331, B330, B329, B328, B327, B326, B264, B263, B262, B261,
    B260, B259, B197, B196, B195, B194, B193, B192, B130, B129, B128, B127,
    B126, B125, B63, B62, B61, B60, B59, B58, A9995, A9994, A9993, A9992,
    A9991, A9990, A9928, A9927, A9926, A9925, A9924, A9923, A9861, A9860,
    A9859, A9858, A9857, A9856, A9794, A9793, A9792, A9791, A9790, A9789,
    A9727, A9726, A9725, A9724, A9723, A9722, A9660, A9659, A9658, A9657,
    A9656, A9655, A9593, A9592, A9591, A9590, A9589, A9588, A9526, A9525,
    A9524, A9523, A9522, A9521, A9459, A9458, A9457, A9456, A9455, A9454,
    A9392, A9391, A9390, A9389, A9388, A9387, A9325, A9324, A9323, A9322,
    A9321, A9320, A9258, A9257, A9256, A9255, A9254, A9253, A9191, A9190,
    A9189, A9188, A9187, A9186, A9124, A9123, A9122, A9121, A9120, A9119,
    A9057, A9056, A9055, A9054, A9053, A9052, A8990, A8989, A8988, A8987,
    A8986, A8985, A8923, A8922, A8921, A8920, A8919, A8918, A8856, A8855,
    A8854, A8853, A8852, A8851, A8789, A8788, A8787, A8786, A8785, A8784,
    A8722, A8721, A8720, A8719, A8718, A8717, A8655, A8654, A8653, A8652,
    A8651, A8650, A8588, A8587, A8586, A8585, A8584, A8583, A8521, A8520,
    A8519, A8518, A8517, A8516, A8454, A8453, A8452, A8451, A8450, A8449,
    A8387, A8386, A8385, A8384, A8383, A8382, A8320, A8319, A8318, A8317,
    A8316, A8315, A8253, A8252, A8251, A8250, A8249, A8248, A8186, A8185,
    A8184, A8183, A8182, A8181, A8119, A8118, A8117, A8116, A8115, A8114,
    A8047, A8048, A8049, A8050, A8051, A8052  );
  input  G5873, G5872, G5871, G5870, G5869, G5868, G5806, G5805, G5804,
    G5803, G5802, G5801, G5739, G5738, G5737, G5736, G5735, G5734, G5672,
    G5671, G5670, G5669, G5668, G5667, G5605, G5604, G5603, G5602, G5601,
    G5600, G5538, G5537, G5536, G5535, G5534, G5533, G5471, G5470, G5469,
    G5468, G5467, G5466, G5404, G5403, G5402, G5401, G5400, G5399, G5337,
    G5336, G5335, G5334, G5333, G5332, G5270, G5269, G5268, G5267, G5266,
    G5265, G5203, G5202, G5201, G5200, G5199, G5198, G5136, G5135, G5134,
    G5133, G5132, G5131, G5069, G5068, G5067, G5066, G5065, G5064, G5002,
    G5001, G5000, G4999, G4998, G4997, G4935, G4934, G4933, G4932, G4931,
    G4930, G4868, G4867, G4866, G4865, G4864, G4863, G4801, G4800, G4799,
    G4798, G4797, G4796, G4734, G4733, G4732, G4731, G4730, G4729, G4667,
    G4666, G4665, G4664, G4663, G4662, G4600, G4599, G4598, G4597, G4596,
    G4595, G4533, G4532, G4531, G4530, G4529, G4528, G4466, G4465, G4464,
    G4463, G4462, G4461, G4399, G4398, G4397, G4396, G4395, G4394, G4332,
    G4331, G4330, G4329, G4328, G4327, G4265, G4264, G4263, G4262, G4261,
    G4260, G4198, G4197, G4196, G4195, G4194, G4193, G4131, G4130, G4129,
    G4128, G4127, G4126, G4064, G4063, G4062, G4061, G4060, G4059, G3997,
    G3996, G3995, G3994, G3993, G3992, G3930, G3929, G3928, G3927, G3926,
    G3925, G3863, G3862, G3861, G3860, G3859, G3858, G3796, G3795, G3794,
    G3793, G3792, G3791, G3729, G3728, G3727, G3726, G3725, G3724, G3662,
    G3661, G3660, G3659, G3658, G3657, G3595, G3594, G3593, G3592, G3591,
    G3590, G3528, G3527, G3526, G3525, G3524, G3523, G3461, G3460, G3459,
    G3458, G3457, G3456, G3394, G3393, G3392, G3391, G3390, G3389, G3327,
    G3326, G3325, G3324, G3323, G3322, G3260, G3259, G3258, G3257, G3256,
    G3255, G3193, G3192, G3191, G3190, G3189, G3188, G3126, G3125, G3124,
    G3123, G3122, G3121, G3059, G3058, G3057, G3056, G3055, G3054, G2992,
    G2991, G2990, G2989, G2988, G2987, G2925, G2924, G2923, G2922, G2921,
    G2920, G2858, G2857, G2856, G2855, G2854, G2853, G2791, G2790, G2789,
    G2788, G2787, G2786, G2724, G2723, G2722, G2721, G2720, G2719, G2657,
    G2656, G2655, G2654, G2653, G2652, G2590, G2589, G2588, G2587, G2586,
    G2585, G2523, G2522, G2521, G2520, G2519, G2518, G2456, G2455, G2454,
    G2453, G2452, G2451, G2389, G2388, G2387, G2386, G2385, G2384, G2322,
    G2321, G2320, G2319, G2318, G2317, G2255, G2254, G2253, G2252, G2251,
    G2250, G2188, G2187, G2186, G2185, G2184, G2183, G2121, G2120, G2119,
    G2118, G2117, G2116, G2054, G2053, G2052, G2051, G2050, G2049, G1987,
    G1986, G1985, G1984, G1983, G1982, G1920, G1919, G1918, G1917, G1916,
    G1915, G1853, G1852, G1851, G1850, G1849, G1848, G1786, G1785, G1784,
    G1783, G1782, G1781, G1719, G1718, G1717, G1716, G1715, G1714, G1652,
    G1651, G1650, G1649, G1648, G1647, G1585, G1584, G1583, G1582, G1581,
    G1580, G1518, G1517, G1516, G1515, G1514, G1513, G1451, G1450, G1449,
    G1448, G1447, G1446, G1384, G1383, G1382, G1381, G1380, G1379, G1317,
    G1316, G1315, G1314, G1313, G1312, G1250, G1249, G1248, G1247, G1246,
    G1245, G1183, G1182, G1181, G1180, G1179, G1178, G1116, G1115, G1114,
    G1113, G1112, G1111, G1049, G1048, G1047, G1046, G1045, G1044, G982,
    G981, G980, G979, G978, G977, G915, G914, G913, G912, G911, G910, G848,
    G847, G846, G845, G844, G843, G781, G780, G779, G778, G777, G776, G714,
    G713, G712, G711, G710, G709, G647, G646, G645, G644, G643, G642, G580,
    G579, G578, G577, G576, G575, G513, G512, G511, G510, G509, G508, G446,
    G445, G444, G443, G442, G441, G379, G378, G377, G376, G375, G374, G312,
    G311, G310, G309, G308, G307, G245, G244, G243, G242, G241, G240, G178,
    G177, G176, G175, G174, G173, G111, G110, G109, G108, G107, G106, G44,
    G43, G42, G41, G40, G39, F9976, F9975, F9974, F9973, F9972, F9971,
    F9909, F9908, F9907, F9906, F9905, F9904, F9842, F9841, F9840, F9839,
    F9838, F9837, F9775, F9774, F9773, F9772, F9771, F9770, F9708, F9707,
    F9706, F9705, F9704, F9703, F9641, F9640, F9639, F9638, F9637, F9636,
    F9574, F9573, F9572, F9571, F9570, F9569, F9507, F9506, F9505, F9504,
    F9503, F9502, F9440, F9439, F9438, F9437, F9436, F9435, F9373, F9372,
    F9371, F9370, F9369, F9368, F9306, F9305, F9304, F9303, F9302, F9301,
    F9239, F9238, F9237, F9236, F9235, F9234, F9172, F9171, F9170, F9169,
    F9168, F9167, F9105, F9104, F9103, F9102, F9101, F9100, F9038, F9037,
    F9036, F9035, F9034, F9033, F8971, F8970, F8969, F8968, F8967, F8966,
    F8904, F8903, F8902, F8901, F8900, F8899, F8837, F8836, F8835, F8834,
    F8833, F8832, F8770, F8769, F8768, F8767, F8766, F8765, F8703, F8702,
    F8701, F8700, F8699, F8698, F8636, F8635, F8634, F8633, F8632, F8631,
    F8569, F8568, F8567, F8566, F8565, F8564, F8502, F8501, F8500, F8499,
    F8498, F8497, F8435, F8434, F8433, F8432, F8431, F8430, F8368, F8367,
    F8366, F8365, F8364, F8363, F8301, F8300, F8299, F8298, F8297, F8296,
    F8234, F8233, F8232, F8231, F8230, F8229, F8167, F8166, F8165, F8164,
    F8163, F8162, F8100, F8099, F8098, F8097, F8096, F8095, F8033, F8032,
    F8031, F8030, F8029, F8028, F7966, F7965, F7964, F7963, F7962, F7961,
    F7899, F7898, F7897, F7896, F7895, F7894, F7832, F7831, F7830, F7829,
    F7828, F7827, F7765, F7764, F7763, F7762, F7761, F7760, F7698, F7697,
    F7696, F7695, F7694, F7693, F7631, F7630, F7629, F7628, F7627, F7626,
    F7564, F7563, F7562, F7561, F7560, F7559, F7497, F7496, F7495, F7494,
    F7493, F7492, F7430, F7429, F7428, F7427, F7426, F7425, F7363, F7362,
    F7361, F7360, F7359, F7358, F7296, F7295, F7294, F7293, F7292, F7291,
    F7229, F7228, F7227, F7226, F7225, F7224, F7162, F7161, F7160, F7159,
    F7158, F7157, F7095, F7094, F7093, F7092, F7091, F7090, F7028, F7027,
    F7026, F7025, F7024, F7023, F6961, F6960, F6959, F6958, F6957, F6956,
    F6894, F6893, F6892, F6891, F6890, F6889, F6827, F6826, F6825, F6824,
    F6823, F6822, F6760, F6759, F6758, F6757, F6756, F6755, F6693, F6692,
    F6691, F6690, F6689, F6688, F6626, F6625, F6624, F6623, F6622, F6621,
    F6559, F6558, F6557, F6556, F6555, F6554, F6492, F6491, F6490, F6489,
    F6488, F6487, F6425, F6424, F6423, F6422, F6421, F6420, F6358, F6357,
    F6356, F6355, F6354, F6353, F6291, F6290, F6289, F6288, F6287, F6286,
    F6224, F6223, F6222, F6221, F6220, F6219, F6157, F6156, F6155, F6154,
    F6153, F6152, F6090, F6089, F6088, F6087, F6086, F6085, F6023, F6022,
    F6021, F6020, F6019, F6018, F5956, F5955, F5954, F5953, F5952, F5951,
    F5889, F5888, F5887, F5886, F5885, F5884, F5822, F5821, F5820, F5819,
    F5818, F5817, F5755, F5754, F5753, F5752, F5751, F5750, F5688, F5687,
    F5686, F5685, F5684, F5683, F5621, F5620, F5619, F5618, F5617, F5616,
    F5554, F5553, F5552, F5551, F5550, F5549, F5487, F5486, F5485, F5484,
    F5483, F5482, F5420, F5419, F5418, F5417, F5416, F5415, F5353, F5352,
    F5351, F5350, F5349, F5348, F5286, F5285, F5284, F5283, F5282, F5281,
    F5219, F5218, F5217, F5216, F5215, F5214, F5152, F5151, F5150, F5149,
    F5148, F5147, F5085, F5084, F5083, F5082, F5081, F5080, F5018, F5017,
    F5016, F5015, F5014, F5013, F4951, F4950, F4949, F4948, F4947, F4946,
    F4884, F4883, F4882, F4881, F4880, F4879, F4817, F4816, F4815, F4814,
    F4813, F4812, F4750, F4749, F4748, F4747, F4746, F4745, F4683, F4682,
    F4681, F4680, F4679, F4678, F4616, F4615, F4614, F4613, F4612, F4611,
    F4549, F4548, F4547, F4546, F4545, F4544, F4482, F4481, F4480, F4479,
    F4478, F4477, F4415, F4414, F4413, F4412, F4411, F4410, F4348, F4347,
    F4346, F4345, F4344, F4343, F4281, F4280, F4279, F4278, F4277, F4276,
    F4214, F4213, F4212, F4211, F4210, F4209, F4147, F4146, F4145, F4144,
    F4143, F4142, F4080, F4079, F4078, F4077, F4076, F4075, F4013, F4012,
    F4011, F4010, F4009, F4008, F3946, F3945, F3944, F3943, F3942, F3941,
    F3879, F3878, F3877, F3876, F3875, F3874, F3812, F3811, F3810, F3809,
    F3808, F3807, F3745, F3744, F3743, F3742, F3741, F3740, F3678, F3677,
    F3676, F3675, F3674, F3673, F3611, F3610, F3609, F3608, F3607, F3606,
    F3544, F3543, F3542, F3541, F3540, F3539, F3477, F3476, F3475, F3474,
    F3473, F3472, F3410, F3409, F3408, F3407, F3406, F3405, F3343, F3342,
    F3341, F3340, F3339, F3338, F3276, F3275, F3274, F3273, F3272, F3271,
    F3209, F3208, F3207, F3206, F3205, F3204, F3142, F3141, F3140, F3139,
    F3138, F3137, F3075, F3074, F3073, F3072, F3071, F3070, F3008, F3007,
    F3006, F3005, F3004, F3003, F2941, F2940, F2939, F2938, F2937, F2936,
    F2874, F2873, F2872, F2871, F2870, F2869, F2807, F2806, F2805, F2804,
    F2803, F2802, F2740, F2739, F2738, F2737, F2736, F2735, F2673, F2672,
    F2671, F2670, F2669, F2668, F2606, F2605, F2604, F2603, F2602, F2601,
    F2539, F2538, F2537, F2536, F2535, F2534, F2472, F2471, F2470, F2469,
    F2468, F2467, F2405, F2404, F2403, F2402, F2401, F2400, F2338, F2337,
    F2336, F2335, F2334, F2333, F2271, F2270, F2269, F2268, F2267, F2266,
    F2204, F2203, F2202, F2201, F2200, F2199, F2137, F2136, F2135, F2134,
    F2133, F2132, F2070, F2069, F2068, F2067, F2066, F2065, F2003, F2002,
    F2001, F2000, F1999, F1998, F1936, F1935, F1934, F1933, F1932, F1931,
    F1869, F1868, F1867, F1866, F1865, F1864, F1802, F1801, F1800, F1799,
    F1798, F1797, F1735, F1734, F1733, F1732, F1731, F1730, F1668, F1667,
    F1666, F1665, F1664, F1663, F1601, F1600, F1599, F1598, F1597, F1596,
    F1534, F1533, F1532, F1531, F1530, F1529, F1462, F1463, F1464, F1465,
    F1466, F1467;
  output C2459, C2458, C2457, C2456, C2455, C2454, C2392, C2391, C2390, C2389,
    C2388, C2387, C2325, C2324, C2323, C2322, C2321, C2320, C2258, C2257,
    C2256, C2255, C2254, C2253, C2191, C2190, C2189, C2188, C2187, C2186,
    C2124, C2123, C2122, C2121, C2120, C2119, C2057, C2056, C2055, C2054,
    C2053, C2052, C1990, C1989, C1988, C1987, C1986, C1985, C1923, C1922,
    C1921, C1920, C1919, C1918, C1856, C1855, C1854, C1853, C1852, C1851,
    C1789, C1788, C1787, C1786, C1785, C1784, C1722, C1721, C1720, C1719,
    C1718, C1717, C1655, C1654, C1653, C1652, C1651, C1650, C1588, C1587,
    C1586, C1585, C1584, C1583, C1521, C1520, C1519, C1518, C1517, C1516,
    C1454, C1453, C1452, C1451, C1450, C1449, C1387, C1386, C1385, C1384,
    C1383, C1382, C1320, C1319, C1318, C1317, C1316, C1315, C1253, C1252,
    C1251, C1250, C1249, C1248, C1186, C1185, C1184, C1183, C1182, C1181,
    C1119, C1118, C1117, C1116, C1115, C1114, C1052, C1051, C1050, C1049,
    C1048, C1047, C985, C984, C983, C982, C981, C980, C918, C917, C916,
    C915, C914, C913, C851, C850, C849, C848, C847, C846, C784, C783, C782,
    C781, C780, C779, C717, C716, C715, C714, C713, C712, C650, C649, C648,
    C647, C646, C645, C583, C582, C581, C580, C579, C578, C516, C515, C514,
    C513, C512, C511, C449, C448, C447, C446, C445, C444, C382, C381, C380,
    C379, C378, C377, C315, C314, C313, C312, C311, C310, C248, C247, C246,
    C245, C244, C243, C181, C180, C179, C178, C177, C176, C114, C113, C112,
    C111, C110, C109, C47, C46, C45, C44, C43, C42, B9979, B9978, B9977,
    B9976, B9975, B9974, B9912, B9911, B9910, B9909, B9908, B9907, B9845,
    B9844, B9843, B9842, B9841, B9840, B9778, B9777, B9776, B9775, B9774,
    B9773, B9711, B9710, B9709, B9708, B9707, B9706, B9644, B9643, B9642,
    B9641, B9640, B9639, B9577, B9576, B9575, B9574, B9573, B9572, B9510,
    B9509, B9508, B9507, B9506, B9505, B9443, B9442, B9441, B9440, B9439,
    B9438, B9376, B9375, B9374, B9373, B9372, B9371, B9309, B9308, B9307,
    B9306, B9305, B9304, B9242, B9241, B9240, B9239, B9238, B9237, B9175,
    B9174, B9173, B9172, B9171, B9170, B9108, B9107, B9106, B9105, B9104,
    B9103, B9041, B9040, B9039, B9038, B9037, B9036, B8974, B8973, B8972,
    B8971, B8970, B8969, B8907, B8906, B8905, B8904, B8903, B8902, B8840,
    B8839, B8838, B8837, B8836, B8835, B8773, B8772, B8771, B8770, B8769,
    B8768, B8706, B8705, B8704, B8703, B8702, B8701, B8639, B8638, B8637,
    B8636, B8635, B8634, B8572, B8571, B8570, B8569, B8568, B8567, B8505,
    B8504, B8503, B8502, B8501, B8500, B8438, B8437, B8436, B8435, B8434,
    B8433, B8371, B8370, B8369, B8368, B8367, B8366, B8304, B8303, B8302,
    B8301, B8300, B8299, B8237, B8236, B8235, B8234, B8233, B8232, B8170,
    B8169, B8168, B8167, B8166, B8165, B8103, B8102, B8101, B8100, B8099,
    B8098, B8036, B8035, B8034, B8033, B8032, B8031, B7969, B7968, B7967,
    B7966, B7965, B7964, B7902, B7901, B7900, B7899, B7898, B7897, B7835,
    B7834, B7833, B7832, B7831, B7830, B7768, B7767, B7766, B7765, B7764,
    B7763, B7701, B7700, B7699, B7698, B7697, B7696, B7634, B7633, B7632,
    B7631, B7630, B7629, B7567, B7566, B7565, B7564, B7563, B7562, B7500,
    B7499, B7498, B7497, B7496, B7495, B7433, B7432, B7431, B7430, B7429,
    B7428, B7366, B7365, B7364, B7363, B7362, B7361, B7299, B7298, B7297,
    B7296, B7295, B7294, B7232, B7231, B7230, B7229, B7228, B7227, B7165,
    B7164, B7163, B7162, B7161, B7160, B7098, B7097, B7096, B7095, B7094,
    B7093, B7031, B7030, B7029, B7028, B7027, B7026, B6964, B6963, B6962,
    B6961, B6960, B6959, B6897, B6896, B6895, B6894, B6893, B6892, B6830,
    B6829, B6828, B6827, B6826, B6825, B6763, B6762, B6761, B6760, B6759,
    B6758, B6696, B6695, B6694, B6693, B6692, B6691, B6629, B6628, B6627,
    B6626, B6625, B6624, B6562, B6561, B6560, B6559, B6558, B6557, B6495,
    B6494, B6493, B6492, B6491, B6490, B6428, B6427, B6426, B6425, B6424,
    B6423, B6361, B6360, B6359, B6358, B6357, B6356, B6294, B6293, B6292,
    B6291, B6290, B6289, B6227, B6226, B6225, B6224, B6223, B6222, B6160,
    B6159, B6158, B6157, B6156, B6155, B6093, B6092, B6091, B6090, B6089,
    B6088, B6026, B6025, B6024, B6023, B6022, B6021, B5959, B5958, B5957,
    B5956, B5955, B5954, B5892, B5891, B5890, B5889, B5888, B5887, B5825,
    B5824, B5823, B5822, B5821, B5820, B5758, B5757, B5756, B5755, B5754,
    B5753, B5691, B5690, B5689, B5688, B5687, B5686, B5624, B5623, B5622,
    B5621, B5620, B5619, B5557, B5556, B5555, B5554, B5553, B5552, B5490,
    B5489, B5488, B5487, B5486, B5485, B5423, B5422, B5421, B5420, B5419,
    B5418, B5356, B5355, B5354, B5353, B5352, B5351, B5289, B5288, B5287,
    B5286, B5285, B5284, B5222, B5221, B5220, B5219, B5218, B5217, B5155,
    B5154, B5153, B5152, B5151, B5150, B5088, B5087, B5086, B5085, B5084,
    B5083, B5021, B5020, B5019, B5018, B5017, B5016, B4954, B4953, B4952,
    B4951, B4950, B4949, B4887, B4886, B4885, B4884, B4883, B4882, B4820,
    B4819, B4818, B4817, B4816, B4815, B4753, B4752, B4751, B4750, B4749,
    B4748, B4686, B4685, B4684, B4683, B4682, B4681, B4619, B4618, B4617,
    B4616, B4615, B4614, B4552, B4551, B4550, B4549, B4548, B4547, B4485,
    B4484, B4483, B4482, B4481, B4480, B4418, B4417, B4416, B4415, B4414,
    B4413, B4351, B4350, B4349, B4348, B4347, B4346, B4284, B4283, B4282,
    B4281, B4280, B4279, B4217, B4216, B4215, B4214, B4213, B4212, B4150,
    B4149, B4148, B4147, B4146, B4145, B4083, B4082, B4081, B4080, B4079,
    B4078, B4016, B4015, B4014, B4013, B4012, B4011, B3949, B3948, B3947,
    B3946, B3945, B3944, B3882, B3881, B3880, B3879, B3878, B3877, B3815,
    B3814, B3813, B3812, B3811, B3810, B3748, B3747, B3746, B3745, B3744,
    B3743, B3681, B3680, B3679, B3678, B3677, B3676, B3614, B3613, B3612,
    B3611, B3610, B3609, B3547, B3546, B3545, B3544, B3543, B3542, B3480,
    B3479, B3478, B3477, B3476, B3475, B3413, B3412, B3411, B3410, B3409,
    B3408, B3346, B3345, B3344, B3343, B3342, B3341, B3279, B3278, B3277,
    B3276, B3275, B3274, B3212, B3211, B3210, B3209, B3208, B3207, B3145,
    B3144, B3143, B3142, B3141, B3140, B3078, B3077, B3076, B3075, B3074,
    B3073, B3011, B3010, B3009, B3008, B3007, B3006, B2944, B2943, B2942,
    B2941, B2940, B2939, B2877, B2876, B2875, B2874, B2873, B2872, B2810,
    B2809, B2808, B2807, B2806, B2805, B2743, B2742, B2741, B2740, B2739,
    B2738, B2676, B2675, B2674, B2673, B2672, B2671, B2609, B2608, B2607,
    B2606, B2605, B2604, B2542, B2541, B2540, B2539, B2538, B2537, B2475,
    B2474, B2473, B2472, B2471, B2470, B2408, B2407, B2406, B2405, B2404,
    B2403, B2341, B2340, B2339, B2338, B2337, B2336, B2274, B2273, B2272,
    B2271, B2270, B2269, B2207, B2206, B2205, B2204, B2203, B2202, B2140,
    B2139, B2138, B2137, B2136, B2135, B2073, B2072, B2071, B2070, B2069,
    B2068, B2006, B2005, B2004, B2003, B2002, B2001, B1939, B1938, B1937,
    B1936, B1935, B1934, B1872, B1871, B1870, B1869, B1868, B1867, B1805,
    B1804, B1803, B1802, B1801, B1800, B1738, B1737, B1736, B1735, B1734,
    B1733, B1671, B1670, B1669, B1668, B1667, B1666, B1604, B1603, B1602,
    B1601, B1600, B1599, B1537, B1536, B1535, B1534, B1533, B1532, B1470,
    B1469, B1468, B1467, B1466, B1465, B1403, B1402, B1401, B1400, B1399,
    B1398, B1336, B1335, B1334, B1333, B1332, B1331, B1269, B1268, B1267,
    B1266, B1265, B1264, B1202, B1201, B1200, B1199, B1198, B1197, B1135,
    B1134, B1133, B1132, B1131, B1130, B1068, B1067, B1066, B1065, B1064,
    B1063, B1001, B1000, B999, B998, B997, B996, B934, B933, B932, B931,
    B930, B929, B867, B866, B865, B864, B863, B862, B800, B799, B798, B797,
    B796, B795, B733, B732, B731, B730, B729, B728, B666, B665, B664, B663,
    B662, B661, B599, B598, B597, B596, B595, B594, B532, B531, B530, B529,
    B528, B527, B465, B464, B463, B462, B461, B460, B398, B397, B396, B395,
    B394, B393, B331, B330, B329, B328, B327, B326, B264, B263, B262, B261,
    B260, B259, B197, B196, B195, B194, B193, B192, B130, B129, B128, B127,
    B126, B125, B63, B62, B61, B60, B59, B58, A9995, A9994, A9993, A9992,
    A9991, A9990, A9928, A9927, A9926, A9925, A9924, A9923, A9861, A9860,
    A9859, A9858, A9857, A9856, A9794, A9793, A9792, A9791, A9790, A9789,
    A9727, A9726, A9725, A9724, A9723, A9722, A9660, A9659, A9658, A9657,
    A9656, A9655, A9593, A9592, A9591, A9590, A9589, A9588, A9526, A9525,
    A9524, A9523, A9522, A9521, A9459, A9458, A9457, A9456, A9455, A9454,
    A9392, A9391, A9390, A9389, A9388, A9387, A9325, A9324, A9323, A9322,
    A9321, A9320, A9258, A9257, A9256, A9255, A9254, A9253, A9191, A9190,
    A9189, A9188, A9187, A9186, A9124, A9123, A9122, A9121, A9120, A9119,
    A9057, A9056, A9055, A9054, A9053, A9052, A8990, A8989, A8988, A8987,
    A8986, A8985, A8923, A8922, A8921, A8920, A8919, A8918, A8856, A8855,
    A8854, A8853, A8852, A8851, A8789, A8788, A8787, A8786, A8785, A8784,
    A8722, A8721, A8720, A8719, A8718, A8717, A8655, A8654, A8653, A8652,
    A8651, A8650, A8588, A8587, A8586, A8585, A8584, A8583, A8521, A8520,
    A8519, A8518, A8517, A8516, A8454, A8453, A8452, A8451, A8450, A8449,
    A8387, A8386, A8385, A8384, A8383, A8382, A8320, A8319, A8318, A8317,
    A8316, A8315, A8253, A8252, A8251, A8250, A8249, A8248, A8186, A8185,
    A8184, A8183, A8182, A8181, A8119, A8118, A8117, A8116, A8115, A8114,
    A8047, A8048, A8049, A8050, A8051, A8052;
  wire new_F1528_, new_F1527_, new_F1526_, new_F1525_, new_F1524_,
    new_F1523_, new_F1522_, new_F1521_, new_F1520_, new_F1519_, new_F1518_,
    new_F1517_, new_F1516_, new_F1515_, new_F1514_, new_F1513_, new_F1512_,
    new_F1511_, new_F1510_, new_F1509_, new_F1508_, new_F1507_, new_F1506_,
    new_F1505_, new_F1504_, new_F1503_, new_F1502_, new_F1501_, new_F1500_,
    new_F1499_, new_F1498_, new_F1497_, new_F1496_, new_F1495_, new_F1494_,
    new_F1493_, new_F1492_, new_F1491_, new_F1490_, new_F1489_, new_F1488_,
    new_F1487_, new_F1486_, new_F1485_, new_F1484_, new_F1483_, new_F1482_,
    new_F1481_, new_F1480_, new_F1479_, new_F1478_, new_F1477_, new_F1476_,
    new_F1475_, new_F1474_, new_F1473_, new_F1472_, new_F1471_, new_F1470_,
    new_F1469_, new_F1468_, new_F1535_, new_F1536_, new_F1537_, new_F1538_,
    new_F1539_, new_F1540_, new_F1541_, new_F1542_, new_F1543_, new_F1544_,
    new_F1545_, new_F1546_, new_F1547_, new_F1548_, new_F1549_, new_F1550_,
    new_F1551_, new_F1552_, new_F1553_, new_F1554_, new_F1555_, new_F1556_,
    new_F1557_, new_F1558_, new_F1559_, new_F1560_, new_F1561_, new_F1562_,
    new_F1563_, new_F1564_, new_F1565_, new_F1566_, new_F1567_, new_F1568_,
    new_F1569_, new_F1570_, new_F1571_, new_F1572_, new_F1573_, new_F1574_,
    new_F1575_, new_F1576_, new_F1577_, new_F1578_, new_F1579_, new_F1580_,
    new_F1581_, new_F1582_, new_F1583_, new_F1584_, new_F1585_, new_F1586_,
    new_F1587_, new_F1588_, new_F1589_, new_F1590_, new_F1591_, new_F1592_,
    new_F1593_, new_F1594_, new_F1595_, new_F1602_, new_F1603_, new_F1604_,
    new_F1605_, new_F1606_, new_F1607_, new_F1608_, new_F1609_, new_F1610_,
    new_F1611_, new_F1612_, new_F1613_, new_F1614_, new_F1615_, new_F1616_,
    new_F1617_, new_F1618_, new_F1619_, new_F1620_, new_F1621_, new_F1622_,
    new_F1623_, new_F1624_, new_F1625_, new_F1626_, new_F1627_, new_F1628_,
    new_F1629_, new_F1630_, new_F1631_, new_F1632_, new_F1633_, new_F1634_,
    new_F1635_, new_F1636_, new_F1637_, new_F1638_, new_F1639_, new_F1640_,
    new_F1641_, new_F1642_, new_F1643_, new_F1644_, new_F1645_, new_F1646_,
    new_F1647_, new_F1648_, new_F1649_, new_F1650_, new_F1651_, new_F1652_,
    new_F1653_, new_F1654_, new_F1655_, new_F1656_, new_F1657_, new_F1658_,
    new_F1659_, new_F1660_, new_F1661_, new_F1662_, new_F1669_, new_F1670_,
    new_F1671_, new_F1672_, new_F1673_, new_F1674_, new_F1675_, new_F1676_,
    new_F1677_, new_F1678_, new_F1679_, new_F1680_, new_F1681_, new_F1682_,
    new_F1683_, new_F1684_, new_F1685_, new_F1686_, new_F1687_, new_F1688_,
    new_F1689_, new_F1690_, new_F1691_, new_F1692_, new_F1693_, new_F1694_,
    new_F1695_, new_F1696_, new_F1697_, new_F1698_, new_F1699_, new_F1700_,
    new_F1701_, new_F1702_, new_F1703_, new_F1704_, new_F1705_, new_F1706_,
    new_F1707_, new_F1708_, new_F1709_, new_F1710_, new_F1711_, new_F1712_,
    new_F1713_, new_F1714_, new_F1715_, new_F1716_, new_F1717_, new_F1718_,
    new_F1719_, new_F1720_, new_F1721_, new_F1722_, new_F1723_, new_F1724_,
    new_F1725_, new_F1726_, new_F1727_, new_F1728_, new_F1729_, new_F1736_,
    new_F1737_, new_F1738_, new_F1739_, new_F1740_, new_F1741_, new_F1742_,
    new_F1743_, new_F1744_, new_F1745_, new_F1746_, new_F1747_, new_F1748_,
    new_F1749_, new_F1750_, new_F1751_, new_F1752_, new_F1753_, new_F1754_,
    new_F1755_, new_F1756_, new_F1757_, new_F1758_, new_F1759_, new_F1760_,
    new_F1761_, new_F1762_, new_F1763_, new_F1764_, new_F1765_, new_F1766_,
    new_F1767_, new_F1768_, new_F1769_, new_F1770_, new_F1771_, new_F1772_,
    new_F1773_, new_F1774_, new_F1775_, new_F1776_, new_F1777_, new_F1778_,
    new_F1779_, new_F1780_, new_F1781_, new_F1782_, new_F1783_, new_F1784_,
    new_F1785_, new_F1786_, new_F1787_, new_F1788_, new_F1789_, new_F1790_,
    new_F1791_, new_F1792_, new_F1793_, new_F1794_, new_F1795_, new_F1796_,
    new_F1803_, new_F1804_, new_F1805_, new_F1806_, new_F1807_, new_F1808_,
    new_F1809_, new_F1810_, new_F1811_, new_F1812_, new_F1813_, new_F1814_,
    new_F1815_, new_F1816_, new_F1817_, new_F1818_, new_F1819_, new_F1820_,
    new_F1821_, new_F1822_, new_F1823_, new_F1824_, new_F1825_, new_F1826_,
    new_F1827_, new_F1828_, new_F1829_, new_F1830_, new_F1831_, new_F1832_,
    new_F1833_, new_F1834_, new_F1835_, new_F1836_, new_F1837_, new_F1838_,
    new_F1839_, new_F1840_, new_F1841_, new_F1842_, new_F1843_, new_F1844_,
    new_F1845_, new_F1846_, new_F1847_, new_F1848_, new_F1849_, new_F1850_,
    new_F1851_, new_F1852_, new_F1853_, new_F1854_, new_F1855_, new_F1856_,
    new_F1857_, new_F1858_, new_F1859_, new_F1860_, new_F1861_, new_F1862_,
    new_F1863_, new_F1870_, new_F1871_, new_F1872_, new_F1873_, new_F1874_,
    new_F1875_, new_F1876_, new_F1877_, new_F1878_, new_F1879_, new_F1880_,
    new_F1881_, new_F1882_, new_F1883_, new_F1884_, new_F1885_, new_F1886_,
    new_F1887_, new_F1888_, new_F1889_, new_F1890_, new_F1891_, new_F1892_,
    new_F1893_, new_F1894_, new_F1895_, new_F1896_, new_F1897_, new_F1898_,
    new_F1899_, new_F1900_, new_F1901_, new_F1902_, new_F1903_, new_F1904_,
    new_F1905_, new_F1906_, new_F1907_, new_F1908_, new_F1909_, new_F1910_,
    new_F1911_, new_F1912_, new_F1913_, new_F1914_, new_F1915_, new_F1916_,
    new_F1917_, new_F1918_, new_F1919_, new_F1920_, new_F1921_, new_F1922_,
    new_F1923_, new_F1924_, new_F1925_, new_F1926_, new_F1927_, new_F1928_,
    new_F1929_, new_F1930_, new_F1937_, new_F1938_, new_F1939_, new_F1940_,
    new_F1941_, new_F1942_, new_F1943_, new_F1944_, new_F1945_, new_F1946_,
    new_F1947_, new_F1948_, new_F1949_, new_F1950_, new_F1951_, new_F1952_,
    new_F1953_, new_F1954_, new_F1955_, new_F1956_, new_F1957_, new_F1958_,
    new_F1959_, new_F1960_, new_F1961_, new_F1962_, new_F1963_, new_F1964_,
    new_F1965_, new_F1966_, new_F1967_, new_F1968_, new_F1969_, new_F1970_,
    new_F1971_, new_F1972_, new_F1973_, new_F1974_, new_F1975_, new_F1976_,
    new_F1977_, new_F1978_, new_F1979_, new_F1980_, new_F1981_, new_F1982_,
    new_F1983_, new_F1984_, new_F1985_, new_F1986_, new_F1987_, new_F1988_,
    new_F1989_, new_F1990_, new_F1991_, new_F1992_, new_F1993_, new_F1994_,
    new_F1995_, new_F1996_, new_F1997_, new_F2004_, new_F2005_, new_F2006_,
    new_F2007_, new_F2008_, new_F2009_, new_F2010_, new_F2011_, new_F2012_,
    new_F2013_, new_F2014_, new_F2015_, new_F2016_, new_F2017_, new_F2018_,
    new_F2019_, new_F2020_, new_F2021_, new_F2022_, new_F2023_, new_F2024_,
    new_F2025_, new_F2026_, new_F2027_, new_F2028_, new_F2029_, new_F2030_,
    new_F2031_, new_F2032_, new_F2033_, new_F2034_, new_F2035_, new_F2036_,
    new_F2037_, new_F2038_, new_F2039_, new_F2040_, new_F2041_, new_F2042_,
    new_F2043_, new_F2044_, new_F2045_, new_F2046_, new_F2047_, new_F2048_,
    new_F2049_, new_F2050_, new_F2051_, new_F2052_, new_F2053_, new_F2054_,
    new_F2055_, new_F2056_, new_F2057_, new_F2058_, new_F2059_, new_F2060_,
    new_F2061_, new_F2062_, new_F2063_, new_F2064_, new_F2071_, new_F2072_,
    new_F2073_, new_F2074_, new_F2075_, new_F2076_, new_F2077_, new_F2078_,
    new_F2079_, new_F2080_, new_F2081_, new_F2082_, new_F2083_, new_F2084_,
    new_F2085_, new_F2086_, new_F2087_, new_F2088_, new_F2089_, new_F2090_,
    new_F2091_, new_F2092_, new_F2093_, new_F2094_, new_F2095_, new_F2096_,
    new_F2097_, new_F2098_, new_F2099_, new_F2100_, new_F2101_, new_F2102_,
    new_F2103_, new_F2104_, new_F2105_, new_F2106_, new_F2107_, new_F2108_,
    new_F2109_, new_F2110_, new_F2111_, new_F2112_, new_F2113_, new_F2114_,
    new_F2115_, new_F2116_, new_F2117_, new_F2118_, new_F2119_, new_F2120_,
    new_F2121_, new_F2122_, new_F2123_, new_F2124_, new_F2125_, new_F2126_,
    new_F2127_, new_F2128_, new_F2129_, new_F2130_, new_F2131_, new_F2138_,
    new_F2139_, new_F2140_, new_F2141_, new_F2142_, new_F2143_, new_F2144_,
    new_F2145_, new_F2146_, new_F2147_, new_F2148_, new_F2149_, new_F2150_,
    new_F2151_, new_F2152_, new_F2153_, new_F2154_, new_F2155_, new_F2156_,
    new_F2157_, new_F2158_, new_F2159_, new_F2160_, new_F2161_, new_F2162_,
    new_F2163_, new_F2164_, new_F2165_, new_F2166_, new_F2167_, new_F2168_,
    new_F2169_, new_F2170_, new_F2171_, new_F2172_, new_F2173_, new_F2174_,
    new_F2175_, new_F2176_, new_F2177_, new_F2178_, new_F2179_, new_F2180_,
    new_F2181_, new_F2182_, new_F2183_, new_F2184_, new_F2185_, new_F2186_,
    new_F2187_, new_F2188_, new_F2189_, new_F2190_, new_F2191_, new_F2192_,
    new_F2193_, new_F2194_, new_F2195_, new_F2196_, new_F2197_, new_F2198_,
    new_F2205_, new_F2206_, new_F2207_, new_F2208_, new_F2209_, new_F2210_,
    new_F2211_, new_F2212_, new_F2213_, new_F2214_, new_F2215_, new_F2216_,
    new_F2217_, new_F2218_, new_F2219_, new_F2220_, new_F2221_, new_F2222_,
    new_F2223_, new_F2224_, new_F2225_, new_F2226_, new_F2227_, new_F2228_,
    new_F2229_, new_F2230_, new_F2231_, new_F2232_, new_F2233_, new_F2234_,
    new_F2235_, new_F2236_, new_F2237_, new_F2238_, new_F2239_, new_F2240_,
    new_F2241_, new_F2242_, new_F2243_, new_F2244_, new_F2245_, new_F2246_,
    new_F2247_, new_F2248_, new_F2249_, new_F2250_, new_F2251_, new_F2252_,
    new_F2253_, new_F2254_, new_F2255_, new_F2256_, new_F2257_, new_F2258_,
    new_F2259_, new_F2260_, new_F2261_, new_F2262_, new_F2263_, new_F2264_,
    new_F2265_, new_F2272_, new_F2273_, new_F2274_, new_F2275_, new_F2276_,
    new_F2277_, new_F2278_, new_F2279_, new_F2280_, new_F2281_, new_F2282_,
    new_F2283_, new_F2284_, new_F2285_, new_F2286_, new_F2287_, new_F2288_,
    new_F2289_, new_F2290_, new_F2291_, new_F2292_, new_F2293_, new_F2294_,
    new_F2295_, new_F2296_, new_F2297_, new_F2298_, new_F2299_, new_F2300_,
    new_F2301_, new_F2302_, new_F2303_, new_F2304_, new_F2305_, new_F2306_,
    new_F2307_, new_F2308_, new_F2309_, new_F2310_, new_F2311_, new_F2312_,
    new_F2313_, new_F2314_, new_F2315_, new_F2316_, new_F2317_, new_F2318_,
    new_F2319_, new_F2320_, new_F2321_, new_F2322_, new_F2323_, new_F2324_,
    new_F2325_, new_F2326_, new_F2327_, new_F2328_, new_F2329_, new_F2330_,
    new_F2331_, new_F2332_, new_F2339_, new_F2340_, new_F2341_, new_F2342_,
    new_F2343_, new_F2344_, new_F2345_, new_F2346_, new_F2347_, new_F2348_,
    new_F2349_, new_F2350_, new_F2351_, new_F2352_, new_F2353_, new_F2354_,
    new_F2355_, new_F2356_, new_F2357_, new_F2358_, new_F2359_, new_F2360_,
    new_F2361_, new_F2362_, new_F2363_, new_F2364_, new_F2365_, new_F2366_,
    new_F2367_, new_F2368_, new_F2369_, new_F2370_, new_F2371_, new_F2372_,
    new_F2373_, new_F2374_, new_F2375_, new_F2376_, new_F2377_, new_F2378_,
    new_F2379_, new_F2380_, new_F2381_, new_F2382_, new_F2383_, new_F2384_,
    new_F2385_, new_F2386_, new_F2387_, new_F2388_, new_F2389_, new_F2390_,
    new_F2391_, new_F2392_, new_F2393_, new_F2394_, new_F2395_, new_F2396_,
    new_F2397_, new_F2398_, new_F2399_, new_F2406_, new_F2407_, new_F2408_,
    new_F2409_, new_F2410_, new_F2411_, new_F2412_, new_F2413_, new_F2414_,
    new_F2415_, new_F2416_, new_F2417_, new_F2418_, new_F2419_, new_F2420_,
    new_F2421_, new_F2422_, new_F2423_, new_F2424_, new_F2425_, new_F2426_,
    new_F2427_, new_F2428_, new_F2429_, new_F2430_, new_F2431_, new_F2432_,
    new_F2433_, new_F2434_, new_F2435_, new_F2436_, new_F2437_, new_F2438_,
    new_F2439_, new_F2440_, new_F2441_, new_F2442_, new_F2443_, new_F2444_,
    new_F2445_, new_F2446_, new_F2447_, new_F2448_, new_F2449_, new_F2450_,
    new_F2451_, new_F2452_, new_F2453_, new_F2454_, new_F2455_, new_F2456_,
    new_F2457_, new_F2458_, new_F2459_, new_F2460_, new_F2461_, new_F2462_,
    new_F2463_, new_F2464_, new_F2465_, new_F2466_, new_F2473_, new_F2474_,
    new_F2475_, new_F2476_, new_F2477_, new_F2478_, new_F2479_, new_F2480_,
    new_F2481_, new_F2482_, new_F2483_, new_F2484_, new_F2485_, new_F2486_,
    new_F2487_, new_F2488_, new_F2489_, new_F2490_, new_F2491_, new_F2492_,
    new_F2493_, new_F2494_, new_F2495_, new_F2496_, new_F2497_, new_F2498_,
    new_F2499_, new_F2500_, new_F2501_, new_F2502_, new_F2503_, new_F2504_,
    new_F2505_, new_F2506_, new_F2507_, new_F2508_, new_F2509_, new_F2510_,
    new_F2511_, new_F2512_, new_F2513_, new_F2514_, new_F2515_, new_F2516_,
    new_F2517_, new_F2518_, new_F2519_, new_F2520_, new_F2521_, new_F2522_,
    new_F2523_, new_F2524_, new_F2525_, new_F2526_, new_F2527_, new_F2528_,
    new_F2529_, new_F2530_, new_F2531_, new_F2532_, new_F2533_, new_F2540_,
    new_F2541_, new_F2542_, new_F2543_, new_F2544_, new_F2545_, new_F2546_,
    new_F2547_, new_F2548_, new_F2549_, new_F2550_, new_F2551_, new_F2552_,
    new_F2553_, new_F2554_, new_F2555_, new_F2556_, new_F2557_, new_F2558_,
    new_F2559_, new_F2560_, new_F2561_, new_F2562_, new_F2563_, new_F2564_,
    new_F2565_, new_F2566_, new_F2567_, new_F2568_, new_F2569_, new_F2570_,
    new_F2571_, new_F2572_, new_F2573_, new_F2574_, new_F2575_, new_F2576_,
    new_F2577_, new_F2578_, new_F2579_, new_F2580_, new_F2581_, new_F2582_,
    new_F2583_, new_F2584_, new_F2585_, new_F2586_, new_F2587_, new_F2588_,
    new_F2589_, new_F2590_, new_F2591_, new_F2592_, new_F2593_, new_F2594_,
    new_F2595_, new_F2596_, new_F2597_, new_F2598_, new_F2599_, new_F2600_,
    new_F2607_, new_F2608_, new_F2609_, new_F2610_, new_F2611_, new_F2612_,
    new_F2613_, new_F2614_, new_F2615_, new_F2616_, new_F2617_, new_F2618_,
    new_F2619_, new_F2620_, new_F2621_, new_F2622_, new_F2623_, new_F2624_,
    new_F2625_, new_F2626_, new_F2627_, new_F2628_, new_F2629_, new_F2630_,
    new_F2631_, new_F2632_, new_F2633_, new_F2634_, new_F2635_, new_F2636_,
    new_F2637_, new_F2638_, new_F2639_, new_F2640_, new_F2641_, new_F2642_,
    new_F2643_, new_F2644_, new_F2645_, new_F2646_, new_F2647_, new_F2648_,
    new_F2649_, new_F2650_, new_F2651_, new_F2652_, new_F2653_, new_F2654_,
    new_F2655_, new_F2656_, new_F2657_, new_F2658_, new_F2659_, new_F2660_,
    new_F2661_, new_F2662_, new_F2663_, new_F2664_, new_F2665_, new_F2666_,
    new_F2667_, new_F2674_, new_F2675_, new_F2676_, new_F2677_, new_F2678_,
    new_F2679_, new_F2680_, new_F2681_, new_F2682_, new_F2683_, new_F2684_,
    new_F2685_, new_F2686_, new_F2687_, new_F2688_, new_F2689_, new_F2690_,
    new_F2691_, new_F2692_, new_F2693_, new_F2694_, new_F2695_, new_F2696_,
    new_F2697_, new_F2698_, new_F2699_, new_F2700_, new_F2701_, new_F2702_,
    new_F2703_, new_F2704_, new_F2705_, new_F2706_, new_F2707_, new_F2708_,
    new_F2709_, new_F2710_, new_F2711_, new_F2712_, new_F2713_, new_F2714_,
    new_F2715_, new_F2716_, new_F2717_, new_F2718_, new_F2719_, new_F2720_,
    new_F2721_, new_F2722_, new_F2723_, new_F2724_, new_F2725_, new_F2726_,
    new_F2727_, new_F2728_, new_F2729_, new_F2730_, new_F2731_, new_F2732_,
    new_F2733_, new_F2734_, new_F2741_, new_F2742_, new_F2743_, new_F2744_,
    new_F2745_, new_F2746_, new_F2747_, new_F2748_, new_F2749_, new_F2750_,
    new_F2751_, new_F2752_, new_F2753_, new_F2754_, new_F2755_, new_F2756_,
    new_F2757_, new_F2758_, new_F2759_, new_F2760_, new_F2761_, new_F2762_,
    new_F2763_, new_F2764_, new_F2765_, new_F2766_, new_F2767_, new_F2768_,
    new_F2769_, new_F2770_, new_F2771_, new_F2772_, new_F2773_, new_F2774_,
    new_F2775_, new_F2776_, new_F2777_, new_F2778_, new_F2779_, new_F2780_,
    new_F2781_, new_F2782_, new_F2783_, new_F2784_, new_F2785_, new_F2786_,
    new_F2787_, new_F2788_, new_F2789_, new_F2790_, new_F2791_, new_F2792_,
    new_F2793_, new_F2794_, new_F2795_, new_F2796_, new_F2797_, new_F2798_,
    new_F2799_, new_F2800_, new_F2801_, new_F2808_, new_F2809_, new_F2810_,
    new_F2811_, new_F2812_, new_F2813_, new_F2814_, new_F2815_, new_F2816_,
    new_F2817_, new_F2818_, new_F2819_, new_F2820_, new_F2821_, new_F2822_,
    new_F2823_, new_F2824_, new_F2825_, new_F2826_, new_F2827_, new_F2828_,
    new_F2829_, new_F2830_, new_F2831_, new_F2832_, new_F2833_, new_F2834_,
    new_F2835_, new_F2836_, new_F2837_, new_F2838_, new_F2839_, new_F2840_,
    new_F2841_, new_F2842_, new_F2843_, new_F2844_, new_F2845_, new_F2846_,
    new_F2847_, new_F2848_, new_F2849_, new_F2850_, new_F2851_, new_F2852_,
    new_F2853_, new_F2854_, new_F2855_, new_F2856_, new_F2857_, new_F2858_,
    new_F2859_, new_F2860_, new_F2861_, new_F2862_, new_F2863_, new_F2864_,
    new_F2865_, new_F2866_, new_F2867_, new_F2868_, new_F2875_, new_F2876_,
    new_F2877_, new_F2878_, new_F2879_, new_F2880_, new_F2881_, new_F2882_,
    new_F2883_, new_F2884_, new_F2885_, new_F2886_, new_F2887_, new_F2888_,
    new_F2889_, new_F2890_, new_F2891_, new_F2892_, new_F2893_, new_F2894_,
    new_F2895_, new_F2896_, new_F2897_, new_F2898_, new_F2899_, new_F2900_,
    new_F2901_, new_F2902_, new_F2903_, new_F2904_, new_F2905_, new_F2906_,
    new_F2907_, new_F2908_, new_F2909_, new_F2910_, new_F2911_, new_F2912_,
    new_F2913_, new_F2914_, new_F2915_, new_F2916_, new_F2917_, new_F2918_,
    new_F2919_, new_F2920_, new_F2921_, new_F2922_, new_F2923_, new_F2924_,
    new_F2925_, new_F2926_, new_F2927_, new_F2928_, new_F2929_, new_F2930_,
    new_F2931_, new_F2932_, new_F2933_, new_F2934_, new_F2935_, new_F2942_,
    new_F2943_, new_F2944_, new_F2945_, new_F2946_, new_F2947_, new_F2948_,
    new_F2949_, new_F2950_, new_F2951_, new_F2952_, new_F2953_, new_F2954_,
    new_F2955_, new_F2956_, new_F2957_, new_F2958_, new_F2959_, new_F2960_,
    new_F2961_, new_F2962_, new_F2963_, new_F2964_, new_F2965_, new_F2966_,
    new_F2967_, new_F2968_, new_F2969_, new_F2970_, new_F2971_, new_F2972_,
    new_F2973_, new_F2974_, new_F2975_, new_F2976_, new_F2977_, new_F2978_,
    new_F2979_, new_F2980_, new_F2981_, new_F2982_, new_F2983_, new_F2984_,
    new_F2985_, new_F2986_, new_F2987_, new_F2988_, new_F2989_, new_F2990_,
    new_F2991_, new_F2992_, new_F2993_, new_F2994_, new_F2995_, new_F2996_,
    new_F2997_, new_F2998_, new_F2999_, new_F3000_, new_F3001_, new_F3002_,
    new_F3009_, new_F3010_, new_F3011_, new_F3012_, new_F3013_, new_F3014_,
    new_F3015_, new_F3016_, new_F3017_, new_F3018_, new_F3019_, new_F3020_,
    new_F3021_, new_F3022_, new_F3023_, new_F3024_, new_F3025_, new_F3026_,
    new_F3027_, new_F3028_, new_F3029_, new_F3030_, new_F3031_, new_F3032_,
    new_F3033_, new_F3034_, new_F3035_, new_F3036_, new_F3037_, new_F3038_,
    new_F3039_, new_F3040_, new_F3041_, new_F3042_, new_F3043_, new_F3044_,
    new_F3045_, new_F3046_, new_F3047_, new_F3048_, new_F3049_, new_F3050_,
    new_F3051_, new_F3052_, new_F3053_, new_F3054_, new_F3055_, new_F3056_,
    new_F3057_, new_F3058_, new_F3059_, new_F3060_, new_F3061_, new_F3062_,
    new_F3063_, new_F3064_, new_F3065_, new_F3066_, new_F3067_, new_F3068_,
    new_F3069_, new_F3076_, new_F3077_, new_F3078_, new_F3079_, new_F3080_,
    new_F3081_, new_F3082_, new_F3083_, new_F3084_, new_F3085_, new_F3086_,
    new_F3087_, new_F3088_, new_F3089_, new_F3090_, new_F3091_, new_F3092_,
    new_F3093_, new_F3094_, new_F3095_, new_F3096_, new_F3097_, new_F3098_,
    new_F3099_, new_F3100_, new_F3101_, new_F3102_, new_F3103_, new_F3104_,
    new_F3105_, new_F3106_, new_F3107_, new_F3108_, new_F3109_, new_F3110_,
    new_F3111_, new_F3112_, new_F3113_, new_F3114_, new_F3115_, new_F3116_,
    new_F3117_, new_F3118_, new_F3119_, new_F3120_, new_F3121_, new_F3122_,
    new_F3123_, new_F3124_, new_F3125_, new_F3126_, new_F3127_, new_F3128_,
    new_F3129_, new_F3130_, new_F3131_, new_F3132_, new_F3133_, new_F3134_,
    new_F3135_, new_F3136_, new_F3143_, new_F3144_, new_F3145_, new_F3146_,
    new_F3147_, new_F3148_, new_F3149_, new_F3150_, new_F3151_, new_F3152_,
    new_F3153_, new_F3154_, new_F3155_, new_F3156_, new_F3157_, new_F3158_,
    new_F3159_, new_F3160_, new_F3161_, new_F3162_, new_F3163_, new_F3164_,
    new_F3165_, new_F3166_, new_F3167_, new_F3168_, new_F3169_, new_F3170_,
    new_F3171_, new_F3172_, new_F3173_, new_F3174_, new_F3175_, new_F3176_,
    new_F3177_, new_F3178_, new_F3179_, new_F3180_, new_F3181_, new_F3182_,
    new_F3183_, new_F3184_, new_F3185_, new_F3186_, new_F3187_, new_F3188_,
    new_F3189_, new_F3190_, new_F3191_, new_F3192_, new_F3193_, new_F3194_,
    new_F3195_, new_F3196_, new_F3197_, new_F3198_, new_F3199_, new_F3200_,
    new_F3201_, new_F3202_, new_F3203_, new_F3210_, new_F3211_, new_F3212_,
    new_F3213_, new_F3214_, new_F3215_, new_F3216_, new_F3217_, new_F3218_,
    new_F3219_, new_F3220_, new_F3221_, new_F3222_, new_F3223_, new_F3224_,
    new_F3225_, new_F3226_, new_F3227_, new_F3228_, new_F3229_, new_F3230_,
    new_F3231_, new_F3232_, new_F3233_, new_F3234_, new_F3235_, new_F3236_,
    new_F3237_, new_F3238_, new_F3239_, new_F3240_, new_F3241_, new_F3242_,
    new_F3243_, new_F3244_, new_F3245_, new_F3246_, new_F3247_, new_F3248_,
    new_F3249_, new_F3250_, new_F3251_, new_F3252_, new_F3253_, new_F3254_,
    new_F3255_, new_F3256_, new_F3257_, new_F3258_, new_F3259_, new_F3260_,
    new_F3261_, new_F3262_, new_F3263_, new_F3264_, new_F3265_, new_F3266_,
    new_F3267_, new_F3268_, new_F3269_, new_F3270_, new_F3277_, new_F3278_,
    new_F3279_, new_F3280_, new_F3281_, new_F3282_, new_F3283_, new_F3284_,
    new_F3285_, new_F3286_, new_F3287_, new_F3288_, new_F3289_, new_F3290_,
    new_F3291_, new_F3292_, new_F3293_, new_F3294_, new_F3295_, new_F3296_,
    new_F3297_, new_F3298_, new_F3299_, new_F3300_, new_F3301_, new_F3302_,
    new_F3303_, new_F3304_, new_F3305_, new_F3306_, new_F3307_, new_F3308_,
    new_F3309_, new_F3310_, new_F3311_, new_F3312_, new_F3313_, new_F3314_,
    new_F3315_, new_F3316_, new_F3317_, new_F3318_, new_F3319_, new_F3320_,
    new_F3321_, new_F3322_, new_F3323_, new_F3324_, new_F3325_, new_F3326_,
    new_F3327_, new_F3328_, new_F3329_, new_F3330_, new_F3331_, new_F3332_,
    new_F3333_, new_F3334_, new_F3335_, new_F3336_, new_F3337_, new_F3344_,
    new_F3345_, new_F3346_, new_F3347_, new_F3348_, new_F3349_, new_F3350_,
    new_F3351_, new_F3352_, new_F3353_, new_F3354_, new_F3355_, new_F3356_,
    new_F3357_, new_F3358_, new_F3359_, new_F3360_, new_F3361_, new_F3362_,
    new_F3363_, new_F3364_, new_F3365_, new_F3366_, new_F3367_, new_F3368_,
    new_F3369_, new_F3370_, new_F3371_, new_F3372_, new_F3373_, new_F3374_,
    new_F3375_, new_F3376_, new_F3377_, new_F3378_, new_F3379_, new_F3380_,
    new_F3381_, new_F3382_, new_F3383_, new_F3384_, new_F3385_, new_F3386_,
    new_F3387_, new_F3388_, new_F3389_, new_F3390_, new_F3391_, new_F3392_,
    new_F3393_, new_F3394_, new_F3395_, new_F3396_, new_F3397_, new_F3398_,
    new_F3399_, new_F3400_, new_F3401_, new_F3402_, new_F3403_, new_F3404_,
    new_F3411_, new_F3412_, new_F3413_, new_F3414_, new_F3415_, new_F3416_,
    new_F3417_, new_F3418_, new_F3419_, new_F3420_, new_F3421_, new_F3422_,
    new_F3423_, new_F3424_, new_F3425_, new_F3426_, new_F3427_, new_F3428_,
    new_F3429_, new_F3430_, new_F3431_, new_F3432_, new_F3433_, new_F3434_,
    new_F3435_, new_F3436_, new_F3437_, new_F3438_, new_F3439_, new_F3440_,
    new_F3441_, new_F3442_, new_F3443_, new_F3444_, new_F3445_, new_F3446_,
    new_F3447_, new_F3448_, new_F3449_, new_F3450_, new_F3451_, new_F3452_,
    new_F3453_, new_F3454_, new_F3455_, new_F3456_, new_F3457_, new_F3458_,
    new_F3459_, new_F3460_, new_F3461_, new_F3462_, new_F3463_, new_F3464_,
    new_F3465_, new_F3466_, new_F3467_, new_F3468_, new_F3469_, new_F3470_,
    new_F3471_, new_F3478_, new_F3479_, new_F3480_, new_F3481_, new_F3482_,
    new_F3483_, new_F3484_, new_F3485_, new_F3486_, new_F3487_, new_F3488_,
    new_F3489_, new_F3490_, new_F3491_, new_F3492_, new_F3493_, new_F3494_,
    new_F3495_, new_F3496_, new_F3497_, new_F3498_, new_F3499_, new_F3500_,
    new_F3501_, new_F3502_, new_F3503_, new_F3504_, new_F3505_, new_F3506_,
    new_F3507_, new_F3508_, new_F3509_, new_F3510_, new_F3511_, new_F3512_,
    new_F3513_, new_F3514_, new_F3515_, new_F3516_, new_F3517_, new_F3518_,
    new_F3519_, new_F3520_, new_F3521_, new_F3522_, new_F3523_, new_F3524_,
    new_F3525_, new_F3526_, new_F3527_, new_F3528_, new_F3529_, new_F3530_,
    new_F3531_, new_F3532_, new_F3533_, new_F3534_, new_F3535_, new_F3536_,
    new_F3537_, new_F3538_, new_F3545_, new_F3546_, new_F3547_, new_F3548_,
    new_F3549_, new_F3550_, new_F3551_, new_F3552_, new_F3553_, new_F3554_,
    new_F3555_, new_F3556_, new_F3557_, new_F3558_, new_F3559_, new_F3560_,
    new_F3561_, new_F3562_, new_F3563_, new_F3564_, new_F3565_, new_F3566_,
    new_F3567_, new_F3568_, new_F3569_, new_F3570_, new_F3571_, new_F3572_,
    new_F3573_, new_F3574_, new_F3575_, new_F3576_, new_F3577_, new_F3578_,
    new_F3579_, new_F3580_, new_F3581_, new_F3582_, new_F3583_, new_F3584_,
    new_F3585_, new_F3586_, new_F3587_, new_F3588_, new_F3589_, new_F3590_,
    new_F3591_, new_F3592_, new_F3593_, new_F3594_, new_F3595_, new_F3596_,
    new_F3597_, new_F3598_, new_F3599_, new_F3600_, new_F3601_, new_F3602_,
    new_F3603_, new_F3604_, new_F3605_, new_F3612_, new_F3613_, new_F3614_,
    new_F3615_, new_F3616_, new_F3617_, new_F3618_, new_F3619_, new_F3620_,
    new_F3621_, new_F3622_, new_F3623_, new_F3624_, new_F3625_, new_F3626_,
    new_F3627_, new_F3628_, new_F3629_, new_F3630_, new_F3631_, new_F3632_,
    new_F3633_, new_F3634_, new_F3635_, new_F3636_, new_F3637_, new_F3638_,
    new_F3639_, new_F3640_, new_F3641_, new_F3642_, new_F3643_, new_F3644_,
    new_F3645_, new_F3646_, new_F3647_, new_F3648_, new_F3649_, new_F3650_,
    new_F3651_, new_F3652_, new_F3653_, new_F3654_, new_F3655_, new_F3656_,
    new_F3657_, new_F3658_, new_F3659_, new_F3660_, new_F3661_, new_F3662_,
    new_F3663_, new_F3664_, new_F3665_, new_F3666_, new_F3667_, new_F3668_,
    new_F3669_, new_F3670_, new_F3671_, new_F3672_, new_F3679_, new_F3680_,
    new_F3681_, new_F3682_, new_F3683_, new_F3684_, new_F3685_, new_F3686_,
    new_F3687_, new_F3688_, new_F3689_, new_F3690_, new_F3691_, new_F3692_,
    new_F3693_, new_F3694_, new_F3695_, new_F3696_, new_F3697_, new_F3698_,
    new_F3699_, new_F3700_, new_F3701_, new_F3702_, new_F3703_, new_F3704_,
    new_F3705_, new_F3706_, new_F3707_, new_F3708_, new_F3709_, new_F3710_,
    new_F3711_, new_F3712_, new_F3713_, new_F3714_, new_F3715_, new_F3716_,
    new_F3717_, new_F3718_, new_F3719_, new_F3720_, new_F3721_, new_F3722_,
    new_F3723_, new_F3724_, new_F3725_, new_F3726_, new_F3727_, new_F3728_,
    new_F3729_, new_F3730_, new_F3731_, new_F3732_, new_F3733_, new_F3734_,
    new_F3735_, new_F3736_, new_F3737_, new_F3738_, new_F3739_, new_F3746_,
    new_F3747_, new_F3748_, new_F3749_, new_F3750_, new_F3751_, new_F3752_,
    new_F3753_, new_F3754_, new_F3755_, new_F3756_, new_F3757_, new_F3758_,
    new_F3759_, new_F3760_, new_F3761_, new_F3762_, new_F3763_, new_F3764_,
    new_F3765_, new_F3766_, new_F3767_, new_F3768_, new_F3769_, new_F3770_,
    new_F3771_, new_F3772_, new_F3773_, new_F3774_, new_F3775_, new_F3776_,
    new_F3777_, new_F3778_, new_F3779_, new_F3780_, new_F3781_, new_F3782_,
    new_F3783_, new_F3784_, new_F3785_, new_F3786_, new_F3787_, new_F3788_,
    new_F3789_, new_F3790_, new_F3791_, new_F3792_, new_F3793_, new_F3794_,
    new_F3795_, new_F3796_, new_F3797_, new_F3798_, new_F3799_, new_F3800_,
    new_F3801_, new_F3802_, new_F3803_, new_F3804_, new_F3805_, new_F3806_,
    new_F3813_, new_F3814_, new_F3815_, new_F3816_, new_F3817_, new_F3818_,
    new_F3819_, new_F3820_, new_F3821_, new_F3822_, new_F3823_, new_F3824_,
    new_F3825_, new_F3826_, new_F3827_, new_F3828_, new_F3829_, new_F3830_,
    new_F3831_, new_F3832_, new_F3833_, new_F3834_, new_F3835_, new_F3836_,
    new_F3837_, new_F3838_, new_F3839_, new_F3840_, new_F3841_, new_F3842_,
    new_F3843_, new_F3844_, new_F3845_, new_F3846_, new_F3847_, new_F3848_,
    new_F3849_, new_F3850_, new_F3851_, new_F3852_, new_F3853_, new_F3854_,
    new_F3855_, new_F3856_, new_F3857_, new_F3858_, new_F3859_, new_F3860_,
    new_F3861_, new_F3862_, new_F3863_, new_F3864_, new_F3865_, new_F3866_,
    new_F3867_, new_F3868_, new_F3869_, new_F3870_, new_F3871_, new_F3872_,
    new_F3873_, new_F3880_, new_F3881_, new_F3882_, new_F3883_, new_F3884_,
    new_F3885_, new_F3886_, new_F3887_, new_F3888_, new_F3889_, new_F3890_,
    new_F3891_, new_F3892_, new_F3893_, new_F3894_, new_F3895_, new_F3896_,
    new_F3897_, new_F3898_, new_F3899_, new_F3900_, new_F3901_, new_F3902_,
    new_F3903_, new_F3904_, new_F3905_, new_F3906_, new_F3907_, new_F3908_,
    new_F3909_, new_F3910_, new_F3911_, new_F3912_, new_F3913_, new_F3914_,
    new_F3915_, new_F3916_, new_F3917_, new_F3918_, new_F3919_, new_F3920_,
    new_F3921_, new_F3922_, new_F3923_, new_F3924_, new_F3925_, new_F3926_,
    new_F3927_, new_F3928_, new_F3929_, new_F3930_, new_F3931_, new_F3932_,
    new_F3933_, new_F3934_, new_F3935_, new_F3936_, new_F3937_, new_F3938_,
    new_F3939_, new_F3940_, new_F3947_, new_F3948_, new_F3949_, new_F3950_,
    new_F3951_, new_F3952_, new_F3953_, new_F3954_, new_F3955_, new_F3956_,
    new_F3957_, new_F3958_, new_F3959_, new_F3960_, new_F3961_, new_F3962_,
    new_F3963_, new_F3964_, new_F3965_, new_F3966_, new_F3967_, new_F3968_,
    new_F3969_, new_F3970_, new_F3971_, new_F3972_, new_F3973_, new_F3974_,
    new_F3975_, new_F3976_, new_F3977_, new_F3978_, new_F3979_, new_F3980_,
    new_F3981_, new_F3982_, new_F3983_, new_F3984_, new_F3985_, new_F3986_,
    new_F3987_, new_F3988_, new_F3989_, new_F3990_, new_F3991_, new_F3992_,
    new_F3993_, new_F3994_, new_F3995_, new_F3996_, new_F3997_, new_F3998_,
    new_F3999_, new_F4000_, new_F4001_, new_F4002_, new_F4003_, new_F4004_,
    new_F4005_, new_F4006_, new_F4007_, new_F4014_, new_F4015_, new_F4016_,
    new_F4017_, new_F4018_, new_F4019_, new_F4020_, new_F4021_, new_F4022_,
    new_F4023_, new_F4024_, new_F4025_, new_F4026_, new_F4027_, new_F4028_,
    new_F4029_, new_F4030_, new_F4031_, new_F4032_, new_F4033_, new_F4034_,
    new_F4035_, new_F4036_, new_F4037_, new_F4038_, new_F4039_, new_F4040_,
    new_F4041_, new_F4042_, new_F4043_, new_F4044_, new_F4045_, new_F4046_,
    new_F4047_, new_F4048_, new_F4049_, new_F4050_, new_F4051_, new_F4052_,
    new_F4053_, new_F4054_, new_F4055_, new_F4056_, new_F4057_, new_F4058_,
    new_F4059_, new_F4060_, new_F4061_, new_F4062_, new_F4063_, new_F4064_,
    new_F4065_, new_F4066_, new_F4067_, new_F4068_, new_F4069_, new_F4070_,
    new_F4071_, new_F4072_, new_F4073_, new_F4074_, new_F4081_, new_F4082_,
    new_F4083_, new_F4084_, new_F4085_, new_F4086_, new_F4087_, new_F4088_,
    new_F4089_, new_F4090_, new_F4091_, new_F4092_, new_F4093_, new_F4094_,
    new_F4095_, new_F4096_, new_F4097_, new_F4098_, new_F4099_, new_F4100_,
    new_F4101_, new_F4102_, new_F4103_, new_F4104_, new_F4105_, new_F4106_,
    new_F4107_, new_F4108_, new_F4109_, new_F4110_, new_F4111_, new_F4112_,
    new_F4113_, new_F4114_, new_F4115_, new_F4116_, new_F4117_, new_F4118_,
    new_F4119_, new_F4120_, new_F4121_, new_F4122_, new_F4123_, new_F4124_,
    new_F4125_, new_F4126_, new_F4127_, new_F4128_, new_F4129_, new_F4130_,
    new_F4131_, new_F4132_, new_F4133_, new_F4134_, new_F4135_, new_F4136_,
    new_F4137_, new_F4138_, new_F4139_, new_F4140_, new_F4141_, new_F4148_,
    new_F4149_, new_F4150_, new_F4151_, new_F4152_, new_F4153_, new_F4154_,
    new_F4155_, new_F4156_, new_F4157_, new_F4158_, new_F4159_, new_F4160_,
    new_F4161_, new_F4162_, new_F4163_, new_F4164_, new_F4165_, new_F4166_,
    new_F4167_, new_F4168_, new_F4169_, new_F4170_, new_F4171_, new_F4172_,
    new_F4173_, new_F4174_, new_F4175_, new_F4176_, new_F4177_, new_F4178_,
    new_F4179_, new_F4180_, new_F4181_, new_F4182_, new_F4183_, new_F4184_,
    new_F4185_, new_F4186_, new_F4187_, new_F4188_, new_F4189_, new_F4190_,
    new_F4191_, new_F4192_, new_F4193_, new_F4194_, new_F4195_, new_F4196_,
    new_F4197_, new_F4198_, new_F4199_, new_F4200_, new_F4201_, new_F4202_,
    new_F4203_, new_F4204_, new_F4205_, new_F4206_, new_F4207_, new_F4208_,
    new_F4215_, new_F4216_, new_F4217_, new_F4218_, new_F4219_, new_F4220_,
    new_F4221_, new_F4222_, new_F4223_, new_F4224_, new_F4225_, new_F4226_,
    new_F4227_, new_F4228_, new_F4229_, new_F4230_, new_F4231_, new_F4232_,
    new_F4233_, new_F4234_, new_F4235_, new_F4236_, new_F4237_, new_F4238_,
    new_F4239_, new_F4240_, new_F4241_, new_F4242_, new_F4243_, new_F4244_,
    new_F4245_, new_F4246_, new_F4247_, new_F4248_, new_F4249_, new_F4250_,
    new_F4251_, new_F4252_, new_F4253_, new_F4254_, new_F4255_, new_F4256_,
    new_F4257_, new_F4258_, new_F4259_, new_F4260_, new_F4261_, new_F4262_,
    new_F4263_, new_F4264_, new_F4265_, new_F4266_, new_F4267_, new_F4268_,
    new_F4269_, new_F4270_, new_F4271_, new_F4272_, new_F4273_, new_F4274_,
    new_F4275_, new_F4282_, new_F4283_, new_F4284_, new_F4285_, new_F4286_,
    new_F4287_, new_F4288_, new_F4289_, new_F4290_, new_F4291_, new_F4292_,
    new_F4293_, new_F4294_, new_F4295_, new_F4296_, new_F4297_, new_F4298_,
    new_F4299_, new_F4300_, new_F4301_, new_F4302_, new_F4303_, new_F4304_,
    new_F4305_, new_F4306_, new_F4307_, new_F4308_, new_F4309_, new_F4310_,
    new_F4311_, new_F4312_, new_F4313_, new_F4314_, new_F4315_, new_F4316_,
    new_F4317_, new_F4318_, new_F4319_, new_F4320_, new_F4321_, new_F4322_,
    new_F4323_, new_F4324_, new_F4325_, new_F4326_, new_F4327_, new_F4328_,
    new_F4329_, new_F4330_, new_F4331_, new_F4332_, new_F4333_, new_F4334_,
    new_F4335_, new_F4336_, new_F4337_, new_F4338_, new_F4339_, new_F4340_,
    new_F4341_, new_F4342_, new_F4349_, new_F4350_, new_F4351_, new_F4352_,
    new_F4353_, new_F4354_, new_F4355_, new_F4356_, new_F4357_, new_F4358_,
    new_F4359_, new_F4360_, new_F4361_, new_F4362_, new_F4363_, new_F4364_,
    new_F4365_, new_F4366_, new_F4367_, new_F4368_, new_F4369_, new_F4370_,
    new_F4371_, new_F4372_, new_F4373_, new_F4374_, new_F4375_, new_F4376_,
    new_F4377_, new_F4378_, new_F4379_, new_F4380_, new_F4381_, new_F4382_,
    new_F4383_, new_F4384_, new_F4385_, new_F4386_, new_F4387_, new_F4388_,
    new_F4389_, new_F4390_, new_F4391_, new_F4392_, new_F4393_, new_F4394_,
    new_F4395_, new_F4396_, new_F4397_, new_F4398_, new_F4399_, new_F4400_,
    new_F4401_, new_F4402_, new_F4403_, new_F4404_, new_F4405_, new_F4406_,
    new_F4407_, new_F4408_, new_F4409_, new_F4416_, new_F4417_, new_F4418_,
    new_F4419_, new_F4420_, new_F4421_, new_F4422_, new_F4423_, new_F4424_,
    new_F4425_, new_F4426_, new_F4427_, new_F4428_, new_F4429_, new_F4430_,
    new_F4431_, new_F4432_, new_F4433_, new_F4434_, new_F4435_, new_F4436_,
    new_F4437_, new_F4438_, new_F4439_, new_F4440_, new_F4441_, new_F4442_,
    new_F4443_, new_F4444_, new_F4445_, new_F4446_, new_F4447_, new_F4448_,
    new_F4449_, new_F4450_, new_F4451_, new_F4452_, new_F4453_, new_F4454_,
    new_F4455_, new_F4456_, new_F4457_, new_F4458_, new_F4459_, new_F4460_,
    new_F4461_, new_F4462_, new_F4463_, new_F4464_, new_F4465_, new_F4466_,
    new_F4467_, new_F4468_, new_F4469_, new_F4470_, new_F4471_, new_F4472_,
    new_F4473_, new_F4474_, new_F4475_, new_F4476_, new_F4483_, new_F4484_,
    new_F4485_, new_F4486_, new_F4487_, new_F4488_, new_F4489_, new_F4490_,
    new_F4491_, new_F4492_, new_F4493_, new_F4494_, new_F4495_, new_F4496_,
    new_F4497_, new_F4498_, new_F4499_, new_F4500_, new_F4501_, new_F4502_,
    new_F4503_, new_F4504_, new_F4505_, new_F4506_, new_F4507_, new_F4508_,
    new_F4509_, new_F4510_, new_F4511_, new_F4512_, new_F4513_, new_F4514_,
    new_F4515_, new_F4516_, new_F4517_, new_F4518_, new_F4519_, new_F4520_,
    new_F4521_, new_F4522_, new_F4523_, new_F4524_, new_F4525_, new_F4526_,
    new_F4527_, new_F4528_, new_F4529_, new_F4530_, new_F4531_, new_F4532_,
    new_F4533_, new_F4534_, new_F4535_, new_F4536_, new_F4537_, new_F4538_,
    new_F4539_, new_F4540_, new_F4541_, new_F4542_, new_F4543_, new_F4550_,
    new_F4551_, new_F4552_, new_F4553_, new_F4554_, new_F4555_, new_F4556_,
    new_F4557_, new_F4558_, new_F4559_, new_F4560_, new_F4561_, new_F4562_,
    new_F4563_, new_F4564_, new_F4565_, new_F4566_, new_F4567_, new_F4568_,
    new_F4569_, new_F4570_, new_F4571_, new_F4572_, new_F4573_, new_F4574_,
    new_F4575_, new_F4576_, new_F4577_, new_F4578_, new_F4579_, new_F4580_,
    new_F4581_, new_F4582_, new_F4583_, new_F4584_, new_F4585_, new_F4586_,
    new_F4587_, new_F4588_, new_F4589_, new_F4590_, new_F4591_, new_F4592_,
    new_F4593_, new_F4594_, new_F4595_, new_F4596_, new_F4597_, new_F4598_,
    new_F4599_, new_F4600_, new_F4601_, new_F4602_, new_F4603_, new_F4604_,
    new_F4605_, new_F4606_, new_F4607_, new_F4608_, new_F4609_, new_F4610_,
    new_F4617_, new_F4618_, new_F4619_, new_F4620_, new_F4621_, new_F4622_,
    new_F4623_, new_F4624_, new_F4625_, new_F4626_, new_F4627_, new_F4628_,
    new_F4629_, new_F4630_, new_F4631_, new_F4632_, new_F4633_, new_F4634_,
    new_F4635_, new_F4636_, new_F4637_, new_F4638_, new_F4639_, new_F4640_,
    new_F4641_, new_F4642_, new_F4643_, new_F4644_, new_F4645_, new_F4646_,
    new_F4647_, new_F4648_, new_F4649_, new_F4650_, new_F4651_, new_F4652_,
    new_F4653_, new_F4654_, new_F4655_, new_F4656_, new_F4657_, new_F4658_,
    new_F4659_, new_F4660_, new_F4661_, new_F4662_, new_F4663_, new_F4664_,
    new_F4665_, new_F4666_, new_F4667_, new_F4668_, new_F4669_, new_F4670_,
    new_F4671_, new_F4672_, new_F4673_, new_F4674_, new_F4675_, new_F4676_,
    new_F4677_, new_F4684_, new_F4685_, new_F4686_, new_F4687_, new_F4688_,
    new_F4689_, new_F4690_, new_F4691_, new_F4692_, new_F4693_, new_F4694_,
    new_F4695_, new_F4696_, new_F4697_, new_F4698_, new_F4699_, new_F4700_,
    new_F4701_, new_F4702_, new_F4703_, new_F4704_, new_F4705_, new_F4706_,
    new_F4707_, new_F4708_, new_F4709_, new_F4710_, new_F4711_, new_F4712_,
    new_F4713_, new_F4714_, new_F4715_, new_F4716_, new_F4717_, new_F4718_,
    new_F4719_, new_F4720_, new_F4721_, new_F4722_, new_F4723_, new_F4724_,
    new_F4725_, new_F4726_, new_F4727_, new_F4728_, new_F4729_, new_F4730_,
    new_F4731_, new_F4732_, new_F4733_, new_F4734_, new_F4735_, new_F4736_,
    new_F4737_, new_F4738_, new_F4739_, new_F4740_, new_F4741_, new_F4742_,
    new_F4743_, new_F4744_, new_F4751_, new_F4752_, new_F4753_, new_F4754_,
    new_F4755_, new_F4756_, new_F4757_, new_F4758_, new_F4759_, new_F4760_,
    new_F4761_, new_F4762_, new_F4763_, new_F4764_, new_F4765_, new_F4766_,
    new_F4767_, new_F4768_, new_F4769_, new_F4770_, new_F4771_, new_F4772_,
    new_F4773_, new_F4774_, new_F4775_, new_F4776_, new_F4777_, new_F4778_,
    new_F4779_, new_F4780_, new_F4781_, new_F4782_, new_F4783_, new_F4784_,
    new_F4785_, new_F4786_, new_F4787_, new_F4788_, new_F4789_, new_F4790_,
    new_F4791_, new_F4792_, new_F4793_, new_F4794_, new_F4795_, new_F4796_,
    new_F4797_, new_F4798_, new_F4799_, new_F4800_, new_F4801_, new_F4802_,
    new_F4803_, new_F4804_, new_F4805_, new_F4806_, new_F4807_, new_F4808_,
    new_F4809_, new_F4810_, new_F4811_, new_F4818_, new_F4819_, new_F4820_,
    new_F4821_, new_F4822_, new_F4823_, new_F4824_, new_F4825_, new_F4826_,
    new_F4827_, new_F4828_, new_F4829_, new_F4830_, new_F4831_, new_F4832_,
    new_F4833_, new_F4834_, new_F4835_, new_F4836_, new_F4837_, new_F4838_,
    new_F4839_, new_F4840_, new_F4841_, new_F4842_, new_F4843_, new_F4844_,
    new_F4845_, new_F4846_, new_F4847_, new_F4848_, new_F4849_, new_F4850_,
    new_F4851_, new_F4852_, new_F4853_, new_F4854_, new_F4855_, new_F4856_,
    new_F4857_, new_F4858_, new_F4859_, new_F4860_, new_F4861_, new_F4862_,
    new_F4863_, new_F4864_, new_F4865_, new_F4866_, new_F4867_, new_F4868_,
    new_F4869_, new_F4870_, new_F4871_, new_F4872_, new_F4873_, new_F4874_,
    new_F4875_, new_F4876_, new_F4877_, new_F4878_, new_F4885_, new_F4886_,
    new_F4887_, new_F4888_, new_F4889_, new_F4890_, new_F4891_, new_F4892_,
    new_F4893_, new_F4894_, new_F4895_, new_F4896_, new_F4897_, new_F4898_,
    new_F4899_, new_F4900_, new_F4901_, new_F4902_, new_F4903_, new_F4904_,
    new_F4905_, new_F4906_, new_F4907_, new_F4908_, new_F4909_, new_F4910_,
    new_F4911_, new_F4912_, new_F4913_, new_F4914_, new_F4915_, new_F4916_,
    new_F4917_, new_F4918_, new_F4919_, new_F4920_, new_F4921_, new_F4922_,
    new_F4923_, new_F4924_, new_F4925_, new_F4926_, new_F4927_, new_F4928_,
    new_F4929_, new_F4930_, new_F4931_, new_F4932_, new_F4933_, new_F4934_,
    new_F4935_, new_F4936_, new_F4937_, new_F4938_, new_F4939_, new_F4940_,
    new_F4941_, new_F4942_, new_F4943_, new_F4944_, new_F4945_, new_F4952_,
    new_F4953_, new_F4954_, new_F4955_, new_F4956_, new_F4957_, new_F4958_,
    new_F4959_, new_F4960_, new_F4961_, new_F4962_, new_F4963_, new_F4964_,
    new_F4965_, new_F4966_, new_F4967_, new_F4968_, new_F4969_, new_F4970_,
    new_F4971_, new_F4972_, new_F4973_, new_F4974_, new_F4975_, new_F4976_,
    new_F4977_, new_F4978_, new_F4979_, new_F4980_, new_F4981_, new_F4982_,
    new_F4983_, new_F4984_, new_F4985_, new_F4986_, new_F4987_, new_F4988_,
    new_F4989_, new_F4990_, new_F4991_, new_F4992_, new_F4993_, new_F4994_,
    new_F4995_, new_F4996_, new_F4997_, new_F4998_, new_F4999_, new_F5000_,
    new_F5001_, new_F5002_, new_F5003_, new_F5004_, new_F5005_, new_F5006_,
    new_F5007_, new_F5008_, new_F5009_, new_F5010_, new_F5011_, new_F5012_,
    new_F5019_, new_F5020_, new_F5021_, new_F5022_, new_F5023_, new_F5024_,
    new_F5025_, new_F5026_, new_F5027_, new_F5028_, new_F5029_, new_F5030_,
    new_F5031_, new_F5032_, new_F5033_, new_F5034_, new_F5035_, new_F5036_,
    new_F5037_, new_F5038_, new_F5039_, new_F5040_, new_F5041_, new_F5042_,
    new_F5043_, new_F5044_, new_F5045_, new_F5046_, new_F5047_, new_F5048_,
    new_F5049_, new_F5050_, new_F5051_, new_F5052_, new_F5053_, new_F5054_,
    new_F5055_, new_F5056_, new_F5057_, new_F5058_, new_F5059_, new_F5060_,
    new_F5061_, new_F5062_, new_F5063_, new_F5064_, new_F5065_, new_F5066_,
    new_F5067_, new_F5068_, new_F5069_, new_F5070_, new_F5071_, new_F5072_,
    new_F5073_, new_F5074_, new_F5075_, new_F5076_, new_F5077_, new_F5078_,
    new_F5079_, new_F5086_, new_F5087_, new_F5088_, new_F5089_, new_F5090_,
    new_F5091_, new_F5092_, new_F5093_, new_F5094_, new_F5095_, new_F5096_,
    new_F5097_, new_F5098_, new_F5099_, new_F5100_, new_F5101_, new_F5102_,
    new_F5103_, new_F5104_, new_F5105_, new_F5106_, new_F5107_, new_F5108_,
    new_F5109_, new_F5110_, new_F5111_, new_F5112_, new_F5113_, new_F5114_,
    new_F5115_, new_F5116_, new_F5117_, new_F5118_, new_F5119_, new_F5120_,
    new_F5121_, new_F5122_, new_F5123_, new_F5124_, new_F5125_, new_F5126_,
    new_F5127_, new_F5128_, new_F5129_, new_F5130_, new_F5131_, new_F5132_,
    new_F5133_, new_F5134_, new_F5135_, new_F5136_, new_F5137_, new_F5138_,
    new_F5139_, new_F5140_, new_F5141_, new_F5142_, new_F5143_, new_F5144_,
    new_F5145_, new_F5146_, new_F5153_, new_F5154_, new_F5155_, new_F5156_,
    new_F5157_, new_F5158_, new_F5159_, new_F5160_, new_F5161_, new_F5162_,
    new_F5163_, new_F5164_, new_F5165_, new_F5166_, new_F5167_, new_F5168_,
    new_F5169_, new_F5170_, new_F5171_, new_F5172_, new_F5173_, new_F5174_,
    new_F5175_, new_F5176_, new_F5177_, new_F5178_, new_F5179_, new_F5180_,
    new_F5181_, new_F5182_, new_F5183_, new_F5184_, new_F5185_, new_F5186_,
    new_F5187_, new_F5188_, new_F5189_, new_F5190_, new_F5191_, new_F5192_,
    new_F5193_, new_F5194_, new_F5195_, new_F5196_, new_F5197_, new_F5198_,
    new_F5199_, new_F5200_, new_F5201_, new_F5202_, new_F5203_, new_F5204_,
    new_F5205_, new_F5206_, new_F5207_, new_F5208_, new_F5209_, new_F5210_,
    new_F5211_, new_F5212_, new_F5213_, new_F5220_, new_F5221_, new_F5222_,
    new_F5223_, new_F5224_, new_F5225_, new_F5226_, new_F5227_, new_F5228_,
    new_F5229_, new_F5230_, new_F5231_, new_F5232_, new_F5233_, new_F5234_,
    new_F5235_, new_F5236_, new_F5237_, new_F5238_, new_F5239_, new_F5240_,
    new_F5241_, new_F5242_, new_F5243_, new_F5244_, new_F5245_, new_F5246_,
    new_F5247_, new_F5248_, new_F5249_, new_F5250_, new_F5251_, new_F5252_,
    new_F5253_, new_F5254_, new_F5255_, new_F5256_, new_F5257_, new_F5258_,
    new_F5259_, new_F5260_, new_F5261_, new_F5262_, new_F5263_, new_F5264_,
    new_F5265_, new_F5266_, new_F5267_, new_F5268_, new_F5269_, new_F5270_,
    new_F5271_, new_F5272_, new_F5273_, new_F5274_, new_F5275_, new_F5276_,
    new_F5277_, new_F5278_, new_F5279_, new_F5280_, new_F5287_, new_F5288_,
    new_F5289_, new_F5290_, new_F5291_, new_F5292_, new_F5293_, new_F5294_,
    new_F5295_, new_F5296_, new_F5297_, new_F5298_, new_F5299_, new_F5300_,
    new_F5301_, new_F5302_, new_F5303_, new_F5304_, new_F5305_, new_F5306_,
    new_F5307_, new_F5308_, new_F5309_, new_F5310_, new_F5311_, new_F5312_,
    new_F5313_, new_F5314_, new_F5315_, new_F5316_, new_F5317_, new_F5318_,
    new_F5319_, new_F5320_, new_F5321_, new_F5322_, new_F5323_, new_F5324_,
    new_F5325_, new_F5326_, new_F5327_, new_F5328_, new_F5329_, new_F5330_,
    new_F5331_, new_F5332_, new_F5333_, new_F5334_, new_F5335_, new_F5336_,
    new_F5337_, new_F5338_, new_F5339_, new_F5340_, new_F5341_, new_F5342_,
    new_F5343_, new_F5344_, new_F5345_, new_F5346_, new_F5347_, new_F5354_,
    new_F5355_, new_F5356_, new_F5357_, new_F5358_, new_F5359_, new_F5360_,
    new_F5361_, new_F5362_, new_F5363_, new_F5364_, new_F5365_, new_F5366_,
    new_F5367_, new_F5368_, new_F5369_, new_F5370_, new_F5371_, new_F5372_,
    new_F5373_, new_F5374_, new_F5375_, new_F5376_, new_F5377_, new_F5378_,
    new_F5379_, new_F5380_, new_F5381_, new_F5382_, new_F5383_, new_F5384_,
    new_F5385_, new_F5386_, new_F5387_, new_F5388_, new_F5389_, new_F5390_,
    new_F5391_, new_F5392_, new_F5393_, new_F5394_, new_F5395_, new_F5396_,
    new_F5397_, new_F5398_, new_F5399_, new_F5400_, new_F5401_, new_F5402_,
    new_F5403_, new_F5404_, new_F5405_, new_F5406_, new_F5407_, new_F5408_,
    new_F5409_, new_F5410_, new_F5411_, new_F5412_, new_F5413_, new_F5414_,
    new_F5421_, new_F5422_, new_F5423_, new_F5424_, new_F5425_, new_F5426_,
    new_F5427_, new_F5428_, new_F5429_, new_F5430_, new_F5431_, new_F5432_,
    new_F5433_, new_F5434_, new_F5435_, new_F5436_, new_F5437_, new_F5438_,
    new_F5439_, new_F5440_, new_F5441_, new_F5442_, new_F5443_, new_F5444_,
    new_F5445_, new_F5446_, new_F5447_, new_F5448_, new_F5449_, new_F5450_,
    new_F5451_, new_F5452_, new_F5453_, new_F5454_, new_F5455_, new_F5456_,
    new_F5457_, new_F5458_, new_F5459_, new_F5460_, new_F5461_, new_F5462_,
    new_F5463_, new_F5464_, new_F5465_, new_F5466_, new_F5467_, new_F5468_,
    new_F5469_, new_F5470_, new_F5471_, new_F5472_, new_F5473_, new_F5474_,
    new_F5475_, new_F5476_, new_F5477_, new_F5478_, new_F5479_, new_F5480_,
    new_F5481_, new_F5488_, new_F5489_, new_F5490_, new_F5491_, new_F5492_,
    new_F5493_, new_F5494_, new_F5495_, new_F5496_, new_F5497_, new_F5498_,
    new_F5499_, new_F5500_, new_F5501_, new_F5502_, new_F5503_, new_F5504_,
    new_F5505_, new_F5506_, new_F5507_, new_F5508_, new_F5509_, new_F5510_,
    new_F5511_, new_F5512_, new_F5513_, new_F5514_, new_F5515_, new_F5516_,
    new_F5517_, new_F5518_, new_F5519_, new_F5520_, new_F5521_, new_F5522_,
    new_F5523_, new_F5524_, new_F5525_, new_F5526_, new_F5527_, new_F5528_,
    new_F5529_, new_F5530_, new_F5531_, new_F5532_, new_F5533_, new_F5534_,
    new_F5535_, new_F5536_, new_F5537_, new_F5538_, new_F5539_, new_F5540_,
    new_F5541_, new_F5542_, new_F5543_, new_F5544_, new_F5545_, new_F5546_,
    new_F5547_, new_F5548_, new_F5555_, new_F5556_, new_F5557_, new_F5558_,
    new_F5559_, new_F5560_, new_F5561_, new_F5562_, new_F5563_, new_F5564_,
    new_F5565_, new_F5566_, new_F5567_, new_F5568_, new_F5569_, new_F5570_,
    new_F5571_, new_F5572_, new_F5573_, new_F5574_, new_F5575_, new_F5576_,
    new_F5577_, new_F5578_, new_F5579_, new_F5580_, new_F5581_, new_F5582_,
    new_F5583_, new_F5584_, new_F5585_, new_F5586_, new_F5587_, new_F5588_,
    new_F5589_, new_F5590_, new_F5591_, new_F5592_, new_F5593_, new_F5594_,
    new_F5595_, new_F5596_, new_F5597_, new_F5598_, new_F5599_, new_F5600_,
    new_F5601_, new_F5602_, new_F5603_, new_F5604_, new_F5605_, new_F5606_,
    new_F5607_, new_F5608_, new_F5609_, new_F5610_, new_F5611_, new_F5612_,
    new_F5613_, new_F5614_, new_F5615_, new_F5622_, new_F5623_, new_F5624_,
    new_F5625_, new_F5626_, new_F5627_, new_F5628_, new_F5629_, new_F5630_,
    new_F5631_, new_F5632_, new_F5633_, new_F5634_, new_F5635_, new_F5636_,
    new_F5637_, new_F5638_, new_F5639_, new_F5640_, new_F5641_, new_F5642_,
    new_F5643_, new_F5644_, new_F5645_, new_F5646_, new_F5647_, new_F5648_,
    new_F5649_, new_F5650_, new_F5651_, new_F5652_, new_F5653_, new_F5654_,
    new_F5655_, new_F5656_, new_F5657_, new_F5658_, new_F5659_, new_F5660_,
    new_F5661_, new_F5662_, new_F5663_, new_F5664_, new_F5665_, new_F5666_,
    new_F5667_, new_F5668_, new_F5669_, new_F5670_, new_F5671_, new_F5672_,
    new_F5673_, new_F5674_, new_F5675_, new_F5676_, new_F5677_, new_F5678_,
    new_F5679_, new_F5680_, new_F5681_, new_F5682_, new_F5689_, new_F5690_,
    new_F5691_, new_F5692_, new_F5693_, new_F5694_, new_F5695_, new_F5696_,
    new_F5697_, new_F5698_, new_F5699_, new_F5700_, new_F5701_, new_F5702_,
    new_F5703_, new_F5704_, new_F5705_, new_F5706_, new_F5707_, new_F5708_,
    new_F5709_, new_F5710_, new_F5711_, new_F5712_, new_F5713_, new_F5714_,
    new_F5715_, new_F5716_, new_F5717_, new_F5718_, new_F5719_, new_F5720_,
    new_F5721_, new_F5722_, new_F5723_, new_F5724_, new_F5725_, new_F5726_,
    new_F5727_, new_F5728_, new_F5729_, new_F5730_, new_F5731_, new_F5732_,
    new_F5733_, new_F5734_, new_F5735_, new_F5736_, new_F5737_, new_F5738_,
    new_F5739_, new_F5740_, new_F5741_, new_F5742_, new_F5743_, new_F5744_,
    new_F5745_, new_F5746_, new_F5747_, new_F5748_, new_F5749_, new_F5756_,
    new_F5757_, new_F5758_, new_F5759_, new_F5760_, new_F5761_, new_F5762_,
    new_F5763_, new_F5764_, new_F5765_, new_F5766_, new_F5767_, new_F5768_,
    new_F5769_, new_F5770_, new_F5771_, new_F5772_, new_F5773_, new_F5774_,
    new_F5775_, new_F5776_, new_F5777_, new_F5778_, new_F5779_, new_F5780_,
    new_F5781_, new_F5782_, new_F5783_, new_F5784_, new_F5785_, new_F5786_,
    new_F5787_, new_F5788_, new_F5789_, new_F5790_, new_F5791_, new_F5792_,
    new_F5793_, new_F5794_, new_F5795_, new_F5796_, new_F5797_, new_F5798_,
    new_F5799_, new_F5800_, new_F5801_, new_F5802_, new_F5803_, new_F5804_,
    new_F5805_, new_F5806_, new_F5807_, new_F5808_, new_F5809_, new_F5810_,
    new_F5811_, new_F5812_, new_F5813_, new_F5814_, new_F5815_, new_F5816_,
    new_F5823_, new_F5824_, new_F5825_, new_F5826_, new_F5827_, new_F5828_,
    new_F5829_, new_F5830_, new_F5831_, new_F5832_, new_F5833_, new_F5834_,
    new_F5835_, new_F5836_, new_F5837_, new_F5838_, new_F5839_, new_F5840_,
    new_F5841_, new_F5842_, new_F5843_, new_F5844_, new_F5845_, new_F5846_,
    new_F5847_, new_F5848_, new_F5849_, new_F5850_, new_F5851_, new_F5852_,
    new_F5853_, new_F5854_, new_F5855_, new_F5856_, new_F5857_, new_F5858_,
    new_F5859_, new_F5860_, new_F5861_, new_F5862_, new_F5863_, new_F5864_,
    new_F5865_, new_F5866_, new_F5867_, new_F5868_, new_F5869_, new_F5870_,
    new_F5871_, new_F5872_, new_F5873_, new_F5874_, new_F5875_, new_F5876_,
    new_F5877_, new_F5878_, new_F5879_, new_F5880_, new_F5881_, new_F5882_,
    new_F5883_, new_F5890_, new_F5891_, new_F5892_, new_F5893_, new_F5894_,
    new_F5895_, new_F5896_, new_F5897_, new_F5898_, new_F5899_, new_F5900_,
    new_F5901_, new_F5902_, new_F5903_, new_F5904_, new_F5905_, new_F5906_,
    new_F5907_, new_F5908_, new_F5909_, new_F5910_, new_F5911_, new_F5912_,
    new_F5913_, new_F5914_, new_F5915_, new_F5916_, new_F5917_, new_F5918_,
    new_F5919_, new_F5920_, new_F5921_, new_F5922_, new_F5923_, new_F5924_,
    new_F5925_, new_F5926_, new_F5927_, new_F5928_, new_F5929_, new_F5930_,
    new_F5931_, new_F5932_, new_F5933_, new_F5934_, new_F5935_, new_F5936_,
    new_F5937_, new_F5938_, new_F5939_, new_F5940_, new_F5941_, new_F5942_,
    new_F5943_, new_F5944_, new_F5945_, new_F5946_, new_F5947_, new_F5948_,
    new_F5949_, new_F5950_, new_F5957_, new_F5958_, new_F5959_, new_F5960_,
    new_F5961_, new_F5962_, new_F5963_, new_F5964_, new_F5965_, new_F5966_,
    new_F5967_, new_F5968_, new_F5969_, new_F5970_, new_F5971_, new_F5972_,
    new_F5973_, new_F5974_, new_F5975_, new_F5976_, new_F5977_, new_F5978_,
    new_F5979_, new_F5980_, new_F5981_, new_F5982_, new_F5983_, new_F5984_,
    new_F5985_, new_F5986_, new_F5987_, new_F5988_, new_F5989_, new_F5990_,
    new_F5991_, new_F5992_, new_F5993_, new_F5994_, new_F5995_, new_F5996_,
    new_F5997_, new_F5998_, new_F5999_, new_F6000_, new_F6001_, new_F6002_,
    new_F6003_, new_F6004_, new_F6005_, new_F6006_, new_F6007_, new_F6008_,
    new_F6009_, new_F6010_, new_F6011_, new_F6012_, new_F6013_, new_F6014_,
    new_F6015_, new_F6016_, new_F6017_, new_F6024_, new_F6025_, new_F6026_,
    new_F6027_, new_F6028_, new_F6029_, new_F6030_, new_F6031_, new_F6032_,
    new_F6033_, new_F6034_, new_F6035_, new_F6036_, new_F6037_, new_F6038_,
    new_F6039_, new_F6040_, new_F6041_, new_F6042_, new_F6043_, new_F6044_,
    new_F6045_, new_F6046_, new_F6047_, new_F6048_, new_F6049_, new_F6050_,
    new_F6051_, new_F6052_, new_F6053_, new_F6054_, new_F6055_, new_F6056_,
    new_F6057_, new_F6058_, new_F6059_, new_F6060_, new_F6061_, new_F6062_,
    new_F6063_, new_F6064_, new_F6065_, new_F6066_, new_F6067_, new_F6068_,
    new_F6069_, new_F6070_, new_F6071_, new_F6072_, new_F6073_, new_F6074_,
    new_F6075_, new_F6076_, new_F6077_, new_F6078_, new_F6079_, new_F6080_,
    new_F6081_, new_F6082_, new_F6083_, new_F6084_, new_F6091_, new_F6092_,
    new_F6093_, new_F6094_, new_F6095_, new_F6096_, new_F6097_, new_F6098_,
    new_F6099_, new_F6100_, new_F6101_, new_F6102_, new_F6103_, new_F6104_,
    new_F6105_, new_F6106_, new_F6107_, new_F6108_, new_F6109_, new_F6110_,
    new_F6111_, new_F6112_, new_F6113_, new_F6114_, new_F6115_, new_F6116_,
    new_F6117_, new_F6118_, new_F6119_, new_F6120_, new_F6121_, new_F6122_,
    new_F6123_, new_F6124_, new_F6125_, new_F6126_, new_F6127_, new_F6128_,
    new_F6129_, new_F6130_, new_F6131_, new_F6132_, new_F6133_, new_F6134_,
    new_F6135_, new_F6136_, new_F6137_, new_F6138_, new_F6139_, new_F6140_,
    new_F6141_, new_F6142_, new_F6143_, new_F6144_, new_F6145_, new_F6146_,
    new_F6147_, new_F6148_, new_F6149_, new_F6150_, new_F6151_, new_F6158_,
    new_F6159_, new_F6160_, new_F6161_, new_F6162_, new_F6163_, new_F6164_,
    new_F6165_, new_F6166_, new_F6167_, new_F6168_, new_F6169_, new_F6170_,
    new_F6171_, new_F6172_, new_F6173_, new_F6174_, new_F6175_, new_F6176_,
    new_F6177_, new_F6178_, new_F6179_, new_F6180_, new_F6181_, new_F6182_,
    new_F6183_, new_F6184_, new_F6185_, new_F6186_, new_F6187_, new_F6188_,
    new_F6189_, new_F6190_, new_F6191_, new_F6192_, new_F6193_, new_F6194_,
    new_F6195_, new_F6196_, new_F6197_, new_F6198_, new_F6199_, new_F6200_,
    new_F6201_, new_F6202_, new_F6203_, new_F6204_, new_F6205_, new_F6206_,
    new_F6207_, new_F6208_, new_F6209_, new_F6210_, new_F6211_, new_F6212_,
    new_F6213_, new_F6214_, new_F6215_, new_F6216_, new_F6217_, new_F6218_,
    new_F6225_, new_F6226_, new_F6227_, new_F6228_, new_F6229_, new_F6230_,
    new_F6231_, new_F6232_, new_F6233_, new_F6234_, new_F6235_, new_F6236_,
    new_F6237_, new_F6238_, new_F6239_, new_F6240_, new_F6241_, new_F6242_,
    new_F6243_, new_F6244_, new_F6245_, new_F6246_, new_F6247_, new_F6248_,
    new_F6249_, new_F6250_, new_F6251_, new_F6252_, new_F6253_, new_F6254_,
    new_F6255_, new_F6256_, new_F6257_, new_F6258_, new_F6259_, new_F6260_,
    new_F6261_, new_F6262_, new_F6263_, new_F6264_, new_F6265_, new_F6266_,
    new_F6267_, new_F6268_, new_F6269_, new_F6270_, new_F6271_, new_F6272_,
    new_F6273_, new_F6274_, new_F6275_, new_F6276_, new_F6277_, new_F6278_,
    new_F6279_, new_F6280_, new_F6281_, new_F6282_, new_F6283_, new_F6284_,
    new_F6285_, new_F6292_, new_F6293_, new_F6294_, new_F6295_, new_F6296_,
    new_F6297_, new_F6298_, new_F6299_, new_F6300_, new_F6301_, new_F6302_,
    new_F6303_, new_F6304_, new_F6305_, new_F6306_, new_F6307_, new_F6308_,
    new_F6309_, new_F6310_, new_F6311_, new_F6312_, new_F6313_, new_F6314_,
    new_F6315_, new_F6316_, new_F6317_, new_F6318_, new_F6319_, new_F6320_,
    new_F6321_, new_F6322_, new_F6323_, new_F6324_, new_F6325_, new_F6326_,
    new_F6327_, new_F6328_, new_F6329_, new_F6330_, new_F6331_, new_F6332_,
    new_F6333_, new_F6334_, new_F6335_, new_F6336_, new_F6337_, new_F6338_,
    new_F6339_, new_F6340_, new_F6341_, new_F6342_, new_F6343_, new_F6344_,
    new_F6345_, new_F6346_, new_F6347_, new_F6348_, new_F6349_, new_F6350_,
    new_F6351_, new_F6352_, new_F6359_, new_F6360_, new_F6361_, new_F6362_,
    new_F6363_, new_F6364_, new_F6365_, new_F6366_, new_F6367_, new_F6368_,
    new_F6369_, new_F6370_, new_F6371_, new_F6372_, new_F6373_, new_F6374_,
    new_F6375_, new_F6376_, new_F6377_, new_F6378_, new_F6379_, new_F6380_,
    new_F6381_, new_F6382_, new_F6383_, new_F6384_, new_F6385_, new_F6386_,
    new_F6387_, new_F6388_, new_F6389_, new_F6390_, new_F6391_, new_F6392_,
    new_F6393_, new_F6394_, new_F6395_, new_F6396_, new_F6397_, new_F6398_,
    new_F6399_, new_F6400_, new_F6401_, new_F6402_, new_F6403_, new_F6404_,
    new_F6405_, new_F6406_, new_F6407_, new_F6408_, new_F6409_, new_F6410_,
    new_F6411_, new_F6412_, new_F6413_, new_F6414_, new_F6415_, new_F6416_,
    new_F6417_, new_F6418_, new_F6419_, new_F6426_, new_F6427_, new_F6428_,
    new_F6429_, new_F6430_, new_F6431_, new_F6432_, new_F6433_, new_F6434_,
    new_F6435_, new_F6436_, new_F6437_, new_F6438_, new_F6439_, new_F6440_,
    new_F6441_, new_F6442_, new_F6443_, new_F6444_, new_F6445_, new_F6446_,
    new_F6447_, new_F6448_, new_F6449_, new_F6450_, new_F6451_, new_F6452_,
    new_F6453_, new_F6454_, new_F6455_, new_F6456_, new_F6457_, new_F6458_,
    new_F6459_, new_F6460_, new_F6461_, new_F6462_, new_F6463_, new_F6464_,
    new_F6465_, new_F6466_, new_F6467_, new_F6468_, new_F6469_, new_F6470_,
    new_F6471_, new_F6472_, new_F6473_, new_F6474_, new_F6475_, new_F6476_,
    new_F6477_, new_F6478_, new_F6479_, new_F6480_, new_F6481_, new_F6482_,
    new_F6483_, new_F6484_, new_F6485_, new_F6486_, new_F6493_, new_F6494_,
    new_F6495_, new_F6496_, new_F6497_, new_F6498_, new_F6499_, new_F6500_,
    new_F6501_, new_F6502_, new_F6503_, new_F6504_, new_F6505_, new_F6506_,
    new_F6507_, new_F6508_, new_F6509_, new_F6510_, new_F6511_, new_F6512_,
    new_F6513_, new_F6514_, new_F6515_, new_F6516_, new_F6517_, new_F6518_,
    new_F6519_, new_F6520_, new_F6521_, new_F6522_, new_F6523_, new_F6524_,
    new_F6525_, new_F6526_, new_F6527_, new_F6528_, new_F6529_, new_F6530_,
    new_F6531_, new_F6532_, new_F6533_, new_F6534_, new_F6535_, new_F6536_,
    new_F6537_, new_F6538_, new_F6539_, new_F6540_, new_F6541_, new_F6542_,
    new_F6543_, new_F6544_, new_F6545_, new_F6546_, new_F6547_, new_F6548_,
    new_F6549_, new_F6550_, new_F6551_, new_F6552_, new_F6553_, new_F6560_,
    new_F6561_, new_F6562_, new_F6563_, new_F6564_, new_F6565_, new_F6566_,
    new_F6567_, new_F6568_, new_F6569_, new_F6570_, new_F6571_, new_F6572_,
    new_F6573_, new_F6574_, new_F6575_, new_F6576_, new_F6577_, new_F6578_,
    new_F6579_, new_F6580_, new_F6581_, new_F6582_, new_F6583_, new_F6584_,
    new_F6585_, new_F6586_, new_F6587_, new_F6588_, new_F6589_, new_F6590_,
    new_F6591_, new_F6592_, new_F6593_, new_F6594_, new_F6595_, new_F6596_,
    new_F6597_, new_F6598_, new_F6599_, new_F6600_, new_F6601_, new_F6602_,
    new_F6603_, new_F6604_, new_F6605_, new_F6606_, new_F6607_, new_F6608_,
    new_F6609_, new_F6610_, new_F6611_, new_F6612_, new_F6613_, new_F6614_,
    new_F6615_, new_F6616_, new_F6617_, new_F6618_, new_F6619_, new_F6620_,
    new_F6627_, new_F6628_, new_F6629_, new_F6630_, new_F6631_, new_F6632_,
    new_F6633_, new_F6634_, new_F6635_, new_F6636_, new_F6637_, new_F6638_,
    new_F6639_, new_F6640_, new_F6641_, new_F6642_, new_F6643_, new_F6644_,
    new_F6645_, new_F6646_, new_F6647_, new_F6648_, new_F6649_, new_F6650_,
    new_F6651_, new_F6652_, new_F6653_, new_F6654_, new_F6655_, new_F6656_,
    new_F6657_, new_F6658_, new_F6659_, new_F6660_, new_F6661_, new_F6662_,
    new_F6663_, new_F6664_, new_F6665_, new_F6666_, new_F6667_, new_F6668_,
    new_F6669_, new_F6670_, new_F6671_, new_F6672_, new_F6673_, new_F6674_,
    new_F6675_, new_F6676_, new_F6677_, new_F6678_, new_F6679_, new_F6680_,
    new_F6681_, new_F6682_, new_F6683_, new_F6684_, new_F6685_, new_F6686_,
    new_F6687_, new_F6694_, new_F6695_, new_F6696_, new_F6697_, new_F6698_,
    new_F6699_, new_F6700_, new_F6701_, new_F6702_, new_F6703_, new_F6704_,
    new_F6705_, new_F6706_, new_F6707_, new_F6708_, new_F6709_, new_F6710_,
    new_F6711_, new_F6712_, new_F6713_, new_F6714_, new_F6715_, new_F6716_,
    new_F6717_, new_F6718_, new_F6719_, new_F6720_, new_F6721_, new_F6722_,
    new_F6723_, new_F6724_, new_F6725_, new_F6726_, new_F6727_, new_F6728_,
    new_F6729_, new_F6730_, new_F6731_, new_F6732_, new_F6733_, new_F6734_,
    new_F6735_, new_F6736_, new_F6737_, new_F6738_, new_F6739_, new_F6740_,
    new_F6741_, new_F6742_, new_F6743_, new_F6744_, new_F6745_, new_F6746_,
    new_F6747_, new_F6748_, new_F6749_, new_F6750_, new_F6751_, new_F6752_,
    new_F6753_, new_F6754_, new_F6761_, new_F6762_, new_F6763_, new_F6764_,
    new_F6765_, new_F6766_, new_F6767_, new_F6768_, new_F6769_, new_F6770_,
    new_F6771_, new_F6772_, new_F6773_, new_F6774_, new_F6775_, new_F6776_,
    new_F6777_, new_F6778_, new_F6779_, new_F6780_, new_F6781_, new_F6782_,
    new_F6783_, new_F6784_, new_F6785_, new_F6786_, new_F6787_, new_F6788_,
    new_F6789_, new_F6790_, new_F6791_, new_F6792_, new_F6793_, new_F6794_,
    new_F6795_, new_F6796_, new_F6797_, new_F6798_, new_F6799_, new_F6800_,
    new_F6801_, new_F6802_, new_F6803_, new_F6804_, new_F6805_, new_F6806_,
    new_F6807_, new_F6808_, new_F6809_, new_F6810_, new_F6811_, new_F6812_,
    new_F6813_, new_F6814_, new_F6815_, new_F6816_, new_F6817_, new_F6818_,
    new_F6819_, new_F6820_, new_F6821_, new_F6828_, new_F6829_, new_F6830_,
    new_F6831_, new_F6832_, new_F6833_, new_F6834_, new_F6835_, new_F6836_,
    new_F6837_, new_F6838_, new_F6839_, new_F6840_, new_F6841_, new_F6842_,
    new_F6843_, new_F6844_, new_F6845_, new_F6846_, new_F6847_, new_F6848_,
    new_F6849_, new_F6850_, new_F6851_, new_F6852_, new_F6853_, new_F6854_,
    new_F6855_, new_F6856_, new_F6857_, new_F6858_, new_F6859_, new_F6860_,
    new_F6861_, new_F6862_, new_F6863_, new_F6864_, new_F6865_, new_F6866_,
    new_F6867_, new_F6868_, new_F6869_, new_F6870_, new_F6871_, new_F6872_,
    new_F6873_, new_F6874_, new_F6875_, new_F6876_, new_F6877_, new_F6878_,
    new_F6879_, new_F6880_, new_F6881_, new_F6882_, new_F6883_, new_F6884_,
    new_F6885_, new_F6886_, new_F6887_, new_F6888_, new_F6895_, new_F6896_,
    new_F6897_, new_F6898_, new_F6899_, new_F6900_, new_F6901_, new_F6902_,
    new_F6903_, new_F6904_, new_F6905_, new_F6906_, new_F6907_, new_F6908_,
    new_F6909_, new_F6910_, new_F6911_, new_F6912_, new_F6913_, new_F6914_,
    new_F6915_, new_F6916_, new_F6917_, new_F6918_, new_F6919_, new_F6920_,
    new_F6921_, new_F6922_, new_F6923_, new_F6924_, new_F6925_, new_F6926_,
    new_F6927_, new_F6928_, new_F6929_, new_F6930_, new_F6931_, new_F6932_,
    new_F6933_, new_F6934_, new_F6935_, new_F6936_, new_F6937_, new_F6938_,
    new_F6939_, new_F6940_, new_F6941_, new_F6942_, new_F6943_, new_F6944_,
    new_F6945_, new_F6946_, new_F6947_, new_F6948_, new_F6949_, new_F6950_,
    new_F6951_, new_F6952_, new_F6953_, new_F6954_, new_F6955_, new_F6962_,
    new_F6963_, new_F6964_, new_F6965_, new_F6966_, new_F6967_, new_F6968_,
    new_F6969_, new_F6970_, new_F6971_, new_F6972_, new_F6973_, new_F6974_,
    new_F6975_, new_F6976_, new_F6977_, new_F6978_, new_F6979_, new_F6980_,
    new_F6981_, new_F6982_, new_F6983_, new_F6984_, new_F6985_, new_F6986_,
    new_F6987_, new_F6988_, new_F6989_, new_F6990_, new_F6991_, new_F6992_,
    new_F6993_, new_F6994_, new_F6995_, new_F6996_, new_F6997_, new_F6998_,
    new_F6999_, new_F7000_, new_F7001_, new_F7002_, new_F7003_, new_F7004_,
    new_F7005_, new_F7006_, new_F7007_, new_F7008_, new_F7009_, new_F7010_,
    new_F7011_, new_F7012_, new_F7013_, new_F7014_, new_F7015_, new_F7016_,
    new_F7017_, new_F7018_, new_F7019_, new_F7020_, new_F7021_, new_F7022_,
    new_F7029_, new_F7030_, new_F7031_, new_F7032_, new_F7033_, new_F7034_,
    new_F7035_, new_F7036_, new_F7037_, new_F7038_, new_F7039_, new_F7040_,
    new_F7041_, new_F7042_, new_F7043_, new_F7044_, new_F7045_, new_F7046_,
    new_F7047_, new_F7048_, new_F7049_, new_F7050_, new_F7051_, new_F7052_,
    new_F7053_, new_F7054_, new_F7055_, new_F7056_, new_F7057_, new_F7058_,
    new_F7059_, new_F7060_, new_F7061_, new_F7062_, new_F7063_, new_F7064_,
    new_F7065_, new_F7066_, new_F7067_, new_F7068_, new_F7069_, new_F7070_,
    new_F7071_, new_F7072_, new_F7073_, new_F7074_, new_F7075_, new_F7076_,
    new_F7077_, new_F7078_, new_F7079_, new_F7080_, new_F7081_, new_F7082_,
    new_F7083_, new_F7084_, new_F7085_, new_F7086_, new_F7087_, new_F7088_,
    new_F7089_, new_F7096_, new_F7097_, new_F7098_, new_F7099_, new_F7100_,
    new_F7101_, new_F7102_, new_F7103_, new_F7104_, new_F7105_, new_F7106_,
    new_F7107_, new_F7108_, new_F7109_, new_F7110_, new_F7111_, new_F7112_,
    new_F7113_, new_F7114_, new_F7115_, new_F7116_, new_F7117_, new_F7118_,
    new_F7119_, new_F7120_, new_F7121_, new_F7122_, new_F7123_, new_F7124_,
    new_F7125_, new_F7126_, new_F7127_, new_F7128_, new_F7129_, new_F7130_,
    new_F7131_, new_F7132_, new_F7133_, new_F7134_, new_F7135_, new_F7136_,
    new_F7137_, new_F7138_, new_F7139_, new_F7140_, new_F7141_, new_F7142_,
    new_F7143_, new_F7144_, new_F7145_, new_F7146_, new_F7147_, new_F7148_,
    new_F7149_, new_F7150_, new_F7151_, new_F7152_, new_F7153_, new_F7154_,
    new_F7155_, new_F7156_, new_F7163_, new_F7164_, new_F7165_, new_F7166_,
    new_F7167_, new_F7168_, new_F7169_, new_F7170_, new_F7171_, new_F7172_,
    new_F7173_, new_F7174_, new_F7175_, new_F7176_, new_F7177_, new_F7178_,
    new_F7179_, new_F7180_, new_F7181_, new_F7182_, new_F7183_, new_F7184_,
    new_F7185_, new_F7186_, new_F7187_, new_F7188_, new_F7189_, new_F7190_,
    new_F7191_, new_F7192_, new_F7193_, new_F7194_, new_F7195_, new_F7196_,
    new_F7197_, new_F7198_, new_F7199_, new_F7200_, new_F7201_, new_F7202_,
    new_F7203_, new_F7204_, new_F7205_, new_F7206_, new_F7207_, new_F7208_,
    new_F7209_, new_F7210_, new_F7211_, new_F7212_, new_F7213_, new_F7214_,
    new_F7215_, new_F7216_, new_F7217_, new_F7218_, new_F7219_, new_F7220_,
    new_F7221_, new_F7222_, new_F7223_, new_F7230_, new_F7231_, new_F7232_,
    new_F7233_, new_F7234_, new_F7235_, new_F7236_, new_F7237_, new_F7238_,
    new_F7239_, new_F7240_, new_F7241_, new_F7242_, new_F7243_, new_F7244_,
    new_F7245_, new_F7246_, new_F7247_, new_F7248_, new_F7249_, new_F7250_,
    new_F7251_, new_F7252_, new_F7253_, new_F7254_, new_F7255_, new_F7256_,
    new_F7257_, new_F7258_, new_F7259_, new_F7260_, new_F7261_, new_F7262_,
    new_F7263_, new_F7264_, new_F7265_, new_F7266_, new_F7267_, new_F7268_,
    new_F7269_, new_F7270_, new_F7271_, new_F7272_, new_F7273_, new_F7274_,
    new_F7275_, new_F7276_, new_F7277_, new_F7278_, new_F7279_, new_F7280_,
    new_F7281_, new_F7282_, new_F7283_, new_F7284_, new_F7285_, new_F7286_,
    new_F7287_, new_F7288_, new_F7289_, new_F7290_, new_F7297_, new_F7298_,
    new_F7299_, new_F7300_, new_F7301_, new_F7302_, new_F7303_, new_F7304_,
    new_F7305_, new_F7306_, new_F7307_, new_F7308_, new_F7309_, new_F7310_,
    new_F7311_, new_F7312_, new_F7313_, new_F7314_, new_F7315_, new_F7316_,
    new_F7317_, new_F7318_, new_F7319_, new_F7320_, new_F7321_, new_F7322_,
    new_F7323_, new_F7324_, new_F7325_, new_F7326_, new_F7327_, new_F7328_,
    new_F7329_, new_F7330_, new_F7331_, new_F7332_, new_F7333_, new_F7334_,
    new_F7335_, new_F7336_, new_F7337_, new_F7338_, new_F7339_, new_F7340_,
    new_F7341_, new_F7342_, new_F7343_, new_F7344_, new_F7345_, new_F7346_,
    new_F7347_, new_F7348_, new_F7349_, new_F7350_, new_F7351_, new_F7352_,
    new_F7353_, new_F7354_, new_F7355_, new_F7356_, new_F7357_, new_F7364_,
    new_F7365_, new_F7366_, new_F7367_, new_F7368_, new_F7369_, new_F7370_,
    new_F7371_, new_F7372_, new_F7373_, new_F7374_, new_F7375_, new_F7376_,
    new_F7377_, new_F7378_, new_F7379_, new_F7380_, new_F7381_, new_F7382_,
    new_F7383_, new_F7384_, new_F7385_, new_F7386_, new_F7387_, new_F7388_,
    new_F7389_, new_F7390_, new_F7391_, new_F7392_, new_F7393_, new_F7394_,
    new_F7395_, new_F7396_, new_F7397_, new_F7398_, new_F7399_, new_F7400_,
    new_F7401_, new_F7402_, new_F7403_, new_F7404_, new_F7405_, new_F7406_,
    new_F7407_, new_F7408_, new_F7409_, new_F7410_, new_F7411_, new_F7412_,
    new_F7413_, new_F7414_, new_F7415_, new_F7416_, new_F7417_, new_F7418_,
    new_F7419_, new_F7420_, new_F7421_, new_F7422_, new_F7423_, new_F7424_,
    new_F7431_, new_F7432_, new_F7433_, new_F7434_, new_F7435_, new_F7436_,
    new_F7437_, new_F7438_, new_F7439_, new_F7440_, new_F7441_, new_F7442_,
    new_F7443_, new_F7444_, new_F7445_, new_F7446_, new_F7447_, new_F7448_,
    new_F7449_, new_F7450_, new_F7451_, new_F7452_, new_F7453_, new_F7454_,
    new_F7455_, new_F7456_, new_F7457_, new_F7458_, new_F7459_, new_F7460_,
    new_F7461_, new_F7462_, new_F7463_, new_F7464_, new_F7465_, new_F7466_,
    new_F7467_, new_F7468_, new_F7469_, new_F7470_, new_F7471_, new_F7472_,
    new_F7473_, new_F7474_, new_F7475_, new_F7476_, new_F7477_, new_F7478_,
    new_F7479_, new_F7480_, new_F7481_, new_F7482_, new_F7483_, new_F7484_,
    new_F7485_, new_F7486_, new_F7487_, new_F7488_, new_F7489_, new_F7490_,
    new_F7491_, new_F7498_, new_F7499_, new_F7500_, new_F7501_, new_F7502_,
    new_F7503_, new_F7504_, new_F7505_, new_F7506_, new_F7507_, new_F7508_,
    new_F7509_, new_F7510_, new_F7511_, new_F7512_, new_F7513_, new_F7514_,
    new_F7515_, new_F7516_, new_F7517_, new_F7518_, new_F7519_, new_F7520_,
    new_F7521_, new_F7522_, new_F7523_, new_F7524_, new_F7525_, new_F7526_,
    new_F7527_, new_F7528_, new_F7529_, new_F7530_, new_F7531_, new_F7532_,
    new_F7533_, new_F7534_, new_F7535_, new_F7536_, new_F7537_, new_F7538_,
    new_F7539_, new_F7540_, new_F7541_, new_F7542_, new_F7543_, new_F7544_,
    new_F7545_, new_F7546_, new_F7547_, new_F7548_, new_F7549_, new_F7550_,
    new_F7551_, new_F7552_, new_F7553_, new_F7554_, new_F7555_, new_F7556_,
    new_F7557_, new_F7558_, new_F7565_, new_F7566_, new_F7567_, new_F7568_,
    new_F7569_, new_F7570_, new_F7571_, new_F7572_, new_F7573_, new_F7574_,
    new_F7575_, new_F7576_, new_F7577_, new_F7578_, new_F7579_, new_F7580_,
    new_F7581_, new_F7582_, new_F7583_, new_F7584_, new_F7585_, new_F7586_,
    new_F7587_, new_F7588_, new_F7589_, new_F7590_, new_F7591_, new_F7592_,
    new_F7593_, new_F7594_, new_F7595_, new_F7596_, new_F7597_, new_F7598_,
    new_F7599_, new_F7600_, new_F7601_, new_F7602_, new_F7603_, new_F7604_,
    new_F7605_, new_F7606_, new_F7607_, new_F7608_, new_F7609_, new_F7610_,
    new_F7611_, new_F7612_, new_F7613_, new_F7614_, new_F7615_, new_F7616_,
    new_F7617_, new_F7618_, new_F7619_, new_F7620_, new_F7621_, new_F7622_,
    new_F7623_, new_F7624_, new_F7625_, new_F7632_, new_F7633_, new_F7634_,
    new_F7635_, new_F7636_, new_F7637_, new_F7638_, new_F7639_, new_F7640_,
    new_F7641_, new_F7642_, new_F7643_, new_F7644_, new_F7645_, new_F7646_,
    new_F7647_, new_F7648_, new_F7649_, new_F7650_, new_F7651_, new_F7652_,
    new_F7653_, new_F7654_, new_F7655_, new_F7656_, new_F7657_, new_F7658_,
    new_F7659_, new_F7660_, new_F7661_, new_F7662_, new_F7663_, new_F7664_,
    new_F7665_, new_F7666_, new_F7667_, new_F7668_, new_F7669_, new_F7670_,
    new_F7671_, new_F7672_, new_F7673_, new_F7674_, new_F7675_, new_F7676_,
    new_F7677_, new_F7678_, new_F7679_, new_F7680_, new_F7681_, new_F7682_,
    new_F7683_, new_F7684_, new_F7685_, new_F7686_, new_F7687_, new_F7688_,
    new_F7689_, new_F7690_, new_F7691_, new_F7692_, new_F7699_, new_F7700_,
    new_F7701_, new_F7702_, new_F7703_, new_F7704_, new_F7705_, new_F7706_,
    new_F7707_, new_F7708_, new_F7709_, new_F7710_, new_F7711_, new_F7712_,
    new_F7713_, new_F7714_, new_F7715_, new_F7716_, new_F7717_, new_F7718_,
    new_F7719_, new_F7720_, new_F7721_, new_F7722_, new_F7723_, new_F7724_,
    new_F7725_, new_F7726_, new_F7727_, new_F7728_, new_F7729_, new_F7730_,
    new_F7731_, new_F7732_, new_F7733_, new_F7734_, new_F7735_, new_F7736_,
    new_F7737_, new_F7738_, new_F7739_, new_F7740_, new_F7741_, new_F7742_,
    new_F7743_, new_F7744_, new_F7745_, new_F7746_, new_F7747_, new_F7748_,
    new_F7749_, new_F7750_, new_F7751_, new_F7752_, new_F7753_, new_F7754_,
    new_F7755_, new_F7756_, new_F7757_, new_F7758_, new_F7759_, new_F7766_,
    new_F7767_, new_F7768_, new_F7769_, new_F7770_, new_F7771_, new_F7772_,
    new_F7773_, new_F7774_, new_F7775_, new_F7776_, new_F7777_, new_F7778_,
    new_F7779_, new_F7780_, new_F7781_, new_F7782_, new_F7783_, new_F7784_,
    new_F7785_, new_F7786_, new_F7787_, new_F7788_, new_F7789_, new_F7790_,
    new_F7791_, new_F7792_, new_F7793_, new_F7794_, new_F7795_, new_F7796_,
    new_F7797_, new_F7798_, new_F7799_, new_F7800_, new_F7801_, new_F7802_,
    new_F7803_, new_F7804_, new_F7805_, new_F7806_, new_F7807_, new_F7808_,
    new_F7809_, new_F7810_, new_F7811_, new_F7812_, new_F7813_, new_F7814_,
    new_F7815_, new_F7816_, new_F7817_, new_F7818_, new_F7819_, new_F7820_,
    new_F7821_, new_F7822_, new_F7823_, new_F7824_, new_F7825_, new_F7826_,
    new_F7833_, new_F7834_, new_F7835_, new_F7836_, new_F7837_, new_F7838_,
    new_F7839_, new_F7840_, new_F7841_, new_F7842_, new_F7843_, new_F7844_,
    new_F7845_, new_F7846_, new_F7847_, new_F7848_, new_F7849_, new_F7850_,
    new_F7851_, new_F7852_, new_F7853_, new_F7854_, new_F7855_, new_F7856_,
    new_F7857_, new_F7858_, new_F7859_, new_F7860_, new_F7861_, new_F7862_,
    new_F7863_, new_F7864_, new_F7865_, new_F7866_, new_F7867_, new_F7868_,
    new_F7869_, new_F7870_, new_F7871_, new_F7872_, new_F7873_, new_F7874_,
    new_F7875_, new_F7876_, new_F7877_, new_F7878_, new_F7879_, new_F7880_,
    new_F7881_, new_F7882_, new_F7883_, new_F7884_, new_F7885_, new_F7886_,
    new_F7887_, new_F7888_, new_F7889_, new_F7890_, new_F7891_, new_F7892_,
    new_F7893_, new_F7900_, new_F7901_, new_F7902_, new_F7903_, new_F7904_,
    new_F7905_, new_F7906_, new_F7907_, new_F7908_, new_F7909_, new_F7910_,
    new_F7911_, new_F7912_, new_F7913_, new_F7914_, new_F7915_, new_F7916_,
    new_F7917_, new_F7918_, new_F7919_, new_F7920_, new_F7921_, new_F7922_,
    new_F7923_, new_F7924_, new_F7925_, new_F7926_, new_F7927_, new_F7928_,
    new_F7929_, new_F7930_, new_F7931_, new_F7932_, new_F7933_, new_F7934_,
    new_F7935_, new_F7936_, new_F7937_, new_F7938_, new_F7939_, new_F7940_,
    new_F7941_, new_F7942_, new_F7943_, new_F7944_, new_F7945_, new_F7946_,
    new_F7947_, new_F7948_, new_F7949_, new_F7950_, new_F7951_, new_F7952_,
    new_F7953_, new_F7954_, new_F7955_, new_F7956_, new_F7957_, new_F7958_,
    new_F7959_, new_F7960_, new_F7967_, new_F7968_, new_F7969_, new_F7970_,
    new_F7971_, new_F7972_, new_F7973_, new_F7974_, new_F7975_, new_F7976_,
    new_F7977_, new_F7978_, new_F7979_, new_F7980_, new_F7981_, new_F7982_,
    new_F7983_, new_F7984_, new_F7985_, new_F7986_, new_F7987_, new_F7988_,
    new_F7989_, new_F7990_, new_F7991_, new_F7992_, new_F7993_, new_F7994_,
    new_F7995_, new_F7996_, new_F7997_, new_F7998_, new_F7999_, new_F8000_,
    new_F8001_, new_F8002_, new_F8003_, new_F8004_, new_F8005_, new_F8006_,
    new_F8007_, new_F8008_, new_F8009_, new_F8010_, new_F8011_, new_F8012_,
    new_F8013_, new_F8014_, new_F8015_, new_F8016_, new_F8017_, new_F8018_,
    new_F8019_, new_F8020_, new_F8021_, new_F8022_, new_F8023_, new_F8024_,
    new_F8025_, new_F8026_, new_F8027_, new_F8034_, new_F8035_, new_F8036_,
    new_F8037_, new_F8038_, new_F8039_, new_F8040_, new_F8041_, new_F8042_,
    new_F8043_, new_F8044_, new_F8045_, new_F8046_, new_F8047_, new_F8048_,
    new_F8049_, new_F8050_, new_F8051_, new_F8052_, new_F8053_, new_F8054_,
    new_F8055_, new_F8056_, new_F8057_, new_F8058_, new_F8059_, new_F8060_,
    new_F8061_, new_F8062_, new_F8063_, new_F8064_, new_F8065_, new_F8066_,
    new_F8067_, new_F8068_, new_F8069_, new_F8070_, new_F8071_, new_F8072_,
    new_F8073_, new_F8074_, new_F8075_, new_F8076_, new_F8077_, new_F8078_,
    new_F8079_, new_F8080_, new_F8081_, new_F8082_, new_F8083_, new_F8084_,
    new_F8085_, new_F8086_, new_F8087_, new_F8088_, new_F8089_, new_F8090_,
    new_F8091_, new_F8092_, new_F8093_, new_F8094_, new_F8101_, new_F8102_,
    new_F8103_, new_F8104_, new_F8105_, new_F8106_, new_F8107_, new_F8108_,
    new_F8109_, new_F8110_, new_F8111_, new_F8112_, new_F8113_, new_F8114_,
    new_F8115_, new_F8116_, new_F8117_, new_F8118_, new_F8119_, new_F8120_,
    new_F8121_, new_F8122_, new_F8123_, new_F8124_, new_F8125_, new_F8126_,
    new_F8127_, new_F8128_, new_F8129_, new_F8130_, new_F8131_, new_F8132_,
    new_F8133_, new_F8134_, new_F8135_, new_F8136_, new_F8137_, new_F8138_,
    new_F8139_, new_F8140_, new_F8141_, new_F8142_, new_F8143_, new_F8144_,
    new_F8145_, new_F8146_, new_F8147_, new_F8148_, new_F8149_, new_F8150_,
    new_F8151_, new_F8152_, new_F8153_, new_F8154_, new_F8155_, new_F8156_,
    new_F8157_, new_F8158_, new_F8159_, new_F8160_, new_F8161_, new_F8168_,
    new_F8169_, new_F8170_, new_F8171_, new_F8172_, new_F8173_, new_F8174_,
    new_F8175_, new_F8176_, new_F8177_, new_F8178_, new_F8179_, new_F8180_,
    new_F8181_, new_F8182_, new_F8183_, new_F8184_, new_F8185_, new_F8186_,
    new_F8187_, new_F8188_, new_F8189_, new_F8190_, new_F8191_, new_F8192_,
    new_F8193_, new_F8194_, new_F8195_, new_F8196_, new_F8197_, new_F8198_,
    new_F8199_, new_F8200_, new_F8201_, new_F8202_, new_F8203_, new_F8204_,
    new_F8205_, new_F8206_, new_F8207_, new_F8208_, new_F8209_, new_F8210_,
    new_F8211_, new_F8212_, new_F8213_, new_F8214_, new_F8215_, new_F8216_,
    new_F8217_, new_F8218_, new_F8219_, new_F8220_, new_F8221_, new_F8222_,
    new_F8223_, new_F8224_, new_F8225_, new_F8226_, new_F8227_, new_F8228_,
    new_F8235_, new_F8236_, new_F8237_, new_F8238_, new_F8239_, new_F8240_,
    new_F8241_, new_F8242_, new_F8243_, new_F8244_, new_F8245_, new_F8246_,
    new_F8247_, new_F8248_, new_F8249_, new_F8250_, new_F8251_, new_F8252_,
    new_F8253_, new_F8254_, new_F8255_, new_F8256_, new_F8257_, new_F8258_,
    new_F8259_, new_F8260_, new_F8261_, new_F8262_, new_F8263_, new_F8264_,
    new_F8265_, new_F8266_, new_F8267_, new_F8268_, new_F8269_, new_F8270_,
    new_F8271_, new_F8272_, new_F8273_, new_F8274_, new_F8275_, new_F8276_,
    new_F8277_, new_F8278_, new_F8279_, new_F8280_, new_F8281_, new_F8282_,
    new_F8283_, new_F8284_, new_F8285_, new_F8286_, new_F8287_, new_F8288_,
    new_F8289_, new_F8290_, new_F8291_, new_F8292_, new_F8293_, new_F8294_,
    new_F8295_, new_F8302_, new_F8303_, new_F8304_, new_F8305_, new_F8306_,
    new_F8307_, new_F8308_, new_F8309_, new_F8310_, new_F8311_, new_F8312_,
    new_F8313_, new_F8314_, new_F8315_, new_F8316_, new_F8317_, new_F8318_,
    new_F8319_, new_F8320_, new_F8321_, new_F8322_, new_F8323_, new_F8324_,
    new_F8325_, new_F8326_, new_F8327_, new_F8328_, new_F8329_, new_F8330_,
    new_F8331_, new_F8332_, new_F8333_, new_F8334_, new_F8335_, new_F8336_,
    new_F8337_, new_F8338_, new_F8339_, new_F8340_, new_F8341_, new_F8342_,
    new_F8343_, new_F8344_, new_F8345_, new_F8346_, new_F8347_, new_F8348_,
    new_F8349_, new_F8350_, new_F8351_, new_F8352_, new_F8353_, new_F8354_,
    new_F8355_, new_F8356_, new_F8357_, new_F8358_, new_F8359_, new_F8360_,
    new_F8361_, new_F8362_, new_F8369_, new_F8370_, new_F8371_, new_F8372_,
    new_F8373_, new_F8374_, new_F8375_, new_F8376_, new_F8377_, new_F8378_,
    new_F8379_, new_F8380_, new_F8381_, new_F8382_, new_F8383_, new_F8384_,
    new_F8385_, new_F8386_, new_F8387_, new_F8388_, new_F8389_, new_F8390_,
    new_F8391_, new_F8392_, new_F8393_, new_F8394_, new_F8395_, new_F8396_,
    new_F8397_, new_F8398_, new_F8399_, new_F8400_, new_F8401_, new_F8402_,
    new_F8403_, new_F8404_, new_F8405_, new_F8406_, new_F8407_, new_F8408_,
    new_F8409_, new_F8410_, new_F8411_, new_F8412_, new_F8413_, new_F8414_,
    new_F8415_, new_F8416_, new_F8417_, new_F8418_, new_F8419_, new_F8420_,
    new_F8421_, new_F8422_, new_F8423_, new_F8424_, new_F8425_, new_F8426_,
    new_F8427_, new_F8428_, new_F8429_, new_F8436_, new_F8437_, new_F8438_,
    new_F8439_, new_F8440_, new_F8441_, new_F8442_, new_F8443_, new_F8444_,
    new_F8445_, new_F8446_, new_F8447_, new_F8448_, new_F8449_, new_F8450_,
    new_F8451_, new_F8452_, new_F8453_, new_F8454_, new_F8455_, new_F8456_,
    new_F8457_, new_F8458_, new_F8459_, new_F8460_, new_F8461_, new_F8462_,
    new_F8463_, new_F8464_, new_F8465_, new_F8466_, new_F8467_, new_F8468_,
    new_F8469_, new_F8470_, new_F8471_, new_F8472_, new_F8473_, new_F8474_,
    new_F8475_, new_F8476_, new_F8477_, new_F8478_, new_F8479_, new_F8480_,
    new_F8481_, new_F8482_, new_F8483_, new_F8484_, new_F8485_, new_F8486_,
    new_F8487_, new_F8488_, new_F8489_, new_F8490_, new_F8491_, new_F8492_,
    new_F8493_, new_F8494_, new_F8495_, new_F8496_, new_F8503_, new_F8504_,
    new_F8505_, new_F8506_, new_F8507_, new_F8508_, new_F8509_, new_F8510_,
    new_F8511_, new_F8512_, new_F8513_, new_F8514_, new_F8515_, new_F8516_,
    new_F8517_, new_F8518_, new_F8519_, new_F8520_, new_F8521_, new_F8522_,
    new_F8523_, new_F8524_, new_F8525_, new_F8526_, new_F8527_, new_F8528_,
    new_F8529_, new_F8530_, new_F8531_, new_F8532_, new_F8533_, new_F8534_,
    new_F8535_, new_F8536_, new_F8537_, new_F8538_, new_F8539_, new_F8540_,
    new_F8541_, new_F8542_, new_F8543_, new_F8544_, new_F8545_, new_F8546_,
    new_F8547_, new_F8548_, new_F8549_, new_F8550_, new_F8551_, new_F8552_,
    new_F8553_, new_F8554_, new_F8555_, new_F8556_, new_F8557_, new_F8558_,
    new_F8559_, new_F8560_, new_F8561_, new_F8562_, new_F8563_, new_F8570_,
    new_F8571_, new_F8572_, new_F8573_, new_F8574_, new_F8575_, new_F8576_,
    new_F8577_, new_F8578_, new_F8579_, new_F8580_, new_F8581_, new_F8582_,
    new_F8583_, new_F8584_, new_F8585_, new_F8586_, new_F8587_, new_F8588_,
    new_F8589_, new_F8590_, new_F8591_, new_F8592_, new_F8593_, new_F8594_,
    new_F8595_, new_F8596_, new_F8597_, new_F8598_, new_F8599_, new_F8600_,
    new_F8601_, new_F8602_, new_F8603_, new_F8604_, new_F8605_, new_F8606_,
    new_F8607_, new_F8608_, new_F8609_, new_F8610_, new_F8611_, new_F8612_,
    new_F8613_, new_F8614_, new_F8615_, new_F8616_, new_F8617_, new_F8618_,
    new_F8619_, new_F8620_, new_F8621_, new_F8622_, new_F8623_, new_F8624_,
    new_F8625_, new_F8626_, new_F8627_, new_F8628_, new_F8629_, new_F8630_,
    new_F8637_, new_F8638_, new_F8639_, new_F8640_, new_F8641_, new_F8642_,
    new_F8643_, new_F8644_, new_F8645_, new_F8646_, new_F8647_, new_F8648_,
    new_F8649_, new_F8650_, new_F8651_, new_F8652_, new_F8653_, new_F8654_,
    new_F8655_, new_F8656_, new_F8657_, new_F8658_, new_F8659_, new_F8660_,
    new_F8661_, new_F8662_, new_F8663_, new_F8664_, new_F8665_, new_F8666_,
    new_F8667_, new_F8668_, new_F8669_, new_F8670_, new_F8671_, new_F8672_,
    new_F8673_, new_F8674_, new_F8675_, new_F8676_, new_F8677_, new_F8678_,
    new_F8679_, new_F8680_, new_F8681_, new_F8682_, new_F8683_, new_F8684_,
    new_F8685_, new_F8686_, new_F8687_, new_F8688_, new_F8689_, new_F8690_,
    new_F8691_, new_F8692_, new_F8693_, new_F8694_, new_F8695_, new_F8696_,
    new_F8697_, new_F8704_, new_F8705_, new_F8706_, new_F8707_, new_F8708_,
    new_F8709_, new_F8710_, new_F8711_, new_F8712_, new_F8713_, new_F8714_,
    new_F8715_, new_F8716_, new_F8717_, new_F8718_, new_F8719_, new_F8720_,
    new_F8721_, new_F8722_, new_F8723_, new_F8724_, new_F8725_, new_F8726_,
    new_F8727_, new_F8728_, new_F8729_, new_F8730_, new_F8731_, new_F8732_,
    new_F8733_, new_F8734_, new_F8735_, new_F8736_, new_F8737_, new_F8738_,
    new_F8739_, new_F8740_, new_F8741_, new_F8742_, new_F8743_, new_F8744_,
    new_F8745_, new_F8746_, new_F8747_, new_F8748_, new_F8749_, new_F8750_,
    new_F8751_, new_F8752_, new_F8753_, new_F8754_, new_F8755_, new_F8756_,
    new_F8757_, new_F8758_, new_F8759_, new_F8760_, new_F8761_, new_F8762_,
    new_F8763_, new_F8764_, new_F8771_, new_F8772_, new_F8773_, new_F8774_,
    new_F8775_, new_F8776_, new_F8777_, new_F8778_, new_F8779_, new_F8780_,
    new_F8781_, new_F8782_, new_F8783_, new_F8784_, new_F8785_, new_F8786_,
    new_F8787_, new_F8788_, new_F8789_, new_F8790_, new_F8791_, new_F8792_,
    new_F8793_, new_F8794_, new_F8795_, new_F8796_, new_F8797_, new_F8798_,
    new_F8799_, new_F8800_, new_F8801_, new_F8802_, new_F8803_, new_F8804_,
    new_F8805_, new_F8806_, new_F8807_, new_F8808_, new_F8809_, new_F8810_,
    new_F8811_, new_F8812_, new_F8813_, new_F8814_, new_F8815_, new_F8816_,
    new_F8817_, new_F8818_, new_F8819_, new_F8820_, new_F8821_, new_F8822_,
    new_F8823_, new_F8824_, new_F8825_, new_F8826_, new_F8827_, new_F8828_,
    new_F8829_, new_F8830_, new_F8831_, new_F8838_, new_F8839_, new_F8840_,
    new_F8841_, new_F8842_, new_F8843_, new_F8844_, new_F8845_, new_F8846_,
    new_F8847_, new_F8848_, new_F8849_, new_F8850_, new_F8851_, new_F8852_,
    new_F8853_, new_F8854_, new_F8855_, new_F8856_, new_F8857_, new_F8858_,
    new_F8859_, new_F8860_, new_F8861_, new_F8862_, new_F8863_, new_F8864_,
    new_F8865_, new_F8866_, new_F8867_, new_F8868_, new_F8869_, new_F8870_,
    new_F8871_, new_F8872_, new_F8873_, new_F8874_, new_F8875_, new_F8876_,
    new_F8877_, new_F8878_, new_F8879_, new_F8880_, new_F8881_, new_F8882_,
    new_F8883_, new_F8884_, new_F8885_, new_F8886_, new_F8887_, new_F8888_,
    new_F8889_, new_F8890_, new_F8891_, new_F8892_, new_F8893_, new_F8894_,
    new_F8895_, new_F8896_, new_F8897_, new_F8898_, new_F8905_, new_F8906_,
    new_F8907_, new_F8908_, new_F8909_, new_F8910_, new_F8911_, new_F8912_,
    new_F8913_, new_F8914_, new_F8915_, new_F8916_, new_F8917_, new_F8918_,
    new_F8919_, new_F8920_, new_F8921_, new_F8922_, new_F8923_, new_F8924_,
    new_F8925_, new_F8926_, new_F8927_, new_F8928_, new_F8929_, new_F8930_,
    new_F8931_, new_F8932_, new_F8933_, new_F8934_, new_F8935_, new_F8936_,
    new_F8937_, new_F8938_, new_F8939_, new_F8940_, new_F8941_, new_F8942_,
    new_F8943_, new_F8944_, new_F8945_, new_F8946_, new_F8947_, new_F8948_,
    new_F8949_, new_F8950_, new_F8951_, new_F8952_, new_F8953_, new_F8954_,
    new_F8955_, new_F8956_, new_F8957_, new_F8958_, new_F8959_, new_F8960_,
    new_F8961_, new_F8962_, new_F8963_, new_F8964_, new_F8965_, new_F8972_,
    new_F8973_, new_F8974_, new_F8975_, new_F8976_, new_F8977_, new_F8978_,
    new_F8979_, new_F8980_, new_F8981_, new_F8982_, new_F8983_, new_F8984_,
    new_F8985_, new_F8986_, new_F8987_, new_F8988_, new_F8989_, new_F8990_,
    new_F8991_, new_F8992_, new_F8993_, new_F8994_, new_F8995_, new_F8996_,
    new_F8997_, new_F8998_, new_F8999_, new_F9000_, new_F9001_, new_F9002_,
    new_F9003_, new_F9004_, new_F9005_, new_F9006_, new_F9007_, new_F9008_,
    new_F9009_, new_F9010_, new_F9011_, new_F9012_, new_F9013_, new_F9014_,
    new_F9015_, new_F9016_, new_F9017_, new_F9018_, new_F9019_, new_F9020_,
    new_F9021_, new_F9022_, new_F9023_, new_F9024_, new_F9025_, new_F9026_,
    new_F9027_, new_F9028_, new_F9029_, new_F9030_, new_F9031_, new_F9032_,
    new_F9039_, new_F9040_, new_F9041_, new_F9042_, new_F9043_, new_F9044_,
    new_F9045_, new_F9046_, new_F9047_, new_F9048_, new_F9049_, new_F9050_,
    new_F9051_, new_F9052_, new_F9053_, new_F9054_, new_F9055_, new_F9056_,
    new_F9057_, new_F9058_, new_F9059_, new_F9060_, new_F9061_, new_F9062_,
    new_F9063_, new_F9064_, new_F9065_, new_F9066_, new_F9067_, new_F9068_,
    new_F9069_, new_F9070_, new_F9071_, new_F9072_, new_F9073_, new_F9074_,
    new_F9075_, new_F9076_, new_F9077_, new_F9078_, new_F9079_, new_F9080_,
    new_F9081_, new_F9082_, new_F9083_, new_F9084_, new_F9085_, new_F9086_,
    new_F9087_, new_F9088_, new_F9089_, new_F9090_, new_F9091_, new_F9092_,
    new_F9093_, new_F9094_, new_F9095_, new_F9096_, new_F9097_, new_F9098_,
    new_F9099_, new_F9106_, new_F9107_, new_F9108_, new_F9109_, new_F9110_,
    new_F9111_, new_F9112_, new_F9113_, new_F9114_, new_F9115_, new_F9116_,
    new_F9117_, new_F9118_, new_F9119_, new_F9120_, new_F9121_, new_F9122_,
    new_F9123_, new_F9124_, new_F9125_, new_F9126_, new_F9127_, new_F9128_,
    new_F9129_, new_F9130_, new_F9131_, new_F9132_, new_F9133_, new_F9134_,
    new_F9135_, new_F9136_, new_F9137_, new_F9138_, new_F9139_, new_F9140_,
    new_F9141_, new_F9142_, new_F9143_, new_F9144_, new_F9145_, new_F9146_,
    new_F9147_, new_F9148_, new_F9149_, new_F9150_, new_F9151_, new_F9152_,
    new_F9153_, new_F9154_, new_F9155_, new_F9156_, new_F9157_, new_F9158_,
    new_F9159_, new_F9160_, new_F9161_, new_F9162_, new_F9163_, new_F9164_,
    new_F9165_, new_F9166_, new_F9173_, new_F9174_, new_F9175_, new_F9176_,
    new_F9177_, new_F9178_, new_F9179_, new_F9180_, new_F9181_, new_F9182_,
    new_F9183_, new_F9184_, new_F9185_, new_F9186_, new_F9187_, new_F9188_,
    new_F9189_, new_F9190_, new_F9191_, new_F9192_, new_F9193_, new_F9194_,
    new_F9195_, new_F9196_, new_F9197_, new_F9198_, new_F9199_, new_F9200_,
    new_F9201_, new_F9202_, new_F9203_, new_F9204_, new_F9205_, new_F9206_,
    new_F9207_, new_F9208_, new_F9209_, new_F9210_, new_F9211_, new_F9212_,
    new_F9213_, new_F9214_, new_F9215_, new_F9216_, new_F9217_, new_F9218_,
    new_F9219_, new_F9220_, new_F9221_, new_F9222_, new_F9223_, new_F9224_,
    new_F9225_, new_F9226_, new_F9227_, new_F9228_, new_F9229_, new_F9230_,
    new_F9231_, new_F9232_, new_F9233_, new_F9240_, new_F9241_, new_F9242_,
    new_F9243_, new_F9244_, new_F9245_, new_F9246_, new_F9247_, new_F9248_,
    new_F9249_, new_F9250_, new_F9251_, new_F9252_, new_F9253_, new_F9254_,
    new_F9255_, new_F9256_, new_F9257_, new_F9258_, new_F9259_, new_F9260_,
    new_F9261_, new_F9262_, new_F9263_, new_F9264_, new_F9265_, new_F9266_,
    new_F9267_, new_F9268_, new_F9269_, new_F9270_, new_F9271_, new_F9272_,
    new_F9273_, new_F9274_, new_F9275_, new_F9276_, new_F9277_, new_F9278_,
    new_F9279_, new_F9280_, new_F9281_, new_F9282_, new_F9283_, new_F9284_,
    new_F9285_, new_F9286_, new_F9287_, new_F9288_, new_F9289_, new_F9290_,
    new_F9291_, new_F9292_, new_F9293_, new_F9294_, new_F9295_, new_F9296_,
    new_F9297_, new_F9298_, new_F9299_, new_F9300_, new_F9307_, new_F9308_,
    new_F9309_, new_F9310_, new_F9311_, new_F9312_, new_F9313_, new_F9314_,
    new_F9315_, new_F9316_, new_F9317_, new_F9318_, new_F9319_, new_F9320_,
    new_F9321_, new_F9322_, new_F9323_, new_F9324_, new_F9325_, new_F9326_,
    new_F9327_, new_F9328_, new_F9329_, new_F9330_, new_F9331_, new_F9332_,
    new_F9333_, new_F9334_, new_F9335_, new_F9336_, new_F9337_, new_F9338_,
    new_F9339_, new_F9340_, new_F9341_, new_F9342_, new_F9343_, new_F9344_,
    new_F9345_, new_F9346_, new_F9347_, new_F9348_, new_F9349_, new_F9350_,
    new_F9351_, new_F9352_, new_F9353_, new_F9354_, new_F9355_, new_F9356_,
    new_F9357_, new_F9358_, new_F9359_, new_F9360_, new_F9361_, new_F9362_,
    new_F9363_, new_F9364_, new_F9365_, new_F9366_, new_F9367_, new_F9374_,
    new_F9375_, new_F9376_, new_F9377_, new_F9378_, new_F9379_, new_F9380_,
    new_F9381_, new_F9382_, new_F9383_, new_F9384_, new_F9385_, new_F9386_,
    new_F9387_, new_F9388_, new_F9389_, new_F9390_, new_F9391_, new_F9392_,
    new_F9393_, new_F9394_, new_F9395_, new_F9396_, new_F9397_, new_F9398_,
    new_F9399_, new_F9400_, new_F9401_, new_F9402_, new_F9403_, new_F9404_,
    new_F9405_, new_F9406_, new_F9407_, new_F9408_, new_F9409_, new_F9410_,
    new_F9411_, new_F9412_, new_F9413_, new_F9414_, new_F9415_, new_F9416_,
    new_F9417_, new_F9418_, new_F9419_, new_F9420_, new_F9421_, new_F9422_,
    new_F9423_, new_F9424_, new_F9425_, new_F9426_, new_F9427_, new_F9428_,
    new_F9429_, new_F9430_, new_F9431_, new_F9432_, new_F9433_, new_F9434_,
    new_F9441_, new_F9442_, new_F9443_, new_F9444_, new_F9445_, new_F9446_,
    new_F9447_, new_F9448_, new_F9449_, new_F9450_, new_F9451_, new_F9452_,
    new_F9453_, new_F9454_, new_F9455_, new_F9456_, new_F9457_, new_F9458_,
    new_F9459_, new_F9460_, new_F9461_, new_F9462_, new_F9463_, new_F9464_,
    new_F9465_, new_F9466_, new_F9467_, new_F9468_, new_F9469_, new_F9470_,
    new_F9471_, new_F9472_, new_F9473_, new_F9474_, new_F9475_, new_F9476_,
    new_F9477_, new_F9478_, new_F9479_, new_F9480_, new_F9481_, new_F9482_,
    new_F9483_, new_F9484_, new_F9485_, new_F9486_, new_F9487_, new_F9488_,
    new_F9489_, new_F9490_, new_F9491_, new_F9492_, new_F9493_, new_F9494_,
    new_F9495_, new_F9496_, new_F9497_, new_F9498_, new_F9499_, new_F9500_,
    new_F9501_, new_F9508_, new_F9509_, new_F9510_, new_F9511_, new_F9512_,
    new_F9513_, new_F9514_, new_F9515_, new_F9516_, new_F9517_, new_F9518_,
    new_F9519_, new_F9520_, new_F9521_, new_F9522_, new_F9523_, new_F9524_,
    new_F9525_, new_F9526_, new_F9527_, new_F9528_, new_F9529_, new_F9530_,
    new_F9531_, new_F9532_, new_F9533_, new_F9534_, new_F9535_, new_F9536_,
    new_F9537_, new_F9538_, new_F9539_, new_F9540_, new_F9541_, new_F9542_,
    new_F9543_, new_F9544_, new_F9545_, new_F9546_, new_F9547_, new_F9548_,
    new_F9549_, new_F9550_, new_F9551_, new_F9552_, new_F9553_, new_F9554_,
    new_F9555_, new_F9556_, new_F9557_, new_F9558_, new_F9559_, new_F9560_,
    new_F9561_, new_F9562_, new_F9563_, new_F9564_, new_F9565_, new_F9566_,
    new_F9567_, new_F9568_, new_F9575_, new_F9576_, new_F9577_, new_F9578_,
    new_F9579_, new_F9580_, new_F9581_, new_F9582_, new_F9583_, new_F9584_,
    new_F9585_, new_F9586_, new_F9587_, new_F9588_, new_F9589_, new_F9590_,
    new_F9591_, new_F9592_, new_F9593_, new_F9594_, new_F9595_, new_F9596_,
    new_F9597_, new_F9598_, new_F9599_, new_F9600_, new_F9601_, new_F9602_,
    new_F9603_, new_F9604_, new_F9605_, new_F9606_, new_F9607_, new_F9608_,
    new_F9609_, new_F9610_, new_F9611_, new_F9612_, new_F9613_, new_F9614_,
    new_F9615_, new_F9616_, new_F9617_, new_F9618_, new_F9619_, new_F9620_,
    new_F9621_, new_F9622_, new_F9623_, new_F9624_, new_F9625_, new_F9626_,
    new_F9627_, new_F9628_, new_F9629_, new_F9630_, new_F9631_, new_F9632_,
    new_F9633_, new_F9634_, new_F9635_, new_F9642_, new_F9643_, new_F9644_,
    new_F9645_, new_F9646_, new_F9647_, new_F9648_, new_F9649_, new_F9650_,
    new_F9651_, new_F9652_, new_F9653_, new_F9654_, new_F9655_, new_F9656_,
    new_F9657_, new_F9658_, new_F9659_, new_F9660_, new_F9661_, new_F9662_,
    new_F9663_, new_F9664_, new_F9665_, new_F9666_, new_F9667_, new_F9668_,
    new_F9669_, new_F9670_, new_F9671_, new_F9672_, new_F9673_, new_F9674_,
    new_F9675_, new_F9676_, new_F9677_, new_F9678_, new_F9679_, new_F9680_,
    new_F9681_, new_F9682_, new_F9683_, new_F9684_, new_F9685_, new_F9686_,
    new_F9687_, new_F9688_, new_F9689_, new_F9690_, new_F9691_, new_F9692_,
    new_F9693_, new_F9694_, new_F9695_, new_F9696_, new_F9697_, new_F9698_,
    new_F9699_, new_F9700_, new_F9701_, new_F9702_, new_F9709_, new_F9710_,
    new_F9711_, new_F9712_, new_F9713_, new_F9714_, new_F9715_, new_F9716_,
    new_F9717_, new_F9718_, new_F9719_, new_F9720_, new_F9721_, new_F9722_,
    new_F9723_, new_F9724_, new_F9725_, new_F9726_, new_F9727_, new_F9728_,
    new_F9729_, new_F9730_, new_F9731_, new_F9732_, new_F9733_, new_F9734_,
    new_F9735_, new_F9736_, new_F9737_, new_F9738_, new_F9739_, new_F9740_,
    new_F9741_, new_F9742_, new_F9743_, new_F9744_, new_F9745_, new_F9746_,
    new_F9747_, new_F9748_, new_F9749_, new_F9750_, new_F9751_, new_F9752_,
    new_F9753_, new_F9754_, new_F9755_, new_F9756_, new_F9757_, new_F9758_,
    new_F9759_, new_F9760_, new_F9761_, new_F9762_, new_F9763_, new_F9764_,
    new_F9765_, new_F9766_, new_F9767_, new_F9768_, new_F9769_, new_F9776_,
    new_F9777_, new_F9778_, new_F9779_, new_F9780_, new_F9781_, new_F9782_,
    new_F9783_, new_F9784_, new_F9785_, new_F9786_, new_F9787_, new_F9788_,
    new_F9789_, new_F9790_, new_F9791_, new_F9792_, new_F9793_, new_F9794_,
    new_F9795_, new_F9796_, new_F9797_, new_F9798_, new_F9799_, new_F9800_,
    new_F9801_, new_F9802_, new_F9803_, new_F9804_, new_F9805_, new_F9806_,
    new_F9807_, new_F9808_, new_F9809_, new_F9810_, new_F9811_, new_F9812_,
    new_F9813_, new_F9814_, new_F9815_, new_F9816_, new_F9817_, new_F9818_,
    new_F9819_, new_F9820_, new_F9821_, new_F9822_, new_F9823_, new_F9824_,
    new_F9825_, new_F9826_, new_F9827_, new_F9828_, new_F9829_, new_F9830_,
    new_F9831_, new_F9832_, new_F9833_, new_F9834_, new_F9835_, new_F9836_,
    new_F9843_, new_F9844_, new_F9845_, new_F9846_, new_F9847_, new_F9848_,
    new_F9849_, new_F9850_, new_F9851_, new_F9852_, new_F9853_, new_F9854_,
    new_F9855_, new_F9856_, new_F9857_, new_F9858_, new_F9859_, new_F9860_,
    new_F9861_, new_F9862_, new_F9863_, new_F9864_, new_F9865_, new_F9866_,
    new_F9867_, new_F9868_, new_F9869_, new_F9870_, new_F9871_, new_F9872_,
    new_F9873_, new_F9874_, new_F9875_, new_F9876_, new_F9877_, new_F9878_,
    new_F9879_, new_F9880_, new_F9881_, new_F9882_, new_F9883_, new_F9884_,
    new_F9885_, new_F9886_, new_F9887_, new_F9888_, new_F9889_, new_F9890_,
    new_F9891_, new_F9892_, new_F9893_, new_F9894_, new_F9895_, new_F9896_,
    new_F9897_, new_F9898_, new_F9899_, new_F9900_, new_F9901_, new_F9902_,
    new_F9903_, new_F9910_, new_F9911_, new_F9912_, new_F9913_, new_F9914_,
    new_F9915_, new_F9916_, new_F9917_, new_F9918_, new_F9919_, new_F9920_,
    new_F9921_, new_F9922_, new_F9923_, new_F9924_, new_F9925_, new_F9926_,
    new_F9927_, new_F9928_, new_F9929_, new_F9930_, new_F9931_, new_F9932_,
    new_F9933_, new_F9934_, new_F9935_, new_F9936_, new_F9937_, new_F9938_,
    new_F9939_, new_F9940_, new_F9941_, new_F9942_, new_F9943_, new_F9944_,
    new_F9945_, new_F9946_, new_F9947_, new_F9948_, new_F9949_, new_F9950_,
    new_F9951_, new_F9952_, new_F9953_, new_F9954_, new_F9955_, new_F9956_,
    new_F9957_, new_F9958_, new_F9959_, new_F9960_, new_F9961_, new_F9962_,
    new_F9963_, new_F9964_, new_F9965_, new_F9966_, new_F9967_, new_F9968_,
    new_F9969_, new_F9970_, new_F9977_, new_F9978_, new_F9979_, new_F9980_,
    new_F9981_, new_F9982_, new_F9983_, new_F9984_, new_F9985_, new_F9986_,
    new_F9987_, new_F9988_, new_F9989_, new_F9990_, new_F9991_, new_F9992_,
    new_F9993_, new_F9994_, new_F9995_, new_F9996_, new_F9997_, new_F9998_,
    new_F9999_, new_G1_, new_G2_, new_G3_, new_G4_, new_G5_, new_G6_,
    new_G7_, new_G8_, new_G9_, new_G10_, new_G11_, new_G12_, new_G13_,
    new_G14_, new_G15_, new_G16_, new_G17_, new_G18_, new_G19_, new_G20_,
    new_G21_, new_G22_, new_G23_, new_G24_, new_G25_, new_G26_, new_G27_,
    new_G28_, new_G29_, new_G30_, new_G31_, new_G32_, new_G33_, new_G34_,
    new_G35_, new_G36_, new_G37_, new_G38_, new_G45_, new_G46_, new_G47_,
    new_G48_, new_G49_, new_G50_, new_G51_, new_G52_, new_G53_, new_G54_,
    new_G55_, new_G56_, new_G57_, new_G58_, new_G59_, new_G60_, new_G61_,
    new_G62_, new_G63_, new_G64_, new_G65_, new_G66_, new_G67_, new_G68_,
    new_G69_, new_G70_, new_G71_, new_G72_, new_G73_, new_G74_, new_G75_,
    new_G76_, new_G77_, new_G78_, new_G79_, new_G80_, new_G81_, new_G82_,
    new_G83_, new_G84_, new_G85_, new_G86_, new_G87_, new_G88_, new_G89_,
    new_G90_, new_G91_, new_G92_, new_G93_, new_G94_, new_G95_, new_G96_,
    new_G97_, new_G98_, new_G99_, new_G100_, new_G101_, new_G102_,
    new_G103_, new_G104_, new_G105_, new_G112_, new_G113_, new_G114_,
    new_G115_, new_G116_, new_G117_, new_G118_, new_G119_, new_G120_,
    new_G121_, new_G122_, new_G123_, new_G124_, new_G125_, new_G126_,
    new_G127_, new_G128_, new_G129_, new_G130_, new_G131_, new_G132_,
    new_G133_, new_G134_, new_G135_, new_G136_, new_G137_, new_G138_,
    new_G139_, new_G140_, new_G141_, new_G142_, new_G143_, new_G144_,
    new_G145_, new_G146_, new_G147_, new_G148_, new_G149_, new_G150_,
    new_G151_, new_G152_, new_G153_, new_G154_, new_G155_, new_G156_,
    new_G157_, new_G158_, new_G159_, new_G160_, new_G161_, new_G162_,
    new_G163_, new_G164_, new_G165_, new_G166_, new_G167_, new_G168_,
    new_G169_, new_G170_, new_G171_, new_G172_, new_G179_, new_G180_,
    new_G181_, new_G182_, new_G183_, new_G184_, new_G185_, new_G186_,
    new_G187_, new_G188_, new_G189_, new_G190_, new_G191_, new_G192_,
    new_G193_, new_G194_, new_G195_, new_G196_, new_G197_, new_G198_,
    new_G199_, new_G200_, new_G201_, new_G202_, new_G203_, new_G204_,
    new_G205_, new_G206_, new_G207_, new_G208_, new_G209_, new_G210_,
    new_G211_, new_G212_, new_G213_, new_G214_, new_G215_, new_G216_,
    new_G217_, new_G218_, new_G219_, new_G220_, new_G221_, new_G222_,
    new_G223_, new_G224_, new_G225_, new_G226_, new_G227_, new_G228_,
    new_G229_, new_G230_, new_G231_, new_G232_, new_G233_, new_G234_,
    new_G235_, new_G236_, new_G237_, new_G238_, new_G239_, new_G246_,
    new_G247_, new_G248_, new_G249_, new_G250_, new_G251_, new_G252_,
    new_G253_, new_G254_, new_G255_, new_G256_, new_G257_, new_G258_,
    new_G259_, new_G260_, new_G261_, new_G262_, new_G263_, new_G264_,
    new_G265_, new_G266_, new_G267_, new_G268_, new_G269_, new_G270_,
    new_G271_, new_G272_, new_G273_, new_G274_, new_G275_, new_G276_,
    new_G277_, new_G278_, new_G279_, new_G280_, new_G281_, new_G282_,
    new_G283_, new_G284_, new_G285_, new_G286_, new_G287_, new_G288_,
    new_G289_, new_G290_, new_G291_, new_G292_, new_G293_, new_G294_,
    new_G295_, new_G296_, new_G297_, new_G298_, new_G299_, new_G300_,
    new_G301_, new_G302_, new_G303_, new_G304_, new_G305_, new_G306_,
    new_G313_, new_G314_, new_G315_, new_G316_, new_G317_, new_G318_,
    new_G319_, new_G320_, new_G321_, new_G322_, new_G323_, new_G324_,
    new_G325_, new_G326_, new_G327_, new_G328_, new_G329_, new_G330_,
    new_G331_, new_G332_, new_G333_, new_G334_, new_G335_, new_G336_,
    new_G337_, new_G338_, new_G339_, new_G340_, new_G341_, new_G342_,
    new_G343_, new_G344_, new_G345_, new_G346_, new_G347_, new_G348_,
    new_G349_, new_G350_, new_G351_, new_G352_, new_G353_, new_G354_,
    new_G355_, new_G356_, new_G357_, new_G358_, new_G359_, new_G360_,
    new_G361_, new_G362_, new_G363_, new_G364_, new_G365_, new_G366_,
    new_G367_, new_G368_, new_G369_, new_G370_, new_G371_, new_G372_,
    new_G373_, new_G380_, new_G381_, new_G382_, new_G383_, new_G384_,
    new_G385_, new_G386_, new_G387_, new_G388_, new_G389_, new_G390_,
    new_G391_, new_G392_, new_G393_, new_G394_, new_G395_, new_G396_,
    new_G397_, new_G398_, new_G399_, new_G400_, new_G401_, new_G402_,
    new_G403_, new_G404_, new_G405_, new_G406_, new_G407_, new_G408_,
    new_G409_, new_G410_, new_G411_, new_G412_, new_G413_, new_G414_,
    new_G415_, new_G416_, new_G417_, new_G418_, new_G419_, new_G420_,
    new_G421_, new_G422_, new_G423_, new_G424_, new_G425_, new_G426_,
    new_G427_, new_G428_, new_G429_, new_G430_, new_G431_, new_G432_,
    new_G433_, new_G434_, new_G435_, new_G436_, new_G437_, new_G438_,
    new_G439_, new_G440_, new_G447_, new_G448_, new_G449_, new_G450_,
    new_G451_, new_G452_, new_G453_, new_G454_, new_G455_, new_G456_,
    new_G457_, new_G458_, new_G459_, new_G460_, new_G461_, new_G462_,
    new_G463_, new_G464_, new_G465_, new_G466_, new_G467_, new_G468_,
    new_G469_, new_G470_, new_G471_, new_G472_, new_G473_, new_G474_,
    new_G475_, new_G476_, new_G477_, new_G478_, new_G479_, new_G480_,
    new_G481_, new_G482_, new_G483_, new_G484_, new_G485_, new_G486_,
    new_G487_, new_G488_, new_G489_, new_G490_, new_G491_, new_G492_,
    new_G493_, new_G494_, new_G495_, new_G496_, new_G497_, new_G498_,
    new_G499_, new_G500_, new_G501_, new_G502_, new_G503_, new_G504_,
    new_G505_, new_G506_, new_G507_, new_G514_, new_G515_, new_G516_,
    new_G517_, new_G518_, new_G519_, new_G520_, new_G521_, new_G522_,
    new_G523_, new_G524_, new_G525_, new_G526_, new_G527_, new_G528_,
    new_G529_, new_G530_, new_G531_, new_G532_, new_G533_, new_G534_,
    new_G535_, new_G536_, new_G537_, new_G538_, new_G539_, new_G540_,
    new_G541_, new_G542_, new_G543_, new_G544_, new_G545_, new_G546_,
    new_G547_, new_G548_, new_G549_, new_G550_, new_G551_, new_G552_,
    new_G553_, new_G554_, new_G555_, new_G556_, new_G557_, new_G558_,
    new_G559_, new_G560_, new_G561_, new_G562_, new_G563_, new_G564_,
    new_G565_, new_G566_, new_G567_, new_G568_, new_G569_, new_G570_,
    new_G571_, new_G572_, new_G573_, new_G574_, new_G581_, new_G582_,
    new_G583_, new_G584_, new_G585_, new_G586_, new_G587_, new_G588_,
    new_G589_, new_G590_, new_G591_, new_G592_, new_G593_, new_G594_,
    new_G595_, new_G596_, new_G597_, new_G598_, new_G599_, new_G600_,
    new_G601_, new_G602_, new_G603_, new_G604_, new_G605_, new_G606_,
    new_G607_, new_G608_, new_G609_, new_G610_, new_G611_, new_G612_,
    new_G613_, new_G614_, new_G615_, new_G616_, new_G617_, new_G618_,
    new_G619_, new_G620_, new_G621_, new_G622_, new_G623_, new_G624_,
    new_G625_, new_G626_, new_G627_, new_G628_, new_G629_, new_G630_,
    new_G631_, new_G632_, new_G633_, new_G634_, new_G635_, new_G636_,
    new_G637_, new_G638_, new_G639_, new_G640_, new_G641_, new_G648_,
    new_G649_, new_G650_, new_G651_, new_G652_, new_G653_, new_G654_,
    new_G655_, new_G656_, new_G657_, new_G658_, new_G659_, new_G660_,
    new_G661_, new_G662_, new_G663_, new_G664_, new_G665_, new_G666_,
    new_G667_, new_G668_, new_G669_, new_G670_, new_G671_, new_G672_,
    new_G673_, new_G674_, new_G675_, new_G676_, new_G677_, new_G678_,
    new_G679_, new_G680_, new_G681_, new_G682_, new_G683_, new_G684_,
    new_G685_, new_G686_, new_G687_, new_G688_, new_G689_, new_G690_,
    new_G691_, new_G692_, new_G693_, new_G694_, new_G695_, new_G696_,
    new_G697_, new_G698_, new_G699_, new_G700_, new_G701_, new_G702_,
    new_G703_, new_G704_, new_G705_, new_G706_, new_G707_, new_G708_,
    new_G715_, new_G716_, new_G717_, new_G718_, new_G719_, new_G720_,
    new_G721_, new_G722_, new_G723_, new_G724_, new_G725_, new_G726_,
    new_G727_, new_G728_, new_G729_, new_G730_, new_G731_, new_G732_,
    new_G733_, new_G734_, new_G735_, new_G736_, new_G737_, new_G738_,
    new_G739_, new_G740_, new_G741_, new_G742_, new_G743_, new_G744_,
    new_G745_, new_G746_, new_G747_, new_G748_, new_G749_, new_G750_,
    new_G751_, new_G752_, new_G753_, new_G754_, new_G755_, new_G756_,
    new_G757_, new_G758_, new_G759_, new_G760_, new_G761_, new_G762_,
    new_G763_, new_G764_, new_G765_, new_G766_, new_G767_, new_G768_,
    new_G769_, new_G770_, new_G771_, new_G772_, new_G773_, new_G774_,
    new_G775_, new_G782_, new_G783_, new_G784_, new_G785_, new_G786_,
    new_G787_, new_G788_, new_G789_, new_G790_, new_G791_, new_G792_,
    new_G793_, new_G794_, new_G795_, new_G796_, new_G797_, new_G798_,
    new_G799_, new_G800_, new_G801_, new_G802_, new_G803_, new_G804_,
    new_G805_, new_G806_, new_G807_, new_G808_, new_G809_, new_G810_,
    new_G811_, new_G812_, new_G813_, new_G814_, new_G815_, new_G816_,
    new_G817_, new_G818_, new_G819_, new_G820_, new_G821_, new_G822_,
    new_G823_, new_G824_, new_G825_, new_G826_, new_G827_, new_G828_,
    new_G829_, new_G830_, new_G831_, new_G832_, new_G833_, new_G834_,
    new_G835_, new_G836_, new_G837_, new_G838_, new_G839_, new_G840_,
    new_G841_, new_G842_, new_G849_, new_G850_, new_G851_, new_G852_,
    new_G853_, new_G854_, new_G855_, new_G856_, new_G857_, new_G858_,
    new_G859_, new_G860_, new_G861_, new_G862_, new_G863_, new_G864_,
    new_G865_, new_G866_, new_G867_, new_G868_, new_G869_, new_G870_,
    new_G871_, new_G872_, new_G873_, new_G874_, new_G875_, new_G876_,
    new_G877_, new_G878_, new_G879_, new_G880_, new_G881_, new_G882_,
    new_G883_, new_G884_, new_G885_, new_G886_, new_G887_, new_G888_,
    new_G889_, new_G890_, new_G891_, new_G892_, new_G893_, new_G894_,
    new_G895_, new_G896_, new_G897_, new_G898_, new_G899_, new_G900_,
    new_G901_, new_G902_, new_G903_, new_G904_, new_G905_, new_G906_,
    new_G907_, new_G908_, new_G909_, new_G916_, new_G917_, new_G918_,
    new_G919_, new_G920_, new_G921_, new_G922_, new_G923_, new_G924_,
    new_G925_, new_G926_, new_G927_, new_G928_, new_G929_, new_G930_,
    new_G931_, new_G932_, new_G933_, new_G934_, new_G935_, new_G936_,
    new_G937_, new_G938_, new_G939_, new_G940_, new_G941_, new_G942_,
    new_G943_, new_G944_, new_G945_, new_G946_, new_G947_, new_G948_,
    new_G949_, new_G950_, new_G951_, new_G952_, new_G953_, new_G954_,
    new_G955_, new_G956_, new_G957_, new_G958_, new_G959_, new_G960_,
    new_G961_, new_G962_, new_G963_, new_G964_, new_G965_, new_G966_,
    new_G967_, new_G968_, new_G969_, new_G970_, new_G971_, new_G972_,
    new_G973_, new_G974_, new_G975_, new_G976_, new_G983_, new_G984_,
    new_G985_, new_G986_, new_G987_, new_G988_, new_G989_, new_G990_,
    new_G991_, new_G992_, new_G993_, new_G994_, new_G995_, new_G996_,
    new_G997_, new_G998_, new_G999_, new_G1000_, new_G1001_, new_G1002_,
    new_G1003_, new_G1004_, new_G1005_, new_G1006_, new_G1007_, new_G1008_,
    new_G1009_, new_G1010_, new_G1011_, new_G1012_, new_G1013_, new_G1014_,
    new_G1015_, new_G1016_, new_G1017_, new_G1018_, new_G1019_, new_G1020_,
    new_G1021_, new_G1022_, new_G1023_, new_G1024_, new_G1025_, new_G1026_,
    new_G1027_, new_G1028_, new_G1029_, new_G1030_, new_G1031_, new_G1032_,
    new_G1033_, new_G1034_, new_G1035_, new_G1036_, new_G1037_, new_G1038_,
    new_G1039_, new_G1040_, new_G1041_, new_G1042_, new_G1043_, new_G1050_,
    new_G1051_, new_G1052_, new_G1053_, new_G1054_, new_G1055_, new_G1056_,
    new_G1057_, new_G1058_, new_G1059_, new_G1060_, new_G1061_, new_G1062_,
    new_G1063_, new_G1064_, new_G1065_, new_G1066_, new_G1067_, new_G1068_,
    new_G1069_, new_G1070_, new_G1071_, new_G1072_, new_G1073_, new_G1074_,
    new_G1075_, new_G1076_, new_G1077_, new_G1078_, new_G1079_, new_G1080_,
    new_G1081_, new_G1082_, new_G1083_, new_G1084_, new_G1085_, new_G1086_,
    new_G1087_, new_G1088_, new_G1089_, new_G1090_, new_G1091_, new_G1092_,
    new_G1093_, new_G1094_, new_G1095_, new_G1096_, new_G1097_, new_G1098_,
    new_G1099_, new_G1100_, new_G1101_, new_G1102_, new_G1103_, new_G1104_,
    new_G1105_, new_G1106_, new_G1107_, new_G1108_, new_G1109_, new_G1110_,
    new_G1117_, new_G1118_, new_G1119_, new_G1120_, new_G1121_, new_G1122_,
    new_G1123_, new_G1124_, new_G1125_, new_G1126_, new_G1127_, new_G1128_,
    new_G1129_, new_G1130_, new_G1131_, new_G1132_, new_G1133_, new_G1134_,
    new_G1135_, new_G1136_, new_G1137_, new_G1138_, new_G1139_, new_G1140_,
    new_G1141_, new_G1142_, new_G1143_, new_G1144_, new_G1145_, new_G1146_,
    new_G1147_, new_G1148_, new_G1149_, new_G1150_, new_G1151_, new_G1152_,
    new_G1153_, new_G1154_, new_G1155_, new_G1156_, new_G1157_, new_G1158_,
    new_G1159_, new_G1160_, new_G1161_, new_G1162_, new_G1163_, new_G1164_,
    new_G1165_, new_G1166_, new_G1167_, new_G1168_, new_G1169_, new_G1170_,
    new_G1171_, new_G1172_, new_G1173_, new_G1174_, new_G1175_, new_G1176_,
    new_G1177_, new_G1184_, new_G1185_, new_G1186_, new_G1187_, new_G1188_,
    new_G1189_, new_G1190_, new_G1191_, new_G1192_, new_G1193_, new_G1194_,
    new_G1195_, new_G1196_, new_G1197_, new_G1198_, new_G1199_, new_G1200_,
    new_G1201_, new_G1202_, new_G1203_, new_G1204_, new_G1205_, new_G1206_,
    new_G1207_, new_G1208_, new_G1209_, new_G1210_, new_G1211_, new_G1212_,
    new_G1213_, new_G1214_, new_G1215_, new_G1216_, new_G1217_, new_G1218_,
    new_G1219_, new_G1220_, new_G1221_, new_G1222_, new_G1223_, new_G1224_,
    new_G1225_, new_G1226_, new_G1227_, new_G1228_, new_G1229_, new_G1230_,
    new_G1231_, new_G1232_, new_G1233_, new_G1234_, new_G1235_, new_G1236_,
    new_G1237_, new_G1238_, new_G1239_, new_G1240_, new_G1241_, new_G1242_,
    new_G1243_, new_G1244_, new_G1251_, new_G1252_, new_G1253_, new_G1254_,
    new_G1255_, new_G1256_, new_G1257_, new_G1258_, new_G1259_, new_G1260_,
    new_G1261_, new_G1262_, new_G1263_, new_G1264_, new_G1265_, new_G1266_,
    new_G1267_, new_G1268_, new_G1269_, new_G1270_, new_G1271_, new_G1272_,
    new_G1273_, new_G1274_, new_G1275_, new_G1276_, new_G1277_, new_G1278_,
    new_G1279_, new_G1280_, new_G1281_, new_G1282_, new_G1283_, new_G1284_,
    new_G1285_, new_G1286_, new_G1287_, new_G1288_, new_G1289_, new_G1290_,
    new_G1291_, new_G1292_, new_G1293_, new_G1294_, new_G1295_, new_G1296_,
    new_G1297_, new_G1298_, new_G1299_, new_G1300_, new_G1301_, new_G1302_,
    new_G1303_, new_G1304_, new_G1305_, new_G1306_, new_G1307_, new_G1308_,
    new_G1309_, new_G1310_, new_G1311_, new_G1318_, new_G1319_, new_G1320_,
    new_G1321_, new_G1322_, new_G1323_, new_G1324_, new_G1325_, new_G1326_,
    new_G1327_, new_G1328_, new_G1329_, new_G1330_, new_G1331_, new_G1332_,
    new_G1333_, new_G1334_, new_G1335_, new_G1336_, new_G1337_, new_G1338_,
    new_G1339_, new_G1340_, new_G1341_, new_G1342_, new_G1343_, new_G1344_,
    new_G1345_, new_G1346_, new_G1347_, new_G1348_, new_G1349_, new_G1350_,
    new_G1351_, new_G1352_, new_G1353_, new_G1354_, new_G1355_, new_G1356_,
    new_G1357_, new_G1358_, new_G1359_, new_G1360_, new_G1361_, new_G1362_,
    new_G1363_, new_G1364_, new_G1365_, new_G1366_, new_G1367_, new_G1368_,
    new_G1369_, new_G1370_, new_G1371_, new_G1372_, new_G1373_, new_G1374_,
    new_G1375_, new_G1376_, new_G1377_, new_G1378_, new_G1385_, new_G1386_,
    new_G1387_, new_G1388_, new_G1389_, new_G1390_, new_G1391_, new_G1392_,
    new_G1393_, new_G1394_, new_G1395_, new_G1396_, new_G1397_, new_G1398_,
    new_G1399_, new_G1400_, new_G1401_, new_G1402_, new_G1403_, new_G1404_,
    new_G1405_, new_G1406_, new_G1407_, new_G1408_, new_G1409_, new_G1410_,
    new_G1411_, new_G1412_, new_G1413_, new_G1414_, new_G1415_, new_G1416_,
    new_G1417_, new_G1418_, new_G1419_, new_G1420_, new_G1421_, new_G1422_,
    new_G1423_, new_G1424_, new_G1425_, new_G1426_, new_G1427_, new_G1428_,
    new_G1429_, new_G1430_, new_G1431_, new_G1432_, new_G1433_, new_G1434_,
    new_G1435_, new_G1436_, new_G1437_, new_G1438_, new_G1439_, new_G1440_,
    new_G1441_, new_G1442_, new_G1443_, new_G1444_, new_G1445_, new_G1452_,
    new_G1453_, new_G1454_, new_G1455_, new_G1456_, new_G1457_, new_G1458_,
    new_G1459_, new_G1460_, new_G1461_, new_G1462_, new_G1463_, new_G1464_,
    new_G1465_, new_G1466_, new_G1467_, new_G1468_, new_G1469_, new_G1470_,
    new_G1471_, new_G1472_, new_G1473_, new_G1474_, new_G1475_, new_G1476_,
    new_G1477_, new_G1478_, new_G1479_, new_G1480_, new_G1481_, new_G1482_,
    new_G1483_, new_G1484_, new_G1485_, new_G1486_, new_G1487_, new_G1488_,
    new_G1489_, new_G1490_, new_G1491_, new_G1492_, new_G1493_, new_G1494_,
    new_G1495_, new_G1496_, new_G1497_, new_G1498_, new_G1499_, new_G1500_,
    new_G1501_, new_G1502_, new_G1503_, new_G1504_, new_G1505_, new_G1506_,
    new_G1507_, new_G1508_, new_G1509_, new_G1510_, new_G1511_, new_G1512_,
    new_G1519_, new_G1520_, new_G1521_, new_G1522_, new_G1523_, new_G1524_,
    new_G1525_, new_G1526_, new_G1527_, new_G1528_, new_G1529_, new_G1530_,
    new_G1531_, new_G1532_, new_G1533_, new_G1534_, new_G1535_, new_G1536_,
    new_G1537_, new_G1538_, new_G1539_, new_G1540_, new_G1541_, new_G1542_,
    new_G1543_, new_G1544_, new_G1545_, new_G1546_, new_G1547_, new_G1548_,
    new_G1549_, new_G1550_, new_G1551_, new_G1552_, new_G1553_, new_G1554_,
    new_G1555_, new_G1556_, new_G1557_, new_G1558_, new_G1559_, new_G1560_,
    new_G1561_, new_G1562_, new_G1563_, new_G1564_, new_G1565_, new_G1566_,
    new_G1567_, new_G1568_, new_G1569_, new_G1570_, new_G1571_, new_G1572_,
    new_G1573_, new_G1574_, new_G1575_, new_G1576_, new_G1577_, new_G1578_,
    new_G1579_, new_G1586_, new_G1587_, new_G1588_, new_G1589_, new_G1590_,
    new_G1591_, new_G1592_, new_G1593_, new_G1594_, new_G1595_, new_G1596_,
    new_G1597_, new_G1598_, new_G1599_, new_G1600_, new_G1601_, new_G1602_,
    new_G1603_, new_G1604_, new_G1605_, new_G1606_, new_G1607_, new_G1608_,
    new_G1609_, new_G1610_, new_G1611_, new_G1612_, new_G1613_, new_G1614_,
    new_G1615_, new_G1616_, new_G1617_, new_G1618_, new_G1619_, new_G1620_,
    new_G1621_, new_G1622_, new_G1623_, new_G1624_, new_G1625_, new_G1626_,
    new_G1627_, new_G1628_, new_G1629_, new_G1630_, new_G1631_, new_G1632_,
    new_G1633_, new_G1634_, new_G1635_, new_G1636_, new_G1637_, new_G1638_,
    new_G1639_, new_G1640_, new_G1641_, new_G1642_, new_G1643_, new_G1644_,
    new_G1645_, new_G1646_, new_G1653_, new_G1654_, new_G1655_, new_G1656_,
    new_G1657_, new_G1658_, new_G1659_, new_G1660_, new_G1661_, new_G1662_,
    new_G1663_, new_G1664_, new_G1665_, new_G1666_, new_G1667_, new_G1668_,
    new_G1669_, new_G1670_, new_G1671_, new_G1672_, new_G1673_, new_G1674_,
    new_G1675_, new_G1676_, new_G1677_, new_G1678_, new_G1679_, new_G1680_,
    new_G1681_, new_G1682_, new_G1683_, new_G1684_, new_G1685_, new_G1686_,
    new_G1687_, new_G1688_, new_G1689_, new_G1690_, new_G1691_, new_G1692_,
    new_G1693_, new_G1694_, new_G1695_, new_G1696_, new_G1697_, new_G1698_,
    new_G1699_, new_G1700_, new_G1701_, new_G1702_, new_G1703_, new_G1704_,
    new_G1705_, new_G1706_, new_G1707_, new_G1708_, new_G1709_, new_G1710_,
    new_G1711_, new_G1712_, new_G1713_, new_G1720_, new_G1721_, new_G1722_,
    new_G1723_, new_G1724_, new_G1725_, new_G1726_, new_G1727_, new_G1728_,
    new_G1729_, new_G1730_, new_G1731_, new_G1732_, new_G1733_, new_G1734_,
    new_G1735_, new_G1736_, new_G1737_, new_G1738_, new_G1739_, new_G1740_,
    new_G1741_, new_G1742_, new_G1743_, new_G1744_, new_G1745_, new_G1746_,
    new_G1747_, new_G1748_, new_G1749_, new_G1750_, new_G1751_, new_G1752_,
    new_G1753_, new_G1754_, new_G1755_, new_G1756_, new_G1757_, new_G1758_,
    new_G1759_, new_G1760_, new_G1761_, new_G1762_, new_G1763_, new_G1764_,
    new_G1765_, new_G1766_, new_G1767_, new_G1768_, new_G1769_, new_G1770_,
    new_G1771_, new_G1772_, new_G1773_, new_G1774_, new_G1775_, new_G1776_,
    new_G1777_, new_G1778_, new_G1779_, new_G1780_, new_G1787_, new_G1788_,
    new_G1789_, new_G1790_, new_G1791_, new_G1792_, new_G1793_, new_G1794_,
    new_G1795_, new_G1796_, new_G1797_, new_G1798_, new_G1799_, new_G1800_,
    new_G1801_, new_G1802_, new_G1803_, new_G1804_, new_G1805_, new_G1806_,
    new_G1807_, new_G1808_, new_G1809_, new_G1810_, new_G1811_, new_G1812_,
    new_G1813_, new_G1814_, new_G1815_, new_G1816_, new_G1817_, new_G1818_,
    new_G1819_, new_G1820_, new_G1821_, new_G1822_, new_G1823_, new_G1824_,
    new_G1825_, new_G1826_, new_G1827_, new_G1828_, new_G1829_, new_G1830_,
    new_G1831_, new_G1832_, new_G1833_, new_G1834_, new_G1835_, new_G1836_,
    new_G1837_, new_G1838_, new_G1839_, new_G1840_, new_G1841_, new_G1842_,
    new_G1843_, new_G1844_, new_G1845_, new_G1846_, new_G1847_, new_G1854_,
    new_G1855_, new_G1856_, new_G1857_, new_G1858_, new_G1859_, new_G1860_,
    new_G1861_, new_G1862_, new_G1863_, new_G1864_, new_G1865_, new_G1866_,
    new_G1867_, new_G1868_, new_G1869_, new_G1870_, new_G1871_, new_G1872_,
    new_G1873_, new_G1874_, new_G1875_, new_G1876_, new_G1877_, new_G1878_,
    new_G1879_, new_G1880_, new_G1881_, new_G1882_, new_G1883_, new_G1884_,
    new_G1885_, new_G1886_, new_G1887_, new_G1888_, new_G1889_, new_G1890_,
    new_G1891_, new_G1892_, new_G1893_, new_G1894_, new_G1895_, new_G1896_,
    new_G1897_, new_G1898_, new_G1899_, new_G1900_, new_G1901_, new_G1902_,
    new_G1903_, new_G1904_, new_G1905_, new_G1906_, new_G1907_, new_G1908_,
    new_G1909_, new_G1910_, new_G1911_, new_G1912_, new_G1913_, new_G1914_,
    new_G1921_, new_G1922_, new_G1923_, new_G1924_, new_G1925_, new_G1926_,
    new_G1927_, new_G1928_, new_G1929_, new_G1930_, new_G1931_, new_G1932_,
    new_G1933_, new_G1934_, new_G1935_, new_G1936_, new_G1937_, new_G1938_,
    new_G1939_, new_G1940_, new_G1941_, new_G1942_, new_G1943_, new_G1944_,
    new_G1945_, new_G1946_, new_G1947_, new_G1948_, new_G1949_, new_G1950_,
    new_G1951_, new_G1952_, new_G1953_, new_G1954_, new_G1955_, new_G1956_,
    new_G1957_, new_G1958_, new_G1959_, new_G1960_, new_G1961_, new_G1962_,
    new_G1963_, new_G1964_, new_G1965_, new_G1966_, new_G1967_, new_G1968_,
    new_G1969_, new_G1970_, new_G1971_, new_G1972_, new_G1973_, new_G1974_,
    new_G1975_, new_G1976_, new_G1977_, new_G1978_, new_G1979_, new_G1980_,
    new_G1981_, new_G1988_, new_G1989_, new_G1990_, new_G1991_, new_G1992_,
    new_G1993_, new_G1994_, new_G1995_, new_G1996_, new_G1997_, new_G1998_,
    new_G1999_, new_G2000_, new_G2001_, new_G2002_, new_G2003_, new_G2004_,
    new_G2005_, new_G2006_, new_G2007_, new_G2008_, new_G2009_, new_G2010_,
    new_G2011_, new_G2012_, new_G2013_, new_G2014_, new_G2015_, new_G2016_,
    new_G2017_, new_G2018_, new_G2019_, new_G2020_, new_G2021_, new_G2022_,
    new_G2023_, new_G2024_, new_G2025_, new_G2026_, new_G2027_, new_G2028_,
    new_G2029_, new_G2030_, new_G2031_, new_G2032_, new_G2033_, new_G2034_,
    new_G2035_, new_G2036_, new_G2037_, new_G2038_, new_G2039_, new_G2040_,
    new_G2041_, new_G2042_, new_G2043_, new_G2044_, new_G2045_, new_G2046_,
    new_G2047_, new_G2048_, new_G2055_, new_G2056_, new_G2057_, new_G2058_,
    new_G2059_, new_G2060_, new_G2061_, new_G2062_, new_G2063_, new_G2064_,
    new_G2065_, new_G2066_, new_G2067_, new_G2068_, new_G2069_, new_G2070_,
    new_G2071_, new_G2072_, new_G2073_, new_G2074_, new_G2075_, new_G2076_,
    new_G2077_, new_G2078_, new_G2079_, new_G2080_, new_G2081_, new_G2082_,
    new_G2083_, new_G2084_, new_G2085_, new_G2086_, new_G2087_, new_G2088_,
    new_G2089_, new_G2090_, new_G2091_, new_G2092_, new_G2093_, new_G2094_,
    new_G2095_, new_G2096_, new_G2097_, new_G2098_, new_G2099_, new_G2100_,
    new_G2101_, new_G2102_, new_G2103_, new_G2104_, new_G2105_, new_G2106_,
    new_G2107_, new_G2108_, new_G2109_, new_G2110_, new_G2111_, new_G2112_,
    new_G2113_, new_G2114_, new_G2115_, new_G2122_, new_G2123_, new_G2124_,
    new_G2125_, new_G2126_, new_G2127_, new_G2128_, new_G2129_, new_G2130_,
    new_G2131_, new_G2132_, new_G2133_, new_G2134_, new_G2135_, new_G2136_,
    new_G2137_, new_G2138_, new_G2139_, new_G2140_, new_G2141_, new_G2142_,
    new_G2143_, new_G2144_, new_G2145_, new_G2146_, new_G2147_, new_G2148_,
    new_G2149_, new_G2150_, new_G2151_, new_G2152_, new_G2153_, new_G2154_,
    new_G2155_, new_G2156_, new_G2157_, new_G2158_, new_G2159_, new_G2160_,
    new_G2161_, new_G2162_, new_G2163_, new_G2164_, new_G2165_, new_G2166_,
    new_G2167_, new_G2168_, new_G2169_, new_G2170_, new_G2171_, new_G2172_,
    new_G2173_, new_G2174_, new_G2175_, new_G2176_, new_G2177_, new_G2178_,
    new_G2179_, new_G2180_, new_G2181_, new_G2182_, new_G2189_, new_G2190_,
    new_G2191_, new_G2192_, new_G2193_, new_G2194_, new_G2195_, new_G2196_,
    new_G2197_, new_G2198_, new_G2199_, new_G2200_, new_G2201_, new_G2202_,
    new_G2203_, new_G2204_, new_G2205_, new_G2206_, new_G2207_, new_G2208_,
    new_G2209_, new_G2210_, new_G2211_, new_G2212_, new_G2213_, new_G2214_,
    new_G2215_, new_G2216_, new_G2217_, new_G2218_, new_G2219_, new_G2220_,
    new_G2221_, new_G2222_, new_G2223_, new_G2224_, new_G2225_, new_G2226_,
    new_G2227_, new_G2228_, new_G2229_, new_G2230_, new_G2231_, new_G2232_,
    new_G2233_, new_G2234_, new_G2235_, new_G2236_, new_G2237_, new_G2238_,
    new_G2239_, new_G2240_, new_G2241_, new_G2242_, new_G2243_, new_G2244_,
    new_G2245_, new_G2246_, new_G2247_, new_G2248_, new_G2249_, new_G2256_,
    new_G2257_, new_G2258_, new_G2259_, new_G2260_, new_G2261_, new_G2262_,
    new_G2263_, new_G2264_, new_G2265_, new_G2266_, new_G2267_, new_G2268_,
    new_G2269_, new_G2270_, new_G2271_, new_G2272_, new_G2273_, new_G2274_,
    new_G2275_, new_G2276_, new_G2277_, new_G2278_, new_G2279_, new_G2280_,
    new_G2281_, new_G2282_, new_G2283_, new_G2284_, new_G2285_, new_G2286_,
    new_G2287_, new_G2288_, new_G2289_, new_G2290_, new_G2291_, new_G2292_,
    new_G2293_, new_G2294_, new_G2295_, new_G2296_, new_G2297_, new_G2298_,
    new_G2299_, new_G2300_, new_G2301_, new_G2302_, new_G2303_, new_G2304_,
    new_G2305_, new_G2306_, new_G2307_, new_G2308_, new_G2309_, new_G2310_,
    new_G2311_, new_G2312_, new_G2313_, new_G2314_, new_G2315_, new_G2316_,
    new_G2323_, new_G2324_, new_G2325_, new_G2326_, new_G2327_, new_G2328_,
    new_G2329_, new_G2330_, new_G2331_, new_G2332_, new_G2333_, new_G2334_,
    new_G2335_, new_G2336_, new_G2337_, new_G2338_, new_G2339_, new_G2340_,
    new_G2341_, new_G2342_, new_G2343_, new_G2344_, new_G2345_, new_G2346_,
    new_G2347_, new_G2348_, new_G2349_, new_G2350_, new_G2351_, new_G2352_,
    new_G2353_, new_G2354_, new_G2355_, new_G2356_, new_G2357_, new_G2358_,
    new_G2359_, new_G2360_, new_G2361_, new_G2362_, new_G2363_, new_G2364_,
    new_G2365_, new_G2366_, new_G2367_, new_G2368_, new_G2369_, new_G2370_,
    new_G2371_, new_G2372_, new_G2373_, new_G2374_, new_G2375_, new_G2376_,
    new_G2377_, new_G2378_, new_G2379_, new_G2380_, new_G2381_, new_G2382_,
    new_G2383_, new_G2390_, new_G2391_, new_G2392_, new_G2393_, new_G2394_,
    new_G2395_, new_G2396_, new_G2397_, new_G2398_, new_G2399_, new_G2400_,
    new_G2401_, new_G2402_, new_G2403_, new_G2404_, new_G2405_, new_G2406_,
    new_G2407_, new_G2408_, new_G2409_, new_G2410_, new_G2411_, new_G2412_,
    new_G2413_, new_G2414_, new_G2415_, new_G2416_, new_G2417_, new_G2418_,
    new_G2419_, new_G2420_, new_G2421_, new_G2422_, new_G2423_, new_G2424_,
    new_G2425_, new_G2426_, new_G2427_, new_G2428_, new_G2429_, new_G2430_,
    new_G2431_, new_G2432_, new_G2433_, new_G2434_, new_G2435_, new_G2436_,
    new_G2437_, new_G2438_, new_G2439_, new_G2440_, new_G2441_, new_G2442_,
    new_G2443_, new_G2444_, new_G2445_, new_G2446_, new_G2447_, new_G2448_,
    new_G2449_, new_G2450_, new_G2457_, new_G2458_, new_G2459_, new_G2460_,
    new_G2461_, new_G2462_, new_G2463_, new_G2464_, new_G2465_, new_G2466_,
    new_G2467_, new_G2468_, new_G2469_, new_G2470_, new_G2471_, new_G2472_,
    new_G2473_, new_G2474_, new_G2475_, new_G2476_, new_G2477_, new_G2478_,
    new_G2479_, new_G2480_, new_G2481_, new_G2482_, new_G2483_, new_G2484_,
    new_G2485_, new_G2486_, new_G2487_, new_G2488_, new_G2489_, new_G2490_,
    new_G2491_, new_G2492_, new_G2493_, new_G2494_, new_G2495_, new_G2496_,
    new_G2497_, new_G2498_, new_G2499_, new_G2500_, new_G2501_, new_G2502_,
    new_G2503_, new_G2504_, new_G2505_, new_G2506_, new_G2507_, new_G2508_,
    new_G2509_, new_G2510_, new_G2511_, new_G2512_, new_G2513_, new_G2514_,
    new_G2515_, new_G2516_, new_G2517_, new_G2524_, new_G2525_, new_G2526_,
    new_G2527_, new_G2528_, new_G2529_, new_G2530_, new_G2531_, new_G2532_,
    new_G2533_, new_G2534_, new_G2535_, new_G2536_, new_G2537_, new_G2538_,
    new_G2539_, new_G2540_, new_G2541_, new_G2542_, new_G2543_, new_G2544_,
    new_G2545_, new_G2546_, new_G2547_, new_G2548_, new_G2549_, new_G2550_,
    new_G2551_, new_G2552_, new_G2553_, new_G2554_, new_G2555_, new_G2556_,
    new_G2557_, new_G2558_, new_G2559_, new_G2560_, new_G2561_, new_G2562_,
    new_G2563_, new_G2564_, new_G2565_, new_G2566_, new_G2567_, new_G2568_,
    new_G2569_, new_G2570_, new_G2571_, new_G2572_, new_G2573_, new_G2574_,
    new_G2575_, new_G2576_, new_G2577_, new_G2578_, new_G2579_, new_G2580_,
    new_G2581_, new_G2582_, new_G2583_, new_G2584_, new_G2591_, new_G2592_,
    new_G2593_, new_G2594_, new_G2595_, new_G2596_, new_G2597_, new_G2598_,
    new_G2599_, new_G2600_, new_G2601_, new_G2602_, new_G2603_, new_G2604_,
    new_G2605_, new_G2606_, new_G2607_, new_G2608_, new_G2609_, new_G2610_,
    new_G2611_, new_G2612_, new_G2613_, new_G2614_, new_G2615_, new_G2616_,
    new_G2617_, new_G2618_, new_G2619_, new_G2620_, new_G2621_, new_G2622_,
    new_G2623_, new_G2624_, new_G2625_, new_G2626_, new_G2627_, new_G2628_,
    new_G2629_, new_G2630_, new_G2631_, new_G2632_, new_G2633_, new_G2634_,
    new_G2635_, new_G2636_, new_G2637_, new_G2638_, new_G2639_, new_G2640_,
    new_G2641_, new_G2642_, new_G2643_, new_G2644_, new_G2645_, new_G2646_,
    new_G2647_, new_G2648_, new_G2649_, new_G2650_, new_G2651_, new_G2658_,
    new_G2659_, new_G2660_, new_G2661_, new_G2662_, new_G2663_, new_G2664_,
    new_G2665_, new_G2666_, new_G2667_, new_G2668_, new_G2669_, new_G2670_,
    new_G2671_, new_G2672_, new_G2673_, new_G2674_, new_G2675_, new_G2676_,
    new_G2677_, new_G2678_, new_G2679_, new_G2680_, new_G2681_, new_G2682_,
    new_G2683_, new_G2684_, new_G2685_, new_G2686_, new_G2687_, new_G2688_,
    new_G2689_, new_G2690_, new_G2691_, new_G2692_, new_G2693_, new_G2694_,
    new_G2695_, new_G2696_, new_G2697_, new_G2698_, new_G2699_, new_G2700_,
    new_G2701_, new_G2702_, new_G2703_, new_G2704_, new_G2705_, new_G2706_,
    new_G2707_, new_G2708_, new_G2709_, new_G2710_, new_G2711_, new_G2712_,
    new_G2713_, new_G2714_, new_G2715_, new_G2716_, new_G2717_, new_G2718_,
    new_G2725_, new_G2726_, new_G2727_, new_G2728_, new_G2729_, new_G2730_,
    new_G2731_, new_G2732_, new_G2733_, new_G2734_, new_G2735_, new_G2736_,
    new_G2737_, new_G2738_, new_G2739_, new_G2740_, new_G2741_, new_G2742_,
    new_G2743_, new_G2744_, new_G2745_, new_G2746_, new_G2747_, new_G2748_,
    new_G2749_, new_G2750_, new_G2751_, new_G2752_, new_G2753_, new_G2754_,
    new_G2755_, new_G2756_, new_G2757_, new_G2758_, new_G2759_, new_G2760_,
    new_G2761_, new_G2762_, new_G2763_, new_G2764_, new_G2765_, new_G2766_,
    new_G2767_, new_G2768_, new_G2769_, new_G2770_, new_G2771_, new_G2772_,
    new_G2773_, new_G2774_, new_G2775_, new_G2776_, new_G2777_, new_G2778_,
    new_G2779_, new_G2780_, new_G2781_, new_G2782_, new_G2783_, new_G2784_,
    new_G2785_, new_G2792_, new_G2793_, new_G2794_, new_G2795_, new_G2796_,
    new_G2797_, new_G2798_, new_G2799_, new_G2800_, new_G2801_, new_G2802_,
    new_G2803_, new_G2804_, new_G2805_, new_G2806_, new_G2807_, new_G2808_,
    new_G2809_, new_G2810_, new_G2811_, new_G2812_, new_G2813_, new_G2814_,
    new_G2815_, new_G2816_, new_G2817_, new_G2818_, new_G2819_, new_G2820_,
    new_G2821_, new_G2822_, new_G2823_, new_G2824_, new_G2825_, new_G2826_,
    new_G2827_, new_G2828_, new_G2829_, new_G2830_, new_G2831_, new_G2832_,
    new_G2833_, new_G2834_, new_G2835_, new_G2836_, new_G2837_, new_G2838_,
    new_G2839_, new_G2840_, new_G2841_, new_G2842_, new_G2843_, new_G2844_,
    new_G2845_, new_G2846_, new_G2847_, new_G2848_, new_G2849_, new_G2850_,
    new_G2851_, new_G2852_, new_G2859_, new_G2860_, new_G2861_, new_G2862_,
    new_G2863_, new_G2864_, new_G2865_, new_G2866_, new_G2867_, new_G2868_,
    new_G2869_, new_G2870_, new_G2871_, new_G2872_, new_G2873_, new_G2874_,
    new_G2875_, new_G2876_, new_G2877_, new_G2878_, new_G2879_, new_G2880_,
    new_G2881_, new_G2882_, new_G2883_, new_G2884_, new_G2885_, new_G2886_,
    new_G2887_, new_G2888_, new_G2889_, new_G2890_, new_G2891_, new_G2892_,
    new_G2893_, new_G2894_, new_G2895_, new_G2896_, new_G2897_, new_G2898_,
    new_G2899_, new_G2900_, new_G2901_, new_G2902_, new_G2903_, new_G2904_,
    new_G2905_, new_G2906_, new_G2907_, new_G2908_, new_G2909_, new_G2910_,
    new_G2911_, new_G2912_, new_G2913_, new_G2914_, new_G2915_, new_G2916_,
    new_G2917_, new_G2918_, new_G2919_, new_G2926_, new_G2927_, new_G2928_,
    new_G2929_, new_G2930_, new_G2931_, new_G2932_, new_G2933_, new_G2934_,
    new_G2935_, new_G2936_, new_G2937_, new_G2938_, new_G2939_, new_G2940_,
    new_G2941_, new_G2942_, new_G2943_, new_G2944_, new_G2945_, new_G2946_,
    new_G2947_, new_G2948_, new_G2949_, new_G2950_, new_G2951_, new_G2952_,
    new_G2953_, new_G2954_, new_G2955_, new_G2956_, new_G2957_, new_G2958_,
    new_G2959_, new_G2960_, new_G2961_, new_G2962_, new_G2963_, new_G2964_,
    new_G2965_, new_G2966_, new_G2967_, new_G2968_, new_G2969_, new_G2970_,
    new_G2971_, new_G2972_, new_G2973_, new_G2974_, new_G2975_, new_G2976_,
    new_G2977_, new_G2978_, new_G2979_, new_G2980_, new_G2981_, new_G2982_,
    new_G2983_, new_G2984_, new_G2985_, new_G2986_, new_G2993_, new_G2994_,
    new_G2995_, new_G2996_, new_G2997_, new_G2998_, new_G2999_, new_G3000_,
    new_G3001_, new_G3002_, new_G3003_, new_G3004_, new_G3005_, new_G3006_,
    new_G3007_, new_G3008_, new_G3009_, new_G3010_, new_G3011_, new_G3012_,
    new_G3013_, new_G3014_, new_G3015_, new_G3016_, new_G3017_, new_G3018_,
    new_G3019_, new_G3020_, new_G3021_, new_G3022_, new_G3023_, new_G3024_,
    new_G3025_, new_G3026_, new_G3027_, new_G3028_, new_G3029_, new_G3030_,
    new_G3031_, new_G3032_, new_G3033_, new_G3034_, new_G3035_, new_G3036_,
    new_G3037_, new_G3038_, new_G3039_, new_G3040_, new_G3041_, new_G3042_,
    new_G3043_, new_G3044_, new_G3045_, new_G3046_, new_G3047_, new_G3048_,
    new_G3049_, new_G3050_, new_G3051_, new_G3052_, new_G3053_, new_G3060_,
    new_G3061_, new_G3062_, new_G3063_, new_G3064_, new_G3065_, new_G3066_,
    new_G3067_, new_G3068_, new_G3069_, new_G3070_, new_G3071_, new_G3072_,
    new_G3073_, new_G3074_, new_G3075_, new_G3076_, new_G3077_, new_G3078_,
    new_G3079_, new_G3080_, new_G3081_, new_G3082_, new_G3083_, new_G3084_,
    new_G3085_, new_G3086_, new_G3087_, new_G3088_, new_G3089_, new_G3090_,
    new_G3091_, new_G3092_, new_G3093_, new_G3094_, new_G3095_, new_G3096_,
    new_G3097_, new_G3098_, new_G3099_, new_G3100_, new_G3101_, new_G3102_,
    new_G3103_, new_G3104_, new_G3105_, new_G3106_, new_G3107_, new_G3108_,
    new_G3109_, new_G3110_, new_G3111_, new_G3112_, new_G3113_, new_G3114_,
    new_G3115_, new_G3116_, new_G3117_, new_G3118_, new_G3119_, new_G3120_,
    new_G3127_, new_G3128_, new_G3129_, new_G3130_, new_G3131_, new_G3132_,
    new_G3133_, new_G3134_, new_G3135_, new_G3136_, new_G3137_, new_G3138_,
    new_G3139_, new_G3140_, new_G3141_, new_G3142_, new_G3143_, new_G3144_,
    new_G3145_, new_G3146_, new_G3147_, new_G3148_, new_G3149_, new_G3150_,
    new_G3151_, new_G3152_, new_G3153_, new_G3154_, new_G3155_, new_G3156_,
    new_G3157_, new_G3158_, new_G3159_, new_G3160_, new_G3161_, new_G3162_,
    new_G3163_, new_G3164_, new_G3165_, new_G3166_, new_G3167_, new_G3168_,
    new_G3169_, new_G3170_, new_G3171_, new_G3172_, new_G3173_, new_G3174_,
    new_G3175_, new_G3176_, new_G3177_, new_G3178_, new_G3179_, new_G3180_,
    new_G3181_, new_G3182_, new_G3183_, new_G3184_, new_G3185_, new_G3186_,
    new_G3187_, new_G3194_, new_G3195_, new_G3196_, new_G3197_, new_G3198_,
    new_G3199_, new_G3200_, new_G3201_, new_G3202_, new_G3203_, new_G3204_,
    new_G3205_, new_G3206_, new_G3207_, new_G3208_, new_G3209_, new_G3210_,
    new_G3211_, new_G3212_, new_G3213_, new_G3214_, new_G3215_, new_G3216_,
    new_G3217_, new_G3218_, new_G3219_, new_G3220_, new_G3221_, new_G3222_,
    new_G3223_, new_G3224_, new_G3225_, new_G3226_, new_G3227_, new_G3228_,
    new_G3229_, new_G3230_, new_G3231_, new_G3232_, new_G3233_, new_G3234_,
    new_G3235_, new_G3236_, new_G3237_, new_G3238_, new_G3239_, new_G3240_,
    new_G3241_, new_G3242_, new_G3243_, new_G3244_, new_G3245_, new_G3246_,
    new_G3247_, new_G3248_, new_G3249_, new_G3250_, new_G3251_, new_G3252_,
    new_G3253_, new_G3254_, new_G3261_, new_G3262_, new_G3263_, new_G3264_,
    new_G3265_, new_G3266_, new_G3267_, new_G3268_, new_G3269_, new_G3270_,
    new_G3271_, new_G3272_, new_G3273_, new_G3274_, new_G3275_, new_G3276_,
    new_G3277_, new_G3278_, new_G3279_, new_G3280_, new_G3281_, new_G3282_,
    new_G3283_, new_G3284_, new_G3285_, new_G3286_, new_G3287_, new_G3288_,
    new_G3289_, new_G3290_, new_G3291_, new_G3292_, new_G3293_, new_G3294_,
    new_G3295_, new_G3296_, new_G3297_, new_G3298_, new_G3299_, new_G3300_,
    new_G3301_, new_G3302_, new_G3303_, new_G3304_, new_G3305_, new_G3306_,
    new_G3307_, new_G3308_, new_G3309_, new_G3310_, new_G3311_, new_G3312_,
    new_G3313_, new_G3314_, new_G3315_, new_G3316_, new_G3317_, new_G3318_,
    new_G3319_, new_G3320_, new_G3321_, new_G3328_, new_G3329_, new_G3330_,
    new_G3331_, new_G3332_, new_G3333_, new_G3334_, new_G3335_, new_G3336_,
    new_G3337_, new_G3338_, new_G3339_, new_G3340_, new_G3341_, new_G3342_,
    new_G3343_, new_G3344_, new_G3345_, new_G3346_, new_G3347_, new_G3348_,
    new_G3349_, new_G3350_, new_G3351_, new_G3352_, new_G3353_, new_G3354_,
    new_G3355_, new_G3356_, new_G3357_, new_G3358_, new_G3359_, new_G3360_,
    new_G3361_, new_G3362_, new_G3363_, new_G3364_, new_G3365_, new_G3366_,
    new_G3367_, new_G3368_, new_G3369_, new_G3370_, new_G3371_, new_G3372_,
    new_G3373_, new_G3374_, new_G3375_, new_G3376_, new_G3377_, new_G3378_,
    new_G3379_, new_G3380_, new_G3381_, new_G3382_, new_G3383_, new_G3384_,
    new_G3385_, new_G3386_, new_G3387_, new_G3388_, new_G3395_, new_G3396_,
    new_G3397_, new_G3398_, new_G3399_, new_G3400_, new_G3401_, new_G3402_,
    new_G3403_, new_G3404_, new_G3405_, new_G3406_, new_G3407_, new_G3408_,
    new_G3409_, new_G3410_, new_G3411_, new_G3412_, new_G3413_, new_G3414_,
    new_G3415_, new_G3416_, new_G3417_, new_G3418_, new_G3419_, new_G3420_,
    new_G3421_, new_G3422_, new_G3423_, new_G3424_, new_G3425_, new_G3426_,
    new_G3427_, new_G3428_, new_G3429_, new_G3430_, new_G3431_, new_G3432_,
    new_G3433_, new_G3434_, new_G3435_, new_G3436_, new_G3437_, new_G3438_,
    new_G3439_, new_G3440_, new_G3441_, new_G3442_, new_G3443_, new_G3444_,
    new_G3445_, new_G3446_, new_G3447_, new_G3448_, new_G3449_, new_G3450_,
    new_G3451_, new_G3452_, new_G3453_, new_G3454_, new_G3455_, new_G3462_,
    new_G3463_, new_G3464_, new_G3465_, new_G3466_, new_G3467_, new_G3468_,
    new_G3469_, new_G3470_, new_G3471_, new_G3472_, new_G3473_, new_G3474_,
    new_G3475_, new_G3476_, new_G3477_, new_G3478_, new_G3479_, new_G3480_,
    new_G3481_, new_G3482_, new_G3483_, new_G3484_, new_G3485_, new_G3486_,
    new_G3487_, new_G3488_, new_G3489_, new_G3490_, new_G3491_, new_G3492_,
    new_G3493_, new_G3494_, new_G3495_, new_G3496_, new_G3497_, new_G3498_,
    new_G3499_, new_G3500_, new_G3501_, new_G3502_, new_G3503_, new_G3504_,
    new_G3505_, new_G3506_, new_G3507_, new_G3508_, new_G3509_, new_G3510_,
    new_G3511_, new_G3512_, new_G3513_, new_G3514_, new_G3515_, new_G3516_,
    new_G3517_, new_G3518_, new_G3519_, new_G3520_, new_G3521_, new_G3522_,
    new_G3529_, new_G3530_, new_G3531_, new_G3532_, new_G3533_, new_G3534_,
    new_G3535_, new_G3536_, new_G3537_, new_G3538_, new_G3539_, new_G3540_,
    new_G3541_, new_G3542_, new_G3543_, new_G3544_, new_G3545_, new_G3546_,
    new_G3547_, new_G3548_, new_G3549_, new_G3550_, new_G3551_, new_G3552_,
    new_G3553_, new_G3554_, new_G3555_, new_G3556_, new_G3557_, new_G3558_,
    new_G3559_, new_G3560_, new_G3561_, new_G3562_, new_G3563_, new_G3564_,
    new_G3565_, new_G3566_, new_G3567_, new_G3568_, new_G3569_, new_G3570_,
    new_G3571_, new_G3572_, new_G3573_, new_G3574_, new_G3575_, new_G3576_,
    new_G3577_, new_G3578_, new_G3579_, new_G3580_, new_G3581_, new_G3582_,
    new_G3583_, new_G3584_, new_G3585_, new_G3586_, new_G3587_, new_G3588_,
    new_G3589_, new_G3596_, new_G3597_, new_G3598_, new_G3599_, new_G3600_,
    new_G3601_, new_G3602_, new_G3603_, new_G3604_, new_G3605_, new_G3606_,
    new_G3607_, new_G3608_, new_G3609_, new_G3610_, new_G3611_, new_G3612_,
    new_G3613_, new_G3614_, new_G3615_, new_G3616_, new_G3617_, new_G3618_,
    new_G3619_, new_G3620_, new_G3621_, new_G3622_, new_G3623_, new_G3624_,
    new_G3625_, new_G3626_, new_G3627_, new_G3628_, new_G3629_, new_G3630_,
    new_G3631_, new_G3632_, new_G3633_, new_G3634_, new_G3635_, new_G3636_,
    new_G3637_, new_G3638_, new_G3639_, new_G3640_, new_G3641_, new_G3642_,
    new_G3643_, new_G3644_, new_G3645_, new_G3646_, new_G3647_, new_G3648_,
    new_G3649_, new_G3650_, new_G3651_, new_G3652_, new_G3653_, new_G3654_,
    new_G3655_, new_G3656_, new_G3663_, new_G3664_, new_G3665_, new_G3666_,
    new_G3667_, new_G3668_, new_G3669_, new_G3670_, new_G3671_, new_G3672_,
    new_G3673_, new_G3674_, new_G3675_, new_G3676_, new_G3677_, new_G3678_,
    new_G3679_, new_G3680_, new_G3681_, new_G3682_, new_G3683_, new_G3684_,
    new_G3685_, new_G3686_, new_G3687_, new_G3688_, new_G3689_, new_G3690_,
    new_G3691_, new_G3692_, new_G3693_, new_G3694_, new_G3695_, new_G3696_,
    new_G3697_, new_G3698_, new_G3699_, new_G3700_, new_G3701_, new_G3702_,
    new_G3703_, new_G3704_, new_G3705_, new_G3706_, new_G3707_, new_G3708_,
    new_G3709_, new_G3710_, new_G3711_, new_G3712_, new_G3713_, new_G3714_,
    new_G3715_, new_G3716_, new_G3717_, new_G3718_, new_G3719_, new_G3720_,
    new_G3721_, new_G3722_, new_G3723_, new_G3730_, new_G3731_, new_G3732_,
    new_G3733_, new_G3734_, new_G3735_, new_G3736_, new_G3737_, new_G3738_,
    new_G3739_, new_G3740_, new_G3741_, new_G3742_, new_G3743_, new_G3744_,
    new_G3745_, new_G3746_, new_G3747_, new_G3748_, new_G3749_, new_G3750_,
    new_G3751_, new_G3752_, new_G3753_, new_G3754_, new_G3755_, new_G3756_,
    new_G3757_, new_G3758_, new_G3759_, new_G3760_, new_G3761_, new_G3762_,
    new_G3763_, new_G3764_, new_G3765_, new_G3766_, new_G3767_, new_G3768_,
    new_G3769_, new_G3770_, new_G3771_, new_G3772_, new_G3773_, new_G3774_,
    new_G3775_, new_G3776_, new_G3777_, new_G3778_, new_G3779_, new_G3780_,
    new_G3781_, new_G3782_, new_G3783_, new_G3784_, new_G3785_, new_G3786_,
    new_G3787_, new_G3788_, new_G3789_, new_G3790_, new_G3797_, new_G3798_,
    new_G3799_, new_G3800_, new_G3801_, new_G3802_, new_G3803_, new_G3804_,
    new_G3805_, new_G3806_, new_G3807_, new_G3808_, new_G3809_, new_G3810_,
    new_G3811_, new_G3812_, new_G3813_, new_G3814_, new_G3815_, new_G3816_,
    new_G3817_, new_G3818_, new_G3819_, new_G3820_, new_G3821_, new_G3822_,
    new_G3823_, new_G3824_, new_G3825_, new_G3826_, new_G3827_, new_G3828_,
    new_G3829_, new_G3830_, new_G3831_, new_G3832_, new_G3833_, new_G3834_,
    new_G3835_, new_G3836_, new_G3837_, new_G3838_, new_G3839_, new_G3840_,
    new_G3841_, new_G3842_, new_G3843_, new_G3844_, new_G3845_, new_G3846_,
    new_G3847_, new_G3848_, new_G3849_, new_G3850_, new_G3851_, new_G3852_,
    new_G3853_, new_G3854_, new_G3855_, new_G3856_, new_G3857_, new_G3864_,
    new_G3865_, new_G3866_, new_G3867_, new_G3868_, new_G3869_, new_G3870_,
    new_G3871_, new_G3872_, new_G3873_, new_G3874_, new_G3875_, new_G3876_,
    new_G3877_, new_G3878_, new_G3879_, new_G3880_, new_G3881_, new_G3882_,
    new_G3883_, new_G3884_, new_G3885_, new_G3886_, new_G3887_, new_G3888_,
    new_G3889_, new_G3890_, new_G3891_, new_G3892_, new_G3893_, new_G3894_,
    new_G3895_, new_G3896_, new_G3897_, new_G3898_, new_G3899_, new_G3900_,
    new_G3901_, new_G3902_, new_G3903_, new_G3904_, new_G3905_, new_G3906_,
    new_G3907_, new_G3908_, new_G3909_, new_G3910_, new_G3911_, new_G3912_,
    new_G3913_, new_G3914_, new_G3915_, new_G3916_, new_G3917_, new_G3918_,
    new_G3919_, new_G3920_, new_G3921_, new_G3922_, new_G3923_, new_G3924_,
    new_G3931_, new_G3932_, new_G3933_, new_G3934_, new_G3935_, new_G3936_,
    new_G3937_, new_G3938_, new_G3939_, new_G3940_, new_G3941_, new_G3942_,
    new_G3943_, new_G3944_, new_G3945_, new_G3946_, new_G3947_, new_G3948_,
    new_G3949_, new_G3950_, new_G3951_, new_G3952_, new_G3953_, new_G3954_,
    new_G3955_, new_G3956_, new_G3957_, new_G3958_, new_G3959_, new_G3960_,
    new_G3961_, new_G3962_, new_G3963_, new_G3964_, new_G3965_, new_G3966_,
    new_G3967_, new_G3968_, new_G3969_, new_G3970_, new_G3971_, new_G3972_,
    new_G3973_, new_G3974_, new_G3975_, new_G3976_, new_G3977_, new_G3978_,
    new_G3979_, new_G3980_, new_G3981_, new_G3982_, new_G3983_, new_G3984_,
    new_G3985_, new_G3986_, new_G3987_, new_G3988_, new_G3989_, new_G3990_,
    new_G3991_, new_G3998_, new_G3999_, new_G4000_, new_G4001_, new_G4002_,
    new_G4003_, new_G4004_, new_G4005_, new_G4006_, new_G4007_, new_G4008_,
    new_G4009_, new_G4010_, new_G4011_, new_G4012_, new_G4013_, new_G4014_,
    new_G4015_, new_G4016_, new_G4017_, new_G4018_, new_G4019_, new_G4020_,
    new_G4021_, new_G4022_, new_G4023_, new_G4024_, new_G4025_, new_G4026_,
    new_G4027_, new_G4028_, new_G4029_, new_G4030_, new_G4031_, new_G4032_,
    new_G4033_, new_G4034_, new_G4035_, new_G4036_, new_G4037_, new_G4038_,
    new_G4039_, new_G4040_, new_G4041_, new_G4042_, new_G4043_, new_G4044_,
    new_G4045_, new_G4046_, new_G4047_, new_G4048_, new_G4049_, new_G4050_,
    new_G4051_, new_G4052_, new_G4053_, new_G4054_, new_G4055_, new_G4056_,
    new_G4057_, new_G4058_, new_G4065_, new_G4066_, new_G4067_, new_G4068_,
    new_G4069_, new_G4070_, new_G4071_, new_G4072_, new_G4073_, new_G4074_,
    new_G4075_, new_G4076_, new_G4077_, new_G4078_, new_G4079_, new_G4080_,
    new_G4081_, new_G4082_, new_G4083_, new_G4084_, new_G4085_, new_G4086_,
    new_G4087_, new_G4088_, new_G4089_, new_G4090_, new_G4091_, new_G4092_,
    new_G4093_, new_G4094_, new_G4095_, new_G4096_, new_G4097_, new_G4098_,
    new_G4099_, new_G4100_, new_G4101_, new_G4102_, new_G4103_, new_G4104_,
    new_G4105_, new_G4106_, new_G4107_, new_G4108_, new_G4109_, new_G4110_,
    new_G4111_, new_G4112_, new_G4113_, new_G4114_, new_G4115_, new_G4116_,
    new_G4117_, new_G4118_, new_G4119_, new_G4120_, new_G4121_, new_G4122_,
    new_G4123_, new_G4124_, new_G4125_, new_G4132_, new_G4133_, new_G4134_,
    new_G4135_, new_G4136_, new_G4137_, new_G4138_, new_G4139_, new_G4140_,
    new_G4141_, new_G4142_, new_G4143_, new_G4144_, new_G4145_, new_G4146_,
    new_G4147_, new_G4148_, new_G4149_, new_G4150_, new_G4151_, new_G4152_,
    new_G4153_, new_G4154_, new_G4155_, new_G4156_, new_G4157_, new_G4158_,
    new_G4159_, new_G4160_, new_G4161_, new_G4162_, new_G4163_, new_G4164_,
    new_G4165_, new_G4166_, new_G4167_, new_G4168_, new_G4169_, new_G4170_,
    new_G4171_, new_G4172_, new_G4173_, new_G4174_, new_G4175_, new_G4176_,
    new_G4177_, new_G4178_, new_G4179_, new_G4180_, new_G4181_, new_G4182_,
    new_G4183_, new_G4184_, new_G4185_, new_G4186_, new_G4187_, new_G4188_,
    new_G4189_, new_G4190_, new_G4191_, new_G4192_, new_G4199_, new_G4200_,
    new_G4201_, new_G4202_, new_G4203_, new_G4204_, new_G4205_, new_G4206_,
    new_G4207_, new_G4208_, new_G4209_, new_G4210_, new_G4211_, new_G4212_,
    new_G4213_, new_G4214_, new_G4215_, new_G4216_, new_G4217_, new_G4218_,
    new_G4219_, new_G4220_, new_G4221_, new_G4222_, new_G4223_, new_G4224_,
    new_G4225_, new_G4226_, new_G4227_, new_G4228_, new_G4229_, new_G4230_,
    new_G4231_, new_G4232_, new_G4233_, new_G4234_, new_G4235_, new_G4236_,
    new_G4237_, new_G4238_, new_G4239_, new_G4240_, new_G4241_, new_G4242_,
    new_G4243_, new_G4244_, new_G4245_, new_G4246_, new_G4247_, new_G4248_,
    new_G4249_, new_G4250_, new_G4251_, new_G4252_, new_G4253_, new_G4254_,
    new_G4255_, new_G4256_, new_G4257_, new_G4258_, new_G4259_, new_G4266_,
    new_G4267_, new_G4268_, new_G4269_, new_G4270_, new_G4271_, new_G4272_,
    new_G4273_, new_G4274_, new_G4275_, new_G4276_, new_G4277_, new_G4278_,
    new_G4279_, new_G4280_, new_G4281_, new_G4282_, new_G4283_, new_G4284_,
    new_G4285_, new_G4286_, new_G4287_, new_G4288_, new_G4289_, new_G4290_,
    new_G4291_, new_G4292_, new_G4293_, new_G4294_, new_G4295_, new_G4296_,
    new_G4297_, new_G4298_, new_G4299_, new_G4300_, new_G4301_, new_G4302_,
    new_G4303_, new_G4304_, new_G4305_, new_G4306_, new_G4307_, new_G4308_,
    new_G4309_, new_G4310_, new_G4311_, new_G4312_, new_G4313_, new_G4314_,
    new_G4315_, new_G4316_, new_G4317_, new_G4318_, new_G4319_, new_G4320_,
    new_G4321_, new_G4322_, new_G4323_, new_G4324_, new_G4325_, new_G4326_,
    new_G4333_, new_G4334_, new_G4335_, new_G4336_, new_G4337_, new_G4338_,
    new_G4339_, new_G4340_, new_G4341_, new_G4342_, new_G4343_, new_G4344_,
    new_G4345_, new_G4346_, new_G4347_, new_G4348_, new_G4349_, new_G4350_,
    new_G4351_, new_G4352_, new_G4353_, new_G4354_, new_G4355_, new_G4356_,
    new_G4357_, new_G4358_, new_G4359_, new_G4360_, new_G4361_, new_G4362_,
    new_G4363_, new_G4364_, new_G4365_, new_G4366_, new_G4367_, new_G4368_,
    new_G4369_, new_G4370_, new_G4371_, new_G4372_, new_G4373_, new_G4374_,
    new_G4375_, new_G4376_, new_G4377_, new_G4378_, new_G4379_, new_G4380_,
    new_G4381_, new_G4382_, new_G4383_, new_G4384_, new_G4385_, new_G4386_,
    new_G4387_, new_G4388_, new_G4389_, new_G4390_, new_G4391_, new_G4392_,
    new_G4393_, new_G4400_, new_G4401_, new_G4402_, new_G4403_, new_G4404_,
    new_G4405_, new_G4406_, new_G4407_, new_G4408_, new_G4409_, new_G4410_,
    new_G4411_, new_G4412_, new_G4413_, new_G4414_, new_G4415_, new_G4416_,
    new_G4417_, new_G4418_, new_G4419_, new_G4420_, new_G4421_, new_G4422_,
    new_G4423_, new_G4424_, new_G4425_, new_G4426_, new_G4427_, new_G4428_,
    new_G4429_, new_G4430_, new_G4431_, new_G4432_, new_G4433_, new_G4434_,
    new_G4435_, new_G4436_, new_G4437_, new_G4438_, new_G4439_, new_G4440_,
    new_G4441_, new_G4442_, new_G4443_, new_G4444_, new_G4445_, new_G4446_,
    new_G4447_, new_G4448_, new_G4449_, new_G4450_, new_G4451_, new_G4452_,
    new_G4453_, new_G4454_, new_G4455_, new_G4456_, new_G4457_, new_G4458_,
    new_G4459_, new_G4460_, new_G4467_, new_G4468_, new_G4469_, new_G4470_,
    new_G4471_, new_G4472_, new_G4473_, new_G4474_, new_G4475_, new_G4476_,
    new_G4477_, new_G4478_, new_G4479_, new_G4480_, new_G4481_, new_G4482_,
    new_G4483_, new_G4484_, new_G4485_, new_G4486_, new_G4487_, new_G4488_,
    new_G4489_, new_G4490_, new_G4491_, new_G4492_, new_G4493_, new_G4494_,
    new_G4495_, new_G4496_, new_G4497_, new_G4498_, new_G4499_, new_G4500_,
    new_G4501_, new_G4502_, new_G4503_, new_G4504_, new_G4505_, new_G4506_,
    new_G4507_, new_G4508_, new_G4509_, new_G4510_, new_G4511_, new_G4512_,
    new_G4513_, new_G4514_, new_G4515_, new_G4516_, new_G4517_, new_G4518_,
    new_G4519_, new_G4520_, new_G4521_, new_G4522_, new_G4523_, new_G4524_,
    new_G4525_, new_G4526_, new_G4527_, new_G4534_, new_G4535_, new_G4536_,
    new_G4537_, new_G4538_, new_G4539_, new_G4540_, new_G4541_, new_G4542_,
    new_G4543_, new_G4544_, new_G4545_, new_G4546_, new_G4547_, new_G4548_,
    new_G4549_, new_G4550_, new_G4551_, new_G4552_, new_G4553_, new_G4554_,
    new_G4555_, new_G4556_, new_G4557_, new_G4558_, new_G4559_, new_G4560_,
    new_G4561_, new_G4562_, new_G4563_, new_G4564_, new_G4565_, new_G4566_,
    new_G4567_, new_G4568_, new_G4569_, new_G4570_, new_G4571_, new_G4572_,
    new_G4573_, new_G4574_, new_G4575_, new_G4576_, new_G4577_, new_G4578_,
    new_G4579_, new_G4580_, new_G4581_, new_G4582_, new_G4583_, new_G4584_,
    new_G4585_, new_G4586_, new_G4587_, new_G4588_, new_G4589_, new_G4590_,
    new_G4591_, new_G4592_, new_G4593_, new_G4594_, new_G4601_, new_G4602_,
    new_G4603_, new_G4604_, new_G4605_, new_G4606_, new_G4607_, new_G4608_,
    new_G4609_, new_G4610_, new_G4611_, new_G4612_, new_G4613_, new_G4614_,
    new_G4615_, new_G4616_, new_G4617_, new_G4618_, new_G4619_, new_G4620_,
    new_G4621_, new_G4622_, new_G4623_, new_G4624_, new_G4625_, new_G4626_,
    new_G4627_, new_G4628_, new_G4629_, new_G4630_, new_G4631_, new_G4632_,
    new_G4633_, new_G4634_, new_G4635_, new_G4636_, new_G4637_, new_G4638_,
    new_G4639_, new_G4640_, new_G4641_, new_G4642_, new_G4643_, new_G4644_,
    new_G4645_, new_G4646_, new_G4647_, new_G4648_, new_G4649_, new_G4650_,
    new_G4651_, new_G4652_, new_G4653_, new_G4654_, new_G4655_, new_G4656_,
    new_G4657_, new_G4658_, new_G4659_, new_G4660_, new_G4661_, new_G4668_,
    new_G4669_, new_G4670_, new_G4671_, new_G4672_, new_G4673_, new_G4674_,
    new_G4675_, new_G4676_, new_G4677_, new_G4678_, new_G4679_, new_G4680_,
    new_G4681_, new_G4682_, new_G4683_, new_G4684_, new_G4685_, new_G4686_,
    new_G4687_, new_G4688_, new_G4689_, new_G4690_, new_G4691_, new_G4692_,
    new_G4693_, new_G4694_, new_G4695_, new_G4696_, new_G4697_, new_G4698_,
    new_G4699_, new_G4700_, new_G4701_, new_G4702_, new_G4703_, new_G4704_,
    new_G4705_, new_G4706_, new_G4707_, new_G4708_, new_G4709_, new_G4710_,
    new_G4711_, new_G4712_, new_G4713_, new_G4714_, new_G4715_, new_G4716_,
    new_G4717_, new_G4718_, new_G4719_, new_G4720_, new_G4721_, new_G4722_,
    new_G4723_, new_G4724_, new_G4725_, new_G4726_, new_G4727_, new_G4728_,
    new_G4735_, new_G4736_, new_G4737_, new_G4738_, new_G4739_, new_G4740_,
    new_G4741_, new_G4742_, new_G4743_, new_G4744_, new_G4745_, new_G4746_,
    new_G4747_, new_G4748_, new_G4749_, new_G4750_, new_G4751_, new_G4752_,
    new_G4753_, new_G4754_, new_G4755_, new_G4756_, new_G4757_, new_G4758_,
    new_G4759_, new_G4760_, new_G4761_, new_G4762_, new_G4763_, new_G4764_,
    new_G4765_, new_G4766_, new_G4767_, new_G4768_, new_G4769_, new_G4770_,
    new_G4771_, new_G4772_, new_G4773_, new_G4774_, new_G4775_, new_G4776_,
    new_G4777_, new_G4778_, new_G4779_, new_G4780_, new_G4781_, new_G4782_,
    new_G4783_, new_G4784_, new_G4785_, new_G4786_, new_G4787_, new_G4788_,
    new_G4789_, new_G4790_, new_G4791_, new_G4792_, new_G4793_, new_G4794_,
    new_G4795_, new_G4802_, new_G4803_, new_G4804_, new_G4805_, new_G4806_,
    new_G4807_, new_G4808_, new_G4809_, new_G4810_, new_G4811_, new_G4812_,
    new_G4813_, new_G4814_, new_G4815_, new_G4816_, new_G4817_, new_G4818_,
    new_G4819_, new_G4820_, new_G4821_, new_G4822_, new_G4823_, new_G4824_,
    new_G4825_, new_G4826_, new_G4827_, new_G4828_, new_G4829_, new_G4830_,
    new_G4831_, new_G4832_, new_G4833_, new_G4834_, new_G4835_, new_G4836_,
    new_G4837_, new_G4838_, new_G4839_, new_G4840_, new_G4841_, new_G4842_,
    new_G4843_, new_G4844_, new_G4845_, new_G4846_, new_G4847_, new_G4848_,
    new_G4849_, new_G4850_, new_G4851_, new_G4852_, new_G4853_, new_G4854_,
    new_G4855_, new_G4856_, new_G4857_, new_G4858_, new_G4859_, new_G4860_,
    new_G4861_, new_G4862_, new_G4869_, new_G4870_, new_G4871_, new_G4872_,
    new_G4873_, new_G4874_, new_G4875_, new_G4876_, new_G4877_, new_G4878_,
    new_G4879_, new_G4880_, new_G4881_, new_G4882_, new_G4883_, new_G4884_,
    new_G4885_, new_G4886_, new_G4887_, new_G4888_, new_G4889_, new_G4890_,
    new_G4891_, new_G4892_, new_G4893_, new_G4894_, new_G4895_, new_G4896_,
    new_G4897_, new_G4898_, new_G4899_, new_G4900_, new_G4901_, new_G4902_,
    new_G4903_, new_G4904_, new_G4905_, new_G4906_, new_G4907_, new_G4908_,
    new_G4909_, new_G4910_, new_G4911_, new_G4912_, new_G4913_, new_G4914_,
    new_G4915_, new_G4916_, new_G4917_, new_G4918_, new_G4919_, new_G4920_,
    new_G4921_, new_G4922_, new_G4923_, new_G4924_, new_G4925_, new_G4926_,
    new_G4927_, new_G4928_, new_G4929_, new_G4936_, new_G4937_, new_G4938_,
    new_G4939_, new_G4940_, new_G4941_, new_G4942_, new_G4943_, new_G4944_,
    new_G4945_, new_G4946_, new_G4947_, new_G4948_, new_G4949_, new_G4950_,
    new_G4951_, new_G4952_, new_G4953_, new_G4954_, new_G4955_, new_G4956_,
    new_G4957_, new_G4958_, new_G4959_, new_G4960_, new_G4961_, new_G4962_,
    new_G4963_, new_G4964_, new_G4965_, new_G4966_, new_G4967_, new_G4968_,
    new_G4969_, new_G4970_, new_G4971_, new_G4972_, new_G4973_, new_G4974_,
    new_G4975_, new_G4976_, new_G4977_, new_G4978_, new_G4979_, new_G4980_,
    new_G4981_, new_G4982_, new_G4983_, new_G4984_, new_G4985_, new_G4986_,
    new_G4987_, new_G4988_, new_G4989_, new_G4990_, new_G4991_, new_G4992_,
    new_G4993_, new_G4994_, new_G4995_, new_G4996_, new_G5003_, new_G5004_,
    new_G5005_, new_G5006_, new_G5007_, new_G5008_, new_G5009_, new_G5010_,
    new_G5011_, new_G5012_, new_G5013_, new_G5014_, new_G5015_, new_G5016_,
    new_G5017_, new_G5018_, new_G5019_, new_G5020_, new_G5021_, new_G5022_,
    new_G5023_, new_G5024_, new_G5025_, new_G5026_, new_G5027_, new_G5028_,
    new_G5029_, new_G5030_, new_G5031_, new_G5032_, new_G5033_, new_G5034_,
    new_G5035_, new_G5036_, new_G5037_, new_G5038_, new_G5039_, new_G5040_,
    new_G5041_, new_G5042_, new_G5043_, new_G5044_, new_G5045_, new_G5046_,
    new_G5047_, new_G5048_, new_G5049_, new_G5050_, new_G5051_, new_G5052_,
    new_G5053_, new_G5054_, new_G5055_, new_G5056_, new_G5057_, new_G5058_,
    new_G5059_, new_G5060_, new_G5061_, new_G5062_, new_G5063_, new_G5070_,
    new_G5071_, new_G5072_, new_G5073_, new_G5074_, new_G5075_, new_G5076_,
    new_G5077_, new_G5078_, new_G5079_, new_G5080_, new_G5081_, new_G5082_,
    new_G5083_, new_G5084_, new_G5085_, new_G5086_, new_G5087_, new_G5088_,
    new_G5089_, new_G5090_, new_G5091_, new_G5092_, new_G5093_, new_G5094_,
    new_G5095_, new_G5096_, new_G5097_, new_G5098_, new_G5099_, new_G5100_,
    new_G5101_, new_G5102_, new_G5103_, new_G5104_, new_G5105_, new_G5106_,
    new_G5107_, new_G5108_, new_G5109_, new_G5110_, new_G5111_, new_G5112_,
    new_G5113_, new_G5114_, new_G5115_, new_G5116_, new_G5117_, new_G5118_,
    new_G5119_, new_G5120_, new_G5121_, new_G5122_, new_G5123_, new_G5124_,
    new_G5125_, new_G5126_, new_G5127_, new_G5128_, new_G5129_, new_G5130_,
    new_G5137_, new_G5138_, new_G5139_, new_G5140_, new_G5141_, new_G5142_,
    new_G5143_, new_G5144_, new_G5145_, new_G5146_, new_G5147_, new_G5148_,
    new_G5149_, new_G5150_, new_G5151_, new_G5152_, new_G5153_, new_G5154_,
    new_G5155_, new_G5156_, new_G5157_, new_G5158_, new_G5159_, new_G5160_,
    new_G5161_, new_G5162_, new_G5163_, new_G5164_, new_G5165_, new_G5166_,
    new_G5167_, new_G5168_, new_G5169_, new_G5170_, new_G5171_, new_G5172_,
    new_G5173_, new_G5174_, new_G5175_, new_G5176_, new_G5177_, new_G5178_,
    new_G5179_, new_G5180_, new_G5181_, new_G5182_, new_G5183_, new_G5184_,
    new_G5185_, new_G5186_, new_G5187_, new_G5188_, new_G5189_, new_G5190_,
    new_G5191_, new_G5192_, new_G5193_, new_G5194_, new_G5195_, new_G5196_,
    new_G5197_, new_G5204_, new_G5205_, new_G5206_, new_G5207_, new_G5208_,
    new_G5209_, new_G5210_, new_G5211_, new_G5212_, new_G5213_, new_G5214_,
    new_G5215_, new_G5216_, new_G5217_, new_G5218_, new_G5219_, new_G5220_,
    new_G5221_, new_G5222_, new_G5223_, new_G5224_, new_G5225_, new_G5226_,
    new_G5227_, new_G5228_, new_G5229_, new_G5230_, new_G5231_, new_G5232_,
    new_G5233_, new_G5234_, new_G5235_, new_G5236_, new_G5237_, new_G5238_,
    new_G5239_, new_G5240_, new_G5241_, new_G5242_, new_G5243_, new_G5244_,
    new_G5245_, new_G5246_, new_G5247_, new_G5248_, new_G5249_, new_G5250_,
    new_G5251_, new_G5252_, new_G5253_, new_G5254_, new_G5255_, new_G5256_,
    new_G5257_, new_G5258_, new_G5259_, new_G5260_, new_G5261_, new_G5262_,
    new_G5263_, new_G5264_, new_G5271_, new_G5272_, new_G5273_, new_G5274_,
    new_G5275_, new_G5276_, new_G5277_, new_G5278_, new_G5279_, new_G5280_,
    new_G5281_, new_G5282_, new_G5283_, new_G5284_, new_G5285_, new_G5286_,
    new_G5287_, new_G5288_, new_G5289_, new_G5290_, new_G5291_, new_G5292_,
    new_G5293_, new_G5294_, new_G5295_, new_G5296_, new_G5297_, new_G5298_,
    new_G5299_, new_G5300_, new_G5301_, new_G5302_, new_G5303_, new_G5304_,
    new_G5305_, new_G5306_, new_G5307_, new_G5308_, new_G5309_, new_G5310_,
    new_G5311_, new_G5312_, new_G5313_, new_G5314_, new_G5315_, new_G5316_,
    new_G5317_, new_G5318_, new_G5319_, new_G5320_, new_G5321_, new_G5322_,
    new_G5323_, new_G5324_, new_G5325_, new_G5326_, new_G5327_, new_G5328_,
    new_G5329_, new_G5330_, new_G5331_, new_G5338_, new_G5339_, new_G5340_,
    new_G5341_, new_G5342_, new_G5343_, new_G5344_, new_G5345_, new_G5346_,
    new_G5347_, new_G5348_, new_G5349_, new_G5350_, new_G5351_, new_G5352_,
    new_G5353_, new_G5354_, new_G5355_, new_G5356_, new_G5357_, new_G5358_,
    new_G5359_, new_G5360_, new_G5361_, new_G5362_, new_G5363_, new_G5364_,
    new_G5365_, new_G5366_, new_G5367_, new_G5368_, new_G5369_, new_G5370_,
    new_G5371_, new_G5372_, new_G5373_, new_G5374_, new_G5375_, new_G5376_,
    new_G5377_, new_G5378_, new_G5379_, new_G5380_, new_G5381_, new_G5382_,
    new_G5383_, new_G5384_, new_G5385_, new_G5386_, new_G5387_, new_G5388_,
    new_G5389_, new_G5390_, new_G5391_, new_G5392_, new_G5393_, new_G5394_,
    new_G5395_, new_G5396_, new_G5397_, new_G5398_, new_G5405_, new_G5406_,
    new_G5407_, new_G5408_, new_G5409_, new_G5410_, new_G5411_, new_G5412_,
    new_G5413_, new_G5414_, new_G5415_, new_G5416_, new_G5417_, new_G5418_,
    new_G5419_, new_G5420_, new_G5421_, new_G5422_, new_G5423_, new_G5424_,
    new_G5425_, new_G5426_, new_G5427_, new_G5428_, new_G5429_, new_G5430_,
    new_G5431_, new_G5432_, new_G5433_, new_G5434_, new_G5435_, new_G5436_,
    new_G5437_, new_G5438_, new_G5439_, new_G5440_, new_G5441_, new_G5442_,
    new_G5443_, new_G5444_, new_G5445_, new_G5446_, new_G5447_, new_G5448_,
    new_G5449_, new_G5450_, new_G5451_, new_G5452_, new_G5453_, new_G5454_,
    new_G5455_, new_G5456_, new_G5457_, new_G5458_, new_G5459_, new_G5460_,
    new_G5461_, new_G5462_, new_G5463_, new_G5464_, new_G5465_, new_G5472_,
    new_G5473_, new_G5474_, new_G5475_, new_G5476_, new_G5477_, new_G5478_,
    new_G5479_, new_G5480_, new_G5481_, new_G5482_, new_G5483_, new_G5484_,
    new_G5485_, new_G5486_, new_G5487_, new_G5488_, new_G5489_, new_G5490_,
    new_G5491_, new_G5492_, new_G5493_, new_G5494_, new_G5495_, new_G5496_,
    new_G5497_, new_G5498_, new_G5499_, new_G5500_, new_G5501_, new_G5502_,
    new_G5503_, new_G5504_, new_G5505_, new_G5506_, new_G5507_, new_G5508_,
    new_G5509_, new_G5510_, new_G5511_, new_G5512_, new_G5513_, new_G5514_,
    new_G5515_, new_G5516_, new_G5517_, new_G5518_, new_G5519_, new_G5520_,
    new_G5521_, new_G5522_, new_G5523_, new_G5524_, new_G5525_, new_G5526_,
    new_G5527_, new_G5528_, new_G5529_, new_G5530_, new_G5531_, new_G5532_,
    new_G5539_, new_G5540_, new_G5541_, new_G5542_, new_G5543_, new_G5544_,
    new_G5545_, new_G5546_, new_G5547_, new_G5548_, new_G5549_, new_G5550_,
    new_G5551_, new_G5552_, new_G5553_, new_G5554_, new_G5555_, new_G5556_,
    new_G5557_, new_G5558_, new_G5559_, new_G5560_, new_G5561_, new_G5562_,
    new_G5563_, new_G5564_, new_G5565_, new_G5566_, new_G5567_, new_G5568_,
    new_G5569_, new_G5570_, new_G5571_, new_G5572_, new_G5573_, new_G5574_,
    new_G5575_, new_G5576_, new_G5577_, new_G5578_, new_G5579_, new_G5580_,
    new_G5581_, new_G5582_, new_G5583_, new_G5584_, new_G5585_, new_G5586_,
    new_G5587_, new_G5588_, new_G5589_, new_G5590_, new_G5591_, new_G5592_,
    new_G5593_, new_G5594_, new_G5595_, new_G5596_, new_G5597_, new_G5598_,
    new_G5599_, new_G5606_, new_G5607_, new_G5608_, new_G5609_, new_G5610_,
    new_G5611_, new_G5612_, new_G5613_, new_G5614_, new_G5615_, new_G5616_,
    new_G5617_, new_G5618_, new_G5619_, new_G5620_, new_G5621_, new_G5622_,
    new_G5623_, new_G5624_, new_G5625_, new_G5626_, new_G5627_, new_G5628_,
    new_G5629_, new_G5630_, new_G5631_, new_G5632_, new_G5633_, new_G5634_,
    new_G5635_, new_G5636_, new_G5637_, new_G5638_, new_G5639_, new_G5640_,
    new_G5641_, new_G5642_, new_G5643_, new_G5644_, new_G5645_, new_G5646_,
    new_G5647_, new_G5648_, new_G5649_, new_G5650_, new_G5651_, new_G5652_,
    new_G5653_, new_G5654_, new_G5655_, new_G5656_, new_G5657_, new_G5658_,
    new_G5659_, new_G5660_, new_G5661_, new_G5662_, new_G5663_, new_G5664_,
    new_G5665_, new_G5666_, new_G5673_, new_G5674_, new_G5675_, new_G5676_,
    new_G5677_, new_G5678_, new_G5679_, new_G5680_, new_G5681_, new_G5682_,
    new_G5683_, new_G5684_, new_G5685_, new_G5686_, new_G5687_, new_G5688_,
    new_G5689_, new_G5690_, new_G5691_, new_G5692_, new_G5693_, new_G5694_,
    new_G5695_, new_G5696_, new_G5697_, new_G5698_, new_G5699_, new_G5700_,
    new_G5701_, new_G5702_, new_G5703_, new_G5704_, new_G5705_, new_G5706_,
    new_G5707_, new_G5708_, new_G5709_, new_G5710_, new_G5711_, new_G5712_,
    new_G5713_, new_G5714_, new_G5715_, new_G5716_, new_G5717_, new_G5718_,
    new_G5719_, new_G5720_, new_G5721_, new_G5722_, new_G5723_, new_G5724_,
    new_G5725_, new_G5726_, new_G5727_, new_G5728_, new_G5729_, new_G5730_,
    new_G5731_, new_G5732_, new_G5733_, new_G5740_, new_G5741_, new_G5742_,
    new_G5743_, new_G5744_, new_G5745_, new_G5746_, new_G5747_, new_G5748_,
    new_G5749_, new_G5750_, new_G5751_, new_G5752_, new_G5753_, new_G5754_,
    new_G5755_, new_G5756_, new_G5757_, new_G5758_, new_G5759_, new_G5760_,
    new_G5761_, new_G5762_, new_G5763_, new_G5764_, new_G5765_, new_G5766_,
    new_G5767_, new_G5768_, new_G5769_, new_G5770_, new_G5771_, new_G5772_,
    new_G5773_, new_G5774_, new_G5775_, new_G5776_, new_G5777_, new_G5778_,
    new_G5779_, new_G5780_, new_G5781_, new_G5782_, new_G5783_, new_G5784_,
    new_G5785_, new_G5786_, new_G5787_, new_G5788_, new_G5789_, new_G5790_,
    new_G5791_, new_G5792_, new_G5793_, new_G5794_, new_G5795_, new_G5796_,
    new_G5797_, new_G5798_, new_G5799_, new_G5800_, new_G5807_, new_G5808_,
    new_G5809_, new_G5810_, new_G5811_, new_G5812_, new_G5813_, new_G5814_,
    new_G5815_, new_G5816_, new_G5817_, new_G5818_, new_G5819_, new_G5820_,
    new_G5821_, new_G5822_, new_G5823_, new_G5824_, new_G5825_, new_G5826_,
    new_G5827_, new_G5828_, new_G5829_, new_G5830_, new_G5831_, new_G5832_,
    new_G5833_, new_G5834_, new_G5835_, new_G5836_, new_G5837_, new_G5838_,
    new_G5839_, new_G5840_, new_G5841_, new_G5842_, new_G5843_, new_G5844_,
    new_G5845_, new_G5846_, new_G5847_, new_G5848_, new_G5849_, new_G5850_,
    new_G5851_, new_G5852_, new_G5853_, new_G5854_, new_G5855_, new_G5856_,
    new_G5857_, new_G5858_, new_G5859_, new_G5860_, new_G5861_, new_G5862_,
    new_G5863_, new_G5864_, new_G5865_, new_G5866_, new_G5867_, new_G5874_,
    new_G5875_, new_G5876_, new_G5877_, new_G5878_, new_G5879_, new_G5880_,
    new_G5881_, new_G5882_, new_G5883_, new_G5884_, new_G5885_, new_G5886_,
    new_G5887_, new_G5888_, new_G5889_, new_G5890_, new_G5891_, new_G5892_,
    new_G5893_, new_G5894_, new_G5895_, new_G5896_, new_G5897_, new_G5898_,
    new_G5899_, new_G5900_, new_G5901_, new_G5902_, new_G5903_, new_G5904_,
    new_G5905_, new_G5906_, new_G5907_, new_G5908_, new_G5909_, new_G5910_,
    new_G5911_, new_G5912_, new_G5913_, new_G5914_, new_G5915_, new_G5916_,
    new_G5917_, new_G5918_, new_G5919_, new_G5920_, new_G5921_, new_G5922_,
    new_G5923_, new_G5924_, new_G5925_, new_G5926_, new_G5927_, new_G5928_,
    new_G5929_, new_G5930_, new_G5931_, new_G5932_, new_G5933_, new_G5934_,
    new_D7054_, new_D7053_, new_D7052_, new_D7051_, new_D7050_, new_D7049_,
    new_D7048_, new_D7047_, new_D7046_, new_D7045_, new_D7044_, new_D7043_,
    new_D7042_, new_D7041_, new_D7040_, new_D7039_, new_D7038_, new_D7037_,
    new_D7036_, new_D7035_, new_D7034_, new_D7033_, new_D7032_, new_D7031_,
    new_D7030_, new_D7029_, new_D7028_, new_D7027_, new_D7026_, new_D7025_,
    new_D7024_, new_D7023_, new_D7022_, new_D7021_, new_D7020_, new_D7019_,
    new_D7018_, new_D7017_, new_D7016_, new_D7015_, new_D7014_, new_D7013_,
    new_D7012_, new_D7011_, new_D7010_, new_D7009_, new_D7008_, new_D7007_,
    new_D7006_, new_D7005_, new_D7004_, new_D7003_, new_D7002_, new_D7001_,
    new_D7000_, new_D6999_, new_D6998_, new_D6997_, new_D6996_, new_D6995_,
    new_D6994_, new_D6993_, new_D6992_, new_D6991_, new_D6990_, new_D6989_,
    new_D6988_, new_D7055_, new_D7056_, new_D7057_, new_D7058_, new_D7059_,
    new_D7060_, new_D7061_, new_D7062_, new_D7063_, new_D7064_, new_D7065_,
    new_D7066_, new_D7067_, new_D7068_, new_D7069_, new_D7070_, new_D7071_,
    new_D7072_, new_D7073_, new_D7074_, new_D7075_, new_D7076_, new_D7077_,
    new_D7078_, new_D7079_, new_D7080_, new_D7081_, new_D7082_, new_D7083_,
    new_D7084_, new_D7085_, new_D7086_, new_D7087_, new_D7088_, new_D7089_,
    new_D7090_, new_D7091_, new_D7092_, new_D7093_, new_D7094_, new_D7095_,
    new_D7096_, new_D7097_, new_D7098_, new_D7099_, new_D7100_, new_D7101_,
    new_D7102_, new_D7103_, new_D7104_, new_D7105_, new_D7106_, new_D7107_,
    new_D7108_, new_D7109_, new_D7110_, new_D7111_, new_D7112_, new_D7113_,
    new_D7114_, new_D7115_, new_D7116_, new_D7117_, new_D7118_, new_D7119_,
    new_D7120_, new_D7121_, new_D7122_, new_D7123_, new_D7124_, new_D7125_,
    new_D7126_, new_D7127_, new_D7128_, new_D7129_, new_D7130_, new_D7131_,
    new_D7132_, new_D7133_, new_D7134_, new_D7135_, new_D7136_, new_D7137_,
    new_D7138_, new_D7139_, new_D7140_, new_D7141_, new_D7142_, new_D7143_,
    new_D7144_, new_D7145_, new_D7146_, new_D7147_, new_D7148_, new_D7149_,
    new_D7150_, new_D7151_, new_D7152_, new_D7153_, new_D7154_, new_D7155_,
    new_D7156_, new_D7157_, new_D7158_, new_D7159_, new_D7160_, new_D7161_,
    new_D7162_, new_D7163_, new_D7164_, new_D7165_, new_D7166_, new_D7167_,
    new_D7168_, new_D7169_, new_D7170_, new_D7171_, new_D7172_, new_D7173_,
    new_D7174_, new_D7175_, new_D7176_, new_D7177_, new_D7178_, new_D7179_,
    new_D7180_, new_D7181_, new_D7182_, new_D7183_, new_D7184_, new_D7185_,
    new_D7186_, new_D7187_, new_D7188_, new_D7189_, new_D7190_, new_D7191_,
    new_D7192_, new_D7193_, new_D7194_, new_D7195_, new_D7196_, new_D7197_,
    new_D7198_, new_D7199_, new_D7200_, new_D7201_, new_D7202_, new_D7203_,
    new_D7204_, new_D7205_, new_D7206_, new_D7207_, new_D7208_, new_D7209_,
    new_D7210_, new_D7211_, new_D7212_, new_D7213_, new_D7214_, new_D7215_,
    new_D7216_, new_D7217_, new_D7218_, new_D7219_, new_D7220_, new_D7221_,
    new_D7222_, new_D7223_, new_D7224_, new_D7225_, new_D7226_, new_D7227_,
    new_D7228_, new_D7229_, new_D7230_, new_D7231_, new_D7232_, new_D7233_,
    new_D7234_, new_D7235_, new_D7236_, new_D7237_, new_D7238_, new_D7239_,
    new_D7240_, new_D7241_, new_D7242_, new_D7243_, new_D7244_, new_D7245_,
    new_D7246_, new_D7247_, new_D7248_, new_D7249_, new_D7250_, new_D7251_,
    new_D7252_, new_D7253_, new_D7254_, new_D7255_, new_D7256_, new_D7257_,
    new_D7258_, new_D7259_, new_D7260_, new_D7261_, new_D7262_, new_D7263_,
    new_D7264_, new_D7265_, new_D7266_, new_D7267_, new_D7268_, new_D7269_,
    new_D7270_, new_D7271_, new_D7272_, new_D7273_, new_D7274_, new_D7275_,
    new_D7276_, new_D7277_, new_D7278_, new_D7279_, new_D7280_, new_D7281_,
    new_D7282_, new_D7283_, new_D7284_, new_D7285_, new_D7286_, new_D7287_,
    new_D7288_, new_D7289_, new_D7290_, new_D7291_, new_D7292_, new_D7293_,
    new_D7294_, new_D7295_, new_D7296_, new_D7297_, new_D7298_, new_D7299_,
    new_D7300_, new_D7301_, new_D7302_, new_D7303_, new_D7304_, new_D7305_,
    new_D7306_, new_D7307_, new_D7308_, new_D7309_, new_D7310_, new_D7311_,
    new_D7312_, new_D7313_, new_D7314_, new_D7315_, new_D7316_, new_D7317_,
    new_D7318_, new_D7319_, new_D7320_, new_D7321_, new_D7322_, new_D7323_,
    new_D7324_, new_D7325_, new_D7326_, new_D7327_, new_D7328_, new_D7329_,
    new_D7330_, new_D7331_, new_D7332_, new_D7333_, new_D7334_, new_D7335_,
    new_D7336_, new_D7337_, new_D7338_, new_D7339_, new_D7340_, new_D7341_,
    new_D7342_, new_D7343_, new_D7344_, new_D7345_, new_D7346_, new_D7347_,
    new_D7348_, new_D7349_, new_D7350_, new_D7351_, new_D7352_, new_D7353_,
    new_D7354_, new_D7355_, new_D7356_, new_D7357_, new_D7358_, new_D7359_,
    new_D7360_, new_D7361_, new_D7362_, new_D7363_, new_D7364_, new_D7365_,
    new_D7366_, new_D7367_, new_D7368_, new_D7369_, new_D7370_, new_D7371_,
    new_D7372_, new_D7373_, new_D7374_, new_D7375_, new_D7376_, new_D7377_,
    new_D7378_, new_D7379_, new_D7380_, new_D7381_, new_D7382_, new_D7383_,
    new_D7384_, new_D7385_, new_D7386_, new_D7387_, new_D7388_, new_D7389_,
    new_D7390_, new_D7391_, new_D7392_, new_D7393_, new_D7394_, new_D7395_,
    new_D7396_, new_D7397_, new_D7398_, new_D7399_, new_D7400_, new_D7401_,
    new_D7402_, new_D7403_, new_D7404_, new_D7405_, new_D7406_, new_D7407_,
    new_D7408_, new_D7409_, new_D7410_, new_D7411_, new_D7412_, new_D7413_,
    new_D7414_, new_D7415_, new_D7416_, new_D7417_, new_D7418_, new_D7419_,
    new_D7420_, new_D7421_, new_D7422_, new_D7423_, new_D7424_, new_D7425_,
    new_D7426_, new_D7427_, new_D7428_, new_D7429_, new_D7430_, new_D7431_,
    new_D7432_, new_D7433_, new_D7434_, new_D7435_, new_D7436_, new_D7437_,
    new_D7438_, new_D7439_, new_D7440_, new_D7441_, new_D7442_, new_D7443_,
    new_D7444_, new_D7445_, new_D7446_, new_D7447_, new_D7448_, new_D7449_,
    new_D7450_, new_D7451_, new_D7452_, new_D7453_, new_D7454_, new_D7455_,
    new_D7456_, new_D7457_, new_D7458_, new_D7459_, new_D7460_, new_D7461_,
    new_D7462_, new_D7463_, new_D7464_, new_D7465_, new_D7466_, new_D7467_,
    new_D7468_, new_D7469_, new_D7470_, new_D7471_, new_D7472_, new_D7473_,
    new_D7474_, new_D7475_, new_D7476_, new_D7477_, new_D7478_, new_D7479_,
    new_D7480_, new_D7481_, new_D7482_, new_D7483_, new_D7484_, new_D7485_,
    new_D7486_, new_D7487_, new_D7488_, new_D7489_, new_D7490_, new_D7491_,
    new_D7492_, new_D7493_, new_D7494_, new_D7495_, new_D7496_, new_D7497_,
    new_D7498_, new_D7499_, new_D7500_, new_D7501_, new_D7502_, new_D7503_,
    new_D7504_, new_D7505_, new_D7506_, new_D7507_, new_D7508_, new_D7509_,
    new_D7510_, new_D7511_, new_D7512_, new_D7513_, new_D7514_, new_D7515_,
    new_D7516_, new_D7517_, new_D7518_, new_D7519_, new_D7520_, new_D7521_,
    new_D7522_, new_D7523_, new_D7524_, new_D7525_, new_D7526_, new_D7527_,
    new_D7528_, new_D7529_, new_D7530_, new_D7531_, new_D7532_, new_D7533_,
    new_D7534_, new_D7535_, new_D7536_, new_D7537_, new_D7538_, new_D7539_,
    new_D7540_, new_D7541_, new_D7542_, new_D7543_, new_D7544_, new_D7545_,
    new_D7546_, new_D7547_, new_D7548_, new_D7549_, new_D7550_, new_D7551_,
    new_D7552_, new_D7553_, new_D7554_, new_D7555_, new_D7556_, new_D7557_,
    new_D7558_, new_D7559_, new_D7560_, new_D7561_, new_D7562_, new_D7563_,
    new_D7564_, new_D7565_, new_D7566_, new_D7567_, new_D7568_, new_D7569_,
    new_D7570_, new_D7571_, new_D7572_, new_D7573_, new_D7574_, new_D7575_,
    new_D7576_, new_D7577_, new_D7578_, new_D7579_, new_D7580_, new_D7581_,
    new_D7582_, new_D7583_, new_D7584_, new_D7585_, new_D7586_, new_D7587_,
    new_D7588_, new_D7589_, new_D7590_, new_D7591_, new_D7592_, new_D7593_,
    new_D7594_, new_D7595_, new_D7596_, new_D7597_, new_D7598_, new_D7599_,
    new_D7600_, new_D7601_, new_D7602_, new_D7603_, new_D7604_, new_D7605_,
    new_D7606_, new_D7607_, new_D7608_, new_D7609_, new_D7610_, new_D7611_,
    new_D7612_, new_D7613_, new_D7614_, new_D7615_, new_D7616_, new_D7617_,
    new_D7618_, new_D7619_, new_D7620_, new_D7621_, new_D7622_, new_D7623_,
    new_D7624_, new_D7625_, new_D7626_, new_D7627_, new_D7628_, new_D7629_,
    new_D7630_, new_D7631_, new_D7632_, new_D7633_, new_D7634_, new_D7635_,
    new_D7636_, new_D7637_, new_D7638_, new_D7639_, new_D7640_, new_D7641_,
    new_D7642_, new_D7643_, new_D7644_, new_D7645_, new_D7646_, new_D7647_,
    new_D7648_, new_D7649_, new_D7650_, new_D7651_, new_D7652_, new_D7653_,
    new_D7654_, new_D7655_, new_D7656_, new_D7657_, new_D7658_, new_D7659_,
    new_D7660_, new_D7661_, new_D7662_, new_D7663_, new_D7664_, new_D7665_,
    new_D7666_, new_D7667_, new_D7668_, new_D7669_, new_D7670_, new_D7671_,
    new_D7672_, new_D7673_, new_D7674_, new_D7675_, new_D7676_, new_D7677_,
    new_D7678_, new_D7679_, new_D7680_, new_D7681_, new_D7682_, new_D7683_,
    new_D7684_, new_D7685_, new_D7686_, new_D7687_, new_D7688_, new_D7689_,
    new_D7690_, new_D7691_, new_D7692_, new_D7693_, new_D7694_, new_D7695_,
    new_D7696_, new_D7697_, new_D7698_, new_D7699_, new_D7700_, new_D7701_,
    new_D7702_, new_D7703_, new_D7704_, new_D7705_, new_D7706_, new_D7707_,
    new_D7708_, new_D7709_, new_D7710_, new_D7711_, new_D7712_, new_D7713_,
    new_D7714_, new_D7715_, new_D7716_, new_D7717_, new_D7718_, new_D7719_,
    new_D7720_, new_D7721_, new_D7722_, new_D7723_, new_D7724_, new_D7725_,
    new_D7726_, new_D7727_, new_D7728_, new_D7729_, new_D7730_, new_D7731_,
    new_D7732_, new_D7733_, new_D7734_, new_D7735_, new_D7736_, new_D7737_,
    new_D7738_, new_D7739_, new_D7740_, new_D7741_, new_D7742_, new_D7743_,
    new_D7744_, new_D7745_, new_D7746_, new_D7747_, new_D7748_, new_D7749_,
    new_D7750_, new_D7751_, new_D7752_, new_D7753_, new_D7754_, new_D7755_,
    new_D7756_, new_D7757_, new_D7758_, new_D7759_, new_D7760_, new_D7761_,
    new_D7762_, new_D7763_, new_D7764_, new_D7765_, new_D7766_, new_D7767_,
    new_D7768_, new_D7769_, new_D7770_, new_D7771_, new_D7772_, new_D7773_,
    new_D7774_, new_D7775_, new_D7776_, new_D7777_, new_D7778_, new_D7779_,
    new_D7780_, new_D7781_, new_D7782_, new_D7783_, new_D7784_, new_D7785_,
    new_D7786_, new_D7787_, new_D7788_, new_D7789_, new_D7790_, new_D7791_,
    new_D7792_, new_D7793_, new_D7794_, new_D7795_, new_D7796_, new_D7797_,
    new_D7798_, new_D7799_, new_D7800_, new_D7801_, new_D7802_, new_D7803_,
    new_D7804_, new_D7805_, new_D7806_, new_D7807_, new_D7808_, new_D7809_,
    new_D7810_, new_D7811_, new_D7812_, new_D7813_, new_D7814_, new_D7815_,
    new_D7816_, new_D7817_, new_D7818_, new_D7819_, new_D7820_, new_D7821_,
    new_D7822_, new_D7823_, new_D7824_, new_D7825_, new_D7826_, new_D7827_,
    new_D7828_, new_D7829_, new_D7830_, new_D7831_, new_D7832_, new_D7833_,
    new_D7834_, new_D7835_, new_D7836_, new_D7837_, new_D7838_, new_D7839_,
    new_D7840_, new_D7841_, new_D7842_, new_D7843_, new_D7844_, new_D7845_,
    new_D7846_, new_D7847_, new_D7848_, new_D7849_, new_D7850_, new_D7851_,
    new_D7852_, new_D7853_, new_D7854_, new_D7855_, new_D7856_, new_D7857_,
    new_D7858_, new_D7859_, new_D7860_, new_D7861_, new_D7862_, new_D7863_,
    new_D7864_, new_D7865_, new_D7866_, new_D7867_, new_D7868_, new_D7869_,
    new_D7870_, new_D7871_, new_D7872_, new_D7873_, new_D7874_, new_D7875_,
    new_D7876_, new_D7877_, new_D7878_, new_D7879_, new_D7880_, new_D7881_,
    new_D7882_, new_D7883_, new_D7884_, new_D7885_, new_D7886_, new_D7887_,
    new_D7888_, new_D7889_, new_D7890_, new_D7891_, new_D7892_, new_D7893_,
    new_D7894_, new_D7895_, new_D7896_, new_D7897_, new_D7898_, new_D7899_,
    new_D7900_, new_D7901_, new_D7902_, new_D7903_, new_D7904_, new_D7905_,
    new_D7906_, new_D7907_, new_D7908_, new_D7909_, new_D7910_, new_D7911_,
    new_D7912_, new_D7913_, new_D7914_, new_D7915_, new_D7916_, new_D7917_,
    new_D7918_, new_D7919_, new_D7920_, new_D7921_, new_D7922_, new_D7923_,
    new_D7924_, new_D7925_, new_D7926_, new_D7927_, new_D7928_, new_D7929_,
    new_D7930_, new_D7931_, new_D7932_, new_D7933_, new_D7934_, new_D7935_,
    new_D7936_, new_D7937_, new_D7938_, new_D7939_, new_D7940_, new_D7941_,
    new_D7942_, new_D7943_, new_D7944_, new_D7945_, new_D7946_, new_D7947_,
    new_D7948_, new_D7949_, new_D7950_, new_D7951_, new_D7952_, new_D7953_,
    new_D7954_, new_D7955_, new_D7956_, new_D7957_, new_D7958_, new_D7959_,
    new_D7960_, new_D7961_, new_D7962_, new_D7963_, new_D7964_, new_D7965_,
    new_D7966_, new_D7967_, new_D7968_, new_D7969_, new_D7970_, new_D7971_,
    new_D7972_, new_D7973_, new_D7974_, new_D7975_, new_D7976_, new_D7977_,
    new_D7978_, new_D7979_, new_D7980_, new_D7981_, new_D7982_, new_D7983_,
    new_D7984_, new_D7985_, new_D7986_, new_D7987_, new_D7988_, new_D7989_,
    new_D7990_, new_D7991_, new_D7992_, new_D7993_, new_D7994_, new_D7995_,
    new_D7996_, new_D7997_, new_D7998_, new_D7999_, new_D8000_, new_D8001_,
    new_D8002_, new_D8003_, new_D8004_, new_D8005_, new_D8006_, new_D8007_,
    new_D8008_, new_D8009_, new_D8010_, new_D8011_, new_D8012_, new_D8013_,
    new_D8014_, new_D8015_, new_D8016_, new_D8017_, new_D8018_, new_D8019_,
    new_D8020_, new_D8021_, new_D8022_, new_D8023_, new_D8024_, new_D8025_,
    new_D8026_, new_D8027_, new_D8028_, new_D8029_, new_D8030_, new_D8031_,
    new_D8032_, new_D8033_, new_D8034_, new_D8035_, new_D8036_, new_D8037_,
    new_D8038_, new_D8039_, new_D8040_, new_D8041_, new_D8042_, new_D8043_,
    new_D8044_, new_D8045_, new_D8046_, new_D8047_, new_D8048_, new_D8049_,
    new_D8050_, new_D8051_, new_D8052_, new_D8053_, new_D8054_, new_D8055_,
    new_D8056_, new_D8057_, new_D8058_, new_D8059_, new_D8060_, new_D8061_,
    new_D8062_, new_D8063_, new_D8064_, new_D8065_, new_D8066_, new_D8067_,
    new_D8068_, new_D8069_, new_D8070_, new_D8071_, new_D8072_, new_D8073_,
    new_D8074_, new_D8075_, new_D8076_, new_D8077_, new_D8078_, new_D8079_,
    new_D8080_, new_D8081_, new_D8082_, new_D8083_, new_D8084_, new_D8085_,
    new_D8086_, new_D8087_, new_D8088_, new_D8089_, new_D8090_, new_D8091_,
    new_D8092_, new_D8093_, new_D8094_, new_D8095_, new_D8096_, new_D8097_,
    new_D8098_, new_D8099_, new_D8100_, new_D8101_, new_D8102_, new_D8103_,
    new_D8104_, new_D8105_, new_D8106_, new_D8107_, new_D8108_, new_D8109_,
    new_D8110_, new_D8111_, new_D8112_, new_D8113_, new_D8114_, new_D8115_,
    new_D8116_, new_D8117_, new_D8118_, new_D8119_, new_D8120_, new_D8121_,
    new_D8122_, new_D8123_, new_D8124_, new_D8125_, new_D8126_, new_D8127_,
    new_D8128_, new_D8129_, new_D8130_, new_D8131_, new_D8132_, new_D8133_,
    new_D8134_, new_D8135_, new_D8136_, new_D8137_, new_D8138_, new_D8139_,
    new_D8140_, new_D8141_, new_D8142_, new_D8143_, new_D8144_, new_D8145_,
    new_D8146_, new_D8147_, new_D8148_, new_D8149_, new_D8150_, new_D8151_,
    new_D8152_, new_D8153_, new_D8154_, new_D8155_, new_D8156_, new_D8157_,
    new_D8158_, new_D8159_, new_D8160_, new_D8161_, new_D8162_, new_D8163_,
    new_D8164_, new_D8165_, new_D8166_, new_D8167_, new_D8168_, new_D8169_,
    new_D8170_, new_D8171_, new_D8172_, new_D8173_, new_D8174_, new_D8175_,
    new_D8176_, new_D8177_, new_D8178_, new_D8179_, new_D8180_, new_D8181_,
    new_D8182_, new_D8183_, new_D8184_, new_D8185_, new_D8186_, new_D8187_,
    new_D8188_, new_D8189_, new_D8190_, new_D8191_, new_D8192_, new_D8193_,
    new_D8194_, new_D8195_, new_D8196_, new_D8197_, new_D8198_, new_D8199_,
    new_D8200_, new_D8201_, new_D8202_, new_D8203_, new_D8204_, new_D8205_,
    new_D8206_, new_D8207_, new_D8208_, new_D8209_, new_D8210_, new_D8211_,
    new_D8212_, new_D8213_, new_D8214_, new_D8215_, new_D8216_, new_D8217_,
    new_D8218_, new_D8219_, new_D8220_, new_D8221_, new_D8222_, new_D8223_,
    new_D8224_, new_D8225_, new_D8226_, new_D8227_, new_D8228_, new_D8229_,
    new_D8230_, new_D8231_, new_D8232_, new_D8233_, new_D8234_, new_D8235_,
    new_D8236_, new_D8237_, new_D8238_, new_D8239_, new_D8240_, new_D8241_,
    new_D8242_, new_D8243_, new_D8244_, new_D8245_, new_D8246_, new_D8247_,
    new_D8248_, new_D8249_, new_D8250_, new_D8251_, new_D8252_, new_D8253_,
    new_D8254_, new_D8255_, new_D8256_, new_D8257_, new_D8258_, new_D8259_,
    new_D8260_, new_D8261_, new_D8262_, new_D8263_, new_D8264_, new_D8265_,
    new_D8266_, new_D8267_, new_D8268_, new_D8269_, new_D8270_, new_D8271_,
    new_D8272_, new_D8273_, new_D8274_, new_D8275_, new_D8276_, new_D8277_,
    new_D8278_, new_D8279_, new_D8280_, new_D8281_, new_D8282_, new_D8283_,
    new_D8284_, new_D8285_, new_D8286_, new_D8287_, new_D8288_, new_D8289_,
    new_D8290_, new_D8291_, new_D8292_, new_D8293_, new_D8294_, new_D8295_,
    new_D8296_, new_D8297_, new_D8298_, new_D8299_, new_D8300_, new_D8301_,
    new_D8302_, new_D8303_, new_D8304_, new_D8305_, new_D8306_, new_D8307_,
    new_D8308_, new_D8309_, new_D8310_, new_D8311_, new_D8312_, new_D8313_,
    new_D8314_, new_D8315_, new_D8316_, new_D8317_, new_D8318_, new_D8319_,
    new_D8320_, new_D8321_, new_D8322_, new_D8323_, new_D8324_, new_D8325_,
    new_D8326_, new_D8327_, new_D8328_, new_D8329_, new_D8330_, new_D8331_,
    new_D8332_, new_D8333_, new_D8334_, new_D8335_, new_D8336_, new_D8337_,
    new_D8338_, new_D8339_, new_D8340_, new_D8341_, new_D8342_, new_D8343_,
    new_D8344_, new_D8345_, new_D8346_, new_D8347_, new_D8348_, new_D8349_,
    new_D8350_, new_D8351_, new_D8352_, new_D8353_, new_D8354_, new_D8355_,
    new_D8356_, new_D8357_, new_D8358_, new_D8359_, new_D8360_, new_D8361_,
    new_D8362_, new_D8363_, new_D8364_, new_D8365_, new_D8366_, new_D8367_,
    new_D8368_, new_D8369_, new_D8370_, new_D8371_, new_D8372_, new_D8373_,
    new_D8374_, new_D8375_, new_D8376_, new_D8377_, new_D8378_, new_D8379_,
    new_D8380_, new_D8381_, new_D8382_, new_D8383_, new_D8384_, new_D8385_,
    new_D8386_, new_D8387_, new_D8388_, new_D8389_, new_D8390_, new_D8391_,
    new_D8392_, new_D8393_, new_D8394_, new_D8395_, new_D8396_, new_D8397_,
    new_D8398_, new_D8399_, new_D8400_, new_D8401_, new_D8402_, new_D8403_,
    new_D8404_, new_D8405_, new_D8406_, new_D8407_, new_D8408_, new_D8409_,
    new_D8410_, new_D8411_, new_D8412_, new_D8413_, new_D8414_, new_D8415_,
    new_D8416_, new_D8417_, new_D8418_, new_D8419_, new_D8420_, new_D8421_,
    new_D8422_, new_D8423_, new_D8424_, new_D8425_, new_D8426_, new_D8427_,
    new_D8428_, new_D8429_, new_D8430_, new_D8431_, new_D8432_, new_D8433_,
    new_D8434_, new_D8435_, new_D8436_, new_D8437_, new_D8438_, new_D8439_,
    new_D8440_, new_D8441_, new_D8442_, new_D8443_, new_D8444_, new_D8445_,
    new_D8446_, new_D8447_, new_D8448_, new_D8449_, new_D8450_, new_D8451_,
    new_D8452_, new_D8453_, new_D8454_, new_D8455_, new_D8456_, new_D8457_,
    new_D8458_, new_D8459_, new_D8460_, new_D8461_, new_D8462_, new_D8463_,
    new_D8464_, new_D8465_, new_D8466_, new_D8467_, new_D8468_, new_D8469_,
    new_D8470_, new_D8471_, new_D8472_, new_D8473_, new_D8474_, new_D8475_,
    new_D8476_, new_D8477_, new_D8478_, new_D8479_, new_D8480_, new_D8481_,
    new_D8482_, new_D8483_, new_D8484_, new_D8485_, new_D8486_, new_D8487_,
    new_D8488_, new_D8489_, new_D8490_, new_D8491_, new_D8492_, new_D8493_,
    new_D8494_, new_D8495_, new_D8496_, new_D8497_, new_D8498_, new_D8499_,
    new_D8500_, new_D8501_, new_D8502_, new_D8503_, new_D8504_, new_D8505_,
    new_D8506_, new_D8507_, new_D8508_, new_D8509_, new_D8510_, new_D8511_,
    new_D8512_, new_D8513_, new_D8514_, new_D8515_, new_D8516_, new_D8517_,
    new_D8518_, new_D8519_, new_D8520_, new_D8521_, new_D8522_, new_D8523_,
    new_D8524_, new_D8525_, new_D8526_, new_D8527_, new_D8528_, new_D8529_,
    new_D8530_, new_D8531_, new_D8532_, new_D8533_, new_D8534_, new_D8535_,
    new_D8536_, new_D8537_, new_D8538_, new_D8539_, new_D8540_, new_D8541_,
    new_D8542_, new_D8543_, new_D8544_, new_D8545_, new_D8546_, new_D8547_,
    new_D8548_, new_D8549_, new_D8550_, new_D8551_, new_D8552_, new_D8553_,
    new_D8554_, new_D8555_, new_D8556_, new_D8557_, new_D8558_, new_D8559_,
    new_D8560_, new_D8561_, new_D8562_, new_D8563_, new_D8564_, new_D8565_,
    new_D8566_, new_D8567_, new_D8568_, new_D8569_, new_D8570_, new_D8571_,
    new_D8572_, new_D8573_, new_D8574_, new_D8575_, new_D8576_, new_D8577_,
    new_D8578_, new_D8579_, new_D8580_, new_D8581_, new_D8582_, new_D8583_,
    new_D8584_, new_D8585_, new_D8586_, new_D8587_, new_D8588_, new_D8589_,
    new_D8590_, new_D8591_, new_D8592_, new_D8593_, new_D8594_, new_D8595_,
    new_D8596_, new_D8597_, new_D8598_, new_D8599_, new_D8600_, new_D8601_,
    new_D8602_, new_D8603_, new_D8604_, new_D8605_, new_D8606_, new_D8607_,
    new_D8608_, new_D8609_, new_D8610_, new_D8611_, new_D8612_, new_D8613_,
    new_D8614_, new_D8615_, new_D8616_, new_D8617_, new_D8618_, new_D8619_,
    new_D8620_, new_D8621_, new_D8622_, new_D8623_, new_D8624_, new_D8625_,
    new_D8626_, new_D8627_, new_D8628_, new_D8629_, new_D8630_, new_D8631_,
    new_D8632_, new_D8633_, new_D8634_, new_D8635_, new_D8636_, new_D8637_,
    new_D8638_, new_D8639_, new_D8640_, new_D8641_, new_D8642_, new_D8643_,
    new_D8644_, new_D8645_, new_D8646_, new_D8647_, new_D8648_, new_D8649_,
    new_D8650_, new_D8651_, new_D8652_, new_D8653_, new_D8654_, new_D8655_,
    new_D8656_, new_D8657_, new_D8658_, new_D8659_, new_D8660_, new_D8661_,
    new_D8662_, new_D8663_, new_D8664_, new_D8665_, new_D8666_, new_D8667_,
    new_D8668_, new_D8669_, new_D8670_, new_D8671_, new_D8672_, new_D8673_,
    new_D8674_, new_D8675_, new_D8676_, new_D8677_, new_D8678_, new_D8679_,
    new_D8680_, new_D8681_, new_D8682_, new_D8683_, new_D8684_, new_D8685_,
    new_D8686_, new_D8687_, new_D8688_, new_D8689_, new_D8690_, new_D8691_,
    new_D8692_, new_D8693_, new_D8694_, new_D8695_, new_D8696_, new_D8697_,
    new_D8698_, new_D8699_, new_D8700_, new_D8701_, new_D8702_, new_D8703_,
    new_D8704_, new_D8705_, new_D8706_, new_D8707_, new_D8708_, new_D8709_,
    new_D8710_, new_D8711_, new_D8712_, new_D8713_, new_D8714_, new_D8715_,
    new_D8716_, new_D8717_, new_D8718_, new_D8719_, new_D8720_, new_D8721_,
    new_D8722_, new_D8723_, new_D8724_, new_D8725_, new_D8726_, new_D8727_,
    new_D8728_, new_D8729_, new_D8730_, new_D8731_, new_D8732_, new_D8733_,
    new_D8734_, new_D8735_, new_D8736_, new_D8737_, new_D8738_, new_D8739_,
    new_D8740_, new_D8741_, new_D8742_, new_D8743_, new_D8744_, new_D8745_,
    new_D8746_, new_D8747_, new_D8748_, new_D8749_, new_D8750_, new_D8751_,
    new_D8752_, new_D8753_, new_D8754_, new_D8755_, new_D8756_, new_D8757_,
    new_D8758_, new_D8759_, new_D8760_, new_D8761_, new_D8762_, new_D8763_,
    new_D8764_, new_D8765_, new_D8766_, new_D8767_, new_D8768_, new_D8769_,
    new_D8770_, new_D8771_, new_D8772_, new_D8773_, new_D8774_, new_D8775_,
    new_D8776_, new_D8777_, new_D8778_, new_D8779_, new_D8780_, new_D8781_,
    new_D8782_, new_D8783_, new_D8784_, new_D8785_, new_D8786_, new_D8787_,
    new_D8788_, new_D8789_, new_D8790_, new_D8791_, new_D8792_, new_D8793_,
    new_D8794_, new_D8795_, new_D8796_, new_D8797_, new_D8798_, new_D8799_,
    new_D8800_, new_D8801_, new_D8802_, new_D8803_, new_D8804_, new_D8805_,
    new_D8806_, new_D8807_, new_D8808_, new_D8809_, new_D8810_, new_D8811_,
    new_D8812_, new_D8813_, new_D8814_, new_D8815_, new_D8816_, new_D8817_,
    new_D8818_, new_D8819_, new_D8820_, new_D8821_, new_D8822_, new_D8823_,
    new_D8824_, new_D8825_, new_D8826_, new_D8827_, new_D8828_, new_D8829_,
    new_D8830_, new_D8831_, new_D8832_, new_D8833_, new_D8834_, new_D8835_,
    new_D8836_, new_D8837_, new_D8838_, new_D8839_, new_D8840_, new_D8841_,
    new_D8842_, new_D8843_, new_D8844_, new_D8845_, new_D8846_, new_D8847_,
    new_D8848_, new_D8849_, new_D8850_, new_D8851_, new_D8852_, new_D8853_,
    new_D8854_, new_D8855_, new_D8856_, new_D8857_, new_D8858_, new_D8859_,
    new_D8860_, new_D8861_, new_D8862_, new_D8863_, new_D8864_, new_D8865_,
    new_D8866_, new_D8867_, new_D8868_, new_D8869_, new_D8870_, new_D8871_,
    new_D8872_, new_D8873_, new_D8874_, new_D8875_, new_D8876_, new_D8877_,
    new_D8878_, new_D8879_, new_D8880_, new_D8881_, new_D8882_, new_D8883_,
    new_D8884_, new_D8885_, new_D8886_, new_D8887_, new_D8888_, new_D8889_,
    new_D8890_, new_D8891_, new_D8892_, new_D8893_, new_D8894_, new_D8895_,
    new_D8896_, new_D8897_, new_D8898_, new_D8899_, new_D8900_, new_D8901_,
    new_D8902_, new_D8903_, new_D8904_, new_D8905_, new_D8906_, new_D8907_,
    new_D8908_, new_D8909_, new_D8910_, new_D8911_, new_D8912_, new_D8913_,
    new_D8914_, new_D8915_, new_D8916_, new_D8917_, new_D8918_, new_D8919_,
    new_D8920_, new_D8921_, new_D8922_, new_D8923_, new_D8924_, new_D8925_,
    new_D8926_, new_D8927_, new_D8928_, new_D8929_, new_D8930_, new_D8931_,
    new_D8932_, new_D8933_, new_D8934_, new_D8935_, new_D8936_, new_D8937_,
    new_D8938_, new_D8939_, new_D8940_, new_D8941_, new_D8942_, new_D8943_,
    new_D8944_, new_D8945_, new_D8946_, new_D8947_, new_D8948_, new_D8949_,
    new_D8950_, new_D8951_, new_D8952_, new_D8953_, new_D8954_, new_D8955_,
    new_D8956_, new_D8957_, new_D8958_, new_D8959_, new_D8960_, new_D8961_,
    new_D8962_, new_D8963_, new_D8964_, new_D8965_, new_D8966_, new_D8967_,
    new_D8968_, new_D8969_, new_D8970_, new_D8971_, new_D8972_, new_D8973_,
    new_D8974_, new_D8975_, new_D8976_, new_D8977_, new_D8978_, new_D8979_,
    new_D8980_, new_D8981_, new_D8982_, new_D8983_, new_D8984_, new_D8985_,
    new_D8986_, new_D8987_, new_D8988_, new_D8989_, new_D8990_, new_D8991_,
    new_D8992_, new_D8993_, new_D8994_, new_D8995_, new_D8996_, new_D8997_,
    new_D8998_, new_D8999_, new_D9000_, new_D9001_, new_D9002_, new_D9003_,
    new_D9004_, new_D9005_, new_D9006_, new_D9007_, new_D9008_, new_D9009_,
    new_D9010_, new_D9011_, new_D9012_, new_D9013_, new_D9014_, new_D9015_,
    new_D9016_, new_D9017_, new_D9018_, new_D9019_, new_D9020_, new_D9021_,
    new_D9022_, new_D9023_, new_D9024_, new_D9025_, new_D9026_, new_D9027_,
    new_D9028_, new_D9029_, new_D9030_, new_D9031_, new_D9032_, new_D9033_,
    new_D9034_, new_D9035_, new_D9036_, new_D9037_, new_D9038_, new_D9039_,
    new_D9040_, new_D9041_, new_D9042_, new_D9043_, new_D9044_, new_D9045_,
    new_D9046_, new_D9047_, new_D9048_, new_D9049_, new_D9050_, new_D9051_,
    new_D9052_, new_D9053_, new_D9054_, new_D9055_, new_D9056_, new_D9057_,
    new_D9058_, new_D9059_, new_D9060_, new_D9061_, new_D9062_, new_D9063_,
    new_D9064_, new_D9065_, new_D9066_, new_D9067_, new_D9068_, new_D9069_,
    new_D9070_, new_D9071_, new_D9072_, new_D9073_, new_D9074_, new_D9075_,
    new_D9076_, new_D9077_, new_D9078_, new_D9079_, new_D9080_, new_D9081_,
    new_D9082_, new_D9083_, new_D9084_, new_D9085_, new_D9086_, new_D9087_,
    new_D9088_, new_D9089_, new_D9090_, new_D9091_, new_D9092_, new_D9093_,
    new_D9094_, new_D9095_, new_D9096_, new_D9097_, new_D9098_, new_D9099_,
    new_D9100_, new_D9101_, new_D9102_, new_D9103_, new_D9104_, new_D9105_,
    new_D9106_, new_D9107_, new_D9108_, new_D9109_, new_D9110_, new_D9111_,
    new_D9112_, new_D9113_, new_D9114_, new_D9115_, new_D9116_, new_D9117_,
    new_D9118_, new_D9119_, new_D9120_, new_D9121_, new_D9122_, new_D9123_,
    new_D9124_, new_D9125_, new_D9126_, new_D9127_, new_D9128_, new_D9129_,
    new_D9130_, new_D9131_, new_D9132_, new_D9133_, new_D9134_, new_D9135_,
    new_D9136_, new_D9137_, new_D9138_, new_D9139_, new_D9140_, new_D9141_,
    new_D9142_, new_D9143_, new_D9144_, new_D9145_, new_D9146_, new_D9147_,
    new_D9148_, new_D9149_, new_D9150_, new_D9151_, new_D9152_, new_D9153_,
    new_D9154_, new_D9155_, new_D9156_, new_D9157_, new_D9158_, new_D9159_,
    new_D9160_, new_D9161_, new_D9162_, new_D9163_, new_D9164_, new_D9165_,
    new_D9166_, new_D9167_, new_D9168_, new_D9169_, new_D9170_, new_D9171_,
    new_D9172_, new_D9173_, new_D9174_, new_D9175_, new_D9176_, new_D9177_,
    new_D9178_, new_D9179_, new_D9180_, new_D9181_, new_D9182_, new_D9183_,
    new_D9184_, new_D9185_, new_D9186_, new_D9187_, new_D9188_, new_D9189_,
    new_D9190_, new_D9191_, new_D9192_, new_D9193_, new_D9194_, new_D9195_,
    new_D9196_, new_D9197_, new_D9198_, new_D9199_, new_D9200_, new_D9201_,
    new_D9202_, new_D9203_, new_D9204_, new_D9205_, new_D9206_, new_D9207_,
    new_D9208_, new_D9209_, new_D9210_, new_D9211_, new_D9212_, new_D9213_,
    new_D9214_, new_D9215_, new_D9216_, new_D9217_, new_D9218_, new_D9219_,
    new_D9220_, new_D9221_, new_D9222_, new_D9223_, new_D9224_, new_D9225_,
    new_D9226_, new_D9227_, new_D9228_, new_D9229_, new_D9230_, new_D9231_,
    new_D9232_, new_D9233_, new_D9234_, new_D9235_, new_D9236_, new_D9237_,
    new_D9238_, new_D9239_, new_D9240_, new_D9241_, new_D9242_, new_D9243_,
    new_D9244_, new_D9245_, new_D9246_, new_D9247_, new_D9248_, new_D9249_,
    new_D9250_, new_D9251_, new_D9252_, new_D9253_, new_D9254_, new_D9255_,
    new_D9256_, new_D9257_, new_D9258_, new_D9259_, new_D9260_, new_D9261_,
    new_D9262_, new_D9263_, new_D9264_, new_D9265_, new_D9266_, new_D9267_,
    new_D9268_, new_D9269_, new_D9270_, new_D9271_, new_D9272_, new_D9273_,
    new_D9274_, new_D9275_, new_D9276_, new_D9277_, new_D9278_, new_D9279_,
    new_D9280_, new_D9281_, new_D9282_, new_D9283_, new_D9284_, new_D9285_,
    new_D9286_, new_D9287_, new_D9288_, new_D9289_, new_D9290_, new_D9291_,
    new_D9292_, new_D9293_, new_D9294_, new_D9295_, new_D9296_, new_D9297_,
    new_D9298_, new_D9299_, new_D9300_, new_D9301_, new_D9302_, new_D9303_,
    new_D9304_, new_D9305_, new_D9306_, new_D9307_, new_D9308_, new_D9309_,
    new_D9310_, new_D9311_, new_D9312_, new_D9313_, new_D9314_, new_D9315_,
    new_D9316_, new_D9317_, new_D9318_, new_D9319_, new_D9320_, new_D9321_,
    new_D9322_, new_D9323_, new_D9324_, new_D9325_, new_D9326_, new_D9327_,
    new_D9328_, new_D9329_, new_D9330_, new_D9331_, new_D9332_, new_D9333_,
    new_D9334_, new_D9335_, new_D9336_, new_D9337_, new_D9338_, new_D9339_,
    new_D9340_, new_D9341_, new_D9342_, new_D9343_, new_D9344_, new_D9345_,
    new_D9346_, new_D9347_, new_D9348_, new_D9349_, new_D9350_, new_D9351_,
    new_D9352_, new_D9353_, new_D9354_, new_D9355_, new_D9356_, new_D9357_,
    new_D9358_, new_D9359_, new_D9360_, new_D9361_, new_D9362_, new_D9363_,
    new_D9364_, new_D9365_, new_D9366_, new_D9367_, new_D9368_, new_D9369_,
    new_D9370_, new_D9371_, new_D9372_, new_D9373_, new_D9374_, new_D9375_,
    new_D9376_, new_D9377_, new_D9378_, new_D9379_, new_D9380_, new_D9381_,
    new_D9382_, new_D9383_, new_D9384_, new_D9385_, new_D9386_, new_D9387_,
    new_D9388_, new_D9389_, new_D9390_, new_D9391_, new_D9392_, new_D9393_,
    new_D9394_, new_D9395_, new_D9396_, new_D9397_, new_D9398_, new_D9399_,
    new_D9400_, new_D9401_, new_D9402_, new_D9403_, new_D9404_, new_D9405_,
    new_D9406_, new_D9407_, new_D9408_, new_D9409_, new_D9410_, new_D9411_,
    new_D9412_, new_D9413_, new_D9414_, new_D9415_, new_D9416_, new_D9417_,
    new_D9418_, new_D9419_, new_D9420_, new_D9421_, new_D9422_, new_D9423_,
    new_D9424_, new_D9425_, new_D9426_, new_D9427_, new_D9428_, new_D9429_,
    new_D9430_, new_D9431_, new_D9432_, new_D9433_, new_D9434_, new_D9435_,
    new_D9436_, new_D9437_, new_D9438_, new_D9439_, new_D9440_, new_D9441_,
    new_D9442_, new_D9443_, new_D9444_, new_D9445_, new_D9446_, new_D9447_,
    new_D9448_, new_D9449_, new_D9450_, new_D9451_, new_D9452_, new_D9453_,
    new_D9454_, new_D9455_, new_D9456_, new_D9457_, new_D9458_, new_D9459_,
    new_D9460_, new_D9461_, new_D9462_, new_D9463_, new_D9464_, new_D9465_,
    new_D9466_, new_D9467_, new_D9468_, new_D9469_, new_D9470_, new_D9471_,
    new_D9472_, new_D9473_, new_D9474_, new_D9475_, new_D9476_, new_D9477_,
    new_D9478_, new_D9479_, new_D9480_, new_D9481_, new_D9482_, new_D9483_,
    new_D9484_, new_D9485_, new_D9486_, new_D9487_, new_D9488_, new_D9489_,
    new_D9490_, new_D9491_, new_D9492_, new_D9493_, new_D9494_, new_D9495_,
    new_D9496_, new_D9497_, new_D9498_, new_D9499_, new_D9500_, new_D9501_,
    new_D9502_, new_D9503_, new_D9504_, new_D9505_, new_D9506_, new_D9507_,
    new_D9508_, new_D9509_, new_D9510_, new_D9511_, new_D9512_, new_D9513_,
    new_D9514_, new_D9515_, new_D9516_, new_D9517_, new_D9518_, new_D9519_,
    new_D9520_, new_D9521_, new_D9522_, new_D9523_, new_D9524_, new_D9525_,
    new_D9526_, new_D9527_, new_D9528_, new_D9529_, new_D9530_, new_D9531_,
    new_D9532_, new_D9533_, new_D9534_, new_D9535_, new_D9536_, new_D9537_,
    new_D9538_, new_D9539_, new_D9540_, new_D9541_, new_D9542_, new_D9543_,
    new_D9544_, new_D9545_, new_D9546_, new_D9547_, new_D9548_, new_D9549_,
    new_D9550_, new_D9551_, new_D9552_, new_D9553_, new_D9554_, new_D9555_,
    new_D9556_, new_D9557_, new_D9558_, new_D9559_, new_D9560_, new_D9561_,
    new_D9562_, new_D9563_, new_D9564_, new_D9565_, new_D9566_, new_D9567_,
    new_D9568_, new_D9569_, new_D9570_, new_D9571_, new_D9572_, new_D9573_,
    new_D9574_, new_D9575_, new_D9576_, new_D9577_, new_D9578_, new_D9579_,
    new_D9580_, new_D9581_, new_D9582_, new_D9583_, new_D9584_, new_D9585_,
    new_D9586_, new_D9587_, new_D9588_, new_D9589_, new_D9590_, new_D9591_,
    new_D9592_, new_D9593_, new_D9594_, new_D9595_, new_D9596_, new_D9597_,
    new_D9598_, new_D9599_, new_D9600_, new_D9601_, new_D9602_, new_D9603_,
    new_D9604_, new_D9605_, new_D9606_, new_D9607_, new_D9608_, new_D9609_,
    new_D9610_, new_D9611_, new_D9612_, new_D9613_, new_D9614_, new_D9615_,
    new_D9616_, new_D9617_, new_D9618_, new_D9619_, new_D9620_, new_D9621_,
    new_D9622_, new_D9623_, new_D9624_, new_D9625_, new_D9626_, new_D9627_,
    new_D9628_, new_D9629_, new_D9630_, new_D9631_, new_D9632_, new_D9633_,
    new_D9634_, new_D9635_, new_D9636_, new_D9637_, new_D9638_, new_D9639_,
    new_D9640_, new_D9641_, new_D9642_, new_D9643_, new_D9644_, new_D9645_,
    new_D9646_, new_D9647_, new_D9648_, new_D9649_, new_D9650_, new_D9651_,
    new_D9652_, new_D9653_, new_D9654_, new_D9655_, new_D9656_, new_D9657_,
    new_D9658_, new_D9659_, new_D9660_, new_D9661_, new_D9662_, new_D9663_,
    new_D9664_, new_D9665_, new_D9666_, new_D9667_, new_D9668_, new_D9669_,
    new_D9670_, new_D9671_, new_D9672_, new_D9673_, new_D9674_, new_D9675_,
    new_D9676_, new_D9677_, new_D9678_, new_D9679_, new_D9680_, new_D9681_,
    new_D9682_, new_D9683_, new_D9684_, new_D9685_, new_D9686_, new_D9687_,
    new_D9688_, new_D9689_, new_D9690_, new_D9691_, new_D9692_, new_D9693_,
    new_D9694_, new_D9695_, new_D9696_, new_D9697_, new_D9698_, new_D9699_,
    new_D9700_, new_D9701_, new_D9702_, new_D9703_, new_D9704_, new_D9705_,
    new_D9706_, new_D9707_, new_D9708_, new_D9709_, new_D9710_, new_D9711_,
    new_D9712_, new_D9713_, new_D9714_, new_D9715_, new_D9716_, new_D9717_,
    new_D9718_, new_D9719_, new_D9720_, new_D9721_, new_D9722_, new_D9723_,
    new_D9724_, new_D9725_, new_D9726_, new_D9727_, new_D9728_, new_D9729_,
    new_D9730_, new_D9731_, new_D9732_, new_D9733_, new_D9734_, new_D9735_,
    new_D9736_, new_D9737_, new_D9738_, new_D9739_, new_D9740_, new_D9741_,
    new_D9742_, new_D9743_, new_D9744_, new_D9745_, new_D9746_, new_D9747_,
    new_D9748_, new_D9749_, new_D9750_, new_D9751_, new_D9752_, new_D9753_,
    new_D9754_, new_D9755_, new_D9756_, new_D9757_, new_D9758_, new_D9759_,
    new_D9760_, new_D9761_, new_D9762_, new_D9763_, new_D9764_, new_D9765_,
    new_D9766_, new_D9767_, new_D9768_, new_D9769_, new_D9770_, new_D9771_,
    new_D9772_, new_D9773_, new_D9774_, new_D9775_, new_D9776_, new_D9777_,
    new_D9778_, new_D9779_, new_D9780_, new_D9781_, new_D9782_, new_D9783_,
    new_D9784_, new_D9785_, new_D9786_, new_D9787_, new_D9788_, new_D9789_,
    new_D9790_, new_D9791_, new_D9792_, new_D9793_, new_D9794_, new_D9795_,
    new_D9796_, new_D9797_, new_D9798_, new_D9799_, new_D9800_, new_D9801_,
    new_D9802_, new_D9803_, new_D9804_, new_D9805_, new_D9806_, new_D9807_,
    new_D9808_, new_D9809_, new_D9810_, new_D9811_, new_D9812_, new_D9813_,
    new_D9814_, new_D9815_, new_D9816_, new_D9817_, new_D9818_, new_D9819_,
    new_D9820_, new_D9821_, new_D9822_, new_D9823_, new_D9824_, new_D9825_,
    new_D9826_, new_D9827_, new_D9828_, new_D9829_, new_D9830_, new_D9831_,
    new_D9832_, new_D9833_, new_D9834_, new_D9835_, new_D9836_, new_D9837_,
    new_D9838_, new_D9839_, new_D9840_, new_D9841_, new_D9842_, new_D9843_,
    new_D9844_, new_D9845_, new_D9846_, new_D9847_, new_D9848_, new_D9849_,
    new_D9850_, new_D9851_, new_D9852_, new_D9853_, new_D9854_, new_D9855_,
    new_D9856_, new_D9857_, new_D9858_, new_D9859_, new_D9860_, new_D9861_,
    new_D9862_, new_D9863_, new_D9864_, new_D9865_, new_D9866_, new_D9867_,
    new_D9868_, new_D9869_, new_D9870_, new_D9871_, new_D9872_, new_D9873_,
    new_D9874_, new_D9875_, new_D9876_, new_D9877_, new_D9878_, new_D9879_,
    new_D9880_, new_D9881_, new_D9882_, new_D9883_, new_D9884_, new_D9885_,
    new_D9886_, new_D9887_, new_D9888_, new_D9889_, new_D9890_, new_D9891_,
    new_D9892_, new_D9893_, new_D9894_, new_D9895_, new_D9896_, new_D9897_,
    new_D9898_, new_D9899_, new_D9900_, new_D9901_, new_D9902_, new_D9903_,
    new_D9904_, new_D9905_, new_D9906_, new_D9907_, new_D9908_, new_D9909_,
    new_D9910_, new_D9911_, new_D9912_, new_D9913_, new_D9914_, new_D9915_,
    new_D9916_, new_D9917_, new_D9918_, new_D9919_, new_D9920_, new_D9921_,
    new_D9922_, new_D9923_, new_D9924_, new_D9925_, new_D9926_, new_D9927_,
    new_D9928_, new_D9929_, new_D9930_, new_D9931_, new_D9932_, new_D9933_,
    new_D9934_, new_D9935_, new_D9936_, new_D9937_, new_D9938_, new_D9939_,
    new_D9940_, new_D9941_, new_D9942_, new_D9943_, new_D9944_, new_D9945_,
    new_D9946_, new_D9947_, new_D9948_, new_D9949_, new_D9950_, new_D9951_,
    new_D9952_, new_D9953_, new_D9954_, new_D9955_, new_D9956_, new_D9957_,
    new_D9958_, new_D9959_, new_D9960_, new_D9961_, new_D9962_, new_D9963_,
    new_D9964_, new_D9965_, new_D9966_, new_D9967_, new_D9968_, new_D9969_,
    new_D9970_, new_D9971_, new_D9972_, new_D9973_, new_D9974_, new_D9975_,
    new_D9976_, new_D9977_, new_D9978_, new_D9979_, new_D9980_, new_D9981_,
    new_D9982_, new_D9983_, new_D9984_, new_D9985_, new_D9986_, new_D9987_,
    new_D9988_, new_D9989_, new_D9990_, new_D9991_, new_D9992_, new_D9993_,
    new_D9994_, new_D9995_, new_D9996_, new_D9997_, new_D9998_, new_D9999_,
    new_E1_, new_E2_, new_E3_, new_E4_, new_E5_, new_E6_, new_E7_, new_E8_,
    new_E9_, new_E10_, new_E11_, new_E12_, new_E13_, new_E14_, new_E15_,
    new_E16_, new_E17_, new_E18_, new_E19_, new_E20_, new_E21_, new_E22_,
    new_E23_, new_E24_, new_E25_, new_E26_, new_E27_, new_E28_, new_E29_,
    new_E30_, new_E31_, new_E32_, new_E33_, new_E34_, new_E35_, new_E36_,
    new_E37_, new_E38_, new_E39_, new_E40_, new_E41_, new_E42_, new_E43_,
    new_E44_, new_E45_, new_E46_, new_E47_, new_E48_, new_E49_, new_E50_,
    new_E51_, new_E52_, new_E53_, new_E54_, new_E55_, new_E56_, new_E57_,
    new_E58_, new_E59_, new_E60_, new_E61_, new_E62_, new_E63_, new_E64_,
    new_E65_, new_E66_, new_E67_, new_E68_, new_E69_, new_E70_, new_E71_,
    new_E72_, new_E73_, new_E74_, new_E75_, new_E76_, new_E77_, new_E78_,
    new_E79_, new_E80_, new_E81_, new_E82_, new_E83_, new_E84_, new_E85_,
    new_E86_, new_E87_, new_E88_, new_E89_, new_E90_, new_E91_, new_E92_,
    new_E93_, new_E94_, new_E95_, new_E96_, new_E97_, new_E98_, new_E99_,
    new_E100_, new_E101_, new_E102_, new_E103_, new_E104_, new_E105_,
    new_E106_, new_E107_, new_E108_, new_E109_, new_E110_, new_E111_,
    new_E112_, new_E113_, new_E114_, new_E115_, new_E116_, new_E117_,
    new_E118_, new_E119_, new_E120_, new_E121_, new_E122_, new_E123_,
    new_E124_, new_E125_, new_E126_, new_E127_, new_E128_, new_E129_,
    new_E130_, new_E131_, new_E132_, new_E133_, new_E134_, new_E135_,
    new_E136_, new_E137_, new_E138_, new_E139_, new_E140_, new_E141_,
    new_E142_, new_E143_, new_E144_, new_E145_, new_E146_, new_E147_,
    new_E148_, new_E149_, new_E150_, new_E151_, new_E152_, new_E153_,
    new_E154_, new_E155_, new_E156_, new_E157_, new_E158_, new_E159_,
    new_E160_, new_E161_, new_E162_, new_E163_, new_E164_, new_E165_,
    new_E166_, new_E167_, new_E168_, new_E169_, new_E170_, new_E171_,
    new_E172_, new_E173_, new_E174_, new_E175_, new_E176_, new_E177_,
    new_E178_, new_E179_, new_E180_, new_E181_, new_E182_, new_E183_,
    new_E184_, new_E185_, new_E186_, new_E187_, new_E188_, new_E189_,
    new_E190_, new_E191_, new_E192_, new_E193_, new_E194_, new_E195_,
    new_E196_, new_E197_, new_E198_, new_E199_, new_E200_, new_E201_,
    new_E202_, new_E203_, new_E204_, new_E205_, new_E206_, new_E207_,
    new_E208_, new_E209_, new_E210_, new_E211_, new_E212_, new_E213_,
    new_E214_, new_E215_, new_E216_, new_E217_, new_E218_, new_E219_,
    new_E220_, new_E221_, new_E222_, new_E223_, new_E224_, new_E225_,
    new_E226_, new_E227_, new_E228_, new_E229_, new_E230_, new_E231_,
    new_E232_, new_E233_, new_E234_, new_E235_, new_E236_, new_E237_,
    new_E238_, new_E239_, new_E240_, new_E241_, new_E242_, new_E243_,
    new_E244_, new_E245_, new_E246_, new_E247_, new_E248_, new_E249_,
    new_E250_, new_E251_, new_E252_, new_E253_, new_E254_, new_E255_,
    new_E256_, new_E257_, new_E258_, new_E259_, new_E260_, new_E261_,
    new_E262_, new_E263_, new_E264_, new_E265_, new_E266_, new_E267_,
    new_E268_, new_E269_, new_E270_, new_E271_, new_E272_, new_E273_,
    new_E274_, new_E275_, new_E276_, new_E277_, new_E278_, new_E279_,
    new_E280_, new_E281_, new_E282_, new_E283_, new_E284_, new_E285_,
    new_E286_, new_E287_, new_E288_, new_E289_, new_E290_, new_E291_,
    new_E292_, new_E293_, new_E294_, new_E295_, new_E296_, new_E297_,
    new_E298_, new_E299_, new_E300_, new_E301_, new_E302_, new_E303_,
    new_E304_, new_E305_, new_E306_, new_E307_, new_E308_, new_E309_,
    new_E310_, new_E311_, new_E312_, new_E313_, new_E314_, new_E315_,
    new_E316_, new_E317_, new_E318_, new_E319_, new_E320_, new_E321_,
    new_E322_, new_E323_, new_E324_, new_E325_, new_E326_, new_E327_,
    new_E328_, new_E329_, new_E330_, new_E331_, new_E332_, new_E333_,
    new_E334_, new_E335_, new_E336_, new_E337_, new_E338_, new_E339_,
    new_E340_, new_E341_, new_E342_, new_E343_, new_E344_, new_E345_,
    new_E346_, new_E347_, new_E348_, new_E349_, new_E350_, new_E351_,
    new_E352_, new_E353_, new_E354_, new_E355_, new_E356_, new_E357_,
    new_E358_, new_E359_, new_E360_, new_E361_, new_E362_, new_E363_,
    new_E364_, new_E365_, new_E366_, new_E367_, new_E368_, new_E369_,
    new_E370_, new_E371_, new_E372_, new_E373_, new_E374_, new_E375_,
    new_E376_, new_E377_, new_E378_, new_E379_, new_E380_, new_E381_,
    new_E382_, new_E383_, new_E384_, new_E385_, new_E386_, new_E387_,
    new_E388_, new_E389_, new_E390_, new_E391_, new_E392_, new_E393_,
    new_E394_, new_E395_, new_E396_, new_E397_, new_E398_, new_E399_,
    new_E400_, new_E401_, new_E402_, new_E403_, new_E404_, new_E405_,
    new_E406_, new_E407_, new_E408_, new_E409_, new_E410_, new_E411_,
    new_E412_, new_E413_, new_E414_, new_E415_, new_E416_, new_E417_,
    new_E418_, new_E419_, new_E420_, new_E421_, new_E422_, new_E423_,
    new_E424_, new_E425_, new_E426_, new_E427_, new_E428_, new_E429_,
    new_E430_, new_E431_, new_E432_, new_E433_, new_E434_, new_E435_,
    new_E436_, new_E437_, new_E438_, new_E439_, new_E440_, new_E441_,
    new_E442_, new_E443_, new_E444_, new_E445_, new_E446_, new_E447_,
    new_E448_, new_E449_, new_E450_, new_E451_, new_E452_, new_E453_,
    new_E454_, new_E455_, new_E456_, new_E457_, new_E458_, new_E459_,
    new_E460_, new_E461_, new_E462_, new_E463_, new_E464_, new_E465_,
    new_E466_, new_E467_, new_E468_, new_E469_, new_E470_, new_E471_,
    new_E472_, new_E473_, new_E474_, new_E475_, new_E476_, new_E477_,
    new_E478_, new_E479_, new_E480_, new_E481_, new_E482_, new_E483_,
    new_E484_, new_E485_, new_E486_, new_E487_, new_E488_, new_E489_,
    new_E490_, new_E491_, new_E492_, new_E493_, new_E494_, new_E495_,
    new_E496_, new_E497_, new_E498_, new_E499_, new_E500_, new_E501_,
    new_E502_, new_E503_, new_E504_, new_E505_, new_E506_, new_E507_,
    new_E508_, new_E509_, new_E510_, new_E511_, new_E512_, new_E513_,
    new_E514_, new_E515_, new_E516_, new_E517_, new_E518_, new_E519_,
    new_E520_, new_E521_, new_E522_, new_E523_, new_E524_, new_E525_,
    new_E526_, new_E527_, new_E528_, new_E529_, new_E530_, new_E531_,
    new_E532_, new_E533_, new_E534_, new_E535_, new_E536_, new_E537_,
    new_E538_, new_E539_, new_E540_, new_E541_, new_E542_, new_E543_,
    new_E544_, new_E545_, new_E546_, new_E547_, new_E548_, new_E549_,
    new_E550_, new_E551_, new_E552_, new_E553_, new_E554_, new_E555_,
    new_E556_, new_E557_, new_E558_, new_E559_, new_E560_, new_E561_,
    new_E562_, new_E563_, new_E564_, new_E565_, new_E566_, new_E567_,
    new_E568_, new_E569_, new_E570_, new_E571_, new_E572_, new_E573_,
    new_E574_, new_E575_, new_E576_, new_E577_, new_E578_, new_E579_,
    new_E580_, new_E581_, new_E582_, new_E583_, new_E584_, new_E585_,
    new_E586_, new_E587_, new_E588_, new_E589_, new_E590_, new_E591_,
    new_E592_, new_E593_, new_E594_, new_E595_, new_E596_, new_E597_,
    new_E598_, new_E599_, new_E600_, new_E601_, new_E602_, new_E603_,
    new_E604_, new_E605_, new_E606_, new_E607_, new_E608_, new_E609_,
    new_E610_, new_E611_, new_E612_, new_E613_, new_E614_, new_E615_,
    new_E616_, new_E617_, new_E618_, new_E619_, new_E620_, new_E621_,
    new_E622_, new_E623_, new_E624_, new_E625_, new_E626_, new_E627_,
    new_E628_, new_E629_, new_E630_, new_E631_, new_E632_, new_E633_,
    new_E634_, new_E635_, new_E636_, new_E637_, new_E638_, new_E639_,
    new_E640_, new_E641_, new_E642_, new_E643_, new_E644_, new_E645_,
    new_E646_, new_E647_, new_E648_, new_E649_, new_E650_, new_E651_,
    new_E652_, new_E653_, new_E654_, new_E655_, new_E656_, new_E657_,
    new_E658_, new_E659_, new_E660_, new_E661_, new_E662_, new_E663_,
    new_E664_, new_E665_, new_E666_, new_E667_, new_E668_, new_E669_,
    new_E670_, new_E671_, new_E672_, new_E673_, new_E674_, new_E675_,
    new_E676_, new_E677_, new_E678_, new_E679_, new_E680_, new_E681_,
    new_E682_, new_E683_, new_E684_, new_E685_, new_E686_, new_E687_,
    new_E688_, new_E689_, new_E690_, new_E691_, new_E692_, new_E693_,
    new_E694_, new_E695_, new_E696_, new_E697_, new_E698_, new_E699_,
    new_E700_, new_E701_, new_E702_, new_E703_, new_E704_, new_E705_,
    new_E706_, new_E707_, new_E708_, new_E709_, new_E710_, new_E711_,
    new_E712_, new_E713_, new_E714_, new_E715_, new_E716_, new_E717_,
    new_E718_, new_E719_, new_E720_, new_E721_, new_E722_, new_E723_,
    new_E724_, new_E725_, new_E726_, new_E727_, new_E728_, new_E729_,
    new_E730_, new_E731_, new_E732_, new_E733_, new_E734_, new_E735_,
    new_E736_, new_E737_, new_E738_, new_E739_, new_E740_, new_E741_,
    new_E742_, new_E743_, new_E744_, new_E745_, new_E746_, new_E747_,
    new_E748_, new_E749_, new_E750_, new_E751_, new_E752_, new_E753_,
    new_E754_, new_E755_, new_E756_, new_E757_, new_E758_, new_E759_,
    new_E760_, new_E761_, new_E762_, new_E763_, new_E764_, new_E765_,
    new_E766_, new_E767_, new_E768_, new_E769_, new_E770_, new_E771_,
    new_E772_, new_E773_, new_E774_, new_E775_, new_E776_, new_E777_,
    new_E778_, new_E779_, new_E780_, new_E781_, new_E782_, new_E783_,
    new_E784_, new_E785_, new_E786_, new_E787_, new_E788_, new_E789_,
    new_E790_, new_E791_, new_E792_, new_E793_, new_E794_, new_E795_,
    new_E796_, new_E797_, new_E798_, new_E799_, new_E800_, new_E801_,
    new_E802_, new_E803_, new_E804_, new_E805_, new_E806_, new_E807_,
    new_E808_, new_E809_, new_E810_, new_E811_, new_E812_, new_E813_,
    new_E814_, new_E815_, new_E816_, new_E817_, new_E818_, new_E819_,
    new_E820_, new_E821_, new_E822_, new_E823_, new_E824_, new_E825_,
    new_E826_, new_E827_, new_E828_, new_E829_, new_E830_, new_E831_,
    new_E832_, new_E833_, new_E834_, new_E835_, new_E836_, new_E837_,
    new_E838_, new_E839_, new_E840_, new_E841_, new_E842_, new_E843_,
    new_E844_, new_E845_, new_E846_, new_E847_, new_E848_, new_E849_,
    new_E850_, new_E851_, new_E852_, new_E853_, new_E854_, new_E855_,
    new_E856_, new_E857_, new_E858_, new_E859_, new_E860_, new_E861_,
    new_E862_, new_E863_, new_E864_, new_E865_, new_E866_, new_E867_,
    new_E868_, new_E869_, new_E870_, new_E871_, new_E872_, new_E873_,
    new_E874_, new_E875_, new_E876_, new_E877_, new_E878_, new_E879_,
    new_E880_, new_E881_, new_E882_, new_E883_, new_E884_, new_E885_,
    new_E886_, new_E887_, new_E888_, new_E889_, new_E890_, new_E891_,
    new_E892_, new_E893_, new_E894_, new_E895_, new_E896_, new_E897_,
    new_E898_, new_E899_, new_E900_, new_E901_, new_E902_, new_E903_,
    new_E904_, new_E905_, new_E906_, new_E907_, new_E908_, new_E909_,
    new_E910_, new_E911_, new_E912_, new_E913_, new_E914_, new_E915_,
    new_E916_, new_E917_, new_E918_, new_E919_, new_E920_, new_E921_,
    new_E922_, new_E923_, new_E924_, new_E925_, new_E926_, new_E927_,
    new_E928_, new_E929_, new_E930_, new_E931_, new_E932_, new_E933_,
    new_E934_, new_E935_, new_E936_, new_E937_, new_E938_, new_E939_,
    new_E940_, new_E941_, new_E942_, new_E943_, new_E944_, new_E945_,
    new_E946_, new_E947_, new_E948_, new_E949_, new_E950_, new_E951_,
    new_E952_, new_E953_, new_E954_, new_E955_, new_E956_, new_E957_,
    new_E958_, new_E959_, new_E960_, new_E961_, new_E962_, new_E963_,
    new_E964_, new_E965_, new_E966_, new_E967_, new_E968_, new_E969_,
    new_E970_, new_E971_, new_E972_, new_E973_, new_E974_, new_E975_,
    new_E976_, new_E977_, new_E978_, new_E979_, new_E980_, new_E981_,
    new_E982_, new_E983_, new_E984_, new_E985_, new_E986_, new_E987_,
    new_E988_, new_E989_, new_E990_, new_E991_, new_E992_, new_E993_,
    new_E994_, new_E995_, new_E996_, new_E997_, new_E998_, new_E999_,
    new_E1000_, new_E1001_, new_E1002_, new_E1003_, new_E1004_, new_E1005_,
    new_E1006_, new_E1007_, new_E1008_, new_E1009_, new_E1010_, new_E1011_,
    new_E1012_, new_E1013_, new_E1014_, new_E1015_, new_E1016_, new_E1017_,
    new_E1018_, new_E1019_, new_E1020_, new_E1021_, new_E1022_, new_E1023_,
    new_E1024_, new_E1025_, new_E1026_, new_E1027_, new_E1028_, new_E1029_,
    new_E1030_, new_E1031_, new_E1032_, new_E1033_, new_E1034_, new_E1035_,
    new_E1036_, new_E1037_, new_E1038_, new_E1039_, new_E1040_, new_E1041_,
    new_E1042_, new_E1043_, new_E1044_, new_E1045_, new_E1046_, new_E1047_,
    new_E1048_, new_E1049_, new_E1050_, new_E1051_, new_E1052_, new_E1053_,
    new_E1054_, new_E1055_, new_E1056_, new_E1057_, new_E1058_, new_E1059_,
    new_E1060_, new_E1061_, new_E1062_, new_E1063_, new_E1064_, new_E1065_,
    new_E1066_, new_E1067_, new_E1068_, new_E1069_, new_E1070_, new_E1071_,
    new_E1072_, new_E1073_, new_E1074_, new_E1075_, new_E1076_, new_E1077_,
    new_E1078_, new_E1079_, new_E1080_, new_E1081_, new_E1082_, new_E1083_,
    new_E1084_, new_E1085_, new_E1086_, new_E1087_, new_E1088_, new_E1089_,
    new_E1090_, new_E1091_, new_E1092_, new_E1093_, new_E1094_, new_E1095_,
    new_E1096_, new_E1097_, new_E1098_, new_E1099_, new_E1100_, new_E1101_,
    new_E1102_, new_E1103_, new_E1104_, new_E1105_, new_E1106_, new_E1107_,
    new_E1108_, new_E1109_, new_E1110_, new_E1111_, new_E1112_, new_E1113_,
    new_E1114_, new_E1115_, new_E1116_, new_E1117_, new_E1118_, new_E1119_,
    new_E1120_, new_E1121_, new_E1122_, new_E1123_, new_E1124_, new_E1125_,
    new_E1126_, new_E1127_, new_E1128_, new_E1129_, new_E1130_, new_E1131_,
    new_E1132_, new_E1133_, new_E1134_, new_E1135_, new_E1136_, new_E1137_,
    new_E1138_, new_E1139_, new_E1140_, new_E1141_, new_E1142_, new_E1143_,
    new_E1144_, new_E1145_, new_E1146_, new_E1147_, new_E1148_, new_E1149_,
    new_E1150_, new_E1151_, new_E1152_, new_E1153_, new_E1154_, new_E1155_,
    new_E1156_, new_E1157_, new_E1158_, new_E1159_, new_E1160_, new_E1161_,
    new_E1162_, new_E1163_, new_E1164_, new_E1165_, new_E1166_, new_E1167_,
    new_E1168_, new_E1169_, new_E1170_, new_E1171_, new_E1172_, new_E1173_,
    new_E1174_, new_E1175_, new_E1176_, new_E1177_, new_E1178_, new_E1179_,
    new_E1180_, new_E1181_, new_E1182_, new_E1183_, new_E1184_, new_E1185_,
    new_E1186_, new_E1187_, new_E1188_, new_E1189_, new_E1190_, new_E1191_,
    new_E1192_, new_E1193_, new_E1194_, new_E1195_, new_E1196_, new_E1197_,
    new_E1198_, new_E1199_, new_E1200_, new_E1201_, new_E1202_, new_E1203_,
    new_E1204_, new_E1205_, new_E1206_, new_E1207_, new_E1208_, new_E1209_,
    new_E1210_, new_E1211_, new_E1212_, new_E1213_, new_E1214_, new_E1215_,
    new_E1216_, new_E1217_, new_E1218_, new_E1219_, new_E1220_, new_E1221_,
    new_E1222_, new_E1223_, new_E1224_, new_E1225_, new_E1226_, new_E1227_,
    new_E1228_, new_E1229_, new_E1230_, new_E1231_, new_E1232_, new_E1233_,
    new_E1234_, new_E1235_, new_E1236_, new_E1237_, new_E1238_, new_E1239_,
    new_E1240_, new_E1241_, new_E1242_, new_E1243_, new_E1244_, new_E1245_,
    new_E1246_, new_E1247_, new_E1248_, new_E1249_, new_E1250_, new_E1251_,
    new_E1252_, new_E1253_, new_E1254_, new_E1255_, new_E1256_, new_E1257_,
    new_E1258_, new_E1259_, new_E1260_, new_E1261_, new_E1262_, new_E1263_,
    new_E1264_, new_E1265_, new_E1266_, new_E1267_, new_E1268_, new_E1269_,
    new_E1270_, new_E1271_, new_E1272_, new_E1273_, new_E1274_, new_E1275_,
    new_E1276_, new_E1277_, new_E1278_, new_E1279_, new_E1280_, new_E1281_,
    new_E1282_, new_E1283_, new_E1284_, new_E1285_, new_E1286_, new_E1287_,
    new_E1288_, new_E1289_, new_E1290_, new_E1291_, new_E1292_, new_E1293_,
    new_E1294_, new_E1295_, new_E1296_, new_E1297_, new_E1298_, new_E1299_,
    new_E1300_, new_E1301_, new_E1302_, new_E1303_, new_E1304_, new_E1305_,
    new_E1306_, new_E1307_, new_E1308_, new_E1309_, new_E1310_, new_E1311_,
    new_E1312_, new_E1313_, new_E1314_, new_E1315_, new_E1316_, new_E1317_,
    new_E1318_, new_E1319_, new_E1320_, new_E1321_, new_E1322_, new_E1323_,
    new_E1324_, new_E1325_, new_E1326_, new_E1327_, new_E1328_, new_E1329_,
    new_E1330_, new_E1331_, new_E1332_, new_E1333_, new_E1334_, new_E1335_,
    new_E1336_, new_E1337_, new_E1338_, new_E1339_, new_E1340_, new_E1341_,
    new_E1342_, new_E1343_, new_E1344_, new_E1345_, new_E1346_, new_E1347_,
    new_E1348_, new_E1349_, new_E1350_, new_E1351_, new_E1352_, new_E1353_,
    new_E1354_, new_E1355_, new_E1356_, new_E1357_, new_E1358_, new_E1359_,
    new_E1360_, new_E1361_, new_E1362_, new_E1363_, new_E1364_, new_E1365_,
    new_E1366_, new_E1367_, new_E1368_, new_E1369_, new_E1370_, new_E1371_,
    new_E1372_, new_E1373_, new_E1374_, new_E1375_, new_E1376_, new_E1377_,
    new_E1378_, new_E1379_, new_E1380_, new_E1381_, new_E1382_, new_E1383_,
    new_E1384_, new_E1385_, new_E1386_, new_E1387_, new_E1388_, new_E1389_,
    new_E1390_, new_E1391_, new_E1392_, new_E1393_, new_E1394_, new_E1395_,
    new_E1396_, new_E1397_, new_E1398_, new_E1399_, new_E1400_, new_E1401_,
    new_E1402_, new_E1403_, new_E1404_, new_E1405_, new_E1406_, new_E1407_,
    new_E1408_, new_E1409_, new_E1410_, new_E1411_, new_E1412_, new_E1413_,
    new_E1414_, new_E1415_, new_E1416_, new_E1417_, new_E1418_, new_E1419_,
    new_E1420_, new_E1421_, new_E1422_, new_E1423_, new_E1424_, new_E1425_,
    new_E1426_, new_E1427_, new_E1428_, new_E1429_, new_E1430_, new_E1431_,
    new_E1432_, new_E1433_, new_E1434_, new_E1435_, new_E1436_, new_E1437_,
    new_E1438_, new_E1439_, new_E1440_, new_E1441_, new_E1442_, new_E1443_,
    new_E1444_, new_E1445_, new_E1446_, new_E1447_, new_E1448_, new_E1449_,
    new_E1450_, new_E1451_, new_E1452_, new_E1453_, new_E1454_, new_E1455_,
    new_E1456_, new_E1457_, new_E1458_, new_E1459_, new_E1460_, new_E1461_,
    new_E1462_, new_E1463_, new_E1464_, new_E1465_, new_E1466_, new_E1467_,
    new_E1468_, new_E1469_, new_E1470_, new_E1471_, new_E1472_, new_E1473_,
    new_E1474_, new_E1475_, new_E1476_, new_E1477_, new_E1478_, new_E1479_,
    new_E1480_, new_E1481_, new_E1482_, new_E1483_, new_E1484_, new_E1485_,
    new_E1486_, new_E1487_, new_E1488_, new_E1489_, new_E1490_, new_E1491_,
    new_E1492_, new_E1493_, new_E1494_, new_E1495_, new_E1496_, new_E1497_,
    new_E1498_, new_E1499_, new_E1500_, new_E1501_, new_E1502_, new_E1503_,
    new_E1504_, new_E1505_, new_E1506_, new_E1507_, new_E1508_, new_E1509_,
    new_E1510_, new_E1511_, new_E1512_, new_E1513_, new_E1514_, new_E1515_,
    new_E1516_, new_E1517_, new_E1518_, new_E1519_, new_E1520_, new_E1521_,
    new_E1522_, new_E1523_, new_E1524_, new_E1525_, new_E1526_, new_E1527_,
    new_E1528_, new_E1529_, new_E1530_, new_E1531_, new_E1532_, new_E1533_,
    new_E1534_, new_E1535_, new_E1536_, new_E1537_, new_E1538_, new_E1539_,
    new_E1540_, new_E1541_, new_E1542_, new_E1543_, new_E1544_, new_E1545_,
    new_E1546_, new_E1547_, new_E1548_, new_E1549_, new_E1550_, new_E1551_,
    new_E1552_, new_E1553_, new_E1554_, new_E1555_, new_E1556_, new_E1557_,
    new_E1558_, new_E1559_, new_E1560_, new_E1561_, new_E1562_, new_E1563_,
    new_E1564_, new_E1565_, new_E1566_, new_E1567_, new_E1568_, new_E1569_,
    new_E1570_, new_E1571_, new_E1572_, new_E1573_, new_E1574_, new_E1575_,
    new_E1576_, new_E1577_, new_E1578_, new_E1579_, new_E1580_, new_E1581_,
    new_E1582_, new_E1583_, new_E1584_, new_E1585_, new_E1586_, new_E1587_,
    new_E1588_, new_E1589_, new_E1590_, new_E1591_, new_E1592_, new_E1593_,
    new_E1594_, new_E1595_, new_E1596_, new_E1597_, new_E1598_, new_E1599_,
    new_E1600_, new_E1601_, new_E1602_, new_E1603_, new_E1604_, new_E1605_,
    new_E1606_, new_E1607_, new_E1608_, new_E1609_, new_E1610_, new_E1611_,
    new_E1612_, new_E1613_, new_E1614_, new_E1615_, new_E1616_, new_E1617_,
    new_E1618_, new_E1619_, new_E1620_, new_E1621_, new_E1622_, new_E1623_,
    new_E1624_, new_E1625_, new_E1626_, new_E1627_, new_E1628_, new_E1629_,
    new_E1630_, new_E1631_, new_E1632_, new_E1633_, new_E1634_, new_E1635_,
    new_E1636_, new_E1637_, new_E1638_, new_E1639_, new_E1640_, new_E1641_,
    new_E1642_, new_E1643_, new_E1644_, new_E1645_, new_E1646_, new_E1647_,
    new_E1648_, new_E1649_, new_E1650_, new_E1651_, new_E1652_, new_E1653_,
    new_E1654_, new_E1655_, new_E1656_, new_E1657_, new_E1658_, new_E1659_,
    new_E1660_, new_E1661_, new_E1662_, new_E1663_, new_E1664_, new_E1665_,
    new_E1666_, new_E1667_, new_E1668_, new_E1669_, new_E1670_, new_E1671_,
    new_E1672_, new_E1673_, new_E1674_, new_E1675_, new_E1676_, new_E1677_,
    new_E1678_, new_E1679_, new_E1680_, new_E1681_, new_E1682_, new_E1683_,
    new_E1684_, new_E1685_, new_E1686_, new_E1687_, new_E1688_, new_E1689_,
    new_E1690_, new_E1691_, new_E1692_, new_E1693_, new_E1694_, new_E1695_,
    new_E1696_, new_E1697_, new_E1698_, new_E1699_, new_E1700_, new_E1701_,
    new_E1702_, new_E1703_, new_E1704_, new_E1705_, new_E1706_, new_E1707_,
    new_E1708_, new_E1709_, new_E1710_, new_E1711_, new_E1712_, new_E1713_,
    new_E1714_, new_E1715_, new_E1716_, new_E1717_, new_E1718_, new_E1719_,
    new_E1720_, new_E1721_, new_E1722_, new_E1723_, new_E1724_, new_E1725_,
    new_E1726_, new_E1727_, new_E1728_, new_E1729_, new_E1730_, new_E1731_,
    new_E1732_, new_E1733_, new_E1734_, new_E1735_, new_E1736_, new_E1737_,
    new_E1738_, new_E1739_, new_E1740_, new_E1741_, new_E1742_, new_E1743_,
    new_E1744_, new_E1745_, new_E1746_, new_E1747_, new_E1748_, new_E1749_,
    new_E1750_, new_E1751_, new_E1752_, new_E1753_, new_E1754_, new_E1755_,
    new_E1756_, new_E1757_, new_E1758_, new_E1759_, new_E1760_, new_E1761_,
    new_E1762_, new_E1763_, new_E1764_, new_E1765_, new_E1766_, new_E1767_,
    new_E1768_, new_E1769_, new_E1770_, new_E1771_, new_E1772_, new_E1773_,
    new_E1774_, new_E1775_, new_E1776_, new_E1777_, new_E1778_, new_E1779_,
    new_E1780_, new_E1781_, new_E1782_, new_E1783_, new_E1784_, new_E1785_,
    new_E1786_, new_E1787_, new_E1788_, new_E1789_, new_E1790_, new_E1791_,
    new_E1792_, new_E1793_, new_E1794_, new_E1795_, new_E1796_, new_E1797_,
    new_E1798_, new_E1799_, new_E1800_, new_E1801_, new_E1802_, new_E1803_,
    new_E1804_, new_E1805_, new_E1806_, new_E1807_, new_E1808_, new_E1809_,
    new_E1810_, new_E1811_, new_E1812_, new_E1813_, new_E1814_, new_E1815_,
    new_E1816_, new_E1817_, new_E1818_, new_E1819_, new_E1820_, new_E1821_,
    new_E1822_, new_E1823_, new_E1824_, new_E1825_, new_E1826_, new_E1827_,
    new_E1828_, new_E1829_, new_E1830_, new_E1831_, new_E1832_, new_E1833_,
    new_E1834_, new_E1835_, new_E1836_, new_E1837_, new_E1838_, new_E1839_,
    new_E1840_, new_E1841_, new_E1842_, new_E1843_, new_E1844_, new_E1845_,
    new_E1846_, new_E1847_, new_E1848_, new_E1849_, new_E1850_, new_E1851_,
    new_E1852_, new_E1853_, new_E1854_, new_E1855_, new_E1856_, new_E1857_,
    new_E1858_, new_E1859_, new_E1860_, new_E1861_, new_E1862_, new_E1863_,
    new_E1864_, new_E1865_, new_E1866_, new_E1867_, new_E1868_, new_E1869_,
    new_E1870_, new_E1871_, new_E1872_, new_E1873_, new_E1874_, new_E1875_,
    new_E1876_, new_E1877_, new_E1878_, new_E1879_, new_E1880_, new_E1881_,
    new_E1882_, new_E1883_, new_E1884_, new_E1885_, new_E1886_, new_E1887_,
    new_E1888_, new_E1889_, new_E1890_, new_E1891_, new_E1892_, new_E1893_,
    new_E1894_, new_E1895_, new_E1896_, new_E1897_, new_E1898_, new_E1899_,
    new_E1900_, new_E1901_, new_E1902_, new_E1903_, new_E1904_, new_E1905_,
    new_E1906_, new_E1907_, new_E1908_, new_E1909_, new_E1910_, new_E1911_,
    new_E1912_, new_E1913_, new_E1914_, new_E1915_, new_E1916_, new_E1917_,
    new_E1918_, new_E1919_, new_E1920_, new_E1921_, new_E1922_, new_E1923_,
    new_E1924_, new_E1925_, new_E1926_, new_E1927_, new_E1928_, new_E1929_,
    new_E1930_, new_E1931_, new_E1932_, new_E1933_, new_E1934_, new_E1935_,
    new_E1936_, new_E1937_, new_E1938_, new_E1939_, new_E1940_, new_E1941_,
    new_E1942_, new_E1943_, new_E1944_, new_E1945_, new_E1946_, new_E1947_,
    new_E1948_, new_E1949_, new_E1950_, new_E1951_, new_E1952_, new_E1953_,
    new_E1954_, new_E1955_, new_E1956_, new_E1957_, new_E1958_, new_E1959_,
    new_E1960_, new_E1961_, new_E1962_, new_E1963_, new_E1964_, new_E1965_,
    new_E1966_, new_E1967_, new_E1968_, new_E1969_, new_E1970_, new_E1971_,
    new_E1972_, new_E1973_, new_E1974_, new_E1975_, new_E1976_, new_E1977_,
    new_E1978_, new_E1979_, new_E1980_, new_E1981_, new_E1982_, new_E1983_,
    new_E1984_, new_E1985_, new_E1986_, new_E1987_, new_E1988_, new_E1989_,
    new_E1990_, new_E1991_, new_E1992_, new_E1993_, new_E1994_, new_E1995_,
    new_E1996_, new_E1997_, new_E1998_, new_E1999_, new_E2000_, new_E2001_,
    new_E2002_, new_E2003_, new_E2004_, new_E2005_, new_E2006_, new_E2007_,
    new_E2008_, new_E2009_, new_E2010_, new_E2011_, new_E2012_, new_E2013_,
    new_E2014_, new_E2015_, new_E2016_, new_E2017_, new_E2018_, new_E2019_,
    new_E2020_, new_E2021_, new_E2022_, new_E2023_, new_E2024_, new_E2025_,
    new_E2026_, new_E2027_, new_E2028_, new_E2029_, new_E2030_, new_E2031_,
    new_E2032_, new_E2033_, new_E2034_, new_E2035_, new_E2036_, new_E2037_,
    new_E2038_, new_E2039_, new_E2040_, new_E2041_, new_E2042_, new_E2043_,
    new_E2044_, new_E2045_, new_E2046_, new_E2047_, new_E2048_, new_E2049_,
    new_E2050_, new_E2051_, new_E2052_, new_E2053_, new_E2054_, new_E2055_,
    new_E2056_, new_E2057_, new_E2058_, new_E2059_, new_E2060_, new_E2061_,
    new_E2062_, new_E2063_, new_E2064_, new_E2065_, new_E2066_, new_E2067_,
    new_E2068_, new_E2069_, new_E2070_, new_E2071_, new_E2072_, new_E2073_,
    new_E2074_, new_E2075_, new_E2076_, new_E2077_, new_E2078_, new_E2079_,
    new_E2080_, new_E2081_, new_E2082_, new_E2083_, new_E2084_, new_E2085_,
    new_E2086_, new_E2087_, new_E2088_, new_E2089_, new_E2090_, new_E2091_,
    new_E2092_, new_E2093_, new_E2094_, new_E2095_, new_E2096_, new_E2097_,
    new_E2098_, new_E2099_, new_E2100_, new_E2101_, new_E2102_, new_E2103_,
    new_E2104_, new_E2105_, new_E2106_, new_E2107_, new_E2108_, new_E2109_,
    new_E2110_, new_E2111_, new_E2112_, new_E2113_, new_E2114_, new_E2115_,
    new_E2116_, new_E2117_, new_E2118_, new_E2119_, new_E2120_, new_E2121_,
    new_E2122_, new_E2123_, new_E2124_, new_E2125_, new_E2126_, new_E2127_,
    new_E2128_, new_E2129_, new_E2130_, new_E2131_, new_E2132_, new_E2133_,
    new_E2134_, new_E2135_, new_E2136_, new_E2137_, new_E2138_, new_E2139_,
    new_E2140_, new_E2141_, new_E2142_, new_E2143_, new_E2144_, new_E2145_,
    new_E2146_, new_E2147_, new_E2148_, new_E2149_, new_E2150_, new_E2151_,
    new_E2152_, new_E2153_, new_E2154_, new_E2155_, new_E2156_, new_E2157_,
    new_E2158_, new_E2159_, new_E2160_, new_E2161_, new_E2162_, new_E2163_,
    new_E2164_, new_E2165_, new_E2166_, new_E2167_, new_E2168_, new_E2169_,
    new_E2170_, new_E2171_, new_E2172_, new_E2173_, new_E2174_, new_E2175_,
    new_E2176_, new_E2177_, new_E2178_, new_E2179_, new_E2180_, new_E2181_,
    new_E2182_, new_E2183_, new_E2184_, new_E2185_, new_E2186_, new_E2187_,
    new_E2188_, new_E2189_, new_E2190_, new_E2191_, new_E2192_, new_E2193_,
    new_E2194_, new_E2195_, new_E2196_, new_E2197_, new_E2198_, new_E2199_,
    new_E2200_, new_E2201_, new_E2202_, new_E2203_, new_E2204_, new_E2205_,
    new_E2206_, new_E2207_, new_E2208_, new_E2209_, new_E2210_, new_E2211_,
    new_E2212_, new_E2213_, new_E2214_, new_E2215_, new_E2216_, new_E2217_,
    new_E2218_, new_E2219_, new_E2220_, new_E2221_, new_E2222_, new_E2223_,
    new_E2224_, new_E2225_, new_E2226_, new_E2227_, new_E2228_, new_E2229_,
    new_E2230_, new_E2231_, new_E2232_, new_E2233_, new_E2234_, new_E2235_,
    new_E2236_, new_E2237_, new_E2238_, new_E2239_, new_E2240_, new_E2241_,
    new_E2242_, new_E2243_, new_E2244_, new_E2245_, new_E2246_, new_E2247_,
    new_E2248_, new_E2249_, new_E2250_, new_E2251_, new_E2252_, new_E2253_,
    new_E2254_, new_E2255_, new_E2256_, new_E2257_, new_E2258_, new_E2259_,
    new_E2260_, new_E2261_, new_E2262_, new_E2263_, new_E2264_, new_E2265_,
    new_E2266_, new_E2267_, new_E2268_, new_E2269_, new_E2270_, new_E2271_,
    new_E2272_, new_E2273_, new_E2274_, new_E2275_, new_E2276_, new_E2277_,
    new_E2278_, new_E2279_, new_E2280_, new_E2281_, new_E2282_, new_E2283_,
    new_E2284_, new_E2285_, new_E2286_, new_E2287_, new_E2288_, new_E2289_,
    new_E2290_, new_E2291_, new_E2292_, new_E2293_, new_E2294_, new_E2295_,
    new_E2296_, new_E2297_, new_E2298_, new_E2299_, new_E2300_, new_E2301_,
    new_E2302_, new_E2303_, new_E2304_, new_E2305_, new_E2306_, new_E2307_,
    new_E2308_, new_E2309_, new_E2310_, new_E2311_, new_E2312_, new_E2313_,
    new_E2314_, new_E2315_, new_E2316_, new_E2317_, new_E2318_, new_E2319_,
    new_E2320_, new_E2321_, new_E2322_, new_E2323_, new_E2324_, new_E2325_,
    new_E2326_, new_E2327_, new_E2328_, new_E2329_, new_E2330_, new_E2331_,
    new_E2332_, new_E2333_, new_E2334_, new_E2335_, new_E2336_, new_E2337_,
    new_E2338_, new_E2339_, new_E2340_, new_E2341_, new_E2342_, new_E2343_,
    new_E2344_, new_E2345_, new_E2346_, new_E2347_, new_E2348_, new_E2349_,
    new_E2350_, new_E2351_, new_E2352_, new_E2353_, new_E2354_, new_E2355_,
    new_E2356_, new_E2357_, new_E2358_, new_E2359_, new_E2360_, new_E2361_,
    new_E2362_, new_E2363_, new_E2364_, new_E2365_, new_E2366_, new_E2367_,
    new_E2368_, new_E2369_, new_E2370_, new_E2371_, new_E2372_, new_E2373_,
    new_E2374_, new_E2375_, new_E2376_, new_E2377_, new_E2378_, new_E2379_,
    new_E2380_, new_E2381_, new_E2382_, new_E2383_, new_E2384_, new_E2385_,
    new_E2386_, new_E2387_, new_E2388_, new_E2389_, new_E2390_, new_E2391_,
    new_E2392_, new_E2393_, new_E2394_, new_E2395_, new_E2396_, new_E2397_,
    new_E2398_, new_E2399_, new_E2400_, new_E2401_, new_E2402_, new_E2403_,
    new_E2404_, new_E2405_, new_E2406_, new_E2407_, new_E2408_, new_E2409_,
    new_E2410_, new_E2411_, new_E2412_, new_E2413_, new_E2414_, new_E2415_,
    new_E2416_, new_E2417_, new_E2418_, new_E2419_, new_E2420_, new_E2421_,
    new_E2422_, new_E2423_, new_E2424_, new_E2425_, new_E2426_, new_E2427_,
    new_E2428_, new_E2429_, new_E2430_, new_E2431_, new_E2432_, new_E2433_,
    new_E2434_, new_E2435_, new_E2436_, new_E2437_, new_E2438_, new_E2439_,
    new_E2440_, new_E2441_, new_E2442_, new_E2443_, new_E2444_, new_E2445_,
    new_E2446_, new_E2447_, new_E2448_, new_E2449_, new_E2450_, new_E2451_,
    new_E2452_, new_E2453_, new_E2454_, new_E2455_, new_E2456_, new_E2457_,
    new_E2458_, new_E2459_, new_E2460_, new_E2461_, new_E2462_, new_E2463_,
    new_E2464_, new_E2465_, new_E2466_, new_E2467_, new_E2468_, new_E2469_,
    new_E2470_, new_E2471_, new_E2472_, new_E2473_, new_E2474_, new_E2475_,
    new_E2476_, new_E2477_, new_E2478_, new_E2479_, new_E2480_, new_E2481_,
    new_E2482_, new_E2483_, new_E2484_, new_E2485_, new_E2486_, new_E2487_,
    new_E2488_, new_E2489_, new_E2490_, new_E2491_, new_E2492_, new_E2493_,
    new_E2494_, new_E2495_, new_E2496_, new_E2497_, new_E2498_, new_E2499_,
    new_E2500_, new_E2501_, new_E2502_, new_E2503_, new_E2504_, new_E2505_,
    new_E2506_, new_E2507_, new_E2508_, new_E2509_, new_E2510_, new_E2511_,
    new_E2512_, new_E2513_, new_E2514_, new_E2515_, new_E2516_, new_E2517_,
    new_E2518_, new_E2519_, new_E2520_, new_E2521_, new_E2522_, new_E2523_,
    new_E2524_, new_E2525_, new_E2526_, new_E2527_, new_E2528_, new_E2529_,
    new_E2530_, new_E2531_, new_E2532_, new_E2533_, new_E2534_, new_E2535_,
    new_E2536_, new_E2537_, new_E2538_, new_E2539_, new_E2540_, new_E2541_,
    new_E2542_, new_E2543_, new_E2544_, new_E2545_, new_E2546_, new_E2547_,
    new_E2548_, new_E2549_, new_E2550_, new_E2551_, new_E2552_, new_E2553_,
    new_E2554_, new_E2555_, new_E2556_, new_E2557_, new_E2558_, new_E2559_,
    new_E2560_, new_E2561_, new_E2562_, new_E2563_, new_E2564_, new_E2565_,
    new_E2566_, new_E2567_, new_E2568_, new_E2569_, new_E2570_, new_E2571_,
    new_E2572_, new_E2573_, new_E2574_, new_E2575_, new_E2576_, new_E2577_,
    new_E2578_, new_E2579_, new_E2580_, new_E2581_, new_E2582_, new_E2583_,
    new_E2584_, new_E2585_, new_E2586_, new_E2587_, new_E2588_, new_E2589_,
    new_E2590_, new_E2591_, new_E2592_, new_E2593_, new_E2594_, new_E2595_,
    new_E2596_, new_E2597_, new_E2598_, new_E2599_, new_E2600_, new_E2601_,
    new_E2602_, new_E2603_, new_E2604_, new_E2605_, new_E2606_, new_E2607_,
    new_E2608_, new_E2609_, new_E2610_, new_E2611_, new_E2612_, new_E2613_,
    new_E2614_, new_E2615_, new_E2616_, new_E2617_, new_E2618_, new_E2619_,
    new_E2620_, new_E2621_, new_E2622_, new_E2623_, new_E2624_, new_E2625_,
    new_E2626_, new_E2627_, new_E2628_, new_E2629_, new_E2630_, new_E2631_,
    new_E2632_, new_E2633_, new_E2634_, new_E2635_, new_E2636_, new_E2637_,
    new_E2638_, new_E2639_, new_E2640_, new_E2641_, new_E2642_, new_E2643_,
    new_E2644_, new_E2645_, new_E2646_, new_E2647_, new_E2648_, new_E2649_,
    new_E2650_, new_E2651_, new_E2652_, new_E2653_, new_E2654_, new_E2655_,
    new_E2656_, new_E2657_, new_E2658_, new_E2659_, new_E2660_, new_E2661_,
    new_E2662_, new_E2663_, new_E2664_, new_E2665_, new_E2666_, new_E2667_,
    new_E2668_, new_E2669_, new_E2670_, new_E2671_, new_E2672_, new_E2673_,
    new_E2674_, new_E2675_, new_E2676_, new_E2677_, new_E2678_, new_E2679_,
    new_E2680_, new_E2681_, new_E2682_, new_E2683_, new_E2684_, new_E2685_,
    new_E2686_, new_E2687_, new_E2688_, new_E2689_, new_E2690_, new_E2691_,
    new_E2692_, new_E2693_, new_E2694_, new_E2695_, new_E2696_, new_E2697_,
    new_E2698_, new_E2699_, new_E2700_, new_E2701_, new_E2702_, new_E2703_,
    new_E2704_, new_E2705_, new_E2706_, new_E2707_, new_E2708_, new_E2709_,
    new_E2710_, new_E2711_, new_E2712_, new_E2713_, new_E2714_, new_E2715_,
    new_E2716_, new_E2717_, new_E2718_, new_E2719_, new_E2720_, new_E2721_,
    new_E2722_, new_E2723_, new_E2724_, new_E2725_, new_E2726_, new_E2727_,
    new_E2728_, new_E2729_, new_E2730_, new_E2731_, new_E2732_, new_E2733_,
    new_E2734_, new_E2735_, new_E2736_, new_E2737_, new_E2738_, new_E2739_,
    new_E2740_, new_E2741_, new_E2742_, new_E2743_, new_E2744_, new_E2745_,
    new_E2746_, new_E2747_, new_E2748_, new_E2749_, new_E2750_, new_E2751_,
    new_E2752_, new_E2753_, new_E2754_, new_E2755_, new_E2756_, new_E2757_,
    new_E2758_, new_E2759_, new_E2760_, new_E2761_, new_E2762_, new_E2763_,
    new_E2764_, new_E2765_, new_E2766_, new_E2767_, new_E2768_, new_E2769_,
    new_E2770_, new_E2771_, new_E2772_, new_E2773_, new_E2774_, new_E2775_,
    new_E2776_, new_E2777_, new_E2778_, new_E2779_, new_E2780_, new_E2781_,
    new_E2782_, new_E2783_, new_E2784_, new_E2785_, new_E2786_, new_E2787_,
    new_E2788_, new_E2789_, new_E2790_, new_E2791_, new_E2792_, new_E2793_,
    new_E2794_, new_E2795_, new_E2796_, new_E2797_, new_E2798_, new_E2799_,
    new_E2800_, new_E2801_, new_E2802_, new_E2803_, new_E2804_, new_E2805_,
    new_E2806_, new_E2807_, new_E2808_, new_E2809_, new_E2810_, new_E2811_,
    new_E2812_, new_E2813_, new_E2814_, new_E2815_, new_E2816_, new_E2817_,
    new_E2818_, new_E2819_, new_E2820_, new_E2821_, new_E2822_, new_E2823_,
    new_E2824_, new_E2825_, new_E2826_, new_E2827_, new_E2828_, new_E2829_,
    new_E2830_, new_E2831_, new_E2832_, new_E2833_, new_E2834_, new_E2835_,
    new_E2836_, new_E2837_, new_E2838_, new_E2839_, new_E2840_, new_E2841_,
    new_E2842_, new_E2843_, new_E2844_, new_E2845_, new_E2846_, new_E2847_,
    new_E2848_, new_E2849_, new_E2850_, new_E2851_, new_E2852_, new_E2853_,
    new_E2854_, new_E2855_, new_E2856_, new_E2857_, new_E2858_, new_E2859_,
    new_E2860_, new_E2861_, new_E2862_, new_E2863_, new_E2864_, new_E2865_,
    new_E2866_, new_E2867_, new_E2868_, new_E2869_, new_E2870_, new_E2871_,
    new_E2872_, new_E2873_, new_E2874_, new_E2875_, new_E2876_, new_E2877_,
    new_E2878_, new_E2879_, new_E2880_, new_E2881_, new_E2882_, new_E2883_,
    new_E2884_, new_E2885_, new_E2886_, new_E2887_, new_E2888_, new_E2889_,
    new_E2890_, new_E2891_, new_E2892_, new_E2893_, new_E2894_, new_E2895_,
    new_E2896_, new_E2897_, new_E2898_, new_E2899_, new_E2900_, new_E2901_,
    new_E2902_, new_E2903_, new_E2904_, new_E2905_, new_E2906_, new_E2907_,
    new_E2908_, new_E2909_, new_E2910_, new_E2911_, new_E2912_, new_E2913_,
    new_E2914_, new_E2915_, new_E2916_, new_E2917_, new_E2918_, new_E2919_,
    new_E2920_, new_E2921_, new_E2922_, new_E2923_, new_E2924_, new_E2925_,
    new_E2926_, new_E2927_, new_E2928_, new_E2929_, new_E2930_, new_E2931_,
    new_E2932_, new_E2933_, new_E2934_, new_E2935_, new_E2936_, new_E2937_,
    new_E2938_, new_E2939_, new_E2940_, new_E2941_, new_E2942_, new_E2943_,
    new_E2944_, new_E2945_, new_E2946_, new_E2947_, new_E2948_, new_E2949_,
    new_E2950_, new_E2951_, new_E2952_, new_E2953_, new_E2954_, new_E2955_,
    new_E2956_, new_E2957_, new_E2958_, new_E2959_, new_E2960_, new_E2961_,
    new_E2962_, new_E2963_, new_E2964_, new_E2965_, new_E2966_, new_E2967_,
    new_E2968_, new_E2969_, new_E2970_, new_E2971_, new_E2972_, new_E2973_,
    new_E2974_, new_E2975_, new_E2976_, new_E2977_, new_E2978_, new_E2979_,
    new_E2980_, new_E2981_, new_E2982_, new_E2983_, new_E2984_, new_E2985_,
    new_E2986_, new_E2987_, new_E2988_, new_E2989_, new_E2990_, new_E2991_,
    new_E2992_, new_E2993_, new_E2994_, new_E2995_, new_E2996_, new_E2997_,
    new_E2998_, new_E2999_, new_E3000_, new_E3001_, new_E3002_, new_E3003_,
    new_E3004_, new_E3005_, new_E3006_, new_E3007_, new_E3008_, new_E3009_,
    new_E3010_, new_E3011_, new_E3012_, new_E3013_, new_E3014_, new_E3015_,
    new_E3016_, new_E3017_, new_E3018_, new_E3019_, new_E3020_, new_E3021_,
    new_E3022_, new_E3023_, new_E3024_, new_E3025_, new_E3026_, new_E3027_,
    new_E3028_, new_E3029_, new_E3030_, new_E3031_, new_E3032_, new_E3033_,
    new_E3034_, new_E3035_, new_E3036_, new_E3037_, new_E3038_, new_E3039_,
    new_E3040_, new_E3041_, new_E3042_, new_E3043_, new_E3044_, new_E3045_,
    new_E3046_, new_E3047_, new_E3048_, new_E3049_, new_E3050_, new_E3051_,
    new_E3052_, new_E3053_, new_E3054_, new_E3055_, new_E3056_, new_E3057_,
    new_E3058_, new_E3059_, new_E3060_, new_E3061_, new_E3062_, new_E3063_,
    new_E3064_, new_E3065_, new_E3066_, new_E3067_, new_E3068_, new_E3069_,
    new_E3070_, new_E3071_, new_E3072_, new_E3073_, new_E3074_, new_E3075_,
    new_E3076_, new_E3077_, new_E3078_, new_E3079_, new_E3080_, new_E3081_,
    new_E3082_, new_E3083_, new_E3084_, new_E3085_, new_E3086_, new_E3087_,
    new_E3088_, new_E3089_, new_E3090_, new_E3091_, new_E3092_, new_E3093_,
    new_E3094_, new_E3095_, new_E3096_, new_E3097_, new_E3098_, new_E3099_,
    new_E3100_, new_E3101_, new_E3102_, new_E3103_, new_E3104_, new_E3105_,
    new_E3106_, new_E3107_, new_E3108_, new_E3109_, new_E3110_, new_E3111_,
    new_E3112_, new_E3113_, new_E3114_, new_E3115_, new_E3116_, new_E3117_,
    new_E3118_, new_E3119_, new_E3120_, new_E3121_, new_E3122_, new_E3123_,
    new_E3124_, new_E3125_, new_E3126_, new_E3127_, new_E3128_, new_E3129_,
    new_E3130_, new_E3131_, new_E3132_, new_E3133_, new_E3134_, new_E3135_,
    new_E3136_, new_E3137_, new_E3138_, new_E3139_, new_E3140_, new_E3141_,
    new_E3142_, new_E3143_, new_E3144_, new_E3145_, new_E3146_, new_E3147_,
    new_E3148_, new_E3149_, new_E3150_, new_E3151_, new_E3152_, new_E3153_,
    new_E3154_, new_E3155_, new_E3156_, new_E3157_, new_E3158_, new_E3159_,
    new_E3160_, new_E3161_, new_E3162_, new_E3163_, new_E3164_, new_E3165_,
    new_E3166_, new_E3167_, new_E3168_, new_E3169_, new_E3170_, new_E3171_,
    new_E3172_, new_E3173_, new_E3174_, new_E3175_, new_E3176_, new_E3177_,
    new_E3178_, new_E3179_, new_E3180_, new_E3181_, new_E3182_, new_E3183_,
    new_E3184_, new_E3185_, new_E3186_, new_E3187_, new_E3188_, new_E3189_,
    new_E3190_, new_E3191_, new_E3192_, new_E3193_, new_E3194_, new_E3195_,
    new_E3196_, new_E3197_, new_E3198_, new_E3199_, new_E3200_, new_E3201_,
    new_E3202_, new_E3203_, new_E3204_, new_E3205_, new_E3206_, new_E3207_,
    new_E3208_, new_E3209_, new_E3210_, new_E3211_, new_E3212_, new_E3213_,
    new_E3214_, new_E3215_, new_E3216_, new_E3217_, new_E3218_, new_E3219_,
    new_E3220_, new_E3221_, new_E3222_, new_E3223_, new_E3224_, new_E3225_,
    new_E3226_, new_E3227_, new_E3228_, new_E3229_, new_E3230_, new_E3231_,
    new_E3232_, new_E3233_, new_E3234_, new_E3235_, new_E3236_, new_E3237_,
    new_E3238_, new_E3239_, new_E3240_, new_E3241_, new_E3242_, new_E3243_,
    new_E3244_, new_E3245_, new_E3246_, new_E3247_, new_E3248_, new_E3249_,
    new_E3250_, new_E3251_, new_E3252_, new_E3253_, new_E3254_, new_E3255_,
    new_E3256_, new_E3257_, new_E3258_, new_E3259_, new_E3260_, new_E3261_,
    new_E3262_, new_E3263_, new_E3264_, new_E3265_, new_E3266_, new_E3267_,
    new_E3268_, new_E3269_, new_E3270_, new_E3271_, new_E3272_, new_E3273_,
    new_E3274_, new_E3275_, new_E3276_, new_E3277_, new_E3278_, new_E3279_,
    new_E3280_, new_E3281_, new_E3282_, new_E3283_, new_E3284_, new_E3285_,
    new_E3286_, new_E3287_, new_E3288_, new_E3289_, new_E3290_, new_E3291_,
    new_E3292_, new_E3293_, new_E3294_, new_E3295_, new_E3296_, new_E3297_,
    new_E3298_, new_E3299_, new_E3300_, new_E3301_, new_E3302_, new_E3303_,
    new_E3304_, new_E3305_, new_E3306_, new_E3307_, new_E3308_, new_E3309_,
    new_E3310_, new_E3311_, new_E3312_, new_E3313_, new_E3314_, new_E3315_,
    new_E3316_, new_E3317_, new_E3318_, new_E3319_, new_E3320_, new_E3321_,
    new_E3322_, new_E3323_, new_E3324_, new_E3325_, new_E3326_, new_E3327_,
    new_E3328_, new_E3329_, new_E3330_, new_E3331_, new_E3332_, new_E3333_,
    new_E3334_, new_E3335_, new_E3336_, new_E3337_, new_E3338_, new_E3339_,
    new_E3340_, new_E3341_, new_E3342_, new_E3343_, new_E3344_, new_E3345_,
    new_E3346_, new_E3347_, new_E3348_, new_E3349_, new_E3350_, new_E3351_,
    new_E3352_, new_E3353_, new_E3354_, new_E3355_, new_E3356_, new_E3357_,
    new_E3358_, new_E3359_, new_E3360_, new_E3361_, new_E3362_, new_E3363_,
    new_E3364_, new_E3365_, new_E3366_, new_E3367_, new_E3368_, new_E3369_,
    new_E3370_, new_E3371_, new_E3372_, new_E3373_, new_E3374_, new_E3375_,
    new_E3376_, new_E3377_, new_E3378_, new_E3379_, new_E3380_, new_E3381_,
    new_E3382_, new_E3383_, new_E3384_, new_E3385_, new_E3386_, new_E3387_,
    new_E3388_, new_E3389_, new_E3390_, new_E3391_, new_E3392_, new_E3393_,
    new_E3394_, new_E3395_, new_E3396_, new_E3397_, new_E3398_, new_E3399_,
    new_E3400_, new_E3401_, new_E3402_, new_E3403_, new_E3404_, new_E3405_,
    new_E3406_, new_E3407_, new_E3408_, new_E3409_, new_E3410_, new_E3411_,
    new_E3412_, new_E3413_, new_E3414_, new_E3415_, new_E3416_, new_E3417_,
    new_E3418_, new_E3419_, new_E3420_, new_E3421_, new_E3422_, new_E3423_,
    new_E3424_, new_E3425_, new_E3426_, new_E3427_, new_E3428_, new_E3429_,
    new_E3430_, new_E3431_, new_E3432_, new_E3433_, new_E3434_, new_E3435_,
    new_E3436_, new_E3437_, new_E3438_, new_E3439_, new_E3440_, new_E3441_,
    new_E3442_, new_E3443_, new_E3444_, new_E3445_, new_E3446_, new_E3447_,
    new_E3448_, new_E3449_, new_E3450_, new_E3451_, new_E3452_, new_E3453_,
    new_E3454_, new_E3455_, new_E3456_, new_E3457_, new_E3458_, new_E3459_,
    new_E3460_, new_E3461_, new_E3462_, new_E3463_, new_E3464_, new_E3465_,
    new_E3466_, new_E3467_, new_E3468_, new_E3469_, new_E3470_, new_E3471_,
    new_E3472_, new_E3473_, new_E3474_, new_E3475_, new_E3476_, new_E3477_,
    new_E3478_, new_E3479_, new_E3480_, new_E3481_, new_E3482_, new_E3483_,
    new_E3484_, new_E3485_, new_E3486_, new_E3487_, new_E3488_, new_E3489_,
    new_E3490_, new_E3491_, new_E3492_, new_E3493_, new_E3494_, new_E3495_,
    new_E3496_, new_E3497_, new_E3498_, new_E3499_, new_E3500_, new_E3501_,
    new_E3502_, new_E3503_, new_E3504_, new_E3505_, new_E3506_, new_E3507_,
    new_E3508_, new_E3509_, new_E3510_, new_E3511_, new_E3512_, new_E3513_,
    new_E3514_, new_E3515_, new_E3516_, new_E3517_, new_E3518_, new_E3519_,
    new_E3520_, new_E3521_, new_E3522_, new_E3523_, new_E3524_, new_E3525_,
    new_E3526_, new_E3527_, new_E3528_, new_E3529_, new_E3530_, new_E3531_,
    new_E3532_, new_E3533_, new_E3534_, new_E3535_, new_E3536_, new_E3537_,
    new_E3538_, new_E3539_, new_E3540_, new_E3541_, new_E3542_, new_E3543_,
    new_E3544_, new_E3545_, new_E3546_, new_E3547_, new_E3548_, new_E3549_,
    new_E3550_, new_E3551_, new_E3552_, new_E3553_, new_E3554_, new_E3555_,
    new_E3556_, new_E3557_, new_E3558_, new_E3559_, new_E3560_, new_E3561_,
    new_E3562_, new_E3563_, new_E3564_, new_E3565_, new_E3566_, new_E3567_,
    new_E3568_, new_E3569_, new_E3570_, new_E3571_, new_E3572_, new_E3573_,
    new_E3574_, new_E3575_, new_E3576_, new_E3577_, new_E3578_, new_E3579_,
    new_E3580_, new_E3581_, new_E3582_, new_E3583_, new_E3584_, new_E3585_,
    new_E3586_, new_E3587_, new_E3588_, new_E3589_, new_E3590_, new_E3591_,
    new_E3592_, new_E3593_, new_E3594_, new_E3595_, new_E3596_, new_E3597_,
    new_E3598_, new_E3599_, new_E3600_, new_E3601_, new_E3602_, new_E3603_,
    new_E3604_, new_E3605_, new_E3606_, new_E3607_, new_E3608_, new_E3609_,
    new_E3610_, new_E3611_, new_E3612_, new_E3613_, new_E3614_, new_E3615_,
    new_E3616_, new_E3617_, new_E3618_, new_E3619_, new_E3620_, new_E3621_,
    new_E3622_, new_E3623_, new_E3624_, new_E3625_, new_E3626_, new_E3627_,
    new_E3628_, new_E3629_, new_E3630_, new_E3631_, new_E3632_, new_E3633_,
    new_E3634_, new_E3635_, new_E3636_, new_E3637_, new_E3638_, new_E3639_,
    new_E3640_, new_E3641_, new_E3642_, new_E3643_, new_E3644_, new_E3645_,
    new_E3646_, new_E3647_, new_E3648_, new_E3649_, new_E3650_, new_E3651_,
    new_E3652_, new_E3653_, new_E3654_, new_E3655_, new_E3656_, new_E3657_,
    new_E3658_, new_E3659_, new_E3660_, new_E3661_, new_E3662_, new_E3663_,
    new_E3664_, new_E3665_, new_E3666_, new_E3667_, new_E3668_, new_E3669_,
    new_E3670_, new_E3671_, new_E3672_, new_E3673_, new_E3674_, new_E3675_,
    new_E3676_, new_E3677_, new_E3678_, new_E3679_, new_E3680_, new_E3681_,
    new_E3682_, new_E3683_, new_E3684_, new_E3685_, new_E3686_, new_E3687_,
    new_E3688_, new_E3689_, new_E3690_, new_E3691_, new_E3692_, new_E3693_,
    new_E3694_, new_E3695_, new_E3696_, new_E3697_, new_E3698_, new_E3699_,
    new_E3700_, new_E3701_, new_E3702_, new_E3703_, new_E3704_, new_E3705_,
    new_E3706_, new_E3707_, new_E3708_, new_E3709_, new_E3710_, new_E3711_,
    new_E3712_, new_E3713_, new_E3714_, new_E3715_, new_E3716_, new_E3717_,
    new_E3718_, new_E3719_, new_E3720_, new_E3721_, new_E3722_, new_E3723_,
    new_E3724_, new_E3725_, new_E3726_, new_E3727_, new_E3728_, new_E3729_,
    new_E3730_, new_E3731_, new_E3732_, new_E3733_, new_E3734_, new_E3735_,
    new_E3736_, new_E3737_, new_E3738_, new_E3739_, new_E3740_, new_E3741_,
    new_E3742_, new_E3743_, new_E3744_, new_E3745_, new_E3746_, new_E3747_,
    new_E3748_, new_E3749_, new_E3750_, new_E3751_, new_E3752_, new_E3753_,
    new_E3754_, new_E3755_, new_E3756_, new_E3757_, new_E3758_, new_E3759_,
    new_E3760_, new_E3761_, new_E3762_, new_E3763_, new_E3764_, new_E3765_,
    new_E3766_, new_E3767_, new_E3768_, new_E3769_, new_E3770_, new_E3771_,
    new_E3772_, new_E3773_, new_E3774_, new_E3775_, new_E3776_, new_E3777_,
    new_E3778_, new_E3779_, new_E3780_, new_E3781_, new_E3782_, new_E3783_,
    new_E3784_, new_E3785_, new_E3786_, new_E3787_, new_E3788_, new_E3789_,
    new_E3790_, new_E3791_, new_E3792_, new_E3793_, new_E3794_, new_E3795_,
    new_E3796_, new_E3797_, new_E3798_, new_E3799_, new_E3800_, new_E3801_,
    new_E3802_, new_E3803_, new_E3804_, new_E3805_, new_E3806_, new_E3807_,
    new_E3808_, new_E3809_, new_E3810_, new_E3811_, new_E3812_, new_E3813_,
    new_E3814_, new_E3815_, new_E3816_, new_E3817_, new_E3818_, new_E3819_,
    new_E3820_, new_E3821_, new_E3822_, new_E3823_, new_E3824_, new_E3825_,
    new_E3826_, new_E3827_, new_E3828_, new_E3829_, new_E3830_, new_E3831_,
    new_E3832_, new_E3833_, new_E3834_, new_E3835_, new_E3836_, new_E3837_,
    new_E3838_, new_E3839_, new_E3840_, new_E3841_, new_E3842_, new_E3843_,
    new_E3844_, new_E3845_, new_E3846_, new_E3847_, new_E3848_, new_E3849_,
    new_E3850_, new_E3851_, new_E3852_, new_E3853_, new_E3854_, new_E3855_,
    new_E3856_, new_E3857_, new_E3858_, new_E3859_, new_E3860_, new_E3861_,
    new_E3862_, new_E3863_, new_E3864_, new_E3865_, new_E3866_, new_E3867_,
    new_E3868_, new_E3869_, new_E3870_, new_E3871_, new_E3872_, new_E3873_,
    new_E3874_, new_E3875_, new_E3876_, new_E3877_, new_E3878_, new_E3879_,
    new_E3880_, new_E3881_, new_E3882_, new_E3883_, new_E3884_, new_E3885_,
    new_E3886_, new_E3887_, new_E3888_, new_E3889_, new_E3890_, new_E3891_,
    new_E3892_, new_E3893_, new_E3894_, new_E3895_, new_E3896_, new_E3897_,
    new_E3898_, new_E3899_, new_E3900_, new_E3901_, new_E3902_, new_E3903_,
    new_E3904_, new_E3905_, new_E3906_, new_E3907_, new_E3908_, new_E3909_,
    new_E3910_, new_E3911_, new_E3912_, new_E3913_, new_E3914_, new_E3915_,
    new_E3916_, new_E3917_, new_E3918_, new_E3919_, new_E3920_, new_E3921_,
    new_E3922_, new_E3923_, new_E3924_, new_E3925_, new_E3926_, new_E3927_,
    new_E3928_, new_E3929_, new_E3930_, new_E3931_, new_E3932_, new_E3933_,
    new_E3934_, new_E3935_, new_E3936_, new_E3937_, new_E3938_, new_E3939_,
    new_E3940_, new_E3941_, new_E3942_, new_E3943_, new_E3944_, new_E3945_,
    new_E3946_, new_E3947_, new_E3948_, new_E3949_, new_E3950_, new_E3951_,
    new_E3952_, new_E3953_, new_E3954_, new_E3955_, new_E3956_, new_E3957_,
    new_E3958_, new_E3959_, new_E3960_, new_E3961_, new_E3962_, new_E3963_,
    new_E3964_, new_E3965_, new_E3966_, new_E3967_, new_E3968_, new_E3969_,
    new_E3970_, new_E3971_, new_E3972_, new_E3973_, new_E3974_, new_E3975_,
    new_E3976_, new_E3977_, new_E3978_, new_E3979_, new_E3980_, new_E3981_,
    new_E3982_, new_E3983_, new_E3984_, new_E3985_, new_E3986_, new_E3987_,
    new_E3988_, new_E3989_, new_E3990_, new_E3991_, new_E3992_, new_E3993_,
    new_E3994_, new_E3995_, new_E3996_, new_E3997_, new_E3998_, new_E3999_,
    new_E4000_, new_E4001_, new_E4002_, new_E4003_, new_E4004_, new_E4005_,
    new_E4006_, new_E4007_, new_E4008_, new_E4009_, new_E4010_, new_E4011_,
    new_E4012_, new_E4013_, new_E4014_, new_E4015_, new_E4016_, new_E4017_,
    new_E4018_, new_E4019_, new_E4020_, new_E4021_, new_E4022_, new_E4023_,
    new_E4024_, new_E4025_, new_E4026_, new_E4027_, new_E4028_, new_E4029_,
    new_E4030_, new_E4031_, new_E4032_, new_E4033_, new_E4034_, new_E4035_,
    new_E4036_, new_E4037_, new_E4038_, new_E4039_, new_E4040_, new_E4041_,
    new_E4042_, new_E4043_, new_E4044_, new_E4045_, new_E4046_, new_E4047_,
    new_E4048_, new_E4049_, new_E4050_, new_E4051_, new_E4052_, new_E4053_,
    new_E4054_, new_E4055_, new_E4056_, new_E4057_, new_E4058_, new_E4059_,
    new_E4060_, new_E4061_, new_E4062_, new_E4063_, new_E4064_, new_E4065_,
    new_E4066_, new_E4067_, new_E4068_, new_E4069_, new_E4070_, new_E4071_,
    new_E4072_, new_E4073_, new_E4074_, new_E4075_, new_E4076_, new_E4077_,
    new_E4078_, new_E4079_, new_E4080_, new_E4081_, new_E4082_, new_E4083_,
    new_E4084_, new_E4085_, new_E4086_, new_E4087_, new_E4088_, new_E4089_,
    new_E4090_, new_E4091_, new_E4092_, new_E4093_, new_E4094_, new_E4095_,
    new_E4096_, new_E4097_, new_E4098_, new_E4099_, new_E4100_, new_E4101_,
    new_E4102_, new_E4103_, new_E4104_, new_E4105_, new_E4106_, new_E4107_,
    new_E4108_, new_E4109_, new_E4110_, new_E4111_, new_E4112_, new_E4113_,
    new_E4114_, new_E4115_, new_E4116_, new_E4117_, new_E4118_, new_E4119_,
    new_E4120_, new_E4121_, new_E4122_, new_E4123_, new_E4124_, new_E4125_,
    new_E4126_, new_E4127_, new_E4128_, new_E4129_, new_E4130_, new_E4131_,
    new_E4132_, new_E4133_, new_E4134_, new_E4135_, new_E4136_, new_E4137_,
    new_E4138_, new_E4139_, new_E4140_, new_E4141_, new_E4142_, new_E4143_,
    new_E4144_, new_E4145_, new_E4146_, new_E4147_, new_E4148_, new_E4149_,
    new_E4150_, new_E4151_, new_E4152_, new_E4153_, new_E4154_, new_E4155_,
    new_E4156_, new_E4157_, new_E4158_, new_E4159_, new_E4160_, new_E4161_,
    new_E4162_, new_E4163_, new_E4164_, new_E4165_, new_E4166_, new_E4167_,
    new_E4168_, new_E4169_, new_E4170_, new_E4171_, new_E4172_, new_E4173_,
    new_E4174_, new_E4175_, new_E4176_, new_E4177_, new_E4178_, new_E4179_,
    new_E4180_, new_E4181_, new_E4182_, new_E4183_, new_E4184_, new_E4185_,
    new_E4186_, new_E4187_, new_E4188_, new_E4189_, new_E4190_, new_E4191_,
    new_E4192_, new_E4193_, new_E4194_, new_E4195_, new_E4196_, new_E4197_,
    new_E4198_, new_E4199_, new_E4200_, new_E4201_, new_E4202_, new_E4203_,
    new_E4204_, new_E4205_, new_E4206_, new_E4207_, new_E4208_, new_E4209_,
    new_E4210_, new_E4211_, new_E4212_, new_E4213_, new_E4214_, new_E4215_,
    new_E4216_, new_E4217_, new_E4218_, new_E4219_, new_E4220_, new_E4221_,
    new_E4222_, new_E4223_, new_E4224_, new_E4225_, new_E4226_, new_E4227_,
    new_E4228_, new_E4229_, new_E4230_, new_E4231_, new_E4232_, new_E4233_,
    new_E4234_, new_E4235_, new_E4236_, new_E4237_, new_E4238_, new_E4239_,
    new_E4240_, new_E4241_, new_E4242_, new_E4243_, new_E4244_, new_E4245_,
    new_E4246_, new_E4247_, new_E4248_, new_E4249_, new_E4250_, new_E4251_,
    new_E4252_, new_E4253_, new_E4254_, new_E4255_, new_E4256_, new_E4257_,
    new_E4258_, new_E4259_, new_E4260_, new_E4261_, new_E4262_, new_E4263_,
    new_E4264_, new_E4265_, new_E4266_, new_E4267_, new_E4268_, new_E4269_,
    new_E4270_, new_E4271_, new_E4272_, new_E4273_, new_E4274_, new_E4275_,
    new_E4276_, new_E4277_, new_E4278_, new_E4279_, new_E4280_, new_E4281_,
    new_E4282_, new_E4283_, new_E4284_, new_E4285_, new_E4286_, new_E4287_,
    new_E4288_, new_E4289_, new_E4290_, new_E4291_, new_E4292_, new_E4293_,
    new_E4294_, new_E4295_, new_E4296_, new_E4297_, new_E4298_, new_E4299_,
    new_E4300_, new_E4301_, new_E4302_, new_E4303_, new_E4304_, new_E4305_,
    new_E4306_, new_E4307_, new_E4308_, new_E4309_, new_E4310_, new_E4311_,
    new_E4312_, new_E4313_, new_E4314_, new_E4315_, new_E4316_, new_E4317_,
    new_E4318_, new_E4319_, new_E4320_, new_E4321_, new_E4322_, new_E4323_,
    new_E4324_, new_E4325_, new_E4326_, new_E4327_, new_E4328_, new_E4329_,
    new_E4330_, new_E4331_, new_E4332_, new_E4333_, new_E4334_, new_E4335_,
    new_E4336_, new_E4337_, new_E4338_, new_E4339_, new_E4340_, new_E4341_,
    new_E4342_, new_E4343_, new_E4344_, new_E4345_, new_E4346_, new_E4347_,
    new_E4348_, new_E4349_, new_E4350_, new_E4351_, new_E4352_, new_E4353_,
    new_E4354_, new_E4355_, new_E4356_, new_E4357_, new_E4358_, new_E4359_,
    new_E4360_, new_E4361_, new_E4362_, new_E4363_, new_E4364_, new_E4365_,
    new_E4366_, new_E4367_, new_E4368_, new_E4369_, new_E4370_, new_E4371_,
    new_E4372_, new_E4373_, new_E4374_, new_E4375_, new_E4376_, new_E4377_,
    new_E4378_, new_E4379_, new_E4380_, new_E4381_, new_E4382_, new_E4383_,
    new_E4384_, new_E4385_, new_E4386_, new_E4387_, new_E4388_, new_E4389_,
    new_E4390_, new_E4391_, new_E4392_, new_E4393_, new_E4394_, new_E4395_,
    new_E4396_, new_E4397_, new_E4398_, new_E4399_, new_E4400_, new_E4401_,
    new_E4402_, new_E4403_, new_E4404_, new_E4405_, new_E4406_, new_E4407_,
    new_E4408_, new_E4409_, new_E4410_, new_E4411_, new_E4412_, new_E4413_,
    new_E4414_, new_E4415_, new_E4416_, new_E4417_, new_E4418_, new_E4419_,
    new_E4420_, new_E4421_, new_E4422_, new_E4423_, new_E4424_, new_E4425_,
    new_E4426_, new_E4427_, new_E4428_, new_E4429_, new_E4430_, new_E4431_,
    new_E4432_, new_E4433_, new_E4434_, new_E4435_, new_E4436_, new_E4437_,
    new_E4438_, new_E4439_, new_E4440_, new_E4441_, new_E4442_, new_E4443_,
    new_E4444_, new_E4445_, new_E4446_, new_E4447_, new_E4448_, new_E4449_,
    new_E4450_, new_E4451_, new_E4452_, new_E4453_, new_E4454_, new_E4455_,
    new_E4456_, new_E4457_, new_E4458_, new_E4459_, new_E4460_, new_E4461_,
    new_E4462_, new_E4463_, new_E4464_, new_E4465_, new_E4466_, new_E4467_,
    new_E4468_, new_E4469_, new_E4470_, new_E4471_, new_E4472_, new_E4473_,
    new_E4474_, new_E4475_, new_E4476_, new_E4477_, new_E4478_, new_E4479_,
    new_E4480_, new_E4481_, new_E4482_, new_E4483_, new_E4484_, new_E4485_,
    new_E4486_, new_E4487_, new_E4488_, new_E4489_, new_E4490_, new_E4491_,
    new_E4492_, new_E4493_, new_E4494_, new_E4495_, new_E4496_, new_E4497_,
    new_E4498_, new_E4499_, new_E4500_, new_E4501_, new_E4502_, new_E4503_,
    new_E4504_, new_E4505_, new_E4506_, new_E4507_, new_E4508_, new_E4509_,
    new_E4510_, new_E4511_, new_E4512_, new_E4513_, new_E4514_, new_E4515_,
    new_E4516_, new_E4517_, new_E4518_, new_E4519_, new_E4520_, new_E4521_,
    new_E4522_, new_E4523_, new_E4524_, new_E4525_, new_E4526_, new_E4527_,
    new_E4528_, new_E4529_, new_E4530_, new_E4531_, new_E4532_, new_E4533_,
    new_E4534_, new_E4535_, new_E4536_, new_E4537_, new_E4538_, new_E4539_,
    new_E4540_, new_E4541_, new_E4542_, new_E4543_, new_E4544_, new_E4545_,
    new_E4546_, new_E4547_, new_E4548_, new_E4549_, new_E4550_, new_E4551_,
    new_E4552_, new_E4553_, new_E4554_, new_E4555_, new_E4556_, new_E4557_,
    new_E4558_, new_E4559_, new_E4560_, new_E4561_, new_E4562_, new_E4563_,
    new_E4564_, new_E4565_, new_E4566_, new_E4567_, new_E4568_, new_E4569_,
    new_E4570_, new_E4571_, new_E4572_, new_E4573_, new_E4574_, new_E4575_,
    new_E4576_, new_E4577_, new_E4578_, new_E4579_, new_E4580_, new_E4581_,
    new_E4582_, new_E4583_, new_E4584_, new_E4585_, new_E4586_, new_E4587_,
    new_E4588_, new_E4589_, new_E4590_, new_E4591_, new_E4592_, new_E4593_,
    new_E4594_, new_E4595_, new_E4596_, new_E4597_, new_E4598_, new_E4599_,
    new_E4600_, new_E4601_, new_E4602_, new_E4603_, new_E4604_, new_E4605_,
    new_E4606_, new_E4607_, new_E4608_, new_E4609_, new_E4610_, new_E4611_,
    new_E4612_, new_E4613_, new_E4614_, new_E4615_, new_E4616_, new_E4617_,
    new_E4618_, new_E4619_, new_E4620_, new_E4621_, new_E4622_, new_E4623_,
    new_E4624_, new_E4625_, new_E4626_, new_E4627_, new_E4628_, new_E4629_,
    new_E4630_, new_E4631_, new_E4632_, new_E4633_, new_E4634_, new_E4635_,
    new_E4636_, new_E4637_, new_E4638_, new_E4639_, new_E4640_, new_E4641_,
    new_E4642_, new_E4643_, new_E4644_, new_E4645_, new_E4646_, new_E4647_,
    new_E4648_, new_E4649_, new_E4650_, new_E4651_, new_E4652_, new_E4653_,
    new_E4654_, new_E4655_, new_E4656_, new_E4657_, new_E4658_, new_E4659_,
    new_E4660_, new_E4661_, new_E4662_, new_E4663_, new_E4664_, new_E4665_,
    new_E4666_, new_E4667_, new_E4668_, new_E4669_, new_E4670_, new_E4671_,
    new_E4672_, new_E4673_, new_E4674_, new_E4675_, new_E4676_, new_E4677_,
    new_E4678_, new_E4679_, new_E4680_, new_E4681_, new_E4682_, new_E4683_,
    new_E4684_, new_E4685_, new_E4686_, new_E4687_, new_E4688_, new_E4689_,
    new_E4690_, new_E4691_, new_E4692_, new_E4693_, new_E4694_, new_E4695_,
    new_E4696_, new_E4697_, new_E4698_, new_E4699_, new_E4700_, new_E4701_,
    new_E4702_, new_E4703_, new_E4704_, new_E4705_, new_E4706_, new_E4707_,
    new_E4708_, new_E4709_, new_E4710_, new_E4711_, new_E4712_, new_E4713_,
    new_E4714_, new_E4715_, new_E4716_, new_E4717_, new_E4718_, new_E4719_,
    new_E4720_, new_E4721_, new_E4722_, new_E4723_, new_E4724_, new_E4725_,
    new_E4726_, new_E4727_, new_E4728_, new_E4729_, new_E4730_, new_E4731_,
    new_E4732_, new_E4733_, new_E4734_, new_E4735_, new_E4736_, new_E4737_,
    new_E4738_, new_E4739_, new_E4740_, new_E4741_, new_E4742_, new_E4743_,
    new_E4744_, new_E4745_, new_E4746_, new_E4747_, new_E4748_, new_E4749_,
    new_E4750_, new_E4751_, new_E4752_, new_E4753_, new_E4754_, new_E4755_,
    new_E4756_, new_E4757_, new_E4758_, new_E4759_, new_E4760_, new_E4761_,
    new_E4762_, new_E4763_, new_E4764_, new_E4765_, new_E4766_, new_E4767_,
    new_E4768_, new_E4769_, new_E4770_, new_E4771_, new_E4772_, new_E4773_,
    new_E4774_, new_E4775_, new_E4776_, new_E4777_, new_E4778_, new_E4779_,
    new_E4780_, new_E4781_, new_E4782_, new_E4783_, new_E4784_, new_E4785_,
    new_E4786_, new_E4787_, new_E4788_, new_E4789_, new_E4790_, new_E4791_,
    new_E4792_, new_E4793_, new_E4794_, new_E4795_, new_E4796_, new_E4797_,
    new_E4798_, new_E4799_, new_E4800_, new_E4801_, new_E4802_, new_E4803_,
    new_E4804_, new_E4805_, new_E4806_, new_E4807_, new_E4808_, new_E4809_,
    new_E4810_, new_E4811_, new_E4812_, new_E4813_, new_E4814_, new_E4815_,
    new_E4816_, new_E4817_, new_E4818_, new_E4819_, new_E4820_, new_E4821_,
    new_E4822_, new_E4823_, new_E4824_, new_E4825_, new_E4826_, new_E4827_,
    new_E4828_, new_E4829_, new_E4830_, new_E4831_, new_E4832_, new_E4833_,
    new_E4834_, new_E4835_, new_E4836_, new_E4837_, new_E4838_, new_E4839_,
    new_E4840_, new_E4841_, new_E4842_, new_E4843_, new_E4844_, new_E4845_,
    new_E4846_, new_E4847_, new_E4848_, new_E4849_, new_E4850_, new_E4851_,
    new_E4852_, new_E4853_, new_E4854_, new_E4855_, new_E4856_, new_E4857_,
    new_E4858_, new_E4859_, new_E4860_, new_E4861_, new_E4862_, new_E4863_,
    new_E4864_, new_E4865_, new_E4866_, new_E4867_, new_E4868_, new_E4869_,
    new_E4870_, new_E4871_, new_E4872_, new_E4873_, new_E4874_, new_E4875_,
    new_E4876_, new_E4877_, new_E4878_, new_E4879_, new_E4880_, new_E4881_,
    new_E4882_, new_E4883_, new_E4884_, new_E4885_, new_E4886_, new_E4887_,
    new_E4888_, new_E4889_, new_E4890_, new_E4891_, new_E4892_, new_E4893_,
    new_E4894_, new_E4895_, new_E4896_, new_E4897_, new_E4898_, new_E4899_,
    new_E4900_, new_E4901_, new_E4902_, new_E4903_, new_E4904_, new_E4905_,
    new_E4906_, new_E4907_, new_E4908_, new_E4909_, new_E4910_, new_E4911_,
    new_E4912_, new_E4913_, new_E4914_, new_E4915_, new_E4916_, new_E4917_,
    new_E4918_, new_E4919_, new_E4920_, new_E4921_, new_E4922_, new_E4923_,
    new_E4924_, new_E4925_, new_E4926_, new_E4927_, new_E4928_, new_E4929_,
    new_E4930_, new_E4931_, new_E4932_, new_E4933_, new_E4934_, new_E4935_,
    new_E4936_, new_E4937_, new_E4938_, new_E4939_, new_E4940_, new_E4941_,
    new_E4942_, new_E4943_, new_E4944_, new_E4945_, new_E4946_, new_E4947_,
    new_E4948_, new_E4949_, new_E4950_, new_E4951_, new_E4952_, new_E4953_,
    new_E4954_, new_E4955_, new_E4956_, new_E4957_, new_E4958_, new_E4959_,
    new_E4960_, new_E4961_, new_E4962_, new_E4963_, new_E4964_, new_E4965_,
    new_E4966_, new_E4967_, new_E4968_, new_E4969_, new_E4970_, new_E4971_,
    new_E4972_, new_E4973_, new_E4974_, new_E4975_, new_E4976_, new_E4977_,
    new_E4978_, new_E4979_, new_E4980_, new_E4981_, new_E4982_, new_E4983_,
    new_E4984_, new_E4985_, new_E4986_, new_E4987_, new_E4988_, new_E4989_,
    new_E4990_, new_E4991_, new_E4992_, new_E4993_, new_E4994_, new_E4995_,
    new_E4996_, new_E4997_, new_E4998_, new_E4999_, new_E5000_, new_E5001_,
    new_E5002_, new_E5003_, new_E5004_, new_E5005_, new_E5006_, new_E5007_,
    new_E5008_, new_E5009_, new_E5010_, new_E5011_, new_E5012_, new_E5013_,
    new_E5014_, new_E5015_, new_E5016_, new_E5017_, new_E5018_, new_E5019_,
    new_E5020_, new_E5021_, new_E5022_, new_E5023_, new_E5024_, new_E5025_,
    new_E5026_, new_E5027_, new_E5028_, new_E5029_, new_E5030_, new_E5031_,
    new_E5032_, new_E5033_, new_E5034_, new_E5035_, new_E5036_, new_E5037_,
    new_E5038_, new_E5039_, new_E5040_, new_E5041_, new_E5042_, new_E5043_,
    new_E5044_, new_E5045_, new_E5046_, new_E5047_, new_E5048_, new_E5049_,
    new_E5050_, new_E5051_, new_E5052_, new_E5053_, new_E5054_, new_E5055_,
    new_E5056_, new_E5057_, new_E5058_, new_E5059_, new_E5060_, new_E5061_,
    new_E5062_, new_E5063_, new_E5064_, new_E5065_, new_E5066_, new_E5067_,
    new_E5068_, new_E5069_, new_E5070_, new_E5071_, new_E5072_, new_E5073_,
    new_E5074_, new_E5075_, new_E5076_, new_E5077_, new_E5078_, new_E5079_,
    new_E5080_, new_E5081_, new_E5082_, new_E5083_, new_E5084_, new_E5085_,
    new_E5086_, new_E5087_, new_E5088_, new_E5089_, new_E5090_, new_E5091_,
    new_E5092_, new_E5093_, new_E5094_, new_E5095_, new_E5096_, new_E5097_,
    new_E5098_, new_E5099_, new_E5100_, new_E5101_, new_E5102_, new_E5103_,
    new_E5104_, new_E5105_, new_E5106_, new_E5107_, new_E5108_, new_E5109_,
    new_E5110_, new_E5111_, new_E5112_, new_E5113_, new_E5114_, new_E5115_,
    new_E5116_, new_E5117_, new_E5118_, new_E5119_, new_E5120_, new_E5121_,
    new_E5122_, new_E5123_, new_E5124_, new_E5125_, new_E5126_, new_E5127_,
    new_E5128_, new_E5129_, new_E5130_, new_E5131_, new_E5132_, new_E5133_,
    new_E5134_, new_E5135_, new_E5136_, new_E5137_, new_E5138_, new_E5139_,
    new_E5140_, new_E5141_, new_E5142_, new_E5143_, new_E5144_, new_E5145_,
    new_E5146_, new_E5147_, new_E5148_, new_E5149_, new_E5150_, new_E5151_,
    new_E5152_, new_E5153_, new_E5154_, new_E5155_, new_E5156_, new_E5157_,
    new_E5158_, new_E5159_, new_E5160_, new_E5161_, new_E5162_, new_E5163_,
    new_E5164_, new_E5165_, new_E5166_, new_E5167_, new_E5168_, new_E5169_,
    new_E5170_, new_E5171_, new_E5172_, new_E5173_, new_E5174_, new_E5175_,
    new_E5176_, new_E5177_, new_E5178_, new_E5179_, new_E5180_, new_E5181_,
    new_E5182_, new_E5183_, new_E5184_, new_E5185_, new_E5186_, new_E5187_,
    new_E5188_, new_E5189_, new_E5190_, new_E5191_, new_E5192_, new_E5193_,
    new_E5194_, new_E5195_, new_E5196_, new_E5197_, new_E5198_, new_E5199_,
    new_E5200_, new_E5201_, new_E5202_, new_E5203_, new_E5204_, new_E5205_,
    new_E5206_, new_E5207_, new_E5208_, new_E5209_, new_E5210_, new_E5211_,
    new_E5212_, new_E5213_, new_E5214_, new_E5215_, new_E5216_, new_E5217_,
    new_E5218_, new_E5219_, new_E5220_, new_E5221_, new_E5222_, new_E5223_,
    new_E5224_, new_E5225_, new_E5226_, new_E5227_, new_E5228_, new_E5229_,
    new_E5230_, new_E5231_, new_E5232_, new_E5233_, new_E5234_, new_E5235_,
    new_E5236_, new_E5237_, new_E5238_, new_E5239_, new_E5240_, new_E5241_,
    new_E5242_, new_E5243_, new_E5244_, new_E5245_, new_E5246_, new_E5247_,
    new_E5248_, new_E5249_, new_E5250_, new_E5251_, new_E5252_, new_E5253_,
    new_E5254_, new_E5255_, new_E5256_, new_E5257_, new_E5258_, new_E5259_,
    new_E5260_, new_E5261_, new_E5262_, new_E5263_, new_E5264_, new_E5265_,
    new_E5266_, new_E5267_, new_E5268_, new_E5269_, new_E5270_, new_E5271_,
    new_E5272_, new_E5273_, new_E5274_, new_E5275_, new_E5276_, new_E5277_,
    new_E5278_, new_E5279_, new_E5280_, new_E5281_, new_E5282_, new_E5283_,
    new_E5284_, new_E5285_, new_E5286_, new_E5287_, new_E5288_, new_E5289_,
    new_E5290_, new_E5291_, new_E5292_, new_E5293_, new_E5294_, new_E5295_,
    new_E5296_, new_E5297_, new_E5298_, new_E5299_, new_E5300_, new_E5301_,
    new_E5302_, new_E5303_, new_E5304_, new_E5305_, new_E5306_, new_E5307_,
    new_E5308_, new_E5309_, new_E5310_, new_E5311_, new_E5312_, new_E5313_,
    new_E5314_, new_E5315_, new_E5316_, new_E5317_, new_E5318_, new_E5319_,
    new_E5320_, new_E5321_, new_E5322_, new_E5323_, new_E5324_, new_E5325_,
    new_E5326_, new_E5327_, new_E5328_, new_E5329_, new_E5330_, new_E5331_,
    new_E5332_, new_E5333_, new_E5334_, new_E5335_, new_E5336_, new_E5337_,
    new_E5338_, new_E5339_, new_E5340_, new_E5341_, new_E5342_, new_E5343_,
    new_E5344_, new_E5345_, new_E5346_, new_E5347_, new_E5348_, new_E5349_,
    new_E5350_, new_E5351_, new_E5352_, new_E5353_, new_E5354_, new_E5355_,
    new_E5356_, new_E5357_, new_E5358_, new_E5359_, new_E5360_, new_E5361_,
    new_E5362_, new_E5363_, new_E5364_, new_E5365_, new_E5366_, new_E5367_,
    new_E5368_, new_E5369_, new_E5370_, new_E5371_, new_E5372_, new_E5373_,
    new_E5374_, new_E5375_, new_E5376_, new_E5377_, new_E5378_, new_E5379_,
    new_E5380_, new_E5381_, new_E5382_, new_E5383_, new_E5384_, new_E5385_,
    new_E5386_, new_E5387_, new_E5388_, new_E5389_, new_E5390_, new_E5391_,
    new_E5392_, new_E5393_, new_E5394_, new_E5395_, new_E5396_, new_E5397_,
    new_E5398_, new_E5399_, new_E5400_, new_E5401_, new_E5402_, new_E5403_,
    new_E5404_, new_E5405_, new_E5406_, new_E5407_, new_E5408_, new_E5409_,
    new_E5410_, new_E5411_, new_E5412_, new_E5413_, new_E5414_, new_E5415_,
    new_E5416_, new_E5417_, new_E5418_, new_E5419_, new_E5420_, new_E5421_,
    new_E5422_, new_E5423_, new_E5424_, new_E5425_, new_E5426_, new_E5427_,
    new_E5428_, new_E5429_, new_E5430_, new_E5431_, new_E5432_, new_E5433_,
    new_E5434_, new_E5435_, new_E5436_, new_E5437_, new_E5438_, new_E5439_,
    new_E5440_, new_E5441_, new_E5442_, new_E5443_, new_E5444_, new_E5445_,
    new_E5446_, new_E5447_, new_E5448_, new_E5449_, new_E5450_, new_E5451_,
    new_E5452_, new_E5453_, new_E5454_, new_E5455_, new_E5456_, new_E5457_,
    new_E5458_, new_E5459_, new_E5460_, new_E5461_, new_E5462_, new_E5463_,
    new_E5464_, new_E5465_, new_E5466_, new_E5467_, new_E5468_, new_E5469_,
    new_E5470_, new_E5471_, new_E5472_, new_E5473_, new_E5474_, new_E5475_,
    new_E5476_, new_E5477_, new_E5478_, new_E5479_, new_E5480_, new_E5481_,
    new_E5482_, new_E5483_, new_E5484_, new_E5485_, new_E5486_, new_E5487_,
    new_E5488_, new_E5489_, new_E5490_, new_E5491_, new_E5492_, new_E5493_,
    new_E5494_, new_E5495_, new_E5496_, new_E5497_, new_E5498_, new_E5499_,
    new_E5500_, new_E5501_, new_E5502_, new_E5503_, new_E5504_, new_E5505_,
    new_E5506_, new_E5507_, new_E5508_, new_E5509_, new_E5510_, new_E5511_,
    new_E5512_, new_E5513_, new_E5514_, new_E5515_, new_E5516_, new_E5517_,
    new_E5518_, new_E5519_, new_E5520_, new_E5521_, new_E5522_, new_E5523_,
    new_E5524_, new_E5525_, new_E5526_, new_E5527_, new_E5528_, new_E5529_,
    new_E5530_, new_E5531_, new_E5532_, new_E5533_, new_E5534_, new_E5535_,
    new_E5536_, new_E5537_, new_E5538_, new_E5539_, new_E5540_, new_E5541_,
    new_E5542_, new_E5543_, new_E5544_, new_E5545_, new_E5546_, new_E5547_,
    new_E5548_, new_E5549_, new_E5550_, new_E5551_, new_E5552_, new_E5553_,
    new_E5554_, new_E5555_, new_E5556_, new_E5557_, new_E5558_, new_E5559_,
    new_E5560_, new_E5561_, new_E5562_, new_E5563_, new_E5564_, new_E5565_,
    new_E5566_, new_E5567_, new_E5568_, new_E5569_, new_E5570_, new_E5571_,
    new_E5572_, new_E5573_, new_E5574_, new_E5575_, new_E5576_, new_E5577_,
    new_E5578_, new_E5579_, new_E5580_, new_E5581_, new_E5582_, new_E5583_,
    new_E5584_, new_E5585_, new_E5586_, new_E5587_, new_E5588_, new_E5589_,
    new_E5590_, new_E5591_, new_E5592_, new_E5593_, new_E5594_, new_E5595_,
    new_E5596_, new_E5597_, new_E5598_, new_E5599_, new_E5600_, new_E5601_,
    new_E5602_, new_E5603_, new_E5604_, new_E5605_, new_E5606_, new_E5607_,
    new_E5608_, new_E5609_, new_E5610_, new_E5611_, new_E5612_, new_E5613_,
    new_E5614_, new_E5615_, new_E5616_, new_E5617_, new_E5618_, new_E5619_,
    new_E5620_, new_E5621_, new_E5622_, new_E5623_, new_E5624_, new_E5625_,
    new_E5626_, new_E5627_, new_E5628_, new_E5629_, new_E5630_, new_E5631_,
    new_E5632_, new_E5633_, new_E5634_, new_E5635_, new_E5636_, new_E5637_,
    new_E5638_, new_E5639_, new_E5640_, new_E5641_, new_E5642_, new_E5643_,
    new_E5644_, new_E5645_, new_E5646_, new_E5647_, new_E5648_, new_E5649_,
    new_E5650_, new_E5651_, new_E5652_, new_E5653_, new_E5654_, new_E5655_,
    new_E5656_, new_E5657_, new_E5658_, new_E5659_, new_E5660_, new_E5661_,
    new_E5662_, new_E5663_, new_E5664_, new_E5665_, new_E5666_, new_E5667_,
    new_E5668_, new_E5669_, new_E5670_, new_E5671_, new_E5672_, new_E5673_,
    new_E5674_, new_E5675_, new_E5676_, new_E5677_, new_E5678_, new_E5679_,
    new_E5680_, new_E5681_, new_E5682_, new_E5683_, new_E5684_, new_E5685_,
    new_E5686_, new_E5687_, new_E5688_, new_E5689_, new_E5690_, new_E5691_,
    new_E5692_, new_E5693_, new_E5694_, new_E5695_, new_E5696_, new_E5697_,
    new_E5698_, new_E5699_, new_E5700_, new_E5701_, new_E5702_, new_E5703_,
    new_E5704_, new_E5705_, new_E5706_, new_E5707_, new_E5708_, new_E5709_,
    new_E5710_, new_E5711_, new_E5712_, new_E5713_, new_E5714_, new_E5715_,
    new_E5716_, new_E5717_, new_E5718_, new_E5719_, new_E5720_, new_E5721_,
    new_E5722_, new_E5723_, new_E5724_, new_E5725_, new_E5726_, new_E5727_,
    new_E5728_, new_E5729_, new_E5730_, new_E5731_, new_E5732_, new_E5733_,
    new_E5734_, new_E5735_, new_E5736_, new_E5737_, new_E5738_, new_E5739_,
    new_E5740_, new_E5741_, new_E5742_, new_E5743_, new_E5744_, new_E5745_,
    new_E5746_, new_E5747_, new_E5748_, new_E5749_, new_E5750_, new_E5751_,
    new_E5752_, new_E5753_, new_E5754_, new_E5755_, new_E5756_, new_E5757_,
    new_E5758_, new_E5759_, new_E5760_, new_E5761_, new_E5762_, new_E5763_,
    new_E5764_, new_E5765_, new_E5766_, new_E5767_, new_E5768_, new_E5769_,
    new_E5770_, new_E5771_, new_E5772_, new_E5773_, new_E5774_, new_E5775_,
    new_E5776_, new_E5777_, new_E5778_, new_E5779_, new_E5780_, new_E5781_,
    new_E5782_, new_E5783_, new_E5784_, new_E5785_, new_E5786_, new_E5787_,
    new_E5788_, new_E5789_, new_E5790_, new_E5791_, new_E5792_, new_E5793_,
    new_E5794_, new_E5795_, new_E5796_, new_E5797_, new_E5798_, new_E5799_,
    new_E5800_, new_E5801_, new_E5802_, new_E5803_, new_E5804_, new_E5805_,
    new_E5806_, new_E5807_, new_E5808_, new_E5809_, new_E5810_, new_E5811_,
    new_E5812_, new_E5813_, new_E5814_, new_E5815_, new_E5816_, new_E5817_,
    new_E5818_, new_E5819_, new_E5820_, new_E5821_, new_E5822_, new_E5823_,
    new_E5824_, new_E5825_, new_E5826_, new_E5827_, new_E5828_, new_E5829_,
    new_E5830_, new_E5831_, new_E5832_, new_E5833_, new_E5834_, new_E5835_,
    new_E5836_, new_E5837_, new_E5838_, new_E5839_, new_E5840_, new_E5841_,
    new_E5842_, new_E5843_, new_E5844_, new_E5845_, new_E5846_, new_E5847_,
    new_E5848_, new_E5849_, new_E5850_, new_E5851_, new_E5852_, new_E5853_,
    new_E5854_, new_E5855_, new_E5856_, new_E5857_, new_E5858_, new_E5859_,
    new_E5860_, new_E5861_, new_E5862_, new_E5863_, new_E5864_, new_E5865_,
    new_E5866_, new_E5867_, new_E5868_, new_E5869_, new_E5870_, new_E5871_,
    new_E5872_, new_E5873_, new_E5874_, new_E5875_, new_E5876_, new_E5877_,
    new_E5878_, new_E5879_, new_E5880_, new_E5881_, new_E5882_, new_E5883_,
    new_E5884_, new_E5885_, new_E5886_, new_E5887_, new_E5888_, new_E5889_,
    new_E5890_, new_E5891_, new_E5892_, new_E5893_, new_E5894_, new_E5895_,
    new_E5896_, new_E5897_, new_E5898_, new_E5899_, new_E5900_, new_E5901_,
    new_E5902_, new_E5903_, new_E5904_, new_E5905_, new_E5906_, new_E5907_,
    new_E5908_, new_E5909_, new_E5910_, new_E5911_, new_E5912_, new_E5913_,
    new_E5914_, new_E5915_, new_E5916_, new_E5917_, new_E5918_, new_E5919_,
    new_E5920_, new_E5921_, new_E5922_, new_E5923_, new_E5924_, new_E5925_,
    new_E5926_, new_E5927_, new_E5928_, new_E5929_, new_E5930_, new_E5931_,
    new_E5932_, new_E5933_, new_E5934_, new_E5935_, new_E5936_, new_E5937_,
    new_E5938_, new_E5939_, new_E5940_, new_E5941_, new_E5942_, new_E5943_,
    new_E5944_, new_E5945_, new_E5946_, new_E5947_, new_E5948_, new_E5949_,
    new_E5950_, new_E5951_, new_E5952_, new_E5953_, new_E5954_, new_E5955_,
    new_E5956_, new_E5957_, new_E5958_, new_E5959_, new_E5960_, new_E5961_,
    new_E5962_, new_E5963_, new_E5964_, new_E5965_, new_E5966_, new_E5967_,
    new_E5968_, new_E5969_, new_E5970_, new_E5971_, new_E5972_, new_E5973_,
    new_E5974_, new_E5975_, new_E5976_, new_E5977_, new_E5978_, new_E5979_,
    new_E5980_, new_E5981_, new_E5982_, new_E5983_, new_E5984_, new_E5985_,
    new_E5986_, new_E5987_, new_E5988_, new_E5989_, new_E5990_, new_E5991_,
    new_E5992_, new_E5993_, new_E5994_, new_E5995_, new_E5996_, new_E5997_,
    new_E5998_, new_E5999_, new_E6000_, new_E6001_, new_E6002_, new_E6003_,
    new_E6004_, new_E6005_, new_E6006_, new_E6007_, new_E6008_, new_E6009_,
    new_E6010_, new_E6011_, new_E6012_, new_E6013_, new_E6014_, new_E6015_,
    new_E6016_, new_E6017_, new_E6018_, new_E6019_, new_E6020_, new_E6021_,
    new_E6022_, new_E6023_, new_E6024_, new_E6025_, new_E6026_, new_E6027_,
    new_E6028_, new_E6029_, new_E6030_, new_E6031_, new_E6032_, new_E6033_,
    new_E6034_, new_E6035_, new_E6036_, new_E6037_, new_E6038_, new_E6039_,
    new_E6040_, new_E6041_, new_E6042_, new_E6043_, new_E6044_, new_E6045_,
    new_E6046_, new_E6047_, new_E6048_, new_E6049_, new_E6050_, new_E6051_,
    new_E6052_, new_E6053_, new_E6054_, new_E6055_, new_E6056_, new_E6057_,
    new_E6058_, new_E6059_, new_E6060_, new_E6061_, new_E6062_, new_E6063_,
    new_E6064_, new_E6065_, new_E6066_, new_E6067_, new_E6068_, new_E6069_,
    new_E6070_, new_E6071_, new_E6072_, new_E6073_, new_E6074_, new_E6075_,
    new_E6076_, new_E6077_, new_E6078_, new_E6079_, new_E6080_, new_E6081_,
    new_E6082_, new_E6083_, new_E6084_, new_E6085_, new_E6086_, new_E6087_,
    new_E6088_, new_E6089_, new_E6090_, new_E6091_, new_E6092_, new_E6093_,
    new_E6094_, new_E6095_, new_E6096_, new_E6097_, new_E6098_, new_E6099_,
    new_E6100_, new_E6101_, new_E6102_, new_E6103_, new_E6104_, new_E6105_,
    new_E6106_, new_E6107_, new_E6108_, new_E6109_, new_E6110_, new_E6111_,
    new_E6112_, new_E6113_, new_E6114_, new_E6115_, new_E6116_, new_E6117_,
    new_E6118_, new_E6119_, new_E6120_, new_E6121_, new_E6122_, new_E6123_,
    new_E6124_, new_E6125_, new_E6126_, new_E6127_, new_E6128_, new_E6129_,
    new_E6130_, new_E6131_, new_E6132_, new_E6133_, new_E6134_, new_E6135_,
    new_E6136_, new_E6137_, new_E6138_, new_E6139_, new_E6140_, new_E6141_,
    new_E6142_, new_E6143_, new_E6144_, new_E6145_, new_E6146_, new_E6147_,
    new_E6148_, new_E6149_, new_E6150_, new_E6151_, new_E6152_, new_E6153_,
    new_E6154_, new_E6155_, new_E6156_, new_E6157_, new_E6158_, new_E6159_,
    new_E6160_, new_E6161_, new_E6162_, new_E6163_, new_E6164_, new_E6165_,
    new_E6166_, new_E6167_, new_E6168_, new_E6169_, new_E6170_, new_E6171_,
    new_E6172_, new_E6173_, new_E6174_, new_E6175_, new_E6176_, new_E6177_,
    new_E6178_, new_E6179_, new_E6180_, new_E6181_, new_E6182_, new_E6183_,
    new_E6184_, new_E6185_, new_E6186_, new_E6187_, new_E6188_, new_E6189_,
    new_E6190_, new_E6191_, new_E6192_, new_E6193_, new_E6194_, new_E6195_,
    new_E6196_, new_E6197_, new_E6198_, new_E6199_, new_E6200_, new_E6201_,
    new_E6202_, new_E6203_, new_E6204_, new_E6205_, new_E6206_, new_E6207_,
    new_E6208_, new_E6209_, new_E6210_, new_E6211_, new_E6212_, new_E6213_,
    new_E6214_, new_E6215_, new_E6216_, new_E6217_, new_E6218_, new_E6219_,
    new_E6220_, new_E6221_, new_E6222_, new_E6223_, new_E6224_, new_E6225_,
    new_E6226_, new_E6227_, new_E6228_, new_E6229_, new_E6230_, new_E6231_,
    new_E6232_, new_E6233_, new_E6234_, new_E6235_, new_E6236_, new_E6237_,
    new_E6238_, new_E6239_, new_E6240_, new_E6241_, new_E6242_, new_E6243_,
    new_E6244_, new_E6245_, new_E6246_, new_E6247_, new_E6248_, new_E6249_,
    new_E6250_, new_E6251_, new_E6252_, new_E6253_, new_E6254_, new_E6255_,
    new_E6256_, new_E6257_, new_E6258_, new_E6259_, new_E6260_, new_E6261_,
    new_E6262_, new_E6263_, new_E6264_, new_E6265_, new_E6266_, new_E6267_,
    new_E6268_, new_E6269_, new_E6270_, new_E6271_, new_E6272_, new_E6273_,
    new_E6274_, new_E6275_, new_E6276_, new_E6277_, new_E6278_, new_E6279_,
    new_E6280_, new_E6281_, new_E6282_, new_E6283_, new_E6284_, new_E6285_,
    new_E6286_, new_E6287_, new_E6288_, new_E6289_, new_E6290_, new_E6291_,
    new_E6292_, new_E6293_, new_E6294_, new_E6295_, new_E6296_, new_E6297_,
    new_E6298_, new_E6299_, new_E6300_, new_E6301_, new_E6302_, new_E6303_,
    new_E6304_, new_E6305_, new_E6306_, new_E6307_, new_E6308_, new_E6309_,
    new_E6310_, new_E6311_, new_E6312_, new_E6313_, new_E6314_, new_E6315_,
    new_E6316_, new_E6317_, new_E6318_, new_E6319_, new_E6320_, new_E6321_,
    new_E6322_, new_E6323_, new_E6324_, new_E6325_, new_E6326_, new_E6327_,
    new_E6328_, new_E6329_, new_E6330_, new_E6331_, new_E6332_, new_E6333_,
    new_E6334_, new_E6335_, new_E6336_, new_E6337_, new_E6338_, new_E6339_,
    new_E6340_, new_E6341_, new_E6342_, new_E6343_, new_E6344_, new_E6345_,
    new_E6346_, new_E6347_, new_E6348_, new_E6349_, new_E6350_, new_E6351_,
    new_E6352_, new_E6353_, new_E6354_, new_E6355_, new_E6356_, new_E6357_,
    new_E6358_, new_E6359_, new_E6360_, new_E6361_, new_E6362_, new_E6363_,
    new_E6364_, new_E6365_, new_E6366_, new_E6367_, new_E6368_, new_E6369_,
    new_E6370_, new_E6371_, new_E6372_, new_E6373_, new_E6374_, new_E6375_,
    new_E6376_, new_E6377_, new_E6378_, new_E6379_, new_E6380_, new_E6381_,
    new_E6382_, new_E6383_, new_E6384_, new_E6385_, new_E6386_, new_E6387_,
    new_E6388_, new_E6389_, new_E6390_, new_E6391_, new_E6392_, new_E6393_,
    new_E6394_, new_E6395_, new_E6396_, new_E6397_, new_E6398_, new_E6399_,
    new_E6400_, new_E6401_, new_E6402_, new_E6403_, new_E6404_, new_E6405_,
    new_E6406_, new_E6407_, new_E6408_, new_E6409_, new_E6410_, new_E6411_,
    new_E6412_, new_E6413_, new_E6414_, new_E6415_, new_E6416_, new_E6417_,
    new_E6418_, new_E6419_, new_E6420_, new_E6421_, new_E6422_, new_E6423_,
    new_E6424_, new_E6425_, new_E6426_, new_E6427_, new_E6428_, new_E6429_,
    new_E6430_, new_E6431_, new_E6432_, new_E6433_, new_E6434_, new_E6435_,
    new_E6436_, new_E6437_, new_E6438_, new_E6439_, new_E6440_, new_E6441_,
    new_E6442_, new_E6443_, new_E6444_, new_E6445_, new_E6446_, new_E6447_,
    new_E6448_, new_E6449_, new_E6450_, new_E6451_, new_E6452_, new_E6453_,
    new_E6454_, new_E6455_, new_E6456_, new_E6457_, new_E6458_, new_E6459_,
    new_E6460_, new_E6461_, new_E6462_, new_E6463_, new_E6464_, new_E6465_,
    new_E6466_, new_E6467_, new_E6468_, new_E6469_, new_E6470_, new_E6471_,
    new_E6472_, new_E6473_, new_E6474_, new_E6475_, new_E6476_, new_E6477_,
    new_E6478_, new_E6479_, new_E6480_, new_E6481_, new_E6482_, new_E6483_,
    new_E6484_, new_E6485_, new_E6486_, new_E6487_, new_E6488_, new_E6489_,
    new_E6490_, new_E6491_, new_E6492_, new_E6493_, new_E6494_, new_E6495_,
    new_E6496_, new_E6497_, new_E6498_, new_E6499_, new_E6500_, new_E6501_,
    new_E6502_, new_E6503_, new_E6504_, new_E6505_, new_E6506_, new_E6507_,
    new_E6508_, new_E6509_, new_E6510_, new_E6511_, new_E6512_, new_E6513_,
    new_E6514_, new_E6515_, new_E6516_, new_E6517_, new_E6518_, new_E6519_,
    new_E6520_, new_E6521_, new_E6522_, new_E6523_, new_E6524_, new_E6525_,
    new_E6526_, new_E6527_, new_E6528_, new_E6529_, new_E6530_, new_E6531_,
    new_E6532_, new_E6533_, new_E6534_, new_E6535_, new_E6536_, new_E6537_,
    new_E6538_, new_E6539_, new_E6540_, new_E6541_, new_E6542_, new_E6543_,
    new_E6544_, new_E6545_, new_E6546_, new_E6547_, new_E6548_, new_E6549_,
    new_E6550_, new_E6551_, new_E6552_, new_E6553_, new_E6554_, new_E6555_,
    new_E6556_, new_E6557_, new_E6558_, new_E6559_, new_E6560_, new_E6561_,
    new_E6562_, new_E6563_, new_E6564_, new_E6565_, new_E6566_, new_E6567_,
    new_E6568_, new_E6569_, new_E6570_, new_E6571_, new_E6572_, new_E6573_,
    new_E6574_, new_E6575_, new_E6576_, new_E6577_, new_E6578_, new_E6579_,
    new_E6580_, new_E6581_, new_E6582_, new_E6583_, new_E6584_, new_E6585_,
    new_E6586_, new_E6587_, new_E6588_, new_E6589_, new_E6590_, new_E6591_,
    new_E6592_, new_E6593_, new_E6594_, new_E6595_, new_E6596_, new_E6597_,
    new_E6598_, new_E6599_, new_E6600_, new_E6601_, new_E6602_, new_E6603_,
    new_E6604_, new_E6605_, new_E6606_, new_E6607_, new_E6608_, new_E6609_,
    new_E6610_, new_E6611_, new_E6612_, new_E6613_, new_E6614_, new_E6615_,
    new_E6616_, new_E6617_, new_E6618_, new_E6619_, new_E6620_, new_E6621_,
    new_E6622_, new_E6623_, new_E6624_, new_E6625_, new_E6626_, new_E6627_,
    new_E6628_, new_E6629_, new_E6630_, new_E6631_, new_E6632_, new_E6633_,
    new_E6634_, new_E6635_, new_E6636_, new_E6637_, new_E6638_, new_E6639_,
    new_E6640_, new_E6641_, new_E6642_, new_E6643_, new_E6644_, new_E6645_,
    new_E6646_, new_E6647_, new_E6648_, new_E6649_, new_E6650_, new_E6651_,
    new_E6652_, new_E6653_, new_E6654_, new_E6655_, new_E6656_, new_E6657_,
    new_E6658_, new_E6659_, new_E6660_, new_E6661_, new_E6662_, new_E6663_,
    new_E6664_, new_E6665_, new_E6666_, new_E6667_, new_E6668_, new_E6669_,
    new_E6670_, new_E6671_, new_E6672_, new_E6673_, new_E6674_, new_E6675_,
    new_E6676_, new_E6677_, new_E6678_, new_E6679_, new_E6680_, new_E6681_,
    new_E6682_, new_E6683_, new_E6684_, new_E6685_, new_E6686_, new_E6687_,
    new_E6688_, new_E6689_, new_E6690_, new_E6691_, new_E6692_, new_E6693_,
    new_E6694_, new_E6695_, new_E6696_, new_E6697_, new_E6698_, new_E6699_,
    new_E6700_, new_E6701_, new_E6702_, new_E6703_, new_E6704_, new_E6705_,
    new_E6706_, new_E6707_, new_E6708_, new_E6709_, new_E6710_, new_E6711_,
    new_E6712_, new_E6713_, new_E6714_, new_E6715_, new_E6716_, new_E6717_,
    new_E6718_, new_E6719_, new_E6720_, new_E6721_, new_E6722_, new_E6723_,
    new_E6724_, new_E6725_, new_E6726_, new_E6727_, new_E6728_, new_E6729_,
    new_E6730_, new_E6731_, new_E6732_, new_E6733_, new_E6734_, new_E6735_,
    new_E6736_, new_E6737_, new_E6738_, new_E6739_, new_E6740_, new_E6741_,
    new_E6742_, new_E6743_, new_E6744_, new_E6745_, new_E6746_, new_E6747_,
    new_E6748_, new_E6749_, new_E6750_, new_E6751_, new_E6752_, new_E6753_,
    new_E6754_, new_E6755_, new_E6756_, new_E6757_, new_E6758_, new_E6759_,
    new_E6760_, new_E6761_, new_E6762_, new_E6763_, new_E6764_, new_E6765_,
    new_E6766_, new_E6767_, new_E6768_, new_E6769_, new_E6770_, new_E6771_,
    new_E6772_, new_E6773_, new_E6774_, new_E6775_, new_E6776_, new_E6777_,
    new_E6778_, new_E6779_, new_E6780_, new_E6781_, new_E6782_, new_E6783_,
    new_E6784_, new_E6785_, new_E6786_, new_E6787_, new_E6788_, new_E6789_,
    new_E6790_, new_E6791_, new_E6792_, new_E6793_, new_E6794_, new_E6795_,
    new_E6796_, new_E6797_, new_E6798_, new_E6799_, new_E6800_, new_E6801_,
    new_E6802_, new_E6803_, new_E6804_, new_E6805_, new_E6806_, new_E6807_,
    new_E6808_, new_E6809_, new_E6810_, new_E6811_, new_E6812_, new_E6813_,
    new_E6814_, new_E6815_, new_E6816_, new_E6817_, new_E6818_, new_E6819_,
    new_E6820_, new_E6821_, new_E6822_, new_E6823_, new_E6824_, new_E6825_,
    new_E6826_, new_E6827_, new_E6828_, new_E6829_, new_E6830_, new_E6831_,
    new_E6832_, new_E6833_, new_E6834_, new_E6835_, new_E6836_, new_E6837_,
    new_E6838_, new_E6839_, new_E6840_, new_E6841_, new_E6842_, new_E6843_,
    new_E6844_, new_E6845_, new_E6846_, new_E6847_, new_E6848_, new_E6849_,
    new_E6850_, new_E6851_, new_E6852_, new_E6853_, new_E6854_, new_E6855_,
    new_E6856_, new_E6857_, new_E6858_, new_E6859_, new_E6860_, new_E6861_,
    new_E6862_, new_E6863_, new_E6864_, new_E6865_, new_E6866_, new_E6867_,
    new_E6868_, new_E6869_, new_E6870_, new_E6871_, new_E6872_, new_E6873_,
    new_E6874_, new_E6875_, new_E6876_, new_E6877_, new_E6878_, new_E6879_,
    new_E6880_, new_E6881_, new_E6882_, new_E6883_, new_E6884_, new_E6885_,
    new_E6886_, new_E6887_, new_E6888_, new_E6889_, new_E6890_, new_E6891_,
    new_E6892_, new_E6893_, new_E6894_, new_E6895_, new_E6896_, new_E6897_,
    new_E6898_, new_E6899_, new_E6900_, new_E6901_, new_E6902_, new_E6903_,
    new_E6904_, new_E6905_, new_E6906_, new_E6907_, new_E6908_, new_E6909_,
    new_E6910_, new_E6911_, new_E6912_, new_E6913_, new_E6914_, new_E6915_,
    new_E6916_, new_E6917_, new_E6918_, new_E6919_, new_E6920_, new_E6921_,
    new_E6922_, new_E6923_, new_E6924_, new_E6925_, new_E6926_, new_E6927_,
    new_E6928_, new_E6929_, new_E6930_, new_E6931_, new_E6932_, new_E6933_,
    new_E6934_, new_E6935_, new_E6936_, new_E6937_, new_E6938_, new_E6939_,
    new_E6940_, new_E6941_, new_E6942_, new_E6943_, new_E6944_, new_E6945_,
    new_E6946_, new_E6947_, new_E6948_, new_E6949_, new_E6950_, new_E6951_,
    new_E6952_, new_E6953_, new_E6954_, new_E6955_, new_E6956_, new_E6957_,
    new_E6958_, new_E6959_, new_E6960_, new_E6961_, new_E6962_, new_E6963_,
    new_E6964_, new_E6965_, new_E6966_, new_E6967_, new_E6968_, new_E6969_,
    new_E6970_, new_E6971_, new_E6972_, new_E6973_, new_E6974_, new_E6975_,
    new_E6976_, new_E6977_, new_E6978_, new_E6979_, new_E6980_, new_E6981_,
    new_E6982_, new_E6983_, new_E6984_, new_E6985_, new_E6986_, new_E6987_,
    new_E6988_, new_E6989_, new_E6990_, new_E6991_, new_E6992_, new_E6993_,
    new_E6994_, new_E6995_, new_E6996_, new_E6997_, new_E6998_, new_E6999_,
    new_E7000_, new_E7001_, new_E7002_, new_E7003_, new_E7004_, new_E7005_,
    new_E7006_, new_E7007_, new_E7008_, new_E7009_, new_E7010_, new_E7011_,
    new_E7012_, new_E7013_, new_E7014_, new_E7015_, new_E7016_, new_E7017_,
    new_E7018_, new_E7019_, new_E7020_, new_E7021_, new_E7022_, new_E7023_,
    new_E7024_, new_E7025_, new_E7026_, new_E7027_, new_E7028_, new_E7029_,
    new_E7030_, new_E7031_, new_E7032_, new_E7033_, new_E7034_, new_E7035_,
    new_E7036_, new_E7037_, new_E7038_, new_E7039_, new_E7040_, new_E7041_,
    new_E7042_, new_E7043_, new_E7044_, new_E7045_, new_E7046_, new_E7047_,
    new_E7048_, new_E7049_, new_E7050_, new_E7051_, new_E7052_, new_E7053_,
    new_E7054_, new_E7055_, new_E7056_, new_E7057_, new_E7058_, new_E7059_,
    new_E7060_, new_E7061_, new_E7062_, new_E7063_, new_E7064_, new_E7065_,
    new_E7066_, new_E7067_, new_E7068_, new_E7069_, new_E7070_, new_E7071_,
    new_E7072_, new_E7073_, new_E7074_, new_E7075_, new_E7076_, new_E7077_,
    new_E7078_, new_E7079_, new_E7080_, new_E7081_, new_E7082_, new_E7083_,
    new_E7084_, new_E7085_, new_E7086_, new_E7087_, new_E7088_, new_E7089_,
    new_E7090_, new_E7091_, new_E7092_, new_E7093_, new_E7094_, new_E7095_,
    new_E7096_, new_E7097_, new_E7098_, new_E7099_, new_E7100_, new_E7101_,
    new_E7102_, new_E7103_, new_E7104_, new_E7105_, new_E7106_, new_E7107_,
    new_E7108_, new_E7109_, new_E7110_, new_E7111_, new_E7112_, new_E7113_,
    new_E7114_, new_E7115_, new_E7116_, new_E7117_, new_E7118_, new_E7119_,
    new_E7120_, new_E7121_, new_E7122_, new_E7123_, new_E7124_, new_E7125_,
    new_E7126_, new_E7127_, new_E7128_, new_E7129_, new_E7130_, new_E7131_,
    new_E7132_, new_E7133_, new_E7134_, new_E7135_, new_E7136_, new_E7137_,
    new_E7138_, new_E7139_, new_E7140_, new_E7141_, new_E7142_, new_E7143_,
    new_E7144_, new_E7145_, new_E7146_, new_E7147_, new_E7148_, new_E7149_,
    new_E7150_, new_E7151_, new_E7152_, new_E7153_, new_E7154_, new_E7155_,
    new_E7156_, new_E7157_, new_E7158_, new_E7159_, new_E7160_, new_E7161_,
    new_E7162_, new_E7163_, new_E7164_, new_E7165_, new_E7166_, new_E7167_,
    new_E7168_, new_E7169_, new_E7170_, new_E7171_, new_E7172_, new_E7173_,
    new_E7174_, new_E7175_, new_E7176_, new_E7177_, new_E7178_, new_E7179_,
    new_E7180_, new_E7181_, new_E7182_, new_E7183_, new_E7184_, new_E7185_,
    new_E7186_, new_E7187_, new_E7188_, new_E7189_, new_E7190_, new_E7191_,
    new_E7192_, new_E7193_, new_E7194_, new_E7195_, new_E7196_, new_E7197_,
    new_E7198_, new_E7199_, new_E7200_, new_E7201_, new_E7202_, new_E7203_,
    new_E7204_, new_E7205_, new_E7206_, new_E7207_, new_E7208_, new_E7209_,
    new_E7210_, new_E7211_, new_E7212_, new_E7213_, new_E7214_, new_E7215_,
    new_E7216_, new_E7217_, new_E7218_, new_E7219_, new_E7220_, new_E7221_,
    new_E7222_, new_E7223_, new_E7224_, new_E7225_, new_E7226_, new_E7227_,
    new_E7228_, new_E7229_, new_E7230_, new_E7231_, new_E7232_, new_E7233_,
    new_E7234_, new_E7235_, new_E7236_, new_E7237_, new_E7238_, new_E7239_,
    new_E7240_, new_E7241_, new_E7242_, new_E7243_, new_E7244_, new_E7245_,
    new_E7246_, new_E7247_, new_E7248_, new_E7249_, new_E7250_, new_E7251_,
    new_E7252_, new_E7253_, new_E7254_, new_E7255_, new_E7256_, new_E7257_,
    new_E7258_, new_E7259_, new_E7260_, new_E7261_, new_E7262_, new_E7263_,
    new_E7264_, new_E7265_, new_E7266_, new_E7267_, new_E7268_, new_E7269_,
    new_E7270_, new_E7271_, new_E7272_, new_E7273_, new_E7274_, new_E7275_,
    new_E7276_, new_E7277_, new_E7278_, new_E7279_, new_E7280_, new_E7281_,
    new_E7282_, new_E7283_, new_E7284_, new_E7285_, new_E7286_, new_E7287_,
    new_E7288_, new_E7289_, new_E7290_, new_E7291_, new_E7292_, new_E7293_,
    new_E7294_, new_E7295_, new_E7296_, new_E7297_, new_E7298_, new_E7299_,
    new_E7300_, new_E7301_, new_E7302_, new_E7303_, new_E7304_, new_E7305_,
    new_E7306_, new_E7307_, new_E7308_, new_E7309_, new_E7310_, new_E7311_,
    new_E7312_, new_E7313_, new_E7314_, new_E7315_, new_E7316_, new_E7317_,
    new_E7318_, new_E7319_, new_E7320_, new_E7321_, new_E7322_, new_E7323_,
    new_E7324_, new_E7325_, new_E7326_, new_E7327_, new_E7328_, new_E7329_,
    new_E7330_, new_E7331_, new_E7332_, new_E7333_, new_E7334_, new_E7335_,
    new_E7336_, new_E7337_, new_E7338_, new_E7339_, new_E7340_, new_E7341_,
    new_E7342_, new_E7343_, new_E7344_, new_E7345_, new_E7346_, new_E7347_,
    new_E7348_, new_E7349_, new_E7350_, new_E7351_, new_E7352_, new_E7353_,
    new_E7354_, new_E7355_, new_E7356_, new_E7357_, new_E7358_, new_E7359_,
    new_E7360_, new_E7361_, new_E7362_, new_E7363_, new_E7364_, new_E7365_,
    new_E7366_, new_E7367_, new_E7368_, new_E7369_, new_E7370_, new_E7371_,
    new_E7372_, new_E7373_, new_E7374_, new_E7375_, new_E7376_, new_E7377_,
    new_E7378_, new_E7379_, new_E7380_, new_E7381_, new_E7382_, new_E7383_,
    new_E7384_, new_E7385_, new_E7386_, new_E7387_, new_E7388_, new_E7389_,
    new_E7390_, new_E7391_, new_E7392_, new_E7393_, new_E7394_, new_E7395_,
    new_E7396_, new_E7397_, new_E7398_, new_E7399_, new_E7400_, new_E7401_,
    new_E7402_, new_E7403_, new_E7404_, new_E7405_, new_E7406_, new_E7407_,
    new_E7408_, new_E7409_, new_E7410_, new_E7411_, new_E7412_, new_E7413_,
    new_E7414_, new_E7415_, new_E7416_, new_E7417_, new_E7418_, new_E7419_,
    new_E7420_, new_E7421_, new_E7422_, new_E7423_, new_E7424_, new_E7425_,
    new_E7426_, new_E7427_, new_E7428_, new_E7429_, new_E7430_, new_E7431_,
    new_E7432_, new_E7433_, new_E7434_, new_E7435_, new_E7436_, new_E7437_,
    new_E7438_, new_E7439_, new_E7440_, new_E7441_, new_E7442_, new_E7443_,
    new_E7444_, new_E7445_, new_E7446_, new_E7447_, new_E7448_, new_E7449_,
    new_E7450_, new_E7451_, new_E7452_, new_E7453_, new_E7454_, new_E7455_,
    new_E7456_, new_E7457_, new_E7458_, new_E7459_, new_E7460_, new_E7461_,
    new_E7462_, new_E7463_, new_E7464_, new_E7465_, new_E7466_, new_E7467_,
    new_E7468_, new_E7469_, new_E7470_, new_E7471_, new_E7472_, new_E7473_,
    new_E7474_, new_E7475_, new_E7476_, new_E7477_, new_E7478_, new_E7479_,
    new_E7480_, new_E7481_, new_E7482_, new_E7483_, new_E7484_, new_E7485_,
    new_E7486_, new_E7487_, new_E7488_, new_E7489_, new_E7490_, new_E7491_,
    new_E7492_, new_E7493_, new_E7494_, new_E7495_, new_E7496_, new_E7497_,
    new_E7498_, new_E7499_, new_E7500_, new_E7501_, new_E7502_, new_E7503_,
    new_E7504_, new_E7505_, new_E7506_, new_E7507_, new_E7508_, new_E7509_,
    new_E7510_, new_E7511_, new_E7512_, new_E7513_, new_E7514_, new_E7515_,
    new_E7516_, new_E7517_, new_E7518_, new_E7519_, new_E7520_, new_E7521_,
    new_E7522_, new_E7523_, new_E7524_, new_E7525_, new_E7526_, new_E7527_,
    new_E7528_, new_E7529_, new_E7530_, new_E7531_, new_E7532_, new_E7533_,
    new_E7534_, new_E7535_, new_E7536_, new_E7537_, new_E7538_, new_E7539_,
    new_E7540_, new_E7541_, new_E7542_, new_E7543_, new_E7544_, new_E7545_,
    new_E7546_, new_E7547_, new_E7548_, new_E7549_, new_E7550_, new_E7551_,
    new_E7552_, new_E7553_, new_E7554_, new_E7555_, new_E7556_, new_E7557_,
    new_E7558_, new_E7559_, new_E7560_, new_E7561_, new_E7562_, new_E7563_,
    new_E7564_, new_E7565_, new_E7566_, new_E7567_, new_E7568_, new_E7569_,
    new_E7570_, new_E7571_, new_E7572_, new_E7573_, new_E7574_, new_E7575_,
    new_E7576_, new_E7577_, new_E7578_, new_E7579_, new_E7580_, new_E7581_,
    new_E7582_, new_E7583_, new_E7584_, new_E7585_, new_E7586_, new_E7587_,
    new_E7588_, new_E7589_, new_E7590_, new_E7591_, new_E7592_, new_E7593_,
    new_E7594_, new_E7595_, new_E7596_, new_E7597_, new_E7598_, new_E7599_,
    new_E7600_, new_E7601_, new_E7602_, new_E7603_, new_E7604_, new_E7605_,
    new_E7606_, new_E7607_, new_E7608_, new_E7609_, new_E7610_, new_E7611_,
    new_E7612_, new_E7613_, new_E7614_, new_E7615_, new_E7616_, new_E7617_,
    new_E7618_, new_E7619_, new_E7620_, new_E7621_, new_E7622_, new_E7623_,
    new_E7624_, new_E7625_, new_E7626_, new_E7627_, new_E7628_, new_E7629_,
    new_E7630_, new_E7631_, new_E7632_, new_E7633_, new_E7634_, new_E7635_,
    new_E7636_, new_E7637_, new_E7638_, new_E7639_, new_E7640_, new_E7641_,
    new_E7642_, new_E7643_, new_E7644_, new_E7645_, new_E7646_, new_E7647_,
    new_E7648_, new_E7649_, new_E7650_, new_E7651_, new_E7652_, new_E7653_,
    new_E7654_, new_E7655_, new_E7656_, new_E7657_, new_E7658_, new_E7659_,
    new_E7660_, new_E7661_, new_E7662_, new_E7663_, new_E7664_, new_E7665_,
    new_E7666_, new_E7667_, new_E7668_, new_E7669_, new_E7670_, new_E7671_,
    new_E7672_, new_E7673_, new_E7674_, new_E7675_, new_E7676_, new_E7677_,
    new_E7678_, new_E7679_, new_E7680_, new_E7681_, new_E7682_, new_E7683_,
    new_E7684_, new_E7685_, new_E7686_, new_E7687_, new_E7688_, new_E7689_,
    new_E7690_, new_E7691_, new_E7692_, new_E7693_, new_E7694_, new_E7695_,
    new_E7696_, new_E7697_, new_E7698_, new_E7699_, new_E7700_, new_E7701_,
    new_E7702_, new_E7703_, new_E7704_, new_E7705_, new_E7706_, new_E7707_,
    new_E7708_, new_E7709_, new_E7710_, new_E7711_, new_E7712_, new_E7713_,
    new_E7714_, new_E7715_, new_E7716_, new_E7717_, new_E7718_, new_E7719_,
    new_E7720_, new_E7721_, new_E7722_, new_E7723_, new_E7724_, new_E7725_,
    new_E7726_, new_E7727_, new_E7728_, new_E7729_, new_E7730_, new_E7731_,
    new_E7732_, new_E7733_, new_E7734_, new_E7735_, new_E7736_, new_E7737_,
    new_E7738_, new_E7739_, new_E7740_, new_E7741_, new_E7742_, new_E7743_,
    new_E7744_, new_E7745_, new_E7746_, new_E7747_, new_E7748_, new_E7749_,
    new_E7750_, new_E7751_, new_E7752_, new_E7753_, new_E7754_, new_E7755_,
    new_E7756_, new_E7757_, new_E7758_, new_E7759_, new_E7760_, new_E7761_,
    new_E7762_, new_E7763_, new_E7764_, new_E7765_, new_E7766_, new_E7767_,
    new_E7768_, new_E7769_, new_E7770_, new_E7771_, new_E7772_, new_E7773_,
    new_E7774_, new_E7775_, new_E7776_, new_E7777_, new_E7778_, new_E7779_,
    new_E7780_, new_E7781_, new_E7782_, new_E7783_, new_E7784_, new_E7785_,
    new_E7786_, new_E7787_, new_E7788_, new_E7789_, new_E7790_, new_E7791_,
    new_E7792_, new_E7793_, new_E7794_, new_E7795_, new_E7796_, new_E7797_,
    new_E7798_, new_E7799_, new_E7800_, new_E7801_, new_E7802_, new_E7803_,
    new_E7804_, new_E7805_, new_E7806_, new_E7807_, new_E7808_, new_E7809_,
    new_E7810_, new_E7811_, new_E7812_, new_E7813_, new_E7814_, new_E7815_,
    new_E7816_, new_E7817_, new_E7818_, new_E7819_, new_E7820_, new_E7821_,
    new_E7822_, new_E7823_, new_E7824_, new_E7825_, new_E7826_, new_E7827_,
    new_E7828_, new_E7829_, new_E7830_, new_E7831_, new_E7832_, new_E7833_,
    new_E7834_, new_E7835_, new_E7836_, new_E7837_, new_E7838_, new_E7839_,
    new_E7840_, new_E7841_, new_E7842_, new_E7843_, new_E7844_, new_E7845_,
    new_E7846_, new_E7847_, new_E7848_, new_E7849_, new_E7850_, new_E7851_,
    new_E7852_, new_E7853_, new_E7854_, new_E7855_, new_E7856_, new_E7857_,
    new_E7858_, new_E7859_, new_E7860_, new_E7861_, new_E7862_, new_E7863_,
    new_E7864_, new_E7865_, new_E7866_, new_E7867_, new_E7868_, new_E7869_,
    new_E7870_, new_E7871_, new_E7872_, new_E7873_, new_E7874_, new_E7875_,
    new_E7876_, new_E7877_, new_E7878_, new_E7879_, new_E7880_, new_E7881_,
    new_E7882_, new_E7883_, new_E7884_, new_E7885_, new_E7886_, new_E7887_,
    new_E7888_, new_E7889_, new_E7890_, new_E7891_, new_E7892_, new_E7893_,
    new_E7894_, new_E7895_, new_E7896_, new_E7897_, new_E7898_, new_E7899_,
    new_E7900_, new_E7901_, new_E7902_, new_E7903_, new_E7904_, new_E7905_,
    new_E7906_, new_E7907_, new_E7908_, new_E7909_, new_E7910_, new_E7911_,
    new_E7912_, new_E7913_, new_E7914_, new_E7915_, new_E7916_, new_E7917_,
    new_E7918_, new_E7919_, new_E7920_, new_E7921_, new_E7922_, new_E7923_,
    new_E7924_, new_E7925_, new_E7926_, new_E7927_, new_E7928_, new_E7929_,
    new_E7930_, new_E7931_, new_E7932_, new_E7933_, new_E7934_, new_E7935_,
    new_E7936_, new_E7937_, new_E7938_, new_E7939_, new_E7940_, new_E7941_,
    new_E7942_, new_E7943_, new_E7944_, new_E7945_, new_E7946_, new_E7947_,
    new_E7948_, new_E7949_, new_E7950_, new_E7951_, new_E7952_, new_E7953_,
    new_E7954_, new_E7955_, new_E7956_, new_E7957_, new_E7958_, new_E7959_,
    new_E7960_, new_E7961_, new_E7962_, new_E7963_, new_E7964_, new_E7965_,
    new_E7966_, new_E7967_, new_E7968_, new_E7969_, new_E7970_, new_E7971_,
    new_E7972_, new_E7973_, new_E7974_, new_E7975_, new_E7976_, new_E7977_,
    new_E7978_, new_E7979_, new_E7980_, new_E7981_, new_E7982_, new_E7983_,
    new_E7984_, new_E7985_, new_E7986_, new_E7987_, new_E7988_, new_E7989_,
    new_E7990_, new_E7991_, new_E7992_, new_E7993_, new_E7994_, new_E7995_,
    new_E7996_, new_E7997_, new_E7998_, new_E7999_, new_E8000_, new_E8001_,
    new_E8002_, new_E8003_, new_E8004_, new_E8005_, new_E8006_, new_E8007_,
    new_E8008_, new_E8009_, new_E8010_, new_E8011_, new_E8012_, new_E8013_,
    new_E8014_, new_E8015_, new_E8016_, new_E8017_, new_E8018_, new_E8019_,
    new_E8020_, new_E8021_, new_E8022_, new_E8023_, new_E8024_, new_E8025_,
    new_E8026_, new_E8027_, new_E8028_, new_E8029_, new_E8030_, new_E8031_,
    new_E8032_, new_E8033_, new_E8034_, new_E8035_, new_E8036_, new_E8037_,
    new_E8038_, new_E8039_, new_E8040_, new_E8041_, new_E8042_, new_E8043_,
    new_E8044_, new_E8045_, new_E8046_, new_E8047_, new_E8048_, new_E8049_,
    new_E8050_, new_E8051_, new_E8052_, new_E8053_, new_E8054_, new_E8055_,
    new_E8056_, new_E8057_, new_E8058_, new_E8059_, new_E8060_, new_E8061_,
    new_E8062_, new_E8063_, new_E8064_, new_E8065_, new_E8066_, new_E8067_,
    new_E8068_, new_E8069_, new_E8070_, new_E8071_, new_E8072_, new_E8073_,
    new_E8074_, new_E8075_, new_E8076_, new_E8077_, new_E8078_, new_E8079_,
    new_E8080_, new_E8081_, new_E8082_, new_E8083_, new_E8084_, new_E8085_,
    new_E8086_, new_E8087_, new_E8088_, new_E8089_, new_E8090_, new_E8091_,
    new_E8092_, new_E8093_, new_E8094_, new_E8095_, new_E8096_, new_E8097_,
    new_E8098_, new_E8099_, new_E8100_, new_E8101_, new_E8102_, new_E8103_,
    new_E8104_, new_E8105_, new_E8106_, new_E8107_, new_E8108_, new_E8109_,
    new_E8110_, new_E8111_, new_E8112_, new_E8113_, new_E8114_, new_E8115_,
    new_E8116_, new_E8117_, new_E8118_, new_E8119_, new_E8120_, new_E8121_,
    new_E8122_, new_E8123_, new_E8124_, new_E8125_, new_E8126_, new_E8127_,
    new_E8128_, new_E8129_, new_E8130_, new_E8131_, new_E8132_, new_E8133_,
    new_E8134_, new_E8135_, new_E8136_, new_E8137_, new_E8138_, new_E8139_,
    new_E8140_, new_E8141_, new_E8142_, new_E8143_, new_E8144_, new_E8145_,
    new_E8146_, new_E8147_, new_E8148_, new_E8149_, new_E8150_, new_E8151_,
    new_E8152_, new_E8153_, new_E8154_, new_E8155_, new_E8156_, new_E8157_,
    new_E8158_, new_E8159_, new_E8160_, new_E8161_, new_E8162_, new_E8163_,
    new_E8164_, new_E8165_, new_E8166_, new_E8167_, new_E8168_, new_E8169_,
    new_E8170_, new_E8171_, new_E8172_, new_E8173_, new_E8174_, new_E8175_,
    new_E8176_, new_E8177_, new_E8178_, new_E8179_, new_E8180_, new_E8181_,
    new_E8182_, new_E8183_, new_E8184_, new_E8185_, new_E8186_, new_E8187_,
    new_E8188_, new_E8189_, new_E8190_, new_E8191_, new_E8192_, new_E8193_,
    new_E8194_, new_E8195_, new_E8196_, new_E8197_, new_E8198_, new_E8199_,
    new_E8200_, new_E8201_, new_E8202_, new_E8203_, new_E8204_, new_E8205_,
    new_E8206_, new_E8207_, new_E8208_, new_E8209_, new_E8210_, new_E8211_,
    new_E8212_, new_E8213_, new_E8214_, new_E8215_, new_E8216_, new_E8217_,
    new_E8218_, new_E8219_, new_E8220_, new_E8221_, new_E8222_, new_E8223_,
    new_E8224_, new_E8225_, new_E8226_, new_E8227_, new_E8228_, new_E8229_,
    new_E8230_, new_E8231_, new_E8232_, new_E8233_, new_E8234_, new_E8235_,
    new_E8236_, new_E8237_, new_E8238_, new_E8239_, new_E8240_, new_E8241_,
    new_E8242_, new_E8243_, new_E8244_, new_E8245_, new_E8246_, new_E8247_,
    new_E8248_, new_E8249_, new_E8250_, new_E8251_, new_E8252_, new_E8253_,
    new_E8254_, new_E8255_, new_E8256_, new_E8257_, new_E8258_, new_E8259_,
    new_E8260_, new_E8261_, new_E8262_, new_E8263_, new_E8264_, new_E8265_,
    new_E8266_, new_E8267_, new_E8268_, new_E8269_, new_E8270_, new_E8271_,
    new_E8272_, new_E8273_, new_E8274_, new_E8275_, new_E8276_, new_E8277_,
    new_E8278_, new_E8279_, new_E8280_, new_E8281_, new_E8282_, new_E8283_,
    new_E8284_, new_E8285_, new_E8286_, new_E8287_, new_E8288_, new_E8289_,
    new_E8290_, new_E8291_, new_E8292_, new_E8293_, new_E8294_, new_E8295_,
    new_E8296_, new_E8297_, new_E8298_, new_E8299_, new_E8300_, new_E8301_,
    new_E8302_, new_E8303_, new_E8304_, new_E8305_, new_E8306_, new_E8307_,
    new_E8308_, new_E8309_, new_E8310_, new_E8311_, new_E8312_, new_E8313_,
    new_E8314_, new_E8315_, new_E8316_, new_E8317_, new_E8318_, new_E8319_,
    new_E8320_, new_E8321_, new_E8322_, new_E8323_, new_E8324_, new_E8325_,
    new_E8326_, new_E8327_, new_E8328_, new_E8329_, new_E8330_, new_E8331_,
    new_E8332_, new_E8333_, new_E8334_, new_E8335_, new_E8336_, new_E8337_,
    new_E8338_, new_E8339_, new_E8340_, new_E8341_, new_E8342_, new_E8343_,
    new_E8344_, new_E8345_, new_E8346_, new_E8347_, new_E8348_, new_E8349_,
    new_E8350_, new_E8351_, new_E8352_, new_E8353_, new_E8354_, new_E8355_,
    new_E8356_, new_E8357_, new_E8358_, new_E8359_, new_E8360_, new_E8361_,
    new_E8362_, new_E8363_, new_E8364_, new_E8365_, new_E8366_, new_E8367_,
    new_E8368_, new_E8369_, new_E8370_, new_E8371_, new_E8372_, new_E8373_,
    new_E8374_, new_E8375_, new_E8376_, new_E8377_, new_E8378_, new_E8379_,
    new_E8380_, new_E8381_, new_E8382_, new_E8383_, new_E8384_, new_E8385_,
    new_E8386_, new_E8387_, new_E8388_, new_E8389_, new_E8390_, new_E8391_,
    new_E8392_, new_E8393_, new_E8394_, new_E8395_, new_E8396_, new_E8397_,
    new_E8398_, new_E8399_, new_E8400_, new_E8401_, new_E8402_, new_E8403_,
    new_E8404_, new_E8405_, new_E8406_, new_E8407_, new_E8408_, new_E8409_,
    new_E8410_, new_E8411_, new_E8412_, new_E8413_, new_E8414_, new_E8415_,
    new_E8416_, new_E8417_, new_E8418_, new_E8419_, new_E8420_, new_E8421_,
    new_E8422_, new_E8423_, new_E8424_, new_E8425_, new_E8426_, new_E8427_,
    new_E8428_, new_E8429_, new_E8430_, new_E8431_, new_E8432_, new_E8433_,
    new_E8434_, new_E8435_, new_E8436_, new_E8437_, new_E8438_, new_E8439_,
    new_E8440_, new_E8441_, new_E8442_, new_E8443_, new_E8444_, new_E8445_,
    new_E8446_, new_E8447_, new_E8448_, new_E8449_, new_E8450_, new_E8451_,
    new_E8452_, new_E8453_, new_E8454_, new_E8455_, new_E8456_, new_E8457_,
    new_E8458_, new_E8459_, new_E8460_, new_E8461_, new_E8462_, new_E8463_,
    new_E8464_, new_E8465_, new_E8466_, new_E8467_, new_E8468_, new_E8469_,
    new_E8470_, new_E8471_, new_E8472_, new_E8473_, new_E8474_, new_E8475_,
    new_E8476_, new_E8477_, new_E8478_, new_E8479_, new_E8480_, new_E8481_,
    new_E8482_, new_E8483_, new_E8484_, new_E8485_, new_E8486_, new_E8487_,
    new_E8488_, new_E8489_, new_E8490_, new_E8491_, new_E8492_, new_E8493_,
    new_E8494_, new_E8495_, new_E8496_, new_E8497_, new_E8498_, new_E8499_,
    new_E8500_, new_E8501_, new_E8502_, new_E8503_, new_E8504_, new_E8505_,
    new_E8506_, new_E8507_, new_E8508_, new_E8509_, new_E8510_, new_E8511_,
    new_E8512_, new_E8513_, new_E8514_, new_E8515_, new_E8516_, new_E8517_,
    new_E8518_, new_E8519_, new_E8520_, new_E8521_, new_E8522_, new_E8523_,
    new_E8524_, new_E8525_, new_E8526_, new_E8527_, new_E8528_, new_E8529_,
    new_E8530_, new_E8531_, new_E8532_, new_E8533_, new_E8534_, new_E8535_,
    new_E8536_, new_E8537_, new_E8538_, new_E8539_, new_E8540_, new_E8541_,
    new_E8542_, new_E8543_, new_E8544_, new_E8545_, new_E8546_, new_E8547_,
    new_E8548_, new_E8549_, new_E8550_, new_E8551_, new_E8552_, new_E8553_,
    new_E8554_, new_E8555_, new_E8556_, new_E8557_, new_E8558_, new_E8559_,
    new_E8560_, new_E8561_, new_E8562_, new_E8563_, new_E8564_, new_E8565_,
    new_E8566_, new_E8567_, new_E8568_, new_E8569_, new_E8570_, new_E8571_,
    new_E8572_, new_E8573_, new_E8574_, new_E8575_, new_E8576_, new_E8577_,
    new_E8578_, new_E8579_, new_E8580_, new_E8581_, new_E8582_, new_E8583_,
    new_E8584_, new_E8585_, new_E8586_, new_E8587_, new_E8588_, new_E8589_,
    new_E8590_, new_E8591_, new_E8592_, new_E8593_, new_E8594_, new_E8595_,
    new_E8596_, new_E8597_, new_E8598_, new_E8599_, new_E8600_, new_E8601_,
    new_E8602_, new_E8603_, new_E8604_, new_E8605_, new_E8606_, new_E8607_,
    new_E8608_, new_E8609_, new_E8610_, new_E8611_, new_E8612_, new_E8613_,
    new_E8614_, new_E8615_, new_E8616_, new_E8617_, new_E8618_, new_E8619_,
    new_E8620_, new_E8621_, new_E8622_, new_E8623_, new_E8624_, new_E8625_,
    new_E8626_, new_E8627_, new_E8628_, new_E8629_, new_E8630_, new_E8631_,
    new_E8632_, new_E8633_, new_E8634_, new_E8635_, new_E8636_, new_E8637_,
    new_E8638_, new_E8639_, new_E8640_, new_E8641_, new_E8642_, new_E8643_,
    new_E8644_, new_E8645_, new_E8646_, new_E8647_, new_E8648_, new_E8649_,
    new_E8650_, new_E8651_, new_E8652_, new_E8653_, new_E8654_, new_E8655_,
    new_E8656_, new_E8657_, new_E8658_, new_E8659_, new_E8660_, new_E8661_,
    new_E8662_, new_E8663_, new_E8664_, new_E8665_, new_E8666_, new_E8667_,
    new_E8668_, new_E8669_, new_E8670_, new_E8671_, new_E8672_, new_E8673_,
    new_E8674_, new_E8675_, new_E8676_, new_E8677_, new_E8678_, new_E8679_,
    new_E8680_, new_E8681_, new_E8682_, new_E8683_, new_E8684_, new_E8685_,
    new_E8686_, new_E8687_, new_E8688_, new_E8689_, new_E8690_, new_E8691_,
    new_E8692_, new_E8693_, new_E8694_, new_E8695_, new_E8696_, new_E8697_,
    new_E8698_, new_E8699_, new_E8700_, new_E8701_, new_E8702_, new_E8703_,
    new_E8704_, new_E8705_, new_E8706_, new_E8707_, new_E8708_, new_E8709_,
    new_E8710_, new_E8711_, new_E8712_, new_E8713_, new_E8714_, new_E8715_,
    new_E8716_, new_E8717_, new_E8718_, new_E8719_, new_E8720_, new_E8721_,
    new_E8722_, new_E8723_, new_E8724_, new_E8725_, new_E8726_, new_E8727_,
    new_E8728_, new_E8729_, new_E8730_, new_E8731_, new_E8732_, new_E8733_,
    new_E8734_, new_E8735_, new_E8736_, new_E8737_, new_E8738_, new_E8739_,
    new_E8740_, new_E8741_, new_E8742_, new_E8743_, new_E8744_, new_E8745_,
    new_E8746_, new_E8747_, new_E8748_, new_E8749_, new_E8750_, new_E8751_,
    new_E8752_, new_E8753_, new_E8754_, new_E8755_, new_E8756_, new_E8757_,
    new_E8758_, new_E8759_, new_E8760_, new_E8761_, new_E8762_, new_E8763_,
    new_E8764_, new_E8765_, new_E8766_, new_E8767_, new_E8768_, new_E8769_,
    new_E8770_, new_E8771_, new_E8772_, new_E8773_, new_E8774_, new_E8775_,
    new_E8776_, new_E8777_, new_E8778_, new_E8779_, new_E8780_, new_E8781_,
    new_E8782_, new_E8783_, new_E8784_, new_E8785_, new_E8786_, new_E8787_,
    new_E8788_, new_E8789_, new_E8790_, new_E8791_, new_E8792_, new_E8793_,
    new_E8794_, new_E8795_, new_E8796_, new_E8797_, new_E8798_, new_E8799_,
    new_E8800_, new_E8801_, new_E8802_, new_E8803_, new_E8804_, new_E8805_,
    new_E8806_, new_E8807_, new_E8808_, new_E8809_, new_E8810_, new_E8811_,
    new_E8812_, new_E8813_, new_E8814_, new_E8815_, new_E8816_, new_E8817_,
    new_E8818_, new_E8819_, new_E8820_, new_E8821_, new_E8822_, new_E8823_,
    new_E8824_, new_E8825_, new_E8826_, new_E8827_, new_E8828_, new_E8829_,
    new_E8830_, new_E8831_, new_E8832_, new_E8833_, new_E8834_, new_E8835_,
    new_E8836_, new_E8837_, new_E8838_, new_E8839_, new_E8840_, new_E8841_,
    new_E8842_, new_E8843_, new_E8844_, new_E8845_, new_E8846_, new_E8847_,
    new_E8848_, new_E8849_, new_E8850_, new_E8851_, new_E8852_, new_E8853_,
    new_E8854_, new_E8855_, new_E8856_, new_E8857_, new_E8858_, new_E8859_,
    new_E8860_, new_E8861_, new_E8862_, new_E8863_, new_E8864_, new_E8865_,
    new_E8866_, new_E8867_, new_E8868_, new_E8869_, new_E8870_, new_E8871_,
    new_E8872_, new_E8873_, new_E8874_, new_E8875_, new_E8876_, new_E8877_,
    new_E8878_, new_E8879_, new_E8880_, new_E8881_, new_E8882_, new_E8883_,
    new_E8884_, new_E8885_, new_E8886_, new_E8887_, new_E8888_, new_E8889_,
    new_E8890_, new_E8891_, new_E8892_, new_E8893_, new_E8894_, new_E8895_,
    new_E8896_, new_E8897_, new_E8898_, new_E8899_, new_E8900_, new_E8901_,
    new_E8902_, new_E8903_, new_E8904_, new_E8905_, new_E8906_, new_E8907_,
    new_E8908_, new_E8909_, new_E8910_, new_E8911_, new_E8912_, new_E8913_,
    new_E8914_, new_E8915_, new_E8916_, new_E8917_, new_E8918_, new_E8919_,
    new_E8920_, new_E8921_, new_E8922_, new_E8923_, new_E8924_, new_E8925_,
    new_E8926_, new_E8927_, new_E8928_, new_E8929_, new_E8930_, new_E8931_,
    new_E8932_, new_E8933_, new_E8934_, new_E8935_, new_E8936_, new_E8937_,
    new_E8938_, new_E8939_, new_E8940_, new_E8941_, new_E8942_, new_E8943_,
    new_E8944_, new_E8945_, new_E8946_, new_E8947_, new_E8948_, new_E8949_,
    new_E8950_, new_E8951_, new_E8952_, new_E8953_, new_E8954_, new_E8955_,
    new_E8956_, new_E8957_, new_E8958_, new_E8959_, new_E8960_, new_E8961_,
    new_E8962_, new_E8963_, new_E8964_, new_E8965_, new_E8966_, new_E8967_,
    new_E8968_, new_E8969_, new_E8970_, new_E8971_, new_E8972_, new_E8973_,
    new_E8974_, new_E8975_, new_E8976_, new_E8977_, new_E8978_, new_E8979_,
    new_E8980_, new_E8981_, new_E8982_, new_E8983_, new_E8984_, new_E8985_,
    new_E8986_, new_E8987_, new_E8988_, new_E8989_, new_E8990_, new_E8991_,
    new_E8992_, new_E8993_, new_E8994_, new_E8995_, new_E8996_, new_E8997_,
    new_E8998_, new_E8999_, new_E9000_, new_E9001_, new_E9002_, new_E9003_,
    new_E9004_, new_E9005_, new_E9006_, new_E9007_, new_E9008_, new_E9009_,
    new_E9010_, new_E9011_, new_E9012_, new_E9013_, new_E9014_, new_E9015_,
    new_E9016_, new_E9017_, new_E9018_, new_E9019_, new_E9020_, new_E9021_,
    new_E9022_, new_E9023_, new_E9024_, new_E9025_, new_E9026_, new_E9027_,
    new_E9028_, new_E9029_, new_E9030_, new_E9031_, new_E9032_, new_E9033_,
    new_E9034_, new_E9035_, new_E9036_, new_E9037_, new_E9038_, new_E9039_,
    new_E9040_, new_E9041_, new_E9042_, new_E9043_, new_E9044_, new_E9045_,
    new_E9046_, new_E9047_, new_E9048_, new_E9049_, new_E9050_, new_E9051_,
    new_E9052_, new_E9053_, new_E9054_, new_E9055_, new_E9056_, new_E9057_,
    new_E9058_, new_E9059_, new_E9060_, new_E9061_, new_E9062_, new_E9063_,
    new_E9064_, new_E9065_, new_E9066_, new_E9067_, new_E9068_, new_E9069_,
    new_E9070_, new_E9071_, new_E9072_, new_E9073_, new_E9074_, new_E9075_,
    new_E9076_, new_E9077_, new_E9078_, new_E9079_, new_E9080_, new_E9081_,
    new_E9082_, new_E9083_, new_E9084_, new_E9085_, new_E9086_, new_E9087_,
    new_E9088_, new_E9089_, new_E9090_, new_E9091_, new_E9092_, new_E9093_,
    new_E9094_, new_E9095_, new_E9096_, new_E9097_, new_E9098_, new_E9099_,
    new_E9100_, new_E9101_, new_E9102_, new_E9103_, new_E9104_, new_E9105_,
    new_E9106_, new_E9107_, new_E9108_, new_E9109_, new_E9110_, new_E9111_,
    new_E9112_, new_E9113_, new_E9114_, new_E9115_, new_E9116_, new_E9117_,
    new_E9118_, new_E9119_, new_E9120_, new_E9121_, new_E9122_, new_E9123_,
    new_E9124_, new_E9125_, new_E9126_, new_E9127_, new_E9128_, new_E9129_,
    new_E9130_, new_E9131_, new_E9132_, new_E9133_, new_E9134_, new_E9135_,
    new_E9136_, new_E9137_, new_E9138_, new_E9139_, new_E9140_, new_E9141_,
    new_E9142_, new_E9143_, new_E9144_, new_E9145_, new_E9146_, new_E9147_,
    new_E9148_, new_E9149_, new_E9150_, new_E9151_, new_E9152_, new_E9153_,
    new_E9154_, new_E9155_, new_E9156_, new_E9157_, new_E9158_, new_E9159_,
    new_E9160_, new_E9161_, new_E9162_, new_E9163_, new_E9164_, new_E9165_,
    new_E9166_, new_E9167_, new_E9168_, new_E9169_, new_E9170_, new_E9171_,
    new_E9172_, new_E9173_, new_E9174_, new_E9175_, new_E9176_, new_E9177_,
    new_E9178_, new_E9179_, new_E9180_, new_E9181_, new_E9182_, new_E9183_,
    new_E9184_, new_E9185_, new_E9186_, new_E9187_, new_E9188_, new_E9189_,
    new_E9190_, new_E9191_, new_E9192_, new_E9193_, new_E9194_, new_E9195_,
    new_E9196_, new_E9197_, new_E9198_, new_E9199_, new_E9200_, new_E9201_,
    new_E9202_, new_E9203_, new_E9204_, new_E9205_, new_E9206_, new_E9207_,
    new_E9208_, new_E9209_, new_E9210_, new_E9211_, new_E9212_, new_E9213_,
    new_E9214_, new_E9215_, new_E9216_, new_E9217_, new_E9218_, new_E9219_,
    new_E9220_, new_E9221_, new_E9222_, new_E9223_, new_E9224_, new_E9225_,
    new_E9226_, new_E9227_, new_E9228_, new_E9229_, new_E9230_, new_E9231_,
    new_E9232_, new_E9233_, new_E9234_, new_E9235_, new_E9236_, new_E9237_,
    new_E9238_, new_E9239_, new_E9240_, new_E9241_, new_E9242_, new_E9243_,
    new_E9244_, new_E9245_, new_E9246_, new_E9247_, new_E9248_, new_E9249_,
    new_E9250_, new_E9251_, new_E9252_, new_E9253_, new_E9254_, new_E9255_,
    new_E9256_, new_E9257_, new_E9258_, new_E9259_, new_E9260_, new_E9261_,
    new_E9262_, new_E9263_, new_E9264_, new_E9265_, new_E9266_, new_E9267_,
    new_E9268_, new_E9269_, new_E9270_, new_E9271_, new_E9272_, new_E9273_,
    new_E9274_, new_E9275_, new_E9276_, new_E9277_, new_E9278_, new_E9279_,
    new_E9280_, new_E9281_, new_E9282_, new_E9283_, new_E9284_, new_E9285_,
    new_E9286_, new_E9287_, new_E9288_, new_E9289_, new_E9290_, new_E9291_,
    new_E9292_, new_E9293_, new_E9294_, new_E9295_, new_E9296_, new_E9297_,
    new_E9298_, new_E9299_, new_E9300_, new_E9301_, new_E9302_, new_E9303_,
    new_E9304_, new_E9305_, new_E9306_, new_E9307_, new_E9308_, new_E9309_,
    new_E9310_, new_E9311_, new_E9312_, new_E9313_, new_E9314_, new_E9315_,
    new_E9316_, new_E9317_, new_E9318_, new_E9319_, new_E9320_, new_E9321_,
    new_E9322_, new_E9323_, new_E9324_, new_E9325_, new_E9326_, new_E9327_,
    new_E9328_, new_E9329_, new_E9330_, new_E9331_, new_E9332_, new_E9333_,
    new_E9334_, new_E9335_, new_E9336_, new_E9337_, new_E9338_, new_E9339_,
    new_E9340_, new_E9341_, new_E9342_, new_E9343_, new_E9344_, new_E9345_,
    new_E9346_, new_E9347_, new_E9348_, new_E9349_, new_E9350_, new_E9351_,
    new_E9352_, new_E9353_, new_E9354_, new_E9355_, new_E9356_, new_E9357_,
    new_E9358_, new_E9359_, new_E9360_, new_E9361_, new_E9362_, new_E9363_,
    new_E9364_, new_E9365_, new_E9366_, new_E9367_, new_E9368_, new_E9369_,
    new_E9370_, new_E9371_, new_E9372_, new_E9373_, new_E9374_, new_E9375_,
    new_E9376_, new_E9377_, new_E9378_, new_E9379_, new_E9380_, new_E9381_,
    new_E9382_, new_E9383_, new_E9384_, new_E9385_, new_E9386_, new_E9387_,
    new_E9388_, new_E9389_, new_E9390_, new_E9391_, new_E9392_, new_E9393_,
    new_E9394_, new_E9395_, new_E9396_, new_E9397_, new_E9398_, new_E9399_,
    new_E9400_, new_E9401_, new_E9402_, new_E9403_, new_E9404_, new_E9405_,
    new_E9406_, new_E9407_, new_E9408_, new_E9409_, new_E9410_, new_E9411_,
    new_E9412_, new_E9413_, new_E9414_, new_E9415_, new_E9416_, new_E9417_,
    new_E9418_, new_E9419_, new_E9420_, new_E9421_, new_E9422_, new_E9423_,
    new_E9424_, new_E9425_, new_E9426_, new_E9427_, new_E9428_, new_E9429_,
    new_E9430_, new_E9431_, new_E9432_, new_E9433_, new_E9434_, new_E9435_,
    new_E9436_, new_E9437_, new_E9438_, new_E9439_, new_E9440_, new_E9441_,
    new_E9442_, new_E9443_, new_E9444_, new_E9445_, new_E9446_, new_E9447_,
    new_E9448_, new_E9449_, new_E9450_, new_E9451_, new_E9452_, new_E9453_,
    new_E9454_, new_E9455_, new_E9456_, new_E9457_, new_E9458_, new_E9459_,
    new_E9460_, new_E9461_, new_E9462_, new_E9463_, new_E9464_, new_E9465_,
    new_E9466_, new_E9467_, new_E9468_, new_E9469_, new_E9470_, new_E9471_,
    new_E9472_, new_E9473_, new_E9474_, new_E9475_, new_E9476_, new_E9477_,
    new_E9478_, new_E9479_, new_E9480_, new_E9481_, new_E9482_, new_E9483_,
    new_E9484_, new_E9485_, new_E9486_, new_E9487_, new_E9488_, new_E9489_,
    new_E9490_, new_E9491_, new_E9492_, new_E9493_, new_E9494_, new_E9495_,
    new_E9496_, new_E9497_, new_E9498_, new_E9499_, new_E9500_, new_E9501_,
    new_E9502_, new_E9503_, new_E9504_, new_E9505_, new_E9506_, new_E9507_,
    new_E9508_, new_E9509_, new_E9510_, new_E9511_, new_E9512_, new_E9513_,
    new_E9514_, new_E9515_, new_E9516_, new_E9517_, new_E9518_, new_E9519_,
    new_E9520_, new_E9521_, new_E9522_, new_E9523_, new_E9524_, new_E9525_,
    new_E9526_, new_E9527_, new_E9528_, new_E9529_, new_E9530_, new_E9531_,
    new_E9532_, new_E9533_, new_E9534_, new_E9535_, new_E9536_, new_E9537_,
    new_E9538_, new_E9539_, new_E9540_, new_E9541_, new_E9542_, new_E9543_,
    new_E9544_, new_E9545_, new_E9546_, new_E9547_, new_E9548_, new_E9549_,
    new_E9550_, new_E9551_, new_E9552_, new_E9553_, new_E9554_, new_E9555_,
    new_E9556_, new_E9557_, new_E9558_, new_E9559_, new_E9560_, new_E9561_,
    new_E9562_, new_E9563_, new_E9564_, new_E9565_, new_E9566_, new_E9567_,
    new_E9568_, new_E9569_, new_E9570_, new_E9571_, new_E9572_, new_E9573_,
    new_E9574_, new_E9575_, new_E9576_, new_E9577_, new_E9578_, new_E9579_,
    new_E9580_, new_E9581_, new_E9582_, new_E9583_, new_E9584_, new_E9585_,
    new_E9586_, new_E9587_, new_E9588_, new_E9589_, new_E9590_, new_E9591_,
    new_E9592_, new_E9593_, new_E9594_, new_E9595_, new_E9596_, new_E9597_,
    new_E9598_, new_E9599_, new_E9600_, new_E9601_, new_E9602_, new_E9603_,
    new_E9604_, new_E9605_, new_E9606_, new_E9607_, new_E9608_, new_E9609_,
    new_E9610_, new_E9611_, new_E9612_, new_E9613_, new_E9614_, new_E9615_,
    new_E9616_, new_E9617_, new_E9618_, new_E9619_, new_E9620_, new_E9621_,
    new_E9622_, new_E9623_, new_E9624_, new_E9625_, new_E9626_, new_E9627_,
    new_E9628_, new_E9629_, new_E9630_, new_E9631_, new_E9632_, new_E9633_,
    new_E9634_, new_E9635_, new_E9636_, new_E9637_, new_E9638_, new_E9639_,
    new_E9640_, new_E9641_, new_E9642_, new_E9643_, new_E9644_, new_E9645_,
    new_E9646_, new_E9647_, new_E9648_, new_E9649_, new_E9650_, new_E9651_,
    new_E9652_, new_E9653_, new_E9654_, new_E9655_, new_E9656_, new_E9657_,
    new_E9658_, new_E9659_, new_E9660_, new_E9661_, new_E9662_, new_E9663_,
    new_E9664_, new_E9665_, new_E9666_, new_E9667_, new_E9668_, new_E9669_,
    new_E9670_, new_E9671_, new_E9672_, new_E9673_, new_E9674_, new_E9675_,
    new_E9676_, new_E9677_, new_E9678_, new_E9679_, new_E9680_, new_E9681_,
    new_E9682_, new_E9683_, new_E9684_, new_E9685_, new_E9686_, new_E9687_,
    new_E9688_, new_E9689_, new_E9690_, new_E9691_, new_E9692_, new_E9693_,
    new_E9694_, new_E9695_, new_E9696_, new_E9697_, new_E9698_, new_E9699_,
    new_E9700_, new_E9701_, new_E9702_, new_E9703_, new_E9704_, new_E9705_,
    new_E9706_, new_E9707_, new_E9708_, new_E9709_, new_E9710_, new_E9711_,
    new_E9712_, new_E9713_, new_E9714_, new_E9715_, new_E9716_, new_E9717_,
    new_E9718_, new_E9719_, new_E9720_, new_E9721_, new_E9722_, new_E9723_,
    new_E9724_, new_E9725_, new_E9726_, new_E9727_, new_E9728_, new_E9729_,
    new_E9730_, new_E9731_, new_E9732_, new_E9733_, new_E9734_, new_E9735_,
    new_E9736_, new_E9737_, new_E9738_, new_E9739_, new_E9740_, new_E9741_,
    new_E9742_, new_E9743_, new_E9744_, new_E9745_, new_E9746_, new_E9747_,
    new_E9748_, new_E9749_, new_E9750_, new_E9751_, new_E9752_, new_E9753_,
    new_E9754_, new_E9755_, new_E9756_, new_E9757_, new_E9758_, new_E9759_,
    new_E9760_, new_E9761_, new_E9762_, new_E9763_, new_E9764_, new_E9765_,
    new_E9766_, new_E9767_, new_E9768_, new_E9769_, new_E9770_, new_E9771_,
    new_E9772_, new_E9773_, new_E9774_, new_E9775_, new_E9776_, new_E9777_,
    new_E9778_, new_E9779_, new_E9780_, new_E9781_, new_E9782_, new_E9783_,
    new_E9784_, new_E9785_, new_E9786_, new_E9787_, new_E9788_, new_E9789_,
    new_E9790_, new_E9791_, new_E9792_, new_E9793_, new_E9794_, new_E9795_,
    new_E9796_, new_E9797_, new_E9798_, new_E9799_, new_E9800_, new_E9801_,
    new_E9802_, new_E9803_, new_E9804_, new_E9805_, new_E9806_, new_E9807_,
    new_E9808_, new_E9809_, new_E9810_, new_E9811_, new_E9812_, new_E9813_,
    new_E9814_, new_E9815_, new_E9816_, new_E9817_, new_E9818_, new_E9819_,
    new_E9820_, new_E9821_, new_E9822_, new_E9823_, new_E9824_, new_E9825_,
    new_E9826_, new_E9827_, new_E9828_, new_E9829_, new_E9830_, new_E9831_,
    new_E9832_, new_E9833_, new_E9834_, new_E9835_, new_E9836_, new_E9837_,
    new_E9838_, new_E9839_, new_E9840_, new_E9841_, new_E9842_, new_E9843_,
    new_E9844_, new_E9845_, new_E9846_, new_E9847_, new_E9848_, new_E9849_,
    new_E9850_, new_E9851_, new_E9852_, new_E9853_, new_E9854_, new_E9855_,
    new_E9856_, new_E9857_, new_E9858_, new_E9859_, new_E9860_, new_E9861_,
    new_E9862_, new_E9863_, new_E9864_, new_E9865_, new_E9866_, new_E9867_,
    new_E9868_, new_E9869_, new_E9870_, new_E9871_, new_E9872_, new_E9873_,
    new_E9874_, new_E9875_, new_E9876_, new_E9877_, new_E9878_, new_E9879_,
    new_E9880_, new_E9881_, new_E9882_, new_E9883_, new_E9884_, new_E9885_,
    new_E9886_, new_E9887_, new_E9888_, new_E9889_, new_E9890_, new_E9891_,
    new_E9892_, new_E9893_, new_E9894_, new_E9895_, new_E9896_, new_E9897_,
    new_E9898_, new_E9899_, new_E9900_, new_E9901_, new_E9902_, new_E9903_,
    new_E9904_, new_E9905_, new_E9906_, new_E9907_, new_E9908_, new_E9909_,
    new_E9910_, new_E9911_, new_E9912_, new_E9913_, new_E9914_, new_E9915_,
    new_E9916_, new_E9917_, new_E9918_, new_E9919_, new_E9920_, new_E9921_,
    new_E9922_, new_E9923_, new_E9924_, new_E9925_, new_E9926_, new_E9927_,
    new_E9928_, new_E9929_, new_E9930_, new_E9931_, new_E9932_, new_E9933_,
    new_E9934_, new_E9935_, new_E9936_, new_E9937_, new_E9938_, new_E9939_,
    new_E9940_, new_E9941_, new_E9942_, new_E9943_, new_E9944_, new_E9945_,
    new_E9946_, new_E9947_, new_E9948_, new_E9949_, new_E9950_, new_E9951_,
    new_E9952_, new_E9953_, new_E9954_, new_E9955_, new_E9956_, new_E9957_,
    new_E9958_, new_E9959_, new_E9960_, new_E9961_, new_E9962_, new_E9963_,
    new_E9964_, new_E9965_, new_E9966_, new_E9967_, new_E9968_, new_E9969_,
    new_E9970_, new_E9971_, new_E9972_, new_E9973_, new_E9974_, new_E9975_,
    new_E9976_, new_E9977_, new_E9978_, new_E9979_, new_E9980_, new_E9981_,
    new_E9982_, new_E9983_, new_E9984_, new_E9985_, new_E9986_, new_E9987_,
    new_E9988_, new_E9989_, new_E9990_, new_E9991_, new_E9992_, new_E9993_,
    new_E9994_, new_E9995_, new_E9996_, new_E9997_, new_E9998_, new_E9999_,
    new_F1_, new_F2_, new_F3_, new_F4_, new_F5_, new_F6_, new_F7_, new_F8_,
    new_F9_, new_F10_, new_F11_, new_F12_, new_F13_, new_F14_, new_F15_,
    new_F16_, new_F17_, new_F18_, new_F19_, new_F20_, new_F21_, new_F22_,
    new_F23_, new_F24_, new_F25_, new_F26_, new_F27_, new_F28_, new_F29_,
    new_F30_, new_F31_, new_F32_, new_F33_, new_F34_, new_F35_, new_F36_,
    new_F37_, new_F38_, new_F39_, new_F40_, new_F41_, new_F42_, new_F43_,
    new_F44_, new_F45_, new_F46_, new_F47_, new_F48_, new_F49_, new_F50_,
    new_F51_, new_F52_, new_F53_, new_F54_, new_F55_, new_F56_, new_F57_,
    new_F58_, new_F59_, new_F60_, new_F61_, new_F62_, new_F63_, new_F64_,
    new_F65_, new_F66_, new_F67_, new_F68_, new_F69_, new_F70_, new_F71_,
    new_F72_, new_F73_, new_F74_, new_F75_, new_F76_, new_F77_, new_F78_,
    new_F79_, new_F80_, new_F81_, new_F82_, new_F83_, new_F84_, new_F85_,
    new_F86_, new_F87_, new_F88_, new_F89_, new_F90_, new_F91_, new_F92_,
    new_F93_, new_F94_, new_F95_, new_F96_, new_F97_, new_F98_, new_F99_,
    new_F100_, new_F101_, new_F102_, new_F103_, new_F104_, new_F105_,
    new_F106_, new_F107_, new_F108_, new_F109_, new_F110_, new_F111_,
    new_F112_, new_F113_, new_F114_, new_F115_, new_F116_, new_F117_,
    new_F118_, new_F119_, new_F120_, new_F121_, new_F122_, new_F123_,
    new_F124_, new_F125_, new_F126_, new_F127_, new_F128_, new_F129_,
    new_F130_, new_F131_, new_F132_, new_F133_, new_F134_, new_F135_,
    new_F136_, new_F137_, new_F138_, new_F139_, new_F140_, new_F141_,
    new_F142_, new_F143_, new_F144_, new_F145_, new_F146_, new_F147_,
    new_F148_, new_F149_, new_F150_, new_F151_, new_F152_, new_F153_,
    new_F154_, new_F155_, new_F156_, new_F157_, new_F158_, new_F159_,
    new_F160_, new_F161_, new_F162_, new_F163_, new_F164_, new_F165_,
    new_F166_, new_F167_, new_F168_, new_F169_, new_F170_, new_F171_,
    new_F172_, new_F173_, new_F174_, new_F175_, new_F176_, new_F177_,
    new_F178_, new_F179_, new_F180_, new_F181_, new_F182_, new_F183_,
    new_F184_, new_F185_, new_F186_, new_F187_, new_F188_, new_F189_,
    new_F190_, new_F191_, new_F192_, new_F193_, new_F194_, new_F195_,
    new_F196_, new_F197_, new_F198_, new_F199_, new_F200_, new_F201_,
    new_F202_, new_F203_, new_F204_, new_F205_, new_F206_, new_F207_,
    new_F208_, new_F209_, new_F210_, new_F211_, new_F212_, new_F213_,
    new_F214_, new_F215_, new_F216_, new_F217_, new_F218_, new_F219_,
    new_F220_, new_F221_, new_F222_, new_F223_, new_F224_, new_F225_,
    new_F226_, new_F227_, new_F228_, new_F229_, new_F230_, new_F231_,
    new_F232_, new_F233_, new_F234_, new_F235_, new_F236_, new_F237_,
    new_F238_, new_F239_, new_F240_, new_F241_, new_F242_, new_F243_,
    new_F244_, new_F245_, new_F246_, new_F247_, new_F248_, new_F249_,
    new_F250_, new_F251_, new_F252_, new_F253_, new_F254_, new_F255_,
    new_F256_, new_F257_, new_F258_, new_F259_, new_F260_, new_F261_,
    new_F262_, new_F263_, new_F264_, new_F265_, new_F266_, new_F267_,
    new_F268_, new_F269_, new_F270_, new_F271_, new_F272_, new_F273_,
    new_F274_, new_F275_, new_F276_, new_F277_, new_F278_, new_F279_,
    new_F280_, new_F281_, new_F282_, new_F283_, new_F284_, new_F285_,
    new_F286_, new_F287_, new_F288_, new_F289_, new_F290_, new_F291_,
    new_F292_, new_F293_, new_F294_, new_F295_, new_F296_, new_F297_,
    new_F298_, new_F299_, new_F300_, new_F301_, new_F302_, new_F303_,
    new_F304_, new_F305_, new_F306_, new_F307_, new_F308_, new_F309_,
    new_F310_, new_F311_, new_F312_, new_F313_, new_F314_, new_F315_,
    new_F316_, new_F317_, new_F318_, new_F319_, new_F320_, new_F321_,
    new_F322_, new_F323_, new_F324_, new_F325_, new_F326_, new_F327_,
    new_F328_, new_F329_, new_F330_, new_F331_, new_F332_, new_F333_,
    new_F334_, new_F335_, new_F336_, new_F337_, new_F338_, new_F339_,
    new_F340_, new_F341_, new_F342_, new_F343_, new_F344_, new_F345_,
    new_F346_, new_F347_, new_F348_, new_F349_, new_F350_, new_F351_,
    new_F352_, new_F353_, new_F354_, new_F355_, new_F356_, new_F357_,
    new_F358_, new_F359_, new_F360_, new_F361_, new_F362_, new_F363_,
    new_F364_, new_F365_, new_F366_, new_F367_, new_F368_, new_F369_,
    new_F370_, new_F371_, new_F372_, new_F373_, new_F374_, new_F375_,
    new_F376_, new_F377_, new_F378_, new_F379_, new_F380_, new_F381_,
    new_F382_, new_F383_, new_F384_, new_F385_, new_F386_, new_F387_,
    new_F388_, new_F389_, new_F390_, new_F391_, new_F392_, new_F393_,
    new_F394_, new_F395_, new_F396_, new_F397_, new_F398_, new_F399_,
    new_F400_, new_F401_, new_F402_, new_F403_, new_F404_, new_F405_,
    new_F406_, new_F407_, new_F408_, new_F409_, new_F410_, new_F411_,
    new_F412_, new_F413_, new_F414_, new_F415_, new_F416_, new_F417_,
    new_F418_, new_F419_, new_F420_, new_F421_, new_F422_, new_F423_,
    new_F424_, new_F425_, new_F426_, new_F427_, new_F428_, new_F429_,
    new_F430_, new_F431_, new_F432_, new_F433_, new_F434_, new_F435_,
    new_F436_, new_F437_, new_F438_, new_F439_, new_F440_, new_F441_,
    new_F442_, new_F443_, new_F444_, new_F445_, new_F446_, new_F447_,
    new_F448_, new_F449_, new_F450_, new_F451_, new_F452_, new_F453_,
    new_F454_, new_F455_, new_F456_, new_F457_, new_F458_, new_F459_,
    new_F460_, new_F461_, new_F462_, new_F463_, new_F464_, new_F465_,
    new_F466_, new_F467_, new_F468_, new_F469_, new_F470_, new_F471_,
    new_F472_, new_F473_, new_F474_, new_F475_, new_F476_, new_F477_,
    new_F478_, new_F479_, new_F480_, new_F481_, new_F482_, new_F483_,
    new_F484_, new_F485_, new_F486_, new_F487_, new_F488_, new_F489_,
    new_F490_, new_F491_, new_F492_, new_F493_, new_F494_, new_F495_,
    new_F496_, new_F497_, new_F498_, new_F499_, new_F500_, new_F501_,
    new_F502_, new_F503_, new_F504_, new_F505_, new_F506_, new_F507_,
    new_F508_, new_F509_, new_F510_, new_F511_, new_F512_, new_F513_,
    new_F514_, new_F515_, new_F516_, new_F517_, new_F518_, new_F519_,
    new_F520_, new_F521_, new_F522_, new_F523_, new_F524_, new_F525_,
    new_F526_, new_F527_, new_F528_, new_F529_, new_F530_, new_F531_,
    new_F532_, new_F533_, new_F534_, new_F535_, new_F536_, new_F537_,
    new_F538_, new_F539_, new_F540_, new_F541_, new_F542_, new_F543_,
    new_F544_, new_F545_, new_F546_, new_F547_, new_F548_, new_F549_,
    new_F550_, new_F551_, new_F552_, new_F553_, new_F554_, new_F555_,
    new_F556_, new_F557_, new_F558_, new_F559_, new_F560_, new_F561_,
    new_F562_, new_F563_, new_F564_, new_F565_, new_F566_, new_F567_,
    new_F568_, new_F569_, new_F570_, new_F571_, new_F572_, new_F573_,
    new_F574_, new_F575_, new_F576_, new_F577_, new_F578_, new_F579_,
    new_F580_, new_F581_, new_F582_, new_F583_, new_F584_, new_F585_,
    new_F586_, new_F587_, new_F588_, new_F589_, new_F590_, new_F591_,
    new_F592_, new_F593_, new_F594_, new_F595_, new_F596_, new_F597_,
    new_F598_, new_F599_, new_F600_, new_F601_, new_F602_, new_F603_,
    new_F604_, new_F605_, new_F606_, new_F607_, new_F608_, new_F609_,
    new_F610_, new_F611_, new_F612_, new_F613_, new_F614_, new_F615_,
    new_F616_, new_F617_, new_F618_, new_F619_, new_F620_, new_F621_,
    new_F622_, new_F623_, new_F624_, new_F625_, new_F626_, new_F627_,
    new_F628_, new_F629_, new_F630_, new_F631_, new_F632_, new_F633_,
    new_F634_, new_F635_, new_F636_, new_F637_, new_F638_, new_F639_,
    new_F640_, new_F641_, new_F642_, new_F643_, new_F644_, new_F645_,
    new_F646_, new_F647_, new_F648_, new_F649_, new_F650_, new_F651_,
    new_F652_, new_F653_, new_F654_, new_F655_, new_F656_, new_F657_,
    new_F658_, new_F659_, new_F660_, new_F661_, new_F662_, new_F663_,
    new_F664_, new_F665_, new_F666_, new_F667_, new_F668_, new_F669_,
    new_F670_, new_F671_, new_F672_, new_F673_, new_F674_, new_F675_,
    new_F676_, new_F677_, new_F678_, new_F679_, new_F680_, new_F681_,
    new_F682_, new_F683_, new_F684_, new_F685_, new_F686_, new_F687_,
    new_F688_, new_F689_, new_F690_, new_F691_, new_F692_, new_F693_,
    new_F694_, new_F695_, new_F696_, new_F697_, new_F698_, new_F699_,
    new_F700_, new_F701_, new_F702_, new_F703_, new_F704_, new_F705_,
    new_F706_, new_F707_, new_F708_, new_F709_, new_F710_, new_F711_,
    new_F712_, new_F713_, new_F714_, new_F715_, new_F716_, new_F717_,
    new_F718_, new_F719_, new_F720_, new_F721_, new_F722_, new_F723_,
    new_F724_, new_F725_, new_F726_, new_F727_, new_F728_, new_F729_,
    new_F730_, new_F731_, new_F732_, new_F733_, new_F734_, new_F735_,
    new_F736_, new_F737_, new_F738_, new_F739_, new_F740_, new_F741_,
    new_F742_, new_F743_, new_F744_, new_F745_, new_F746_, new_F747_,
    new_F748_, new_F749_, new_F750_, new_F751_, new_F752_, new_F753_,
    new_F754_, new_F755_, new_F756_, new_F757_, new_F758_, new_F759_,
    new_F760_, new_F761_, new_F762_, new_F763_, new_F764_, new_F765_,
    new_F766_, new_F767_, new_F768_, new_F769_, new_F770_, new_F771_,
    new_F772_, new_F773_, new_F774_, new_F775_, new_F776_, new_F777_,
    new_F778_, new_F779_, new_F780_, new_F781_, new_F782_, new_F783_,
    new_F784_, new_F785_, new_F786_, new_F787_, new_F788_, new_F789_,
    new_F790_, new_F791_, new_F792_, new_F793_, new_F794_, new_F795_,
    new_F796_, new_F797_, new_F798_, new_F799_, new_F800_, new_F801_,
    new_F802_, new_F803_, new_F804_, new_F805_, new_F806_, new_F807_,
    new_F808_, new_F809_, new_F810_, new_F811_, new_F812_, new_F813_,
    new_F814_, new_F815_, new_F816_, new_F817_, new_F818_, new_F819_,
    new_F820_, new_F821_, new_F822_, new_F823_, new_F824_, new_F825_,
    new_F826_, new_F827_, new_F828_, new_F829_, new_F830_, new_F831_,
    new_F832_, new_F833_, new_F834_, new_F835_, new_F836_, new_F837_,
    new_F838_, new_F839_, new_F840_, new_F841_, new_F842_, new_F843_,
    new_F844_, new_F845_, new_F846_, new_F847_, new_F848_, new_F849_,
    new_F850_, new_F851_, new_F852_, new_F853_, new_F854_, new_F855_,
    new_F856_, new_F857_, new_F858_, new_F859_, new_F860_, new_F861_,
    new_F862_, new_F863_, new_F864_, new_F865_, new_F866_, new_F867_,
    new_F868_, new_F869_, new_F870_, new_F871_, new_F872_, new_F873_,
    new_F874_, new_F875_, new_F876_, new_F877_, new_F878_, new_F879_,
    new_F880_, new_F881_, new_F882_, new_F883_, new_F884_, new_F885_,
    new_F886_, new_F887_, new_F888_, new_F889_, new_F890_, new_F891_,
    new_F892_, new_F893_, new_F894_, new_F895_, new_F896_, new_F897_,
    new_F898_, new_F899_, new_F900_, new_F901_, new_F902_, new_F903_,
    new_F904_, new_F905_, new_F906_, new_F907_, new_F908_, new_F909_,
    new_F910_, new_F911_, new_F912_, new_F913_, new_F914_, new_F915_,
    new_F916_, new_F917_, new_F918_, new_F919_, new_F920_, new_F921_,
    new_F922_, new_F923_, new_F924_, new_F925_, new_F926_, new_F927_,
    new_F928_, new_F929_, new_F930_, new_F931_, new_F932_, new_F933_,
    new_F934_, new_F935_, new_F936_, new_F937_, new_F938_, new_F939_,
    new_F940_, new_F941_, new_F942_, new_F943_, new_F944_, new_F945_,
    new_F946_, new_F947_, new_F948_, new_F949_, new_F950_, new_F951_,
    new_F952_, new_F953_, new_F954_, new_F955_, new_F956_, new_F957_,
    new_F958_, new_F959_, new_F960_, new_F961_, new_F962_, new_F963_,
    new_F964_, new_F965_, new_F966_, new_F967_, new_F968_, new_F969_,
    new_F970_, new_F971_, new_F972_, new_F973_, new_F974_, new_F975_,
    new_F976_, new_F977_, new_F978_, new_F979_, new_F980_, new_F981_,
    new_F982_, new_F983_, new_F984_, new_F985_, new_F986_, new_F987_,
    new_F988_, new_F989_, new_F990_, new_F991_, new_F992_, new_F993_,
    new_F994_, new_F995_, new_F996_, new_F997_, new_F998_, new_F999_,
    new_F1000_, new_F1001_, new_F1002_, new_F1003_, new_F1004_, new_F1005_,
    new_F1006_, new_F1007_, new_F1008_, new_F1009_, new_F1010_, new_F1011_,
    new_F1012_, new_F1013_, new_F1014_, new_F1015_, new_F1016_, new_F1017_,
    new_F1018_, new_F1019_, new_F1020_, new_F1021_, new_F1022_, new_F1023_,
    new_F1024_, new_F1025_, new_F1026_, new_F1027_, new_F1028_, new_F1029_,
    new_F1030_, new_F1031_, new_F1032_, new_F1033_, new_F1034_, new_F1035_,
    new_F1036_, new_F1037_, new_F1038_, new_F1039_, new_F1040_, new_F1041_,
    new_F1042_, new_F1043_, new_F1044_, new_F1045_, new_F1046_, new_F1047_,
    new_F1048_, new_F1049_, new_F1050_, new_F1051_, new_F1052_, new_F1053_,
    new_F1054_, new_F1055_, new_F1056_, new_F1057_, new_F1058_, new_F1059_,
    new_F1060_, new_F1061_, new_F1062_, new_F1063_, new_F1064_, new_F1065_,
    new_F1066_, new_F1067_, new_F1068_, new_F1069_, new_F1070_, new_F1071_,
    new_F1072_, new_F1073_, new_F1074_, new_F1075_, new_F1076_, new_F1077_,
    new_F1078_, new_F1079_, new_F1080_, new_F1081_, new_F1082_, new_F1083_,
    new_F1084_, new_F1085_, new_F1086_, new_F1087_, new_F1088_, new_F1089_,
    new_F1090_, new_F1091_, new_F1092_, new_F1093_, new_F1094_, new_F1095_,
    new_F1096_, new_F1097_, new_F1098_, new_F1099_, new_F1100_, new_F1101_,
    new_F1102_, new_F1103_, new_F1104_, new_F1105_, new_F1106_, new_F1107_,
    new_F1108_, new_F1109_, new_F1110_, new_F1111_, new_F1112_, new_F1113_,
    new_F1114_, new_F1115_, new_F1116_, new_F1117_, new_F1118_, new_F1119_,
    new_F1120_, new_F1121_, new_F1122_, new_F1123_, new_F1124_, new_F1125_,
    new_F1126_, new_F1127_, new_F1128_, new_F1129_, new_F1130_, new_F1131_,
    new_F1132_, new_F1133_, new_F1134_, new_F1135_, new_F1136_, new_F1137_,
    new_F1138_, new_F1139_, new_F1140_, new_F1141_, new_F1142_, new_F1143_,
    new_F1144_, new_F1145_, new_F1146_, new_F1147_, new_F1148_, new_F1149_,
    new_F1150_, new_F1151_, new_F1152_, new_F1153_, new_F1154_, new_F1155_,
    new_F1156_, new_F1157_, new_F1158_, new_F1159_, new_F1160_, new_F1161_,
    new_F1162_, new_F1163_, new_F1164_, new_F1165_, new_F1166_, new_F1167_,
    new_F1168_, new_F1169_, new_F1170_, new_F1171_, new_F1172_, new_F1173_,
    new_F1174_, new_F1175_, new_F1176_, new_F1177_, new_F1178_, new_F1179_,
    new_F1180_, new_F1181_, new_F1182_, new_F1183_, new_F1184_, new_F1185_,
    new_F1186_, new_F1187_, new_F1188_, new_F1189_, new_F1190_, new_F1191_,
    new_F1192_, new_F1193_, new_F1194_, new_F1195_, new_F1196_, new_F1197_,
    new_F1198_, new_F1199_, new_F1200_, new_F1201_, new_F1202_, new_F1203_,
    new_F1204_, new_F1205_, new_F1206_, new_F1207_, new_F1208_, new_F1209_,
    new_F1210_, new_F1211_, new_F1212_, new_F1213_, new_F1214_, new_F1215_,
    new_F1216_, new_F1217_, new_F1218_, new_F1219_, new_F1220_, new_F1221_,
    new_F1222_, new_F1223_, new_F1224_, new_F1225_, new_F1226_, new_F1227_,
    new_F1228_, new_F1229_, new_F1230_, new_F1231_, new_F1232_, new_F1233_,
    new_F1234_, new_F1235_, new_F1236_, new_F1237_, new_F1238_, new_F1239_,
    new_F1240_, new_F1241_, new_F1242_, new_F1243_, new_F1244_, new_F1245_,
    new_F1246_, new_F1247_, new_F1248_, new_F1249_, new_F1250_, new_F1251_,
    new_F1252_, new_F1253_, new_F1254_, new_F1255_, new_F1256_, new_F1257_,
    new_F1258_, new_F1259_, new_F1260_, new_F1261_, new_F1262_, new_F1263_,
    new_F1264_, new_F1265_, new_F1266_, new_F1267_, new_F1268_, new_F1269_,
    new_F1270_, new_F1271_, new_F1272_, new_F1273_, new_F1274_, new_F1275_,
    new_F1276_, new_F1277_, new_F1278_, new_F1279_, new_F1280_, new_F1281_,
    new_F1282_, new_F1283_, new_F1284_, new_F1285_, new_F1286_, new_F1287_,
    new_F1288_, new_F1289_, new_F1290_, new_F1291_, new_F1292_, new_F1293_,
    new_F1294_, new_F1295_, new_F1296_, new_F1297_, new_F1298_, new_F1299_,
    new_F1300_, new_F1301_, new_F1302_, new_F1303_, new_F1304_, new_F1305_,
    new_F1306_, new_F1307_, new_F1308_, new_F1309_, new_F1310_, new_F1311_,
    new_F1312_, new_F1313_, new_F1314_, new_F1315_, new_F1316_, new_F1317_,
    new_F1318_, new_F1319_, new_F1320_, new_F1321_, new_F1322_, new_F1323_,
    new_F1324_, new_F1325_, new_F1326_, new_F1327_, new_F1328_, new_F1329_,
    new_F1330_, new_F1331_, new_F1332_, new_F1333_, new_F1334_, new_F1335_,
    new_F1336_, new_F1337_, new_F1338_, new_F1339_, new_F1340_, new_F1341_,
    new_F1342_, new_F1343_, new_F1344_, new_F1345_, new_F1346_, new_F1347_,
    new_F1348_, new_F1349_, new_F1350_, new_F1351_, new_F1352_, new_F1353_,
    new_F1354_, new_F1355_, new_F1356_, new_F1357_, new_F1358_, new_F1359_,
    new_F1360_, new_F1361_, new_F1362_, new_F1363_, new_F1364_, new_F1365_,
    new_F1366_, new_F1367_, new_F1368_, new_F1369_, new_F1370_, new_F1371_,
    new_F1372_, new_F1373_, new_F1374_, new_F1375_, new_F1376_, new_F1377_,
    new_F1378_, new_F1379_, new_F1380_, new_F1381_, new_F1382_, new_F1383_,
    new_F1384_, new_F1385_, new_F1386_, new_F1387_, new_F1388_, new_F1389_,
    new_F1390_, new_F1391_, new_F1392_, new_F1393_, new_F1394_, new_F1395_,
    new_F1396_, new_F1397_, new_F1398_, new_F1399_, new_F1400_, new_F1401_,
    new_F1402_, new_F1403_, new_F1404_, new_F1405_, new_F1406_, new_F1407_,
    new_F1408_, new_F1409_, new_F1410_, new_F1411_, new_F1412_, new_F1413_,
    new_F1414_, new_F1415_, new_F1416_, new_F1417_, new_F1418_, new_F1419_,
    new_F1420_, new_F1421_, new_F1422_, new_F1423_, new_F1424_, new_F1425_,
    new_F1426_, new_F1427_, new_F1428_, new_F1429_, new_F1430_, new_F1431_,
    new_F1432_, new_F1433_, new_F1434_, new_F1435_, new_F1436_, new_F1437_,
    new_F1438_, new_F1439_, new_F1440_, new_F1441_, new_F1442_, new_F1443_,
    new_F1444_, new_F1445_, new_F1446_, new_F1447_, new_F1448_, new_F1449_,
    new_F1450_, new_F1451_, new_F1452_, new_F1453_, new_F1454_, new_F1455_,
    new_F1456_, new_F1457_, new_F1458_, new_F1459_, new_F1460_, new_F1461_,
    new_C2581_, new_C2580_, new_C2579_, new_C2578_, new_C2577_, new_C2576_,
    new_C2575_, new_C2574_, new_C2573_, new_C2572_, new_C2571_, new_C2570_,
    new_C2569_, new_C2568_, new_C2567_, new_C2566_, new_C2565_, new_C2564_,
    new_C2563_, new_C2562_, new_C2561_, new_C2560_, new_C2559_, new_C2558_,
    new_C2557_, new_C2556_, new_C2555_, new_C2554_, new_C2553_, new_C2552_,
    new_C2551_, new_C2550_, new_C2549_, new_C2548_, new_C2547_, new_C2546_,
    new_C2545_, new_C2544_, new_C2543_, new_C2542_, new_C2541_, new_C2540_,
    new_C2539_, new_C2538_, new_C2537_, new_C2536_, new_C2535_, new_C2534_,
    new_C2533_, new_C2532_, new_C2531_, new_C2530_, new_C2529_, new_C2528_,
    new_C2527_, new_C2526_, new_C2525_, new_C2524_, new_C2523_, new_C2522_,
    new_C2521_, new_C2520_, new_C2519_, new_C2518_, new_C2517_, new_C2516_,
    new_C2515_, new_C2582_, new_C2583_, new_C2584_, new_C2585_, new_C2586_,
    new_C2587_, new_C2588_, new_C2589_, new_C2590_, new_C2591_, new_C2592_,
    new_C2593_, new_C2594_, new_C2595_, new_C2596_, new_C2597_, new_C2598_,
    new_C2599_, new_C2600_, new_C2601_, new_C2602_, new_C2603_, new_C2604_,
    new_C2605_, new_C2606_, new_C2607_, new_C2608_, new_C2609_, new_C2610_,
    new_C2611_, new_C2612_, new_C2613_, new_C2614_, new_C2615_, new_C2616_,
    new_C2617_, new_C2618_, new_C2619_, new_C2620_, new_C2621_, new_C2622_,
    new_C2623_, new_C2624_, new_C2625_, new_C2626_, new_C2627_, new_C2628_,
    new_C2629_, new_C2630_, new_C2631_, new_C2632_, new_C2633_, new_C2634_,
    new_C2635_, new_C2636_, new_C2637_, new_C2638_, new_C2639_, new_C2640_,
    new_C2641_, new_C2642_, new_C2643_, new_C2644_, new_C2645_, new_C2646_,
    new_C2647_, new_C2648_, new_C2649_, new_C2650_, new_C2651_, new_C2652_,
    new_C2653_, new_C2654_, new_C2655_, new_C2656_, new_C2657_, new_C2658_,
    new_C2659_, new_C2660_, new_C2661_, new_C2662_, new_C2663_, new_C2664_,
    new_C2665_, new_C2666_, new_C2667_, new_C2668_, new_C2669_, new_C2670_,
    new_C2671_, new_C2672_, new_C2673_, new_C2674_, new_C2675_, new_C2676_,
    new_C2677_, new_C2678_, new_C2679_, new_C2680_, new_C2681_, new_C2682_,
    new_C2683_, new_C2684_, new_C2685_, new_C2686_, new_C2687_, new_C2688_,
    new_C2689_, new_C2690_, new_C2691_, new_C2692_, new_C2693_, new_C2694_,
    new_C2695_, new_C2696_, new_C2697_, new_C2698_, new_C2699_, new_C2700_,
    new_C2701_, new_C2702_, new_C2703_, new_C2704_, new_C2705_, new_C2706_,
    new_C2707_, new_C2708_, new_C2709_, new_C2710_, new_C2711_, new_C2712_,
    new_C2713_, new_C2714_, new_C2715_, new_C2716_, new_C2717_, new_C2718_,
    new_C2719_, new_C2720_, new_C2721_, new_C2722_, new_C2723_, new_C2724_,
    new_C2725_, new_C2726_, new_C2727_, new_C2728_, new_C2729_, new_C2730_,
    new_C2731_, new_C2732_, new_C2733_, new_C2734_, new_C2735_, new_C2736_,
    new_C2737_, new_C2738_, new_C2739_, new_C2740_, new_C2741_, new_C2742_,
    new_C2743_, new_C2744_, new_C2745_, new_C2746_, new_C2747_, new_C2748_,
    new_C2749_, new_C2750_, new_C2751_, new_C2752_, new_C2753_, new_C2754_,
    new_C2755_, new_C2756_, new_C2757_, new_C2758_, new_C2759_, new_C2760_,
    new_C2761_, new_C2762_, new_C2763_, new_C2764_, new_C2765_, new_C2766_,
    new_C2767_, new_C2768_, new_C2769_, new_C2770_, new_C2771_, new_C2772_,
    new_C2773_, new_C2774_, new_C2775_, new_C2776_, new_C2777_, new_C2778_,
    new_C2779_, new_C2780_, new_C2781_, new_C2782_, new_C2783_, new_C2784_,
    new_C2785_, new_C2786_, new_C2787_, new_C2788_, new_C2789_, new_C2790_,
    new_C2791_, new_C2792_, new_C2793_, new_C2794_, new_C2795_, new_C2796_,
    new_C2797_, new_C2798_, new_C2799_, new_C2800_, new_C2801_, new_C2802_,
    new_C2803_, new_C2804_, new_C2805_, new_C2806_, new_C2807_, new_C2808_,
    new_C2809_, new_C2810_, new_C2811_, new_C2812_, new_C2813_, new_C2814_,
    new_C2815_, new_C2816_, new_C2817_, new_C2818_, new_C2819_, new_C2820_,
    new_C2821_, new_C2822_, new_C2823_, new_C2824_, new_C2825_, new_C2826_,
    new_C2827_, new_C2828_, new_C2829_, new_C2830_, new_C2831_, new_C2832_,
    new_C2833_, new_C2834_, new_C2835_, new_C2836_, new_C2837_, new_C2838_,
    new_C2839_, new_C2840_, new_C2841_, new_C2842_, new_C2843_, new_C2844_,
    new_C2845_, new_C2846_, new_C2847_, new_C2848_, new_C2849_, new_C2850_,
    new_C2851_, new_C2852_, new_C2853_, new_C2854_, new_C2855_, new_C2856_,
    new_C2857_, new_C2858_, new_C2859_, new_C2860_, new_C2861_, new_C2862_,
    new_C2863_, new_C2864_, new_C2865_, new_C2866_, new_C2867_, new_C2868_,
    new_C2869_, new_C2870_, new_C2871_, new_C2872_, new_C2873_, new_C2874_,
    new_C2875_, new_C2876_, new_C2877_, new_C2878_, new_C2879_, new_C2880_,
    new_C2881_, new_C2882_, new_C2883_, new_C2884_, new_C2885_, new_C2886_,
    new_C2887_, new_C2888_, new_C2889_, new_C2890_, new_C2891_, new_C2892_,
    new_C2893_, new_C2894_, new_C2895_, new_C2896_, new_C2897_, new_C2898_,
    new_C2899_, new_C2900_, new_C2901_, new_C2902_, new_C2903_, new_C2904_,
    new_C2905_, new_C2906_, new_C2907_, new_C2908_, new_C2909_, new_C2910_,
    new_C2911_, new_C2912_, new_C2913_, new_C2914_, new_C2915_, new_C2916_,
    new_C2917_, new_C2918_, new_C2919_, new_C2920_, new_C2921_, new_C2922_,
    new_C2923_, new_C2924_, new_C2925_, new_C2926_, new_C2927_, new_C2928_,
    new_C2929_, new_C2930_, new_C2931_, new_C2932_, new_C2933_, new_C2934_,
    new_C2935_, new_C2936_, new_C2937_, new_C2938_, new_C2939_, new_C2940_,
    new_C2941_, new_C2942_, new_C2943_, new_C2944_, new_C2945_, new_C2946_,
    new_C2947_, new_C2948_, new_C2949_, new_C2950_, new_C2951_, new_C2952_,
    new_C2953_, new_C2954_, new_C2955_, new_C2956_, new_C2957_, new_C2958_,
    new_C2959_, new_C2960_, new_C2961_, new_C2962_, new_C2963_, new_C2964_,
    new_C2965_, new_C2966_, new_C2967_, new_C2968_, new_C2969_, new_C2970_,
    new_C2971_, new_C2972_, new_C2973_, new_C2974_, new_C2975_, new_C2976_,
    new_C2977_, new_C2978_, new_C2979_, new_C2980_, new_C2981_, new_C2982_,
    new_C2983_, new_C2984_, new_C2985_, new_C2986_, new_C2987_, new_C2988_,
    new_C2989_, new_C2990_, new_C2991_, new_C2992_, new_C2993_, new_C2994_,
    new_C2995_, new_C2996_, new_C2997_, new_C2998_, new_C2999_, new_C3000_,
    new_C3001_, new_C3002_, new_C3003_, new_C3004_, new_C3005_, new_C3006_,
    new_C3007_, new_C3008_, new_C3009_, new_C3010_, new_C3011_, new_C3012_,
    new_C3013_, new_C3014_, new_C3015_, new_C3016_, new_C3017_, new_C3018_,
    new_C3019_, new_C3020_, new_C3021_, new_C3022_, new_C3023_, new_C3024_,
    new_C3025_, new_C3026_, new_C3027_, new_C3028_, new_C3029_, new_C3030_,
    new_C3031_, new_C3032_, new_C3033_, new_C3034_, new_C3035_, new_C3036_,
    new_C3037_, new_C3038_, new_C3039_, new_C3040_, new_C3041_, new_C3042_,
    new_C3043_, new_C3044_, new_C3045_, new_C3046_, new_C3047_, new_C3048_,
    new_C3049_, new_C3050_, new_C3051_, new_C3052_, new_C3053_, new_C3054_,
    new_C3055_, new_C3056_, new_C3057_, new_C3058_, new_C3059_, new_C3060_,
    new_C3061_, new_C3062_, new_C3063_, new_C3064_, new_C3065_, new_C3066_,
    new_C3067_, new_C3068_, new_C3069_, new_C3070_, new_C3071_, new_C3072_,
    new_C3073_, new_C3074_, new_C3075_, new_C3076_, new_C3077_, new_C3078_,
    new_C3079_, new_C3080_, new_C3081_, new_C3082_, new_C3083_, new_C3084_,
    new_C3085_, new_C3086_, new_C3087_, new_C3088_, new_C3089_, new_C3090_,
    new_C3091_, new_C3092_, new_C3093_, new_C3094_, new_C3095_, new_C3096_,
    new_C3097_, new_C3098_, new_C3099_, new_C3100_, new_C3101_, new_C3102_,
    new_C3103_, new_C3104_, new_C3105_, new_C3106_, new_C3107_, new_C3108_,
    new_C3109_, new_C3110_, new_C3111_, new_C3112_, new_C3113_, new_C3114_,
    new_C3115_, new_C3116_, new_C3117_, new_C3118_, new_C3119_, new_C3120_,
    new_C3121_, new_C3122_, new_C3123_, new_C3124_, new_C3125_, new_C3126_,
    new_C3127_, new_C3128_, new_C3129_, new_C3130_, new_C3131_, new_C3132_,
    new_C3133_, new_C3134_, new_C3135_, new_C3136_, new_C3137_, new_C3138_,
    new_C3139_, new_C3140_, new_C3141_, new_C3142_, new_C3143_, new_C3144_,
    new_C3145_, new_C3146_, new_C3147_, new_C3148_, new_C3149_, new_C3150_,
    new_C3151_, new_C3152_, new_C3153_, new_C3154_, new_C3155_, new_C3156_,
    new_C3157_, new_C3158_, new_C3159_, new_C3160_, new_C3161_, new_C3162_,
    new_C3163_, new_C3164_, new_C3165_, new_C3166_, new_C3167_, new_C3168_,
    new_C3169_, new_C3170_, new_C3171_, new_C3172_, new_C3173_, new_C3174_,
    new_C3175_, new_C3176_, new_C3177_, new_C3178_, new_C3179_, new_C3180_,
    new_C3181_, new_C3182_, new_C3183_, new_C3184_, new_C3185_, new_C3186_,
    new_C3187_, new_C3188_, new_C3189_, new_C3190_, new_C3191_, new_C3192_,
    new_C3193_, new_C3194_, new_C3195_, new_C3196_, new_C3197_, new_C3198_,
    new_C3199_, new_C3200_, new_C3201_, new_C3202_, new_C3203_, new_C3204_,
    new_C3205_, new_C3206_, new_C3207_, new_C3208_, new_C3209_, new_C3210_,
    new_C3211_, new_C3212_, new_C3213_, new_C3214_, new_C3215_, new_C3216_,
    new_C3217_, new_C3218_, new_C3219_, new_C3220_, new_C3221_, new_C3222_,
    new_C3223_, new_C3224_, new_C3225_, new_C3226_, new_C3227_, new_C3228_,
    new_C3229_, new_C3230_, new_C3231_, new_C3232_, new_C3233_, new_C3234_,
    new_C3235_, new_C3236_, new_C3237_, new_C3238_, new_C3239_, new_C3240_,
    new_C3241_, new_C3242_, new_C3243_, new_C3244_, new_C3245_, new_C3246_,
    new_C3247_, new_C3248_, new_C3249_, new_C3250_, new_C3251_, new_C3252_,
    new_C3253_, new_C3254_, new_C3255_, new_C3256_, new_C3257_, new_C3258_,
    new_C3259_, new_C3260_, new_C3261_, new_C3262_, new_C3263_, new_C3264_,
    new_C3265_, new_C3266_, new_C3267_, new_C3268_, new_C3269_, new_C3270_,
    new_C3271_, new_C3272_, new_C3273_, new_C3274_, new_C3275_, new_C3276_,
    new_C3277_, new_C3278_, new_C3279_, new_C3280_, new_C3281_, new_C3282_,
    new_C3283_, new_C3284_, new_C3285_, new_C3286_, new_C3287_, new_C3288_,
    new_C3289_, new_C3290_, new_C3291_, new_C3292_, new_C3293_, new_C3294_,
    new_C3295_, new_C3296_, new_C3297_, new_C3298_, new_C3299_, new_C3300_,
    new_C3301_, new_C3302_, new_C3303_, new_C3304_, new_C3305_, new_C3306_,
    new_C3307_, new_C3308_, new_C3309_, new_C3310_, new_C3311_, new_C3312_,
    new_C3313_, new_C3314_, new_C3315_, new_C3316_, new_C3317_, new_C3318_,
    new_C3319_, new_C3320_, new_C3321_, new_C3322_, new_C3323_, new_C3324_,
    new_C3325_, new_C3326_, new_C3327_, new_C3328_, new_C3329_, new_C3330_,
    new_C3331_, new_C3332_, new_C3333_, new_C3334_, new_C3335_, new_C3336_,
    new_C3337_, new_C3338_, new_C3339_, new_C3340_, new_C3341_, new_C3342_,
    new_C3343_, new_C3344_, new_C3345_, new_C3346_, new_C3347_, new_C3348_,
    new_C3349_, new_C3350_, new_C3351_, new_C3352_, new_C3353_, new_C3354_,
    new_C3355_, new_C3356_, new_C3357_, new_C3358_, new_C3359_, new_C3360_,
    new_C3361_, new_C3362_, new_C3363_, new_C3364_, new_C3365_, new_C3366_,
    new_C3367_, new_C3368_, new_C3369_, new_C3370_, new_C3371_, new_C3372_,
    new_C3373_, new_C3374_, new_C3375_, new_C3376_, new_C3377_, new_C3378_,
    new_C3379_, new_C3380_, new_C3381_, new_C3382_, new_C3383_, new_C3384_,
    new_C3385_, new_C3386_, new_C3387_, new_C3388_, new_C3389_, new_C3390_,
    new_C3391_, new_C3392_, new_C3393_, new_C3394_, new_C3395_, new_C3396_,
    new_C3397_, new_C3398_, new_C3399_, new_C3400_, new_C3401_, new_C3402_,
    new_C3403_, new_C3404_, new_C3405_, new_C3406_, new_C3407_, new_C3408_,
    new_C3409_, new_C3410_, new_C3411_, new_C3412_, new_C3413_, new_C3414_,
    new_C3415_, new_C3416_, new_C3417_, new_C3418_, new_C3419_, new_C3420_,
    new_C3421_, new_C3422_, new_C3423_, new_C3424_, new_C3425_, new_C3426_,
    new_C3427_, new_C3428_, new_C3429_, new_C3430_, new_C3431_, new_C3432_,
    new_C3433_, new_C3434_, new_C3435_, new_C3436_, new_C3437_, new_C3438_,
    new_C3439_, new_C3440_, new_C3441_, new_C3442_, new_C3443_, new_C3444_,
    new_C3445_, new_C3446_, new_C3447_, new_C3448_, new_C3449_, new_C3450_,
    new_C3451_, new_C3452_, new_C3453_, new_C3454_, new_C3455_, new_C3456_,
    new_C3457_, new_C3458_, new_C3459_, new_C3460_, new_C3461_, new_C3462_,
    new_C3463_, new_C3464_, new_C3465_, new_C3466_, new_C3467_, new_C3468_,
    new_C3469_, new_C3470_, new_C3471_, new_C3472_, new_C3473_, new_C3474_,
    new_C3475_, new_C3476_, new_C3477_, new_C3478_, new_C3479_, new_C3480_,
    new_C3481_, new_C3482_, new_C3483_, new_C3484_, new_C3485_, new_C3486_,
    new_C3487_, new_C3488_, new_C3489_, new_C3490_, new_C3491_, new_C3492_,
    new_C3493_, new_C3494_, new_C3495_, new_C3496_, new_C3497_, new_C3498_,
    new_C3499_, new_C3500_, new_C3501_, new_C3502_, new_C3503_, new_C3504_,
    new_C3505_, new_C3506_, new_C3507_, new_C3508_, new_C3509_, new_C3510_,
    new_C3511_, new_C3512_, new_C3513_, new_C3514_, new_C3515_, new_C3516_,
    new_C3517_, new_C3518_, new_C3519_, new_C3520_, new_C3521_, new_C3522_,
    new_C3523_, new_C3524_, new_C3525_, new_C3526_, new_C3527_, new_C3528_,
    new_C3529_, new_C3530_, new_C3531_, new_C3532_, new_C3533_, new_C3534_,
    new_C3535_, new_C3536_, new_C3537_, new_C3538_, new_C3539_, new_C3540_,
    new_C3541_, new_C3542_, new_C3543_, new_C3544_, new_C3545_, new_C3546_,
    new_C3547_, new_C3548_, new_C3549_, new_C3550_, new_C3551_, new_C3552_,
    new_C3553_, new_C3554_, new_C3555_, new_C3556_, new_C3557_, new_C3558_,
    new_C3559_, new_C3560_, new_C3561_, new_C3562_, new_C3563_, new_C3564_,
    new_C3565_, new_C3566_, new_C3567_, new_C3568_, new_C3569_, new_C3570_,
    new_C3571_, new_C3572_, new_C3573_, new_C3574_, new_C3575_, new_C3576_,
    new_C3577_, new_C3578_, new_C3579_, new_C3580_, new_C3581_, new_C3582_,
    new_C3583_, new_C3584_, new_C3585_, new_C3586_, new_C3587_, new_C3588_,
    new_C3589_, new_C3590_, new_C3591_, new_C3592_, new_C3593_, new_C3594_,
    new_C3595_, new_C3596_, new_C3597_, new_C3598_, new_C3599_, new_C3600_,
    new_C3601_, new_C3602_, new_C3603_, new_C3604_, new_C3605_, new_C3606_,
    new_C3607_, new_C3608_, new_C3609_, new_C3610_, new_C3611_, new_C3612_,
    new_C3613_, new_C3614_, new_C3615_, new_C3616_, new_C3617_, new_C3618_,
    new_C3619_, new_C3620_, new_C3621_, new_C3622_, new_C3623_, new_C3624_,
    new_C3625_, new_C3626_, new_C3627_, new_C3628_, new_C3629_, new_C3630_,
    new_C3631_, new_C3632_, new_C3633_, new_C3634_, new_C3635_, new_C3636_,
    new_C3637_, new_C3638_, new_C3639_, new_C3640_, new_C3641_, new_C3642_,
    new_C3643_, new_C3644_, new_C3645_, new_C3646_, new_C3647_, new_C3648_,
    new_C3649_, new_C3650_, new_C3651_, new_C3652_, new_C3653_, new_C3654_,
    new_C3655_, new_C3656_, new_C3657_, new_C3658_, new_C3659_, new_C3660_,
    new_C3661_, new_C3662_, new_C3663_, new_C3664_, new_C3665_, new_C3666_,
    new_C3667_, new_C3668_, new_C3669_, new_C3670_, new_C3671_, new_C3672_,
    new_C3673_, new_C3674_, new_C3675_, new_C3676_, new_C3677_, new_C3678_,
    new_C3679_, new_C3680_, new_C3681_, new_C3682_, new_C3683_, new_C3684_,
    new_C3685_, new_C3686_, new_C3687_, new_C3688_, new_C3689_, new_C3690_,
    new_C3691_, new_C3692_, new_C3693_, new_C3694_, new_C3695_, new_C3696_,
    new_C3697_, new_C3698_, new_C3699_, new_C3700_, new_C3701_, new_C3702_,
    new_C3703_, new_C3704_, new_C3705_, new_C3706_, new_C3707_, new_C3708_,
    new_C3709_, new_C3710_, new_C3711_, new_C3712_, new_C3713_, new_C3714_,
    new_C3715_, new_C3716_, new_C3717_, new_C3718_, new_C3719_, new_C3720_,
    new_C3721_, new_C3722_, new_C3723_, new_C3724_, new_C3725_, new_C3726_,
    new_C3727_, new_C3728_, new_C3729_, new_C3730_, new_C3731_, new_C3732_,
    new_C3733_, new_C3734_, new_C3735_, new_C3736_, new_C3737_, new_C3738_,
    new_C3739_, new_C3740_, new_C3741_, new_C3742_, new_C3743_, new_C3744_,
    new_C3745_, new_C3746_, new_C3747_, new_C3748_, new_C3749_, new_C3750_,
    new_C3751_, new_C3752_, new_C3753_, new_C3754_, new_C3755_, new_C3756_,
    new_C3757_, new_C3758_, new_C3759_, new_C3760_, new_C3761_, new_C3762_,
    new_C3763_, new_C3764_, new_C3765_, new_C3766_, new_C3767_, new_C3768_,
    new_C3769_, new_C3770_, new_C3771_, new_C3772_, new_C3773_, new_C3774_,
    new_C3775_, new_C3776_, new_C3777_, new_C3778_, new_C3779_, new_C3780_,
    new_C3781_, new_C3782_, new_C3783_, new_C3784_, new_C3785_, new_C3786_,
    new_C3787_, new_C3788_, new_C3789_, new_C3790_, new_C3791_, new_C3792_,
    new_C3793_, new_C3794_, new_C3795_, new_C3796_, new_C3797_, new_C3798_,
    new_C3799_, new_C3800_, new_C3801_, new_C3802_, new_C3803_, new_C3804_,
    new_C3805_, new_C3806_, new_C3807_, new_C3808_, new_C3809_, new_C3810_,
    new_C3811_, new_C3812_, new_C3813_, new_C3814_, new_C3815_, new_C3816_,
    new_C3817_, new_C3818_, new_C3819_, new_C3820_, new_C3821_, new_C3822_,
    new_C3823_, new_C3824_, new_C3825_, new_C3826_, new_C3827_, new_C3828_,
    new_C3829_, new_C3830_, new_C3831_, new_C3832_, new_C3833_, new_C3834_,
    new_C3835_, new_C3836_, new_C3837_, new_C3838_, new_C3839_, new_C3840_,
    new_C3841_, new_C3842_, new_C3843_, new_C3844_, new_C3845_, new_C3846_,
    new_C3847_, new_C3848_, new_C3849_, new_C3850_, new_C3851_, new_C3852_,
    new_C3853_, new_C3854_, new_C3855_, new_C3856_, new_C3857_, new_C3858_,
    new_C3859_, new_C3860_, new_C3861_, new_C3862_, new_C3863_, new_C3864_,
    new_C3865_, new_C3866_, new_C3867_, new_C3868_, new_C3869_, new_C3870_,
    new_C3871_, new_C3872_, new_C3873_, new_C3874_, new_C3875_, new_C3876_,
    new_C3877_, new_C3878_, new_C3879_, new_C3880_, new_C3881_, new_C3882_,
    new_C3883_, new_C3884_, new_C3885_, new_C3886_, new_C3887_, new_C3888_,
    new_C3889_, new_C3890_, new_C3891_, new_C3892_, new_C3893_, new_C3894_,
    new_C3895_, new_C3896_, new_C3897_, new_C3898_, new_C3899_, new_C3900_,
    new_C3901_, new_C3902_, new_C3903_, new_C3904_, new_C3905_, new_C3906_,
    new_C3907_, new_C3908_, new_C3909_, new_C3910_, new_C3911_, new_C3912_,
    new_C3913_, new_C3914_, new_C3915_, new_C3916_, new_C3917_, new_C3918_,
    new_C3919_, new_C3920_, new_C3921_, new_C3922_, new_C3923_, new_C3924_,
    new_C3925_, new_C3926_, new_C3927_, new_C3928_, new_C3929_, new_C3930_,
    new_C3931_, new_C3932_, new_C3933_, new_C3934_, new_C3935_, new_C3936_,
    new_C3937_, new_C3938_, new_C3939_, new_C3940_, new_C3941_, new_C3942_,
    new_C3943_, new_C3944_, new_C3945_, new_C3946_, new_C3947_, new_C3948_,
    new_C3949_, new_C3950_, new_C3951_, new_C3952_, new_C3953_, new_C3954_,
    new_C3955_, new_C3956_, new_C3957_, new_C3958_, new_C3959_, new_C3960_,
    new_C3961_, new_C3962_, new_C3963_, new_C3964_, new_C3965_, new_C3966_,
    new_C3967_, new_C3968_, new_C3969_, new_C3970_, new_C3971_, new_C3972_,
    new_C3973_, new_C3974_, new_C3975_, new_C3976_, new_C3977_, new_C3978_,
    new_C3979_, new_C3980_, new_C3981_, new_C3982_, new_C3983_, new_C3984_,
    new_C3985_, new_C3986_, new_C3987_, new_C3988_, new_C3989_, new_C3990_,
    new_C3991_, new_C3992_, new_C3993_, new_C3994_, new_C3995_, new_C3996_,
    new_C3997_, new_C3998_, new_C3999_, new_C4000_, new_C4001_, new_C4002_,
    new_C4003_, new_C4004_, new_C4005_, new_C4006_, new_C4007_, new_C4008_,
    new_C4009_, new_C4010_, new_C4011_, new_C4012_, new_C4013_, new_C4014_,
    new_C4015_, new_C4016_, new_C4017_, new_C4018_, new_C4019_, new_C4020_,
    new_C4021_, new_C4022_, new_C4023_, new_C4024_, new_C4025_, new_C4026_,
    new_C4027_, new_C4028_, new_C4029_, new_C4030_, new_C4031_, new_C4032_,
    new_C4033_, new_C4034_, new_C4035_, new_C4036_, new_C4037_, new_C4038_,
    new_C4039_, new_C4040_, new_C4041_, new_C4042_, new_C4043_, new_C4044_,
    new_C4045_, new_C4046_, new_C4047_, new_C4048_, new_C4049_, new_C4050_,
    new_C4051_, new_C4052_, new_C4053_, new_C4054_, new_C4055_, new_C4056_,
    new_C4057_, new_C4058_, new_C4059_, new_C4060_, new_C4061_, new_C4062_,
    new_C4063_, new_C4064_, new_C4065_, new_C4066_, new_C4067_, new_C4068_,
    new_C4069_, new_C4070_, new_C4071_, new_C4072_, new_C4073_, new_C4074_,
    new_C4075_, new_C4076_, new_C4077_, new_C4078_, new_C4079_, new_C4080_,
    new_C4081_, new_C4082_, new_C4083_, new_C4084_, new_C4085_, new_C4086_,
    new_C4087_, new_C4088_, new_C4089_, new_C4090_, new_C4091_, new_C4092_,
    new_C4093_, new_C4094_, new_C4095_, new_C4096_, new_C4097_, new_C4098_,
    new_C4099_, new_C4100_, new_C4101_, new_C4102_, new_C4103_, new_C4104_,
    new_C4105_, new_C4106_, new_C4107_, new_C4108_, new_C4109_, new_C4110_,
    new_C4111_, new_C4112_, new_C4113_, new_C4114_, new_C4115_, new_C4116_,
    new_C4117_, new_C4118_, new_C4119_, new_C4120_, new_C4121_, new_C4122_,
    new_C4123_, new_C4124_, new_C4125_, new_C4126_, new_C4127_, new_C4128_,
    new_C4129_, new_C4130_, new_C4131_, new_C4132_, new_C4133_, new_C4134_,
    new_C4135_, new_C4136_, new_C4137_, new_C4138_, new_C4139_, new_C4140_,
    new_C4141_, new_C4142_, new_C4143_, new_C4144_, new_C4145_, new_C4146_,
    new_C4147_, new_C4148_, new_C4149_, new_C4150_, new_C4151_, new_C4152_,
    new_C4153_, new_C4154_, new_C4155_, new_C4156_, new_C4157_, new_C4158_,
    new_C4159_, new_C4160_, new_C4161_, new_C4162_, new_C4163_, new_C4164_,
    new_C4165_, new_C4166_, new_C4167_, new_C4168_, new_C4169_, new_C4170_,
    new_C4171_, new_C4172_, new_C4173_, new_C4174_, new_C4175_, new_C4176_,
    new_C4177_, new_C4178_, new_C4179_, new_C4180_, new_C4181_, new_C4182_,
    new_C4183_, new_C4184_, new_C4185_, new_C4186_, new_C4187_, new_C4188_,
    new_C4189_, new_C4190_, new_C4191_, new_C4192_, new_C4193_, new_C4194_,
    new_C4195_, new_C4196_, new_C4197_, new_C4198_, new_C4199_, new_C4200_,
    new_C4201_, new_C4202_, new_C4203_, new_C4204_, new_C4205_, new_C4206_,
    new_C4207_, new_C4208_, new_C4209_, new_C4210_, new_C4211_, new_C4212_,
    new_C4213_, new_C4214_, new_C4215_, new_C4216_, new_C4217_, new_C4218_,
    new_C4219_, new_C4220_, new_C4221_, new_C4222_, new_C4223_, new_C4224_,
    new_C4225_, new_C4226_, new_C4227_, new_C4228_, new_C4229_, new_C4230_,
    new_C4231_, new_C4232_, new_C4233_, new_C4234_, new_C4235_, new_C4236_,
    new_C4237_, new_C4238_, new_C4239_, new_C4240_, new_C4241_, new_C4242_,
    new_C4243_, new_C4244_, new_C4245_, new_C4246_, new_C4247_, new_C4248_,
    new_C4249_, new_C4250_, new_C4251_, new_C4252_, new_C4253_, new_C4254_,
    new_C4255_, new_C4256_, new_C4257_, new_C4258_, new_C4259_, new_C4260_,
    new_C4261_, new_C4262_, new_C4263_, new_C4264_, new_C4265_, new_C4266_,
    new_C4267_, new_C4268_, new_C4269_, new_C4270_, new_C4271_, new_C4272_,
    new_C4273_, new_C4274_, new_C4275_, new_C4276_, new_C4277_, new_C4278_,
    new_C4279_, new_C4280_, new_C4281_, new_C4282_, new_C4283_, new_C4284_,
    new_C4285_, new_C4286_, new_C4287_, new_C4288_, new_C4289_, new_C4290_,
    new_C4291_, new_C4292_, new_C4293_, new_C4294_, new_C4295_, new_C4296_,
    new_C4297_, new_C4298_, new_C4299_, new_C4300_, new_C4301_, new_C4302_,
    new_C4303_, new_C4304_, new_C4305_, new_C4306_, new_C4307_, new_C4308_,
    new_C4309_, new_C4310_, new_C4311_, new_C4312_, new_C4313_, new_C4314_,
    new_C4315_, new_C4316_, new_C4317_, new_C4318_, new_C4319_, new_C4320_,
    new_C4321_, new_C4322_, new_C4323_, new_C4324_, new_C4325_, new_C4326_,
    new_C4327_, new_C4328_, new_C4329_, new_C4330_, new_C4331_, new_C4332_,
    new_C4333_, new_C4334_, new_C4335_, new_C4336_, new_C4337_, new_C4338_,
    new_C4339_, new_C4340_, new_C4341_, new_C4342_, new_C4343_, new_C4344_,
    new_C4345_, new_C4346_, new_C4347_, new_C4348_, new_C4349_, new_C4350_,
    new_C4351_, new_C4352_, new_C4353_, new_C4354_, new_C4355_, new_C4356_,
    new_C4357_, new_C4358_, new_C4359_, new_C4360_, new_C4361_, new_C4362_,
    new_C4363_, new_C4364_, new_C4365_, new_C4366_, new_C4367_, new_C4368_,
    new_C4369_, new_C4370_, new_C4371_, new_C4372_, new_C4373_, new_C4374_,
    new_C4375_, new_C4376_, new_C4377_, new_C4378_, new_C4379_, new_C4380_,
    new_C4381_, new_C4382_, new_C4383_, new_C4384_, new_C4385_, new_C4386_,
    new_C4387_, new_C4388_, new_C4389_, new_C4390_, new_C4391_, new_C4392_,
    new_C4393_, new_C4394_, new_C4395_, new_C4396_, new_C4397_, new_C4398_,
    new_C4399_, new_C4400_, new_C4401_, new_C4402_, new_C4403_, new_C4404_,
    new_C4405_, new_C4406_, new_C4407_, new_C4408_, new_C4409_, new_C4410_,
    new_C4411_, new_C4412_, new_C4413_, new_C4414_, new_C4415_, new_C4416_,
    new_C4417_, new_C4418_, new_C4419_, new_C4420_, new_C4421_, new_C4422_,
    new_C4423_, new_C4424_, new_C4425_, new_C4426_, new_C4427_, new_C4428_,
    new_C4429_, new_C4430_, new_C4431_, new_C4432_, new_C4433_, new_C4434_,
    new_C4435_, new_C4436_, new_C4437_, new_C4438_, new_C4439_, new_C4440_,
    new_C4441_, new_C4442_, new_C4443_, new_C4444_, new_C4445_, new_C4446_,
    new_C4447_, new_C4448_, new_C4449_, new_C4450_, new_C4451_, new_C4452_,
    new_C4453_, new_C4454_, new_C4455_, new_C4456_, new_C4457_, new_C4458_,
    new_C4459_, new_C4460_, new_C4461_, new_C4462_, new_C4463_, new_C4464_,
    new_C4465_, new_C4466_, new_C4467_, new_C4468_, new_C4469_, new_C4470_,
    new_C4471_, new_C4472_, new_C4473_, new_C4474_, new_C4475_, new_C4476_,
    new_C4477_, new_C4478_, new_C4479_, new_C4480_, new_C4481_, new_C4482_,
    new_C4483_, new_C4484_, new_C4485_, new_C4486_, new_C4487_, new_C4488_,
    new_C4489_, new_C4490_, new_C4491_, new_C4492_, new_C4493_, new_C4494_,
    new_C4495_, new_C4496_, new_C4497_, new_C4498_, new_C4499_, new_C4500_,
    new_C4501_, new_C4502_, new_C4503_, new_C4504_, new_C4505_, new_C4506_,
    new_C4507_, new_C4508_, new_C4509_, new_C4510_, new_C4511_, new_C4512_,
    new_C4513_, new_C4514_, new_C4515_, new_C4516_, new_C4517_, new_C4518_,
    new_C4519_, new_C4520_, new_C4521_, new_C4522_, new_C4523_, new_C4524_,
    new_C4525_, new_C4526_, new_C4527_, new_C4528_, new_C4529_, new_C4530_,
    new_C4531_, new_C4532_, new_C4533_, new_C4534_, new_C4535_, new_C4536_,
    new_C4537_, new_C4538_, new_C4539_, new_C4540_, new_C4541_, new_C4542_,
    new_C4543_, new_C4544_, new_C4545_, new_C4546_, new_C4547_, new_C4548_,
    new_C4549_, new_C4550_, new_C4551_, new_C4552_, new_C4553_, new_C4554_,
    new_C4555_, new_C4556_, new_C4557_, new_C4558_, new_C4559_, new_C4560_,
    new_C4561_, new_C4562_, new_C4563_, new_C4564_, new_C4565_, new_C4566_,
    new_C4567_, new_C4568_, new_C4569_, new_C4570_, new_C4571_, new_C4572_,
    new_C4573_, new_C4574_, new_C4575_, new_C4576_, new_C4577_, new_C4578_,
    new_C4579_, new_C4580_, new_C4581_, new_C4582_, new_C4583_, new_C4584_,
    new_C4585_, new_C4586_, new_C4587_, new_C4588_, new_C4589_, new_C4590_,
    new_C4591_, new_C4592_, new_C4593_, new_C4594_, new_C4595_, new_C4596_,
    new_C4597_, new_C4598_, new_C4599_, new_C4600_, new_C4601_, new_C4602_,
    new_C4603_, new_C4604_, new_C4605_, new_C4606_, new_C4607_, new_C4608_,
    new_C4609_, new_C4610_, new_C4611_, new_C4612_, new_C4613_, new_C4614_,
    new_C4615_, new_C4616_, new_C4617_, new_C4618_, new_C4619_, new_C4620_,
    new_C4621_, new_C4622_, new_C4623_, new_C4624_, new_C4625_, new_C4626_,
    new_C4627_, new_C4628_, new_C4629_, new_C4630_, new_C4631_, new_C4632_,
    new_C4633_, new_C4634_, new_C4635_, new_C4636_, new_C4637_, new_C4638_,
    new_C4639_, new_C4640_, new_C4641_, new_C4642_, new_C4643_, new_C4644_,
    new_C4645_, new_C4646_, new_C4647_, new_C4648_, new_C4649_, new_C4650_,
    new_C4651_, new_C4652_, new_C4653_, new_C4654_, new_C4655_, new_C4656_,
    new_C4657_, new_C4658_, new_C4659_, new_C4660_, new_C4661_, new_C4662_,
    new_C4663_, new_C4664_, new_C4665_, new_C4666_, new_C4667_, new_C4668_,
    new_C4669_, new_C4670_, new_C4671_, new_C4672_, new_C4673_, new_C4674_,
    new_C4675_, new_C4676_, new_C4677_, new_C4678_, new_C4679_, new_C4680_,
    new_C4681_, new_C4682_, new_C4683_, new_C4684_, new_C4685_, new_C4686_,
    new_C4687_, new_C4688_, new_C4689_, new_C4690_, new_C4691_, new_C4692_,
    new_C4693_, new_C4694_, new_C4695_, new_C4696_, new_C4697_, new_C4698_,
    new_C4699_, new_C4700_, new_C4701_, new_C4702_, new_C4703_, new_C4704_,
    new_C4705_, new_C4706_, new_C4707_, new_C4708_, new_C4709_, new_C4710_,
    new_C4711_, new_C4712_, new_C4713_, new_C4714_, new_C4715_, new_C4716_,
    new_C4717_, new_C4718_, new_C4719_, new_C4720_, new_C4721_, new_C4722_,
    new_C4723_, new_C4724_, new_C4725_, new_C4726_, new_C4727_, new_C4728_,
    new_C4729_, new_C4730_, new_C4731_, new_C4732_, new_C4733_, new_C4734_,
    new_C4735_, new_C4736_, new_C4737_, new_C4738_, new_C4739_, new_C4740_,
    new_C4741_, new_C4742_, new_C4743_, new_C4744_, new_C4745_, new_C4746_,
    new_C4747_, new_C4748_, new_C4749_, new_C4750_, new_C4751_, new_C4752_,
    new_C4753_, new_C4754_, new_C4755_, new_C4756_, new_C4757_, new_C4758_,
    new_C4759_, new_C4760_, new_C4761_, new_C4762_, new_C4763_, new_C4764_,
    new_C4765_, new_C4766_, new_C4767_, new_C4768_, new_C4769_, new_C4770_,
    new_C4771_, new_C4772_, new_C4773_, new_C4774_, new_C4775_, new_C4776_,
    new_C4777_, new_C4778_, new_C4779_, new_C4780_, new_C4781_, new_C4782_,
    new_C4783_, new_C4784_, new_C4785_, new_C4786_, new_C4787_, new_C4788_,
    new_C4789_, new_C4790_, new_C4791_, new_C4792_, new_C4793_, new_C4794_,
    new_C4795_, new_C4796_, new_C4797_, new_C4798_, new_C4799_, new_C4800_,
    new_C4801_, new_C4802_, new_C4803_, new_C4804_, new_C4805_, new_C4806_,
    new_C4807_, new_C4808_, new_C4809_, new_C4810_, new_C4811_, new_C4812_,
    new_C4813_, new_C4814_, new_C4815_, new_C4816_, new_C4817_, new_C4818_,
    new_C4819_, new_C4820_, new_C4821_, new_C4822_, new_C4823_, new_C4824_,
    new_C4825_, new_C4826_, new_C4827_, new_C4828_, new_C4829_, new_C4830_,
    new_C4831_, new_C4832_, new_C4833_, new_C4834_, new_C4835_, new_C4836_,
    new_C4837_, new_C4838_, new_C4839_, new_C4840_, new_C4841_, new_C4842_,
    new_C4843_, new_C4844_, new_C4845_, new_C4846_, new_C4847_, new_C4848_,
    new_C4849_, new_C4850_, new_C4851_, new_C4852_, new_C4853_, new_C4854_,
    new_C4855_, new_C4856_, new_C4857_, new_C4858_, new_C4859_, new_C4860_,
    new_C4861_, new_C4862_, new_C4863_, new_C4864_, new_C4865_, new_C4866_,
    new_C4867_, new_C4868_, new_C4869_, new_C4870_, new_C4871_, new_C4872_,
    new_C4873_, new_C4874_, new_C4875_, new_C4876_, new_C4877_, new_C4878_,
    new_C4879_, new_C4880_, new_C4881_, new_C4882_, new_C4883_, new_C4884_,
    new_C4885_, new_C4886_, new_C4887_, new_C4888_, new_C4889_, new_C4890_,
    new_C4891_, new_C4892_, new_C4893_, new_C4894_, new_C4895_, new_C4896_,
    new_C4897_, new_C4898_, new_C4899_, new_C4900_, new_C4901_, new_C4902_,
    new_C4903_, new_C4904_, new_C4905_, new_C4906_, new_C4907_, new_C4908_,
    new_C4909_, new_C4910_, new_C4911_, new_C4912_, new_C4913_, new_C4914_,
    new_C4915_, new_C4916_, new_C4917_, new_C4918_, new_C4919_, new_C4920_,
    new_C4921_, new_C4922_, new_C4923_, new_C4924_, new_C4925_, new_C4926_,
    new_C4927_, new_C4928_, new_C4929_, new_C4930_, new_C4931_, new_C4932_,
    new_C4933_, new_C4934_, new_C4935_, new_C4936_, new_C4937_, new_C4938_,
    new_C4939_, new_C4940_, new_C4941_, new_C4942_, new_C4943_, new_C4944_,
    new_C4945_, new_C4946_, new_C4947_, new_C4948_, new_C4949_, new_C4950_,
    new_C4951_, new_C4952_, new_C4953_, new_C4954_, new_C4955_, new_C4956_,
    new_C4957_, new_C4958_, new_C4959_, new_C4960_, new_C4961_, new_C4962_,
    new_C4963_, new_C4964_, new_C4965_, new_C4966_, new_C4967_, new_C4968_,
    new_C4969_, new_C4970_, new_C4971_, new_C4972_, new_C4973_, new_C4974_,
    new_C4975_, new_C4976_, new_C4977_, new_C4978_, new_C4979_, new_C4980_,
    new_C4981_, new_C4982_, new_C4983_, new_C4984_, new_C4985_, new_C4986_,
    new_C4987_, new_C4988_, new_C4989_, new_C4990_, new_C4991_, new_C4992_,
    new_C4993_, new_C4994_, new_C4995_, new_C4996_, new_C4997_, new_C4998_,
    new_C4999_, new_C5000_, new_C5001_, new_C5002_, new_C5003_, new_C5004_,
    new_C5005_, new_C5006_, new_C5007_, new_C5008_, new_C5009_, new_C5010_,
    new_C5011_, new_C5012_, new_C5013_, new_C5014_, new_C5015_, new_C5016_,
    new_C5017_, new_C5018_, new_C5019_, new_C5020_, new_C5021_, new_C5022_,
    new_C5023_, new_C5024_, new_C5025_, new_C5026_, new_C5027_, new_C5028_,
    new_C5029_, new_C5030_, new_C5031_, new_C5032_, new_C5033_, new_C5034_,
    new_C5035_, new_C5036_, new_C5037_, new_C5038_, new_C5039_, new_C5040_,
    new_C5041_, new_C5042_, new_C5043_, new_C5044_, new_C5045_, new_C5046_,
    new_C5047_, new_C5048_, new_C5049_, new_C5050_, new_C5051_, new_C5052_,
    new_C5053_, new_C5054_, new_C5055_, new_C5056_, new_C5057_, new_C5058_,
    new_C5059_, new_C5060_, new_C5061_, new_C5062_, new_C5063_, new_C5064_,
    new_C5065_, new_C5066_, new_C5067_, new_C5068_, new_C5069_, new_C5070_,
    new_C5071_, new_C5072_, new_C5073_, new_C5074_, new_C5075_, new_C5076_,
    new_C5077_, new_C5078_, new_C5079_, new_C5080_, new_C5081_, new_C5082_,
    new_C5083_, new_C5084_, new_C5085_, new_C5086_, new_C5087_, new_C5088_,
    new_C5089_, new_C5090_, new_C5091_, new_C5092_, new_C5093_, new_C5094_,
    new_C5095_, new_C5096_, new_C5097_, new_C5098_, new_C5099_, new_C5100_,
    new_C5101_, new_C5102_, new_C5103_, new_C5104_, new_C5105_, new_C5106_,
    new_C5107_, new_C5108_, new_C5109_, new_C5110_, new_C5111_, new_C5112_,
    new_C5113_, new_C5114_, new_C5115_, new_C5116_, new_C5117_, new_C5118_,
    new_C5119_, new_C5120_, new_C5121_, new_C5122_, new_C5123_, new_C5124_,
    new_C5125_, new_C5126_, new_C5127_, new_C5128_, new_C5129_, new_C5130_,
    new_C5131_, new_C5132_, new_C5133_, new_C5134_, new_C5135_, new_C5136_,
    new_C5137_, new_C5138_, new_C5139_, new_C5140_, new_C5141_, new_C5142_,
    new_C5143_, new_C5144_, new_C5145_, new_C5146_, new_C5147_, new_C5148_,
    new_C5149_, new_C5150_, new_C5151_, new_C5152_, new_C5153_, new_C5154_,
    new_C5155_, new_C5156_, new_C5157_, new_C5158_, new_C5159_, new_C5160_,
    new_C5161_, new_C5162_, new_C5163_, new_C5164_, new_C5165_, new_C5166_,
    new_C5167_, new_C5168_, new_C5169_, new_C5170_, new_C5171_, new_C5172_,
    new_C5173_, new_C5174_, new_C5175_, new_C5176_, new_C5177_, new_C5178_,
    new_C5179_, new_C5180_, new_C5181_, new_C5182_, new_C5183_, new_C5184_,
    new_C5185_, new_C5186_, new_C5187_, new_C5188_, new_C5189_, new_C5190_,
    new_C5191_, new_C5192_, new_C5193_, new_C5194_, new_C5195_, new_C5196_,
    new_C5197_, new_C5198_, new_C5199_, new_C5200_, new_C5201_, new_C5202_,
    new_C5203_, new_C5204_, new_C5205_, new_C5206_, new_C5207_, new_C5208_,
    new_C5209_, new_C5210_, new_C5211_, new_C5212_, new_C5213_, new_C5214_,
    new_C5215_, new_C5216_, new_C5217_, new_C5218_, new_C5219_, new_C5220_,
    new_C5221_, new_C5222_, new_C5223_, new_C5224_, new_C5225_, new_C5226_,
    new_C5227_, new_C5228_, new_C5229_, new_C5230_, new_C5231_, new_C5232_,
    new_C5233_, new_C5234_, new_C5235_, new_C5236_, new_C5237_, new_C5238_,
    new_C5239_, new_C5240_, new_C5241_, new_C5242_, new_C5243_, new_C5244_,
    new_C5245_, new_C5246_, new_C5247_, new_C5248_, new_C5249_, new_C5250_,
    new_C5251_, new_C5252_, new_C5253_, new_C5254_, new_C5255_, new_C5256_,
    new_C5257_, new_C5258_, new_C5259_, new_C5260_, new_C5261_, new_C5262_,
    new_C5263_, new_C5264_, new_C5265_, new_C5266_, new_C5267_, new_C5268_,
    new_C5269_, new_C5270_, new_C5271_, new_C5272_, new_C5273_, new_C5274_,
    new_C5275_, new_C5276_, new_C5277_, new_C5278_, new_C5279_, new_C5280_,
    new_C5281_, new_C5282_, new_C5283_, new_C5284_, new_C5285_, new_C5286_,
    new_C5287_, new_C5288_, new_C5289_, new_C5290_, new_C5291_, new_C5292_,
    new_C5293_, new_C5294_, new_C5295_, new_C5296_, new_C5297_, new_C5298_,
    new_C5299_, new_C5300_, new_C5301_, new_C5302_, new_C5303_, new_C5304_,
    new_C5305_, new_C5306_, new_C5307_, new_C5308_, new_C5309_, new_C5310_,
    new_C5311_, new_C5312_, new_C5313_, new_C5314_, new_C5315_, new_C5316_,
    new_C5317_, new_C5318_, new_C5319_, new_C5320_, new_C5321_, new_C5322_,
    new_C5323_, new_C5324_, new_C5325_, new_C5326_, new_C5327_, new_C5328_,
    new_C5329_, new_C5330_, new_C5331_, new_C5332_, new_C5333_, new_C5334_,
    new_C5335_, new_C5336_, new_C5337_, new_C5338_, new_C5339_, new_C5340_,
    new_C5341_, new_C5342_, new_C5343_, new_C5344_, new_C5345_, new_C5346_,
    new_C5347_, new_C5348_, new_C5349_, new_C5350_, new_C5351_, new_C5352_,
    new_C5353_, new_C5354_, new_C5355_, new_C5356_, new_C5357_, new_C5358_,
    new_C5359_, new_C5360_, new_C5361_, new_C5362_, new_C5363_, new_C5364_,
    new_C5365_, new_C5366_, new_C5367_, new_C5368_, new_C5369_, new_C5370_,
    new_C5371_, new_C5372_, new_C5373_, new_C5374_, new_C5375_, new_C5376_,
    new_C5377_, new_C5378_, new_C5379_, new_C5380_, new_C5381_, new_C5382_,
    new_C5383_, new_C5384_, new_C5385_, new_C5386_, new_C5387_, new_C5388_,
    new_C5389_, new_C5390_, new_C5391_, new_C5392_, new_C5393_, new_C5394_,
    new_C5395_, new_C5396_, new_C5397_, new_C5398_, new_C5399_, new_C5400_,
    new_C5401_, new_C5402_, new_C5403_, new_C5404_, new_C5405_, new_C5406_,
    new_C5407_, new_C5408_, new_C5409_, new_C5410_, new_C5411_, new_C5412_,
    new_C5413_, new_C5414_, new_C5415_, new_C5416_, new_C5417_, new_C5418_,
    new_C5419_, new_C5420_, new_C5421_, new_C5422_, new_C5423_, new_C5424_,
    new_C5425_, new_C5426_, new_C5427_, new_C5428_, new_C5429_, new_C5430_,
    new_C5431_, new_C5432_, new_C5433_, new_C5434_, new_C5435_, new_C5436_,
    new_C5437_, new_C5438_, new_C5439_, new_C5440_, new_C5441_, new_C5442_,
    new_C5443_, new_C5444_, new_C5445_, new_C5446_, new_C5447_, new_C5448_,
    new_C5449_, new_C5450_, new_C5451_, new_C5452_, new_C5453_, new_C5454_,
    new_C5455_, new_C5456_, new_C5457_, new_C5458_, new_C5459_, new_C5460_,
    new_C5461_, new_C5462_, new_C5463_, new_C5464_, new_C5465_, new_C5466_,
    new_C5467_, new_C5468_, new_C5469_, new_C5470_, new_C5471_, new_C5472_,
    new_C5473_, new_C5474_, new_C5475_, new_C5476_, new_C5477_, new_C5478_,
    new_C5479_, new_C5480_, new_C5481_, new_C5482_, new_C5483_, new_C5484_,
    new_C5485_, new_C5486_, new_C5487_, new_C5488_, new_C5489_, new_C5490_,
    new_C5491_, new_C5492_, new_C5493_, new_C5494_, new_C5495_, new_C5496_,
    new_C5497_, new_C5498_, new_C5499_, new_C5500_, new_C5501_, new_C5502_,
    new_C5503_, new_C5504_, new_C5505_, new_C5506_, new_C5507_, new_C5508_,
    new_C5509_, new_C5510_, new_C5511_, new_C5512_, new_C5513_, new_C5514_,
    new_C5515_, new_C5516_, new_C5517_, new_C5518_, new_C5519_, new_C5520_,
    new_C5521_, new_C5522_, new_C5523_, new_C5524_, new_C5525_, new_C5526_,
    new_C5527_, new_C5528_, new_C5529_, new_C5530_, new_C5531_, new_C5532_,
    new_C5533_, new_C5534_, new_C5535_, new_C5536_, new_C5537_, new_C5538_,
    new_C5539_, new_C5540_, new_C5541_, new_C5542_, new_C5543_, new_C5544_,
    new_C5545_, new_C5546_, new_C5547_, new_C5548_, new_C5549_, new_C5550_,
    new_C5551_, new_C5552_, new_C5553_, new_C5554_, new_C5555_, new_C5556_,
    new_C5557_, new_C5558_, new_C5559_, new_C5560_, new_C5561_, new_C5562_,
    new_C5563_, new_C5564_, new_C5565_, new_C5566_, new_C5567_, new_C5568_,
    new_C5569_, new_C5570_, new_C5571_, new_C5572_, new_C5573_, new_C5574_,
    new_C5575_, new_C5576_, new_C5577_, new_C5578_, new_C5579_, new_C5580_,
    new_C5581_, new_C5582_, new_C5583_, new_C5584_, new_C5585_, new_C5586_,
    new_C5587_, new_C5588_, new_C5589_, new_C5590_, new_C5591_, new_C5592_,
    new_C5593_, new_C5594_, new_C5595_, new_C5596_, new_C5597_, new_C5598_,
    new_C5599_, new_C5600_, new_C5601_, new_C5602_, new_C5603_, new_C5604_,
    new_C5605_, new_C5606_, new_C5607_, new_C5608_, new_C5609_, new_C5610_,
    new_C5611_, new_C5612_, new_C5613_, new_C5614_, new_C5615_, new_C5616_,
    new_C5617_, new_C5618_, new_C5619_, new_C5620_, new_C5621_, new_C5622_,
    new_C5623_, new_C5624_, new_C5625_, new_C5626_, new_C5627_, new_C5628_,
    new_C5629_, new_C5630_, new_C5631_, new_C5632_, new_C5633_, new_C5634_,
    new_C5635_, new_C5636_, new_C5637_, new_C5638_, new_C5639_, new_C5640_,
    new_C5641_, new_C5642_, new_C5643_, new_C5644_, new_C5645_, new_C5646_,
    new_C5647_, new_C5648_, new_C5649_, new_C5650_, new_C5651_, new_C5652_,
    new_C5653_, new_C5654_, new_C5655_, new_C5656_, new_C5657_, new_C5658_,
    new_C5659_, new_C5660_, new_C5661_, new_C5662_, new_C5663_, new_C5664_,
    new_C5665_, new_C5666_, new_C5667_, new_C5668_, new_C5669_, new_C5670_,
    new_C5671_, new_C5672_, new_C5673_, new_C5674_, new_C5675_, new_C5676_,
    new_C5677_, new_C5678_, new_C5679_, new_C5680_, new_C5681_, new_C5682_,
    new_C5683_, new_C5684_, new_C5685_, new_C5686_, new_C5687_, new_C5688_,
    new_C5689_, new_C5690_, new_C5691_, new_C5692_, new_C5693_, new_C5694_,
    new_C5695_, new_C5696_, new_C5697_, new_C5698_, new_C5699_, new_C5700_,
    new_C5701_, new_C5702_, new_C5703_, new_C5704_, new_C5705_, new_C5706_,
    new_C5707_, new_C5708_, new_C5709_, new_C5710_, new_C5711_, new_C5712_,
    new_C5713_, new_C5714_, new_C5715_, new_C5716_, new_C5717_, new_C5718_,
    new_C5719_, new_C5720_, new_C5721_, new_C5722_, new_C5723_, new_C5724_,
    new_C5725_, new_C5726_, new_C5727_, new_C5728_, new_C5729_, new_C5730_,
    new_C5731_, new_C5732_, new_C5733_, new_C5734_, new_C5735_, new_C5736_,
    new_C5737_, new_C5738_, new_C5739_, new_C5740_, new_C5741_, new_C5742_,
    new_C5743_, new_C5744_, new_C5745_, new_C5746_, new_C5747_, new_C5748_,
    new_C5749_, new_C5750_, new_C5751_, new_C5752_, new_C5753_, new_C5754_,
    new_C5755_, new_C5756_, new_C5757_, new_C5758_, new_C5759_, new_C5760_,
    new_C5761_, new_C5762_, new_C5763_, new_C5764_, new_C5765_, new_C5766_,
    new_C5767_, new_C5768_, new_C5769_, new_C5770_, new_C5771_, new_C5772_,
    new_C5773_, new_C5774_, new_C5775_, new_C5776_, new_C5777_, new_C5778_,
    new_C5779_, new_C5780_, new_C5781_, new_C5782_, new_C5783_, new_C5784_,
    new_C5785_, new_C5786_, new_C5787_, new_C5788_, new_C5789_, new_C5790_,
    new_C5791_, new_C5792_, new_C5793_, new_C5794_, new_C5795_, new_C5796_,
    new_C5797_, new_C5798_, new_C5799_, new_C5800_, new_C5801_, new_C5802_,
    new_C5803_, new_C5804_, new_C5805_, new_C5806_, new_C5807_, new_C5808_,
    new_C5809_, new_C5810_, new_C5811_, new_C5812_, new_C5813_, new_C5814_,
    new_C5815_, new_C5816_, new_C5817_, new_C5818_, new_C5819_, new_C5820_,
    new_C5821_, new_C5822_, new_C5823_, new_C5824_, new_C5825_, new_C5826_,
    new_C5827_, new_C5828_, new_C5829_, new_C5830_, new_C5831_, new_C5832_,
    new_C5833_, new_C5834_, new_C5835_, new_C5836_, new_C5837_, new_C5838_,
    new_C5839_, new_C5840_, new_C5841_, new_C5842_, new_C5843_, new_C5844_,
    new_C5845_, new_C5846_, new_C5847_, new_C5848_, new_C5849_, new_C5850_,
    new_C5851_, new_C5852_, new_C5853_, new_C5854_, new_C5855_, new_C5856_,
    new_C5857_, new_C5858_, new_C5859_, new_C5860_, new_C5861_, new_C5862_,
    new_C5863_, new_C5864_, new_C5865_, new_C5866_, new_C5867_, new_C5868_,
    new_C5869_, new_C5870_, new_C5871_, new_C5872_, new_C5873_, new_C5874_,
    new_C5875_, new_C5876_, new_C5877_, new_C5878_, new_C5879_, new_C5880_,
    new_C5881_, new_C5882_, new_C5883_, new_C5884_, new_C5885_, new_C5886_,
    new_C5887_, new_C5888_, new_C5889_, new_C5890_, new_C5891_, new_C5892_,
    new_C5893_, new_C5894_, new_C5895_, new_C5896_, new_C5897_, new_C5898_,
    new_C5899_, new_C5900_, new_C5901_, new_C5902_, new_C5903_, new_C5904_,
    new_C5905_, new_C5906_, new_C5907_, new_C5908_, new_C5909_, new_C5910_,
    new_C5911_, new_C5912_, new_C5913_, new_C5914_, new_C5915_, new_C5916_,
    new_C5917_, new_C5918_, new_C5919_, new_C5920_, new_C5921_, new_C5922_,
    new_C5923_, new_C5924_, new_C5925_, new_C5926_, new_C5927_, new_C5928_,
    new_C5929_, new_C5930_, new_C5931_, new_C5932_, new_C5933_, new_C5934_,
    new_C5935_, new_C5936_, new_C5937_, new_C5938_, new_C5939_, new_C5940_,
    new_C5941_, new_C5942_, new_C5943_, new_C5944_, new_C5945_, new_C5946_,
    new_C5947_, new_C5948_, new_C5949_, new_C5950_, new_C5951_, new_C5952_,
    new_C5953_, new_C5954_, new_C5955_, new_C5956_, new_C5957_, new_C5958_,
    new_C5959_, new_C5960_, new_C5961_, new_C5962_, new_C5963_, new_C5964_,
    new_C5965_, new_C5966_, new_C5967_, new_C5968_, new_C5969_, new_C5970_,
    new_C5971_, new_C5972_, new_C5973_, new_C5974_, new_C5975_, new_C5976_,
    new_C5977_, new_C5978_, new_C5979_, new_C5980_, new_C5981_, new_C5982_,
    new_C5983_, new_C5984_, new_C5985_, new_C5986_, new_C5987_, new_C5988_,
    new_C5989_, new_C5990_, new_C5991_, new_C5992_, new_C5993_, new_C5994_,
    new_C5995_, new_C5996_, new_C5997_, new_C5998_, new_C5999_, new_C6000_,
    new_C6001_, new_C6002_, new_C6003_, new_C6004_, new_C6005_, new_C6006_,
    new_C6007_, new_C6008_, new_C6009_, new_C6010_, new_C6011_, new_C6012_,
    new_C6013_, new_C6014_, new_C6015_, new_C6016_, new_C6017_, new_C6018_,
    new_C6019_, new_C6020_, new_C6021_, new_C6022_, new_C6023_, new_C6024_,
    new_C6025_, new_C6026_, new_C6027_, new_C6028_, new_C6029_, new_C6030_,
    new_C6031_, new_C6032_, new_C6033_, new_C6034_, new_C6035_, new_C6036_,
    new_C6037_, new_C6038_, new_C6039_, new_C6040_, new_C6041_, new_C6042_,
    new_C6043_, new_C6044_, new_C6045_, new_C6046_, new_C6047_, new_C6048_,
    new_C6049_, new_C6050_, new_C6051_, new_C6052_, new_C6053_, new_C6054_,
    new_C6055_, new_C6056_, new_C6057_, new_C6058_, new_C6059_, new_C6060_,
    new_C6061_, new_C6062_, new_C6063_, new_C6064_, new_C6065_, new_C6066_,
    new_C6067_, new_C6068_, new_C6069_, new_C6070_, new_C6071_, new_C6072_,
    new_C6073_, new_C6074_, new_C6075_, new_C6076_, new_C6077_, new_C6078_,
    new_C6079_, new_C6080_, new_C6081_, new_C6082_, new_C6083_, new_C6084_,
    new_C6085_, new_C6086_, new_C6087_, new_C6088_, new_C6089_, new_C6090_,
    new_C6091_, new_C6092_, new_C6093_, new_C6094_, new_C6095_, new_C6096_,
    new_C6097_, new_C6098_, new_C6099_, new_C6100_, new_C6101_, new_C6102_,
    new_C6103_, new_C6104_, new_C6105_, new_C6106_, new_C6107_, new_C6108_,
    new_C6109_, new_C6110_, new_C6111_, new_C6112_, new_C6113_, new_C6114_,
    new_C6115_, new_C6116_, new_C6117_, new_C6118_, new_C6119_, new_C6120_,
    new_C6121_, new_C6122_, new_C6123_, new_C6124_, new_C6125_, new_C6126_,
    new_C6127_, new_C6128_, new_C6129_, new_C6130_, new_C6131_, new_C6132_,
    new_C6133_, new_C6134_, new_C6135_, new_C6136_, new_C6137_, new_C6138_,
    new_C6139_, new_C6140_, new_C6141_, new_C6142_, new_C6143_, new_C6144_,
    new_C6145_, new_C6146_, new_C6147_, new_C6148_, new_C6149_, new_C6150_,
    new_C6151_, new_C6152_, new_C6153_, new_C6154_, new_C6155_, new_C6156_,
    new_C6157_, new_C6158_, new_C6159_, new_C6160_, new_C6161_, new_C6162_,
    new_C6163_, new_C6164_, new_C6165_, new_C6166_, new_C6167_, new_C6168_,
    new_C6169_, new_C6170_, new_C6171_, new_C6172_, new_C6173_, new_C6174_,
    new_C6175_, new_C6176_, new_C6177_, new_C6178_, new_C6179_, new_C6180_,
    new_C6181_, new_C6182_, new_C6183_, new_C6184_, new_C6185_, new_C6186_,
    new_C6187_, new_C6188_, new_C6189_, new_C6190_, new_C6191_, new_C6192_,
    new_C6193_, new_C6194_, new_C6195_, new_C6196_, new_C6197_, new_C6198_,
    new_C6199_, new_C6200_, new_C6201_, new_C6202_, new_C6203_, new_C6204_,
    new_C6205_, new_C6206_, new_C6207_, new_C6208_, new_C6209_, new_C6210_,
    new_C6211_, new_C6212_, new_C6213_, new_C6214_, new_C6215_, new_C6216_,
    new_C6217_, new_C6218_, new_C6219_, new_C6220_, new_C6221_, new_C6222_,
    new_C6223_, new_C6224_, new_C6225_, new_C6226_, new_C6227_, new_C6228_,
    new_C6229_, new_C6230_, new_C6231_, new_C6232_, new_C6233_, new_C6234_,
    new_C6235_, new_C6236_, new_C6237_, new_C6238_, new_C6239_, new_C6240_,
    new_C6241_, new_C6242_, new_C6243_, new_C6244_, new_C6245_, new_C6246_,
    new_C6247_, new_C6248_, new_C6249_, new_C6250_, new_C6251_, new_C6252_,
    new_C6253_, new_C6254_, new_C6255_, new_C6256_, new_C6257_, new_C6258_,
    new_C6259_, new_C6260_, new_C6261_, new_C6262_, new_C6263_, new_C6264_,
    new_C6265_, new_C6266_, new_C6267_, new_C6268_, new_C6269_, new_C6270_,
    new_C6271_, new_C6272_, new_C6273_, new_C6274_, new_C6275_, new_C6276_,
    new_C6277_, new_C6278_, new_C6279_, new_C6280_, new_C6281_, new_C6282_,
    new_C6283_, new_C6284_, new_C6285_, new_C6286_, new_C6287_, new_C6288_,
    new_C6289_, new_C6290_, new_C6291_, new_C6292_, new_C6293_, new_C6294_,
    new_C6295_, new_C6296_, new_C6297_, new_C6298_, new_C6299_, new_C6300_,
    new_C6301_, new_C6302_, new_C6303_, new_C6304_, new_C6305_, new_C6306_,
    new_C6307_, new_C6308_, new_C6309_, new_C6310_, new_C6311_, new_C6312_,
    new_C6313_, new_C6314_, new_C6315_, new_C6316_, new_C6317_, new_C6318_,
    new_C6319_, new_C6320_, new_C6321_, new_C6322_, new_C6323_, new_C6324_,
    new_C6325_, new_C6326_, new_C6327_, new_C6328_, new_C6329_, new_C6330_,
    new_C6331_, new_C6332_, new_C6333_, new_C6334_, new_C6335_, new_C6336_,
    new_C6337_, new_C6338_, new_C6339_, new_C6340_, new_C6341_, new_C6342_,
    new_C6343_, new_C6344_, new_C6345_, new_C6346_, new_C6347_, new_C6348_,
    new_C6349_, new_C6350_, new_C6351_, new_C6352_, new_C6353_, new_C6354_,
    new_C6355_, new_C6356_, new_C6357_, new_C6358_, new_C6359_, new_C6360_,
    new_C6361_, new_C6362_, new_C6363_, new_C6364_, new_C6365_, new_C6366_,
    new_C6367_, new_C6368_, new_C6369_, new_C6370_, new_C6371_, new_C6372_,
    new_C6373_, new_C6374_, new_C6375_, new_C6376_, new_C6377_, new_C6378_,
    new_C6379_, new_C6380_, new_C6381_, new_C6382_, new_C6383_, new_C6384_,
    new_C6385_, new_C6386_, new_C6387_, new_C6388_, new_C6389_, new_C6390_,
    new_C6391_, new_C6392_, new_C6393_, new_C6394_, new_C6395_, new_C6396_,
    new_C6397_, new_C6398_, new_C6399_, new_C6400_, new_C6401_, new_C6402_,
    new_C6403_, new_C6404_, new_C6405_, new_C6406_, new_C6407_, new_C6408_,
    new_C6409_, new_C6410_, new_C6411_, new_C6412_, new_C6413_, new_C6414_,
    new_C6415_, new_C6416_, new_C6417_, new_C6418_, new_C6419_, new_C6420_,
    new_C6421_, new_C6422_, new_C6423_, new_C6424_, new_C6425_, new_C6426_,
    new_C6427_, new_C6428_, new_C6429_, new_C6430_, new_C6431_, new_C6432_,
    new_C6433_, new_C6434_, new_C6435_, new_C6436_, new_C6437_, new_C6438_,
    new_C6439_, new_C6440_, new_C6441_, new_C6442_, new_C6443_, new_C6444_,
    new_C6445_, new_C6446_, new_C6447_, new_C6448_, new_C6449_, new_C6450_,
    new_C6451_, new_C6452_, new_C6453_, new_C6454_, new_C6455_, new_C6456_,
    new_C6457_, new_C6458_, new_C6459_, new_C6460_, new_C6461_, new_C6462_,
    new_C6463_, new_C6464_, new_C6465_, new_C6466_, new_C6467_, new_C6468_,
    new_C6469_, new_C6470_, new_C6471_, new_C6472_, new_C6473_, new_C6474_,
    new_C6475_, new_C6476_, new_C6477_, new_C6478_, new_C6479_, new_C6480_,
    new_C6481_, new_C6482_, new_C6483_, new_C6484_, new_C6485_, new_C6486_,
    new_C6487_, new_C6488_, new_C6489_, new_C6490_, new_C6491_, new_C6492_,
    new_C6493_, new_C6494_, new_C6495_, new_C6496_, new_C6497_, new_C6498_,
    new_C6499_, new_C6500_, new_C6501_, new_C6502_, new_C6503_, new_C6504_,
    new_C6505_, new_C6506_, new_C6507_, new_C6508_, new_C6509_, new_C6510_,
    new_C6511_, new_C6512_, new_C6513_, new_C6514_, new_C6515_, new_C6516_,
    new_C6517_, new_C6518_, new_C6519_, new_C6520_, new_C6521_, new_C6522_,
    new_C6523_, new_C6524_, new_C6525_, new_C6526_, new_C6527_, new_C6528_,
    new_C6529_, new_C6530_, new_C6531_, new_C6532_, new_C6533_, new_C6534_,
    new_C6535_, new_C6536_, new_C6537_, new_C6538_, new_C6539_, new_C6540_,
    new_C6541_, new_C6542_, new_C6543_, new_C6544_, new_C6545_, new_C6546_,
    new_C6547_, new_C6548_, new_C6549_, new_C6550_, new_C6551_, new_C6552_,
    new_C6553_, new_C6554_, new_C6555_, new_C6556_, new_C6557_, new_C6558_,
    new_C6559_, new_C6560_, new_C6561_, new_C6562_, new_C6563_, new_C6564_,
    new_C6565_, new_C6566_, new_C6567_, new_C6568_, new_C6569_, new_C6570_,
    new_C6571_, new_C6572_, new_C6573_, new_C6574_, new_C6575_, new_C6576_,
    new_C6577_, new_C6578_, new_C6579_, new_C6580_, new_C6581_, new_C6582_,
    new_C6583_, new_C6584_, new_C6585_, new_C6586_, new_C6587_, new_C6588_,
    new_C6589_, new_C6590_, new_C6591_, new_C6592_, new_C6593_, new_C6594_,
    new_C6595_, new_C6596_, new_C6597_, new_C6598_, new_C6599_, new_C6600_,
    new_C6601_, new_C6602_, new_C6603_, new_C6604_, new_C6605_, new_C6606_,
    new_C6607_, new_C6608_, new_C6609_, new_C6610_, new_C6611_, new_C6612_,
    new_C6613_, new_C6614_, new_C6615_, new_C6616_, new_C6617_, new_C6618_,
    new_C6619_, new_C6620_, new_C6621_, new_C6622_, new_C6623_, new_C6624_,
    new_C6625_, new_C6626_, new_C6627_, new_C6628_, new_C6629_, new_C6630_,
    new_C6631_, new_C6632_, new_C6633_, new_C6634_, new_C6635_, new_C6636_,
    new_C6637_, new_C6638_, new_C6639_, new_C6640_, new_C6641_, new_C6642_,
    new_C6643_, new_C6644_, new_C6645_, new_C6646_, new_C6647_, new_C6648_,
    new_C6649_, new_C6650_, new_C6651_, new_C6652_, new_C6653_, new_C6654_,
    new_C6655_, new_C6656_, new_C6657_, new_C6658_, new_C6659_, new_C6660_,
    new_C6661_, new_C6662_, new_C6663_, new_C6664_, new_C6665_, new_C6666_,
    new_C6667_, new_C6668_, new_C6669_, new_C6670_, new_C6671_, new_C6672_,
    new_C6673_, new_C6674_, new_C6675_, new_C6676_, new_C6677_, new_C6678_,
    new_C6679_, new_C6680_, new_C6681_, new_C6682_, new_C6683_, new_C6684_,
    new_C6685_, new_C6686_, new_C6687_, new_C6688_, new_C6689_, new_C6690_,
    new_C6691_, new_C6692_, new_C6693_, new_C6694_, new_C6695_, new_C6696_,
    new_C6697_, new_C6698_, new_C6699_, new_C6700_, new_C6701_, new_C6702_,
    new_C6703_, new_C6704_, new_C6705_, new_C6706_, new_C6707_, new_C6708_,
    new_C6709_, new_C6710_, new_C6711_, new_C6712_, new_C6713_, new_C6714_,
    new_C6715_, new_C6716_, new_C6717_, new_C6718_, new_C6719_, new_C6720_,
    new_C6721_, new_C6722_, new_C6723_, new_C6724_, new_C6725_, new_C6726_,
    new_C6727_, new_C6728_, new_C6729_, new_C6730_, new_C6731_, new_C6732_,
    new_C6733_, new_C6734_, new_C6735_, new_C6736_, new_C6737_, new_C6738_,
    new_C6739_, new_C6740_, new_C6741_, new_C6742_, new_C6743_, new_C6744_,
    new_C6745_, new_C6746_, new_C6747_, new_C6748_, new_C6749_, new_C6750_,
    new_C6751_, new_C6752_, new_C6753_, new_C6754_, new_C6755_, new_C6756_,
    new_C6757_, new_C6758_, new_C6759_, new_C6760_, new_C6761_, new_C6762_,
    new_C6763_, new_C6764_, new_C6765_, new_C6766_, new_C6767_, new_C6768_,
    new_C6769_, new_C6770_, new_C6771_, new_C6772_, new_C6773_, new_C6774_,
    new_C6775_, new_C6776_, new_C6777_, new_C6778_, new_C6779_, new_C6780_,
    new_C6781_, new_C6782_, new_C6783_, new_C6784_, new_C6785_, new_C6786_,
    new_C6787_, new_C6788_, new_C6789_, new_C6790_, new_C6791_, new_C6792_,
    new_C6793_, new_C6794_, new_C6795_, new_C6796_, new_C6797_, new_C6798_,
    new_C6799_, new_C6800_, new_C6801_, new_C6802_, new_C6803_, new_C6804_,
    new_C6805_, new_C6806_, new_C6807_, new_C6808_, new_C6809_, new_C6810_,
    new_C6811_, new_C6812_, new_C6813_, new_C6814_, new_C6815_, new_C6816_,
    new_C6817_, new_C6818_, new_C6819_, new_C6820_, new_C6821_, new_C6822_,
    new_C6823_, new_C6824_, new_C6825_, new_C6826_, new_C6827_, new_C6828_,
    new_C6829_, new_C6830_, new_C6831_, new_C6832_, new_C6833_, new_C6834_,
    new_C6835_, new_C6836_, new_C6837_, new_C6838_, new_C6839_, new_C6840_,
    new_C6841_, new_C6842_, new_C6843_, new_C6844_, new_C6845_, new_C6846_,
    new_C6847_, new_C6848_, new_C6849_, new_C6850_, new_C6851_, new_C6852_,
    new_C6853_, new_C6854_, new_C6855_, new_C6856_, new_C6857_, new_C6858_,
    new_C6859_, new_C6860_, new_C6861_, new_C6862_, new_C6863_, new_C6864_,
    new_C6865_, new_C6866_, new_C6867_, new_C6868_, new_C6869_, new_C6870_,
    new_C6871_, new_C6872_, new_C6873_, new_C6874_, new_C6875_, new_C6876_,
    new_C6877_, new_C6878_, new_C6879_, new_C6880_, new_C6881_, new_C6882_,
    new_C6883_, new_C6884_, new_C6885_, new_C6886_, new_C6887_, new_C6888_,
    new_C6889_, new_C6890_, new_C6891_, new_C6892_, new_C6893_, new_C6894_,
    new_C6895_, new_C6896_, new_C6897_, new_C6898_, new_C6899_, new_C6900_,
    new_C6901_, new_C6902_, new_C6903_, new_C6904_, new_C6905_, new_C6906_,
    new_C6907_, new_C6908_, new_C6909_, new_C6910_, new_C6911_, new_C6912_,
    new_C6913_, new_C6914_, new_C6915_, new_C6916_, new_C6917_, new_C6918_,
    new_C6919_, new_C6920_, new_C6921_, new_C6922_, new_C6923_, new_C6924_,
    new_C6925_, new_C6926_, new_C6927_, new_C6928_, new_C6929_, new_C6930_,
    new_C6931_, new_C6932_, new_C6933_, new_C6934_, new_C6935_, new_C6936_,
    new_C6937_, new_C6938_, new_C6939_, new_C6940_, new_C6941_, new_C6942_,
    new_C6943_, new_C6944_, new_C6945_, new_C6946_, new_C6947_, new_C6948_,
    new_C6949_, new_C6950_, new_C6951_, new_C6952_, new_C6953_, new_C6954_,
    new_C6955_, new_C6956_, new_C6957_, new_C6958_, new_C6959_, new_C6960_,
    new_C6961_, new_C6962_, new_C6963_, new_C6964_, new_C6965_, new_C6966_,
    new_C6967_, new_C6968_, new_C6969_, new_C6970_, new_C6971_, new_C6972_,
    new_C6973_, new_C6974_, new_C6975_, new_C6976_, new_C6977_, new_C6978_,
    new_C6979_, new_C6980_, new_C6981_, new_C6982_, new_C6983_, new_C6984_,
    new_C6985_, new_C6986_, new_C6987_, new_C6988_, new_C6989_, new_C6990_,
    new_C6991_, new_C6992_, new_C6993_, new_C6994_, new_C6995_, new_C6996_,
    new_C6997_, new_C6998_, new_C6999_, new_C7000_, new_C7001_, new_C7002_,
    new_C7003_, new_C7004_, new_C7005_, new_C7006_, new_C7007_, new_C7008_,
    new_C7009_, new_C7010_, new_C7011_, new_C7012_, new_C7013_, new_C7014_,
    new_C7015_, new_C7016_, new_C7017_, new_C7018_, new_C7019_, new_C7020_,
    new_C7021_, new_C7022_, new_C7023_, new_C7024_, new_C7025_, new_C7026_,
    new_C7027_, new_C7028_, new_C7029_, new_C7030_, new_C7031_, new_C7032_,
    new_C7033_, new_C7034_, new_C7035_, new_C7036_, new_C7037_, new_C7038_,
    new_C7039_, new_C7040_, new_C7041_, new_C7042_, new_C7043_, new_C7044_,
    new_C7045_, new_C7046_, new_C7047_, new_C7048_, new_C7049_, new_C7050_,
    new_C7051_, new_C7052_, new_C7053_, new_C7054_, new_C7055_, new_C7056_,
    new_C7057_, new_C7058_, new_C7059_, new_C7060_, new_C7061_, new_C7062_,
    new_C7063_, new_C7064_, new_C7065_, new_C7066_, new_C7067_, new_C7068_,
    new_C7069_, new_C7070_, new_C7071_, new_C7072_, new_C7073_, new_C7074_,
    new_C7075_, new_C7076_, new_C7077_, new_C7078_, new_C7079_, new_C7080_,
    new_C7081_, new_C7082_, new_C7083_, new_C7084_, new_C7085_, new_C7086_,
    new_C7087_, new_C7088_, new_C7089_, new_C7090_, new_C7091_, new_C7092_,
    new_C7093_, new_C7094_, new_C7095_, new_C7096_, new_C7097_, new_C7098_,
    new_C7099_, new_C7100_, new_C7101_, new_C7102_, new_C7103_, new_C7104_,
    new_C7105_, new_C7106_, new_C7107_, new_C7108_, new_C7109_, new_C7110_,
    new_C7111_, new_C7112_, new_C7113_, new_C7114_, new_C7115_, new_C7116_,
    new_C7117_, new_C7118_, new_C7119_, new_C7120_, new_C7121_, new_C7122_,
    new_C7123_, new_C7124_, new_C7125_, new_C7126_, new_C7127_, new_C7128_,
    new_C7129_, new_C7130_, new_C7131_, new_C7132_, new_C7133_, new_C7134_,
    new_C7135_, new_C7136_, new_C7137_, new_C7138_, new_C7139_, new_C7140_,
    new_C7141_, new_C7142_, new_C7143_, new_C7144_, new_C7145_, new_C7146_,
    new_C7147_, new_C7148_, new_C7149_, new_C7150_, new_C7151_, new_C7152_,
    new_C7153_, new_C7154_, new_C7155_, new_C7156_, new_C7157_, new_C7158_,
    new_C7159_, new_C7160_, new_C7161_, new_C7162_, new_C7163_, new_C7164_,
    new_C7165_, new_C7166_, new_C7167_, new_C7168_, new_C7169_, new_C7170_,
    new_C7171_, new_C7172_, new_C7173_, new_C7174_, new_C7175_, new_C7176_,
    new_C7177_, new_C7178_, new_C7179_, new_C7180_, new_C7181_, new_C7182_,
    new_C7183_, new_C7184_, new_C7185_, new_C7186_, new_C7187_, new_C7188_,
    new_C7189_, new_C7190_, new_C7191_, new_C7192_, new_C7193_, new_C7194_,
    new_C7195_, new_C7196_, new_C7197_, new_C7198_, new_C7199_, new_C7200_,
    new_C7201_, new_C7202_, new_C7203_, new_C7204_, new_C7205_, new_C7206_,
    new_C7207_, new_C7208_, new_C7209_, new_C7210_, new_C7211_, new_C7212_,
    new_C7213_, new_C7214_, new_C7215_, new_C7216_, new_C7217_, new_C7218_,
    new_C7219_, new_C7220_, new_C7221_, new_C7222_, new_C7223_, new_C7224_,
    new_C7225_, new_C7226_, new_C7227_, new_C7228_, new_C7229_, new_C7230_,
    new_C7231_, new_C7232_, new_C7233_, new_C7234_, new_C7235_, new_C7236_,
    new_C7237_, new_C7238_, new_C7239_, new_C7240_, new_C7241_, new_C7242_,
    new_C7243_, new_C7244_, new_C7245_, new_C7246_, new_C7247_, new_C7248_,
    new_C7249_, new_C7250_, new_C7251_, new_C7252_, new_C7253_, new_C7254_,
    new_C7255_, new_C7256_, new_C7257_, new_C7258_, new_C7259_, new_C7260_,
    new_C7261_, new_C7262_, new_C7263_, new_C7264_, new_C7265_, new_C7266_,
    new_C7267_, new_C7268_, new_C7269_, new_C7270_, new_C7271_, new_C7272_,
    new_C7273_, new_C7274_, new_C7275_, new_C7276_, new_C7277_, new_C7278_,
    new_C7279_, new_C7280_, new_C7281_, new_C7282_, new_C7283_, new_C7284_,
    new_C7285_, new_C7286_, new_C7287_, new_C7288_, new_C7289_, new_C7290_,
    new_C7291_, new_C7292_, new_C7293_, new_C7294_, new_C7295_, new_C7296_,
    new_C7297_, new_C7298_, new_C7299_, new_C7300_, new_C7301_, new_C7302_,
    new_C7303_, new_C7304_, new_C7305_, new_C7306_, new_C7307_, new_C7308_,
    new_C7309_, new_C7310_, new_C7311_, new_C7312_, new_C7313_, new_C7314_,
    new_C7315_, new_C7316_, new_C7317_, new_C7318_, new_C7319_, new_C7320_,
    new_C7321_, new_C7322_, new_C7323_, new_C7324_, new_C7325_, new_C7326_,
    new_C7327_, new_C7328_, new_C7329_, new_C7330_, new_C7331_, new_C7332_,
    new_C7333_, new_C7334_, new_C7335_, new_C7336_, new_C7337_, new_C7338_,
    new_C7339_, new_C7340_, new_C7341_, new_C7342_, new_C7343_, new_C7344_,
    new_C7345_, new_C7346_, new_C7347_, new_C7348_, new_C7349_, new_C7350_,
    new_C7351_, new_C7352_, new_C7353_, new_C7354_, new_C7355_, new_C7356_,
    new_C7357_, new_C7358_, new_C7359_, new_C7360_, new_C7361_, new_C7362_,
    new_C7363_, new_C7364_, new_C7365_, new_C7366_, new_C7367_, new_C7368_,
    new_C7369_, new_C7370_, new_C7371_, new_C7372_, new_C7373_, new_C7374_,
    new_C7375_, new_C7376_, new_C7377_, new_C7378_, new_C7379_, new_C7380_,
    new_C7381_, new_C7382_, new_C7383_, new_C7384_, new_C7385_, new_C7386_,
    new_C7387_, new_C7388_, new_C7389_, new_C7390_, new_C7391_, new_C7392_,
    new_C7393_, new_C7394_, new_C7395_, new_C7396_, new_C7397_, new_C7398_,
    new_C7399_, new_C7400_, new_C7401_, new_C7402_, new_C7403_, new_C7404_,
    new_C7405_, new_C7406_, new_C7407_, new_C7408_, new_C7409_, new_C7410_,
    new_C7411_, new_C7412_, new_C7413_, new_C7414_, new_C7415_, new_C7416_,
    new_C7417_, new_C7418_, new_C7419_, new_C7420_, new_C7421_, new_C7422_,
    new_C7423_, new_C7424_, new_C7425_, new_C7426_, new_C7427_, new_C7428_,
    new_C7429_, new_C7430_, new_C7431_, new_C7432_, new_C7433_, new_C7434_,
    new_C7435_, new_C7436_, new_C7437_, new_C7438_, new_C7439_, new_C7440_,
    new_C7441_, new_C7442_, new_C7443_, new_C7444_, new_C7445_, new_C7446_,
    new_C7447_, new_C7448_, new_C7449_, new_C7450_, new_C7451_, new_C7452_,
    new_C7453_, new_C7454_, new_C7455_, new_C7456_, new_C7457_, new_C7458_,
    new_C7459_, new_C7460_, new_C7461_, new_C7462_, new_C7463_, new_C7464_,
    new_C7465_, new_C7466_, new_C7467_, new_C7468_, new_C7469_, new_C7470_,
    new_C7471_, new_C7472_, new_C7473_, new_C7474_, new_C7475_, new_C7476_,
    new_C7477_, new_C7478_, new_C7479_, new_C7480_, new_C7481_, new_C7482_,
    new_C7483_, new_C7484_, new_C7485_, new_C7486_, new_C7487_, new_C7488_,
    new_C7489_, new_C7490_, new_C7491_, new_C7492_, new_C7493_, new_C7494_,
    new_C7495_, new_C7496_, new_C7497_, new_C7498_, new_C7499_, new_C7500_,
    new_C7501_, new_C7502_, new_C7503_, new_C7504_, new_C7505_, new_C7506_,
    new_C7507_, new_C7508_, new_C7509_, new_C7510_, new_C7511_, new_C7512_,
    new_C7513_, new_C7514_, new_C7515_, new_C7516_, new_C7517_, new_C7518_,
    new_C7519_, new_C7520_, new_C7521_, new_C7522_, new_C7523_, new_C7524_,
    new_C7525_, new_C7526_, new_C7527_, new_C7528_, new_C7529_, new_C7530_,
    new_C7531_, new_C7532_, new_C7533_, new_C7534_, new_C7535_, new_C7536_,
    new_C7537_, new_C7538_, new_C7539_, new_C7540_, new_C7541_, new_C7542_,
    new_C7543_, new_C7544_, new_C7545_, new_C7546_, new_C7547_, new_C7548_,
    new_C7549_, new_C7550_, new_C7551_, new_C7552_, new_C7553_, new_C7554_,
    new_C7555_, new_C7556_, new_C7557_, new_C7558_, new_C7559_, new_C7560_,
    new_C7561_, new_C7562_, new_C7563_, new_C7564_, new_C7565_, new_C7566_,
    new_C7567_, new_C7568_, new_C7569_, new_C7570_, new_C7571_, new_C7572_,
    new_C7573_, new_C7574_, new_C7575_, new_C7576_, new_C7577_, new_C7578_,
    new_C7579_, new_C7580_, new_C7581_, new_C7582_, new_C7583_, new_C7584_,
    new_C7585_, new_C7586_, new_C7587_, new_C7588_, new_C7589_, new_C7590_,
    new_C7591_, new_C7592_, new_C7593_, new_C7594_, new_C7595_, new_C7596_,
    new_C7597_, new_C7598_, new_C7599_, new_C7600_, new_C7601_, new_C7602_,
    new_C7603_, new_C7604_, new_C7605_, new_C7606_, new_C7607_, new_C7608_,
    new_C7609_, new_C7610_, new_C7611_, new_C7612_, new_C7613_, new_C7614_,
    new_C7615_, new_C7616_, new_C7617_, new_C7618_, new_C7619_, new_C7620_,
    new_C7621_, new_C7622_, new_C7623_, new_C7624_, new_C7625_, new_C7626_,
    new_C7627_, new_C7628_, new_C7629_, new_C7630_, new_C7631_, new_C7632_,
    new_C7633_, new_C7634_, new_C7635_, new_C7636_, new_C7637_, new_C7638_,
    new_C7639_, new_C7640_, new_C7641_, new_C7642_, new_C7643_, new_C7644_,
    new_C7645_, new_C7646_, new_C7647_, new_C7648_, new_C7649_, new_C7650_,
    new_C7651_, new_C7652_, new_C7653_, new_C7654_, new_C7655_, new_C7656_,
    new_C7657_, new_C7658_, new_C7659_, new_C7660_, new_C7661_, new_C7662_,
    new_C7663_, new_C7664_, new_C7665_, new_C7666_, new_C7667_, new_C7668_,
    new_C7669_, new_C7670_, new_C7671_, new_C7672_, new_C7673_, new_C7674_,
    new_C7675_, new_C7676_, new_C7677_, new_C7678_, new_C7679_, new_C7680_,
    new_C7681_, new_C7682_, new_C7683_, new_C7684_, new_C7685_, new_C7686_,
    new_C7687_, new_C7688_, new_C7689_, new_C7690_, new_C7691_, new_C7692_,
    new_C7693_, new_C7694_, new_C7695_, new_C7696_, new_C7697_, new_C7698_,
    new_C7699_, new_C7700_, new_C7701_, new_C7702_, new_C7703_, new_C7704_,
    new_C7705_, new_C7706_, new_C7707_, new_C7708_, new_C7709_, new_C7710_,
    new_C7711_, new_C7712_, new_C7713_, new_C7714_, new_C7715_, new_C7716_,
    new_C7717_, new_C7718_, new_C7719_, new_C7720_, new_C7721_, new_C7722_,
    new_C7723_, new_C7724_, new_C7725_, new_C7726_, new_C7727_, new_C7728_,
    new_C7729_, new_C7730_, new_C7731_, new_C7732_, new_C7733_, new_C7734_,
    new_C7735_, new_C7736_, new_C7737_, new_C7738_, new_C7739_, new_C7740_,
    new_C7741_, new_C7742_, new_C7743_, new_C7744_, new_C7745_, new_C7746_,
    new_C7747_, new_C7748_, new_C7749_, new_C7750_, new_C7751_, new_C7752_,
    new_C7753_, new_C7754_, new_C7755_, new_C7756_, new_C7757_, new_C7758_,
    new_C7759_, new_C7760_, new_C7761_, new_C7762_, new_C7763_, new_C7764_,
    new_C7765_, new_C7766_, new_C7767_, new_C7768_, new_C7769_, new_C7770_,
    new_C7771_, new_C7772_, new_C7773_, new_C7774_, new_C7775_, new_C7776_,
    new_C7777_, new_C7778_, new_C7779_, new_C7780_, new_C7781_, new_C7782_,
    new_C7783_, new_C7784_, new_C7785_, new_C7786_, new_C7787_, new_C7788_,
    new_C7789_, new_C7790_, new_C7791_, new_C7792_, new_C7793_, new_C7794_,
    new_C7795_, new_C7796_, new_C7797_, new_C7798_, new_C7799_, new_C7800_,
    new_C7801_, new_C7802_, new_C7803_, new_C7804_, new_C7805_, new_C7806_,
    new_C7807_, new_C7808_, new_C7809_, new_C7810_, new_C7811_, new_C7812_,
    new_C7813_, new_C7814_, new_C7815_, new_C7816_, new_C7817_, new_C7818_,
    new_C7819_, new_C7820_, new_C7821_, new_C7822_, new_C7823_, new_C7824_,
    new_C7825_, new_C7826_, new_C7827_, new_C7828_, new_C7829_, new_C7830_,
    new_C7831_, new_C7832_, new_C7833_, new_C7834_, new_C7835_, new_C7836_,
    new_C7837_, new_C7838_, new_C7839_, new_C7840_, new_C7841_, new_C7842_,
    new_C7843_, new_C7844_, new_C7845_, new_C7846_, new_C7847_, new_C7848_,
    new_C7849_, new_C7850_, new_C7851_, new_C7852_, new_C7853_, new_C7854_,
    new_C7855_, new_C7856_, new_C7857_, new_C7858_, new_C7859_, new_C7860_,
    new_C7861_, new_C7862_, new_C7863_, new_C7864_, new_C7865_, new_C7866_,
    new_C7867_, new_C7868_, new_C7869_, new_C7870_, new_C7871_, new_C7872_,
    new_C7873_, new_C7874_, new_C7875_, new_C7876_, new_C7877_, new_C7878_,
    new_C7879_, new_C7880_, new_C7881_, new_C7882_, new_C7883_, new_C7884_,
    new_C7885_, new_C7886_, new_C7887_, new_C7888_, new_C7889_, new_C7890_,
    new_C7891_, new_C7892_, new_C7893_, new_C7894_, new_C7895_, new_C7896_,
    new_C7897_, new_C7898_, new_C7899_, new_C7900_, new_C7901_, new_C7902_,
    new_C7903_, new_C7904_, new_C7905_, new_C7906_, new_C7907_, new_C7908_,
    new_C7909_, new_C7910_, new_C7911_, new_C7912_, new_C7913_, new_C7914_,
    new_C7915_, new_C7916_, new_C7917_, new_C7918_, new_C7919_, new_C7920_,
    new_C7921_, new_C7922_, new_C7923_, new_C7924_, new_C7925_, new_C7926_,
    new_C7927_, new_C7928_, new_C7929_, new_C7930_, new_C7931_, new_C7932_,
    new_C7933_, new_C7934_, new_C7935_, new_C7936_, new_C7937_, new_C7938_,
    new_C7939_, new_C7940_, new_C7941_, new_C7942_, new_C7943_, new_C7944_,
    new_C7945_, new_C7946_, new_C7947_, new_C7948_, new_C7949_, new_C7950_,
    new_C7951_, new_C7952_, new_C7953_, new_C7954_, new_C7955_, new_C7956_,
    new_C7957_, new_C7958_, new_C7959_, new_C7960_, new_C7961_, new_C7962_,
    new_C7963_, new_C7964_, new_C7965_, new_C7966_, new_C7967_, new_C7968_,
    new_C7969_, new_C7970_, new_C7971_, new_C7972_, new_C7973_, new_C7974_,
    new_C7975_, new_C7976_, new_C7977_, new_C7978_, new_C7979_, new_C7980_,
    new_C7981_, new_C7982_, new_C7983_, new_C7984_, new_C7985_, new_C7986_,
    new_C7987_, new_C7988_, new_C7989_, new_C7990_, new_C7991_, new_C7992_,
    new_C7993_, new_C7994_, new_C7995_, new_C7996_, new_C7997_, new_C7998_,
    new_C7999_, new_C8000_, new_C8001_, new_C8002_, new_C8003_, new_C8004_,
    new_C8005_, new_C8006_, new_C8007_, new_C8008_, new_C8009_, new_C8010_,
    new_C8011_, new_C8012_, new_C8013_, new_C8014_, new_C8015_, new_C8016_,
    new_C8017_, new_C8018_, new_C8019_, new_C8020_, new_C8021_, new_C8022_,
    new_C8023_, new_C8024_, new_C8025_, new_C8026_, new_C8027_, new_C8028_,
    new_C8029_, new_C8030_, new_C8031_, new_C8032_, new_C8033_, new_C8034_,
    new_C8035_, new_C8036_, new_C8037_, new_C8038_, new_C8039_, new_C8040_,
    new_C8041_, new_C8042_, new_C8043_, new_C8044_, new_C8045_, new_C8046_,
    new_C8047_, new_C8048_, new_C8049_, new_C8050_, new_C8051_, new_C8052_,
    new_C8053_, new_C8054_, new_C8055_, new_C8056_, new_C8057_, new_C8058_,
    new_C8059_, new_C8060_, new_C8061_, new_C8062_, new_C8063_, new_C8064_,
    new_C8065_, new_C8066_, new_C8067_, new_C8068_, new_C8069_, new_C8070_,
    new_C8071_, new_C8072_, new_C8073_, new_C8074_, new_C8075_, new_C8076_,
    new_C8077_, new_C8078_, new_C8079_, new_C8080_, new_C8081_, new_C8082_,
    new_C8083_, new_C8084_, new_C8085_, new_C8086_, new_C8087_, new_C8088_,
    new_C8089_, new_C8090_, new_C8091_, new_C8092_, new_C8093_, new_C8094_,
    new_C8095_, new_C8096_, new_C8097_, new_C8098_, new_C8099_, new_C8100_,
    new_C8101_, new_C8102_, new_C8103_, new_C8104_, new_C8105_, new_C8106_,
    new_C8107_, new_C8108_, new_C8109_, new_C8110_, new_C8111_, new_C8112_,
    new_C8113_, new_C8114_, new_C8115_, new_C8116_, new_C8117_, new_C8118_,
    new_C8119_, new_C8120_, new_C8121_, new_C8122_, new_C8123_, new_C8124_,
    new_C8125_, new_C8126_, new_C8127_, new_C8128_, new_C8129_, new_C8130_,
    new_C8131_, new_C8132_, new_C8133_, new_C8134_, new_C8135_, new_C8136_,
    new_C8137_, new_C8138_, new_C8139_, new_C8140_, new_C8141_, new_C8142_,
    new_C8143_, new_C8144_, new_C8145_, new_C8146_, new_C8147_, new_C8148_,
    new_C8149_, new_C8150_, new_C8151_, new_C8152_, new_C8153_, new_C8154_,
    new_C8155_, new_C8156_, new_C8157_, new_C8158_, new_C8159_, new_C8160_,
    new_C8161_, new_C8162_, new_C8163_, new_C8164_, new_C8165_, new_C8166_,
    new_C8167_, new_C8168_, new_C8169_, new_C8170_, new_C8171_, new_C8172_,
    new_C8173_, new_C8174_, new_C8175_, new_C8176_, new_C8177_, new_C8178_,
    new_C8179_, new_C8180_, new_C8181_, new_C8182_, new_C8183_, new_C8184_,
    new_C8185_, new_C8186_, new_C8187_, new_C8188_, new_C8189_, new_C8190_,
    new_C8191_, new_C8192_, new_C8193_, new_C8194_, new_C8195_, new_C8196_,
    new_C8197_, new_C8198_, new_C8199_, new_C8200_, new_C8201_, new_C8202_,
    new_C8203_, new_C8204_, new_C8205_, new_C8206_, new_C8207_, new_C8208_,
    new_C8209_, new_C8210_, new_C8211_, new_C8212_, new_C8213_, new_C8214_,
    new_C8215_, new_C8216_, new_C8217_, new_C8218_, new_C8219_, new_C8220_,
    new_C8221_, new_C8222_, new_C8223_, new_C8224_, new_C8225_, new_C8226_,
    new_C8227_, new_C8228_, new_C8229_, new_C8230_, new_C8231_, new_C8232_,
    new_C8233_, new_C8234_, new_C8235_, new_C8236_, new_C8237_, new_C8238_,
    new_C8239_, new_C8240_, new_C8241_, new_C8242_, new_C8243_, new_C8244_,
    new_C8245_, new_C8246_, new_C8247_, new_C8248_, new_C8249_, new_C8250_,
    new_C8251_, new_C8252_, new_C8253_, new_C8254_, new_C8255_, new_C8256_,
    new_C8257_, new_C8258_, new_C8259_, new_C8260_, new_C8261_, new_C8262_,
    new_C8263_, new_C8264_, new_C8265_, new_C8266_, new_C8267_, new_C8268_,
    new_C8269_, new_C8270_, new_C8271_, new_C8272_, new_C8273_, new_C8274_,
    new_C8275_, new_C8276_, new_C8277_, new_C8278_, new_C8279_, new_C8280_,
    new_C8281_, new_C8282_, new_C8283_, new_C8284_, new_C8285_, new_C8286_,
    new_C8287_, new_C8288_, new_C8289_, new_C8290_, new_C8291_, new_C8292_,
    new_C8293_, new_C8294_, new_C8295_, new_C8296_, new_C8297_, new_C8298_,
    new_C8299_, new_C8300_, new_C8301_, new_C8302_, new_C8303_, new_C8304_,
    new_C8305_, new_C8306_, new_C8307_, new_C8308_, new_C8309_, new_C8310_,
    new_C8311_, new_C8312_, new_C8313_, new_C8314_, new_C8315_, new_C8316_,
    new_C8317_, new_C8318_, new_C8319_, new_C8320_, new_C8321_, new_C8322_,
    new_C8323_, new_C8324_, new_C8325_, new_C8326_, new_C8327_, new_C8328_,
    new_C8329_, new_C8330_, new_C8331_, new_C8332_, new_C8333_, new_C8334_,
    new_C8335_, new_C8336_, new_C8337_, new_C8338_, new_C8339_, new_C8340_,
    new_C8341_, new_C8342_, new_C8343_, new_C8344_, new_C8345_, new_C8346_,
    new_C8347_, new_C8348_, new_C8349_, new_C8350_, new_C8351_, new_C8352_,
    new_C8353_, new_C8354_, new_C8355_, new_C8356_, new_C8357_, new_C8358_,
    new_C8359_, new_C8360_, new_C8361_, new_C8362_, new_C8363_, new_C8364_,
    new_C8365_, new_C8366_, new_C8367_, new_C8368_, new_C8369_, new_C8370_,
    new_C8371_, new_C8372_, new_C8373_, new_C8374_, new_C8375_, new_C8376_,
    new_C8377_, new_C8378_, new_C8379_, new_C8380_, new_C8381_, new_C8382_,
    new_C8383_, new_C8384_, new_C8385_, new_C8386_, new_C8387_, new_C8388_,
    new_C8389_, new_C8390_, new_C8391_, new_C8392_, new_C8393_, new_C8394_,
    new_C8395_, new_C8396_, new_C8397_, new_C8398_, new_C8399_, new_C8400_,
    new_C8401_, new_C8402_, new_C8403_, new_C8404_, new_C8405_, new_C8406_,
    new_C8407_, new_C8408_, new_C8409_, new_C8410_, new_C8411_, new_C8412_,
    new_C8413_, new_C8414_, new_C8415_, new_C8416_, new_C8417_, new_C8418_,
    new_C8419_, new_C8420_, new_C8421_, new_C8422_, new_C8423_, new_C8424_,
    new_C8425_, new_C8426_, new_C8427_, new_C8428_, new_C8429_, new_C8430_,
    new_C8431_, new_C8432_, new_C8433_, new_C8434_, new_C8435_, new_C8436_,
    new_C8437_, new_C8438_, new_C8439_, new_C8440_, new_C8441_, new_C8442_,
    new_C8443_, new_C8444_, new_C8445_, new_C8446_, new_C8447_, new_C8448_,
    new_C8449_, new_C8450_, new_C8451_, new_C8452_, new_C8453_, new_C8454_,
    new_C8455_, new_C8456_, new_C8457_, new_C8458_, new_C8459_, new_C8460_,
    new_C8461_, new_C8462_, new_C8463_, new_C8464_, new_C8465_, new_C8466_,
    new_C8467_, new_C8468_, new_C8469_, new_C8470_, new_C8471_, new_C8472_,
    new_C8473_, new_C8474_, new_C8475_, new_C8476_, new_C8477_, new_C8478_,
    new_C8479_, new_C8480_, new_C8481_, new_C8482_, new_C8483_, new_C8484_,
    new_C8485_, new_C8486_, new_C8487_, new_C8488_, new_C8489_, new_C8490_,
    new_C8491_, new_C8492_, new_C8493_, new_C8494_, new_C8495_, new_C8496_,
    new_C8497_, new_C8498_, new_C8499_, new_C8500_, new_C8501_, new_C8502_,
    new_C8503_, new_C8504_, new_C8505_, new_C8506_, new_C8507_, new_C8508_,
    new_C8509_, new_C8510_, new_C8511_, new_C8512_, new_C8513_, new_C8514_,
    new_C8515_, new_C8516_, new_C8517_, new_C8518_, new_C8519_, new_C8520_,
    new_C8521_, new_C8522_, new_C8523_, new_C8524_, new_C8525_, new_C8526_,
    new_C8527_, new_C8528_, new_C8529_, new_C8530_, new_C8531_, new_C8532_,
    new_C8533_, new_C8534_, new_C8535_, new_C8536_, new_C8537_, new_C8538_,
    new_C8539_, new_C8540_, new_C8541_, new_C8542_, new_C8543_, new_C8544_,
    new_C8545_, new_C8546_, new_C8547_, new_C8548_, new_C8549_, new_C8550_,
    new_C8551_, new_C8552_, new_C8553_, new_C8554_, new_C8555_, new_C8556_,
    new_C8557_, new_C8558_, new_C8559_, new_C8560_, new_C8561_, new_C8562_,
    new_C8563_, new_C8564_, new_C8565_, new_C8566_, new_C8567_, new_C8568_,
    new_C8569_, new_C8570_, new_C8571_, new_C8572_, new_C8573_, new_C8574_,
    new_C8575_, new_C8576_, new_C8577_, new_C8578_, new_C8579_, new_C8580_,
    new_C8581_, new_C8582_, new_C8583_, new_C8584_, new_C8585_, new_C8586_,
    new_C8587_, new_C8588_, new_C8589_, new_C8590_, new_C8591_, new_C8592_,
    new_C8593_, new_C8594_, new_C8595_, new_C8596_, new_C8597_, new_C8598_,
    new_C8599_, new_C8600_, new_C8601_, new_C8602_, new_C8603_, new_C8604_,
    new_C8605_, new_C8606_, new_C8607_, new_C8608_, new_C8609_, new_C8610_,
    new_C8611_, new_C8612_, new_C8613_, new_C8614_, new_C8615_, new_C8616_,
    new_C8617_, new_C8618_, new_C8619_, new_C8620_, new_C8621_, new_C8622_,
    new_C8623_, new_C8624_, new_C8625_, new_C8626_, new_C8627_, new_C8628_,
    new_C8629_, new_C8630_, new_C8631_, new_C8632_, new_C8633_, new_C8634_,
    new_C8635_, new_C8636_, new_C8637_, new_C8638_, new_C8639_, new_C8640_,
    new_C8641_, new_C8642_, new_C8643_, new_C8644_, new_C8645_, new_C8646_,
    new_C8647_, new_C8648_, new_C8649_, new_C8650_, new_C8651_, new_C8652_,
    new_C8653_, new_C8654_, new_C8655_, new_C8656_, new_C8657_, new_C8658_,
    new_C8659_, new_C8660_, new_C8661_, new_C8662_, new_C8663_, new_C8664_,
    new_C8665_, new_C8666_, new_C8667_, new_C8668_, new_C8669_, new_C8670_,
    new_C8671_, new_C8672_, new_C8673_, new_C8674_, new_C8675_, new_C8676_,
    new_C8677_, new_C8678_, new_C8679_, new_C8680_, new_C8681_, new_C8682_,
    new_C8683_, new_C8684_, new_C8685_, new_C8686_, new_C8687_, new_C8688_,
    new_C8689_, new_C8690_, new_C8691_, new_C8692_, new_C8693_, new_C8694_,
    new_C8695_, new_C8696_, new_C8697_, new_C8698_, new_C8699_, new_C8700_,
    new_C8701_, new_C8702_, new_C8703_, new_C8704_, new_C8705_, new_C8706_,
    new_C8707_, new_C8708_, new_C8709_, new_C8710_, new_C8711_, new_C8712_,
    new_C8713_, new_C8714_, new_C8715_, new_C8716_, new_C8717_, new_C8718_,
    new_C8719_, new_C8720_, new_C8721_, new_C8722_, new_C8723_, new_C8724_,
    new_C8725_, new_C8726_, new_C8727_, new_C8728_, new_C8729_, new_C8730_,
    new_C8731_, new_C8732_, new_C8733_, new_C8734_, new_C8735_, new_C8736_,
    new_C8737_, new_C8738_, new_C8739_, new_C8740_, new_C8741_, new_C8742_,
    new_C8743_, new_C8744_, new_C8745_, new_C8746_, new_C8747_, new_C8748_,
    new_C8749_, new_C8750_, new_C8751_, new_C8752_, new_C8753_, new_C8754_,
    new_C8755_, new_C8756_, new_C8757_, new_C8758_, new_C8759_, new_C8760_,
    new_C8761_, new_C8762_, new_C8763_, new_C8764_, new_C8765_, new_C8766_,
    new_C8767_, new_C8768_, new_C8769_, new_C8770_, new_C8771_, new_C8772_,
    new_C8773_, new_C8774_, new_C8775_, new_C8776_, new_C8777_, new_C8778_,
    new_C8779_, new_C8780_, new_C8781_, new_C8782_, new_C8783_, new_C8784_,
    new_C8785_, new_C8786_, new_C8787_, new_C8788_, new_C8789_, new_C8790_,
    new_C8791_, new_C8792_, new_C8793_, new_C8794_, new_C8795_, new_C8796_,
    new_C8797_, new_C8798_, new_C8799_, new_C8800_, new_C8801_, new_C8802_,
    new_C8803_, new_C8804_, new_C8805_, new_C8806_, new_C8807_, new_C8808_,
    new_C8809_, new_C8810_, new_C8811_, new_C8812_, new_C8813_, new_C8814_,
    new_C8815_, new_C8816_, new_C8817_, new_C8818_, new_C8819_, new_C8820_,
    new_C8821_, new_C8822_, new_C8823_, new_C8824_, new_C8825_, new_C8826_,
    new_C8827_, new_C8828_, new_C8829_, new_C8830_, new_C8831_, new_C8832_,
    new_C8833_, new_C8834_, new_C8835_, new_C8836_, new_C8837_, new_C8838_,
    new_C8839_, new_C8840_, new_C8841_, new_C8842_, new_C8843_, new_C8844_,
    new_C8845_, new_C8846_, new_C8847_, new_C8848_, new_C8849_, new_C8850_,
    new_C8851_, new_C8852_, new_C8853_, new_C8854_, new_C8855_, new_C8856_,
    new_C8857_, new_C8858_, new_C8859_, new_C8860_, new_C8861_, new_C8862_,
    new_C8863_, new_C8864_, new_C8865_, new_C8866_, new_C8867_, new_C8868_,
    new_C8869_, new_C8870_, new_C8871_, new_C8872_, new_C8873_, new_C8874_,
    new_C8875_, new_C8876_, new_C8877_, new_C8878_, new_C8879_, new_C8880_,
    new_C8881_, new_C8882_, new_C8883_, new_C8884_, new_C8885_, new_C8886_,
    new_C8887_, new_C8888_, new_C8889_, new_C8890_, new_C8891_, new_C8892_,
    new_C8893_, new_C8894_, new_C8895_, new_C8896_, new_C8897_, new_C8898_,
    new_C8899_, new_C8900_, new_C8901_, new_C8902_, new_C8903_, new_C8904_,
    new_C8905_, new_C8906_, new_C8907_, new_C8908_, new_C8909_, new_C8910_,
    new_C8911_, new_C8912_, new_C8913_, new_C8914_, new_C8915_, new_C8916_,
    new_C8917_, new_C8918_, new_C8919_, new_C8920_, new_C8921_, new_C8922_,
    new_C8923_, new_C8924_, new_C8925_, new_C8926_, new_C8927_, new_C8928_,
    new_C8929_, new_C8930_, new_C8931_, new_C8932_, new_C8933_, new_C8934_,
    new_C8935_, new_C8936_, new_C8937_, new_C8938_, new_C8939_, new_C8940_,
    new_C8941_, new_C8942_, new_C8943_, new_C8944_, new_C8945_, new_C8946_,
    new_C8947_, new_C8948_, new_C8949_, new_C8950_, new_C8951_, new_C8952_,
    new_C8953_, new_C8954_, new_C8955_, new_C8956_, new_C8957_, new_C8958_,
    new_C8959_, new_C8960_, new_C8961_, new_C8962_, new_C8963_, new_C8964_,
    new_C8965_, new_C8966_, new_C8967_, new_C8968_, new_C8969_, new_C8970_,
    new_C8971_, new_C8972_, new_C8973_, new_C8974_, new_C8975_, new_C8976_,
    new_C8977_, new_C8978_, new_C8979_, new_C8980_, new_C8981_, new_C8982_,
    new_C8983_, new_C8984_, new_C8985_, new_C8986_, new_C8987_, new_C8988_,
    new_C8989_, new_C8990_, new_C8991_, new_C8992_, new_C8993_, new_C8994_,
    new_C8995_, new_C8996_, new_C8997_, new_C8998_, new_C8999_, new_C9000_,
    new_C9001_, new_C9002_, new_C9003_, new_C9004_, new_C9005_, new_C9006_,
    new_C9007_, new_C9008_, new_C9009_, new_C9010_, new_C9011_, new_C9012_,
    new_C9013_, new_C9014_, new_C9015_, new_C9016_, new_C9017_, new_C9018_,
    new_C9019_, new_C9020_, new_C9021_, new_C9022_, new_C9023_, new_C9024_,
    new_C9025_, new_C9026_, new_C9027_, new_C9028_, new_C9029_, new_C9030_,
    new_C9031_, new_C9032_, new_C9033_, new_C9034_, new_C9035_, new_C9036_,
    new_C9037_, new_C9038_, new_C9039_, new_C9040_, new_C9041_, new_C9042_,
    new_C9043_, new_C9044_, new_C9045_, new_C9046_, new_C9047_, new_C9048_,
    new_C9049_, new_C9050_, new_C9051_, new_C9052_, new_C9053_, new_C9054_,
    new_C9055_, new_C9056_, new_C9057_, new_C9058_, new_C9059_, new_C9060_,
    new_C9061_, new_C9062_, new_C9063_, new_C9064_, new_C9065_, new_C9066_,
    new_C9067_, new_C9068_, new_C9069_, new_C9070_, new_C9071_, new_C9072_,
    new_C9073_, new_C9074_, new_C9075_, new_C9076_, new_C9077_, new_C9078_,
    new_C9079_, new_C9080_, new_C9081_, new_C9082_, new_C9083_, new_C9084_,
    new_C9085_, new_C9086_, new_C9087_, new_C9088_, new_C9089_, new_C9090_,
    new_C9091_, new_C9092_, new_C9093_, new_C9094_, new_C9095_, new_C9096_,
    new_C9097_, new_C9098_, new_C9099_, new_C9100_, new_C9101_, new_C9102_,
    new_C9103_, new_C9104_, new_C9105_, new_C9106_, new_C9107_, new_C9108_,
    new_C9109_, new_C9110_, new_C9111_, new_C9112_, new_C9113_, new_C9114_,
    new_C9115_, new_C9116_, new_C9117_, new_C9118_, new_C9119_, new_C9120_,
    new_C9121_, new_C9122_, new_C9123_, new_C9124_, new_C9125_, new_C9126_,
    new_C9127_, new_C9128_, new_C9129_, new_C9130_, new_C9131_, new_C9132_,
    new_C9133_, new_C9134_, new_C9135_, new_C9136_, new_C9137_, new_C9138_,
    new_C9139_, new_C9140_, new_C9141_, new_C9142_, new_C9143_, new_C9144_,
    new_C9145_, new_C9146_, new_C9147_, new_C9148_, new_C9149_, new_C9150_,
    new_C9151_, new_C9152_, new_C9153_, new_C9154_, new_C9155_, new_C9156_,
    new_C9157_, new_C9158_, new_C9159_, new_C9160_, new_C9161_, new_C9162_,
    new_C9163_, new_C9164_, new_C9165_, new_C9166_, new_C9167_, new_C9168_,
    new_C9169_, new_C9170_, new_C9171_, new_C9172_, new_C9173_, new_C9174_,
    new_C9175_, new_C9176_, new_C9177_, new_C9178_, new_C9179_, new_C9180_,
    new_C9181_, new_C9182_, new_C9183_, new_C9184_, new_C9185_, new_C9186_,
    new_C9187_, new_C9188_, new_C9189_, new_C9190_, new_C9191_, new_C9192_,
    new_C9193_, new_C9194_, new_C9195_, new_C9196_, new_C9197_, new_C9198_,
    new_C9199_, new_C9200_, new_C9201_, new_C9202_, new_C9203_, new_C9204_,
    new_C9205_, new_C9206_, new_C9207_, new_C9208_, new_C9209_, new_C9210_,
    new_C9211_, new_C9212_, new_C9213_, new_C9214_, new_C9215_, new_C9216_,
    new_C9217_, new_C9218_, new_C9219_, new_C9220_, new_C9221_, new_C9222_,
    new_C9223_, new_C9224_, new_C9225_, new_C9226_, new_C9227_, new_C9228_,
    new_C9229_, new_C9230_, new_C9231_, new_C9232_, new_C9233_, new_C9234_,
    new_C9235_, new_C9236_, new_C9237_, new_C9238_, new_C9239_, new_C9240_,
    new_C9241_, new_C9242_, new_C9243_, new_C9244_, new_C9245_, new_C9246_,
    new_C9247_, new_C9248_, new_C9249_, new_C9250_, new_C9251_, new_C9252_,
    new_C9253_, new_C9254_, new_C9255_, new_C9256_, new_C9257_, new_C9258_,
    new_C9259_, new_C9260_, new_C9261_, new_C9262_, new_C9263_, new_C9264_,
    new_C9265_, new_C9266_, new_C9267_, new_C9268_, new_C9269_, new_C9270_,
    new_C9271_, new_C9272_, new_C9273_, new_C9274_, new_C9275_, new_C9276_,
    new_C9277_, new_C9278_, new_C9279_, new_C9280_, new_C9281_, new_C9282_,
    new_C9283_, new_C9284_, new_C9285_, new_C9286_, new_C9287_, new_C9288_,
    new_C9289_, new_C9290_, new_C9291_, new_C9292_, new_C9293_, new_C9294_,
    new_C9295_, new_C9296_, new_C9297_, new_C9298_, new_C9299_, new_C9300_,
    new_C9301_, new_C9302_, new_C9303_, new_C9304_, new_C9305_, new_C9306_,
    new_C9307_, new_C9308_, new_C9309_, new_C9310_, new_C9311_, new_C9312_,
    new_C9313_, new_C9314_, new_C9315_, new_C9316_, new_C9317_, new_C9318_,
    new_C9319_, new_C9320_, new_C9321_, new_C9322_, new_C9323_, new_C9324_,
    new_C9325_, new_C9326_, new_C9327_, new_C9328_, new_C9329_, new_C9330_,
    new_C9331_, new_C9332_, new_C9333_, new_C9334_, new_C9335_, new_C9336_,
    new_C9337_, new_C9338_, new_C9339_, new_C9340_, new_C9341_, new_C9342_,
    new_C9343_, new_C9344_, new_C9345_, new_C9346_, new_C9347_, new_C9348_,
    new_C9349_, new_C9350_, new_C9351_, new_C9352_, new_C9353_, new_C9354_,
    new_C9355_, new_C9356_, new_C9357_, new_C9358_, new_C9359_, new_C9360_,
    new_C9361_, new_C9362_, new_C9363_, new_C9364_, new_C9365_, new_C9366_,
    new_C9367_, new_C9368_, new_C9369_, new_C9370_, new_C9371_, new_C9372_,
    new_C9373_, new_C9374_, new_C9375_, new_C9376_, new_C9377_, new_C9378_,
    new_C9379_, new_C9380_, new_C9381_, new_C9382_, new_C9383_, new_C9384_,
    new_C9385_, new_C9386_, new_C9387_, new_C9388_, new_C9389_, new_C9390_,
    new_C9391_, new_C9392_, new_C9393_, new_C9394_, new_C9395_, new_C9396_,
    new_C9397_, new_C9398_, new_C9399_, new_C9400_, new_C9401_, new_C9402_,
    new_C9403_, new_C9404_, new_C9405_, new_C9406_, new_C9407_, new_C9408_,
    new_C9409_, new_C9410_, new_C9411_, new_C9412_, new_C9413_, new_C9414_,
    new_C9415_, new_C9416_, new_C9417_, new_C9418_, new_C9419_, new_C9420_,
    new_C9421_, new_C9422_, new_C9423_, new_C9424_, new_C9425_, new_C9426_,
    new_C9427_, new_C9428_, new_C9429_, new_C9430_, new_C9431_, new_C9432_,
    new_C9433_, new_C9434_, new_C9435_, new_C9436_, new_C9437_, new_C9438_,
    new_C9439_, new_C9440_, new_C9441_, new_C9442_, new_C9443_, new_C9444_,
    new_C9445_, new_C9446_, new_C9447_, new_C9448_, new_C9449_, new_C9450_,
    new_C9451_, new_C9452_, new_C9453_, new_C9454_, new_C9455_, new_C9456_,
    new_C9457_, new_C9458_, new_C9459_, new_C9460_, new_C9461_, new_C9462_,
    new_C9463_, new_C9464_, new_C9465_, new_C9466_, new_C9467_, new_C9468_,
    new_C9469_, new_C9470_, new_C9471_, new_C9472_, new_C9473_, new_C9474_,
    new_C9475_, new_C9476_, new_C9477_, new_C9478_, new_C9479_, new_C9480_,
    new_C9481_, new_C9482_, new_C9483_, new_C9484_, new_C9485_, new_C9486_,
    new_C9487_, new_C9488_, new_C9489_, new_C9490_, new_C9491_, new_C9492_,
    new_C9493_, new_C9494_, new_C9495_, new_C9496_, new_C9497_, new_C9498_,
    new_C9499_, new_C9500_, new_C9501_, new_C9502_, new_C9503_, new_C9504_,
    new_C9505_, new_C9506_, new_C9507_, new_C9508_, new_C9509_, new_C9510_,
    new_C9511_, new_C9512_, new_C9513_, new_C9514_, new_C9515_, new_C9516_,
    new_C9517_, new_C9518_, new_C9519_, new_C9520_, new_C9521_, new_C9522_,
    new_C9523_, new_C9524_, new_C9525_, new_C9526_, new_C9527_, new_C9528_,
    new_C9529_, new_C9530_, new_C9531_, new_C9532_, new_C9533_, new_C9534_,
    new_C9535_, new_C9536_, new_C9537_, new_C9538_, new_C9539_, new_C9540_,
    new_C9541_, new_C9542_, new_C9543_, new_C9544_, new_C9545_, new_C9546_,
    new_C9547_, new_C9548_, new_C9549_, new_C9550_, new_C9551_, new_C9552_,
    new_C9553_, new_C9554_, new_C9555_, new_C9556_, new_C9557_, new_C9558_,
    new_C9559_, new_C9560_, new_C9561_, new_C9562_, new_C9563_, new_C9564_,
    new_C9565_, new_C9566_, new_C9567_, new_C9568_, new_C9569_, new_C9570_,
    new_C9571_, new_C9572_, new_C9573_, new_C9574_, new_C9575_, new_C9576_,
    new_C9577_, new_C9578_, new_C9579_, new_C9580_, new_C9581_, new_C9582_,
    new_C9583_, new_C9584_, new_C9585_, new_C9586_, new_C9587_, new_C9588_,
    new_C9589_, new_C9590_, new_C9591_, new_C9592_, new_C9593_, new_C9594_,
    new_C9595_, new_C9596_, new_C9597_, new_C9598_, new_C9599_, new_C9600_,
    new_C9601_, new_C9602_, new_C9603_, new_C9604_, new_C9605_, new_C9606_,
    new_C9607_, new_C9608_, new_C9609_, new_C9610_, new_C9611_, new_C9612_,
    new_C9613_, new_C9614_, new_C9615_, new_C9616_, new_C9617_, new_C9618_,
    new_C9619_, new_C9620_, new_C9621_, new_C9622_, new_C9623_, new_C9624_,
    new_C9625_, new_C9626_, new_C9627_, new_C9628_, new_C9629_, new_C9630_,
    new_C9631_, new_C9632_, new_C9633_, new_C9634_, new_C9635_, new_C9636_,
    new_C9637_, new_C9638_, new_C9639_, new_C9640_, new_C9641_, new_C9642_,
    new_C9643_, new_C9644_, new_C9645_, new_C9646_, new_C9647_, new_C9648_,
    new_C9649_, new_C9650_, new_C9651_, new_C9652_, new_C9653_, new_C9654_,
    new_C9655_, new_C9656_, new_C9657_, new_C9658_, new_C9659_, new_C9660_,
    new_C9661_, new_C9662_, new_C9663_, new_C9664_, new_C9665_, new_C9666_,
    new_C9667_, new_C9668_, new_C9669_, new_C9670_, new_C9671_, new_C9672_,
    new_C9673_, new_C9674_, new_C9675_, new_C9676_, new_C9677_, new_C9678_,
    new_C9679_, new_C9680_, new_C9681_, new_C9682_, new_C9683_, new_C9684_,
    new_C9685_, new_C9686_, new_C9687_, new_C9688_, new_C9689_, new_C9690_,
    new_C9691_, new_C9692_, new_C9693_, new_C9694_, new_C9695_, new_C9696_,
    new_C9697_, new_C9698_, new_C9699_, new_C9700_, new_C9701_, new_C9702_,
    new_C9703_, new_C9704_, new_C9705_, new_C9706_, new_C9707_, new_C9708_,
    new_C9709_, new_C9710_, new_C9711_, new_C9712_, new_C9713_, new_C9714_,
    new_C9715_, new_C9716_, new_C9717_, new_C9718_, new_C9719_, new_C9720_,
    new_C9721_, new_C9722_, new_C9723_, new_C9724_, new_C9725_, new_C9726_,
    new_C9727_, new_C9728_, new_C9729_, new_C9730_, new_C9731_, new_C9732_,
    new_C9733_, new_C9734_, new_C9735_, new_C9736_, new_C9737_, new_C9738_,
    new_C9739_, new_C9740_, new_C9741_, new_C9742_, new_C9743_, new_C9744_,
    new_C9745_, new_C9746_, new_C9747_, new_C9748_, new_C9749_, new_C9750_,
    new_C9751_, new_C9752_, new_C9753_, new_C9754_, new_C9755_, new_C9756_,
    new_C9757_, new_C9758_, new_C9759_, new_C9760_, new_C9761_, new_C9762_,
    new_C9763_, new_C9764_, new_C9765_, new_C9766_, new_C9767_, new_C9768_,
    new_C9769_, new_C9770_, new_C9771_, new_C9772_, new_C9773_, new_C9774_,
    new_C9775_, new_C9776_, new_C9777_, new_C9778_, new_C9779_, new_C9780_,
    new_C9781_, new_C9782_, new_C9783_, new_C9784_, new_C9785_, new_C9786_,
    new_C9787_, new_C9788_, new_C9789_, new_C9790_, new_C9791_, new_C9792_,
    new_C9793_, new_C9794_, new_C9795_, new_C9796_, new_C9797_, new_C9798_,
    new_C9799_, new_C9800_, new_C9801_, new_C9802_, new_C9803_, new_C9804_,
    new_C9805_, new_C9806_, new_C9807_, new_C9808_, new_C9809_, new_C9810_,
    new_C9811_, new_C9812_, new_C9813_, new_C9814_, new_C9815_, new_C9816_,
    new_C9817_, new_C9818_, new_C9819_, new_C9820_, new_C9821_, new_C9822_,
    new_C9823_, new_C9824_, new_C9825_, new_C9826_, new_C9827_, new_C9828_,
    new_C9829_, new_C9830_, new_C9831_, new_C9832_, new_C9833_, new_C9834_,
    new_C9835_, new_C9836_, new_C9837_, new_C9838_, new_C9839_, new_C9840_,
    new_C9841_, new_C9842_, new_C9843_, new_C9844_, new_C9845_, new_C9846_,
    new_C9847_, new_C9848_, new_C9849_, new_C9850_, new_C9851_, new_C9852_,
    new_C9853_, new_C9854_, new_C9855_, new_C9856_, new_C9857_, new_C9858_,
    new_C9859_, new_C9860_, new_C9861_, new_C9862_, new_C9863_, new_C9864_,
    new_C9865_, new_C9866_, new_C9867_, new_C9868_, new_C9869_, new_C9870_,
    new_C9871_, new_C9872_, new_C9873_, new_C9874_, new_C9875_, new_C9876_,
    new_C9877_, new_C9878_, new_C9879_, new_C9880_, new_C9881_, new_C9882_,
    new_C9883_, new_C9884_, new_C9885_, new_C9886_, new_C9887_, new_C9888_,
    new_C9889_, new_C9890_, new_C9891_, new_C9892_, new_C9893_, new_C9894_,
    new_C9895_, new_C9896_, new_C9897_, new_C9898_, new_C9899_, new_C9900_,
    new_C9901_, new_C9902_, new_C9903_, new_C9904_, new_C9905_, new_C9906_,
    new_C9907_, new_C9908_, new_C9909_, new_C9910_, new_C9911_, new_C9912_,
    new_C9913_, new_C9914_, new_C9915_, new_C9916_, new_C9917_, new_C9918_,
    new_C9919_, new_C9920_, new_C9921_, new_C9922_, new_C9923_, new_C9924_,
    new_C9925_, new_C9926_, new_C9927_, new_C9928_, new_C9929_, new_C9930_,
    new_C9931_, new_C9932_, new_C9933_, new_C9934_, new_C9935_, new_C9936_,
    new_C9937_, new_C9938_, new_C9939_, new_C9940_, new_C9941_, new_C9942_,
    new_C9943_, new_C9944_, new_C9945_, new_C9946_, new_C9947_, new_C9948_,
    new_C9949_, new_C9950_, new_C9951_, new_C9952_, new_C9953_, new_C9954_,
    new_C9955_, new_C9956_, new_C9957_, new_C9958_, new_C9959_, new_C9960_,
    new_C9961_, new_C9962_, new_C9963_, new_C9964_, new_C9965_, new_C9966_,
    new_C9967_, new_C9968_, new_C9969_, new_C9970_, new_C9971_, new_C9972_,
    new_C9973_, new_C9974_, new_C9975_, new_C9976_, new_C9977_, new_C9978_,
    new_C9979_, new_C9980_, new_C9981_, new_C9982_, new_C9983_, new_C9984_,
    new_C9985_, new_C9986_, new_C9987_, new_C9988_, new_C9989_, new_C9990_,
    new_C9991_, new_C9992_, new_C9993_, new_C9994_, new_C9995_, new_C9996_,
    new_C9997_, new_C9998_, new_C9999_, new_D1_, new_D2_, new_D3_, new_D4_,
    new_D5_, new_D6_, new_D7_, new_D8_, new_D9_, new_D10_, new_D11_,
    new_D12_, new_D13_, new_D14_, new_D15_, new_D16_, new_D17_, new_D18_,
    new_D19_, new_D20_, new_D21_, new_D22_, new_D23_, new_D24_, new_D25_,
    new_D26_, new_D27_, new_D28_, new_D29_, new_D30_, new_D31_, new_D32_,
    new_D33_, new_D34_, new_D35_, new_D36_, new_D37_, new_D38_, new_D39_,
    new_D40_, new_D41_, new_D42_, new_D43_, new_D44_, new_D45_, new_D46_,
    new_D47_, new_D48_, new_D49_, new_D50_, new_D51_, new_D52_, new_D53_,
    new_D54_, new_D55_, new_D56_, new_D57_, new_D58_, new_D59_, new_D60_,
    new_D61_, new_D62_, new_D63_, new_D64_, new_D65_, new_D66_, new_D67_,
    new_D68_, new_D69_, new_D70_, new_D71_, new_D72_, new_D73_, new_D74_,
    new_D75_, new_D76_, new_D77_, new_D78_, new_D79_, new_D80_, new_D81_,
    new_D82_, new_D83_, new_D84_, new_D85_, new_D86_, new_D87_, new_D88_,
    new_D89_, new_D90_, new_D91_, new_D92_, new_D93_, new_D94_, new_D95_,
    new_D96_, new_D97_, new_D98_, new_D99_, new_D100_, new_D101_,
    new_D102_, new_D103_, new_D104_, new_D105_, new_D106_, new_D107_,
    new_D108_, new_D109_, new_D110_, new_D111_, new_D112_, new_D113_,
    new_D114_, new_D115_, new_D116_, new_D117_, new_D118_, new_D119_,
    new_D120_, new_D121_, new_D122_, new_D123_, new_D124_, new_D125_,
    new_D126_, new_D127_, new_D128_, new_D129_, new_D130_, new_D131_,
    new_D132_, new_D133_, new_D134_, new_D135_, new_D136_, new_D137_,
    new_D138_, new_D139_, new_D140_, new_D141_, new_D142_, new_D143_,
    new_D144_, new_D145_, new_D146_, new_D147_, new_D148_, new_D149_,
    new_D150_, new_D151_, new_D152_, new_D153_, new_D154_, new_D155_,
    new_D156_, new_D157_, new_D158_, new_D159_, new_D160_, new_D161_,
    new_D162_, new_D163_, new_D164_, new_D165_, new_D166_, new_D167_,
    new_D168_, new_D169_, new_D170_, new_D171_, new_D172_, new_D173_,
    new_D174_, new_D175_, new_D176_, new_D177_, new_D178_, new_D179_,
    new_D180_, new_D181_, new_D182_, new_D183_, new_D184_, new_D185_,
    new_D186_, new_D187_, new_D188_, new_D189_, new_D190_, new_D191_,
    new_D192_, new_D193_, new_D194_, new_D195_, new_D196_, new_D197_,
    new_D198_, new_D199_, new_D200_, new_D201_, new_D202_, new_D203_,
    new_D204_, new_D205_, new_D206_, new_D207_, new_D208_, new_D209_,
    new_D210_, new_D211_, new_D212_, new_D213_, new_D214_, new_D215_,
    new_D216_, new_D217_, new_D218_, new_D219_, new_D220_, new_D221_,
    new_D222_, new_D223_, new_D224_, new_D225_, new_D226_, new_D227_,
    new_D228_, new_D229_, new_D230_, new_D231_, new_D232_, new_D233_,
    new_D234_, new_D235_, new_D236_, new_D237_, new_D238_, new_D239_,
    new_D240_, new_D241_, new_D242_, new_D243_, new_D244_, new_D245_,
    new_D246_, new_D247_, new_D248_, new_D249_, new_D250_, new_D251_,
    new_D252_, new_D253_, new_D254_, new_D255_, new_D256_, new_D257_,
    new_D258_, new_D259_, new_D260_, new_D261_, new_D262_, new_D263_,
    new_D264_, new_D265_, new_D266_, new_D267_, new_D268_, new_D269_,
    new_D270_, new_D271_, new_D272_, new_D273_, new_D274_, new_D275_,
    new_D276_, new_D277_, new_D278_, new_D279_, new_D280_, new_D281_,
    new_D282_, new_D283_, new_D284_, new_D285_, new_D286_, new_D287_,
    new_D288_, new_D289_, new_D290_, new_D291_, new_D292_, new_D293_,
    new_D294_, new_D295_, new_D296_, new_D297_, new_D298_, new_D299_,
    new_D300_, new_D301_, new_D302_, new_D303_, new_D304_, new_D305_,
    new_D306_, new_D307_, new_D308_, new_D309_, new_D310_, new_D311_,
    new_D312_, new_D313_, new_D314_, new_D315_, new_D316_, new_D317_,
    new_D318_, new_D319_, new_D320_, new_D321_, new_D322_, new_D323_,
    new_D324_, new_D325_, new_D326_, new_D327_, new_D328_, new_D329_,
    new_D330_, new_D331_, new_D332_, new_D333_, new_D334_, new_D335_,
    new_D336_, new_D337_, new_D338_, new_D339_, new_D340_, new_D341_,
    new_D342_, new_D343_, new_D344_, new_D345_, new_D346_, new_D347_,
    new_D348_, new_D349_, new_D350_, new_D351_, new_D352_, new_D353_,
    new_D354_, new_D355_, new_D356_, new_D357_, new_D358_, new_D359_,
    new_D360_, new_D361_, new_D362_, new_D363_, new_D364_, new_D365_,
    new_D366_, new_D367_, new_D368_, new_D369_, new_D370_, new_D371_,
    new_D372_, new_D373_, new_D374_, new_D375_, new_D376_, new_D377_,
    new_D378_, new_D379_, new_D380_, new_D381_, new_D382_, new_D383_,
    new_D384_, new_D385_, new_D386_, new_D387_, new_D388_, new_D389_,
    new_D390_, new_D391_, new_D392_, new_D393_, new_D394_, new_D395_,
    new_D396_, new_D397_, new_D398_, new_D399_, new_D400_, new_D401_,
    new_D402_, new_D403_, new_D404_, new_D405_, new_D406_, new_D407_,
    new_D408_, new_D409_, new_D410_, new_D411_, new_D412_, new_D413_,
    new_D414_, new_D415_, new_D416_, new_D417_, new_D418_, new_D419_,
    new_D420_, new_D421_, new_D422_, new_D423_, new_D424_, new_D425_,
    new_D426_, new_D427_, new_D428_, new_D429_, new_D430_, new_D431_,
    new_D432_, new_D433_, new_D434_, new_D435_, new_D436_, new_D437_,
    new_D438_, new_D439_, new_D440_, new_D441_, new_D442_, new_D443_,
    new_D444_, new_D445_, new_D446_, new_D447_, new_D448_, new_D449_,
    new_D450_, new_D451_, new_D452_, new_D453_, new_D454_, new_D455_,
    new_D456_, new_D457_, new_D458_, new_D459_, new_D460_, new_D461_,
    new_D462_, new_D463_, new_D464_, new_D465_, new_D466_, new_D467_,
    new_D468_, new_D469_, new_D470_, new_D471_, new_D472_, new_D473_,
    new_D474_, new_D475_, new_D476_, new_D477_, new_D478_, new_D479_,
    new_D480_, new_D481_, new_D482_, new_D483_, new_D484_, new_D485_,
    new_D486_, new_D487_, new_D488_, new_D489_, new_D490_, new_D491_,
    new_D492_, new_D493_, new_D494_, new_D495_, new_D496_, new_D497_,
    new_D498_, new_D499_, new_D500_, new_D501_, new_D502_, new_D503_,
    new_D504_, new_D505_, new_D506_, new_D507_, new_D508_, new_D509_,
    new_D510_, new_D511_, new_D512_, new_D513_, new_D514_, new_D515_,
    new_D516_, new_D517_, new_D518_, new_D519_, new_D520_, new_D521_,
    new_D522_, new_D523_, new_D524_, new_D525_, new_D526_, new_D527_,
    new_D528_, new_D529_, new_D530_, new_D531_, new_D532_, new_D533_,
    new_D534_, new_D535_, new_D536_, new_D537_, new_D538_, new_D539_,
    new_D540_, new_D541_, new_D542_, new_D543_, new_D544_, new_D545_,
    new_D546_, new_D547_, new_D548_, new_D549_, new_D550_, new_D551_,
    new_D552_, new_D553_, new_D554_, new_D555_, new_D556_, new_D557_,
    new_D558_, new_D559_, new_D560_, new_D561_, new_D562_, new_D563_,
    new_D564_, new_D565_, new_D566_, new_D567_, new_D568_, new_D569_,
    new_D570_, new_D571_, new_D572_, new_D573_, new_D574_, new_D575_,
    new_D576_, new_D577_, new_D578_, new_D579_, new_D580_, new_D581_,
    new_D582_, new_D583_, new_D584_, new_D585_, new_D586_, new_D587_,
    new_D588_, new_D589_, new_D590_, new_D591_, new_D592_, new_D593_,
    new_D594_, new_D595_, new_D596_, new_D597_, new_D598_, new_D599_,
    new_D600_, new_D601_, new_D602_, new_D603_, new_D604_, new_D605_,
    new_D606_, new_D607_, new_D608_, new_D609_, new_D610_, new_D611_,
    new_D612_, new_D613_, new_D614_, new_D615_, new_D616_, new_D617_,
    new_D618_, new_D619_, new_D620_, new_D621_, new_D622_, new_D623_,
    new_D624_, new_D625_, new_D626_, new_D627_, new_D628_, new_D629_,
    new_D630_, new_D631_, new_D632_, new_D633_, new_D634_, new_D635_,
    new_D636_, new_D637_, new_D638_, new_D639_, new_D640_, new_D641_,
    new_D642_, new_D643_, new_D644_, new_D645_, new_D646_, new_D647_,
    new_D648_, new_D649_, new_D650_, new_D651_, new_D652_, new_D653_,
    new_D654_, new_D655_, new_D656_, new_D657_, new_D658_, new_D659_,
    new_D660_, new_D661_, new_D662_, new_D663_, new_D664_, new_D665_,
    new_D666_, new_D667_, new_D668_, new_D669_, new_D670_, new_D671_,
    new_D672_, new_D673_, new_D674_, new_D675_, new_D676_, new_D677_,
    new_D678_, new_D679_, new_D680_, new_D681_, new_D682_, new_D683_,
    new_D684_, new_D685_, new_D686_, new_D687_, new_D688_, new_D689_,
    new_D690_, new_D691_, new_D692_, new_D693_, new_D694_, new_D695_,
    new_D696_, new_D697_, new_D698_, new_D699_, new_D700_, new_D701_,
    new_D702_, new_D703_, new_D704_, new_D705_, new_D706_, new_D707_,
    new_D708_, new_D709_, new_D710_, new_D711_, new_D712_, new_D713_,
    new_D714_, new_D715_, new_D716_, new_D717_, new_D718_, new_D719_,
    new_D720_, new_D721_, new_D722_, new_D723_, new_D724_, new_D725_,
    new_D726_, new_D727_, new_D728_, new_D729_, new_D730_, new_D731_,
    new_D732_, new_D733_, new_D734_, new_D735_, new_D736_, new_D737_,
    new_D738_, new_D739_, new_D740_, new_D741_, new_D742_, new_D743_,
    new_D744_, new_D745_, new_D746_, new_D747_, new_D748_, new_D749_,
    new_D750_, new_D751_, new_D752_, new_D753_, new_D754_, new_D755_,
    new_D756_, new_D757_, new_D758_, new_D759_, new_D760_, new_D761_,
    new_D762_, new_D763_, new_D764_, new_D765_, new_D766_, new_D767_,
    new_D768_, new_D769_, new_D770_, new_D771_, new_D772_, new_D773_,
    new_D774_, new_D775_, new_D776_, new_D777_, new_D778_, new_D779_,
    new_D780_, new_D781_, new_D782_, new_D783_, new_D784_, new_D785_,
    new_D786_, new_D787_, new_D788_, new_D789_, new_D790_, new_D791_,
    new_D792_, new_D793_, new_D794_, new_D795_, new_D796_, new_D797_,
    new_D798_, new_D799_, new_D800_, new_D801_, new_D802_, new_D803_,
    new_D804_, new_D805_, new_D806_, new_D807_, new_D808_, new_D809_,
    new_D810_, new_D811_, new_D812_, new_D813_, new_D814_, new_D815_,
    new_D816_, new_D817_, new_D818_, new_D819_, new_D820_, new_D821_,
    new_D822_, new_D823_, new_D824_, new_D825_, new_D826_, new_D827_,
    new_D828_, new_D829_, new_D830_, new_D831_, new_D832_, new_D833_,
    new_D834_, new_D835_, new_D836_, new_D837_, new_D838_, new_D839_,
    new_D840_, new_D841_, new_D842_, new_D843_, new_D844_, new_D845_,
    new_D846_, new_D847_, new_D848_, new_D849_, new_D850_, new_D851_,
    new_D852_, new_D853_, new_D854_, new_D855_, new_D856_, new_D857_,
    new_D858_, new_D859_, new_D860_, new_D861_, new_D862_, new_D863_,
    new_D864_, new_D865_, new_D866_, new_D867_, new_D868_, new_D869_,
    new_D870_, new_D871_, new_D872_, new_D873_, new_D874_, new_D875_,
    new_D876_, new_D877_, new_D878_, new_D879_, new_D880_, new_D881_,
    new_D882_, new_D883_, new_D884_, new_D885_, new_D886_, new_D887_,
    new_D888_, new_D889_, new_D890_, new_D891_, new_D892_, new_D893_,
    new_D894_, new_D895_, new_D896_, new_D897_, new_D898_, new_D899_,
    new_D900_, new_D901_, new_D902_, new_D903_, new_D904_, new_D905_,
    new_D906_, new_D907_, new_D908_, new_D909_, new_D910_, new_D911_,
    new_D912_, new_D913_, new_D914_, new_D915_, new_D916_, new_D917_,
    new_D918_, new_D919_, new_D920_, new_D921_, new_D922_, new_D923_,
    new_D924_, new_D925_, new_D926_, new_D927_, new_D928_, new_D929_,
    new_D930_, new_D931_, new_D932_, new_D933_, new_D934_, new_D935_,
    new_D936_, new_D937_, new_D938_, new_D939_, new_D940_, new_D941_,
    new_D942_, new_D943_, new_D944_, new_D945_, new_D946_, new_D947_,
    new_D948_, new_D949_, new_D950_, new_D951_, new_D952_, new_D953_,
    new_D954_, new_D955_, new_D956_, new_D957_, new_D958_, new_D959_,
    new_D960_, new_D961_, new_D962_, new_D963_, new_D964_, new_D965_,
    new_D966_, new_D967_, new_D968_, new_D969_, new_D970_, new_D971_,
    new_D972_, new_D973_, new_D974_, new_D975_, new_D976_, new_D977_,
    new_D978_, new_D979_, new_D980_, new_D981_, new_D982_, new_D983_,
    new_D984_, new_D985_, new_D986_, new_D987_, new_D988_, new_D989_,
    new_D990_, new_D991_, new_D992_, new_D993_, new_D994_, new_D995_,
    new_D996_, new_D997_, new_D998_, new_D999_, new_D1000_, new_D1001_,
    new_D1002_, new_D1003_, new_D1004_, new_D1005_, new_D1006_, new_D1007_,
    new_D1008_, new_D1009_, new_D1010_, new_D1011_, new_D1012_, new_D1013_,
    new_D1014_, new_D1015_, new_D1016_, new_D1017_, new_D1018_, new_D1019_,
    new_D1020_, new_D1021_, new_D1022_, new_D1023_, new_D1024_, new_D1025_,
    new_D1026_, new_D1027_, new_D1028_, new_D1029_, new_D1030_, new_D1031_,
    new_D1032_, new_D1033_, new_D1034_, new_D1035_, new_D1036_, new_D1037_,
    new_D1038_, new_D1039_, new_D1040_, new_D1041_, new_D1042_, new_D1043_,
    new_D1044_, new_D1045_, new_D1046_, new_D1047_, new_D1048_, new_D1049_,
    new_D1050_, new_D1051_, new_D1052_, new_D1053_, new_D1054_, new_D1055_,
    new_D1056_, new_D1057_, new_D1058_, new_D1059_, new_D1060_, new_D1061_,
    new_D1062_, new_D1063_, new_D1064_, new_D1065_, new_D1066_, new_D1067_,
    new_D1068_, new_D1069_, new_D1070_, new_D1071_, new_D1072_, new_D1073_,
    new_D1074_, new_D1075_, new_D1076_, new_D1077_, new_D1078_, new_D1079_,
    new_D1080_, new_D1081_, new_D1082_, new_D1083_, new_D1084_, new_D1085_,
    new_D1086_, new_D1087_, new_D1088_, new_D1089_, new_D1090_, new_D1091_,
    new_D1092_, new_D1093_, new_D1094_, new_D1095_, new_D1096_, new_D1097_,
    new_D1098_, new_D1099_, new_D1100_, new_D1101_, new_D1102_, new_D1103_,
    new_D1104_, new_D1105_, new_D1106_, new_D1107_, new_D1108_, new_D1109_,
    new_D1110_, new_D1111_, new_D1112_, new_D1113_, new_D1114_, new_D1115_,
    new_D1116_, new_D1117_, new_D1118_, new_D1119_, new_D1120_, new_D1121_,
    new_D1122_, new_D1123_, new_D1124_, new_D1125_, new_D1126_, new_D1127_,
    new_D1128_, new_D1129_, new_D1130_, new_D1131_, new_D1132_, new_D1133_,
    new_D1134_, new_D1135_, new_D1136_, new_D1137_, new_D1138_, new_D1139_,
    new_D1140_, new_D1141_, new_D1142_, new_D1143_, new_D1144_, new_D1145_,
    new_D1146_, new_D1147_, new_D1148_, new_D1149_, new_D1150_, new_D1151_,
    new_D1152_, new_D1153_, new_D1154_, new_D1155_, new_D1156_, new_D1157_,
    new_D1158_, new_D1159_, new_D1160_, new_D1161_, new_D1162_, new_D1163_,
    new_D1164_, new_D1165_, new_D1166_, new_D1167_, new_D1168_, new_D1169_,
    new_D1170_, new_D1171_, new_D1172_, new_D1173_, new_D1174_, new_D1175_,
    new_D1176_, new_D1177_, new_D1178_, new_D1179_, new_D1180_, new_D1181_,
    new_D1182_, new_D1183_, new_D1184_, new_D1185_, new_D1186_, new_D1187_,
    new_D1188_, new_D1189_, new_D1190_, new_D1191_, new_D1192_, new_D1193_,
    new_D1194_, new_D1195_, new_D1196_, new_D1197_, new_D1198_, new_D1199_,
    new_D1200_, new_D1201_, new_D1202_, new_D1203_, new_D1204_, new_D1205_,
    new_D1206_, new_D1207_, new_D1208_, new_D1209_, new_D1210_, new_D1211_,
    new_D1212_, new_D1213_, new_D1214_, new_D1215_, new_D1216_, new_D1217_,
    new_D1218_, new_D1219_, new_D1220_, new_D1221_, new_D1222_, new_D1223_,
    new_D1224_, new_D1225_, new_D1226_, new_D1227_, new_D1228_, new_D1229_,
    new_D1230_, new_D1231_, new_D1232_, new_D1233_, new_D1234_, new_D1235_,
    new_D1236_, new_D1237_, new_D1238_, new_D1239_, new_D1240_, new_D1241_,
    new_D1242_, new_D1243_, new_D1244_, new_D1245_, new_D1246_, new_D1247_,
    new_D1248_, new_D1249_, new_D1250_, new_D1251_, new_D1252_, new_D1253_,
    new_D1254_, new_D1255_, new_D1256_, new_D1257_, new_D1258_, new_D1259_,
    new_D1260_, new_D1261_, new_D1262_, new_D1263_, new_D1264_, new_D1265_,
    new_D1266_, new_D1267_, new_D1268_, new_D1269_, new_D1270_, new_D1271_,
    new_D1272_, new_D1273_, new_D1274_, new_D1275_, new_D1276_, new_D1277_,
    new_D1278_, new_D1279_, new_D1280_, new_D1281_, new_D1282_, new_D1283_,
    new_D1284_, new_D1285_, new_D1286_, new_D1287_, new_D1288_, new_D1289_,
    new_D1290_, new_D1291_, new_D1292_, new_D1293_, new_D1294_, new_D1295_,
    new_D1296_, new_D1297_, new_D1298_, new_D1299_, new_D1300_, new_D1301_,
    new_D1302_, new_D1303_, new_D1304_, new_D1305_, new_D1306_, new_D1307_,
    new_D1308_, new_D1309_, new_D1310_, new_D1311_, new_D1312_, new_D1313_,
    new_D1314_, new_D1315_, new_D1316_, new_D1317_, new_D1318_, new_D1319_,
    new_D1320_, new_D1321_, new_D1322_, new_D1323_, new_D1324_, new_D1325_,
    new_D1326_, new_D1327_, new_D1328_, new_D1329_, new_D1330_, new_D1331_,
    new_D1332_, new_D1333_, new_D1334_, new_D1335_, new_D1336_, new_D1337_,
    new_D1338_, new_D1339_, new_D1340_, new_D1341_, new_D1342_, new_D1343_,
    new_D1344_, new_D1345_, new_D1346_, new_D1347_, new_D1348_, new_D1349_,
    new_D1350_, new_D1351_, new_D1352_, new_D1353_, new_D1354_, new_D1355_,
    new_D1356_, new_D1357_, new_D1358_, new_D1359_, new_D1360_, new_D1361_,
    new_D1362_, new_D1363_, new_D1364_, new_D1365_, new_D1366_, new_D1367_,
    new_D1368_, new_D1369_, new_D1370_, new_D1371_, new_D1372_, new_D1373_,
    new_D1374_, new_D1375_, new_D1376_, new_D1377_, new_D1378_, new_D1379_,
    new_D1380_, new_D1381_, new_D1382_, new_D1383_, new_D1384_, new_D1385_,
    new_D1386_, new_D1387_, new_D1388_, new_D1389_, new_D1390_, new_D1391_,
    new_D1392_, new_D1393_, new_D1394_, new_D1395_, new_D1396_, new_D1397_,
    new_D1398_, new_D1399_, new_D1400_, new_D1401_, new_D1402_, new_D1403_,
    new_D1404_, new_D1405_, new_D1406_, new_D1407_, new_D1408_, new_D1409_,
    new_D1410_, new_D1411_, new_D1412_, new_D1413_, new_D1414_, new_D1415_,
    new_D1416_, new_D1417_, new_D1418_, new_D1419_, new_D1420_, new_D1421_,
    new_D1422_, new_D1423_, new_D1424_, new_D1425_, new_D1426_, new_D1427_,
    new_D1428_, new_D1429_, new_D1430_, new_D1431_, new_D1432_, new_D1433_,
    new_D1434_, new_D1435_, new_D1436_, new_D1437_, new_D1438_, new_D1439_,
    new_D1440_, new_D1441_, new_D1442_, new_D1443_, new_D1444_, new_D1445_,
    new_D1446_, new_D1447_, new_D1448_, new_D1449_, new_D1450_, new_D1451_,
    new_D1452_, new_D1453_, new_D1454_, new_D1455_, new_D1456_, new_D1457_,
    new_D1458_, new_D1459_, new_D1460_, new_D1461_, new_D1462_, new_D1463_,
    new_D1464_, new_D1465_, new_D1466_, new_D1467_, new_D1468_, new_D1469_,
    new_D1470_, new_D1471_, new_D1472_, new_D1473_, new_D1474_, new_D1475_,
    new_D1476_, new_D1477_, new_D1478_, new_D1479_, new_D1480_, new_D1481_,
    new_D1482_, new_D1483_, new_D1484_, new_D1485_, new_D1486_, new_D1487_,
    new_D1488_, new_D1489_, new_D1490_, new_D1491_, new_D1492_, new_D1493_,
    new_D1494_, new_D1495_, new_D1496_, new_D1497_, new_D1498_, new_D1499_,
    new_D1500_, new_D1501_, new_D1502_, new_D1503_, new_D1504_, new_D1505_,
    new_D1506_, new_D1507_, new_D1508_, new_D1509_, new_D1510_, new_D1511_,
    new_D1512_, new_D1513_, new_D1514_, new_D1515_, new_D1516_, new_D1517_,
    new_D1518_, new_D1519_, new_D1520_, new_D1521_, new_D1522_, new_D1523_,
    new_D1524_, new_D1525_, new_D1526_, new_D1527_, new_D1528_, new_D1529_,
    new_D1530_, new_D1531_, new_D1532_, new_D1533_, new_D1534_, new_D1535_,
    new_D1536_, new_D1537_, new_D1538_, new_D1539_, new_D1540_, new_D1541_,
    new_D1542_, new_D1543_, new_D1544_, new_D1545_, new_D1546_, new_D1547_,
    new_D1548_, new_D1549_, new_D1550_, new_D1551_, new_D1552_, new_D1553_,
    new_D1554_, new_D1555_, new_D1556_, new_D1557_, new_D1558_, new_D1559_,
    new_D1560_, new_D1561_, new_D1562_, new_D1563_, new_D1564_, new_D1565_,
    new_D1566_, new_D1567_, new_D1568_, new_D1569_, new_D1570_, new_D1571_,
    new_D1572_, new_D1573_, new_D1574_, new_D1575_, new_D1576_, new_D1577_,
    new_D1578_, new_D1579_, new_D1580_, new_D1581_, new_D1582_, new_D1583_,
    new_D1584_, new_D1585_, new_D1586_, new_D1587_, new_D1588_, new_D1589_,
    new_D1590_, new_D1591_, new_D1592_, new_D1593_, new_D1594_, new_D1595_,
    new_D1596_, new_D1597_, new_D1598_, new_D1599_, new_D1600_, new_D1601_,
    new_D1602_, new_D1603_, new_D1604_, new_D1605_, new_D1606_, new_D1607_,
    new_D1608_, new_D1609_, new_D1610_, new_D1611_, new_D1612_, new_D1613_,
    new_D1614_, new_D1615_, new_D1616_, new_D1617_, new_D1618_, new_D1619_,
    new_D1620_, new_D1621_, new_D1622_, new_D1623_, new_D1624_, new_D1625_,
    new_D1626_, new_D1627_, new_D1628_, new_D1629_, new_D1630_, new_D1631_,
    new_D1632_, new_D1633_, new_D1634_, new_D1635_, new_D1636_, new_D1637_,
    new_D1638_, new_D1639_, new_D1640_, new_D1641_, new_D1642_, new_D1643_,
    new_D1644_, new_D1645_, new_D1646_, new_D1647_, new_D1648_, new_D1649_,
    new_D1650_, new_D1651_, new_D1652_, new_D1653_, new_D1654_, new_D1655_,
    new_D1656_, new_D1657_, new_D1658_, new_D1659_, new_D1660_, new_D1661_,
    new_D1662_, new_D1663_, new_D1664_, new_D1665_, new_D1666_, new_D1667_,
    new_D1668_, new_D1669_, new_D1670_, new_D1671_, new_D1672_, new_D1673_,
    new_D1674_, new_D1675_, new_D1676_, new_D1677_, new_D1678_, new_D1679_,
    new_D1680_, new_D1681_, new_D1682_, new_D1683_, new_D1684_, new_D1685_,
    new_D1686_, new_D1687_, new_D1688_, new_D1689_, new_D1690_, new_D1691_,
    new_D1692_, new_D1693_, new_D1694_, new_D1695_, new_D1696_, new_D1697_,
    new_D1698_, new_D1699_, new_D1700_, new_D1701_, new_D1702_, new_D1703_,
    new_D1704_, new_D1705_, new_D1706_, new_D1707_, new_D1708_, new_D1709_,
    new_D1710_, new_D1711_, new_D1712_, new_D1713_, new_D1714_, new_D1715_,
    new_D1716_, new_D1717_, new_D1718_, new_D1719_, new_D1720_, new_D1721_,
    new_D1722_, new_D1723_, new_D1724_, new_D1725_, new_D1726_, new_D1727_,
    new_D1728_, new_D1729_, new_D1730_, new_D1731_, new_D1732_, new_D1733_,
    new_D1734_, new_D1735_, new_D1736_, new_D1737_, new_D1738_, new_D1739_,
    new_D1740_, new_D1741_, new_D1742_, new_D1743_, new_D1744_, new_D1745_,
    new_D1746_, new_D1747_, new_D1748_, new_D1749_, new_D1750_, new_D1751_,
    new_D1752_, new_D1753_, new_D1754_, new_D1755_, new_D1756_, new_D1757_,
    new_D1758_, new_D1759_, new_D1760_, new_D1761_, new_D1762_, new_D1763_,
    new_D1764_, new_D1765_, new_D1766_, new_D1767_, new_D1768_, new_D1769_,
    new_D1770_, new_D1771_, new_D1772_, new_D1773_, new_D1774_, new_D1775_,
    new_D1776_, new_D1777_, new_D1778_, new_D1779_, new_D1780_, new_D1781_,
    new_D1782_, new_D1783_, new_D1784_, new_D1785_, new_D1786_, new_D1787_,
    new_D1788_, new_D1789_, new_D1790_, new_D1791_, new_D1792_, new_D1793_,
    new_D1794_, new_D1795_, new_D1796_, new_D1797_, new_D1798_, new_D1799_,
    new_D1800_, new_D1801_, new_D1802_, new_D1803_, new_D1804_, new_D1805_,
    new_D1806_, new_D1807_, new_D1808_, new_D1809_, new_D1810_, new_D1811_,
    new_D1812_, new_D1813_, new_D1814_, new_D1815_, new_D1816_, new_D1817_,
    new_D1818_, new_D1819_, new_D1820_, new_D1821_, new_D1822_, new_D1823_,
    new_D1824_, new_D1825_, new_D1826_, new_D1827_, new_D1828_, new_D1829_,
    new_D1830_, new_D1831_, new_D1832_, new_D1833_, new_D1834_, new_D1835_,
    new_D1836_, new_D1837_, new_D1838_, new_D1839_, new_D1840_, new_D1841_,
    new_D1842_, new_D1843_, new_D1844_, new_D1845_, new_D1846_, new_D1847_,
    new_D1848_, new_D1849_, new_D1850_, new_D1851_, new_D1852_, new_D1853_,
    new_D1854_, new_D1855_, new_D1856_, new_D1857_, new_D1858_, new_D1859_,
    new_D1860_, new_D1861_, new_D1862_, new_D1863_, new_D1864_, new_D1865_,
    new_D1866_, new_D1867_, new_D1868_, new_D1869_, new_D1870_, new_D1871_,
    new_D1872_, new_D1873_, new_D1874_, new_D1875_, new_D1876_, new_D1877_,
    new_D1878_, new_D1879_, new_D1880_, new_D1881_, new_D1882_, new_D1883_,
    new_D1884_, new_D1885_, new_D1886_, new_D1887_, new_D1888_, new_D1889_,
    new_D1890_, new_D1891_, new_D1892_, new_D1893_, new_D1894_, new_D1895_,
    new_D1896_, new_D1897_, new_D1898_, new_D1899_, new_D1900_, new_D1901_,
    new_D1902_, new_D1903_, new_D1904_, new_D1905_, new_D1906_, new_D1907_,
    new_D1908_, new_D1909_, new_D1910_, new_D1911_, new_D1912_, new_D1913_,
    new_D1914_, new_D1915_, new_D1916_, new_D1917_, new_D1918_, new_D1919_,
    new_D1920_, new_D1921_, new_D1922_, new_D1923_, new_D1924_, new_D1925_,
    new_D1926_, new_D1927_, new_D1928_, new_D1929_, new_D1930_, new_D1931_,
    new_D1932_, new_D1933_, new_D1934_, new_D1935_, new_D1936_, new_D1937_,
    new_D1938_, new_D1939_, new_D1940_, new_D1941_, new_D1942_, new_D1943_,
    new_D1944_, new_D1945_, new_D1946_, new_D1947_, new_D1948_, new_D1949_,
    new_D1950_, new_D1951_, new_D1952_, new_D1953_, new_D1954_, new_D1955_,
    new_D1956_, new_D1957_, new_D1958_, new_D1959_, new_D1960_, new_D1961_,
    new_D1962_, new_D1963_, new_D1964_, new_D1965_, new_D1966_, new_D1967_,
    new_D1968_, new_D1969_, new_D1970_, new_D1971_, new_D1972_, new_D1973_,
    new_D1974_, new_D1975_, new_D1976_, new_D1977_, new_D1978_, new_D1979_,
    new_D1980_, new_D1981_, new_D1982_, new_D1983_, new_D1984_, new_D1985_,
    new_D1986_, new_D1987_, new_D1988_, new_D1989_, new_D1990_, new_D1991_,
    new_D1992_, new_D1993_, new_D1994_, new_D1995_, new_D1996_, new_D1997_,
    new_D1998_, new_D1999_, new_D2000_, new_D2001_, new_D2002_, new_D2003_,
    new_D2004_, new_D2005_, new_D2006_, new_D2007_, new_D2008_, new_D2009_,
    new_D2010_, new_D2011_, new_D2012_, new_D2013_, new_D2014_, new_D2015_,
    new_D2016_, new_D2017_, new_D2018_, new_D2019_, new_D2020_, new_D2021_,
    new_D2022_, new_D2023_, new_D2024_, new_D2025_, new_D2026_, new_D2027_,
    new_D2028_, new_D2029_, new_D2030_, new_D2031_, new_D2032_, new_D2033_,
    new_D2034_, new_D2035_, new_D2036_, new_D2037_, new_D2038_, new_D2039_,
    new_D2040_, new_D2041_, new_D2042_, new_D2043_, new_D2044_, new_D2045_,
    new_D2046_, new_D2047_, new_D2048_, new_D2049_, new_D2050_, new_D2051_,
    new_D2052_, new_D2053_, new_D2054_, new_D2055_, new_D2056_, new_D2057_,
    new_D2058_, new_D2059_, new_D2060_, new_D2061_, new_D2062_, new_D2063_,
    new_D2064_, new_D2065_, new_D2066_, new_D2067_, new_D2068_, new_D2069_,
    new_D2070_, new_D2071_, new_D2072_, new_D2073_, new_D2074_, new_D2075_,
    new_D2076_, new_D2077_, new_D2078_, new_D2079_, new_D2080_, new_D2081_,
    new_D2082_, new_D2083_, new_D2084_, new_D2085_, new_D2086_, new_D2087_,
    new_D2088_, new_D2089_, new_D2090_, new_D2091_, new_D2092_, new_D2093_,
    new_D2094_, new_D2095_, new_D2096_, new_D2097_, new_D2098_, new_D2099_,
    new_D2100_, new_D2101_, new_D2102_, new_D2103_, new_D2104_, new_D2105_,
    new_D2106_, new_D2107_, new_D2108_, new_D2109_, new_D2110_, new_D2111_,
    new_D2112_, new_D2113_, new_D2114_, new_D2115_, new_D2116_, new_D2117_,
    new_D2118_, new_D2119_, new_D2120_, new_D2121_, new_D2122_, new_D2123_,
    new_D2124_, new_D2125_, new_D2126_, new_D2127_, new_D2128_, new_D2129_,
    new_D2130_, new_D2131_, new_D2132_, new_D2133_, new_D2134_, new_D2135_,
    new_D2136_, new_D2137_, new_D2138_, new_D2139_, new_D2140_, new_D2141_,
    new_D2142_, new_D2143_, new_D2144_, new_D2145_, new_D2146_, new_D2147_,
    new_D2148_, new_D2149_, new_D2150_, new_D2151_, new_D2152_, new_D2153_,
    new_D2154_, new_D2155_, new_D2156_, new_D2157_, new_D2158_, new_D2159_,
    new_D2160_, new_D2161_, new_D2162_, new_D2163_, new_D2164_, new_D2165_,
    new_D2166_, new_D2167_, new_D2168_, new_D2169_, new_D2170_, new_D2171_,
    new_D2172_, new_D2173_, new_D2174_, new_D2175_, new_D2176_, new_D2177_,
    new_D2178_, new_D2179_, new_D2180_, new_D2181_, new_D2182_, new_D2183_,
    new_D2184_, new_D2185_, new_D2186_, new_D2187_, new_D2188_, new_D2189_,
    new_D2190_, new_D2191_, new_D2192_, new_D2193_, new_D2194_, new_D2195_,
    new_D2196_, new_D2197_, new_D2198_, new_D2199_, new_D2200_, new_D2201_,
    new_D2202_, new_D2203_, new_D2204_, new_D2205_, new_D2206_, new_D2207_,
    new_D2208_, new_D2209_, new_D2210_, new_D2211_, new_D2212_, new_D2213_,
    new_D2214_, new_D2215_, new_D2216_, new_D2217_, new_D2218_, new_D2219_,
    new_D2220_, new_D2221_, new_D2222_, new_D2223_, new_D2224_, new_D2225_,
    new_D2226_, new_D2227_, new_D2228_, new_D2229_, new_D2230_, new_D2231_,
    new_D2232_, new_D2233_, new_D2234_, new_D2235_, new_D2236_, new_D2237_,
    new_D2238_, new_D2239_, new_D2240_, new_D2241_, new_D2242_, new_D2243_,
    new_D2244_, new_D2245_, new_D2246_, new_D2247_, new_D2248_, new_D2249_,
    new_D2250_, new_D2251_, new_D2252_, new_D2253_, new_D2254_, new_D2255_,
    new_D2256_, new_D2257_, new_D2258_, new_D2259_, new_D2260_, new_D2261_,
    new_D2262_, new_D2263_, new_D2264_, new_D2265_, new_D2266_, new_D2267_,
    new_D2268_, new_D2269_, new_D2270_, new_D2271_, new_D2272_, new_D2273_,
    new_D2274_, new_D2275_, new_D2276_, new_D2277_, new_D2278_, new_D2279_,
    new_D2280_, new_D2281_, new_D2282_, new_D2283_, new_D2284_, new_D2285_,
    new_D2286_, new_D2287_, new_D2288_, new_D2289_, new_D2290_, new_D2291_,
    new_D2292_, new_D2293_, new_D2294_, new_D2295_, new_D2296_, new_D2297_,
    new_D2298_, new_D2299_, new_D2300_, new_D2301_, new_D2302_, new_D2303_,
    new_D2304_, new_D2305_, new_D2306_, new_D2307_, new_D2308_, new_D2309_,
    new_D2310_, new_D2311_, new_D2312_, new_D2313_, new_D2314_, new_D2315_,
    new_D2316_, new_D2317_, new_D2318_, new_D2319_, new_D2320_, new_D2321_,
    new_D2322_, new_D2323_, new_D2324_, new_D2325_, new_D2326_, new_D2327_,
    new_D2328_, new_D2329_, new_D2330_, new_D2331_, new_D2332_, new_D2333_,
    new_D2334_, new_D2335_, new_D2336_, new_D2337_, new_D2338_, new_D2339_,
    new_D2340_, new_D2341_, new_D2342_, new_D2343_, new_D2344_, new_D2345_,
    new_D2346_, new_D2347_, new_D2348_, new_D2349_, new_D2350_, new_D2351_,
    new_D2352_, new_D2353_, new_D2354_, new_D2355_, new_D2356_, new_D2357_,
    new_D2358_, new_D2359_, new_D2360_, new_D2361_, new_D2362_, new_D2363_,
    new_D2364_, new_D2365_, new_D2366_, new_D2367_, new_D2368_, new_D2369_,
    new_D2370_, new_D2371_, new_D2372_, new_D2373_, new_D2374_, new_D2375_,
    new_D2376_, new_D2377_, new_D2378_, new_D2379_, new_D2380_, new_D2381_,
    new_D2382_, new_D2383_, new_D2384_, new_D2385_, new_D2386_, new_D2387_,
    new_D2388_, new_D2389_, new_D2390_, new_D2391_, new_D2392_, new_D2393_,
    new_D2394_, new_D2395_, new_D2396_, new_D2397_, new_D2398_, new_D2399_,
    new_D2400_, new_D2401_, new_D2402_, new_D2403_, new_D2404_, new_D2405_,
    new_D2406_, new_D2407_, new_D2408_, new_D2409_, new_D2410_, new_D2411_,
    new_D2412_, new_D2413_, new_D2414_, new_D2415_, new_D2416_, new_D2417_,
    new_D2418_, new_D2419_, new_D2420_, new_D2421_, new_D2422_, new_D2423_,
    new_D2424_, new_D2425_, new_D2426_, new_D2427_, new_D2428_, new_D2429_,
    new_D2430_, new_D2431_, new_D2432_, new_D2433_, new_D2434_, new_D2435_,
    new_D2436_, new_D2437_, new_D2438_, new_D2439_, new_D2440_, new_D2441_,
    new_D2442_, new_D2443_, new_D2444_, new_D2445_, new_D2446_, new_D2447_,
    new_D2448_, new_D2449_, new_D2450_, new_D2451_, new_D2452_, new_D2453_,
    new_D2454_, new_D2455_, new_D2456_, new_D2457_, new_D2458_, new_D2459_,
    new_D2460_, new_D2461_, new_D2462_, new_D2463_, new_D2464_, new_D2465_,
    new_D2466_, new_D2467_, new_D2468_, new_D2469_, new_D2470_, new_D2471_,
    new_D2472_, new_D2473_, new_D2474_, new_D2475_, new_D2476_, new_D2477_,
    new_D2478_, new_D2479_, new_D2480_, new_D2481_, new_D2482_, new_D2483_,
    new_D2484_, new_D2485_, new_D2486_, new_D2487_, new_D2488_, new_D2489_,
    new_D2490_, new_D2491_, new_D2492_, new_D2493_, new_D2494_, new_D2495_,
    new_D2496_, new_D2497_, new_D2498_, new_D2499_, new_D2500_, new_D2501_,
    new_D2502_, new_D2503_, new_D2504_, new_D2505_, new_D2506_, new_D2507_,
    new_D2508_, new_D2509_, new_D2510_, new_D2511_, new_D2512_, new_D2513_,
    new_D2514_, new_D2515_, new_D2516_, new_D2517_, new_D2518_, new_D2519_,
    new_D2520_, new_D2521_, new_D2522_, new_D2523_, new_D2524_, new_D2525_,
    new_D2526_, new_D2527_, new_D2528_, new_D2529_, new_D2530_, new_D2531_,
    new_D2532_, new_D2533_, new_D2534_, new_D2535_, new_D2536_, new_D2537_,
    new_D2538_, new_D2539_, new_D2540_, new_D2541_, new_D2542_, new_D2543_,
    new_D2544_, new_D2545_, new_D2546_, new_D2547_, new_D2548_, new_D2549_,
    new_D2550_, new_D2551_, new_D2552_, new_D2553_, new_D2554_, new_D2555_,
    new_D2556_, new_D2557_, new_D2558_, new_D2559_, new_D2560_, new_D2561_,
    new_D2562_, new_D2563_, new_D2564_, new_D2565_, new_D2566_, new_D2567_,
    new_D2568_, new_D2569_, new_D2570_, new_D2571_, new_D2572_, new_D2573_,
    new_D2574_, new_D2575_, new_D2576_, new_D2577_, new_D2578_, new_D2579_,
    new_D2580_, new_D2581_, new_D2582_, new_D2583_, new_D2584_, new_D2585_,
    new_D2586_, new_D2587_, new_D2588_, new_D2589_, new_D2590_, new_D2591_,
    new_D2592_, new_D2593_, new_D2594_, new_D2595_, new_D2596_, new_D2597_,
    new_D2598_, new_D2599_, new_D2600_, new_D2601_, new_D2602_, new_D2603_,
    new_D2604_, new_D2605_, new_D2606_, new_D2607_, new_D2608_, new_D2609_,
    new_D2610_, new_D2611_, new_D2612_, new_D2613_, new_D2614_, new_D2615_,
    new_D2616_, new_D2617_, new_D2618_, new_D2619_, new_D2620_, new_D2621_,
    new_D2622_, new_D2623_, new_D2624_, new_D2625_, new_D2626_, new_D2627_,
    new_D2628_, new_D2629_, new_D2630_, new_D2631_, new_D2632_, new_D2633_,
    new_D2634_, new_D2635_, new_D2636_, new_D2637_, new_D2638_, new_D2639_,
    new_D2640_, new_D2641_, new_D2642_, new_D2643_, new_D2644_, new_D2645_,
    new_D2646_, new_D2647_, new_D2648_, new_D2649_, new_D2650_, new_D2651_,
    new_D2652_, new_D2653_, new_D2654_, new_D2655_, new_D2656_, new_D2657_,
    new_D2658_, new_D2659_, new_D2660_, new_D2661_, new_D2662_, new_D2663_,
    new_D2664_, new_D2665_, new_D2666_, new_D2667_, new_D2668_, new_D2669_,
    new_D2670_, new_D2671_, new_D2672_, new_D2673_, new_D2674_, new_D2675_,
    new_D2676_, new_D2677_, new_D2678_, new_D2679_, new_D2680_, new_D2681_,
    new_D2682_, new_D2683_, new_D2684_, new_D2685_, new_D2686_, new_D2687_,
    new_D2688_, new_D2689_, new_D2690_, new_D2691_, new_D2692_, new_D2693_,
    new_D2694_, new_D2695_, new_D2696_, new_D2697_, new_D2698_, new_D2699_,
    new_D2700_, new_D2701_, new_D2702_, new_D2703_, new_D2704_, new_D2705_,
    new_D2706_, new_D2707_, new_D2708_, new_D2709_, new_D2710_, new_D2711_,
    new_D2712_, new_D2713_, new_D2714_, new_D2715_, new_D2716_, new_D2717_,
    new_D2718_, new_D2719_, new_D2720_, new_D2721_, new_D2722_, new_D2723_,
    new_D2724_, new_D2725_, new_D2726_, new_D2727_, new_D2728_, new_D2729_,
    new_D2730_, new_D2731_, new_D2732_, new_D2733_, new_D2734_, new_D2735_,
    new_D2736_, new_D2737_, new_D2738_, new_D2739_, new_D2740_, new_D2741_,
    new_D2742_, new_D2743_, new_D2744_, new_D2745_, new_D2746_, new_D2747_,
    new_D2748_, new_D2749_, new_D2750_, new_D2751_, new_D2752_, new_D2753_,
    new_D2754_, new_D2755_, new_D2756_, new_D2757_, new_D2758_, new_D2759_,
    new_D2760_, new_D2761_, new_D2762_, new_D2763_, new_D2764_, new_D2765_,
    new_D2766_, new_D2767_, new_D2768_, new_D2769_, new_D2770_, new_D2771_,
    new_D2772_, new_D2773_, new_D2774_, new_D2775_, new_D2776_, new_D2777_,
    new_D2778_, new_D2779_, new_D2780_, new_D2781_, new_D2782_, new_D2783_,
    new_D2784_, new_D2785_, new_D2786_, new_D2787_, new_D2788_, new_D2789_,
    new_D2790_, new_D2791_, new_D2792_, new_D2793_, new_D2794_, new_D2795_,
    new_D2796_, new_D2797_, new_D2798_, new_D2799_, new_D2800_, new_D2801_,
    new_D2802_, new_D2803_, new_D2804_, new_D2805_, new_D2806_, new_D2807_,
    new_D2808_, new_D2809_, new_D2810_, new_D2811_, new_D2812_, new_D2813_,
    new_D2814_, new_D2815_, new_D2816_, new_D2817_, new_D2818_, new_D2819_,
    new_D2820_, new_D2821_, new_D2822_, new_D2823_, new_D2824_, new_D2825_,
    new_D2826_, new_D2827_, new_D2828_, new_D2829_, new_D2830_, new_D2831_,
    new_D2832_, new_D2833_, new_D2834_, new_D2835_, new_D2836_, new_D2837_,
    new_D2838_, new_D2839_, new_D2840_, new_D2841_, new_D2842_, new_D2843_,
    new_D2844_, new_D2845_, new_D2846_, new_D2847_, new_D2848_, new_D2849_,
    new_D2850_, new_D2851_, new_D2852_, new_D2853_, new_D2854_, new_D2855_,
    new_D2856_, new_D2857_, new_D2858_, new_D2859_, new_D2860_, new_D2861_,
    new_D2862_, new_D2863_, new_D2864_, new_D2865_, new_D2866_, new_D2867_,
    new_D2868_, new_D2869_, new_D2870_, new_D2871_, new_D2872_, new_D2873_,
    new_D2874_, new_D2875_, new_D2876_, new_D2877_, new_D2878_, new_D2879_,
    new_D2880_, new_D2881_, new_D2882_, new_D2883_, new_D2884_, new_D2885_,
    new_D2886_, new_D2887_, new_D2888_, new_D2889_, new_D2890_, new_D2891_,
    new_D2892_, new_D2893_, new_D2894_, new_D2895_, new_D2896_, new_D2897_,
    new_D2898_, new_D2899_, new_D2900_, new_D2901_, new_D2902_, new_D2903_,
    new_D2904_, new_D2905_, new_D2906_, new_D2907_, new_D2908_, new_D2909_,
    new_D2910_, new_D2911_, new_D2912_, new_D2913_, new_D2914_, new_D2915_,
    new_D2916_, new_D2917_, new_D2918_, new_D2919_, new_D2920_, new_D2921_,
    new_D2922_, new_D2923_, new_D2924_, new_D2925_, new_D2926_, new_D2927_,
    new_D2928_, new_D2929_, new_D2930_, new_D2931_, new_D2932_, new_D2933_,
    new_D2934_, new_D2935_, new_D2936_, new_D2937_, new_D2938_, new_D2939_,
    new_D2940_, new_D2941_, new_D2942_, new_D2943_, new_D2944_, new_D2945_,
    new_D2946_, new_D2947_, new_D2948_, new_D2949_, new_D2950_, new_D2951_,
    new_D2952_, new_D2953_, new_D2954_, new_D2955_, new_D2956_, new_D2957_,
    new_D2958_, new_D2959_, new_D2960_, new_D2961_, new_D2962_, new_D2963_,
    new_D2964_, new_D2965_, new_D2966_, new_D2967_, new_D2968_, new_D2969_,
    new_D2970_, new_D2971_, new_D2972_, new_D2973_, new_D2974_, new_D2975_,
    new_D2976_, new_D2977_, new_D2978_, new_D2979_, new_D2980_, new_D2981_,
    new_D2982_, new_D2983_, new_D2984_, new_D2985_, new_D2986_, new_D2987_,
    new_D2988_, new_D2989_, new_D2990_, new_D2991_, new_D2992_, new_D2993_,
    new_D2994_, new_D2995_, new_D2996_, new_D2997_, new_D2998_, new_D2999_,
    new_D3000_, new_D3001_, new_D3002_, new_D3003_, new_D3004_, new_D3005_,
    new_D3006_, new_D3007_, new_D3008_, new_D3009_, new_D3010_, new_D3011_,
    new_D3012_, new_D3013_, new_D3014_, new_D3015_, new_D3016_, new_D3017_,
    new_D3018_, new_D3019_, new_D3020_, new_D3021_, new_D3022_, new_D3023_,
    new_D3024_, new_D3025_, new_D3026_, new_D3027_, new_D3028_, new_D3029_,
    new_D3030_, new_D3031_, new_D3032_, new_D3033_, new_D3034_, new_D3035_,
    new_D3036_, new_D3037_, new_D3038_, new_D3039_, new_D3040_, new_D3041_,
    new_D3042_, new_D3043_, new_D3044_, new_D3045_, new_D3046_, new_D3047_,
    new_D3048_, new_D3049_, new_D3050_, new_D3051_, new_D3052_, new_D3053_,
    new_D3054_, new_D3055_, new_D3056_, new_D3057_, new_D3058_, new_D3059_,
    new_D3060_, new_D3061_, new_D3062_, new_D3063_, new_D3064_, new_D3065_,
    new_D3066_, new_D3067_, new_D3068_, new_D3069_, new_D3070_, new_D3071_,
    new_D3072_, new_D3073_, new_D3074_, new_D3075_, new_D3076_, new_D3077_,
    new_D3078_, new_D3079_, new_D3080_, new_D3081_, new_D3082_, new_D3083_,
    new_D3084_, new_D3085_, new_D3086_, new_D3087_, new_D3088_, new_D3089_,
    new_D3090_, new_D3091_, new_D3092_, new_D3093_, new_D3094_, new_D3095_,
    new_D3096_, new_D3097_, new_D3098_, new_D3099_, new_D3100_, new_D3101_,
    new_D3102_, new_D3103_, new_D3104_, new_D3105_, new_D3106_, new_D3107_,
    new_D3108_, new_D3109_, new_D3110_, new_D3111_, new_D3112_, new_D3113_,
    new_D3114_, new_D3115_, new_D3116_, new_D3117_, new_D3118_, new_D3119_,
    new_D3120_, new_D3121_, new_D3122_, new_D3123_, new_D3124_, new_D3125_,
    new_D3126_, new_D3127_, new_D3128_, new_D3129_, new_D3130_, new_D3131_,
    new_D3132_, new_D3133_, new_D3134_, new_D3135_, new_D3136_, new_D3137_,
    new_D3138_, new_D3139_, new_D3140_, new_D3141_, new_D3142_, new_D3143_,
    new_D3144_, new_D3145_, new_D3146_, new_D3147_, new_D3148_, new_D3149_,
    new_D3150_, new_D3151_, new_D3152_, new_D3153_, new_D3154_, new_D3155_,
    new_D3156_, new_D3157_, new_D3158_, new_D3159_, new_D3160_, new_D3161_,
    new_D3162_, new_D3163_, new_D3164_, new_D3165_, new_D3166_, new_D3167_,
    new_D3168_, new_D3169_, new_D3170_, new_D3171_, new_D3172_, new_D3173_,
    new_D3174_, new_D3175_, new_D3176_, new_D3177_, new_D3178_, new_D3179_,
    new_D3180_, new_D3181_, new_D3182_, new_D3183_, new_D3184_, new_D3185_,
    new_D3186_, new_D3187_, new_D3188_, new_D3189_, new_D3190_, new_D3191_,
    new_D3192_, new_D3193_, new_D3194_, new_D3195_, new_D3196_, new_D3197_,
    new_D3198_, new_D3199_, new_D3200_, new_D3201_, new_D3202_, new_D3203_,
    new_D3204_, new_D3205_, new_D3206_, new_D3207_, new_D3208_, new_D3209_,
    new_D3210_, new_D3211_, new_D3212_, new_D3213_, new_D3214_, new_D3215_,
    new_D3216_, new_D3217_, new_D3218_, new_D3219_, new_D3220_, new_D3221_,
    new_D3222_, new_D3223_, new_D3224_, new_D3225_, new_D3226_, new_D3227_,
    new_D3228_, new_D3229_, new_D3230_, new_D3231_, new_D3232_, new_D3233_,
    new_D3234_, new_D3235_, new_D3236_, new_D3237_, new_D3238_, new_D3239_,
    new_D3240_, new_D3241_, new_D3242_, new_D3243_, new_D3244_, new_D3245_,
    new_D3246_, new_D3247_, new_D3248_, new_D3249_, new_D3250_, new_D3251_,
    new_D3252_, new_D3253_, new_D3254_, new_D3255_, new_D3256_, new_D3257_,
    new_D3258_, new_D3259_, new_D3260_, new_D3261_, new_D3262_, new_D3263_,
    new_D3264_, new_D3265_, new_D3266_, new_D3267_, new_D3268_, new_D3269_,
    new_D3270_, new_D3271_, new_D3272_, new_D3273_, new_D3274_, new_D3275_,
    new_D3276_, new_D3277_, new_D3278_, new_D3279_, new_D3280_, new_D3281_,
    new_D3282_, new_D3283_, new_D3284_, new_D3285_, new_D3286_, new_D3287_,
    new_D3288_, new_D3289_, new_D3290_, new_D3291_, new_D3292_, new_D3293_,
    new_D3294_, new_D3295_, new_D3296_, new_D3297_, new_D3298_, new_D3299_,
    new_D3300_, new_D3301_, new_D3302_, new_D3303_, new_D3304_, new_D3305_,
    new_D3306_, new_D3307_, new_D3308_, new_D3309_, new_D3310_, new_D3311_,
    new_D3312_, new_D3313_, new_D3314_, new_D3315_, new_D3316_, new_D3317_,
    new_D3318_, new_D3319_, new_D3320_, new_D3321_, new_D3322_, new_D3323_,
    new_D3324_, new_D3325_, new_D3326_, new_D3327_, new_D3328_, new_D3329_,
    new_D3330_, new_D3331_, new_D3332_, new_D3333_, new_D3334_, new_D3335_,
    new_D3336_, new_D3337_, new_D3338_, new_D3339_, new_D3340_, new_D3341_,
    new_D3342_, new_D3343_, new_D3344_, new_D3345_, new_D3346_, new_D3347_,
    new_D3348_, new_D3349_, new_D3350_, new_D3351_, new_D3352_, new_D3353_,
    new_D3354_, new_D3355_, new_D3356_, new_D3357_, new_D3358_, new_D3359_,
    new_D3360_, new_D3361_, new_D3362_, new_D3363_, new_D3364_, new_D3365_,
    new_D3366_, new_D3367_, new_D3368_, new_D3369_, new_D3370_, new_D3371_,
    new_D3372_, new_D3373_, new_D3374_, new_D3375_, new_D3376_, new_D3377_,
    new_D3378_, new_D3379_, new_D3380_, new_D3381_, new_D3382_, new_D3383_,
    new_D3384_, new_D3385_, new_D3386_, new_D3387_, new_D3388_, new_D3389_,
    new_D3390_, new_D3391_, new_D3392_, new_D3393_, new_D3394_, new_D3395_,
    new_D3396_, new_D3397_, new_D3398_, new_D3399_, new_D3400_, new_D3401_,
    new_D3402_, new_D3403_, new_D3404_, new_D3405_, new_D3406_, new_D3407_,
    new_D3408_, new_D3409_, new_D3410_, new_D3411_, new_D3412_, new_D3413_,
    new_D3414_, new_D3415_, new_D3416_, new_D3417_, new_D3418_, new_D3419_,
    new_D3420_, new_D3421_, new_D3422_, new_D3423_, new_D3424_, new_D3425_,
    new_D3426_, new_D3427_, new_D3428_, new_D3429_, new_D3430_, new_D3431_,
    new_D3432_, new_D3433_, new_D3434_, new_D3435_, new_D3436_, new_D3437_,
    new_D3438_, new_D3439_, new_D3440_, new_D3441_, new_D3442_, new_D3443_,
    new_D3444_, new_D3445_, new_D3446_, new_D3447_, new_D3448_, new_D3449_,
    new_D3450_, new_D3451_, new_D3452_, new_D3453_, new_D3454_, new_D3455_,
    new_D3456_, new_D3457_, new_D3458_, new_D3459_, new_D3460_, new_D3461_,
    new_D3462_, new_D3463_, new_D3464_, new_D3465_, new_D3466_, new_D3467_,
    new_D3468_, new_D3469_, new_D3470_, new_D3471_, new_D3472_, new_D3473_,
    new_D3474_, new_D3475_, new_D3476_, new_D3477_, new_D3478_, new_D3479_,
    new_D3480_, new_D3481_, new_D3482_, new_D3483_, new_D3484_, new_D3485_,
    new_D3486_, new_D3487_, new_D3488_, new_D3489_, new_D3490_, new_D3491_,
    new_D3492_, new_D3493_, new_D3494_, new_D3495_, new_D3496_, new_D3497_,
    new_D3498_, new_D3499_, new_D3500_, new_D3501_, new_D3502_, new_D3503_,
    new_D3504_, new_D3505_, new_D3506_, new_D3507_, new_D3508_, new_D3509_,
    new_D3510_, new_D3511_, new_D3512_, new_D3513_, new_D3514_, new_D3515_,
    new_D3516_, new_D3517_, new_D3518_, new_D3519_, new_D3520_, new_D3521_,
    new_D3522_, new_D3523_, new_D3524_, new_D3525_, new_D3526_, new_D3527_,
    new_D3528_, new_D3529_, new_D3530_, new_D3531_, new_D3532_, new_D3533_,
    new_D3534_, new_D3535_, new_D3536_, new_D3537_, new_D3538_, new_D3539_,
    new_D3540_, new_D3541_, new_D3542_, new_D3543_, new_D3544_, new_D3545_,
    new_D3546_, new_D3547_, new_D3548_, new_D3549_, new_D3550_, new_D3551_,
    new_D3552_, new_D3553_, new_D3554_, new_D3555_, new_D3556_, new_D3557_,
    new_D3558_, new_D3559_, new_D3560_, new_D3561_, new_D3562_, new_D3563_,
    new_D3564_, new_D3565_, new_D3566_, new_D3567_, new_D3568_, new_D3569_,
    new_D3570_, new_D3571_, new_D3572_, new_D3573_, new_D3574_, new_D3575_,
    new_D3576_, new_D3577_, new_D3578_, new_D3579_, new_D3580_, new_D3581_,
    new_D3582_, new_D3583_, new_D3584_, new_D3585_, new_D3586_, new_D3587_,
    new_D3588_, new_D3589_, new_D3590_, new_D3591_, new_D3592_, new_D3593_,
    new_D3594_, new_D3595_, new_D3596_, new_D3597_, new_D3598_, new_D3599_,
    new_D3600_, new_D3601_, new_D3602_, new_D3603_, new_D3604_, new_D3605_,
    new_D3606_, new_D3607_, new_D3608_, new_D3609_, new_D3610_, new_D3611_,
    new_D3612_, new_D3613_, new_D3614_, new_D3615_, new_D3616_, new_D3617_,
    new_D3618_, new_D3619_, new_D3620_, new_D3621_, new_D3622_, new_D3623_,
    new_D3624_, new_D3625_, new_D3626_, new_D3627_, new_D3628_, new_D3629_,
    new_D3630_, new_D3631_, new_D3632_, new_D3633_, new_D3634_, new_D3635_,
    new_D3636_, new_D3637_, new_D3638_, new_D3639_, new_D3640_, new_D3641_,
    new_D3642_, new_D3643_, new_D3644_, new_D3645_, new_D3646_, new_D3647_,
    new_D3648_, new_D3649_, new_D3650_, new_D3651_, new_D3652_, new_D3653_,
    new_D3654_, new_D3655_, new_D3656_, new_D3657_, new_D3658_, new_D3659_,
    new_D3660_, new_D3661_, new_D3662_, new_D3663_, new_D3664_, new_D3665_,
    new_D3666_, new_D3667_, new_D3668_, new_D3669_, new_D3670_, new_D3671_,
    new_D3672_, new_D3673_, new_D3674_, new_D3675_, new_D3676_, new_D3677_,
    new_D3678_, new_D3679_, new_D3680_, new_D3681_, new_D3682_, new_D3683_,
    new_D3684_, new_D3685_, new_D3686_, new_D3687_, new_D3688_, new_D3689_,
    new_D3690_, new_D3691_, new_D3692_, new_D3693_, new_D3694_, new_D3695_,
    new_D3696_, new_D3697_, new_D3698_, new_D3699_, new_D3700_, new_D3701_,
    new_D3702_, new_D3703_, new_D3704_, new_D3705_, new_D3706_, new_D3707_,
    new_D3708_, new_D3709_, new_D3710_, new_D3711_, new_D3712_, new_D3713_,
    new_D3714_, new_D3715_, new_D3716_, new_D3717_, new_D3718_, new_D3719_,
    new_D3720_, new_D3721_, new_D3722_, new_D3723_, new_D3724_, new_D3725_,
    new_D3726_, new_D3727_, new_D3728_, new_D3729_, new_D3730_, new_D3731_,
    new_D3732_, new_D3733_, new_D3734_, new_D3735_, new_D3736_, new_D3737_,
    new_D3738_, new_D3739_, new_D3740_, new_D3741_, new_D3742_, new_D3743_,
    new_D3744_, new_D3745_, new_D3746_, new_D3747_, new_D3748_, new_D3749_,
    new_D3750_, new_D3751_, new_D3752_, new_D3753_, new_D3754_, new_D3755_,
    new_D3756_, new_D3757_, new_D3758_, new_D3759_, new_D3760_, new_D3761_,
    new_D3762_, new_D3763_, new_D3764_, new_D3765_, new_D3766_, new_D3767_,
    new_D3768_, new_D3769_, new_D3770_, new_D3771_, new_D3772_, new_D3773_,
    new_D3774_, new_D3775_, new_D3776_, new_D3777_, new_D3778_, new_D3779_,
    new_D3780_, new_D3781_, new_D3782_, new_D3783_, new_D3784_, new_D3785_,
    new_D3786_, new_D3787_, new_D3788_, new_D3789_, new_D3790_, new_D3791_,
    new_D3792_, new_D3793_, new_D3794_, new_D3795_, new_D3796_, new_D3797_,
    new_D3798_, new_D3799_, new_D3800_, new_D3801_, new_D3802_, new_D3803_,
    new_D3804_, new_D3805_, new_D3806_, new_D3807_, new_D3808_, new_D3809_,
    new_D3810_, new_D3811_, new_D3812_, new_D3813_, new_D3814_, new_D3815_,
    new_D3816_, new_D3817_, new_D3818_, new_D3819_, new_D3820_, new_D3821_,
    new_D3822_, new_D3823_, new_D3824_, new_D3825_, new_D3826_, new_D3827_,
    new_D3828_, new_D3829_, new_D3830_, new_D3831_, new_D3832_, new_D3833_,
    new_D3834_, new_D3835_, new_D3836_, new_D3837_, new_D3838_, new_D3839_,
    new_D3840_, new_D3841_, new_D3842_, new_D3843_, new_D3844_, new_D3845_,
    new_D3846_, new_D3847_, new_D3848_, new_D3849_, new_D3850_, new_D3851_,
    new_D3852_, new_D3853_, new_D3854_, new_D3855_, new_D3856_, new_D3857_,
    new_D3858_, new_D3859_, new_D3860_, new_D3861_, new_D3862_, new_D3863_,
    new_D3864_, new_D3865_, new_D3866_, new_D3867_, new_D3868_, new_D3869_,
    new_D3870_, new_D3871_, new_D3872_, new_D3873_, new_D3874_, new_D3875_,
    new_D3876_, new_D3877_, new_D3878_, new_D3879_, new_D3880_, new_D3881_,
    new_D3882_, new_D3883_, new_D3884_, new_D3885_, new_D3886_, new_D3887_,
    new_D3888_, new_D3889_, new_D3890_, new_D3891_, new_D3892_, new_D3893_,
    new_D3894_, new_D3895_, new_D3896_, new_D3897_, new_D3898_, new_D3899_,
    new_D3900_, new_D3901_, new_D3902_, new_D3903_, new_D3904_, new_D3905_,
    new_D3906_, new_D3907_, new_D3908_, new_D3909_, new_D3910_, new_D3911_,
    new_D3912_, new_D3913_, new_D3914_, new_D3915_, new_D3916_, new_D3917_,
    new_D3918_, new_D3919_, new_D3920_, new_D3921_, new_D3922_, new_D3923_,
    new_D3924_, new_D3925_, new_D3926_, new_D3927_, new_D3928_, new_D3929_,
    new_D3930_, new_D3931_, new_D3932_, new_D3933_, new_D3934_, new_D3935_,
    new_D3936_, new_D3937_, new_D3938_, new_D3939_, new_D3940_, new_D3941_,
    new_D3942_, new_D3943_, new_D3944_, new_D3945_, new_D3946_, new_D3947_,
    new_D3948_, new_D3949_, new_D3950_, new_D3951_, new_D3952_, new_D3953_,
    new_D3954_, new_D3955_, new_D3956_, new_D3957_, new_D3958_, new_D3959_,
    new_D3960_, new_D3961_, new_D3962_, new_D3963_, new_D3964_, new_D3965_,
    new_D3966_, new_D3967_, new_D3968_, new_D3969_, new_D3970_, new_D3971_,
    new_D3972_, new_D3973_, new_D3974_, new_D3975_, new_D3976_, new_D3977_,
    new_D3978_, new_D3979_, new_D3980_, new_D3981_, new_D3982_, new_D3983_,
    new_D3984_, new_D3985_, new_D3986_, new_D3987_, new_D3988_, new_D3989_,
    new_D3990_, new_D3991_, new_D3992_, new_D3993_, new_D3994_, new_D3995_,
    new_D3996_, new_D3997_, new_D3998_, new_D3999_, new_D4000_, new_D4001_,
    new_D4002_, new_D4003_, new_D4004_, new_D4005_, new_D4006_, new_D4007_,
    new_D4008_, new_D4009_, new_D4010_, new_D4011_, new_D4012_, new_D4013_,
    new_D4014_, new_D4015_, new_D4016_, new_D4017_, new_D4018_, new_D4019_,
    new_D4020_, new_D4021_, new_D4022_, new_D4023_, new_D4024_, new_D4025_,
    new_D4026_, new_D4027_, new_D4028_, new_D4029_, new_D4030_, new_D4031_,
    new_D4032_, new_D4033_, new_D4034_, new_D4035_, new_D4036_, new_D4037_,
    new_D4038_, new_D4039_, new_D4040_, new_D4041_, new_D4042_, new_D4043_,
    new_D4044_, new_D4045_, new_D4046_, new_D4047_, new_D4048_, new_D4049_,
    new_D4050_, new_D4051_, new_D4052_, new_D4053_, new_D4054_, new_D4055_,
    new_D4056_, new_D4057_, new_D4058_, new_D4059_, new_D4060_, new_D4061_,
    new_D4062_, new_D4063_, new_D4064_, new_D4065_, new_D4066_, new_D4067_,
    new_D4068_, new_D4069_, new_D4070_, new_D4071_, new_D4072_, new_D4073_,
    new_D4074_, new_D4075_, new_D4076_, new_D4077_, new_D4078_, new_D4079_,
    new_D4080_, new_D4081_, new_D4082_, new_D4083_, new_D4084_, new_D4085_,
    new_D4086_, new_D4087_, new_D4088_, new_D4089_, new_D4090_, new_D4091_,
    new_D4092_, new_D4093_, new_D4094_, new_D4095_, new_D4096_, new_D4097_,
    new_D4098_, new_D4099_, new_D4100_, new_D4101_, new_D4102_, new_D4103_,
    new_D4104_, new_D4105_, new_D4106_, new_D4107_, new_D4108_, new_D4109_,
    new_D4110_, new_D4111_, new_D4112_, new_D4113_, new_D4114_, new_D4115_,
    new_D4116_, new_D4117_, new_D4118_, new_D4119_, new_D4120_, new_D4121_,
    new_D4122_, new_D4123_, new_D4124_, new_D4125_, new_D4126_, new_D4127_,
    new_D4128_, new_D4129_, new_D4130_, new_D4131_, new_D4132_, new_D4133_,
    new_D4134_, new_D4135_, new_D4136_, new_D4137_, new_D4138_, new_D4139_,
    new_D4140_, new_D4141_, new_D4142_, new_D4143_, new_D4144_, new_D4145_,
    new_D4146_, new_D4147_, new_D4148_, new_D4149_, new_D4150_, new_D4151_,
    new_D4152_, new_D4153_, new_D4154_, new_D4155_, new_D4156_, new_D4157_,
    new_D4158_, new_D4159_, new_D4160_, new_D4161_, new_D4162_, new_D4163_,
    new_D4164_, new_D4165_, new_D4166_, new_D4167_, new_D4168_, new_D4169_,
    new_D4170_, new_D4171_, new_D4172_, new_D4173_, new_D4174_, new_D4175_,
    new_D4176_, new_D4177_, new_D4178_, new_D4179_, new_D4180_, new_D4181_,
    new_D4182_, new_D4183_, new_D4184_, new_D4185_, new_D4186_, new_D4187_,
    new_D4188_, new_D4189_, new_D4190_, new_D4191_, new_D4192_, new_D4193_,
    new_D4194_, new_D4195_, new_D4196_, new_D4197_, new_D4198_, new_D4199_,
    new_D4200_, new_D4201_, new_D4202_, new_D4203_, new_D4204_, new_D4205_,
    new_D4206_, new_D4207_, new_D4208_, new_D4209_, new_D4210_, new_D4211_,
    new_D4212_, new_D4213_, new_D4214_, new_D4215_, new_D4216_, new_D4217_,
    new_D4218_, new_D4219_, new_D4220_, new_D4221_, new_D4222_, new_D4223_,
    new_D4224_, new_D4225_, new_D4226_, new_D4227_, new_D4228_, new_D4229_,
    new_D4230_, new_D4231_, new_D4232_, new_D4233_, new_D4234_, new_D4235_,
    new_D4236_, new_D4237_, new_D4238_, new_D4239_, new_D4240_, new_D4241_,
    new_D4242_, new_D4243_, new_D4244_, new_D4245_, new_D4246_, new_D4247_,
    new_D4248_, new_D4249_, new_D4250_, new_D4251_, new_D4252_, new_D4253_,
    new_D4254_, new_D4255_, new_D4256_, new_D4257_, new_D4258_, new_D4259_,
    new_D4260_, new_D4261_, new_D4262_, new_D4263_, new_D4264_, new_D4265_,
    new_D4266_, new_D4267_, new_D4268_, new_D4269_, new_D4270_, new_D4271_,
    new_D4272_, new_D4273_, new_D4274_, new_D4275_, new_D4276_, new_D4277_,
    new_D4278_, new_D4279_, new_D4280_, new_D4281_, new_D4282_, new_D4283_,
    new_D4284_, new_D4285_, new_D4286_, new_D4287_, new_D4288_, new_D4289_,
    new_D4290_, new_D4291_, new_D4292_, new_D4293_, new_D4294_, new_D4295_,
    new_D4296_, new_D4297_, new_D4298_, new_D4299_, new_D4300_, new_D4301_,
    new_D4302_, new_D4303_, new_D4304_, new_D4305_, new_D4306_, new_D4307_,
    new_D4308_, new_D4309_, new_D4310_, new_D4311_, new_D4312_, new_D4313_,
    new_D4314_, new_D4315_, new_D4316_, new_D4317_, new_D4318_, new_D4319_,
    new_D4320_, new_D4321_, new_D4322_, new_D4323_, new_D4324_, new_D4325_,
    new_D4326_, new_D4327_, new_D4328_, new_D4329_, new_D4330_, new_D4331_,
    new_D4332_, new_D4333_, new_D4334_, new_D4335_, new_D4336_, new_D4337_,
    new_D4338_, new_D4339_, new_D4340_, new_D4341_, new_D4342_, new_D4343_,
    new_D4344_, new_D4345_, new_D4346_, new_D4347_, new_D4348_, new_D4349_,
    new_D4350_, new_D4351_, new_D4352_, new_D4353_, new_D4354_, new_D4355_,
    new_D4356_, new_D4357_, new_D4358_, new_D4359_, new_D4360_, new_D4361_,
    new_D4362_, new_D4363_, new_D4364_, new_D4365_, new_D4366_, new_D4367_,
    new_D4368_, new_D4369_, new_D4370_, new_D4371_, new_D4372_, new_D4373_,
    new_D4374_, new_D4375_, new_D4376_, new_D4377_, new_D4378_, new_D4379_,
    new_D4380_, new_D4381_, new_D4382_, new_D4383_, new_D4384_, new_D4385_,
    new_D4386_, new_D4387_, new_D4388_, new_D4389_, new_D4390_, new_D4391_,
    new_D4392_, new_D4393_, new_D4394_, new_D4395_, new_D4396_, new_D4397_,
    new_D4398_, new_D4399_, new_D4400_, new_D4401_, new_D4402_, new_D4403_,
    new_D4404_, new_D4405_, new_D4406_, new_D4407_, new_D4408_, new_D4409_,
    new_D4410_, new_D4411_, new_D4412_, new_D4413_, new_D4414_, new_D4415_,
    new_D4416_, new_D4417_, new_D4418_, new_D4419_, new_D4420_, new_D4421_,
    new_D4422_, new_D4423_, new_D4424_, new_D4425_, new_D4426_, new_D4427_,
    new_D4428_, new_D4429_, new_D4430_, new_D4431_, new_D4432_, new_D4433_,
    new_D4434_, new_D4435_, new_D4436_, new_D4437_, new_D4438_, new_D4439_,
    new_D4440_, new_D4441_, new_D4442_, new_D4443_, new_D4444_, new_D4445_,
    new_D4446_, new_D4447_, new_D4448_, new_D4449_, new_D4450_, new_D4451_,
    new_D4452_, new_D4453_, new_D4454_, new_D4455_, new_D4456_, new_D4457_,
    new_D4458_, new_D4459_, new_D4460_, new_D4461_, new_D4462_, new_D4463_,
    new_D4464_, new_D4465_, new_D4466_, new_D4467_, new_D4468_, new_D4469_,
    new_D4470_, new_D4471_, new_D4472_, new_D4473_, new_D4474_, new_D4475_,
    new_D4476_, new_D4477_, new_D4478_, new_D4479_, new_D4480_, new_D4481_,
    new_D4482_, new_D4483_, new_D4484_, new_D4485_, new_D4486_, new_D4487_,
    new_D4488_, new_D4489_, new_D4490_, new_D4491_, new_D4492_, new_D4493_,
    new_D4494_, new_D4495_, new_D4496_, new_D4497_, new_D4498_, new_D4499_,
    new_D4500_, new_D4501_, new_D4502_, new_D4503_, new_D4504_, new_D4505_,
    new_D4506_, new_D4507_, new_D4508_, new_D4509_, new_D4510_, new_D4511_,
    new_D4512_, new_D4513_, new_D4514_, new_D4515_, new_D4516_, new_D4517_,
    new_D4518_, new_D4519_, new_D4520_, new_D4521_, new_D4522_, new_D4523_,
    new_D4524_, new_D4525_, new_D4526_, new_D4527_, new_D4528_, new_D4529_,
    new_D4530_, new_D4531_, new_D4532_, new_D4533_, new_D4534_, new_D4535_,
    new_D4536_, new_D4537_, new_D4538_, new_D4539_, new_D4540_, new_D4541_,
    new_D4542_, new_D4543_, new_D4544_, new_D4545_, new_D4546_, new_D4547_,
    new_D4548_, new_D4549_, new_D4550_, new_D4551_, new_D4552_, new_D4553_,
    new_D4554_, new_D4555_, new_D4556_, new_D4557_, new_D4558_, new_D4559_,
    new_D4560_, new_D4561_, new_D4562_, new_D4563_, new_D4564_, new_D4565_,
    new_D4566_, new_D4567_, new_D4568_, new_D4569_, new_D4570_, new_D4571_,
    new_D4572_, new_D4573_, new_D4574_, new_D4575_, new_D4576_, new_D4577_,
    new_D4578_, new_D4579_, new_D4580_, new_D4581_, new_D4582_, new_D4583_,
    new_D4584_, new_D4585_, new_D4586_, new_D4587_, new_D4588_, new_D4589_,
    new_D4590_, new_D4591_, new_D4592_, new_D4593_, new_D4594_, new_D4595_,
    new_D4596_, new_D4597_, new_D4598_, new_D4599_, new_D4600_, new_D4601_,
    new_D4602_, new_D4603_, new_D4604_, new_D4605_, new_D4606_, new_D4607_,
    new_D4608_, new_D4609_, new_D4610_, new_D4611_, new_D4612_, new_D4613_,
    new_D4614_, new_D4615_, new_D4616_, new_D4617_, new_D4618_, new_D4619_,
    new_D4620_, new_D4621_, new_D4622_, new_D4623_, new_D4624_, new_D4625_,
    new_D4626_, new_D4627_, new_D4628_, new_D4629_, new_D4630_, new_D4631_,
    new_D4632_, new_D4633_, new_D4634_, new_D4635_, new_D4636_, new_D4637_,
    new_D4638_, new_D4639_, new_D4640_, new_D4641_, new_D4642_, new_D4643_,
    new_D4644_, new_D4645_, new_D4646_, new_D4647_, new_D4648_, new_D4649_,
    new_D4650_, new_D4651_, new_D4652_, new_D4653_, new_D4654_, new_D4655_,
    new_D4656_, new_D4657_, new_D4658_, new_D4659_, new_D4660_, new_D4661_,
    new_D4662_, new_D4663_, new_D4664_, new_D4665_, new_D4666_, new_D4667_,
    new_D4668_, new_D4669_, new_D4670_, new_D4671_, new_D4672_, new_D4673_,
    new_D4674_, new_D4675_, new_D4676_, new_D4677_, new_D4678_, new_D4679_,
    new_D4680_, new_D4681_, new_D4682_, new_D4683_, new_D4684_, new_D4685_,
    new_D4686_, new_D4687_, new_D4688_, new_D4689_, new_D4690_, new_D4691_,
    new_D4692_, new_D4693_, new_D4694_, new_D4695_, new_D4696_, new_D4697_,
    new_D4698_, new_D4699_, new_D4700_, new_D4701_, new_D4702_, new_D4703_,
    new_D4704_, new_D4705_, new_D4706_, new_D4707_, new_D4708_, new_D4709_,
    new_D4710_, new_D4711_, new_D4712_, new_D4713_, new_D4714_, new_D4715_,
    new_D4716_, new_D4717_, new_D4718_, new_D4719_, new_D4720_, new_D4721_,
    new_D4722_, new_D4723_, new_D4724_, new_D4725_, new_D4726_, new_D4727_,
    new_D4728_, new_D4729_, new_D4730_, new_D4731_, new_D4732_, new_D4733_,
    new_D4734_, new_D4735_, new_D4736_, new_D4737_, new_D4738_, new_D4739_,
    new_D4740_, new_D4741_, new_D4742_, new_D4743_, new_D4744_, new_D4745_,
    new_D4746_, new_D4747_, new_D4748_, new_D4749_, new_D4750_, new_D4751_,
    new_D4752_, new_D4753_, new_D4754_, new_D4755_, new_D4756_, new_D4757_,
    new_D4758_, new_D4759_, new_D4760_, new_D4761_, new_D4762_, new_D4763_,
    new_D4764_, new_D4765_, new_D4766_, new_D4767_, new_D4768_, new_D4769_,
    new_D4770_, new_D4771_, new_D4772_, new_D4773_, new_D4774_, new_D4775_,
    new_D4776_, new_D4777_, new_D4778_, new_D4779_, new_D4780_, new_D4781_,
    new_D4782_, new_D4783_, new_D4784_, new_D4785_, new_D4786_, new_D4787_,
    new_D4788_, new_D4789_, new_D4790_, new_D4791_, new_D4792_, new_D4793_,
    new_D4794_, new_D4795_, new_D4796_, new_D4797_, new_D4798_, new_D4799_,
    new_D4800_, new_D4801_, new_D4802_, new_D4803_, new_D4804_, new_D4805_,
    new_D4806_, new_D4807_, new_D4808_, new_D4809_, new_D4810_, new_D4811_,
    new_D4812_, new_D4813_, new_D4814_, new_D4815_, new_D4816_, new_D4817_,
    new_D4818_, new_D4819_, new_D4820_, new_D4821_, new_D4822_, new_D4823_,
    new_D4824_, new_D4825_, new_D4826_, new_D4827_, new_D4828_, new_D4829_,
    new_D4830_, new_D4831_, new_D4832_, new_D4833_, new_D4834_, new_D4835_,
    new_D4836_, new_D4837_, new_D4838_, new_D4839_, new_D4840_, new_D4841_,
    new_D4842_, new_D4843_, new_D4844_, new_D4845_, new_D4846_, new_D4847_,
    new_D4848_, new_D4849_, new_D4850_, new_D4851_, new_D4852_, new_D4853_,
    new_D4854_, new_D4855_, new_D4856_, new_D4857_, new_D4858_, new_D4859_,
    new_D4860_, new_D4861_, new_D4862_, new_D4863_, new_D4864_, new_D4865_,
    new_D4866_, new_D4867_, new_D4868_, new_D4869_, new_D4870_, new_D4871_,
    new_D4872_, new_D4873_, new_D4874_, new_D4875_, new_D4876_, new_D4877_,
    new_D4878_, new_D4879_, new_D4880_, new_D4881_, new_D4882_, new_D4883_,
    new_D4884_, new_D4885_, new_D4886_, new_D4887_, new_D4888_, new_D4889_,
    new_D4890_, new_D4891_, new_D4892_, new_D4893_, new_D4894_, new_D4895_,
    new_D4896_, new_D4897_, new_D4898_, new_D4899_, new_D4900_, new_D4901_,
    new_D4902_, new_D4903_, new_D4904_, new_D4905_, new_D4906_, new_D4907_,
    new_D4908_, new_D4909_, new_D4910_, new_D4911_, new_D4912_, new_D4913_,
    new_D4914_, new_D4915_, new_D4916_, new_D4917_, new_D4918_, new_D4919_,
    new_D4920_, new_D4921_, new_D4922_, new_D4923_, new_D4924_, new_D4925_,
    new_D4926_, new_D4927_, new_D4928_, new_D4929_, new_D4930_, new_D4931_,
    new_D4932_, new_D4933_, new_D4934_, new_D4935_, new_D4936_, new_D4937_,
    new_D4938_, new_D4939_, new_D4940_, new_D4941_, new_D4942_, new_D4943_,
    new_D4944_, new_D4945_, new_D4946_, new_D4947_, new_D4948_, new_D4949_,
    new_D4950_, new_D4951_, new_D4952_, new_D4953_, new_D4954_, new_D4955_,
    new_D4956_, new_D4957_, new_D4958_, new_D4959_, new_D4960_, new_D4961_,
    new_D4962_, new_D4963_, new_D4964_, new_D4965_, new_D4966_, new_D4967_,
    new_D4968_, new_D4969_, new_D4970_, new_D4971_, new_D4972_, new_D4973_,
    new_D4974_, new_D4975_, new_D4976_, new_D4977_, new_D4978_, new_D4979_,
    new_D4980_, new_D4981_, new_D4982_, new_D4983_, new_D4984_, new_D4985_,
    new_D4986_, new_D4987_, new_D4988_, new_D4989_, new_D4990_, new_D4991_,
    new_D4992_, new_D4993_, new_D4994_, new_D4995_, new_D4996_, new_D4997_,
    new_D4998_, new_D4999_, new_D5000_, new_D5001_, new_D5002_, new_D5003_,
    new_D5004_, new_D5005_, new_D5006_, new_D5007_, new_D5008_, new_D5009_,
    new_D5010_, new_D5011_, new_D5012_, new_D5013_, new_D5014_, new_D5015_,
    new_D5016_, new_D5017_, new_D5018_, new_D5019_, new_D5020_, new_D5021_,
    new_D5022_, new_D5023_, new_D5024_, new_D5025_, new_D5026_, new_D5027_,
    new_D5028_, new_D5029_, new_D5030_, new_D5031_, new_D5032_, new_D5033_,
    new_D5034_, new_D5035_, new_D5036_, new_D5037_, new_D5038_, new_D5039_,
    new_D5040_, new_D5041_, new_D5042_, new_D5043_, new_D5044_, new_D5045_,
    new_D5046_, new_D5047_, new_D5048_, new_D5049_, new_D5050_, new_D5051_,
    new_D5052_, new_D5053_, new_D5054_, new_D5055_, new_D5056_, new_D5057_,
    new_D5058_, new_D5059_, new_D5060_, new_D5061_, new_D5062_, new_D5063_,
    new_D5064_, new_D5065_, new_D5066_, new_D5067_, new_D5068_, new_D5069_,
    new_D5070_, new_D5071_, new_D5072_, new_D5073_, new_D5074_, new_D5075_,
    new_D5076_, new_D5077_, new_D5078_, new_D5079_, new_D5080_, new_D5081_,
    new_D5082_, new_D5083_, new_D5084_, new_D5085_, new_D5086_, new_D5087_,
    new_D5088_, new_D5089_, new_D5090_, new_D5091_, new_D5092_, new_D5093_,
    new_D5094_, new_D5095_, new_D5096_, new_D5097_, new_D5098_, new_D5099_,
    new_D5100_, new_D5101_, new_D5102_, new_D5103_, new_D5104_, new_D5105_,
    new_D5106_, new_D5107_, new_D5108_, new_D5109_, new_D5110_, new_D5111_,
    new_D5112_, new_D5113_, new_D5114_, new_D5115_, new_D5116_, new_D5117_,
    new_D5118_, new_D5119_, new_D5120_, new_D5121_, new_D5122_, new_D5123_,
    new_D5124_, new_D5125_, new_D5126_, new_D5127_, new_D5128_, new_D5129_,
    new_D5130_, new_D5131_, new_D5132_, new_D5133_, new_D5134_, new_D5135_,
    new_D5136_, new_D5137_, new_D5138_, new_D5139_, new_D5140_, new_D5141_,
    new_D5142_, new_D5143_, new_D5144_, new_D5145_, new_D5146_, new_D5147_,
    new_D5148_, new_D5149_, new_D5150_, new_D5151_, new_D5152_, new_D5153_,
    new_D5154_, new_D5155_, new_D5156_, new_D5157_, new_D5158_, new_D5159_,
    new_D5160_, new_D5161_, new_D5162_, new_D5163_, new_D5164_, new_D5165_,
    new_D5166_, new_D5167_, new_D5168_, new_D5169_, new_D5170_, new_D5171_,
    new_D5172_, new_D5173_, new_D5174_, new_D5175_, new_D5176_, new_D5177_,
    new_D5178_, new_D5179_, new_D5180_, new_D5181_, new_D5182_, new_D5183_,
    new_D5184_, new_D5185_, new_D5186_, new_D5187_, new_D5188_, new_D5189_,
    new_D5190_, new_D5191_, new_D5192_, new_D5193_, new_D5194_, new_D5195_,
    new_D5196_, new_D5197_, new_D5198_, new_D5199_, new_D5200_, new_D5201_,
    new_D5202_, new_D5203_, new_D5204_, new_D5205_, new_D5206_, new_D5207_,
    new_D5208_, new_D5209_, new_D5210_, new_D5211_, new_D5212_, new_D5213_,
    new_D5214_, new_D5215_, new_D5216_, new_D5217_, new_D5218_, new_D5219_,
    new_D5220_, new_D5221_, new_D5222_, new_D5223_, new_D5224_, new_D5225_,
    new_D5226_, new_D5227_, new_D5228_, new_D5229_, new_D5230_, new_D5231_,
    new_D5232_, new_D5233_, new_D5234_, new_D5235_, new_D5236_, new_D5237_,
    new_D5238_, new_D5239_, new_D5240_, new_D5241_, new_D5242_, new_D5243_,
    new_D5244_, new_D5245_, new_D5246_, new_D5247_, new_D5248_, new_D5249_,
    new_D5250_, new_D5251_, new_D5252_, new_D5253_, new_D5254_, new_D5255_,
    new_D5256_, new_D5257_, new_D5258_, new_D5259_, new_D5260_, new_D5261_,
    new_D5262_, new_D5263_, new_D5264_, new_D5265_, new_D5266_, new_D5267_,
    new_D5268_, new_D5269_, new_D5270_, new_D5271_, new_D5272_, new_D5273_,
    new_D5274_, new_D5275_, new_D5276_, new_D5277_, new_D5278_, new_D5279_,
    new_D5280_, new_D5281_, new_D5282_, new_D5283_, new_D5284_, new_D5285_,
    new_D5286_, new_D5287_, new_D5288_, new_D5289_, new_D5290_, new_D5291_,
    new_D5292_, new_D5293_, new_D5294_, new_D5295_, new_D5296_, new_D5297_,
    new_D5298_, new_D5299_, new_D5300_, new_D5301_, new_D5302_, new_D5303_,
    new_D5304_, new_D5305_, new_D5306_, new_D5307_, new_D5308_, new_D5309_,
    new_D5310_, new_D5311_, new_D5312_, new_D5313_, new_D5314_, new_D5315_,
    new_D5316_, new_D5317_, new_D5318_, new_D5319_, new_D5320_, new_D5321_,
    new_D5322_, new_D5323_, new_D5324_, new_D5325_, new_D5326_, new_D5327_,
    new_D5328_, new_D5329_, new_D5330_, new_D5331_, new_D5332_, new_D5333_,
    new_D5334_, new_D5335_, new_D5336_, new_D5337_, new_D5338_, new_D5339_,
    new_D5340_, new_D5341_, new_D5342_, new_D5343_, new_D5344_, new_D5345_,
    new_D5346_, new_D5347_, new_D5348_, new_D5349_, new_D5350_, new_D5351_,
    new_D5352_, new_D5353_, new_D5354_, new_D5355_, new_D5356_, new_D5357_,
    new_D5358_, new_D5359_, new_D5360_, new_D5361_, new_D5362_, new_D5363_,
    new_D5364_, new_D5365_, new_D5366_, new_D5367_, new_D5368_, new_D5369_,
    new_D5370_, new_D5371_, new_D5372_, new_D5373_, new_D5374_, new_D5375_,
    new_D5376_, new_D5377_, new_D5378_, new_D5379_, new_D5380_, new_D5381_,
    new_D5382_, new_D5383_, new_D5384_, new_D5385_, new_D5386_, new_D5387_,
    new_D5388_, new_D5389_, new_D5390_, new_D5391_, new_D5392_, new_D5393_,
    new_D5394_, new_D5395_, new_D5396_, new_D5397_, new_D5398_, new_D5399_,
    new_D5400_, new_D5401_, new_D5402_, new_D5403_, new_D5404_, new_D5405_,
    new_D5406_, new_D5407_, new_D5408_, new_D5409_, new_D5410_, new_D5411_,
    new_D5412_, new_D5413_, new_D5414_, new_D5415_, new_D5416_, new_D5417_,
    new_D5418_, new_D5419_, new_D5420_, new_D5421_, new_D5422_, new_D5423_,
    new_D5424_, new_D5425_, new_D5426_, new_D5427_, new_D5428_, new_D5429_,
    new_D5430_, new_D5431_, new_D5432_, new_D5433_, new_D5434_, new_D5435_,
    new_D5436_, new_D5437_, new_D5438_, new_D5439_, new_D5440_, new_D5441_,
    new_D5442_, new_D5443_, new_D5444_, new_D5445_, new_D5446_, new_D5447_,
    new_D5448_, new_D5449_, new_D5450_, new_D5451_, new_D5452_, new_D5453_,
    new_D5454_, new_D5455_, new_D5456_, new_D5457_, new_D5458_, new_D5459_,
    new_D5460_, new_D5461_, new_D5462_, new_D5463_, new_D5464_, new_D5465_,
    new_D5466_, new_D5467_, new_D5468_, new_D5469_, new_D5470_, new_D5471_,
    new_D5472_, new_D5473_, new_D5474_, new_D5475_, new_D5476_, new_D5477_,
    new_D5478_, new_D5479_, new_D5480_, new_D5481_, new_D5482_, new_D5483_,
    new_D5484_, new_D5485_, new_D5486_, new_D5487_, new_D5488_, new_D5489_,
    new_D5490_, new_D5491_, new_D5492_, new_D5493_, new_D5494_, new_D5495_,
    new_D5496_, new_D5497_, new_D5498_, new_D5499_, new_D5500_, new_D5501_,
    new_D5502_, new_D5503_, new_D5504_, new_D5505_, new_D5506_, new_D5507_,
    new_D5508_, new_D5509_, new_D5510_, new_D5511_, new_D5512_, new_D5513_,
    new_D5514_, new_D5515_, new_D5516_, new_D5517_, new_D5518_, new_D5519_,
    new_D5520_, new_D5521_, new_D5522_, new_D5523_, new_D5524_, new_D5525_,
    new_D5526_, new_D5527_, new_D5528_, new_D5529_, new_D5530_, new_D5531_,
    new_D5532_, new_D5533_, new_D5534_, new_D5535_, new_D5536_, new_D5537_,
    new_D5538_, new_D5539_, new_D5540_, new_D5541_, new_D5542_, new_D5543_,
    new_D5544_, new_D5545_, new_D5546_, new_D5547_, new_D5548_, new_D5549_,
    new_D5550_, new_D5551_, new_D5552_, new_D5553_, new_D5554_, new_D5555_,
    new_D5556_, new_D5557_, new_D5558_, new_D5559_, new_D5560_, new_D5561_,
    new_D5562_, new_D5563_, new_D5564_, new_D5565_, new_D5566_, new_D5567_,
    new_D5568_, new_D5569_, new_D5570_, new_D5571_, new_D5572_, new_D5573_,
    new_D5574_, new_D5575_, new_D5576_, new_D5577_, new_D5578_, new_D5579_,
    new_D5580_, new_D5581_, new_D5582_, new_D5583_, new_D5584_, new_D5585_,
    new_D5586_, new_D5587_, new_D5588_, new_D5589_, new_D5590_, new_D5591_,
    new_D5592_, new_D5593_, new_D5594_, new_D5595_, new_D5596_, new_D5597_,
    new_D5598_, new_D5599_, new_D5600_, new_D5601_, new_D5602_, new_D5603_,
    new_D5604_, new_D5605_, new_D5606_, new_D5607_, new_D5608_, new_D5609_,
    new_D5610_, new_D5611_, new_D5612_, new_D5613_, new_D5614_, new_D5615_,
    new_D5616_, new_D5617_, new_D5618_, new_D5619_, new_D5620_, new_D5621_,
    new_D5622_, new_D5623_, new_D5624_, new_D5625_, new_D5626_, new_D5627_,
    new_D5628_, new_D5629_, new_D5630_, new_D5631_, new_D5632_, new_D5633_,
    new_D5634_, new_D5635_, new_D5636_, new_D5637_, new_D5638_, new_D5639_,
    new_D5640_, new_D5641_, new_D5642_, new_D5643_, new_D5644_, new_D5645_,
    new_D5646_, new_D5647_, new_D5648_, new_D5649_, new_D5650_, new_D5651_,
    new_D5652_, new_D5653_, new_D5654_, new_D5655_, new_D5656_, new_D5657_,
    new_D5658_, new_D5659_, new_D5660_, new_D5661_, new_D5662_, new_D5663_,
    new_D5664_, new_D5665_, new_D5666_, new_D5667_, new_D5668_, new_D5669_,
    new_D5670_, new_D5671_, new_D5672_, new_D5673_, new_D5674_, new_D5675_,
    new_D5676_, new_D5677_, new_D5678_, new_D5679_, new_D5680_, new_D5681_,
    new_D5682_, new_D5683_, new_D5684_, new_D5685_, new_D5686_, new_D5687_,
    new_D5688_, new_D5689_, new_D5690_, new_D5691_, new_D5692_, new_D5693_,
    new_D5694_, new_D5695_, new_D5696_, new_D5697_, new_D5698_, new_D5699_,
    new_D5700_, new_D5701_, new_D5702_, new_D5703_, new_D5704_, new_D5705_,
    new_D5706_, new_D5707_, new_D5708_, new_D5709_, new_D5710_, new_D5711_,
    new_D5712_, new_D5713_, new_D5714_, new_D5715_, new_D5716_, new_D5717_,
    new_D5718_, new_D5719_, new_D5720_, new_D5721_, new_D5722_, new_D5723_,
    new_D5724_, new_D5725_, new_D5726_, new_D5727_, new_D5728_, new_D5729_,
    new_D5730_, new_D5731_, new_D5732_, new_D5733_, new_D5734_, new_D5735_,
    new_D5736_, new_D5737_, new_D5738_, new_D5739_, new_D5740_, new_D5741_,
    new_D5742_, new_D5743_, new_D5744_, new_D5745_, new_D5746_, new_D5747_,
    new_D5748_, new_D5749_, new_D5750_, new_D5751_, new_D5752_, new_D5753_,
    new_D5754_, new_D5755_, new_D5756_, new_D5757_, new_D5758_, new_D5759_,
    new_D5760_, new_D5761_, new_D5762_, new_D5763_, new_D5764_, new_D5765_,
    new_D5766_, new_D5767_, new_D5768_, new_D5769_, new_D5770_, new_D5771_,
    new_D5772_, new_D5773_, new_D5774_, new_D5775_, new_D5776_, new_D5777_,
    new_D5778_, new_D5779_, new_D5780_, new_D5781_, new_D5782_, new_D5783_,
    new_D5784_, new_D5785_, new_D5786_, new_D5787_, new_D5788_, new_D5789_,
    new_D5790_, new_D5791_, new_D5792_, new_D5793_, new_D5794_, new_D5795_,
    new_D5796_, new_D5797_, new_D5798_, new_D5799_, new_D5800_, new_D5801_,
    new_D5802_, new_D5803_, new_D5804_, new_D5805_, new_D5806_, new_D5807_,
    new_D5808_, new_D5809_, new_D5810_, new_D5811_, new_D5812_, new_D5813_,
    new_D5814_, new_D5815_, new_D5816_, new_D5817_, new_D5818_, new_D5819_,
    new_D5820_, new_D5821_, new_D5822_, new_D5823_, new_D5824_, new_D5825_,
    new_D5826_, new_D5827_, new_D5828_, new_D5829_, new_D5830_, new_D5831_,
    new_D5832_, new_D5833_, new_D5834_, new_D5835_, new_D5836_, new_D5837_,
    new_D5838_, new_D5839_, new_D5840_, new_D5841_, new_D5842_, new_D5843_,
    new_D5844_, new_D5845_, new_D5846_, new_D5847_, new_D5848_, new_D5849_,
    new_D5850_, new_D5851_, new_D5852_, new_D5853_, new_D5854_, new_D5855_,
    new_D5856_, new_D5857_, new_D5858_, new_D5859_, new_D5860_, new_D5861_,
    new_D5862_, new_D5863_, new_D5864_, new_D5865_, new_D5866_, new_D5867_,
    new_D5868_, new_D5869_, new_D5870_, new_D5871_, new_D5872_, new_D5873_,
    new_D5874_, new_D5875_, new_D5876_, new_D5877_, new_D5878_, new_D5879_,
    new_D5880_, new_D5881_, new_D5882_, new_D5883_, new_D5884_, new_D5885_,
    new_D5886_, new_D5887_, new_D5888_, new_D5889_, new_D5890_, new_D5891_,
    new_D5892_, new_D5893_, new_D5894_, new_D5895_, new_D5896_, new_D5897_,
    new_D5898_, new_D5899_, new_D5900_, new_D5901_, new_D5902_, new_D5903_,
    new_D5904_, new_D5905_, new_D5906_, new_D5907_, new_D5908_, new_D5909_,
    new_D5910_, new_D5911_, new_D5912_, new_D5913_, new_D5914_, new_D5915_,
    new_D5916_, new_D5917_, new_D5918_, new_D5919_, new_D5920_, new_D5921_,
    new_D5922_, new_D5923_, new_D5924_, new_D5925_, new_D5926_, new_D5927_,
    new_D5928_, new_D5929_, new_D5930_, new_D5931_, new_D5932_, new_D5933_,
    new_D5934_, new_D5935_, new_D5936_, new_D5937_, new_D5938_, new_D5939_,
    new_D5940_, new_D5941_, new_D5942_, new_D5943_, new_D5944_, new_D5945_,
    new_D5946_, new_D5947_, new_D5948_, new_D5949_, new_D5950_, new_D5951_,
    new_D5952_, new_D5953_, new_D5954_, new_D5955_, new_D5956_, new_D5957_,
    new_D5958_, new_D5959_, new_D5960_, new_D5961_, new_D5962_, new_D5963_,
    new_D5964_, new_D5965_, new_D5966_, new_D5967_, new_D5968_, new_D5969_,
    new_D5970_, new_D5971_, new_D5972_, new_D5973_, new_D5974_, new_D5975_,
    new_D5976_, new_D5977_, new_D5978_, new_D5979_, new_D5980_, new_D5981_,
    new_D5982_, new_D5983_, new_D5984_, new_D5985_, new_D5986_, new_D5987_,
    new_D5988_, new_D5989_, new_D5990_, new_D5991_, new_D5992_, new_D5993_,
    new_D5994_, new_D5995_, new_D5996_, new_D5997_, new_D5998_, new_D5999_,
    new_D6000_, new_D6001_, new_D6002_, new_D6003_, new_D6004_, new_D6005_,
    new_D6006_, new_D6007_, new_D6008_, new_D6009_, new_D6010_, new_D6011_,
    new_D6012_, new_D6013_, new_D6014_, new_D6015_, new_D6016_, new_D6017_,
    new_D6018_, new_D6019_, new_D6020_, new_D6021_, new_D6022_, new_D6023_,
    new_D6024_, new_D6025_, new_D6026_, new_D6027_, new_D6028_, new_D6029_,
    new_D6030_, new_D6031_, new_D6032_, new_D6033_, new_D6034_, new_D6035_,
    new_D6036_, new_D6037_, new_D6038_, new_D6039_, new_D6040_, new_D6041_,
    new_D6042_, new_D6043_, new_D6044_, new_D6045_, new_D6046_, new_D6047_,
    new_D6048_, new_D6049_, new_D6050_, new_D6051_, new_D6052_, new_D6053_,
    new_D6054_, new_D6055_, new_D6056_, new_D6057_, new_D6058_, new_D6059_,
    new_D6060_, new_D6061_, new_D6062_, new_D6063_, new_D6064_, new_D6065_,
    new_D6066_, new_D6067_, new_D6068_, new_D6069_, new_D6070_, new_D6071_,
    new_D6072_, new_D6073_, new_D6074_, new_D6075_, new_D6076_, new_D6077_,
    new_D6078_, new_D6079_, new_D6080_, new_D6081_, new_D6082_, new_D6083_,
    new_D6084_, new_D6085_, new_D6086_, new_D6087_, new_D6088_, new_D6089_,
    new_D6090_, new_D6091_, new_D6092_, new_D6093_, new_D6094_, new_D6095_,
    new_D6096_, new_D6097_, new_D6098_, new_D6099_, new_D6100_, new_D6101_,
    new_D6102_, new_D6103_, new_D6104_, new_D6105_, new_D6106_, new_D6107_,
    new_D6108_, new_D6109_, new_D6110_, new_D6111_, new_D6112_, new_D6113_,
    new_D6114_, new_D6115_, new_D6116_, new_D6117_, new_D6118_, new_D6119_,
    new_D6120_, new_D6121_, new_D6122_, new_D6123_, new_D6124_, new_D6125_,
    new_D6126_, new_D6127_, new_D6128_, new_D6129_, new_D6130_, new_D6131_,
    new_D6132_, new_D6133_, new_D6134_, new_D6135_, new_D6136_, new_D6137_,
    new_D6138_, new_D6139_, new_D6140_, new_D6141_, new_D6142_, new_D6143_,
    new_D6144_, new_D6145_, new_D6146_, new_D6147_, new_D6148_, new_D6149_,
    new_D6150_, new_D6151_, new_D6152_, new_D6153_, new_D6154_, new_D6155_,
    new_D6156_, new_D6157_, new_D6158_, new_D6159_, new_D6160_, new_D6161_,
    new_D6162_, new_D6163_, new_D6164_, new_D6165_, new_D6166_, new_D6167_,
    new_D6168_, new_D6169_, new_D6170_, new_D6171_, new_D6172_, new_D6173_,
    new_D6174_, new_D6175_, new_D6176_, new_D6177_, new_D6178_, new_D6179_,
    new_D6180_, new_D6181_, new_D6182_, new_D6183_, new_D6184_, new_D6185_,
    new_D6186_, new_D6187_, new_D6188_, new_D6189_, new_D6190_, new_D6191_,
    new_D6192_, new_D6193_, new_D6194_, new_D6195_, new_D6196_, new_D6197_,
    new_D6198_, new_D6199_, new_D6200_, new_D6201_, new_D6202_, new_D6203_,
    new_D6204_, new_D6205_, new_D6206_, new_D6207_, new_D6208_, new_D6209_,
    new_D6210_, new_D6211_, new_D6212_, new_D6213_, new_D6214_, new_D6215_,
    new_D6216_, new_D6217_, new_D6218_, new_D6219_, new_D6220_, new_D6221_,
    new_D6222_, new_D6223_, new_D6224_, new_D6225_, new_D6226_, new_D6227_,
    new_D6228_, new_D6229_, new_D6230_, new_D6231_, new_D6232_, new_D6233_,
    new_D6234_, new_D6235_, new_D6236_, new_D6237_, new_D6238_, new_D6239_,
    new_D6240_, new_D6241_, new_D6242_, new_D6243_, new_D6244_, new_D6245_,
    new_D6246_, new_D6247_, new_D6248_, new_D6249_, new_D6250_, new_D6251_,
    new_D6252_, new_D6253_, new_D6254_, new_D6255_, new_D6256_, new_D6257_,
    new_D6258_, new_D6259_, new_D6260_, new_D6261_, new_D6262_, new_D6263_,
    new_D6264_, new_D6265_, new_D6266_, new_D6267_, new_D6268_, new_D6269_,
    new_D6270_, new_D6271_, new_D6272_, new_D6273_, new_D6274_, new_D6275_,
    new_D6276_, new_D6277_, new_D6278_, new_D6279_, new_D6280_, new_D6281_,
    new_D6282_, new_D6283_, new_D6284_, new_D6285_, new_D6286_, new_D6287_,
    new_D6288_, new_D6289_, new_D6290_, new_D6291_, new_D6292_, new_D6293_,
    new_D6294_, new_D6295_, new_D6296_, new_D6297_, new_D6298_, new_D6299_,
    new_D6300_, new_D6301_, new_D6302_, new_D6303_, new_D6304_, new_D6305_,
    new_D6306_, new_D6307_, new_D6308_, new_D6309_, new_D6310_, new_D6311_,
    new_D6312_, new_D6313_, new_D6314_, new_D6315_, new_D6316_, new_D6317_,
    new_D6318_, new_D6319_, new_D6320_, new_D6321_, new_D6322_, new_D6323_,
    new_D6324_, new_D6325_, new_D6326_, new_D6327_, new_D6328_, new_D6329_,
    new_D6330_, new_D6331_, new_D6332_, new_D6333_, new_D6334_, new_D6335_,
    new_D6336_, new_D6337_, new_D6338_, new_D6339_, new_D6340_, new_D6341_,
    new_D6342_, new_D6343_, new_D6344_, new_D6345_, new_D6346_, new_D6347_,
    new_D6348_, new_D6349_, new_D6350_, new_D6351_, new_D6352_, new_D6353_,
    new_D6354_, new_D6355_, new_D6356_, new_D6357_, new_D6358_, new_D6359_,
    new_D6360_, new_D6361_, new_D6362_, new_D6363_, new_D6364_, new_D6365_,
    new_D6366_, new_D6367_, new_D6368_, new_D6369_, new_D6370_, new_D6371_,
    new_D6372_, new_D6373_, new_D6374_, new_D6375_, new_D6376_, new_D6377_,
    new_D6378_, new_D6379_, new_D6380_, new_D6381_, new_D6382_, new_D6383_,
    new_D6384_, new_D6385_, new_D6386_, new_D6387_, new_D6388_, new_D6389_,
    new_D6390_, new_D6391_, new_D6392_, new_D6393_, new_D6394_, new_D6395_,
    new_D6396_, new_D6397_, new_D6398_, new_D6399_, new_D6400_, new_D6401_,
    new_D6402_, new_D6403_, new_D6404_, new_D6405_, new_D6406_, new_D6407_,
    new_D6408_, new_D6409_, new_D6410_, new_D6411_, new_D6412_, new_D6413_,
    new_D6414_, new_D6415_, new_D6416_, new_D6417_, new_D6418_, new_D6419_,
    new_D6420_, new_D6421_, new_D6422_, new_D6423_, new_D6424_, new_D6425_,
    new_D6426_, new_D6427_, new_D6428_, new_D6429_, new_D6430_, new_D6431_,
    new_D6432_, new_D6433_, new_D6434_, new_D6435_, new_D6436_, new_D6437_,
    new_D6438_, new_D6439_, new_D6440_, new_D6441_, new_D6442_, new_D6443_,
    new_D6444_, new_D6445_, new_D6446_, new_D6447_, new_D6448_, new_D6449_,
    new_D6450_, new_D6451_, new_D6452_, new_D6453_, new_D6454_, new_D6455_,
    new_D6456_, new_D6457_, new_D6458_, new_D6459_, new_D6460_, new_D6461_,
    new_D6462_, new_D6463_, new_D6464_, new_D6465_, new_D6466_, new_D6467_,
    new_D6468_, new_D6469_, new_D6470_, new_D6471_, new_D6472_, new_D6473_,
    new_D6474_, new_D6475_, new_D6476_, new_D6477_, new_D6478_, new_D6479_,
    new_D6480_, new_D6481_, new_D6482_, new_D6483_, new_D6484_, new_D6485_,
    new_D6486_, new_D6487_, new_D6488_, new_D6489_, new_D6490_, new_D6491_,
    new_D6492_, new_D6493_, new_D6494_, new_D6495_, new_D6496_, new_D6497_,
    new_D6498_, new_D6499_, new_D6500_, new_D6501_, new_D6502_, new_D6503_,
    new_D6504_, new_D6505_, new_D6506_, new_D6507_, new_D6508_, new_D6509_,
    new_D6510_, new_D6511_, new_D6512_, new_D6513_, new_D6514_, new_D6515_,
    new_D6516_, new_D6517_, new_D6518_, new_D6519_, new_D6520_, new_D6521_,
    new_D6522_, new_D6523_, new_D6524_, new_D6525_, new_D6526_, new_D6527_,
    new_D6528_, new_D6529_, new_D6530_, new_D6531_, new_D6532_, new_D6533_,
    new_D6534_, new_D6535_, new_D6536_, new_D6537_, new_D6538_, new_D6539_,
    new_D6540_, new_D6541_, new_D6542_, new_D6543_, new_D6544_, new_D6545_,
    new_D6546_, new_D6547_, new_D6548_, new_D6549_, new_D6550_, new_D6551_,
    new_D6552_, new_D6553_, new_D6554_, new_D6555_, new_D6556_, new_D6557_,
    new_D6558_, new_D6559_, new_D6560_, new_D6561_, new_D6562_, new_D6563_,
    new_D6564_, new_D6565_, new_D6566_, new_D6567_, new_D6568_, new_D6569_,
    new_D6570_, new_D6571_, new_D6572_, new_D6573_, new_D6574_, new_D6575_,
    new_D6576_, new_D6577_, new_D6578_, new_D6579_, new_D6580_, new_D6581_,
    new_D6582_, new_D6583_, new_D6584_, new_D6585_, new_D6586_, new_D6587_,
    new_D6588_, new_D6589_, new_D6590_, new_D6591_, new_D6592_, new_D6593_,
    new_D6594_, new_D6595_, new_D6596_, new_D6597_, new_D6598_, new_D6599_,
    new_D6600_, new_D6601_, new_D6602_, new_D6603_, new_D6604_, new_D6605_,
    new_D6606_, new_D6607_, new_D6608_, new_D6609_, new_D6610_, new_D6611_,
    new_D6612_, new_D6613_, new_D6614_, new_D6615_, new_D6616_, new_D6617_,
    new_D6618_, new_D6619_, new_D6620_, new_D6621_, new_D6622_, new_D6623_,
    new_D6624_, new_D6625_, new_D6626_, new_D6627_, new_D6628_, new_D6629_,
    new_D6630_, new_D6631_, new_D6632_, new_D6633_, new_D6634_, new_D6635_,
    new_D6636_, new_D6637_, new_D6638_, new_D6639_, new_D6640_, new_D6641_,
    new_D6642_, new_D6643_, new_D6644_, new_D6645_, new_D6646_, new_D6647_,
    new_D6648_, new_D6649_, new_D6650_, new_D6651_, new_D6652_, new_D6653_,
    new_D6654_, new_D6655_, new_D6656_, new_D6657_, new_D6658_, new_D6659_,
    new_D6660_, new_D6661_, new_D6662_, new_D6663_, new_D6664_, new_D6665_,
    new_D6666_, new_D6667_, new_D6668_, new_D6669_, new_D6670_, new_D6671_,
    new_D6672_, new_D6673_, new_D6674_, new_D6675_, new_D6676_, new_D6677_,
    new_D6678_, new_D6679_, new_D6680_, new_D6681_, new_D6682_, new_D6683_,
    new_D6684_, new_D6685_, new_D6686_, new_D6687_, new_D6688_, new_D6689_,
    new_D6690_, new_D6691_, new_D6692_, new_D6693_, new_D6694_, new_D6695_,
    new_D6696_, new_D6697_, new_D6698_, new_D6699_, new_D6700_, new_D6701_,
    new_D6702_, new_D6703_, new_D6704_, new_D6705_, new_D6706_, new_D6707_,
    new_D6708_, new_D6709_, new_D6710_, new_D6711_, new_D6712_, new_D6713_,
    new_D6714_, new_D6715_, new_D6716_, new_D6717_, new_D6718_, new_D6719_,
    new_D6720_, new_D6721_, new_D6722_, new_D6723_, new_D6724_, new_D6725_,
    new_D6726_, new_D6727_, new_D6728_, new_D6729_, new_D6730_, new_D6731_,
    new_D6732_, new_D6733_, new_D6734_, new_D6735_, new_D6736_, new_D6737_,
    new_D6738_, new_D6739_, new_D6740_, new_D6741_, new_D6742_, new_D6743_,
    new_D6744_, new_D6745_, new_D6746_, new_D6747_, new_D6748_, new_D6749_,
    new_D6750_, new_D6751_, new_D6752_, new_D6753_, new_D6754_, new_D6755_,
    new_D6756_, new_D6757_, new_D6758_, new_D6759_, new_D6760_, new_D6761_,
    new_D6762_, new_D6763_, new_D6764_, new_D6765_, new_D6766_, new_D6767_,
    new_D6768_, new_D6769_, new_D6770_, new_D6771_, new_D6772_, new_D6773_,
    new_D6774_, new_D6775_, new_D6776_, new_D6777_, new_D6778_, new_D6779_,
    new_D6780_, new_D6781_, new_D6782_, new_D6783_, new_D6784_, new_D6785_,
    new_D6786_, new_D6787_, new_D6788_, new_D6789_, new_D6790_, new_D6791_,
    new_D6792_, new_D6793_, new_D6794_, new_D6795_, new_D6796_, new_D6797_,
    new_D6798_, new_D6799_, new_D6800_, new_D6801_, new_D6802_, new_D6803_,
    new_D6804_, new_D6805_, new_D6806_, new_D6807_, new_D6808_, new_D6809_,
    new_D6810_, new_D6811_, new_D6812_, new_D6813_, new_D6814_, new_D6815_,
    new_D6816_, new_D6817_, new_D6818_, new_D6819_, new_D6820_, new_D6821_,
    new_D6822_, new_D6823_, new_D6824_, new_D6825_, new_D6826_, new_D6827_,
    new_D6828_, new_D6829_, new_D6830_, new_D6831_, new_D6832_, new_D6833_,
    new_D6834_, new_D6835_, new_D6836_, new_D6837_, new_D6838_, new_D6839_,
    new_D6840_, new_D6841_, new_D6842_, new_D6843_, new_D6844_, new_D6845_,
    new_D6846_, new_D6847_, new_D6848_, new_D6849_, new_D6850_, new_D6851_,
    new_D6852_, new_D6853_, new_D6854_, new_D6855_, new_D6856_, new_D6857_,
    new_D6858_, new_D6859_, new_D6860_, new_D6861_, new_D6862_, new_D6863_,
    new_D6864_, new_D6865_, new_D6866_, new_D6867_, new_D6868_, new_D6869_,
    new_D6870_, new_D6871_, new_D6872_, new_D6873_, new_D6874_, new_D6875_,
    new_D6876_, new_D6877_, new_D6878_, new_D6879_, new_D6880_, new_D6881_,
    new_D6882_, new_D6883_, new_D6884_, new_D6885_, new_D6886_, new_D6887_,
    new_D6888_, new_D6889_, new_D6890_, new_D6891_, new_D6892_, new_D6893_,
    new_D6894_, new_D6895_, new_D6896_, new_D6897_, new_D6898_, new_D6899_,
    new_D6900_, new_D6901_, new_D6902_, new_D6903_, new_D6904_, new_D6905_,
    new_D6906_, new_D6907_, new_D6908_, new_D6909_, new_D6910_, new_D6911_,
    new_D6912_, new_D6913_, new_D6914_, new_D6915_, new_D6916_, new_D6917_,
    new_D6918_, new_D6919_, new_D6920_, new_D6921_, new_D6922_, new_D6923_,
    new_D6924_, new_D6925_, new_D6926_, new_D6927_, new_D6928_, new_D6929_,
    new_D6930_, new_D6931_, new_D6932_, new_D6933_, new_D6934_, new_D6935_,
    new_D6936_, new_D6937_, new_D6938_, new_D6939_, new_D6940_, new_D6941_,
    new_D6942_, new_D6943_, new_D6944_, new_D6945_, new_D6946_, new_D6947_,
    new_D6948_, new_D6949_, new_D6950_, new_D6951_, new_D6952_, new_D6953_,
    new_D6954_, new_D6955_, new_D6956_, new_D6957_, new_D6958_, new_D6959_,
    new_D6960_, new_D6961_, new_D6962_, new_D6963_, new_D6964_, new_D6965_,
    new_D6966_, new_D6967_, new_D6968_, new_D6969_, new_D6970_, new_D6971_,
    new_D6972_, new_D6973_, new_D6974_, new_D6975_, new_D6976_, new_D6977_,
    new_D6978_, new_D6979_, new_D6980_, new_D6981_, new_D6982_, new_D6983_,
    new_D6984_, new_D6985_, new_D6986_, new_D6987_, new_C2514_, new_C2513_,
    new_C2512_, new_C2511_, new_C2510_, new_C2509_, new_C2508_, new_C2507_,
    new_C2506_, new_C2505_, new_C2504_, new_C2503_, new_C2502_, new_C2501_,
    new_C2500_, new_C2499_, new_C2498_, new_C2497_, new_C2496_, new_C2495_,
    new_C2494_, new_C2493_, new_C2492_, new_C2491_, new_C2490_, new_C2489_,
    new_C2488_, new_C2487_, new_C2486_, new_C2485_, new_C2484_, new_C2483_,
    new_C2482_, new_C2481_, new_C2480_, new_C2479_, new_C2478_, new_C2477_,
    new_C2476_, new_C2475_, new_C2474_, new_C2473_, new_C2472_, new_C2471_,
    new_C2470_, new_C2469_, new_C2468_, new_C2467_, new_C2466_, new_C2465_,
    new_C2464_, new_C2463_, new_C2462_, new_C2461_, new_C2460_, new_C2453_,
    new_C2452_, new_C2451_, new_C2450_, new_C2449_, new_C2448_, new_C2447_,
    new_C2446_, new_C2445_, new_C2444_, new_C2443_, new_C2442_, new_C2441_,
    new_C2440_, new_C2439_, new_C2438_, new_C2437_, new_C2436_, new_C2435_,
    new_C2434_, new_C2433_, new_C2432_, new_C2431_, new_C2430_, new_C2429_,
    new_C2428_, new_C2427_, new_C2426_, new_C2425_, new_C2424_, new_C2423_,
    new_C2422_, new_C2421_, new_C2420_, new_C2419_, new_C2418_, new_C2417_,
    new_C2416_, new_C2415_, new_C2414_, new_C2413_, new_C2412_, new_C2411_,
    new_C2410_, new_C2409_, new_C2408_, new_C2407_, new_C2406_, new_C2405_,
    new_C2404_, new_C2403_, new_C2402_, new_C2401_, new_C2400_, new_C2399_,
    new_C2398_, new_C2397_, new_C2396_, new_C2395_, new_C2394_, new_C2393_,
    new_C2386_, new_C2385_, new_C2384_, new_C2383_, new_C2382_, new_C2381_,
    new_C2380_, new_C2379_, new_C2378_, new_C2377_, new_C2376_, new_C2375_,
    new_C2374_, new_C2373_, new_C2372_, new_C2371_, new_C2370_, new_C2369_,
    new_C2368_, new_C2367_, new_C2366_, new_C2365_, new_C2364_, new_C2363_,
    new_C2362_, new_C2361_, new_C2360_, new_C2359_, new_C2358_, new_C2357_,
    new_C2356_, new_C2355_, new_C2354_, new_C2353_, new_C2352_, new_C2351_,
    new_C2350_, new_C2349_, new_C2348_, new_C2347_, new_C2346_, new_C2345_,
    new_C2344_, new_C2343_, new_C2342_, new_C2341_, new_C2340_, new_C2339_,
    new_C2338_, new_C2337_, new_C2336_, new_C2335_, new_C2334_, new_C2333_,
    new_C2332_, new_C2331_, new_C2330_, new_C2329_, new_C2328_, new_C2327_,
    new_C2326_, new_C2319_, new_C2318_, new_C2317_, new_C2316_, new_C2315_,
    new_C2314_, new_C2313_, new_C2312_, new_C2311_, new_C2310_, new_C2309_,
    new_C2308_, new_C2307_, new_C2306_, new_C2305_, new_C2304_, new_C2303_,
    new_C2302_, new_C2301_, new_C2300_, new_C2299_, new_C2298_, new_C2297_,
    new_C2296_, new_C2295_, new_C2294_, new_C2293_, new_C2292_, new_C2291_,
    new_C2290_, new_C2289_, new_C2288_, new_C2287_, new_C2286_, new_C2285_,
    new_C2284_, new_C2283_, new_C2282_, new_C2281_, new_C2280_, new_C2279_,
    new_C2278_, new_C2277_, new_C2276_, new_C2275_, new_C2274_, new_C2273_,
    new_C2272_, new_C2271_, new_C2270_, new_C2269_, new_C2268_, new_C2267_,
    new_C2266_, new_C2265_, new_C2264_, new_C2263_, new_C2262_, new_C2261_,
    new_C2260_, new_C2259_, new_C2252_, new_C2251_, new_C2250_, new_C2249_,
    new_C2248_, new_C2247_, new_C2246_, new_C2245_, new_C2244_, new_C2243_,
    new_C2242_, new_C2241_, new_C2240_, new_C2239_, new_C2238_, new_C2237_,
    new_C2236_, new_C2235_, new_C2234_, new_C2233_, new_C2232_, new_C2231_,
    new_C2230_, new_C2229_, new_C2228_, new_C2227_, new_C2226_, new_C2225_,
    new_C2224_, new_C2223_, new_C2222_, new_C2221_, new_C2220_, new_C2219_,
    new_C2218_, new_C2217_, new_C2216_, new_C2215_, new_C2214_, new_C2213_,
    new_C2212_, new_C2211_, new_C2210_, new_C2209_, new_C2208_, new_C2207_,
    new_C2206_, new_C2205_, new_C2204_, new_C2203_, new_C2202_, new_C2201_,
    new_C2200_, new_C2199_, new_C2198_, new_C2197_, new_C2196_, new_C2195_,
    new_C2194_, new_C2193_, new_C2192_, new_C2185_, new_C2184_, new_C2183_,
    new_C2182_, new_C2181_, new_C2180_, new_C2179_, new_C2178_, new_C2177_,
    new_C2176_, new_C2175_, new_C2174_, new_C2173_, new_C2172_, new_C2171_,
    new_C2170_, new_C2169_, new_C2168_, new_C2167_, new_C2166_, new_C2165_,
    new_C2164_, new_C2163_, new_C2162_, new_C2161_, new_C2160_, new_C2159_,
    new_C2158_, new_C2157_, new_C2156_, new_C2155_, new_C2154_, new_C2153_,
    new_C2152_, new_C2151_, new_C2150_, new_C2149_, new_C2148_, new_C2147_,
    new_C2146_, new_C2145_, new_C2144_, new_C2143_, new_C2142_, new_C2141_,
    new_C2140_, new_C2139_, new_C2138_, new_C2137_, new_C2136_, new_C2135_,
    new_C2134_, new_C2133_, new_C2132_, new_C2131_, new_C2130_, new_C2129_,
    new_C2128_, new_C2127_, new_C2126_, new_C2125_, new_C2118_, new_C2117_,
    new_C2116_, new_C2115_, new_C2114_, new_C2113_, new_C2112_, new_C2111_,
    new_C2110_, new_C2109_, new_C2108_, new_C2107_, new_C2106_, new_C2105_,
    new_C2104_, new_C2103_, new_C2102_, new_C2101_, new_C2100_, new_C2099_,
    new_C2098_, new_C2097_, new_C2096_, new_C2095_, new_C2094_, new_C2093_,
    new_C2092_, new_C2091_, new_C2090_, new_C2089_, new_C2088_, new_C2087_,
    new_C2086_, new_C2085_, new_C2084_, new_C2083_, new_C2082_, new_C2081_,
    new_C2080_, new_C2079_, new_C2078_, new_C2077_, new_C2076_, new_C2075_,
    new_C2074_, new_C2073_, new_C2072_, new_C2071_, new_C2070_, new_C2069_,
    new_C2068_, new_C2067_, new_C2066_, new_C2065_, new_C2064_, new_C2063_,
    new_C2062_, new_C2061_, new_C2060_, new_C2059_, new_C2058_, new_C2051_,
    new_C2050_, new_C2049_, new_C2048_, new_C2047_, new_C2046_, new_C2045_,
    new_C2044_, new_C2043_, new_C2042_, new_C2041_, new_C2040_, new_C2039_,
    new_C2038_, new_C2037_, new_C2036_, new_C2035_, new_C2034_, new_C2033_,
    new_C2032_, new_C2031_, new_C2030_, new_C2029_, new_C2028_, new_C2027_,
    new_C2026_, new_C2025_, new_C2024_, new_C2023_, new_C2022_, new_C2021_,
    new_C2020_, new_C2019_, new_C2018_, new_C2017_, new_C2016_, new_C2015_,
    new_C2014_, new_C2013_, new_C2012_, new_C2011_, new_C2010_, new_C2009_,
    new_C2008_, new_C2007_, new_C2006_, new_C2005_, new_C2004_, new_C2003_,
    new_C2002_, new_C2001_, new_C2000_, new_C1999_, new_C1998_, new_C1997_,
    new_C1996_, new_C1995_, new_C1994_, new_C1993_, new_C1992_, new_C1991_,
    new_C1984_, new_C1983_, new_C1982_, new_C1981_, new_C1980_, new_C1979_,
    new_C1978_, new_C1977_, new_C1976_, new_C1975_, new_C1974_, new_C1973_,
    new_C1972_, new_C1971_, new_C1970_, new_C1969_, new_C1968_, new_C1967_,
    new_C1966_, new_C1965_, new_C1964_, new_C1963_, new_C1962_, new_C1961_,
    new_C1960_, new_C1959_, new_C1958_, new_C1957_, new_C1956_, new_C1955_,
    new_C1954_, new_C1953_, new_C1952_, new_C1951_, new_C1950_, new_C1949_,
    new_C1948_, new_C1947_, new_C1946_, new_C1945_, new_C1944_, new_C1943_,
    new_C1942_, new_C1941_, new_C1940_, new_C1939_, new_C1938_, new_C1937_,
    new_C1936_, new_C1935_, new_C1934_, new_C1933_, new_C1932_, new_C1931_,
    new_C1930_, new_C1929_, new_C1928_, new_C1927_, new_C1926_, new_C1925_,
    new_C1924_, new_C1917_, new_C1916_, new_C1915_, new_C1914_, new_C1913_,
    new_C1912_, new_C1911_, new_C1910_, new_C1909_, new_C1908_, new_C1907_,
    new_C1906_, new_C1905_, new_C1904_, new_C1903_, new_C1902_, new_C1901_,
    new_C1900_, new_C1899_, new_C1898_, new_C1897_, new_C1896_, new_C1895_,
    new_C1894_, new_C1893_, new_C1892_, new_C1891_, new_C1890_, new_C1889_,
    new_C1888_, new_C1887_, new_C1886_, new_C1885_, new_C1884_, new_C1883_,
    new_C1882_, new_C1881_, new_C1880_, new_C1879_, new_C1878_, new_C1877_,
    new_C1876_, new_C1875_, new_C1874_, new_C1873_, new_C1872_, new_C1871_,
    new_C1870_, new_C1869_, new_C1868_, new_C1867_, new_C1866_, new_C1865_,
    new_C1864_, new_C1863_, new_C1862_, new_C1861_, new_C1860_, new_C1859_,
    new_C1858_, new_C1857_, new_C1850_, new_C1849_, new_C1848_, new_C1847_,
    new_C1846_, new_C1845_, new_C1844_, new_C1843_, new_C1842_, new_C1841_,
    new_C1840_, new_C1839_, new_C1838_, new_C1837_, new_C1836_, new_C1835_,
    new_C1834_, new_C1833_, new_C1832_, new_C1831_, new_C1830_, new_C1829_,
    new_C1828_, new_C1827_, new_C1826_, new_C1825_, new_C1824_, new_C1823_,
    new_C1822_, new_C1821_, new_C1820_, new_C1819_, new_C1818_, new_C1817_,
    new_C1816_, new_C1815_, new_C1814_, new_C1813_, new_C1812_, new_C1811_,
    new_C1810_, new_C1809_, new_C1808_, new_C1807_, new_C1806_, new_C1805_,
    new_C1804_, new_C1803_, new_C1802_, new_C1801_, new_C1800_, new_C1799_,
    new_C1798_, new_C1797_, new_C1796_, new_C1795_, new_C1794_, new_C1793_,
    new_C1792_, new_C1791_, new_C1790_, new_C1783_, new_C1782_, new_C1781_,
    new_C1780_, new_C1779_, new_C1778_, new_C1777_, new_C1776_, new_C1775_,
    new_C1774_, new_C1773_, new_C1772_, new_C1771_, new_C1770_, new_C1769_,
    new_C1768_, new_C1767_, new_C1766_, new_C1765_, new_C1764_, new_C1763_,
    new_C1762_, new_C1761_, new_C1760_, new_C1759_, new_C1758_, new_C1757_,
    new_C1756_, new_C1755_, new_C1754_, new_C1753_, new_C1752_, new_C1751_,
    new_C1750_, new_C1749_, new_C1748_, new_C1747_, new_C1746_, new_C1745_,
    new_C1744_, new_C1743_, new_C1742_, new_C1741_, new_C1740_, new_C1739_,
    new_C1738_, new_C1737_, new_C1736_, new_C1735_, new_C1734_, new_C1733_,
    new_C1732_, new_C1731_, new_C1730_, new_C1729_, new_C1728_, new_C1727_,
    new_C1726_, new_C1725_, new_C1724_, new_C1723_, new_C1716_, new_C1715_,
    new_C1714_, new_C1713_, new_C1712_, new_C1711_, new_C1710_, new_C1709_,
    new_C1708_, new_C1707_, new_C1706_, new_C1705_, new_C1704_, new_C1703_,
    new_C1702_, new_C1701_, new_C1700_, new_C1699_, new_C1698_, new_C1697_,
    new_C1696_, new_C1695_, new_C1694_, new_C1693_, new_C1692_, new_C1691_,
    new_C1690_, new_C1689_, new_C1688_, new_C1687_, new_C1686_, new_C1685_,
    new_C1684_, new_C1683_, new_C1682_, new_C1681_, new_C1680_, new_C1679_,
    new_C1678_, new_C1677_, new_C1676_, new_C1675_, new_C1674_, new_C1673_,
    new_C1672_, new_C1671_, new_C1670_, new_C1669_, new_C1668_, new_C1667_,
    new_C1666_, new_C1665_, new_C1664_, new_C1663_, new_C1662_, new_C1661_,
    new_C1660_, new_C1659_, new_C1658_, new_C1657_, new_C1656_, new_C1649_,
    new_C1648_, new_C1647_, new_C1646_, new_C1645_, new_C1644_, new_C1643_,
    new_C1642_, new_C1641_, new_C1640_, new_C1639_, new_C1638_, new_C1637_,
    new_C1636_, new_C1635_, new_C1634_, new_C1633_, new_C1632_, new_C1631_,
    new_C1630_, new_C1629_, new_C1628_, new_C1627_, new_C1626_, new_C1625_,
    new_C1624_, new_C1623_, new_C1622_, new_C1621_, new_C1620_, new_C1619_,
    new_C1618_, new_C1617_, new_C1616_, new_C1615_, new_C1614_, new_C1613_,
    new_C1612_, new_C1611_, new_C1610_, new_C1609_, new_C1608_, new_C1607_,
    new_C1606_, new_C1605_, new_C1604_, new_C1603_, new_C1602_, new_C1601_,
    new_C1600_, new_C1599_, new_C1598_, new_C1597_, new_C1596_, new_C1595_,
    new_C1594_, new_C1593_, new_C1592_, new_C1591_, new_C1590_, new_C1589_,
    new_C1582_, new_C1581_, new_C1580_, new_C1579_, new_C1578_, new_C1577_,
    new_C1576_, new_C1575_, new_C1574_, new_C1573_, new_C1572_, new_C1571_,
    new_C1570_, new_C1569_, new_C1568_, new_C1567_, new_C1566_, new_C1565_,
    new_C1564_, new_C1563_, new_C1562_, new_C1561_, new_C1560_, new_C1559_,
    new_C1558_, new_C1557_, new_C1556_, new_C1555_, new_C1554_, new_C1553_,
    new_C1552_, new_C1551_, new_C1550_, new_C1549_, new_C1548_, new_C1547_,
    new_C1546_, new_C1545_, new_C1544_, new_C1543_, new_C1542_, new_C1541_,
    new_C1540_, new_C1539_, new_C1538_, new_C1537_, new_C1536_, new_C1535_,
    new_C1534_, new_C1533_, new_C1532_, new_C1531_, new_C1530_, new_C1529_,
    new_C1528_, new_C1527_, new_C1526_, new_C1525_, new_C1524_, new_C1523_,
    new_C1522_, new_C1515_, new_C1514_, new_C1513_, new_C1512_, new_C1511_,
    new_C1510_, new_C1509_, new_C1508_, new_C1507_, new_C1506_, new_C1505_,
    new_C1504_, new_C1503_, new_C1502_, new_C1501_, new_C1500_, new_C1499_,
    new_C1498_, new_C1497_, new_C1496_, new_C1495_, new_C1494_, new_C1493_,
    new_C1492_, new_C1491_, new_C1490_, new_C1489_, new_C1488_, new_C1487_,
    new_C1486_, new_C1485_, new_C1484_, new_C1483_, new_C1482_, new_C1481_,
    new_C1480_, new_C1479_, new_C1478_, new_C1477_, new_C1476_, new_C1475_,
    new_C1474_, new_C1473_, new_C1472_, new_C1471_, new_C1470_, new_C1469_,
    new_C1468_, new_C1467_, new_C1466_, new_C1465_, new_C1464_, new_C1463_,
    new_C1462_, new_C1461_, new_C1460_, new_C1459_, new_C1458_, new_C1457_,
    new_C1456_, new_C1455_, new_C1448_, new_C1447_, new_C1446_, new_C1445_,
    new_C1444_, new_C1443_, new_C1442_, new_C1441_, new_C1440_, new_C1439_,
    new_C1438_, new_C1437_, new_C1436_, new_C1435_, new_C1434_, new_C1433_,
    new_C1432_, new_C1431_, new_C1430_, new_C1429_, new_C1428_, new_C1427_,
    new_C1426_, new_C1425_, new_C1424_, new_C1423_, new_C1422_, new_C1421_,
    new_C1420_, new_C1419_, new_C1418_, new_C1417_, new_C1416_, new_C1415_,
    new_C1414_, new_C1413_, new_C1412_, new_C1411_, new_C1410_, new_C1409_,
    new_C1408_, new_C1407_, new_C1406_, new_C1405_, new_C1404_, new_C1403_,
    new_C1402_, new_C1401_, new_C1400_, new_C1399_, new_C1398_, new_C1397_,
    new_C1396_, new_C1395_, new_C1394_, new_C1393_, new_C1392_, new_C1391_,
    new_C1390_, new_C1389_, new_C1388_, new_C1381_, new_C1380_, new_C1379_,
    new_C1378_, new_C1377_, new_C1376_, new_C1375_, new_C1374_, new_C1373_,
    new_C1372_, new_C1371_, new_C1370_, new_C1369_, new_C1368_, new_C1367_,
    new_C1366_, new_C1365_, new_C1364_, new_C1363_, new_C1362_, new_C1361_,
    new_C1360_, new_C1359_, new_C1358_, new_C1357_, new_C1356_, new_C1355_,
    new_C1354_, new_C1353_, new_C1352_, new_C1351_, new_C1350_, new_C1349_,
    new_C1348_, new_C1347_, new_C1346_, new_C1345_, new_C1344_, new_C1343_,
    new_C1342_, new_C1341_, new_C1340_, new_C1339_, new_C1338_, new_C1337_,
    new_C1336_, new_C1335_, new_C1334_, new_C1333_, new_C1332_, new_C1331_,
    new_C1330_, new_C1329_, new_C1328_, new_C1327_, new_C1326_, new_C1325_,
    new_C1324_, new_C1323_, new_C1322_, new_C1321_, new_C1314_, new_C1313_,
    new_C1312_, new_C1311_, new_C1310_, new_C1309_, new_C1308_, new_C1307_,
    new_C1306_, new_C1305_, new_C1304_, new_C1303_, new_C1302_, new_C1301_,
    new_C1300_, new_C1299_, new_C1298_, new_C1297_, new_C1296_, new_C1295_,
    new_C1294_, new_C1293_, new_C1292_, new_C1291_, new_C1290_, new_C1289_,
    new_C1288_, new_C1287_, new_C1286_, new_C1285_, new_C1284_, new_C1283_,
    new_C1282_, new_C1281_, new_C1280_, new_C1279_, new_C1278_, new_C1277_,
    new_C1276_, new_C1275_, new_C1274_, new_C1273_, new_C1272_, new_C1271_,
    new_C1270_, new_C1269_, new_C1268_, new_C1267_, new_C1266_, new_C1265_,
    new_C1264_, new_C1263_, new_C1262_, new_C1261_, new_C1260_, new_C1259_,
    new_C1258_, new_C1257_, new_C1256_, new_C1255_, new_C1254_, new_C1247_,
    new_C1246_, new_C1245_, new_C1244_, new_C1243_, new_C1242_, new_C1241_,
    new_C1240_, new_C1239_, new_C1238_, new_C1237_, new_C1236_, new_C1235_,
    new_C1234_, new_C1233_, new_C1232_, new_C1231_, new_C1230_, new_C1229_,
    new_C1228_, new_C1227_, new_C1226_, new_C1225_, new_C1224_, new_C1223_,
    new_C1222_, new_C1221_, new_C1220_, new_C1219_, new_C1218_, new_C1217_,
    new_C1216_, new_C1215_, new_C1214_, new_C1213_, new_C1212_, new_C1211_,
    new_C1210_, new_C1209_, new_C1208_, new_C1207_, new_C1206_, new_C1205_,
    new_C1204_, new_C1203_, new_C1202_, new_C1201_, new_C1200_, new_C1199_,
    new_C1198_, new_C1197_, new_C1196_, new_C1195_, new_C1194_, new_C1193_,
    new_C1192_, new_C1191_, new_C1190_, new_C1189_, new_C1188_, new_C1187_,
    new_C1180_, new_C1179_, new_C1178_, new_C1177_, new_C1176_, new_C1175_,
    new_C1174_, new_C1173_, new_C1172_, new_C1171_, new_C1170_, new_C1169_,
    new_C1168_, new_C1167_, new_C1166_, new_C1165_, new_C1164_, new_C1163_,
    new_C1162_, new_C1161_, new_C1160_, new_C1159_, new_C1158_, new_C1157_,
    new_C1156_, new_C1155_, new_C1154_, new_C1153_, new_C1152_, new_C1151_,
    new_C1150_, new_C1149_, new_C1148_, new_C1147_, new_C1146_, new_C1145_,
    new_C1144_, new_C1143_, new_C1142_, new_C1141_, new_C1140_, new_C1139_,
    new_C1138_, new_C1137_, new_C1136_, new_C1135_, new_C1134_, new_C1133_,
    new_C1132_, new_C1131_, new_C1130_, new_C1129_, new_C1128_, new_C1127_,
    new_C1126_, new_C1125_, new_C1124_, new_C1123_, new_C1122_, new_C1121_,
    new_C1120_, new_C1113_, new_C1112_, new_C1111_, new_C1110_, new_C1109_,
    new_C1108_, new_C1107_, new_C1106_, new_C1105_, new_C1104_, new_C1103_,
    new_C1102_, new_C1101_, new_C1100_, new_C1099_, new_C1098_, new_C1097_,
    new_C1096_, new_C1095_, new_C1094_, new_C1093_, new_C1092_, new_C1091_,
    new_C1090_, new_C1089_, new_C1088_, new_C1087_, new_C1086_, new_C1085_,
    new_C1084_, new_C1083_, new_C1082_, new_C1081_, new_C1080_, new_C1079_,
    new_C1078_, new_C1077_, new_C1076_, new_C1075_, new_C1074_, new_C1073_,
    new_C1072_, new_C1071_, new_C1070_, new_C1069_, new_C1068_, new_C1067_,
    new_C1066_, new_C1065_, new_C1064_, new_C1063_, new_C1062_, new_C1061_,
    new_C1060_, new_C1059_, new_C1058_, new_C1057_, new_C1056_, new_C1055_,
    new_C1054_, new_C1053_, new_C1046_, new_C1045_, new_C1044_, new_C1043_,
    new_C1042_, new_C1041_, new_C1040_, new_C1039_, new_C1038_, new_C1037_,
    new_C1036_, new_C1035_, new_C1034_, new_C1033_, new_C1032_, new_C1031_,
    new_C1030_, new_C1029_, new_C1028_, new_C1027_, new_C1026_, new_C1025_,
    new_C1024_, new_C1023_, new_C1022_, new_C1021_, new_C1020_, new_C1019_,
    new_C1018_, new_C1017_, new_C1016_, new_C1015_, new_C1014_, new_C1013_,
    new_C1012_, new_C1011_, new_C1010_, new_C1009_, new_C1008_, new_C1007_,
    new_C1006_, new_C1005_, new_C1004_, new_C1003_, new_C1002_, new_C1001_,
    new_C1000_, new_C999_, new_C998_, new_C997_, new_C996_, new_C995_,
    new_C994_, new_C993_, new_C992_, new_C991_, new_C990_, new_C989_,
    new_C988_, new_C987_, new_C986_, new_C979_, new_C978_, new_C977_,
    new_C976_, new_C975_, new_C974_, new_C973_, new_C972_, new_C971_,
    new_C970_, new_C969_, new_C968_, new_C967_, new_C966_, new_C965_,
    new_C964_, new_C963_, new_C962_, new_C961_, new_C960_, new_C959_,
    new_C958_, new_C957_, new_C956_, new_C955_, new_C954_, new_C953_,
    new_C952_, new_C951_, new_C950_, new_C949_, new_C948_, new_C947_,
    new_C946_, new_C945_, new_C944_, new_C943_, new_C942_, new_C941_,
    new_C940_, new_C939_, new_C938_, new_C937_, new_C936_, new_C935_,
    new_C934_, new_C933_, new_C932_, new_C931_, new_C930_, new_C929_,
    new_C928_, new_C927_, new_C926_, new_C925_, new_C924_, new_C923_,
    new_C922_, new_C921_, new_C920_, new_C919_, new_C912_, new_C911_,
    new_C910_, new_C909_, new_C908_, new_C907_, new_C906_, new_C905_,
    new_C904_, new_C903_, new_C902_, new_C901_, new_C900_, new_C899_,
    new_C898_, new_C897_, new_C896_, new_C895_, new_C894_, new_C893_,
    new_C892_, new_C891_, new_C890_, new_C889_, new_C888_, new_C887_,
    new_C886_, new_C885_, new_C884_, new_C883_, new_C882_, new_C881_,
    new_C880_, new_C879_, new_C878_, new_C877_, new_C876_, new_C875_,
    new_C874_, new_C873_, new_C872_, new_C871_, new_C870_, new_C869_,
    new_C868_, new_C867_, new_C866_, new_C865_, new_C864_, new_C863_,
    new_C862_, new_C861_, new_C860_, new_C859_, new_C858_, new_C857_,
    new_C856_, new_C855_, new_C854_, new_C853_, new_C852_, new_C845_,
    new_C844_, new_C843_, new_C842_, new_C841_, new_C840_, new_C839_,
    new_C838_, new_C837_, new_C836_, new_C835_, new_C834_, new_C833_,
    new_C832_, new_C831_, new_C830_, new_C829_, new_C828_, new_C827_,
    new_C826_, new_C825_, new_C824_, new_C823_, new_C822_, new_C821_,
    new_C820_, new_C819_, new_C818_, new_C817_, new_C816_, new_C815_,
    new_C814_, new_C813_, new_C812_, new_C811_, new_C810_, new_C809_,
    new_C808_, new_C807_, new_C806_, new_C805_, new_C804_, new_C803_,
    new_C802_, new_C801_, new_C800_, new_C799_, new_C798_, new_C797_,
    new_C796_, new_C795_, new_C794_, new_C793_, new_C792_, new_C791_,
    new_C790_, new_C789_, new_C788_, new_C787_, new_C786_, new_C785_,
    new_C778_, new_C777_, new_C776_, new_C775_, new_C774_, new_C773_,
    new_C772_, new_C771_, new_C770_, new_C769_, new_C768_, new_C767_,
    new_C766_, new_C765_, new_C764_, new_C763_, new_C762_, new_C761_,
    new_C760_, new_C759_, new_C758_, new_C757_, new_C756_, new_C755_,
    new_C754_, new_C753_, new_C752_, new_C751_, new_C750_, new_C749_,
    new_C748_, new_C747_, new_C746_, new_C745_, new_C744_, new_C743_,
    new_C742_, new_C741_, new_C740_, new_C739_, new_C738_, new_C737_,
    new_C736_, new_C735_, new_C734_, new_C733_, new_C732_, new_C731_,
    new_C730_, new_C729_, new_C728_, new_C727_, new_C726_, new_C725_,
    new_C724_, new_C723_, new_C722_, new_C721_, new_C720_, new_C719_,
    new_C718_, new_C711_, new_C710_, new_C709_, new_C708_, new_C707_,
    new_C706_, new_C705_, new_C704_, new_C703_, new_C702_, new_C701_,
    new_C700_, new_C699_, new_C698_, new_C697_, new_C696_, new_C695_,
    new_C694_, new_C693_, new_C692_, new_C691_, new_C690_, new_C689_,
    new_C688_, new_C687_, new_C686_, new_C685_, new_C684_, new_C683_,
    new_C682_, new_C681_, new_C680_, new_C679_, new_C678_, new_C677_,
    new_C676_, new_C675_, new_C674_, new_C673_, new_C672_, new_C671_,
    new_C670_, new_C669_, new_C668_, new_C667_, new_C666_, new_C665_,
    new_C664_, new_C663_, new_C662_, new_C661_, new_C660_, new_C659_,
    new_C658_, new_C657_, new_C656_, new_C655_, new_C654_, new_C653_,
    new_C652_, new_C651_, new_C644_, new_C643_, new_C642_, new_C641_,
    new_C640_, new_C639_, new_C638_, new_C637_, new_C636_, new_C635_,
    new_C634_, new_C633_, new_C632_, new_C631_, new_C630_, new_C629_,
    new_C628_, new_C627_, new_C626_, new_C625_, new_C624_, new_C623_,
    new_C622_, new_C621_, new_C620_, new_C619_, new_C618_, new_C617_,
    new_C616_, new_C615_, new_C614_, new_C613_, new_C612_, new_C611_,
    new_C610_, new_C609_, new_C608_, new_C607_, new_C606_, new_C605_,
    new_C604_, new_C603_, new_C602_, new_C601_, new_C600_, new_C599_,
    new_C598_, new_C597_, new_C596_, new_C595_, new_C594_, new_C593_,
    new_C592_, new_C591_, new_C590_, new_C589_, new_C588_, new_C587_,
    new_C586_, new_C585_, new_C584_, new_C577_, new_C576_, new_C575_,
    new_C574_, new_C573_, new_C572_, new_C571_, new_C570_, new_C569_,
    new_C568_, new_C567_, new_C566_, new_C565_, new_C564_, new_C563_,
    new_C562_, new_C561_, new_C560_, new_C559_, new_C558_, new_C557_,
    new_C556_, new_C555_, new_C554_, new_C553_, new_C552_, new_C551_,
    new_C550_, new_C549_, new_C548_, new_C547_, new_C546_, new_C545_,
    new_C544_, new_C543_, new_C542_, new_C541_, new_C540_, new_C539_,
    new_C538_, new_C537_, new_C536_, new_C535_, new_C534_, new_C533_,
    new_C532_, new_C531_, new_C530_, new_C529_, new_C528_, new_C527_,
    new_C526_, new_C525_, new_C524_, new_C523_, new_C522_, new_C521_,
    new_C520_, new_C519_, new_C518_, new_C517_, new_C510_, new_C509_,
    new_C508_, new_C507_, new_C506_, new_C505_, new_C504_, new_C503_,
    new_C502_, new_C501_, new_C500_, new_C499_, new_C498_, new_C497_,
    new_C496_, new_C495_, new_C494_, new_C493_, new_C492_, new_C491_,
    new_C490_, new_C489_, new_C488_, new_C487_, new_C486_, new_C485_,
    new_C484_, new_C483_, new_C482_, new_C481_, new_C480_, new_C479_,
    new_C478_, new_C477_, new_C476_, new_C475_, new_C474_, new_C473_,
    new_C472_, new_C471_, new_C470_, new_C469_, new_C468_, new_C467_,
    new_C466_, new_C465_, new_C464_, new_C463_, new_C462_, new_C461_,
    new_C460_, new_C459_, new_C458_, new_C457_, new_C456_, new_C455_,
    new_C454_, new_C453_, new_C452_, new_C451_, new_C450_, new_C443_,
    new_C442_, new_C441_, new_C440_, new_C439_, new_C438_, new_C437_,
    new_C436_, new_C435_, new_C434_, new_C433_, new_C432_, new_C431_,
    new_C430_, new_C429_, new_C428_, new_C427_, new_C426_, new_C425_,
    new_C424_, new_C423_, new_C422_, new_C421_, new_C420_, new_C419_,
    new_C418_, new_C417_, new_C416_, new_C415_, new_C414_, new_C413_,
    new_C412_, new_C411_, new_C410_, new_C409_, new_C408_, new_C407_,
    new_C406_, new_C405_, new_C404_, new_C403_, new_C402_, new_C401_,
    new_C400_, new_C399_, new_C398_, new_C397_, new_C396_, new_C395_,
    new_C394_, new_C393_, new_C392_, new_C391_, new_C390_, new_C389_,
    new_C388_, new_C387_, new_C386_, new_C385_, new_C384_, new_C383_,
    new_C376_, new_C375_, new_C374_, new_C373_, new_C372_, new_C371_,
    new_C370_, new_C369_, new_C368_, new_C367_, new_C366_, new_C365_,
    new_C364_, new_C363_, new_C362_, new_C361_, new_C360_, new_C359_,
    new_C358_, new_C357_, new_C356_, new_C355_, new_C354_, new_C353_,
    new_C352_, new_C351_, new_C350_, new_C349_, new_C348_, new_C347_,
    new_C346_, new_C345_, new_C344_, new_C343_, new_C342_, new_C341_,
    new_C340_, new_C339_, new_C338_, new_C337_, new_C336_, new_C335_,
    new_C334_, new_C333_, new_C332_, new_C331_, new_C330_, new_C329_,
    new_C328_, new_C327_, new_C326_, new_C325_, new_C324_, new_C323_,
    new_C322_, new_C321_, new_C320_, new_C319_, new_C318_, new_C317_,
    new_C316_, new_C309_, new_C308_, new_C307_, new_C306_, new_C305_,
    new_C304_, new_C303_, new_C302_, new_C301_, new_C300_, new_C299_,
    new_C298_, new_C297_, new_C296_, new_C295_, new_C294_, new_C293_,
    new_C292_, new_C291_, new_C290_, new_C289_, new_C288_, new_C287_,
    new_C286_, new_C285_, new_C284_, new_C283_, new_C282_, new_C281_,
    new_C280_, new_C279_, new_C278_, new_C277_, new_C276_, new_C275_,
    new_C274_, new_C273_, new_C272_, new_C271_, new_C270_, new_C269_,
    new_C268_, new_C267_, new_C266_, new_C265_, new_C264_, new_C263_,
    new_C262_, new_C261_, new_C260_, new_C259_, new_C258_, new_C257_,
    new_C256_, new_C255_, new_C254_, new_C253_, new_C252_, new_C251_,
    new_C250_, new_C249_, new_C242_, new_C241_, new_C240_, new_C239_,
    new_C238_, new_C237_, new_C236_, new_C235_, new_C234_, new_C233_,
    new_C232_, new_C231_, new_C230_, new_C229_, new_C228_, new_C227_,
    new_C226_, new_C225_, new_C224_, new_C223_, new_C222_, new_C221_,
    new_C220_, new_C219_, new_C218_, new_C217_, new_C216_, new_C215_,
    new_C214_, new_C213_, new_C212_, new_C211_, new_C210_, new_C209_,
    new_C208_, new_C207_, new_C206_, new_C205_, new_C204_, new_C203_,
    new_C202_, new_C201_, new_C200_, new_C199_, new_C198_, new_C197_,
    new_C196_, new_C195_, new_C194_, new_C193_, new_C192_, new_C191_,
    new_C190_, new_C189_, new_C188_, new_C187_, new_C186_, new_C185_,
    new_C184_, new_C183_, new_C182_, new_C175_, new_C174_, new_C173_,
    new_C172_, new_C171_, new_C170_, new_C169_, new_C168_, new_C167_,
    new_C166_, new_C165_, new_C164_, new_C163_, new_C162_, new_C161_,
    new_C160_, new_C159_, new_C158_, new_C157_, new_C156_, new_C155_,
    new_C154_, new_C153_, new_C152_, new_C151_, new_C150_, new_C149_,
    new_C148_, new_C147_, new_C146_, new_C145_, new_C144_, new_C143_,
    new_C142_, new_C141_, new_C140_, new_C139_, new_C138_, new_C137_,
    new_C136_, new_C135_, new_C134_, new_C133_, new_C132_, new_C131_,
    new_C130_, new_C129_, new_C128_, new_C127_, new_C126_, new_C125_,
    new_C124_, new_C123_, new_C122_, new_C121_, new_C120_, new_C119_,
    new_C118_, new_C117_, new_C116_, new_C115_, new_C108_, new_C107_,
    new_C106_, new_C105_, new_C104_, new_C103_, new_C102_, new_C101_,
    new_C100_, new_C99_, new_C98_, new_C97_, new_C96_, new_C95_, new_C94_,
    new_C93_, new_C92_, new_C91_, new_C90_, new_C89_, new_C88_, new_C87_,
    new_C86_, new_C85_, new_C84_, new_C83_, new_C82_, new_C81_, new_C80_,
    new_C79_, new_C78_, new_C77_, new_C76_, new_C75_, new_C74_, new_C73_,
    new_C72_, new_C71_, new_C70_, new_C69_, new_C68_, new_C67_, new_C66_,
    new_C65_, new_C64_, new_C63_, new_C62_, new_C61_, new_C60_, new_C59_,
    new_C58_, new_C57_, new_C56_, new_C55_, new_C54_, new_C53_, new_C52_,
    new_C51_, new_C50_, new_C49_, new_C48_, new_C41_, new_C40_, new_C39_,
    new_C38_, new_C37_, new_C36_, new_C35_, new_C34_, new_C33_, new_C32_,
    new_C31_, new_C30_, new_C29_, new_C28_, new_C27_, new_C26_, new_C25_,
    new_C24_, new_C23_, new_C22_, new_C21_, new_C20_, new_C19_, new_C18_,
    new_C17_, new_C16_, new_C15_, new_C14_, new_C13_, new_C12_, new_C11_,
    new_C10_, new_C9_, new_C8_, new_C7_, new_C6_, new_C5_, new_C4_,
    new_C3_, new_C2_, new_C1_, new_B9999_, new_B9998_, new_B9997_,
    new_B9996_, new_B9995_, new_B9994_, new_B9993_, new_B9992_, new_B9991_,
    new_B9990_, new_B9989_, new_B9988_, new_B9987_, new_B9986_, new_B9985_,
    new_B9984_, new_B9983_, new_B9982_, new_B9981_, new_B9980_, new_B9973_,
    new_B9972_, new_B9971_, new_B9970_, new_B9969_, new_B9968_, new_B9967_,
    new_B9966_, new_B9965_, new_B9964_, new_B9963_, new_B9962_, new_B9961_,
    new_B9960_, new_B9959_, new_B9958_, new_B9957_, new_B9956_, new_B9955_,
    new_B9954_, new_B9953_, new_B9952_, new_B9951_, new_B9950_, new_B9949_,
    new_B9948_, new_B9947_, new_B9946_, new_B9945_, new_B9944_, new_B9943_,
    new_B9942_, new_B9941_, new_B9940_, new_B9939_, new_B9938_, new_B9937_,
    new_B9936_, new_B9935_, new_B9934_, new_B9933_, new_B9932_, new_B9931_,
    new_B9930_, new_B9929_, new_B9928_, new_B9927_, new_B9926_, new_B9925_,
    new_B9924_, new_B9923_, new_B9922_, new_B9921_, new_B9920_, new_B9919_,
    new_B9918_, new_B9917_, new_B9916_, new_B9915_, new_B9914_, new_B9913_,
    new_B9906_, new_B9905_, new_B9904_, new_B9903_, new_B9902_, new_B9901_,
    new_B9900_, new_B9899_, new_B9898_, new_B9897_, new_B9896_, new_B9895_,
    new_B9894_, new_B9893_, new_B9892_, new_B9891_, new_B9890_, new_B9889_,
    new_B9888_, new_B9887_, new_B9886_, new_B9885_, new_B9884_, new_B9883_,
    new_B9882_, new_B9881_, new_B9880_, new_B9879_, new_B9878_, new_B9877_,
    new_B9876_, new_B9875_, new_B9874_, new_B9873_, new_B9872_, new_B9871_,
    new_B9870_, new_B9869_, new_B9868_, new_B9867_, new_B9866_, new_B9865_,
    new_B9864_, new_B9863_, new_B9862_, new_B9861_, new_B9860_, new_B9859_,
    new_B9858_, new_B9857_, new_B9856_, new_B9855_, new_B9854_, new_B9853_,
    new_B9852_, new_B9851_, new_B9850_, new_B9849_, new_B9848_, new_B9847_,
    new_B9846_, new_B9839_, new_B9838_, new_B9837_, new_B9836_, new_B9835_,
    new_B9834_, new_B9833_, new_B9832_, new_B9831_, new_B9830_, new_B9829_,
    new_B9828_, new_B9827_, new_B9826_, new_B9825_, new_B9824_, new_B9823_,
    new_B9822_, new_B9821_, new_B9820_, new_B9819_, new_B9818_, new_B9817_,
    new_B9816_, new_B9815_, new_B9814_, new_B9813_, new_B9812_, new_B9811_,
    new_B9810_, new_B9809_, new_B9808_, new_B9807_, new_B9806_, new_B9805_,
    new_B9804_, new_B9803_, new_B9802_, new_B9801_, new_B9800_, new_B9799_,
    new_B9798_, new_B9797_, new_B9796_, new_B9795_, new_B9794_, new_B9793_,
    new_B9792_, new_B9791_, new_B9790_, new_B9789_, new_B9788_, new_B9787_,
    new_B9786_, new_B9785_, new_B9784_, new_B9783_, new_B9782_, new_B9781_,
    new_B9780_, new_B9779_, new_B9772_, new_B9771_, new_B9770_, new_B9769_,
    new_B9768_, new_B9767_, new_B9766_, new_B9765_, new_B9764_, new_B9763_,
    new_B9762_, new_B9761_, new_B9760_, new_B9759_, new_B9758_, new_B9757_,
    new_B9756_, new_B9755_, new_B9754_, new_B9753_, new_B9752_, new_B9751_,
    new_B9750_, new_B9749_, new_B9748_, new_B9747_, new_B9746_, new_B9745_,
    new_B9744_, new_B9743_, new_B9742_, new_B9741_, new_B9740_, new_B9739_,
    new_B9738_, new_B9737_, new_B9736_, new_B9735_, new_B9734_, new_B9733_,
    new_B9732_, new_B9731_, new_B9730_, new_B9729_, new_B9728_, new_B9727_,
    new_B9726_, new_B9725_, new_B9724_, new_B9723_, new_B9722_, new_B9721_,
    new_B9720_, new_B9719_, new_B9718_, new_B9717_, new_B9716_, new_B9715_,
    new_B9714_, new_B9713_, new_B9712_, new_B9705_, new_B9704_, new_B9703_,
    new_B9702_, new_B9701_, new_B9700_, new_B9699_, new_B9698_, new_B9697_,
    new_B9696_, new_B9695_, new_B9694_, new_B9693_, new_B9692_, new_B9691_,
    new_B9690_, new_B9689_, new_B9688_, new_B9687_, new_B9686_, new_B9685_,
    new_B9684_, new_B9683_, new_B9682_, new_B9681_, new_B9680_, new_B9679_,
    new_B9678_, new_B9677_, new_B9676_, new_B9675_, new_B9674_, new_B9673_,
    new_B9672_, new_B9671_, new_B9670_, new_B9669_, new_B9668_, new_B9667_,
    new_B9666_, new_B9665_, new_B9664_, new_B9663_, new_B9662_, new_B9661_,
    new_B9660_, new_B9659_, new_B9658_, new_B9657_, new_B9656_, new_B9655_,
    new_B9654_, new_B9653_, new_B9652_, new_B9651_, new_B9650_, new_B9649_,
    new_B9648_, new_B9647_, new_B9646_, new_B9645_, new_B9638_, new_B9637_,
    new_B9636_, new_B9635_, new_B9634_, new_B9633_, new_B9632_, new_B9631_,
    new_B9630_, new_B9629_, new_B9628_, new_B9627_, new_B9626_, new_B9625_,
    new_B9624_, new_B9623_, new_B9622_, new_B9621_, new_B9620_, new_B9619_,
    new_B9618_, new_B9617_, new_B9616_, new_B9615_, new_B9614_, new_B9613_,
    new_B9612_, new_B9611_, new_B9610_, new_B9609_, new_B9608_, new_B9607_,
    new_B9606_, new_B9605_, new_B9604_, new_B9603_, new_B9602_, new_B9601_,
    new_B9600_, new_B9599_, new_B9598_, new_B9597_, new_B9596_, new_B9595_,
    new_B9594_, new_B9593_, new_B9592_, new_B9591_, new_B9590_, new_B9589_,
    new_B9588_, new_B9587_, new_B9586_, new_B9585_, new_B9584_, new_B9583_,
    new_B9582_, new_B9581_, new_B9580_, new_B9579_, new_B9578_, new_B9571_,
    new_B9570_, new_B9569_, new_B9568_, new_B9567_, new_B9566_, new_B9565_,
    new_B9564_, new_B9563_, new_B9562_, new_B9561_, new_B9560_, new_B9559_,
    new_B9558_, new_B9557_, new_B9556_, new_B9555_, new_B9554_, new_B9553_,
    new_B9552_, new_B9551_, new_B9550_, new_B9549_, new_B9548_, new_B9547_,
    new_B9546_, new_B9545_, new_B9544_, new_B9543_, new_B9542_, new_B9541_,
    new_B9540_, new_B9539_, new_B9538_, new_B9537_, new_B9536_, new_B9535_,
    new_B9534_, new_B9533_, new_B9532_, new_B9531_, new_B9530_, new_B9529_,
    new_B9528_, new_B9527_, new_B9526_, new_B9525_, new_B9524_, new_B9523_,
    new_B9522_, new_B9521_, new_B9520_, new_B9519_, new_B9518_, new_B9517_,
    new_B9516_, new_B9515_, new_B9514_, new_B9513_, new_B9512_, new_B9511_,
    new_B9504_, new_B9503_, new_B9502_, new_B9501_, new_B9500_, new_B9499_,
    new_B9498_, new_B9497_, new_B9496_, new_B9495_, new_B9494_, new_B9493_,
    new_B9492_, new_B9491_, new_B9490_, new_B9489_, new_B9488_, new_B9487_,
    new_B9486_, new_B9485_, new_B9484_, new_B9483_, new_B9482_, new_B9481_,
    new_B9480_, new_B9479_, new_B9478_, new_B9477_, new_B9476_, new_B9475_,
    new_B9474_, new_B9473_, new_B9472_, new_B9471_, new_B9470_, new_B9469_,
    new_B9468_, new_B9467_, new_B9466_, new_B9465_, new_B9464_, new_B9463_,
    new_B9462_, new_B9461_, new_B9460_, new_B9459_, new_B9458_, new_B9457_,
    new_B9456_, new_B9455_, new_B9454_, new_B9453_, new_B9452_, new_B9451_,
    new_B9450_, new_B9449_, new_B9448_, new_B9447_, new_B9446_, new_B9445_,
    new_B9444_, new_B9437_, new_B9436_, new_B9435_, new_B9434_, new_B9433_,
    new_B9432_, new_B9431_, new_B9430_, new_B9429_, new_B9428_, new_B9427_,
    new_B9426_, new_B9425_, new_B9424_, new_B9423_, new_B9422_, new_B9421_,
    new_B9420_, new_B9419_, new_B9418_, new_B9417_, new_B9416_, new_B9415_,
    new_B9414_, new_B9413_, new_B9412_, new_B9411_, new_B9410_, new_B9409_,
    new_B9408_, new_B9407_, new_B9406_, new_B9405_, new_B9404_, new_B9403_,
    new_B9402_, new_B9401_, new_B9400_, new_B9399_, new_B9398_, new_B9397_,
    new_B9396_, new_B9395_, new_B9394_, new_B9393_, new_B9392_, new_B9391_,
    new_B9390_, new_B9389_, new_B9388_, new_B9387_, new_B9386_, new_B9385_,
    new_B9384_, new_B9383_, new_B9382_, new_B9381_, new_B9380_, new_B9379_,
    new_B9378_, new_B9377_, new_B9370_, new_B9369_, new_B9368_, new_B9367_,
    new_B9366_, new_B9365_, new_B9364_, new_B9363_, new_B9362_, new_B9361_,
    new_B9360_, new_B9359_, new_B9358_, new_B9357_, new_B9356_, new_B9355_,
    new_B9354_, new_B9353_, new_B9352_, new_B9351_, new_B9350_, new_B9349_,
    new_B9348_, new_B9347_, new_B9346_, new_B9345_, new_B9344_, new_B9343_,
    new_B9342_, new_B9341_, new_B9340_, new_B9339_, new_B9338_, new_B9337_,
    new_B9336_, new_B9335_, new_B9334_, new_B9333_, new_B9332_, new_B9331_,
    new_B9330_, new_B9329_, new_B9328_, new_B9327_, new_B9326_, new_B9325_,
    new_B9324_, new_B9323_, new_B9322_, new_B9321_, new_B9320_, new_B9319_,
    new_B9318_, new_B9317_, new_B9316_, new_B9315_, new_B9314_, new_B9313_,
    new_B9312_, new_B9311_, new_B9310_, new_B9303_, new_B9302_, new_B9301_,
    new_B9300_, new_B9299_, new_B9298_, new_B9297_, new_B9296_, new_B9295_,
    new_B9294_, new_B9293_, new_B9292_, new_B9291_, new_B9290_, new_B9289_,
    new_B9288_, new_B9287_, new_B9286_, new_B9285_, new_B9284_, new_B9283_,
    new_B9282_, new_B9281_, new_B9280_, new_B9279_, new_B9278_, new_B9277_,
    new_B9276_, new_B9275_, new_B9274_, new_B9273_, new_B9272_, new_B9271_,
    new_B9270_, new_B9269_, new_B9268_, new_B9267_, new_B9266_, new_B9265_,
    new_B9264_, new_B9263_, new_B9262_, new_B9261_, new_B9260_, new_B9259_,
    new_B9258_, new_B9257_, new_B9256_, new_B9255_, new_B9254_, new_B9253_,
    new_B9252_, new_B9251_, new_B9250_, new_B9249_, new_B9248_, new_B9247_,
    new_B9246_, new_B9245_, new_B9244_, new_B9243_, new_B9236_, new_B9235_,
    new_B9234_, new_B9233_, new_B9232_, new_B9231_, new_B9230_, new_B9229_,
    new_B9228_, new_B9227_, new_B9226_, new_B9225_, new_B9224_, new_B9223_,
    new_B9222_, new_B9221_, new_B9220_, new_B9219_, new_B9218_, new_B9217_,
    new_B9216_, new_B9215_, new_B9214_, new_B9213_, new_B9212_, new_B9211_,
    new_B9210_, new_B9209_, new_B9208_, new_B9207_, new_B9206_, new_B9205_,
    new_B9204_, new_B9203_, new_B9202_, new_B9201_, new_B9200_, new_B9199_,
    new_B9198_, new_B9197_, new_B9196_, new_B9195_, new_B9194_, new_B9193_,
    new_B9192_, new_B9191_, new_B9190_, new_B9189_, new_B9188_, new_B9187_,
    new_B9186_, new_B9185_, new_B9184_, new_B9183_, new_B9182_, new_B9181_,
    new_B9180_, new_B9179_, new_B9178_, new_B9177_, new_B9176_, new_B9169_,
    new_B9168_, new_B9167_, new_B9166_, new_B9165_, new_B9164_, new_B9163_,
    new_B9162_, new_B9161_, new_B9160_, new_B9159_, new_B9158_, new_B9157_,
    new_B9156_, new_B9155_, new_B9154_, new_B9153_, new_B9152_, new_B9151_,
    new_B9150_, new_B9149_, new_B9148_, new_B9147_, new_B9146_, new_B9145_,
    new_B9144_, new_B9143_, new_B9142_, new_B9141_, new_B9140_, new_B9139_,
    new_B9138_, new_B9137_, new_B9136_, new_B9135_, new_B9134_, new_B9133_,
    new_B9132_, new_B9131_, new_B9130_, new_B9129_, new_B9128_, new_B9127_,
    new_B9126_, new_B9125_, new_B9124_, new_B9123_, new_B9122_, new_B9121_,
    new_B9120_, new_B9119_, new_B9118_, new_B9117_, new_B9116_, new_B9115_,
    new_B9114_, new_B9113_, new_B9112_, new_B9111_, new_B9110_, new_B9109_,
    new_B9102_, new_B9101_, new_B9100_, new_B9099_, new_B9098_, new_B9097_,
    new_B9096_, new_B9095_, new_B9094_, new_B9093_, new_B9092_, new_B9091_,
    new_B9090_, new_B9089_, new_B9088_, new_B9087_, new_B9086_, new_B9085_,
    new_B9084_, new_B9083_, new_B9082_, new_B9081_, new_B9080_, new_B9079_,
    new_B9078_, new_B9077_, new_B9076_, new_B9075_, new_B9074_, new_B9073_,
    new_B9072_, new_B9071_, new_B9070_, new_B9069_, new_B9068_, new_B9067_,
    new_B9066_, new_B9065_, new_B9064_, new_B9063_, new_B9062_, new_B9061_,
    new_B9060_, new_B9059_, new_B9058_, new_B9057_, new_B9056_, new_B9055_,
    new_B9054_, new_B9053_, new_B9052_, new_B9051_, new_B9050_, new_B9049_,
    new_B9048_, new_B9047_, new_B9046_, new_B9045_, new_B9044_, new_B9043_,
    new_B9042_, new_B9035_, new_B9034_, new_B9033_, new_B9032_, new_B9031_,
    new_B9030_, new_B9029_, new_B9028_, new_B9027_, new_B9026_, new_B9025_,
    new_B9024_, new_B9023_, new_B9022_, new_B9021_, new_B9020_, new_B9019_,
    new_B9018_, new_B9017_, new_B9016_, new_B9015_, new_B9014_, new_B9013_,
    new_B9012_, new_B9011_, new_B9010_, new_B9009_, new_B9008_, new_B9007_,
    new_B9006_, new_B9005_, new_B9004_, new_B9003_, new_B9002_, new_B9001_,
    new_B9000_, new_B8999_, new_B8998_, new_B8997_, new_B8996_, new_B8995_,
    new_B8994_, new_B8993_, new_B8992_, new_B8991_, new_B8990_, new_B8989_,
    new_B8988_, new_B8987_, new_B8986_, new_B8985_, new_B8984_, new_B8983_,
    new_B8982_, new_B8981_, new_B8980_, new_B8979_, new_B8978_, new_B8977_,
    new_B8976_, new_B8975_, new_B8968_, new_B8967_, new_B8966_, new_B8965_,
    new_B8964_, new_B8963_, new_B8962_, new_B8961_, new_B8960_, new_B8959_,
    new_B8958_, new_B8957_, new_B8956_, new_B8955_, new_B8954_, new_B8953_,
    new_B8952_, new_B8951_, new_B8950_, new_B8949_, new_B8948_, new_B8947_,
    new_B8946_, new_B8945_, new_B8944_, new_B8943_, new_B8942_, new_B8941_,
    new_B8940_, new_B8939_, new_B8938_, new_B8937_, new_B8936_, new_B8935_,
    new_B8934_, new_B8933_, new_B8932_, new_B8931_, new_B8930_, new_B8929_,
    new_B8928_, new_B8927_, new_B8926_, new_B8925_, new_B8924_, new_B8923_,
    new_B8922_, new_B8921_, new_B8920_, new_B8919_, new_B8918_, new_B8917_,
    new_B8916_, new_B8915_, new_B8914_, new_B8913_, new_B8912_, new_B8911_,
    new_B8910_, new_B8909_, new_B8908_, new_B8901_, new_B8900_, new_B8899_,
    new_B8898_, new_B8897_, new_B8896_, new_B8895_, new_B8894_, new_B8893_,
    new_B8892_, new_B8891_, new_B8890_, new_B8889_, new_B8888_, new_B8887_,
    new_B8886_, new_B8885_, new_B8884_, new_B8883_, new_B8882_, new_B8881_,
    new_B8880_, new_B8879_, new_B8878_, new_B8877_, new_B8876_, new_B8875_,
    new_B8874_, new_B8873_, new_B8872_, new_B8871_, new_B8870_, new_B8869_,
    new_B8868_, new_B8867_, new_B8866_, new_B8865_, new_B8864_, new_B8863_,
    new_B8862_, new_B8861_, new_B8860_, new_B8859_, new_B8858_, new_B8857_,
    new_B8856_, new_B8855_, new_B8854_, new_B8853_, new_B8852_, new_B8851_,
    new_B8850_, new_B8849_, new_B8848_, new_B8847_, new_B8846_, new_B8845_,
    new_B8844_, new_B8843_, new_B8842_, new_B8841_, new_B8834_, new_B8833_,
    new_B8832_, new_B8831_, new_B8830_, new_B8829_, new_B8828_, new_B8827_,
    new_B8826_, new_B8825_, new_B8824_, new_B8823_, new_B8822_, new_B8821_,
    new_B8820_, new_B8819_, new_B8818_, new_B8817_, new_B8816_, new_B8815_,
    new_B8814_, new_B8813_, new_B8812_, new_B8811_, new_B8810_, new_B8809_,
    new_B8808_, new_B8807_, new_B8806_, new_B8805_, new_B8804_, new_B8803_,
    new_B8802_, new_B8801_, new_B8800_, new_B8799_, new_B8798_, new_B8797_,
    new_B8796_, new_B8795_, new_B8794_, new_B8793_, new_B8792_, new_B8791_,
    new_B8790_, new_B8789_, new_B8788_, new_B8787_, new_B8786_, new_B8785_,
    new_B8784_, new_B8783_, new_B8782_, new_B8781_, new_B8780_, new_B8779_,
    new_B8778_, new_B8777_, new_B8776_, new_B8775_, new_B8774_, new_B8767_,
    new_B8766_, new_B8765_, new_B8764_, new_B8763_, new_B8762_, new_B8761_,
    new_B8760_, new_B8759_, new_B8758_, new_B8757_, new_B8756_, new_B8755_,
    new_B8754_, new_B8753_, new_B8752_, new_B8751_, new_B8750_, new_B8749_,
    new_B8748_, new_B8747_, new_B8746_, new_B8745_, new_B8744_, new_B8743_,
    new_B8742_, new_B8741_, new_B8740_, new_B8739_, new_B8738_, new_B8737_,
    new_B8736_, new_B8735_, new_B8734_, new_B8733_, new_B8732_, new_B8731_,
    new_B8730_, new_B8729_, new_B8728_, new_B8727_, new_B8726_, new_B8725_,
    new_B8724_, new_B8723_, new_B8722_, new_B8721_, new_B8720_, new_B8719_,
    new_B8718_, new_B8717_, new_B8716_, new_B8715_, new_B8714_, new_B8713_,
    new_B8712_, new_B8711_, new_B8710_, new_B8709_, new_B8708_, new_B8707_,
    new_B8700_, new_B8699_, new_B8698_, new_B8697_, new_B8696_, new_B8695_,
    new_B8694_, new_B8693_, new_B8692_, new_B8691_, new_B8690_, new_B8689_,
    new_B8688_, new_B8687_, new_B8686_, new_B8685_, new_B8684_, new_B8683_,
    new_B8682_, new_B8681_, new_B8680_, new_B8679_, new_B8678_, new_B8677_,
    new_B8676_, new_B8675_, new_B8674_, new_B8673_, new_B8672_, new_B8671_,
    new_B8670_, new_B8669_, new_B8668_, new_B8667_, new_B8666_, new_B8665_,
    new_B8664_, new_B8663_, new_B8662_, new_B8661_, new_B8660_, new_B8659_,
    new_B8658_, new_B8657_, new_B8656_, new_B8655_, new_B8654_, new_B8653_,
    new_B8652_, new_B8651_, new_B8650_, new_B8649_, new_B8648_, new_B8647_,
    new_B8646_, new_B8645_, new_B8644_, new_B8643_, new_B8642_, new_B8641_,
    new_B8640_, new_B8633_, new_B8632_, new_B8631_, new_B8630_, new_B8629_,
    new_B8628_, new_B8627_, new_B8626_, new_B8625_, new_B8624_, new_B8623_,
    new_B8622_, new_B8621_, new_B8620_, new_B8619_, new_B8618_, new_B8617_,
    new_B8616_, new_B8615_, new_B8614_, new_B8613_, new_B8612_, new_B8611_,
    new_B8610_, new_B8609_, new_B8608_, new_B8607_, new_B8606_, new_B8605_,
    new_B8604_, new_B8603_, new_B8602_, new_B8601_, new_B8600_, new_B8599_,
    new_B8598_, new_B8597_, new_B8596_, new_B8595_, new_B8594_, new_B8593_,
    new_B8592_, new_B8591_, new_B8590_, new_B8589_, new_B8588_, new_B8587_,
    new_B8586_, new_B8585_, new_B8584_, new_B8583_, new_B8582_, new_B8581_,
    new_B8580_, new_B8579_, new_B8578_, new_B8577_, new_B8576_, new_B8575_,
    new_B8574_, new_B8573_, new_B8566_, new_B8565_, new_B8564_, new_B8563_,
    new_B8562_, new_B8561_, new_B8560_, new_B8559_, new_B8558_, new_B8557_,
    new_B8556_, new_B8555_, new_B8554_, new_B8553_, new_B8552_, new_B8551_,
    new_B8550_, new_B8549_, new_B8548_, new_B8547_, new_B8546_, new_B8545_,
    new_B8544_, new_B8543_, new_B8542_, new_B8541_, new_B8540_, new_B8539_,
    new_B8538_, new_B8537_, new_B8536_, new_B8535_, new_B8534_, new_B8533_,
    new_B8532_, new_B8531_, new_B8530_, new_B8529_, new_B8528_, new_B8527_,
    new_B8526_, new_B8525_, new_B8524_, new_B8523_, new_B8522_, new_B8521_,
    new_B8520_, new_B8519_, new_B8518_, new_B8517_, new_B8516_, new_B8515_,
    new_B8514_, new_B8513_, new_B8512_, new_B8511_, new_B8510_, new_B8509_,
    new_B8508_, new_B8507_, new_B8506_, new_B8499_, new_B8498_, new_B8497_,
    new_B8496_, new_B8495_, new_B8494_, new_B8493_, new_B8492_, new_B8491_,
    new_B8490_, new_B8489_, new_B8488_, new_B8487_, new_B8486_, new_B8485_,
    new_B8484_, new_B8483_, new_B8482_, new_B8481_, new_B8480_, new_B8479_,
    new_B8478_, new_B8477_, new_B8476_, new_B8475_, new_B8474_, new_B8473_,
    new_B8472_, new_B8471_, new_B8470_, new_B8469_, new_B8468_, new_B8467_,
    new_B8466_, new_B8465_, new_B8464_, new_B8463_, new_B8462_, new_B8461_,
    new_B8460_, new_B8459_, new_B8458_, new_B8457_, new_B8456_, new_B8455_,
    new_B8454_, new_B8453_, new_B8452_, new_B8451_, new_B8450_, new_B8449_,
    new_B8448_, new_B8447_, new_B8446_, new_B8445_, new_B8444_, new_B8443_,
    new_B8442_, new_B8441_, new_B8440_, new_B8439_, new_B8432_, new_B8431_,
    new_B8430_, new_B8429_, new_B8428_, new_B8427_, new_B8426_, new_B8425_,
    new_B8424_, new_B8423_, new_B8422_, new_B8421_, new_B8420_, new_B8419_,
    new_B8418_, new_B8417_, new_B8416_, new_B8415_, new_B8414_, new_B8413_,
    new_B8412_, new_B8411_, new_B8410_, new_B8409_, new_B8408_, new_B8407_,
    new_B8406_, new_B8405_, new_B8404_, new_B8403_, new_B8402_, new_B8401_,
    new_B8400_, new_B8399_, new_B8398_, new_B8397_, new_B8396_, new_B8395_,
    new_B8394_, new_B8393_, new_B8392_, new_B8391_, new_B8390_, new_B8389_,
    new_B8388_, new_B8387_, new_B8386_, new_B8385_, new_B8384_, new_B8383_,
    new_B8382_, new_B8381_, new_B8380_, new_B8379_, new_B8378_, new_B8377_,
    new_B8376_, new_B8375_, new_B8374_, new_B8373_, new_B8372_, new_B8365_,
    new_B8364_, new_B8363_, new_B8362_, new_B8361_, new_B8360_, new_B8359_,
    new_B8358_, new_B8357_, new_B8356_, new_B8355_, new_B8354_, new_B8353_,
    new_B8352_, new_B8351_, new_B8350_, new_B8349_, new_B8348_, new_B8347_,
    new_B8346_, new_B8345_, new_B8344_, new_B8343_, new_B8342_, new_B8341_,
    new_B8340_, new_B8339_, new_B8338_, new_B8337_, new_B8336_, new_B8335_,
    new_B8334_, new_B8333_, new_B8332_, new_B8331_, new_B8330_, new_B8329_,
    new_B8328_, new_B8327_, new_B8326_, new_B8325_, new_B8324_, new_B8323_,
    new_B8322_, new_B8321_, new_B8320_, new_B8319_, new_B8318_, new_B8317_,
    new_B8316_, new_B8315_, new_B8314_, new_B8313_, new_B8312_, new_B8311_,
    new_B8310_, new_B8309_, new_B8308_, new_B8307_, new_B8306_, new_B8305_,
    new_B8298_, new_B8297_, new_B8296_, new_B8295_, new_B8294_, new_B8293_,
    new_B8292_, new_B8291_, new_B8290_, new_B8289_, new_B8288_, new_B8287_,
    new_B8286_, new_B8285_, new_B8284_, new_B8283_, new_B8282_, new_B8281_,
    new_B8280_, new_B8279_, new_B8278_, new_B8277_, new_B8276_, new_B8275_,
    new_B8274_, new_B8273_, new_B8272_, new_B8271_, new_B8270_, new_B8269_,
    new_B8268_, new_B8267_, new_B8266_, new_B8265_, new_B8264_, new_B8263_,
    new_B8262_, new_B8261_, new_B8260_, new_B8259_, new_B8258_, new_B8257_,
    new_B8256_, new_B8255_, new_B8254_, new_B8253_, new_B8252_, new_B8251_,
    new_B8250_, new_B8249_, new_B8248_, new_B8247_, new_B8246_, new_B8245_,
    new_B8244_, new_B8243_, new_B8242_, new_B8241_, new_B8240_, new_B8239_,
    new_B8238_, new_B8231_, new_B8230_, new_B8229_, new_B8228_, new_B8227_,
    new_B8226_, new_B8225_, new_B8224_, new_B8223_, new_B8222_, new_B8221_,
    new_B8220_, new_B8219_, new_B8218_, new_B8217_, new_B8216_, new_B8215_,
    new_B8214_, new_B8213_, new_B8212_, new_B8211_, new_B8210_, new_B8209_,
    new_B8208_, new_B8207_, new_B8206_, new_B8205_, new_B8204_, new_B8203_,
    new_B8202_, new_B8201_, new_B8200_, new_B8199_, new_B8198_, new_B8197_,
    new_B8196_, new_B8195_, new_B8194_, new_B8193_, new_B8192_, new_B8191_,
    new_B8190_, new_B8189_, new_B8188_, new_B8187_, new_B8186_, new_B8185_,
    new_B8184_, new_B8183_, new_B8182_, new_B8181_, new_B8180_, new_B8179_,
    new_B8178_, new_B8177_, new_B8176_, new_B8175_, new_B8174_, new_B8173_,
    new_B8172_, new_B8171_, new_B8164_, new_B8163_, new_B8162_, new_B8161_,
    new_B8160_, new_B8159_, new_B8158_, new_B8157_, new_B8156_, new_B8155_,
    new_B8154_, new_B8153_, new_B8152_, new_B8151_, new_B8150_, new_B8149_,
    new_B8148_, new_B8147_, new_B8146_, new_B8145_, new_B8144_, new_B8143_,
    new_B8142_, new_B8141_, new_B8140_, new_B8139_, new_B8138_, new_B8137_,
    new_B8136_, new_B8135_, new_B8134_, new_B8133_, new_B8132_, new_B8131_,
    new_B8130_, new_B8129_, new_B8128_, new_B8127_, new_B8126_, new_B8125_,
    new_B8124_, new_B8123_, new_B8122_, new_B8121_, new_B8120_, new_B8119_,
    new_B8118_, new_B8117_, new_B8116_, new_B8115_, new_B8114_, new_B8113_,
    new_B8112_, new_B8111_, new_B8110_, new_B8109_, new_B8108_, new_B8107_,
    new_B8106_, new_B8105_, new_B8104_, new_B8097_, new_B8096_, new_B8095_,
    new_B8094_, new_B8093_, new_B8092_, new_B8091_, new_B8090_, new_B8089_,
    new_B8088_, new_B8087_, new_B8086_, new_B8085_, new_B8084_, new_B8083_,
    new_B8082_, new_B8081_, new_B8080_, new_B8079_, new_B8078_, new_B8077_,
    new_B8076_, new_B8075_, new_B8074_, new_B8073_, new_B8072_, new_B8071_,
    new_B8070_, new_B8069_, new_B8068_, new_B8067_, new_B8066_, new_B8065_,
    new_B8064_, new_B8063_, new_B8062_, new_B8061_, new_B8060_, new_B8059_,
    new_B8058_, new_B8057_, new_B8056_, new_B8055_, new_B8054_, new_B8053_,
    new_B8052_, new_B8051_, new_B8050_, new_B8049_, new_B8048_, new_B8047_,
    new_B8046_, new_B8045_, new_B8044_, new_B8043_, new_B8042_, new_B8041_,
    new_B8040_, new_B8039_, new_B8038_, new_B8037_, new_B8030_, new_B8029_,
    new_B8028_, new_B8027_, new_B8026_, new_B8025_, new_B8024_, new_B8023_,
    new_B8022_, new_B8021_, new_B8020_, new_B8019_, new_B8018_, new_B8017_,
    new_B8016_, new_B8015_, new_B8014_, new_B8013_, new_B8012_, new_B8011_,
    new_B8010_, new_B8009_, new_B8008_, new_B8007_, new_B8006_, new_B8005_,
    new_B8004_, new_B8003_, new_B8002_, new_B8001_, new_B8000_, new_B7999_,
    new_B7998_, new_B7997_, new_B7996_, new_B7995_, new_B7994_, new_B7993_,
    new_B7992_, new_B7991_, new_B7990_, new_B7989_, new_B7988_, new_B7987_,
    new_B7986_, new_B7985_, new_B7984_, new_B7983_, new_B7982_, new_B7981_,
    new_B7980_, new_B7979_, new_B7978_, new_B7977_, new_B7976_, new_B7975_,
    new_B7974_, new_B7973_, new_B7972_, new_B7971_, new_B7970_, new_B7963_,
    new_B7962_, new_B7961_, new_B7960_, new_B7959_, new_B7958_, new_B7957_,
    new_B7956_, new_B7955_, new_B7954_, new_B7953_, new_B7952_, new_B7951_,
    new_B7950_, new_B7949_, new_B7948_, new_B7947_, new_B7946_, new_B7945_,
    new_B7944_, new_B7943_, new_B7942_, new_B7941_, new_B7940_, new_B7939_,
    new_B7938_, new_B7937_, new_B7936_, new_B7935_, new_B7934_, new_B7933_,
    new_B7932_, new_B7931_, new_B7930_, new_B7929_, new_B7928_, new_B7927_,
    new_B7926_, new_B7925_, new_B7924_, new_B7923_, new_B7922_, new_B7921_,
    new_B7920_, new_B7919_, new_B7918_, new_B7917_, new_B7916_, new_B7915_,
    new_B7914_, new_B7913_, new_B7912_, new_B7911_, new_B7910_, new_B7909_,
    new_B7908_, new_B7907_, new_B7906_, new_B7905_, new_B7904_, new_B7903_,
    new_B7896_, new_B7895_, new_B7894_, new_B7893_, new_B7892_, new_B7891_,
    new_B7890_, new_B7889_, new_B7888_, new_B7887_, new_B7886_, new_B7885_,
    new_B7884_, new_B7883_, new_B7882_, new_B7881_, new_B7880_, new_B7879_,
    new_B7878_, new_B7877_, new_B7876_, new_B7875_, new_B7874_, new_B7873_,
    new_B7872_, new_B7871_, new_B7870_, new_B7869_, new_B7868_, new_B7867_,
    new_B7866_, new_B7865_, new_B7864_, new_B7863_, new_B7862_, new_B7861_,
    new_B7860_, new_B7859_, new_B7858_, new_B7857_, new_B7856_, new_B7855_,
    new_B7854_, new_B7853_, new_B7852_, new_B7851_, new_B7850_, new_B7849_,
    new_B7848_, new_B7847_, new_B7846_, new_B7845_, new_B7844_, new_B7843_,
    new_B7842_, new_B7841_, new_B7840_, new_B7839_, new_B7838_, new_B7837_,
    new_B7836_, new_B7829_, new_B7828_, new_B7827_, new_B7826_, new_B7825_,
    new_B7824_, new_B7823_, new_B7822_, new_B7821_, new_B7820_, new_B7819_,
    new_B7818_, new_B7817_, new_B7816_, new_B7815_, new_B7814_, new_B7813_,
    new_B7812_, new_B7811_, new_B7810_, new_B7809_, new_B7808_, new_B7807_,
    new_B7806_, new_B7805_, new_B7804_, new_B7803_, new_B7802_, new_B7801_,
    new_B7800_, new_B7799_, new_B7798_, new_B7797_, new_B7796_, new_B7795_,
    new_B7794_, new_B7793_, new_B7792_, new_B7791_, new_B7790_, new_B7789_,
    new_B7788_, new_B7787_, new_B7786_, new_B7785_, new_B7784_, new_B7783_,
    new_B7782_, new_B7781_, new_B7780_, new_B7779_, new_B7778_, new_B7777_,
    new_B7776_, new_B7775_, new_B7774_, new_B7773_, new_B7772_, new_B7771_,
    new_B7770_, new_B7769_, new_B7762_, new_B7761_, new_B7760_, new_B7759_,
    new_B7758_, new_B7757_, new_B7756_, new_B7755_, new_B7754_, new_B7753_,
    new_B7752_, new_B7751_, new_B7750_, new_B7749_, new_B7748_, new_B7747_,
    new_B7746_, new_B7745_, new_B7744_, new_B7743_, new_B7742_, new_B7741_,
    new_B7740_, new_B7739_, new_B7738_, new_B7737_, new_B7736_, new_B7735_,
    new_B7734_, new_B7733_, new_B7732_, new_B7731_, new_B7730_, new_B7729_,
    new_B7728_, new_B7727_, new_B7726_, new_B7725_, new_B7724_, new_B7723_,
    new_B7722_, new_B7721_, new_B7720_, new_B7719_, new_B7718_, new_B7717_,
    new_B7716_, new_B7715_, new_B7714_, new_B7713_, new_B7712_, new_B7711_,
    new_B7710_, new_B7709_, new_B7708_, new_B7707_, new_B7706_, new_B7705_,
    new_B7704_, new_B7703_, new_B7702_, new_B7695_, new_B7694_, new_B7693_,
    new_B7692_, new_B7691_, new_B7690_, new_B7689_, new_B7688_, new_B7687_,
    new_B7686_, new_B7685_, new_B7684_, new_B7683_, new_B7682_, new_B7681_,
    new_B7680_, new_B7679_, new_B7678_, new_B7677_, new_B7676_, new_B7675_,
    new_B7674_, new_B7673_, new_B7672_, new_B7671_, new_B7670_, new_B7669_,
    new_B7668_, new_B7667_, new_B7666_, new_B7665_, new_B7664_, new_B7663_,
    new_B7662_, new_B7661_, new_B7660_, new_B7659_, new_B7658_, new_B7657_,
    new_B7656_, new_B7655_, new_B7654_, new_B7653_, new_B7652_, new_B7651_,
    new_B7650_, new_B7649_, new_B7648_, new_B7647_, new_B7646_, new_B7645_,
    new_B7644_, new_B7643_, new_B7642_, new_B7641_, new_B7640_, new_B7639_,
    new_B7638_, new_B7637_, new_B7636_, new_B7635_, new_B7628_, new_B7627_,
    new_B7626_, new_B7625_, new_B7624_, new_B7623_, new_B7622_, new_B7621_,
    new_B7620_, new_B7619_, new_B7618_, new_B7617_, new_B7616_, new_B7615_,
    new_B7614_, new_B7613_, new_B7612_, new_B7611_, new_B7610_, new_B7609_,
    new_B7608_, new_B7607_, new_B7606_, new_B7605_, new_B7604_, new_B7603_,
    new_B7602_, new_B7601_, new_B7600_, new_B7599_, new_B7598_, new_B7597_,
    new_B7596_, new_B7595_, new_B7594_, new_B7593_, new_B7592_, new_B7591_,
    new_B7590_, new_B7589_, new_B7588_, new_B7587_, new_B7586_, new_B7585_,
    new_B7584_, new_B7583_, new_B7582_, new_B7581_, new_B7580_, new_B7579_,
    new_B7578_, new_B7577_, new_B7576_, new_B7575_, new_B7574_, new_B7573_,
    new_B7572_, new_B7571_, new_B7570_, new_B7569_, new_B7568_, new_B7561_,
    new_B7560_, new_B7559_, new_B7558_, new_B7557_, new_B7556_, new_B7555_,
    new_B7554_, new_B7553_, new_B7552_, new_B7551_, new_B7550_, new_B7549_,
    new_B7548_, new_B7547_, new_B7546_, new_B7545_, new_B7544_, new_B7543_,
    new_B7542_, new_B7541_, new_B7540_, new_B7539_, new_B7538_, new_B7537_,
    new_B7536_, new_B7535_, new_B7534_, new_B7533_, new_B7532_, new_B7531_,
    new_B7530_, new_B7529_, new_B7528_, new_B7527_, new_B7526_, new_B7525_,
    new_B7524_, new_B7523_, new_B7522_, new_B7521_, new_B7520_, new_B7519_,
    new_B7518_, new_B7517_, new_B7516_, new_B7515_, new_B7514_, new_B7513_,
    new_B7512_, new_B7511_, new_B7510_, new_B7509_, new_B7508_, new_B7507_,
    new_B7506_, new_B7505_, new_B7504_, new_B7503_, new_B7502_, new_B7501_,
    new_B7494_, new_B7493_, new_B7492_, new_B7491_, new_B7490_, new_B7489_,
    new_B7488_, new_B7487_, new_B7486_, new_B7485_, new_B7484_, new_B7483_,
    new_B7482_, new_B7481_, new_B7480_, new_B7479_, new_B7478_, new_B7477_,
    new_B7476_, new_B7475_, new_B7474_, new_B7473_, new_B7472_, new_B7471_,
    new_B7470_, new_B7469_, new_B7468_, new_B7467_, new_B7466_, new_B7465_,
    new_B7464_, new_B7463_, new_B7462_, new_B7461_, new_B7460_, new_B7459_,
    new_B7458_, new_B7457_, new_B7456_, new_B7455_, new_B7454_, new_B7453_,
    new_B7452_, new_B7451_, new_B7450_, new_B7449_, new_B7448_, new_B7447_,
    new_B7446_, new_B7445_, new_B7444_, new_B7443_, new_B7442_, new_B7441_,
    new_B7440_, new_B7439_, new_B7438_, new_B7437_, new_B7436_, new_B7435_,
    new_B7434_, new_B7427_, new_B7426_, new_B7425_, new_B7424_, new_B7423_,
    new_B7422_, new_B7421_, new_B7420_, new_B7419_, new_B7418_, new_B7417_,
    new_B7416_, new_B7415_, new_B7414_, new_B7413_, new_B7412_, new_B7411_,
    new_B7410_, new_B7409_, new_B7408_, new_B7407_, new_B7406_, new_B7405_,
    new_B7404_, new_B7403_, new_B7402_, new_B7401_, new_B7400_, new_B7399_,
    new_B7398_, new_B7397_, new_B7396_, new_B7395_, new_B7394_, new_B7393_,
    new_B7392_, new_B7391_, new_B7390_, new_B7389_, new_B7388_, new_B7387_,
    new_B7386_, new_B7385_, new_B7384_, new_B7383_, new_B7382_, new_B7381_,
    new_B7380_, new_B7379_, new_B7378_, new_B7377_, new_B7376_, new_B7375_,
    new_B7374_, new_B7373_, new_B7372_, new_B7371_, new_B7370_, new_B7369_,
    new_B7368_, new_B7367_, new_B7360_, new_B7359_, new_B7358_, new_B7357_,
    new_B7356_, new_B7355_, new_B7354_, new_B7353_, new_B7352_, new_B7351_,
    new_B7350_, new_B7349_, new_B7348_, new_B7347_, new_B7346_, new_B7345_,
    new_B7344_, new_B7343_, new_B7342_, new_B7341_, new_B7340_, new_B7339_,
    new_B7338_, new_B7337_, new_B7336_, new_B7335_, new_B7334_, new_B7333_,
    new_B7332_, new_B7331_, new_B7330_, new_B7329_, new_B7328_, new_B7327_,
    new_B7326_, new_B7325_, new_B7324_, new_B7323_, new_B7322_, new_B7321_,
    new_B7320_, new_B7319_, new_B7318_, new_B7317_, new_B7316_, new_B7315_,
    new_B7314_, new_B7313_, new_B7312_, new_B7311_, new_B7310_, new_B7309_,
    new_B7308_, new_B7307_, new_B7306_, new_B7305_, new_B7304_, new_B7303_,
    new_B7302_, new_B7301_, new_B7300_, new_B7293_, new_B7292_, new_B7291_,
    new_B7290_, new_B7289_, new_B7288_, new_B7287_, new_B7286_, new_B7285_,
    new_B7284_, new_B7283_, new_B7282_, new_B7281_, new_B7280_, new_B7279_,
    new_B7278_, new_B7277_, new_B7276_, new_B7275_, new_B7274_, new_B7273_,
    new_B7272_, new_B7271_, new_B7270_, new_B7269_, new_B7268_, new_B7267_,
    new_B7266_, new_B7265_, new_B7264_, new_B7263_, new_B7262_, new_B7261_,
    new_B7260_, new_B7259_, new_B7258_, new_B7257_, new_B7256_, new_B7255_,
    new_B7254_, new_B7253_, new_B7252_, new_B7251_, new_B7250_, new_B7249_,
    new_B7248_, new_B7247_, new_B7246_, new_B7245_, new_B7244_, new_B7243_,
    new_B7242_, new_B7241_, new_B7240_, new_B7239_, new_B7238_, new_B7237_,
    new_B7236_, new_B7235_, new_B7234_, new_B7233_, new_B7226_, new_B7225_,
    new_B7224_, new_B7223_, new_B7222_, new_B7221_, new_B7220_, new_B7219_,
    new_B7218_, new_B7217_, new_B7216_, new_B7215_, new_B7214_, new_B7213_,
    new_B7212_, new_B7211_, new_B7210_, new_B7209_, new_B7208_, new_B7207_,
    new_B7206_, new_B7205_, new_B7204_, new_B7203_, new_B7202_, new_B7201_,
    new_B7200_, new_B7199_, new_B7198_, new_B7197_, new_B7196_, new_B7195_,
    new_B7194_, new_B7193_, new_B7192_, new_B7191_, new_B7190_, new_B7189_,
    new_B7188_, new_B7187_, new_B7186_, new_B7185_, new_B7184_, new_B7183_,
    new_B7182_, new_B7181_, new_B7180_, new_B7179_, new_B7178_, new_B7177_,
    new_B7176_, new_B7175_, new_B7174_, new_B7173_, new_B7172_, new_B7171_,
    new_B7170_, new_B7169_, new_B7168_, new_B7167_, new_B7166_, new_B7159_,
    new_B7158_, new_B7157_, new_B7156_, new_B7155_, new_B7154_, new_B7153_,
    new_B7152_, new_B7151_, new_B7150_, new_B7149_, new_B7148_, new_B7147_,
    new_B7146_, new_B7145_, new_B7144_, new_B7143_, new_B7142_, new_B7141_,
    new_B7140_, new_B7139_, new_B7138_, new_B7137_, new_B7136_, new_B7135_,
    new_B7134_, new_B7133_, new_B7132_, new_B7131_, new_B7130_, new_B7129_,
    new_B7128_, new_B7127_, new_B7126_, new_B7125_, new_B7124_, new_B7123_,
    new_B7122_, new_B7121_, new_B7120_, new_B7119_, new_B7118_, new_B7117_,
    new_B7116_, new_B7115_, new_B7114_, new_B7113_, new_B7112_, new_B7111_,
    new_B7110_, new_B7109_, new_B7108_, new_B7107_, new_B7106_, new_B7105_,
    new_B7104_, new_B7103_, new_B7102_, new_B7101_, new_B7100_, new_B7099_,
    new_B7092_, new_B7091_, new_B7090_, new_B7089_, new_B7088_, new_B7087_,
    new_B7086_, new_B7085_, new_B7084_, new_B7083_, new_B7082_, new_B7081_,
    new_B7080_, new_B7079_, new_B7078_, new_B7077_, new_B7076_, new_B7075_,
    new_B7074_, new_B7073_, new_B7072_, new_B7071_, new_B7070_, new_B7069_,
    new_B7068_, new_B7067_, new_B7066_, new_B7065_, new_B7064_, new_B7063_,
    new_B7062_, new_B7061_, new_B7060_, new_B7059_, new_B7058_, new_B7057_,
    new_B7056_, new_B7055_, new_B7054_, new_B7053_, new_B7052_, new_B7051_,
    new_B7050_, new_B7049_, new_B7048_, new_B7047_, new_B7046_, new_B7045_,
    new_B7044_, new_B7043_, new_B7042_, new_B7041_, new_B7040_, new_B7039_,
    new_B7038_, new_B7037_, new_B7036_, new_B7035_, new_B7034_, new_B7033_,
    new_B7032_, new_B7025_, new_B7024_, new_B7023_, new_B7022_, new_B7021_,
    new_B7020_, new_B7019_, new_B7018_, new_B7017_, new_B7016_, new_B7015_,
    new_B7014_, new_B7013_, new_B7012_, new_B7011_, new_B7010_, new_B7009_,
    new_B7008_, new_B7007_, new_B7006_, new_B7005_, new_B7004_, new_B7003_,
    new_B7002_, new_B7001_, new_B7000_, new_B6999_, new_B6998_, new_B6997_,
    new_B6996_, new_B6995_, new_B6994_, new_B6993_, new_B6992_, new_B6991_,
    new_B6990_, new_B6989_, new_B6988_, new_B6987_, new_B6986_, new_B6985_,
    new_B6984_, new_B6983_, new_B6982_, new_B6981_, new_B6980_, new_B6979_,
    new_B6978_, new_B6977_, new_B6976_, new_B6975_, new_B6974_, new_B6973_,
    new_B6972_, new_B6971_, new_B6970_, new_B6969_, new_B6968_, new_B6967_,
    new_B6966_, new_B6965_, new_B6958_, new_B6957_, new_B6956_, new_B6955_,
    new_B6954_, new_B6953_, new_B6952_, new_B6951_, new_B6950_, new_B6949_,
    new_B6948_, new_B6947_, new_B6946_, new_B6945_, new_B6944_, new_B6943_,
    new_B6942_, new_B6941_, new_B6940_, new_B6939_, new_B6938_, new_B6937_,
    new_B6936_, new_B6935_, new_B6934_, new_B6933_, new_B6932_, new_B6931_,
    new_B6930_, new_B6929_, new_B6928_, new_B6927_, new_B6926_, new_B6925_,
    new_B6924_, new_B6923_, new_B6922_, new_B6921_, new_B6920_, new_B6919_,
    new_B6918_, new_B6917_, new_B6916_, new_B6915_, new_B6914_, new_B6913_,
    new_B6912_, new_B6911_, new_B6910_, new_B6909_, new_B6908_, new_B6907_,
    new_B6906_, new_B6905_, new_B6904_, new_B6903_, new_B6902_, new_B6901_,
    new_B6900_, new_B6899_, new_B6898_, new_B6891_, new_B6890_, new_B6889_,
    new_B6888_, new_B6887_, new_B6886_, new_B6885_, new_B6884_, new_B6883_,
    new_B6882_, new_B6881_, new_B6880_, new_B6879_, new_B6878_, new_B6877_,
    new_B6876_, new_B6875_, new_B6874_, new_B6873_, new_B6872_, new_B6871_,
    new_B6870_, new_B6869_, new_B6868_, new_B6867_, new_B6866_, new_B6865_,
    new_B6864_, new_B6863_, new_B6862_, new_B6861_, new_B6860_, new_B6859_,
    new_B6858_, new_B6857_, new_B6856_, new_B6855_, new_B6854_, new_B6853_,
    new_B6852_, new_B6851_, new_B6850_, new_B6849_, new_B6848_, new_B6847_,
    new_B6846_, new_B6845_, new_B6844_, new_B6843_, new_B6842_, new_B6841_,
    new_B6840_, new_B6839_, new_B6838_, new_B6837_, new_B6836_, new_B6835_,
    new_B6834_, new_B6833_, new_B6832_, new_B6831_, new_B6824_, new_B6823_,
    new_B6822_, new_B6821_, new_B6820_, new_B6819_, new_B6818_, new_B6817_,
    new_B6816_, new_B6815_, new_B6814_, new_B6813_, new_B6812_, new_B6811_,
    new_B6810_, new_B6809_, new_B6808_, new_B6807_, new_B6806_, new_B6805_,
    new_B6804_, new_B6803_, new_B6802_, new_B6801_, new_B6800_, new_B6799_,
    new_B6798_, new_B6797_, new_B6796_, new_B6795_, new_B6794_, new_B6793_,
    new_B6792_, new_B6791_, new_B6790_, new_B6789_, new_B6788_, new_B6787_,
    new_B6786_, new_B6785_, new_B6784_, new_B6783_, new_B6782_, new_B6781_,
    new_B6780_, new_B6779_, new_B6778_, new_B6777_, new_B6776_, new_B6775_,
    new_B6774_, new_B6773_, new_B6772_, new_B6771_, new_B6770_, new_B6769_,
    new_B6768_, new_B6767_, new_B6766_, new_B6765_, new_B6764_, new_B6757_,
    new_B6756_, new_B6755_, new_B6754_, new_B6753_, new_B6752_, new_B6751_,
    new_B6750_, new_B6749_, new_B6748_, new_B6747_, new_B6746_, new_B6745_,
    new_B6744_, new_B6743_, new_B6742_, new_B6741_, new_B6740_, new_B6739_,
    new_B6738_, new_B6737_, new_B6736_, new_B6735_, new_B6734_, new_B6733_,
    new_B6732_, new_B6731_, new_B6730_, new_B6729_, new_B6728_, new_B6727_,
    new_B6726_, new_B6725_, new_B6724_, new_B6723_, new_B6722_, new_B6721_,
    new_B6720_, new_B6719_, new_B6718_, new_B6717_, new_B6716_, new_B6715_,
    new_B6714_, new_B6713_, new_B6712_, new_B6711_, new_B6710_, new_B6709_,
    new_B6708_, new_B6707_, new_B6706_, new_B6705_, new_B6704_, new_B6703_,
    new_B6702_, new_B6701_, new_B6700_, new_B6699_, new_B6698_, new_B6697_,
    new_B6690_, new_B6689_, new_B6688_, new_B6687_, new_B6686_, new_B6685_,
    new_B6684_, new_B6683_, new_B6682_, new_B6681_, new_B6680_, new_B6679_,
    new_B6678_, new_B6677_, new_B6676_, new_B6675_, new_B6674_, new_B6673_,
    new_B6672_, new_B6671_, new_B6670_, new_B6669_, new_B6668_, new_B6667_,
    new_B6666_, new_B6665_, new_B6664_, new_B6663_, new_B6662_, new_B6661_,
    new_B6660_, new_B6659_, new_B6658_, new_B6657_, new_B6656_, new_B6655_,
    new_B6654_, new_B6653_, new_B6652_, new_B6651_, new_B6650_, new_B6649_,
    new_B6648_, new_B6647_, new_B6646_, new_B6645_, new_B6644_, new_B6643_,
    new_B6642_, new_B6641_, new_B6640_, new_B6639_, new_B6638_, new_B6637_,
    new_B6636_, new_B6635_, new_B6634_, new_B6633_, new_B6632_, new_B6631_,
    new_B6630_, new_B6623_, new_B6622_, new_B6621_, new_B6620_, new_B6619_,
    new_B6618_, new_B6617_, new_B6616_, new_B6615_, new_B6614_, new_B6613_,
    new_B6612_, new_B6611_, new_B6610_, new_B6609_, new_B6608_, new_B6607_,
    new_B6606_, new_B6605_, new_B6604_, new_B6603_, new_B6602_, new_B6601_,
    new_B6600_, new_B6599_, new_B6598_, new_B6597_, new_B6596_, new_B6595_,
    new_B6594_, new_B6593_, new_B6592_, new_B6591_, new_B6590_, new_B6589_,
    new_B6588_, new_B6587_, new_B6586_, new_B6585_, new_B6584_, new_B6583_,
    new_B6582_, new_B6581_, new_B6580_, new_B6579_, new_B6578_, new_B6577_,
    new_B6576_, new_B6575_, new_B6574_, new_B6573_, new_B6572_, new_B6571_,
    new_B6570_, new_B6569_, new_B6568_, new_B6567_, new_B6566_, new_B6565_,
    new_B6564_, new_B6563_, new_B6556_, new_B6555_, new_B6554_, new_B6553_,
    new_B6552_, new_B6551_, new_B6550_, new_B6549_, new_B6548_, new_B6547_,
    new_B6546_, new_B6545_, new_B6544_, new_B6543_, new_B6542_, new_B6541_,
    new_B6540_, new_B6539_, new_B6538_, new_B6537_, new_B6536_, new_B6535_,
    new_B6534_, new_B6533_, new_B6532_, new_B6531_, new_B6530_, new_B6529_,
    new_B6528_, new_B6527_, new_B6526_, new_B6525_, new_B6524_, new_B6523_,
    new_B6522_, new_B6521_, new_B6520_, new_B6519_, new_B6518_, new_B6517_,
    new_B6516_, new_B6515_, new_B6514_, new_B6513_, new_B6512_, new_B6511_,
    new_B6510_, new_B6509_, new_B6508_, new_B6507_, new_B6506_, new_B6505_,
    new_B6504_, new_B6503_, new_B6502_, new_B6501_, new_B6500_, new_B6499_,
    new_B6498_, new_B6497_, new_B6496_, new_B6489_, new_B6488_, new_B6487_,
    new_B6486_, new_B6485_, new_B6484_, new_B6483_, new_B6482_, new_B6481_,
    new_B6480_, new_B6479_, new_B6478_, new_B6477_, new_B6476_, new_B6475_,
    new_B6474_, new_B6473_, new_B6472_, new_B6471_, new_B6470_, new_B6469_,
    new_B6468_, new_B6467_, new_B6466_, new_B6465_, new_B6464_, new_B6463_,
    new_B6462_, new_B6461_, new_B6460_, new_B6459_, new_B6458_, new_B6457_,
    new_B6456_, new_B6455_, new_B6454_, new_B6453_, new_B6452_, new_B6451_,
    new_B6450_, new_B6449_, new_B6448_, new_B6447_, new_B6446_, new_B6445_,
    new_B6444_, new_B6443_, new_B6442_, new_B6441_, new_B6440_, new_B6439_,
    new_B6438_, new_B6437_, new_B6436_, new_B6435_, new_B6434_, new_B6433_,
    new_B6432_, new_B6431_, new_B6430_, new_B6429_, new_B6422_, new_B6421_,
    new_B6420_, new_B6419_, new_B6418_, new_B6417_, new_B6416_, new_B6415_,
    new_B6414_, new_B6413_, new_B6412_, new_B6411_, new_B6410_, new_B6409_,
    new_B6408_, new_B6407_, new_B6406_, new_B6405_, new_B6404_, new_B6403_,
    new_B6402_, new_B6401_, new_B6400_, new_B6399_, new_B6398_, new_B6397_,
    new_B6396_, new_B6395_, new_B6394_, new_B6393_, new_B6392_, new_B6391_,
    new_B6390_, new_B6389_, new_B6388_, new_B6387_, new_B6386_, new_B6385_,
    new_B6384_, new_B6383_, new_B6382_, new_B6381_, new_B6380_, new_B6379_,
    new_B6378_, new_B6377_, new_B6376_, new_B6375_, new_B6374_, new_B6373_,
    new_B6372_, new_B6371_, new_B6370_, new_B6369_, new_B6368_, new_B6367_,
    new_B6366_, new_B6365_, new_B6364_, new_B6363_, new_B6362_, new_B6355_,
    new_B6354_, new_B6353_, new_B6352_, new_B6351_, new_B6350_, new_B6349_,
    new_B6348_, new_B6347_, new_B6346_, new_B6345_, new_B6344_, new_B6343_,
    new_B6342_, new_B6341_, new_B6340_, new_B6339_, new_B6338_, new_B6337_,
    new_B6336_, new_B6335_, new_B6334_, new_B6333_, new_B6332_, new_B6331_,
    new_B6330_, new_B6329_, new_B6328_, new_B6327_, new_B6326_, new_B6325_,
    new_B6324_, new_B6323_, new_B6322_, new_B6321_, new_B6320_, new_B6319_,
    new_B6318_, new_B6317_, new_B6316_, new_B6315_, new_B6314_, new_B6313_,
    new_B6312_, new_B6311_, new_B6310_, new_B6309_, new_B6308_, new_B6307_,
    new_B6306_, new_B6305_, new_B6304_, new_B6303_, new_B6302_, new_B6301_,
    new_B6300_, new_B6299_, new_B6298_, new_B6297_, new_B6296_, new_B6295_,
    new_B6288_, new_B6287_, new_B6286_, new_B6285_, new_B6284_, new_B6283_,
    new_B6282_, new_B6281_, new_B6280_, new_B6279_, new_B6278_, new_B6277_,
    new_B6276_, new_B6275_, new_B6274_, new_B6273_, new_B6272_, new_B6271_,
    new_B6270_, new_B6269_, new_B6268_, new_B6267_, new_B6266_, new_B6265_,
    new_B6264_, new_B6263_, new_B6262_, new_B6261_, new_B6260_, new_B6259_,
    new_B6258_, new_B6257_, new_B6256_, new_B6255_, new_B6254_, new_B6253_,
    new_B6252_, new_B6251_, new_B6250_, new_B6249_, new_B6248_, new_B6247_,
    new_B6246_, new_B6245_, new_B6244_, new_B6243_, new_B6242_, new_B6241_,
    new_B6240_, new_B6239_, new_B6238_, new_B6237_, new_B6236_, new_B6235_,
    new_B6234_, new_B6233_, new_B6232_, new_B6231_, new_B6230_, new_B6229_,
    new_B6228_, new_B6221_, new_B6220_, new_B6219_, new_B6218_, new_B6217_,
    new_B6216_, new_B6215_, new_B6214_, new_B6213_, new_B6212_, new_B6211_,
    new_B6210_, new_B6209_, new_B6208_, new_B6207_, new_B6206_, new_B6205_,
    new_B6204_, new_B6203_, new_B6202_, new_B6201_, new_B6200_, new_B6199_,
    new_B6198_, new_B6197_, new_B6196_, new_B6195_, new_B6194_, new_B6193_,
    new_B6192_, new_B6191_, new_B6190_, new_B6189_, new_B6188_, new_B6187_,
    new_B6186_, new_B6185_, new_B6184_, new_B6183_, new_B6182_, new_B6181_,
    new_B6180_, new_B6179_, new_B6178_, new_B6177_, new_B6176_, new_B6175_,
    new_B6174_, new_B6173_, new_B6172_, new_B6171_, new_B6170_, new_B6169_,
    new_B6168_, new_B6167_, new_B6166_, new_B6165_, new_B6164_, new_B6163_,
    new_B6162_, new_B6161_, new_B6154_, new_B6153_, new_B6152_, new_B6151_,
    new_B6150_, new_B6149_, new_B6148_, new_B6147_, new_B6146_, new_B6145_,
    new_B6144_, new_B6143_, new_B6142_, new_B6141_, new_B6140_, new_B6139_,
    new_B6138_, new_B6137_, new_B6136_, new_B6135_, new_B6134_, new_B6133_,
    new_B6132_, new_B6131_, new_B6130_, new_B6129_, new_B6128_, new_B6127_,
    new_B6126_, new_B6125_, new_B6124_, new_B6123_, new_B6122_, new_B6121_,
    new_B6120_, new_B6119_, new_B6118_, new_B6117_, new_B6116_, new_B6115_,
    new_B6114_, new_B6113_, new_B6112_, new_B6111_, new_B6110_, new_B6109_,
    new_B6108_, new_B6107_, new_B6106_, new_B6105_, new_B6104_, new_B6103_,
    new_B6102_, new_B6101_, new_B6100_, new_B6099_, new_B6098_, new_B6097_,
    new_B6096_, new_B6095_, new_B6094_, new_B6087_, new_B6086_, new_B6085_,
    new_B6084_, new_B6083_, new_B6082_, new_B6081_, new_B6080_, new_B6079_,
    new_B6078_, new_B6077_, new_B6076_, new_B6075_, new_B6074_, new_B6073_,
    new_B6072_, new_B6071_, new_B6070_, new_B6069_, new_B6068_, new_B6067_,
    new_B6066_, new_B6065_, new_B6064_, new_B6063_, new_B6062_, new_B6061_,
    new_B6060_, new_B6059_, new_B6058_, new_B6057_, new_B6056_, new_B6055_,
    new_B6054_, new_B6053_, new_B6052_, new_B6051_, new_B6050_, new_B6049_,
    new_B6048_, new_B6047_, new_B6046_, new_B6045_, new_B6044_, new_B6043_,
    new_B6042_, new_B6041_, new_B6040_, new_B6039_, new_B6038_, new_B6037_,
    new_B6036_, new_B6035_, new_B6034_, new_B6033_, new_B6032_, new_B6031_,
    new_B6030_, new_B6029_, new_B6028_, new_B6027_, new_B6020_, new_B6019_,
    new_B6018_, new_B6017_, new_B6016_, new_B6015_, new_B6014_, new_B6013_,
    new_B6012_, new_B6011_, new_B6010_, new_B6009_, new_B6008_, new_B6007_,
    new_B6006_, new_B6005_, new_B6004_, new_B6003_, new_B6002_, new_B6001_,
    new_B6000_, new_B5999_, new_B5998_, new_B5997_, new_B5996_, new_B5995_,
    new_B5994_, new_B5993_, new_B5992_, new_B5991_, new_B5990_, new_B5989_,
    new_B5988_, new_B5987_, new_B5986_, new_B5985_, new_B5984_, new_B5983_,
    new_B5982_, new_B5981_, new_B5980_, new_B5979_, new_B5978_, new_B5977_,
    new_B5976_, new_B5975_, new_B5974_, new_B5973_, new_B5972_, new_B5971_,
    new_B5970_, new_B5969_, new_B5968_, new_B5967_, new_B5966_, new_B5965_,
    new_B5964_, new_B5963_, new_B5962_, new_B5961_, new_B5960_, new_B5953_,
    new_B5952_, new_B5951_, new_B5950_, new_B5949_, new_B5948_, new_B5947_,
    new_B5946_, new_B5945_, new_B5944_, new_B5943_, new_B5942_, new_B5941_,
    new_B5940_, new_B5939_, new_B5938_, new_B5937_, new_B5936_, new_B5935_,
    new_B5934_, new_B5933_, new_B5932_, new_B5931_, new_B5930_, new_B5929_,
    new_B5928_, new_B5927_, new_B5926_, new_B5925_, new_B5924_, new_B5923_,
    new_B5922_, new_B5921_, new_B5920_, new_B5919_, new_B5918_, new_B5917_,
    new_B5916_, new_B5915_, new_B5914_, new_B5913_, new_B5912_, new_B5911_,
    new_B5910_, new_B5909_, new_B5908_, new_B5907_, new_B5906_, new_B5905_,
    new_B5904_, new_B5903_, new_B5902_, new_B5901_, new_B5900_, new_B5899_,
    new_B5898_, new_B5897_, new_B5896_, new_B5895_, new_B5894_, new_B5893_,
    new_B5886_, new_B5885_, new_B5884_, new_B5883_, new_B5882_, new_B5881_,
    new_B5880_, new_B5879_, new_B5878_, new_B5877_, new_B5876_, new_B5875_,
    new_B5874_, new_B5873_, new_B5872_, new_B5871_, new_B5870_, new_B5869_,
    new_B5868_, new_B5867_, new_B5866_, new_B5865_, new_B5864_, new_B5863_,
    new_B5862_, new_B5861_, new_B5860_, new_B5859_, new_B5858_, new_B5857_,
    new_B5856_, new_B5855_, new_B5854_, new_B5853_, new_B5852_, new_B5851_,
    new_B5850_, new_B5849_, new_B5848_, new_B5847_, new_B5846_, new_B5845_,
    new_B5844_, new_B5843_, new_B5842_, new_B5841_, new_B5840_, new_B5839_,
    new_B5838_, new_B5837_, new_B5836_, new_B5835_, new_B5834_, new_B5833_,
    new_B5832_, new_B5831_, new_B5830_, new_B5829_, new_B5828_, new_B5827_,
    new_B5826_, new_B5819_, new_B5818_, new_B5817_, new_B5816_, new_B5815_,
    new_B5814_, new_B5813_, new_B5812_, new_B5811_, new_B5810_, new_B5809_,
    new_B5808_, new_B5807_, new_B5806_, new_B5805_, new_B5804_, new_B5803_,
    new_B5802_, new_B5801_, new_B5800_, new_B5799_, new_B5798_, new_B5797_,
    new_B5796_, new_B5795_, new_B5794_, new_B5793_, new_B5792_, new_B5791_,
    new_B5790_, new_B5789_, new_B5788_, new_B5787_, new_B5786_, new_B5785_,
    new_B5784_, new_B5783_, new_B5782_, new_B5781_, new_B5780_, new_B5779_,
    new_B5778_, new_B5777_, new_B5776_, new_B5775_, new_B5774_, new_B5773_,
    new_B5772_, new_B5771_, new_B5770_, new_B5769_, new_B5768_, new_B5767_,
    new_B5766_, new_B5765_, new_B5764_, new_B5763_, new_B5762_, new_B5761_,
    new_B5760_, new_B5759_, new_B5752_, new_B5751_, new_B5750_, new_B5749_,
    new_B5748_, new_B5747_, new_B5746_, new_B5745_, new_B5744_, new_B5743_,
    new_B5742_, new_B5741_, new_B5740_, new_B5739_, new_B5738_, new_B5737_,
    new_B5736_, new_B5735_, new_B5734_, new_B5733_, new_B5732_, new_B5731_,
    new_B5730_, new_B5729_, new_B5728_, new_B5727_, new_B5726_, new_B5725_,
    new_B5724_, new_B5723_, new_B5722_, new_B5721_, new_B5720_, new_B5719_,
    new_B5718_, new_B5717_, new_B5716_, new_B5715_, new_B5714_, new_B5713_,
    new_B5712_, new_B5711_, new_B5710_, new_B5709_, new_B5708_, new_B5707_,
    new_B5706_, new_B5705_, new_B5704_, new_B5703_, new_B5702_, new_B5701_,
    new_B5700_, new_B5699_, new_B5698_, new_B5697_, new_B5696_, new_B5695_,
    new_B5694_, new_B5693_, new_B5692_, new_B5685_, new_B5684_, new_B5683_,
    new_B5682_, new_B5681_, new_B5680_, new_B5679_, new_B5678_, new_B5677_,
    new_B5676_, new_B5675_, new_B5674_, new_B5673_, new_B5672_, new_B5671_,
    new_B5670_, new_B5669_, new_B5668_, new_B5667_, new_B5666_, new_B5665_,
    new_B5664_, new_B5663_, new_B5662_, new_B5661_, new_B5660_, new_B5659_,
    new_B5658_, new_B5657_, new_B5656_, new_B5655_, new_B5654_, new_B5653_,
    new_B5652_, new_B5651_, new_B5650_, new_B5649_, new_B5648_, new_B5647_,
    new_B5646_, new_B5645_, new_B5644_, new_B5643_, new_B5642_, new_B5641_,
    new_B5640_, new_B5639_, new_B5638_, new_B5637_, new_B5636_, new_B5635_,
    new_B5634_, new_B5633_, new_B5632_, new_B5631_, new_B5630_, new_B5629_,
    new_B5628_, new_B5627_, new_B5626_, new_B5625_, new_B5618_, new_B5617_,
    new_B5616_, new_B5615_, new_B5614_, new_B5613_, new_B5612_, new_B5611_,
    new_B5610_, new_B5609_, new_B5608_, new_B5607_, new_B5606_, new_B5605_,
    new_B5604_, new_B5603_, new_B5602_, new_B5601_, new_B5600_, new_B5599_,
    new_B5598_, new_B5597_, new_B5596_, new_B5595_, new_B5594_, new_B5593_,
    new_B5592_, new_B5591_, new_B5590_, new_B5589_, new_B5588_, new_B5587_,
    new_B5586_, new_B5585_, new_B5584_, new_B5583_, new_B5582_, new_B5581_,
    new_B5580_, new_B5579_, new_B5578_, new_B5577_, new_B5576_, new_B5575_,
    new_B5574_, new_B5573_, new_B5572_, new_B5571_, new_B5570_, new_B5569_,
    new_B5568_, new_B5567_, new_B5566_, new_B5565_, new_B5564_, new_B5563_,
    new_B5562_, new_B5561_, new_B5560_, new_B5559_, new_B5558_, new_B5551_,
    new_B5550_, new_B5549_, new_B5548_, new_B5547_, new_B5546_, new_B5545_,
    new_B5544_, new_B5543_, new_B5542_, new_B5541_, new_B5540_, new_B5539_,
    new_B5538_, new_B5537_, new_B5536_, new_B5535_, new_B5534_, new_B5533_,
    new_B5532_, new_B5531_, new_B5530_, new_B5529_, new_B5528_, new_B5527_,
    new_B5526_, new_B5525_, new_B5524_, new_B5523_, new_B5522_, new_B5521_,
    new_B5520_, new_B5519_, new_B5518_, new_B5517_, new_B5516_, new_B5515_,
    new_B5514_, new_B5513_, new_B5512_, new_B5511_, new_B5510_, new_B5509_,
    new_B5508_, new_B5507_, new_B5506_, new_B5505_, new_B5504_, new_B5503_,
    new_B5502_, new_B5501_, new_B5500_, new_B5499_, new_B5498_, new_B5497_,
    new_B5496_, new_B5495_, new_B5494_, new_B5493_, new_B5492_, new_B5491_,
    new_B5484_, new_B5483_, new_B5482_, new_B5481_, new_B5480_, new_B5479_,
    new_B5478_, new_B5477_, new_B5476_, new_B5475_, new_B5474_, new_B5473_,
    new_B5472_, new_B5471_, new_B5470_, new_B5469_, new_B5468_, new_B5467_,
    new_B5466_, new_B5465_, new_B5464_, new_B5463_, new_B5462_, new_B5461_,
    new_B5460_, new_B5459_, new_B5458_, new_B5457_, new_B5456_, new_B5455_,
    new_B5454_, new_B5453_, new_B5452_, new_B5451_, new_B5450_, new_B5449_,
    new_B5448_, new_B5447_, new_B5446_, new_B5445_, new_B5444_, new_B5443_,
    new_B5442_, new_B5441_, new_B5440_, new_B5439_, new_B5438_, new_B5437_,
    new_B5436_, new_B5435_, new_B5434_, new_B5433_, new_B5432_, new_B5431_,
    new_B5430_, new_B5429_, new_B5428_, new_B5427_, new_B5426_, new_B5425_,
    new_B5424_, new_B5417_, new_B5416_, new_B5415_, new_B5414_, new_B5413_,
    new_B5412_, new_B5411_, new_B5410_, new_B5409_, new_B5408_, new_B5407_,
    new_B5406_, new_B5405_, new_B5404_, new_B5403_, new_B5402_, new_B5401_,
    new_B5400_, new_B5399_, new_B5398_, new_B5397_, new_B5396_, new_B5395_,
    new_B5394_, new_B5393_, new_B5392_, new_B5391_, new_B5390_, new_B5389_,
    new_B5388_, new_B5387_, new_B5386_, new_B5385_, new_B5384_, new_B5383_,
    new_B5382_, new_B5381_, new_B5380_, new_B5379_, new_B5378_, new_B5377_,
    new_B5376_, new_B5375_, new_B5374_, new_B5373_, new_B5372_, new_B5371_,
    new_B5370_, new_B5369_, new_B5368_, new_B5367_, new_B5366_, new_B5365_,
    new_B5364_, new_B5363_, new_B5362_, new_B5361_, new_B5360_, new_B5359_,
    new_B5358_, new_B5357_, new_B5350_, new_B5349_, new_B5348_, new_B5347_,
    new_B5346_, new_B5345_, new_B5344_, new_B5343_, new_B5342_, new_B5341_,
    new_B5340_, new_B5339_, new_B5338_, new_B5337_, new_B5336_, new_B5335_,
    new_B5334_, new_B5333_, new_B5332_, new_B5331_, new_B5330_, new_B5329_,
    new_B5328_, new_B5327_, new_B5326_, new_B5325_, new_B5324_, new_B5323_,
    new_B5322_, new_B5321_, new_B5320_, new_B5319_, new_B5318_, new_B5317_,
    new_B5316_, new_B5315_, new_B5314_, new_B5313_, new_B5312_, new_B5311_,
    new_B5310_, new_B5309_, new_B5308_, new_B5307_, new_B5306_, new_B5305_,
    new_B5304_, new_B5303_, new_B5302_, new_B5301_, new_B5300_, new_B5299_,
    new_B5298_, new_B5297_, new_B5296_, new_B5295_, new_B5294_, new_B5293_,
    new_B5292_, new_B5291_, new_B5290_, new_B5283_, new_B5282_, new_B5281_,
    new_B5280_, new_B5279_, new_B5278_, new_B5277_, new_B5276_, new_B5275_,
    new_B5274_, new_B5273_, new_B5272_, new_B5271_, new_B5270_, new_B5269_,
    new_B5268_, new_B5267_, new_B5266_, new_B5265_, new_B5264_, new_B5263_,
    new_B5262_, new_B5261_, new_B5260_, new_B5259_, new_B5258_, new_B5257_,
    new_B5256_, new_B5255_, new_B5254_, new_B5253_, new_B5252_, new_B5251_,
    new_B5250_, new_B5249_, new_B5248_, new_B5247_, new_B5246_, new_B5245_,
    new_B5244_, new_B5243_, new_B5242_, new_B5241_, new_B5240_, new_B5239_,
    new_B5238_, new_B5237_, new_B5236_, new_B5235_, new_B5234_, new_B5233_,
    new_B5232_, new_B5231_, new_B5230_, new_B5229_, new_B5228_, new_B5227_,
    new_B5226_, new_B5225_, new_B5224_, new_B5223_, new_B5216_, new_B5215_,
    new_B5214_, new_B5213_, new_B5212_, new_B5211_, new_B5210_, new_B5209_,
    new_B5208_, new_B5207_, new_B5206_, new_B5205_, new_B5204_, new_B5203_,
    new_B5202_, new_B5201_, new_B5200_, new_B5199_, new_B5198_, new_B5197_,
    new_B5196_, new_B5195_, new_B5194_, new_B5193_, new_B5192_, new_B5191_,
    new_B5190_, new_B5189_, new_B5188_, new_B5187_, new_B5186_, new_B5185_,
    new_B5184_, new_B5183_, new_B5182_, new_B5181_, new_B5180_, new_B5179_,
    new_B5178_, new_B5177_, new_B5176_, new_B5175_, new_B5174_, new_B5173_,
    new_B5172_, new_B5171_, new_B5170_, new_B5169_, new_B5168_, new_B5167_,
    new_B5166_, new_B5165_, new_B5164_, new_B5163_, new_B5162_, new_B5161_,
    new_B5160_, new_B5159_, new_B5158_, new_B5157_, new_B5156_, new_B5149_,
    new_B5148_, new_B5147_, new_B5146_, new_B5145_, new_B5144_, new_B5143_,
    new_B5142_, new_B5141_, new_B5140_, new_B5139_, new_B5138_, new_B5137_,
    new_B5136_, new_B5135_, new_B5134_, new_B5133_, new_B5132_, new_B5131_,
    new_B5130_, new_B5129_, new_B5128_, new_B5127_, new_B5126_, new_B5125_,
    new_B5124_, new_B5123_, new_B5122_, new_B5121_, new_B5120_, new_B5119_,
    new_B5118_, new_B5117_, new_B5116_, new_B5115_, new_B5114_, new_B5113_,
    new_B5112_, new_B5111_, new_B5110_, new_B5109_, new_B5108_, new_B5107_,
    new_B5106_, new_B5105_, new_B5104_, new_B5103_, new_B5102_, new_B5101_,
    new_B5100_, new_B5099_, new_B5098_, new_B5097_, new_B5096_, new_B5095_,
    new_B5094_, new_B5093_, new_B5092_, new_B5091_, new_B5090_, new_B5089_,
    new_B5082_, new_B5081_, new_B5080_, new_B5079_, new_B5078_, new_B5077_,
    new_B5076_, new_B5075_, new_B5074_, new_B5073_, new_B5072_, new_B5071_,
    new_B5070_, new_B5069_, new_B5068_, new_B5067_, new_B5066_, new_B5065_,
    new_B5064_, new_B5063_, new_B5062_, new_B5061_, new_B5060_, new_B5059_,
    new_B5058_, new_B5057_, new_B5056_, new_B5055_, new_B5054_, new_B5053_,
    new_B5052_, new_B5051_, new_B5050_, new_B5049_, new_B5048_, new_B5047_,
    new_B5046_, new_B5045_, new_B5044_, new_B5043_, new_B5042_, new_B5041_,
    new_B5040_, new_B5039_, new_B5038_, new_B5037_, new_B5036_, new_B5035_,
    new_B5034_, new_B5033_, new_B5032_, new_B5031_, new_B5030_, new_B5029_,
    new_B5028_, new_B5027_, new_B5026_, new_B5025_, new_B5024_, new_B5023_,
    new_B5022_, new_B5015_, new_B5014_, new_B5013_, new_B5012_, new_B5011_,
    new_B5010_, new_B5009_, new_B5008_, new_B5007_, new_B5006_, new_B5005_,
    new_B5004_, new_B5003_, new_B5002_, new_B5001_, new_B5000_, new_B4999_,
    new_B4998_, new_B4997_, new_B4996_, new_B4995_, new_B4994_, new_B4993_,
    new_B4992_, new_B4991_, new_B4990_, new_B4989_, new_B4988_, new_B4987_,
    new_B4986_, new_B4985_, new_B4984_, new_B4983_, new_B4982_, new_B4981_,
    new_B4980_, new_B4979_, new_B4978_, new_B4977_, new_B4976_, new_B4975_,
    new_B4974_, new_B4973_, new_B4972_, new_B4971_, new_B4970_, new_B4969_,
    new_B4968_, new_B4967_, new_B4966_, new_B4965_, new_B4964_, new_B4963_,
    new_B4962_, new_B4961_, new_B4960_, new_B4959_, new_B4958_, new_B4957_,
    new_B4956_, new_B4955_, new_B4948_, new_B4947_, new_B4946_, new_B4945_,
    new_B4944_, new_B4943_, new_B4942_, new_B4941_, new_B4940_, new_B4939_,
    new_B4938_, new_B4937_, new_B4936_, new_B4935_, new_B4934_, new_B4933_,
    new_B4932_, new_B4931_, new_B4930_, new_B4929_, new_B4928_, new_B4927_,
    new_B4926_, new_B4925_, new_B4924_, new_B4923_, new_B4922_, new_B4921_,
    new_B4920_, new_B4919_, new_B4918_, new_B4917_, new_B4916_, new_B4915_,
    new_B4914_, new_B4913_, new_B4912_, new_B4911_, new_B4910_, new_B4909_,
    new_B4908_, new_B4907_, new_B4906_, new_B4905_, new_B4904_, new_B4903_,
    new_B4902_, new_B4901_, new_B4900_, new_B4899_, new_B4898_, new_B4897_,
    new_B4896_, new_B4895_, new_B4894_, new_B4893_, new_B4892_, new_B4891_,
    new_B4890_, new_B4889_, new_B4888_, new_B4881_, new_B4880_, new_B4879_,
    new_B4878_, new_B4877_, new_B4876_, new_B4875_, new_B4874_, new_B4873_,
    new_B4872_, new_B4871_, new_B4870_, new_B4869_, new_B4868_, new_B4867_,
    new_B4866_, new_B4865_, new_B4864_, new_B4863_, new_B4862_, new_B4861_,
    new_B4860_, new_B4859_, new_B4858_, new_B4857_, new_B4856_, new_B4855_,
    new_B4854_, new_B4853_, new_B4852_, new_B4851_, new_B4850_, new_B4849_,
    new_B4848_, new_B4847_, new_B4846_, new_B4845_, new_B4844_, new_B4843_,
    new_B4842_, new_B4841_, new_B4840_, new_B4839_, new_B4838_, new_B4837_,
    new_B4836_, new_B4835_, new_B4834_, new_B4833_, new_B4832_, new_B4831_,
    new_B4830_, new_B4829_, new_B4828_, new_B4827_, new_B4826_, new_B4825_,
    new_B4824_, new_B4823_, new_B4822_, new_B4821_, new_B4814_, new_B4813_,
    new_B4812_, new_B4811_, new_B4810_, new_B4809_, new_B4808_, new_B4807_,
    new_B4806_, new_B4805_, new_B4804_, new_B4803_, new_B4802_, new_B4801_,
    new_B4800_, new_B4799_, new_B4798_, new_B4797_, new_B4796_, new_B4795_,
    new_B4794_, new_B4793_, new_B4792_, new_B4791_, new_B4790_, new_B4789_,
    new_B4788_, new_B4787_, new_B4786_, new_B4785_, new_B4784_, new_B4783_,
    new_B4782_, new_B4781_, new_B4780_, new_B4779_, new_B4778_, new_B4777_,
    new_B4776_, new_B4775_, new_B4774_, new_B4773_, new_B4772_, new_B4771_,
    new_B4770_, new_B4769_, new_B4768_, new_B4767_, new_B4766_, new_B4765_,
    new_B4764_, new_B4763_, new_B4762_, new_B4761_, new_B4760_, new_B4759_,
    new_B4758_, new_B4757_, new_B4756_, new_B4755_, new_B4754_, new_B4747_,
    new_B4746_, new_B4745_, new_B4744_, new_B4743_, new_B4742_, new_B4741_,
    new_B4740_, new_B4739_, new_B4738_, new_B4737_, new_B4736_, new_B4735_,
    new_B4734_, new_B4733_, new_B4732_, new_B4731_, new_B4730_, new_B4729_,
    new_B4728_, new_B4727_, new_B4726_, new_B4725_, new_B4724_, new_B4723_,
    new_B4722_, new_B4721_, new_B4720_, new_B4719_, new_B4718_, new_B4717_,
    new_B4716_, new_B4715_, new_B4714_, new_B4713_, new_B4712_, new_B4711_,
    new_B4710_, new_B4709_, new_B4708_, new_B4707_, new_B4706_, new_B4705_,
    new_B4704_, new_B4703_, new_B4702_, new_B4701_, new_B4700_, new_B4699_,
    new_B4698_, new_B4697_, new_B4696_, new_B4695_, new_B4694_, new_B4693_,
    new_B4692_, new_B4691_, new_B4690_, new_B4689_, new_B4688_, new_B4687_,
    new_B4680_, new_B4679_, new_B4678_, new_B4677_, new_B4676_, new_B4675_,
    new_B4674_, new_B4673_, new_B4672_, new_B4671_, new_B4670_, new_B4669_,
    new_B4668_, new_B4667_, new_B4666_, new_B4665_, new_B4664_, new_B4663_,
    new_B4662_, new_B4661_, new_B4660_, new_B4659_, new_B4658_, new_B4657_,
    new_B4656_, new_B4655_, new_B4654_, new_B4653_, new_B4652_, new_B4651_,
    new_B4650_, new_B4649_, new_B4648_, new_B4647_, new_B4646_, new_B4645_,
    new_B4644_, new_B4643_, new_B4642_, new_B4641_, new_B4640_, new_B4639_,
    new_B4638_, new_B4637_, new_B4636_, new_B4635_, new_B4634_, new_B4633_,
    new_B4632_, new_B4631_, new_B4630_, new_B4629_, new_B4628_, new_B4627_,
    new_B4626_, new_B4625_, new_B4624_, new_B4623_, new_B4622_, new_B4621_,
    new_B4620_, new_B4613_, new_B4612_, new_B4611_, new_B4610_, new_B4609_,
    new_B4608_, new_B4607_, new_B4606_, new_B4605_, new_B4604_, new_B4603_,
    new_B4602_, new_B4601_, new_B4600_, new_B4599_, new_B4598_, new_B4597_,
    new_B4596_, new_B4595_, new_B4594_, new_B4593_, new_B4592_, new_B4591_,
    new_B4590_, new_B4589_, new_B4588_, new_B4587_, new_B4586_, new_B4585_,
    new_B4584_, new_B4583_, new_B4582_, new_B4581_, new_B4580_, new_B4579_,
    new_B4578_, new_B4577_, new_B4576_, new_B4575_, new_B4574_, new_B4573_,
    new_B4572_, new_B4571_, new_B4570_, new_B4569_, new_B4568_, new_B4567_,
    new_B4566_, new_B4565_, new_B4564_, new_B4563_, new_B4562_, new_B4561_,
    new_B4560_, new_B4559_, new_B4558_, new_B4557_, new_B4556_, new_B4555_,
    new_B4554_, new_B4553_, new_B4546_, new_B4545_, new_B4544_, new_B4543_,
    new_B4542_, new_B4541_, new_B4540_, new_B4539_, new_B4538_, new_B4537_,
    new_B4536_, new_B4535_, new_B4534_, new_B4533_, new_B4532_, new_B4531_,
    new_B4530_, new_B4529_, new_B4528_, new_B4527_, new_B4526_, new_B4525_,
    new_B4524_, new_B4523_, new_B4522_, new_B4521_, new_B4520_, new_B4519_,
    new_B4518_, new_B4517_, new_B4516_, new_B4515_, new_B4514_, new_B4513_,
    new_B4512_, new_B4511_, new_B4510_, new_B4509_, new_B4508_, new_B4507_,
    new_B4506_, new_B4505_, new_B4504_, new_B4503_, new_B4502_, new_B4501_,
    new_B4500_, new_B4499_, new_B4498_, new_B4497_, new_B4496_, new_B4495_,
    new_B4494_, new_B4493_, new_B4492_, new_B4491_, new_B4490_, new_B4489_,
    new_B4488_, new_B4487_, new_B4486_, new_B4479_, new_B4478_, new_B4477_,
    new_B4476_, new_B4475_, new_B4474_, new_B4473_, new_B4472_, new_B4471_,
    new_B4470_, new_B4469_, new_B4468_, new_B4467_, new_B4466_, new_B4465_,
    new_B4464_, new_B4463_, new_B4462_, new_B4461_, new_B4460_, new_B4459_,
    new_B4458_, new_B4457_, new_B4456_, new_B4455_, new_B4454_, new_B4453_,
    new_B4452_, new_B4451_, new_B4450_, new_B4449_, new_B4448_, new_B4447_,
    new_B4446_, new_B4445_, new_B4444_, new_B4443_, new_B4442_, new_B4441_,
    new_B4440_, new_B4439_, new_B4438_, new_B4437_, new_B4436_, new_B4435_,
    new_B4434_, new_B4433_, new_B4432_, new_B4431_, new_B4430_, new_B4429_,
    new_B4428_, new_B4427_, new_B4426_, new_B4425_, new_B4424_, new_B4423_,
    new_B4422_, new_B4421_, new_B4420_, new_B4419_, new_B4412_, new_B4411_,
    new_B4410_, new_B4409_, new_B4408_, new_B4407_, new_B4406_, new_B4405_,
    new_B4404_, new_B4403_, new_B4402_, new_B4401_, new_B4400_, new_B4399_,
    new_B4398_, new_B4397_, new_B4396_, new_B4395_, new_B4394_, new_B4393_,
    new_B4392_, new_B4391_, new_B4390_, new_B4389_, new_B4388_, new_B4387_,
    new_B4386_, new_B4385_, new_B4384_, new_B4383_, new_B4382_, new_B4381_,
    new_B4380_, new_B4379_, new_B4378_, new_B4377_, new_B4376_, new_B4375_,
    new_B4374_, new_B4373_, new_B4372_, new_B4371_, new_B4370_, new_B4369_,
    new_B4368_, new_B4367_, new_B4366_, new_B4365_, new_B4364_, new_B4363_,
    new_B4362_, new_B4361_, new_B4360_, new_B4359_, new_B4358_, new_B4357_,
    new_B4356_, new_B4355_, new_B4354_, new_B4353_, new_B4352_, new_B4345_,
    new_B4344_, new_B4343_, new_B4342_, new_B4341_, new_B4340_, new_B4339_,
    new_B4338_, new_B4337_, new_B4336_, new_B4335_, new_B4334_, new_B4333_,
    new_B4332_, new_B4331_, new_B4330_, new_B4329_, new_B4328_, new_B4327_,
    new_B4326_, new_B4325_, new_B4324_, new_B4323_, new_B4322_, new_B4321_,
    new_B4320_, new_B4319_, new_B4318_, new_B4317_, new_B4316_, new_B4315_,
    new_B4314_, new_B4313_, new_B4312_, new_B4311_, new_B4310_, new_B4309_,
    new_B4308_, new_B4307_, new_B4306_, new_B4305_, new_B4304_, new_B4303_,
    new_B4302_, new_B4301_, new_B4300_, new_B4299_, new_B4298_, new_B4297_,
    new_B4296_, new_B4295_, new_B4294_, new_B4293_, new_B4292_, new_B4291_,
    new_B4290_, new_B4289_, new_B4288_, new_B4287_, new_B4286_, new_B4285_,
    new_B4278_, new_B4277_, new_B4276_, new_B4275_, new_B4274_, new_B4273_,
    new_B4272_, new_B4271_, new_B4270_, new_B4269_, new_B4268_, new_B4267_,
    new_B4266_, new_B4265_, new_B4264_, new_B4263_, new_B4262_, new_B4261_,
    new_B4260_, new_B4259_, new_B4258_, new_B4257_, new_B4256_, new_B4255_,
    new_B4254_, new_B4253_, new_B4252_, new_B4251_, new_B4250_, new_B4249_,
    new_B4248_, new_B4247_, new_B4246_, new_B4245_, new_B4244_, new_B4243_,
    new_B4242_, new_B4241_, new_B4240_, new_B4239_, new_B4238_, new_B4237_,
    new_B4236_, new_B4235_, new_B4234_, new_B4233_, new_B4232_, new_B4231_,
    new_B4230_, new_B4229_, new_B4228_, new_B4227_, new_B4226_, new_B4225_,
    new_B4224_, new_B4223_, new_B4222_, new_B4221_, new_B4220_, new_B4219_,
    new_B4218_, new_B4211_, new_B4210_, new_B4209_, new_B4208_, new_B4207_,
    new_B4206_, new_B4205_, new_B4204_, new_B4203_, new_B4202_, new_B4201_,
    new_B4200_, new_B4199_, new_B4198_, new_B4197_, new_B4196_, new_B4195_,
    new_B4194_, new_B4193_, new_B4192_, new_B4191_, new_B4190_, new_B4189_,
    new_B4188_, new_B4187_, new_B4186_, new_B4185_, new_B4184_, new_B4183_,
    new_B4182_, new_B4181_, new_B4180_, new_B4179_, new_B4178_, new_B4177_,
    new_B4176_, new_B4175_, new_B4174_, new_B4173_, new_B4172_, new_B4171_,
    new_B4170_, new_B4169_, new_B4168_, new_B4167_, new_B4166_, new_B4165_,
    new_B4164_, new_B4163_, new_B4162_, new_B4161_, new_B4160_, new_B4159_,
    new_B4158_, new_B4157_, new_B4156_, new_B4155_, new_B4154_, new_B4153_,
    new_B4152_, new_B4151_, new_B4144_, new_B4143_, new_B4142_, new_B4141_,
    new_B4140_, new_B4139_, new_B4138_, new_B4137_, new_B4136_, new_B4135_,
    new_B4134_, new_B4133_, new_B4132_, new_B4131_, new_B4130_, new_B4129_,
    new_B4128_, new_B4127_, new_B4126_, new_B4125_, new_B4124_, new_B4123_,
    new_B4122_, new_B4121_, new_B4120_, new_B4119_, new_B4118_, new_B4117_,
    new_B4116_, new_B4115_, new_B4114_, new_B4113_, new_B4112_, new_B4111_,
    new_B4110_, new_B4109_, new_B4108_, new_B4107_, new_B4106_, new_B4105_,
    new_B4104_, new_B4103_, new_B4102_, new_B4101_, new_B4100_, new_B4099_,
    new_B4098_, new_B4097_, new_B4096_, new_B4095_, new_B4094_, new_B4093_,
    new_B4092_, new_B4091_, new_B4090_, new_B4089_, new_B4088_, new_B4087_,
    new_B4086_, new_B4085_, new_B4084_, new_B4077_, new_B4076_, new_B4075_,
    new_B4074_, new_B4073_, new_B4072_, new_B4071_, new_B4070_, new_B4069_,
    new_B4068_, new_B4067_, new_B4066_, new_B4065_, new_B4064_, new_B4063_,
    new_B4062_, new_B4061_, new_B4060_, new_B4059_, new_B4058_, new_B4057_,
    new_B4056_, new_B4055_, new_B4054_, new_B4053_, new_B4052_, new_B4051_,
    new_B4050_, new_B4049_, new_B4048_, new_B4047_, new_B4046_, new_B4045_,
    new_B4044_, new_B4043_, new_B4042_, new_B4041_, new_B4040_, new_B4039_,
    new_B4038_, new_B4037_, new_B4036_, new_B4035_, new_B4034_, new_B4033_,
    new_B4032_, new_B4031_, new_B4030_, new_B4029_, new_B4028_, new_B4027_,
    new_B4026_, new_B4025_, new_B4024_, new_B4023_, new_B4022_, new_B4021_,
    new_B4020_, new_B4019_, new_B4018_, new_B4017_, new_B4010_, new_B4009_,
    new_B4008_, new_B4007_, new_B4006_, new_B4005_, new_B4004_, new_B4003_,
    new_B4002_, new_B4001_, new_B4000_, new_B3999_, new_B3998_, new_B3997_,
    new_B3996_, new_B3995_, new_B3994_, new_B3993_, new_B3992_, new_B3991_,
    new_B3990_, new_B3989_, new_B3988_, new_B3987_, new_B3986_, new_B3985_,
    new_B3984_, new_B3983_, new_B3982_, new_B3981_, new_B3980_, new_B3979_,
    new_B3978_, new_B3977_, new_B3976_, new_B3975_, new_B3974_, new_B3973_,
    new_B3972_, new_B3971_, new_B3970_, new_B3969_, new_B3968_, new_B3967_,
    new_B3966_, new_B3965_, new_B3964_, new_B3963_, new_B3962_, new_B3961_,
    new_B3960_, new_B3959_, new_B3958_, new_B3957_, new_B3956_, new_B3955_,
    new_B3954_, new_B3953_, new_B3952_, new_B3951_, new_B3950_, new_B3943_,
    new_B3942_, new_B3941_, new_B3940_, new_B3939_, new_B3938_, new_B3937_,
    new_B3936_, new_B3935_, new_B3934_, new_B3933_, new_B3932_, new_B3931_,
    new_B3930_, new_B3929_, new_B3928_, new_B3927_, new_B3926_, new_B3925_,
    new_B3924_, new_B3923_, new_B3922_, new_B3921_, new_B3920_, new_B3919_,
    new_B3918_, new_B3917_, new_B3916_, new_B3915_, new_B3914_, new_B3913_,
    new_B3912_, new_B3911_, new_B3910_, new_B3909_, new_B3908_, new_B3907_,
    new_B3906_, new_B3905_, new_B3904_, new_B3903_, new_B3902_, new_B3901_,
    new_B3900_, new_B3899_, new_B3898_, new_B3897_, new_B3896_, new_B3895_,
    new_B3894_, new_B3893_, new_B3892_, new_B3891_, new_B3890_, new_B3889_,
    new_B3888_, new_B3887_, new_B3886_, new_B3885_, new_B3884_, new_B3883_,
    new_B3876_, new_B3875_, new_B3874_, new_B3873_, new_B3872_, new_B3871_,
    new_B3870_, new_B3869_, new_B3868_, new_B3867_, new_B3866_, new_B3865_,
    new_B3864_, new_B3863_, new_B3862_, new_B3861_, new_B3860_, new_B3859_,
    new_B3858_, new_B3857_, new_B3856_, new_B3855_, new_B3854_, new_B3853_,
    new_B3852_, new_B3851_, new_B3850_, new_B3849_, new_B3848_, new_B3847_,
    new_B3846_, new_B3845_, new_B3844_, new_B3843_, new_B3842_, new_B3841_,
    new_B3840_, new_B3839_, new_B3838_, new_B3837_, new_B3836_, new_B3835_,
    new_B3834_, new_B3833_, new_B3832_, new_B3831_, new_B3830_, new_B3829_,
    new_B3828_, new_B3827_, new_B3826_, new_B3825_, new_B3824_, new_B3823_,
    new_B3822_, new_B3821_, new_B3820_, new_B3819_, new_B3818_, new_B3817_,
    new_B3816_, new_B3809_, new_B3808_, new_B3807_, new_B3806_, new_B3805_,
    new_B3804_, new_B3803_, new_B3802_, new_B3801_, new_B3800_, new_B3799_,
    new_B3798_, new_B3797_, new_B3796_, new_B3795_, new_B3794_, new_B3793_,
    new_B3792_, new_B3791_, new_B3790_, new_B3789_, new_B3788_, new_B3787_,
    new_B3786_, new_B3785_, new_B3784_, new_B3783_, new_B3782_, new_B3781_,
    new_B3780_, new_B3779_, new_B3778_, new_B3777_, new_B3776_, new_B3775_,
    new_B3774_, new_B3773_, new_B3772_, new_B3771_, new_B3770_, new_B3769_,
    new_B3768_, new_B3767_, new_B3766_, new_B3765_, new_B3764_, new_B3763_,
    new_B3762_, new_B3761_, new_B3760_, new_B3759_, new_B3758_, new_B3757_,
    new_B3756_, new_B3755_, new_B3754_, new_B3753_, new_B3752_, new_B3751_,
    new_B3750_, new_B3749_, new_B3742_, new_B3741_, new_B3740_, new_B3739_,
    new_B3738_, new_B3737_, new_B3736_, new_B3735_, new_B3734_, new_B3733_,
    new_B3732_, new_B3731_, new_B3730_, new_B3729_, new_B3728_, new_B3727_,
    new_B3726_, new_B3725_, new_B3724_, new_B3723_, new_B3722_, new_B3721_,
    new_B3720_, new_B3719_, new_B3718_, new_B3717_, new_B3716_, new_B3715_,
    new_B3714_, new_B3713_, new_B3712_, new_B3711_, new_B3710_, new_B3709_,
    new_B3708_, new_B3707_, new_B3706_, new_B3705_, new_B3704_, new_B3703_,
    new_B3702_, new_B3701_, new_B3700_, new_B3699_, new_B3698_, new_B3697_,
    new_B3696_, new_B3695_, new_B3694_, new_B3693_, new_B3692_, new_B3691_,
    new_B3690_, new_B3689_, new_B3688_, new_B3687_, new_B3686_, new_B3685_,
    new_B3684_, new_B3683_, new_B3682_, new_B3675_, new_B3674_, new_B3673_,
    new_B3672_, new_B3671_, new_B3670_, new_B3669_, new_B3668_, new_B3667_,
    new_B3666_, new_B3665_, new_B3664_, new_B3663_, new_B3662_, new_B3661_,
    new_B3660_, new_B3659_, new_B3658_, new_B3657_, new_B3656_, new_B3655_,
    new_B3654_, new_B3653_, new_B3652_, new_B3651_, new_B3650_, new_B3649_,
    new_B3648_, new_B3647_, new_B3646_, new_B3645_, new_B3644_, new_B3643_,
    new_B3642_, new_B3641_, new_B3640_, new_B3639_, new_B3638_, new_B3637_,
    new_B3636_, new_B3635_, new_B3634_, new_B3633_, new_B3632_, new_B3631_,
    new_B3630_, new_B3629_, new_B3628_, new_B3627_, new_B3626_, new_B3625_,
    new_B3624_, new_B3623_, new_B3622_, new_B3621_, new_B3620_, new_B3619_,
    new_B3618_, new_B3617_, new_B3616_, new_B3615_, new_B3608_, new_B3607_,
    new_B3606_, new_B3605_, new_B3604_, new_B3603_, new_B3602_, new_B3601_,
    new_B3600_, new_B3599_, new_B3598_, new_B3597_, new_B3596_, new_B3595_,
    new_B3594_, new_B3593_, new_B3592_, new_B3591_, new_B3590_, new_B3589_,
    new_B3588_, new_B3587_, new_B3586_, new_B3585_, new_B3584_, new_B3583_,
    new_B3582_, new_B3581_, new_B3580_, new_B3579_, new_B3578_, new_B3577_,
    new_B3576_, new_B3575_, new_B3574_, new_B3573_, new_B3572_, new_B3571_,
    new_B3570_, new_B3569_, new_B3568_, new_B3567_, new_B3566_, new_B3565_,
    new_B3564_, new_B3563_, new_B3562_, new_B3561_, new_B3560_, new_B3559_,
    new_B3558_, new_B3557_, new_B3556_, new_B3555_, new_B3554_, new_B3553_,
    new_B3552_, new_B3551_, new_B3550_, new_B3549_, new_B3548_, new_B3541_,
    new_B3540_, new_B3539_, new_B3538_, new_B3537_, new_B3536_, new_B3535_,
    new_B3534_, new_B3533_, new_B3532_, new_B3531_, new_B3530_, new_B3529_,
    new_B3528_, new_B3527_, new_B3526_, new_B3525_, new_B3524_, new_B3523_,
    new_B3522_, new_B3521_, new_B3520_, new_B3519_, new_B3518_, new_B3517_,
    new_B3516_, new_B3515_, new_B3514_, new_B3513_, new_B3512_, new_B3511_,
    new_B3510_, new_B3509_, new_B3508_, new_B3507_, new_B3506_, new_B3505_,
    new_B3504_, new_B3503_, new_B3502_, new_B3501_, new_B3500_, new_B3499_,
    new_B3498_, new_B3497_, new_B3496_, new_B3495_, new_B3494_, new_B3493_,
    new_B3492_, new_B3491_, new_B3490_, new_B3489_, new_B3488_, new_B3487_,
    new_B3486_, new_B3485_, new_B3484_, new_B3483_, new_B3482_, new_B3481_,
    new_B3474_, new_B3473_, new_B3472_, new_B3471_, new_B3470_, new_B3469_,
    new_B3468_, new_B3467_, new_B3466_, new_B3465_, new_B3464_, new_B3463_,
    new_B3462_, new_B3461_, new_B3460_, new_B3459_, new_B3458_, new_B3457_,
    new_B3456_, new_B3455_, new_B3454_, new_B3453_, new_B3452_, new_B3451_,
    new_B3450_, new_B3449_, new_B3448_, new_B3447_, new_B3446_, new_B3445_,
    new_B3444_, new_B3443_, new_B3442_, new_B3441_, new_B3440_, new_B3439_,
    new_B3438_, new_B3437_, new_B3436_, new_B3435_, new_B3434_, new_B3433_,
    new_B3432_, new_B3431_, new_B3430_, new_B3429_, new_B3428_, new_B3427_,
    new_B3426_, new_B3425_, new_B3424_, new_B3423_, new_B3422_, new_B3421_,
    new_B3420_, new_B3419_, new_B3418_, new_B3417_, new_B3416_, new_B3415_,
    new_B3414_, new_B3407_, new_B3406_, new_B3405_, new_B3404_, new_B3403_,
    new_B3402_, new_B3401_, new_B3400_, new_B3399_, new_B3398_, new_B3397_,
    new_B3396_, new_B3395_, new_B3394_, new_B3393_, new_B3392_, new_B3391_,
    new_B3390_, new_B3389_, new_B3388_, new_B3387_, new_B3386_, new_B3385_,
    new_B3384_, new_B3383_, new_B3382_, new_B3381_, new_B3380_, new_B3379_,
    new_B3378_, new_B3377_, new_B3376_, new_B3375_, new_B3374_, new_B3373_,
    new_B3372_, new_B3371_, new_B3370_, new_B3369_, new_B3368_, new_B3367_,
    new_B3366_, new_B3365_, new_B3364_, new_B3363_, new_B3362_, new_B3361_,
    new_B3360_, new_B3359_, new_B3358_, new_B3357_, new_B3356_, new_B3355_,
    new_B3354_, new_B3353_, new_B3352_, new_B3351_, new_B3350_, new_B3349_,
    new_B3348_, new_B3347_, new_B3340_, new_B3339_, new_B3338_, new_B3337_,
    new_B3336_, new_B3335_, new_B3334_, new_B3333_, new_B3332_, new_B3331_,
    new_B3330_, new_B3329_, new_B3328_, new_B3327_, new_B3326_, new_B3325_,
    new_B3324_, new_B3323_, new_B3322_, new_B3321_, new_B3320_, new_B3319_,
    new_B3318_, new_B3317_, new_B3316_, new_B3315_, new_B3314_, new_B3313_,
    new_B3312_, new_B3311_, new_B3310_, new_B3309_, new_B3308_, new_B3307_,
    new_B3306_, new_B3305_, new_B3304_, new_B3303_, new_B3302_, new_B3301_,
    new_B3300_, new_B3299_, new_B3298_, new_B3297_, new_B3296_, new_B3295_,
    new_B3294_, new_B3293_, new_B3292_, new_B3291_, new_B3290_, new_B3289_,
    new_B3288_, new_B3287_, new_B3286_, new_B3285_, new_B3284_, new_B3283_,
    new_B3282_, new_B3281_, new_B3280_, new_B3273_, new_B3272_, new_B3271_,
    new_B3270_, new_B3269_, new_B3268_, new_B3267_, new_B3266_, new_B3265_,
    new_B3264_, new_B3263_, new_B3262_, new_B3261_, new_B3260_, new_B3259_,
    new_B3258_, new_B3257_, new_B3256_, new_B3255_, new_B3254_, new_B3253_,
    new_B3252_, new_B3251_, new_B3250_, new_B3249_, new_B3248_, new_B3247_,
    new_B3246_, new_B3245_, new_B3244_, new_B3243_, new_B3242_, new_B3241_,
    new_B3240_, new_B3239_, new_B3238_, new_B3237_, new_B3236_, new_B3235_,
    new_B3234_, new_B3233_, new_B3232_, new_B3231_, new_B3230_, new_B3229_,
    new_B3228_, new_B3227_, new_B3226_, new_B3225_, new_B3224_, new_B3223_,
    new_B3222_, new_B3221_, new_B3220_, new_B3219_, new_B3218_, new_B3217_,
    new_B3216_, new_B3215_, new_B3214_, new_B3213_, new_B3206_, new_B3205_,
    new_B3204_, new_B3203_, new_B3202_, new_B3201_, new_B3200_, new_B3199_,
    new_B3198_, new_B3197_, new_B3196_, new_B3195_, new_B3194_, new_B3193_,
    new_B3192_, new_B3191_, new_B3190_, new_B3189_, new_B3188_, new_B3187_,
    new_B3186_, new_B3185_, new_B3184_, new_B3183_, new_B3182_, new_B3181_,
    new_B3180_, new_B3179_, new_B3178_, new_B3177_, new_B3176_, new_B3175_,
    new_B3174_, new_B3173_, new_B3172_, new_B3171_, new_B3170_, new_B3169_,
    new_B3168_, new_B3167_, new_B3166_, new_B3165_, new_B3164_, new_B3163_,
    new_B3162_, new_B3161_, new_B3160_, new_B3159_, new_B3158_, new_B3157_,
    new_B3156_, new_B3155_, new_B3154_, new_B3153_, new_B3152_, new_B3151_,
    new_B3150_, new_B3149_, new_B3148_, new_B3147_, new_B3146_, new_B3139_,
    new_B3138_, new_B3137_, new_B3136_, new_B3135_, new_B3134_, new_B3133_,
    new_B3132_, new_B3131_, new_B3130_, new_B3129_, new_B3128_, new_B3127_,
    new_B3126_, new_B3125_, new_B3124_, new_B3123_, new_B3122_, new_B3121_,
    new_B3120_, new_B3119_, new_B3118_, new_B3117_, new_B3116_, new_B3115_,
    new_B3114_, new_B3113_, new_B3112_, new_B3111_, new_B3110_, new_B3109_,
    new_B3108_, new_B3107_, new_B3106_, new_B3105_, new_B3104_, new_B3103_,
    new_B3102_, new_B3101_, new_B3100_, new_B3099_, new_B3098_, new_B3097_,
    new_B3096_, new_B3095_, new_B3094_, new_B3093_, new_B3092_, new_B3091_,
    new_B3090_, new_B3089_, new_B3088_, new_B3087_, new_B3086_, new_B3085_,
    new_B3084_, new_B3083_, new_B3082_, new_B3081_, new_B3080_, new_B3079_,
    new_B3072_, new_B3071_, new_B3070_, new_B3069_, new_B3068_, new_B3067_,
    new_B3066_, new_B3065_, new_B3064_, new_B3063_, new_B3062_, new_B3061_,
    new_B3060_, new_B3059_, new_B3058_, new_B3057_, new_B3056_, new_B3055_,
    new_B3054_, new_B3053_, new_B3052_, new_B3051_, new_B3050_, new_B3049_,
    new_B3048_, new_B3047_, new_B3046_, new_B3045_, new_B3044_, new_B3043_,
    new_B3042_, new_B3041_, new_B3040_, new_B3039_, new_B3038_, new_B3037_,
    new_B3036_, new_B3035_, new_B3034_, new_B3033_, new_B3032_, new_B3031_,
    new_B3030_, new_B3029_, new_B3028_, new_B3027_, new_B3026_, new_B3025_,
    new_B3024_, new_B3023_, new_B3022_, new_B3021_, new_B3020_, new_B3019_,
    new_B3018_, new_B3017_, new_B3016_, new_B3015_, new_B3014_, new_B3013_,
    new_B3012_, new_B3005_, new_B3004_, new_B3003_, new_B3002_, new_B3001_,
    new_B3000_, new_B2999_, new_B2998_, new_B2997_, new_B2996_, new_B2995_,
    new_B2994_, new_B2993_, new_B2992_, new_B2991_, new_B2990_, new_B2989_,
    new_B2988_, new_B2987_, new_B2986_, new_B2985_, new_B2984_, new_B2983_,
    new_B2982_, new_B2981_, new_B2980_, new_B2979_, new_B2978_, new_B2977_,
    new_B2976_, new_B2975_, new_B2974_, new_B2973_, new_B2972_, new_B2971_,
    new_B2970_, new_B2969_, new_B2968_, new_B2967_, new_B2966_, new_B2965_,
    new_B2964_, new_B2963_, new_B2962_, new_B2961_, new_B2960_, new_B2959_,
    new_B2958_, new_B2957_, new_B2956_, new_B2955_, new_B2954_, new_B2953_,
    new_B2952_, new_B2951_, new_B2950_, new_B2949_, new_B2948_, new_B2947_,
    new_B2946_, new_B2945_, new_B2938_, new_B2937_, new_B2936_, new_B2935_,
    new_B2934_, new_B2933_, new_B2932_, new_B2931_, new_B2930_, new_B2929_,
    new_B2928_, new_B2927_, new_B2926_, new_B2925_, new_B2924_, new_B2923_,
    new_B2922_, new_B2921_, new_B2920_, new_B2919_, new_B2918_, new_B2917_,
    new_B2916_, new_B2915_, new_B2914_, new_B2913_, new_B2912_, new_B2911_,
    new_B2910_, new_B2909_, new_B2908_, new_B2907_, new_B2906_, new_B2905_,
    new_B2904_, new_B2903_, new_B2902_, new_B2901_, new_B2900_, new_B2899_,
    new_B2898_, new_B2897_, new_B2896_, new_B2895_, new_B2894_, new_B2893_,
    new_B2892_, new_B2891_, new_B2890_, new_B2889_, new_B2888_, new_B2887_,
    new_B2886_, new_B2885_, new_B2884_, new_B2883_, new_B2882_, new_B2881_,
    new_B2880_, new_B2879_, new_B2878_, new_B2871_, new_B2870_, new_B2869_,
    new_B2868_, new_B2867_, new_B2866_, new_B2865_, new_B2864_, new_B2863_,
    new_B2862_, new_B2861_, new_B2860_, new_B2859_, new_B2858_, new_B2857_,
    new_B2856_, new_B2855_, new_B2854_, new_B2853_, new_B2852_, new_B2851_,
    new_B2850_, new_B2849_, new_B2848_, new_B2847_, new_B2846_, new_B2845_,
    new_B2844_, new_B2843_, new_B2842_, new_B2841_, new_B2840_, new_B2839_,
    new_B2838_, new_B2837_, new_B2836_, new_B2835_, new_B2834_, new_B2833_,
    new_B2832_, new_B2831_, new_B2830_, new_B2829_, new_B2828_, new_B2827_,
    new_B2826_, new_B2825_, new_B2824_, new_B2823_, new_B2822_, new_B2821_,
    new_B2820_, new_B2819_, new_B2818_, new_B2817_, new_B2816_, new_B2815_,
    new_B2814_, new_B2813_, new_B2812_, new_B2811_, new_B2804_, new_B2803_,
    new_B2802_, new_B2801_, new_B2800_, new_B2799_, new_B2798_, new_B2797_,
    new_B2796_, new_B2795_, new_B2794_, new_B2793_, new_B2792_, new_B2791_,
    new_B2790_, new_B2789_, new_B2788_, new_B2787_, new_B2786_, new_B2785_,
    new_B2784_, new_B2783_, new_B2782_, new_B2781_, new_B2780_, new_B2779_,
    new_B2778_, new_B2777_, new_B2776_, new_B2775_, new_B2774_, new_B2773_,
    new_B2772_, new_B2771_, new_B2770_, new_B2769_, new_B2768_, new_B2767_,
    new_B2766_, new_B2765_, new_B2764_, new_B2763_, new_B2762_, new_B2761_,
    new_B2760_, new_B2759_, new_B2758_, new_B2757_, new_B2756_, new_B2755_,
    new_B2754_, new_B2753_, new_B2752_, new_B2751_, new_B2750_, new_B2749_,
    new_B2748_, new_B2747_, new_B2746_, new_B2745_, new_B2744_, new_B2737_,
    new_B2736_, new_B2735_, new_B2734_, new_B2733_, new_B2732_, new_B2731_,
    new_B2730_, new_B2729_, new_B2728_, new_B2727_, new_B2726_, new_B2725_,
    new_B2724_, new_B2723_, new_B2722_, new_B2721_, new_B2720_, new_B2719_,
    new_B2718_, new_B2717_, new_B2716_, new_B2715_, new_B2714_, new_B2713_,
    new_B2712_, new_B2711_, new_B2710_, new_B2709_, new_B2708_, new_B2707_,
    new_B2706_, new_B2705_, new_B2704_, new_B2703_, new_B2702_, new_B2701_,
    new_B2700_, new_B2699_, new_B2698_, new_B2697_, new_B2696_, new_B2695_,
    new_B2694_, new_B2693_, new_B2692_, new_B2691_, new_B2690_, new_B2689_,
    new_B2688_, new_B2687_, new_B2686_, new_B2685_, new_B2684_, new_B2683_,
    new_B2682_, new_B2681_, new_B2680_, new_B2679_, new_B2678_, new_B2677_,
    new_B2670_, new_B2669_, new_B2668_, new_B2667_, new_B2666_, new_B2665_,
    new_B2664_, new_B2663_, new_B2662_, new_B2661_, new_B2660_, new_B2659_,
    new_B2658_, new_B2657_, new_B2656_, new_B2655_, new_B2654_, new_B2653_,
    new_B2652_, new_B2651_, new_B2650_, new_B2649_, new_B2648_, new_B2647_,
    new_B2646_, new_B2645_, new_B2644_, new_B2643_, new_B2642_, new_B2641_,
    new_B2640_, new_B2639_, new_B2638_, new_B2637_, new_B2636_, new_B2635_,
    new_B2634_, new_B2633_, new_B2632_, new_B2631_, new_B2630_, new_B2629_,
    new_B2628_, new_B2627_, new_B2626_, new_B2625_, new_B2624_, new_B2623_,
    new_B2622_, new_B2621_, new_B2620_, new_B2619_, new_B2618_, new_B2617_,
    new_B2616_, new_B2615_, new_B2614_, new_B2613_, new_B2612_, new_B2611_,
    new_B2610_, new_B2603_, new_B2602_, new_B2601_, new_B2600_, new_B2599_,
    new_B2598_, new_B2597_, new_B2596_, new_B2595_, new_B2594_, new_B2593_,
    new_B2592_, new_B2591_, new_B2590_, new_B2589_, new_B2588_, new_B2587_,
    new_B2586_, new_B2585_, new_B2584_, new_B2583_, new_B2582_, new_B2581_,
    new_B2580_, new_B2579_, new_B2578_, new_B2577_, new_B2576_, new_B2575_,
    new_B2574_, new_B2573_, new_B2572_, new_B2571_, new_B2570_, new_B2569_,
    new_B2568_, new_B2567_, new_B2566_, new_B2565_, new_B2564_, new_B2563_,
    new_B2562_, new_B2561_, new_B2560_, new_B2559_, new_B2558_, new_B2557_,
    new_B2556_, new_B2555_, new_B2554_, new_B2553_, new_B2552_, new_B2551_,
    new_B2550_, new_B2549_, new_B2548_, new_B2547_, new_B2546_, new_B2545_,
    new_B2544_, new_B2543_, new_B2536_, new_B2535_, new_B2534_, new_B2533_,
    new_B2532_, new_B2531_, new_B2530_, new_B2529_, new_B2528_, new_B2527_,
    new_B2526_, new_B2525_, new_B2524_, new_B2523_, new_B2522_, new_B2521_,
    new_B2520_, new_B2519_, new_B2518_, new_B2517_, new_B2516_, new_B2515_,
    new_B2514_, new_B2513_, new_B2512_, new_B2511_, new_B2510_, new_B2509_,
    new_B2508_, new_B2507_, new_B2506_, new_B2505_, new_B2504_, new_B2503_,
    new_B2502_, new_B2501_, new_B2500_, new_B2499_, new_B2498_, new_B2497_,
    new_B2496_, new_B2495_, new_B2494_, new_B2493_, new_B2492_, new_B2491_,
    new_B2490_, new_B2489_, new_B2488_, new_B2487_, new_B2486_, new_B2485_,
    new_B2484_, new_B2483_, new_B2482_, new_B2481_, new_B2480_, new_B2479_,
    new_B2478_, new_B2477_, new_B2476_, new_B2469_, new_B2468_, new_B2467_,
    new_B2466_, new_B2465_, new_B2464_, new_B2463_, new_B2462_, new_B2461_,
    new_B2460_, new_B2459_, new_B2458_, new_B2457_, new_B2456_, new_B2455_,
    new_B2454_, new_B2453_, new_B2452_, new_B2451_, new_B2450_, new_B2449_,
    new_B2448_, new_B2447_, new_B2446_, new_B2445_, new_B2444_, new_B2443_,
    new_B2442_, new_B2441_, new_B2440_, new_B2439_, new_B2438_, new_B2437_,
    new_B2436_, new_B2435_, new_B2434_, new_B2433_, new_B2432_, new_B2431_,
    new_B2430_, new_B2429_, new_B2428_, new_B2427_, new_B2426_, new_B2425_,
    new_B2424_, new_B2423_, new_B2422_, new_B2421_, new_B2420_, new_B2419_,
    new_B2418_, new_B2417_, new_B2416_, new_B2415_, new_B2414_, new_B2413_,
    new_B2412_, new_B2411_, new_B2410_, new_B2409_, new_B2402_, new_B2401_,
    new_B2400_, new_B2399_, new_B2398_, new_B2397_, new_B2396_, new_B2395_,
    new_B2394_, new_B2393_, new_B2392_, new_B2391_, new_B2390_, new_B2389_,
    new_B2388_, new_B2387_, new_B2386_, new_B2385_, new_B2384_, new_B2383_,
    new_B2382_, new_B2381_, new_B2380_, new_B2379_, new_B2378_, new_B2377_,
    new_B2376_, new_B2375_, new_B2374_, new_B2373_, new_B2372_, new_B2371_,
    new_B2370_, new_B2369_, new_B2368_, new_B2367_, new_B2366_, new_B2365_,
    new_B2364_, new_B2363_, new_B2362_, new_B2361_, new_B2360_, new_B2359_,
    new_B2358_, new_B2357_, new_B2356_, new_B2355_, new_B2354_, new_B2353_,
    new_B2352_, new_B2351_, new_B2350_, new_B2349_, new_B2348_, new_B2347_,
    new_B2346_, new_B2345_, new_B2344_, new_B2343_, new_B2342_, new_B2335_,
    new_B2334_, new_B2333_, new_B2332_, new_B2331_, new_B2330_, new_B2329_,
    new_B2328_, new_B2327_, new_B2326_, new_B2325_, new_B2324_, new_B2323_,
    new_B2322_, new_B2321_, new_B2320_, new_B2319_, new_B2318_, new_B2317_,
    new_B2316_, new_B2315_, new_B2314_, new_B2313_, new_B2312_, new_B2311_,
    new_B2310_, new_B2309_, new_B2308_, new_B2307_, new_B2306_, new_B2305_,
    new_B2304_, new_B2303_, new_B2302_, new_B2301_, new_B2300_, new_B2299_,
    new_B2298_, new_B2297_, new_B2296_, new_B2295_, new_B2294_, new_B2293_,
    new_B2292_, new_B2291_, new_B2290_, new_B2289_, new_B2288_, new_B2287_,
    new_B2286_, new_B2285_, new_B2284_, new_B2283_, new_B2282_, new_B2281_,
    new_B2280_, new_B2279_, new_B2278_, new_B2277_, new_B2276_, new_B2275_,
    new_B2268_, new_B2267_, new_B2266_, new_B2265_, new_B2264_, new_B2263_,
    new_B2262_, new_B2261_, new_B2260_, new_B2259_, new_B2258_, new_B2257_,
    new_B2256_, new_B2255_, new_B2254_, new_B2253_, new_B2252_, new_B2251_,
    new_B2250_, new_B2249_, new_B2248_, new_B2247_, new_B2246_, new_B2245_,
    new_B2244_, new_B2243_, new_B2242_, new_B2241_, new_B2240_, new_B2239_,
    new_B2238_, new_B2237_, new_B2236_, new_B2235_, new_B2234_, new_B2233_,
    new_B2232_, new_B2231_, new_B2230_, new_B2229_, new_B2228_, new_B2227_,
    new_B2226_, new_B2225_, new_B2224_, new_B2223_, new_B2222_, new_B2221_,
    new_B2220_, new_B2219_, new_B2218_, new_B2217_, new_B2216_, new_B2215_,
    new_B2214_, new_B2213_, new_B2212_, new_B2211_, new_B2210_, new_B2209_,
    new_B2208_, new_B2201_, new_B2200_, new_B2199_, new_B2198_, new_B2197_,
    new_B2196_, new_B2195_, new_B2194_, new_B2193_, new_B2192_, new_B2191_,
    new_B2190_, new_B2189_, new_B2188_, new_B2187_, new_B2186_, new_B2185_,
    new_B2184_, new_B2183_, new_B2182_, new_B2181_, new_B2180_, new_B2179_,
    new_B2178_, new_B2177_, new_B2176_, new_B2175_, new_B2174_, new_B2173_,
    new_B2172_, new_B2171_, new_B2170_, new_B2169_, new_B2168_, new_B2167_,
    new_B2166_, new_B2165_, new_B2164_, new_B2163_, new_B2162_, new_B2161_,
    new_B2160_, new_B2159_, new_B2158_, new_B2157_, new_B2156_, new_B2155_,
    new_B2154_, new_B2153_, new_B2152_, new_B2151_, new_B2150_, new_B2149_,
    new_B2148_, new_B2147_, new_B2146_, new_B2145_, new_B2144_, new_B2143_,
    new_B2142_, new_B2141_, new_B2134_, new_B2133_, new_B2132_, new_B2131_,
    new_B2130_, new_B2129_, new_B2128_, new_B2127_, new_B2126_, new_B2125_,
    new_B2124_, new_B2123_, new_B2122_, new_B2121_, new_B2120_, new_B2119_,
    new_B2118_, new_B2117_, new_B2116_, new_B2115_, new_B2114_, new_B2113_,
    new_B2112_, new_B2111_, new_B2110_, new_B2109_, new_B2108_, new_B2107_,
    new_B2106_, new_B2105_, new_B2104_, new_B2103_, new_B2102_, new_B2101_,
    new_B2100_, new_B2099_, new_B2098_, new_B2097_, new_B2096_, new_B2095_,
    new_B2094_, new_B2093_, new_B2092_, new_B2091_, new_B2090_, new_B2089_,
    new_B2088_, new_B2087_, new_B2086_, new_B2085_, new_B2084_, new_B2083_,
    new_B2082_, new_B2081_, new_B2080_, new_B2079_, new_B2078_, new_B2077_,
    new_B2076_, new_B2075_, new_B2074_, new_B2067_, new_B2066_, new_B2065_,
    new_B2064_, new_B2063_, new_B2062_, new_B2061_, new_B2060_, new_B2059_,
    new_B2058_, new_B2057_, new_B2056_, new_B2055_, new_B2054_, new_B2053_,
    new_B2052_, new_B2051_, new_B2050_, new_B2049_, new_B2048_, new_B2047_,
    new_B2046_, new_B2045_, new_B2044_, new_B2043_, new_B2042_, new_B2041_,
    new_B2040_, new_B2039_, new_B2038_, new_B2037_, new_B2036_, new_B2035_,
    new_B2034_, new_B2033_, new_B2032_, new_B2031_, new_B2030_, new_B2029_,
    new_B2028_, new_B2027_, new_B2026_, new_B2025_, new_B2024_, new_B2023_,
    new_B2022_, new_B2021_, new_B2020_, new_B2019_, new_B2018_, new_B2017_,
    new_B2016_, new_B2015_, new_B2014_, new_B2013_, new_B2012_, new_B2011_,
    new_B2010_, new_B2009_, new_B2008_, new_B2007_, new_B2000_, new_B1999_,
    new_B1998_, new_B1997_, new_B1996_, new_B1995_, new_B1994_, new_B1993_,
    new_B1992_, new_B1991_, new_B1990_, new_B1989_, new_B1988_, new_B1987_,
    new_B1986_, new_B1985_, new_B1984_, new_B1983_, new_B1982_, new_B1981_,
    new_B1980_, new_B1979_, new_B1978_, new_B1977_, new_B1976_, new_B1975_,
    new_B1974_, new_B1973_, new_B1972_, new_B1971_, new_B1970_, new_B1969_,
    new_B1968_, new_B1967_, new_B1966_, new_B1965_, new_B1964_, new_B1963_,
    new_B1962_, new_B1961_, new_B1960_, new_B1959_, new_B1958_, new_B1957_,
    new_B1956_, new_B1955_, new_B1954_, new_B1953_, new_B1952_, new_B1951_,
    new_B1950_, new_B1949_, new_B1948_, new_B1947_, new_B1946_, new_B1945_,
    new_B1944_, new_B1943_, new_B1942_, new_B1941_, new_B1940_, new_B1933_,
    new_B1932_, new_B1931_, new_B1930_, new_B1929_, new_B1928_, new_B1927_,
    new_B1926_, new_B1925_, new_B1924_, new_B1923_, new_B1922_, new_B1921_,
    new_B1920_, new_B1919_, new_B1918_, new_B1917_, new_B1916_, new_B1915_,
    new_B1914_, new_B1913_, new_B1912_, new_B1911_, new_B1910_, new_B1909_,
    new_B1908_, new_B1907_, new_B1906_, new_B1905_, new_B1904_, new_B1903_,
    new_B1902_, new_B1901_, new_B1900_, new_B1899_, new_B1898_, new_B1897_,
    new_B1896_, new_B1895_, new_B1894_, new_B1893_, new_B1892_, new_B1891_,
    new_B1890_, new_B1889_, new_B1888_, new_B1887_, new_B1886_, new_B1885_,
    new_B1884_, new_B1883_, new_B1882_, new_B1881_, new_B1880_, new_B1879_,
    new_B1878_, new_B1877_, new_B1876_, new_B1875_, new_B1874_, new_B1873_,
    new_B1866_, new_B1865_, new_B1864_, new_B1863_, new_B1862_, new_B1861_,
    new_B1860_, new_B1859_, new_B1858_, new_B1857_, new_B1856_, new_B1855_,
    new_B1854_, new_B1853_, new_B1852_, new_B1851_, new_B1850_, new_B1849_,
    new_B1848_, new_B1847_, new_B1846_, new_B1845_, new_B1844_, new_B1843_,
    new_B1842_, new_B1841_, new_B1840_, new_B1839_, new_B1838_, new_B1837_,
    new_B1836_, new_B1835_, new_B1834_, new_B1833_, new_B1832_, new_B1831_,
    new_B1830_, new_B1829_, new_B1828_, new_B1827_, new_B1826_, new_B1825_,
    new_B1824_, new_B1823_, new_B1822_, new_B1821_, new_B1820_, new_B1819_,
    new_B1818_, new_B1817_, new_B1816_, new_B1815_, new_B1814_, new_B1813_,
    new_B1812_, new_B1811_, new_B1810_, new_B1809_, new_B1808_, new_B1807_,
    new_B1806_, new_B1799_, new_B1798_, new_B1797_, new_B1796_, new_B1795_,
    new_B1794_, new_B1793_, new_B1792_, new_B1791_, new_B1790_, new_B1789_,
    new_B1788_, new_B1787_, new_B1786_, new_B1785_, new_B1784_, new_B1783_,
    new_B1782_, new_B1781_, new_B1780_, new_B1779_, new_B1778_, new_B1777_,
    new_B1776_, new_B1775_, new_B1774_, new_B1773_, new_B1772_, new_B1771_,
    new_B1770_, new_B1769_, new_B1768_, new_B1767_, new_B1766_, new_B1765_,
    new_B1764_, new_B1763_, new_B1762_, new_B1761_, new_B1760_, new_B1759_,
    new_B1758_, new_B1757_, new_B1756_, new_B1755_, new_B1754_, new_B1753_,
    new_B1752_, new_B1751_, new_B1750_, new_B1749_, new_B1748_, new_B1747_,
    new_B1746_, new_B1745_, new_B1744_, new_B1743_, new_B1742_, new_B1741_,
    new_B1740_, new_B1739_, new_B1732_, new_B1731_, new_B1730_, new_B1729_,
    new_B1728_, new_B1727_, new_B1726_, new_B1725_, new_B1724_, new_B1723_,
    new_B1722_, new_B1721_, new_B1720_, new_B1719_, new_B1718_, new_B1717_,
    new_B1716_, new_B1715_, new_B1714_, new_B1713_, new_B1712_, new_B1711_,
    new_B1710_, new_B1709_, new_B1708_, new_B1707_, new_B1706_, new_B1705_,
    new_B1704_, new_B1703_, new_B1702_, new_B1701_, new_B1700_, new_B1699_,
    new_B1698_, new_B1697_, new_B1696_, new_B1695_, new_B1694_, new_B1693_,
    new_B1692_, new_B1691_, new_B1690_, new_B1689_, new_B1688_, new_B1687_,
    new_B1686_, new_B1685_, new_B1684_, new_B1683_, new_B1682_, new_B1681_,
    new_B1680_, new_B1679_, new_B1678_, new_B1677_, new_B1676_, new_B1675_,
    new_B1674_, new_B1673_, new_B1672_, new_B1665_, new_B1664_, new_B1663_,
    new_B1662_, new_B1661_, new_B1660_, new_B1659_, new_B1658_, new_B1657_,
    new_B1656_, new_B1655_, new_B1654_, new_B1653_, new_B1652_, new_B1651_,
    new_B1650_, new_B1649_, new_B1648_, new_B1647_, new_B1646_, new_B1645_,
    new_B1644_, new_B1643_, new_B1642_, new_B1641_, new_B1640_, new_B1639_,
    new_B1638_, new_B1637_, new_B1636_, new_B1635_, new_B1634_, new_B1633_,
    new_B1632_, new_B1631_, new_B1630_, new_B1629_, new_B1628_, new_B1627_,
    new_B1626_, new_B1625_, new_B1624_, new_B1623_, new_B1622_, new_B1621_,
    new_B1620_, new_B1619_, new_B1618_, new_B1617_, new_B1616_, new_B1615_,
    new_B1614_, new_B1613_, new_B1612_, new_B1611_, new_B1610_, new_B1609_,
    new_B1608_, new_B1607_, new_B1606_, new_B1605_, new_B1598_, new_B1597_,
    new_B1596_, new_B1595_, new_B1594_, new_B1593_, new_B1592_, new_B1591_,
    new_B1590_, new_B1589_, new_B1588_, new_B1587_, new_B1586_, new_B1585_,
    new_B1584_, new_B1583_, new_B1582_, new_B1581_, new_B1580_, new_B1579_,
    new_B1578_, new_B1577_, new_B1576_, new_B1575_, new_B1574_, new_B1573_,
    new_B1572_, new_B1571_, new_B1570_, new_B1569_, new_B1568_, new_B1567_,
    new_B1566_, new_B1565_, new_B1564_, new_B1563_, new_B1562_, new_B1561_,
    new_B1560_, new_B1559_, new_B1558_, new_B1557_, new_B1556_, new_B1555_,
    new_B1554_, new_B1553_, new_B1552_, new_B1551_, new_B1550_, new_B1549_,
    new_B1548_, new_B1547_, new_B1546_, new_B1545_, new_B1544_, new_B1543_,
    new_B1542_, new_B1541_, new_B1540_, new_B1539_, new_B1538_, new_B1531_,
    new_B1530_, new_B1529_, new_B1528_, new_B1527_, new_B1526_, new_B1525_,
    new_B1524_, new_B1523_, new_B1522_, new_B1521_, new_B1520_, new_B1519_,
    new_B1518_, new_B1517_, new_B1516_, new_B1515_, new_B1514_, new_B1513_,
    new_B1512_, new_B1511_, new_B1510_, new_B1509_, new_B1508_, new_B1507_,
    new_B1506_, new_B1505_, new_B1504_, new_B1503_, new_B1502_, new_B1501_,
    new_B1500_, new_B1499_, new_B1498_, new_B1497_, new_B1496_, new_B1495_,
    new_B1494_, new_B1493_, new_B1492_, new_B1491_, new_B1490_, new_B1489_,
    new_B1488_, new_B1487_, new_B1486_, new_B1485_, new_B1484_, new_B1483_,
    new_B1482_, new_B1481_, new_B1480_, new_B1479_, new_B1478_, new_B1477_,
    new_B1476_, new_B1475_, new_B1474_, new_B1473_, new_B1472_, new_B1471_,
    new_B1464_, new_B1463_, new_B1462_, new_B1461_, new_B1460_, new_B1459_,
    new_B1458_, new_B1457_, new_B1456_, new_B1455_, new_B1454_, new_B1453_,
    new_B1452_, new_B1451_, new_B1450_, new_B1449_, new_B1448_, new_B1447_,
    new_B1446_, new_B1445_, new_B1444_, new_B1443_, new_B1442_, new_B1441_,
    new_B1440_, new_B1439_, new_B1438_, new_B1437_, new_B1436_, new_B1435_,
    new_B1434_, new_B1433_, new_B1432_, new_B1431_, new_B1430_, new_B1429_,
    new_B1428_, new_B1427_, new_B1426_, new_B1425_, new_B1424_, new_B1423_,
    new_B1422_, new_B1421_, new_B1420_, new_B1419_, new_B1418_, new_B1417_,
    new_B1416_, new_B1415_, new_B1414_, new_B1413_, new_B1412_, new_B1411_,
    new_B1410_, new_B1409_, new_B1408_, new_B1407_, new_B1406_, new_B1405_,
    new_B1404_, new_B1397_, new_B1396_, new_B1395_, new_B1394_, new_B1393_,
    new_B1392_, new_B1391_, new_B1390_, new_B1389_, new_B1388_, new_B1387_,
    new_B1386_, new_B1385_, new_B1384_, new_B1383_, new_B1382_, new_B1381_,
    new_B1380_, new_B1379_, new_B1378_, new_B1377_, new_B1376_, new_B1375_,
    new_B1374_, new_B1373_, new_B1372_, new_B1371_, new_B1370_, new_B1369_,
    new_B1368_, new_B1367_, new_B1366_, new_B1365_, new_B1364_, new_B1363_,
    new_B1362_, new_B1361_, new_B1360_, new_B1359_, new_B1358_, new_B1357_,
    new_B1356_, new_B1355_, new_B1354_, new_B1353_, new_B1352_, new_B1351_,
    new_B1350_, new_B1349_, new_B1348_, new_B1347_, new_B1346_, new_B1345_,
    new_B1344_, new_B1343_, new_B1342_, new_B1341_, new_B1340_, new_B1339_,
    new_B1338_, new_B1337_, new_B1330_, new_B1329_, new_B1328_, new_B1327_,
    new_B1326_, new_B1325_, new_B1324_, new_B1323_, new_B1322_, new_B1321_,
    new_B1320_, new_B1319_, new_B1318_, new_B1317_, new_B1316_, new_B1315_,
    new_B1314_, new_B1313_, new_B1312_, new_B1311_, new_B1310_, new_B1309_,
    new_B1308_, new_B1307_, new_B1306_, new_B1305_, new_B1304_, new_B1303_,
    new_B1302_, new_B1301_, new_B1300_, new_B1299_, new_B1298_, new_B1297_,
    new_B1296_, new_B1295_, new_B1294_, new_B1293_, new_B1292_, new_B1291_,
    new_B1290_, new_B1289_, new_B1288_, new_B1287_, new_B1286_, new_B1285_,
    new_B1284_, new_B1283_, new_B1282_, new_B1281_, new_B1280_, new_B1279_,
    new_B1278_, new_B1277_, new_B1276_, new_B1275_, new_B1274_, new_B1273_,
    new_B1272_, new_B1271_, new_B1270_, new_B1263_, new_B1262_, new_B1261_,
    new_B1260_, new_B1259_, new_B1258_, new_B1257_, new_B1256_, new_B1255_,
    new_B1254_, new_B1253_, new_B1252_, new_B1251_, new_B1250_, new_B1249_,
    new_B1248_, new_B1247_, new_B1246_, new_B1245_, new_B1244_, new_B1243_,
    new_B1242_, new_B1241_, new_B1240_, new_B1239_, new_B1238_, new_B1237_,
    new_B1236_, new_B1235_, new_B1234_, new_B1233_, new_B1232_, new_B1231_,
    new_B1230_, new_B1229_, new_B1228_, new_B1227_, new_B1226_, new_B1225_,
    new_B1224_, new_B1223_, new_B1222_, new_B1221_, new_B1220_, new_B1219_,
    new_B1218_, new_B1217_, new_B1216_, new_B1215_, new_B1214_, new_B1213_,
    new_B1212_, new_B1211_, new_B1210_, new_B1209_, new_B1208_, new_B1207_,
    new_B1206_, new_B1205_, new_B1204_, new_B1203_, new_B1196_, new_B1195_,
    new_B1194_, new_B1193_, new_B1192_, new_B1191_, new_B1190_, new_B1189_,
    new_B1188_, new_B1187_, new_B1186_, new_B1185_, new_B1184_, new_B1183_,
    new_B1182_, new_B1181_, new_B1180_, new_B1179_, new_B1178_, new_B1177_,
    new_B1176_, new_B1175_, new_B1174_, new_B1173_, new_B1172_, new_B1171_,
    new_B1170_, new_B1169_, new_B1168_, new_B1167_, new_B1166_, new_B1165_,
    new_B1164_, new_B1163_, new_B1162_, new_B1161_, new_B1160_, new_B1159_,
    new_B1158_, new_B1157_, new_B1156_, new_B1155_, new_B1154_, new_B1153_,
    new_B1152_, new_B1151_, new_B1150_, new_B1149_, new_B1148_, new_B1147_,
    new_B1146_, new_B1145_, new_B1144_, new_B1143_, new_B1142_, new_B1141_,
    new_B1140_, new_B1139_, new_B1138_, new_B1137_, new_B1136_, new_B1129_,
    new_B1128_, new_B1127_, new_B1126_, new_B1125_, new_B1124_, new_B1123_,
    new_B1122_, new_B1121_, new_B1120_, new_B1119_, new_B1118_, new_B1117_,
    new_B1116_, new_B1115_, new_B1114_, new_B1113_, new_B1112_, new_B1111_,
    new_B1110_, new_B1109_, new_B1108_, new_B1107_, new_B1106_, new_B1105_,
    new_B1104_, new_B1103_, new_B1102_, new_B1101_, new_B1100_, new_B1099_,
    new_B1098_, new_B1097_, new_B1096_, new_B1095_, new_B1094_, new_B1093_,
    new_B1092_, new_B1091_, new_B1090_, new_B1089_, new_B1088_, new_B1087_,
    new_B1086_, new_B1085_, new_B1084_, new_B1083_, new_B1082_, new_B1081_,
    new_B1080_, new_B1079_, new_B1078_, new_B1077_, new_B1076_, new_B1075_,
    new_B1074_, new_B1073_, new_B1072_, new_B1071_, new_B1070_, new_B1069_,
    new_B1062_, new_B1061_, new_B1060_, new_B1059_, new_B1058_, new_B1057_,
    new_B1056_, new_B1055_, new_B1054_, new_B1053_, new_B1052_, new_B1051_,
    new_B1050_, new_B1049_, new_B1048_, new_B1047_, new_B1046_, new_B1045_,
    new_B1044_, new_B1043_, new_B1042_, new_B1041_, new_B1040_, new_B1039_,
    new_B1038_, new_B1037_, new_B1036_, new_B1035_, new_B1034_, new_B1033_,
    new_B1032_, new_B1031_, new_B1030_, new_B1029_, new_B1028_, new_B1027_,
    new_B1026_, new_B1025_, new_B1024_, new_B1023_, new_B1022_, new_B1021_,
    new_B1020_, new_B1019_, new_B1018_, new_B1017_, new_B1016_, new_B1015_,
    new_B1014_, new_B1013_, new_B1012_, new_B1011_, new_B1010_, new_B1009_,
    new_B1008_, new_B1007_, new_B1006_, new_B1005_, new_B1004_, new_B1003_,
    new_B1002_, new_B995_, new_B994_, new_B993_, new_B992_, new_B991_,
    new_B990_, new_B989_, new_B988_, new_B987_, new_B986_, new_B985_,
    new_B984_, new_B983_, new_B982_, new_B981_, new_B980_, new_B979_,
    new_B978_, new_B977_, new_B976_, new_B975_, new_B974_, new_B973_,
    new_B972_, new_B971_, new_B970_, new_B969_, new_B968_, new_B967_,
    new_B966_, new_B965_, new_B964_, new_B963_, new_B962_, new_B961_,
    new_B960_, new_B959_, new_B958_, new_B957_, new_B956_, new_B955_,
    new_B954_, new_B953_, new_B952_, new_B951_, new_B950_, new_B949_,
    new_B948_, new_B947_, new_B946_, new_B945_, new_B944_, new_B943_,
    new_B942_, new_B941_, new_B940_, new_B939_, new_B938_, new_B937_,
    new_B936_, new_B935_, new_B928_, new_B927_, new_B926_, new_B925_,
    new_B924_, new_B923_, new_B922_, new_B921_, new_B920_, new_B919_,
    new_B918_, new_B917_, new_B916_, new_B915_, new_B914_, new_B913_,
    new_B912_, new_B911_, new_B910_, new_B909_, new_B908_, new_B907_,
    new_B906_, new_B905_, new_B904_, new_B903_, new_B902_, new_B901_,
    new_B900_, new_B899_, new_B898_, new_B897_, new_B896_, new_B895_,
    new_B894_, new_B893_, new_B892_, new_B891_, new_B890_, new_B889_,
    new_B888_, new_B887_, new_B886_, new_B885_, new_B884_, new_B883_,
    new_B882_, new_B881_, new_B880_, new_B879_, new_B878_, new_B877_,
    new_B876_, new_B875_, new_B874_, new_B873_, new_B872_, new_B871_,
    new_B870_, new_B869_, new_B868_, new_B861_, new_B860_, new_B859_,
    new_B858_, new_B857_, new_B856_, new_B855_, new_B854_, new_B853_,
    new_B852_, new_B851_, new_B850_, new_B849_, new_B848_, new_B847_,
    new_B846_, new_B845_, new_B844_, new_B843_, new_B842_, new_B841_,
    new_B840_, new_B839_, new_B838_, new_B837_, new_B836_, new_B835_,
    new_B834_, new_B833_, new_B832_, new_B831_, new_B830_, new_B829_,
    new_B828_, new_B827_, new_B826_, new_B825_, new_B824_, new_B823_,
    new_B822_, new_B821_, new_B820_, new_B819_, new_B818_, new_B817_,
    new_B816_, new_B815_, new_B814_, new_B813_, new_B812_, new_B811_,
    new_B810_, new_B809_, new_B808_, new_B807_, new_B806_, new_B805_,
    new_B804_, new_B803_, new_B802_, new_B801_, new_B794_, new_B793_,
    new_B792_, new_B791_, new_B790_, new_B789_, new_B788_, new_B787_,
    new_B786_, new_B785_, new_B784_, new_B783_, new_B782_, new_B781_,
    new_B780_, new_B779_, new_B778_, new_B777_, new_B776_, new_B775_,
    new_B774_, new_B773_, new_B772_, new_B771_, new_B770_, new_B769_,
    new_B768_, new_B767_, new_B766_, new_B765_, new_B764_, new_B763_,
    new_B762_, new_B761_, new_B760_, new_B759_, new_B758_, new_B757_,
    new_B756_, new_B755_, new_B754_, new_B753_, new_B752_, new_B751_,
    new_B750_, new_B749_, new_B748_, new_B747_, new_B746_, new_B745_,
    new_B744_, new_B743_, new_B742_, new_B741_, new_B740_, new_B739_,
    new_B738_, new_B737_, new_B736_, new_B735_, new_B734_, new_B727_,
    new_B726_, new_B725_, new_B724_, new_B723_, new_B722_, new_B721_,
    new_B720_, new_B719_, new_B718_, new_B717_, new_B716_, new_B715_,
    new_B714_, new_B713_, new_B712_, new_B711_, new_B710_, new_B709_,
    new_B708_, new_B707_, new_B706_, new_B705_, new_B704_, new_B703_,
    new_B702_, new_B701_, new_B700_, new_B699_, new_B698_, new_B697_,
    new_B696_, new_B695_, new_B694_, new_B693_, new_B692_, new_B691_,
    new_B690_, new_B689_, new_B688_, new_B687_, new_B686_, new_B685_,
    new_B684_, new_B683_, new_B682_, new_B681_, new_B680_, new_B679_,
    new_B678_, new_B677_, new_B676_, new_B675_, new_B674_, new_B673_,
    new_B672_, new_B671_, new_B670_, new_B669_, new_B668_, new_B667_,
    new_B660_, new_B659_, new_B658_, new_B657_, new_B656_, new_B655_,
    new_B654_, new_B653_, new_B652_, new_B651_, new_B650_, new_B649_,
    new_B648_, new_B647_, new_B646_, new_B645_, new_B644_, new_B643_,
    new_B642_, new_B641_, new_B640_, new_B639_, new_B638_, new_B637_,
    new_B636_, new_B635_, new_B634_, new_B633_, new_B632_, new_B631_,
    new_B630_, new_B629_, new_B628_, new_B627_, new_B626_, new_B625_,
    new_B624_, new_B623_, new_B622_, new_B621_, new_B620_, new_B619_,
    new_B618_, new_B617_, new_B616_, new_B615_, new_B614_, new_B613_,
    new_B612_, new_B611_, new_B610_, new_B609_, new_B608_, new_B607_,
    new_B606_, new_B605_, new_B604_, new_B603_, new_B602_, new_B601_,
    new_B600_, new_B593_, new_B592_, new_B591_, new_B590_, new_B589_,
    new_B588_, new_B587_, new_B586_, new_B585_, new_B584_, new_B583_,
    new_B582_, new_B581_, new_B580_, new_B579_, new_B578_, new_B577_,
    new_B576_, new_B575_, new_B574_, new_B573_, new_B572_, new_B571_,
    new_B570_, new_B569_, new_B568_, new_B567_, new_B566_, new_B565_,
    new_B564_, new_B563_, new_B562_, new_B561_, new_B560_, new_B559_,
    new_B558_, new_B557_, new_B556_, new_B555_, new_B554_, new_B553_,
    new_B552_, new_B551_, new_B550_, new_B549_, new_B548_, new_B547_,
    new_B546_, new_B545_, new_B544_, new_B543_, new_B542_, new_B541_,
    new_B540_, new_B539_, new_B538_, new_B537_, new_B536_, new_B535_,
    new_B534_, new_B533_, new_B526_, new_B525_, new_B524_, new_B523_,
    new_B522_, new_B521_, new_B520_, new_B519_, new_B518_, new_B517_,
    new_B516_, new_B515_, new_B514_, new_B513_, new_B512_, new_B511_,
    new_B510_, new_B509_, new_B508_, new_B507_, new_B506_, new_B505_,
    new_B504_, new_B503_, new_B502_, new_B501_, new_B500_, new_B499_,
    new_B498_, new_B497_, new_B496_, new_B495_, new_B494_, new_B493_,
    new_B492_, new_B491_, new_B490_, new_B489_, new_B488_, new_B487_,
    new_B486_, new_B485_, new_B484_, new_B483_, new_B482_, new_B481_,
    new_B480_, new_B479_, new_B478_, new_B477_, new_B476_, new_B475_,
    new_B474_, new_B473_, new_B472_, new_B471_, new_B470_, new_B469_,
    new_B468_, new_B467_, new_B466_, new_B459_, new_B458_, new_B457_,
    new_B456_, new_B455_, new_B454_, new_B453_, new_B452_, new_B451_,
    new_B450_, new_B449_, new_B448_, new_B447_, new_B446_, new_B445_,
    new_B444_, new_B443_, new_B442_, new_B441_, new_B440_, new_B439_,
    new_B438_, new_B437_, new_B436_, new_B435_, new_B434_, new_B433_,
    new_B432_, new_B431_, new_B430_, new_B429_, new_B428_, new_B427_,
    new_B426_, new_B425_, new_B424_, new_B423_, new_B422_, new_B421_,
    new_B420_, new_B419_, new_B418_, new_B417_, new_B416_, new_B415_,
    new_B414_, new_B413_, new_B412_, new_B411_, new_B410_, new_B409_,
    new_B408_, new_B407_, new_B406_, new_B405_, new_B404_, new_B403_,
    new_B402_, new_B401_, new_B400_, new_B399_, new_B392_, new_B391_,
    new_B390_, new_B389_, new_B388_, new_B387_, new_B386_, new_B385_,
    new_B384_, new_B383_, new_B382_, new_B381_, new_B380_, new_B379_,
    new_B378_, new_B377_, new_B376_, new_B375_, new_B374_, new_B373_,
    new_B372_, new_B371_, new_B370_, new_B369_, new_B368_, new_B367_,
    new_B366_, new_B365_, new_B364_, new_B363_, new_B362_, new_B361_,
    new_B360_, new_B359_, new_B358_, new_B357_, new_B356_, new_B355_,
    new_B354_, new_B353_, new_B352_, new_B351_, new_B350_, new_B349_,
    new_B348_, new_B347_, new_B346_, new_B345_, new_B344_, new_B343_,
    new_B342_, new_B341_, new_B340_, new_B339_, new_B338_, new_B337_,
    new_B336_, new_B335_, new_B334_, new_B333_, new_B332_, new_B325_,
    new_B324_, new_B323_, new_B322_, new_B321_, new_B320_, new_B319_,
    new_B318_, new_B317_, new_B316_, new_B315_, new_B314_, new_B313_,
    new_B312_, new_B311_, new_B310_, new_B309_, new_B308_, new_B307_,
    new_B306_, new_B305_, new_B304_, new_B303_, new_B302_, new_B301_,
    new_B300_, new_B299_, new_B298_, new_B297_, new_B296_, new_B295_,
    new_B294_, new_B293_, new_B292_, new_B291_, new_B290_, new_B289_,
    new_B288_, new_B287_, new_B286_, new_B285_, new_B284_, new_B283_,
    new_B282_, new_B281_, new_B280_, new_B279_, new_B278_, new_B277_,
    new_B276_, new_B275_, new_B274_, new_B273_, new_B272_, new_B271_,
    new_B270_, new_B269_, new_B268_, new_B267_, new_B266_, new_B265_,
    new_B258_, new_B257_, new_B256_, new_B255_, new_B254_, new_B253_,
    new_B252_, new_B251_, new_B250_, new_B249_, new_B248_, new_B247_,
    new_B246_, new_B245_, new_B244_, new_B243_, new_B242_, new_B241_,
    new_B240_, new_B239_, new_B238_, new_B237_, new_B236_, new_B235_,
    new_B234_, new_B233_, new_B232_, new_B231_, new_B230_, new_B229_,
    new_B228_, new_B227_, new_B226_, new_B225_, new_B224_, new_B223_,
    new_B222_, new_B221_, new_B220_, new_B219_, new_B218_, new_B217_,
    new_B216_, new_B215_, new_B214_, new_B213_, new_B212_, new_B211_,
    new_B210_, new_B209_, new_B208_, new_B207_, new_B206_, new_B205_,
    new_B204_, new_B203_, new_B202_, new_B201_, new_B200_, new_B199_,
    new_B198_, new_B191_, new_B190_, new_B189_, new_B188_, new_B187_,
    new_B186_, new_B185_, new_B184_, new_B183_, new_B182_, new_B181_,
    new_B180_, new_B179_, new_B178_, new_B177_, new_B176_, new_B175_,
    new_B174_, new_B173_, new_B172_, new_B171_, new_B170_, new_B169_,
    new_B168_, new_B167_, new_B166_, new_B165_, new_B164_, new_B163_,
    new_B162_, new_B161_, new_B160_, new_B159_, new_B158_, new_B157_,
    new_B156_, new_B155_, new_B154_, new_B153_, new_B152_, new_B151_,
    new_B150_, new_B149_, new_B148_, new_B147_, new_B146_, new_B145_,
    new_B144_, new_B143_, new_B142_, new_B141_, new_B140_, new_B139_,
    new_B138_, new_B137_, new_B136_, new_B135_, new_B134_, new_B133_,
    new_B132_, new_B131_, new_B124_, new_B123_, new_B122_, new_B121_,
    new_B120_, new_B119_, new_B118_, new_B117_, new_B116_, new_B115_,
    new_B114_, new_B113_, new_B112_, new_B111_, new_B110_, new_B109_,
    new_B108_, new_B107_, new_B106_, new_B105_, new_B104_, new_B103_,
    new_B102_, new_B101_, new_B100_, new_B99_, new_B98_, new_B97_,
    new_B96_, new_B95_, new_B94_, new_B93_, new_B92_, new_B91_, new_B90_,
    new_B89_, new_B88_, new_B87_, new_B86_, new_B85_, new_B84_, new_B83_,
    new_B82_, new_B81_, new_B80_, new_B79_, new_B78_, new_B77_, new_B76_,
    new_B75_, new_B74_, new_B73_, new_B72_, new_B71_, new_B70_, new_B69_,
    new_B68_, new_B67_, new_B66_, new_B65_, new_B64_, new_B57_, new_B56_,
    new_B55_, new_B54_, new_B53_, new_B52_, new_B51_, new_B50_, new_B49_,
    new_B48_, new_B47_, new_B46_, new_B45_, new_B44_, new_B43_, new_B42_,
    new_B41_, new_B40_, new_B39_, new_B38_, new_B37_, new_B36_, new_B35_,
    new_B34_, new_B33_, new_B32_, new_B31_, new_B30_, new_B29_, new_B28_,
    new_B27_, new_B26_, new_B25_, new_B24_, new_B23_, new_B22_, new_B21_,
    new_B20_, new_B19_, new_B18_, new_B17_, new_B16_, new_B15_, new_B14_,
    new_B13_, new_B12_, new_B11_, new_B10_, new_B9_, new_B8_, new_B7_,
    new_B6_, new_B5_, new_B4_, new_B3_, new_B2_, new_B1_, new_A9999_,
    new_A9998_, new_A9997_, new_A9996_, new_A9989_, new_A9988_, new_A9987_,
    new_A9986_, new_A9985_, new_A9984_, new_A9983_, new_A9982_, new_A9981_,
    new_A9980_, new_A9979_, new_A9978_, new_A9977_, new_A9976_, new_A9975_,
    new_A9974_, new_A9973_, new_A9972_, new_A9971_, new_A9970_, new_A9969_,
    new_A9968_, new_A9967_, new_A9966_, new_A9965_, new_A9964_, new_A9963_,
    new_A9962_, new_A9961_, new_A9960_, new_A9959_, new_A9958_, new_A9957_,
    new_A9956_, new_A9955_, new_A9954_, new_A9953_, new_A9952_, new_A9951_,
    new_A9950_, new_A9949_, new_A9948_, new_A9947_, new_A9946_, new_A9945_,
    new_A9944_, new_A9943_, new_A9942_, new_A9941_, new_A9940_, new_A9939_,
    new_A9938_, new_A9937_, new_A9936_, new_A9935_, new_A9934_, new_A9933_,
    new_A9932_, new_A9931_, new_A9930_, new_A9929_, new_A9922_, new_A9921_,
    new_A9920_, new_A9919_, new_A9918_, new_A9917_, new_A9916_, new_A9915_,
    new_A9914_, new_A9913_, new_A9912_, new_A9911_, new_A9910_, new_A9909_,
    new_A9908_, new_A9907_, new_A9906_, new_A9905_, new_A9904_, new_A9903_,
    new_A9902_, new_A9901_, new_A9900_, new_A9899_, new_A9898_, new_A9897_,
    new_A9896_, new_A9895_, new_A9894_, new_A9893_, new_A9892_, new_A9891_,
    new_A9890_, new_A9889_, new_A9888_, new_A9887_, new_A9886_, new_A9885_,
    new_A9884_, new_A9883_, new_A9882_, new_A9881_, new_A9880_, new_A9879_,
    new_A9878_, new_A9877_, new_A9876_, new_A9875_, new_A9874_, new_A9873_,
    new_A9872_, new_A9871_, new_A9870_, new_A9869_, new_A9868_, new_A9867_,
    new_A9866_, new_A9865_, new_A9864_, new_A9863_, new_A9862_, new_A9855_,
    new_A9854_, new_A9853_, new_A9852_, new_A9851_, new_A9850_, new_A9849_,
    new_A9848_, new_A9847_, new_A9846_, new_A9845_, new_A9844_, new_A9843_,
    new_A9842_, new_A9841_, new_A9840_, new_A9839_, new_A9838_, new_A9837_,
    new_A9836_, new_A9835_, new_A9834_, new_A9833_, new_A9832_, new_A9831_,
    new_A9830_, new_A9829_, new_A9828_, new_A9827_, new_A9826_, new_A9825_,
    new_A9824_, new_A9823_, new_A9822_, new_A9821_, new_A9820_, new_A9819_,
    new_A9818_, new_A9817_, new_A9816_, new_A9815_, new_A9814_, new_A9813_,
    new_A9812_, new_A9811_, new_A9810_, new_A9809_, new_A9808_, new_A9807_,
    new_A9806_, new_A9805_, new_A9804_, new_A9803_, new_A9802_, new_A9801_,
    new_A9800_, new_A9799_, new_A9798_, new_A9797_, new_A9796_, new_A9795_,
    new_A9788_, new_A9787_, new_A9786_, new_A9785_, new_A9784_, new_A9783_,
    new_A9782_, new_A9781_, new_A9780_, new_A9779_, new_A9778_, new_A9777_,
    new_A9776_, new_A9775_, new_A9774_, new_A9773_, new_A9772_, new_A9771_,
    new_A9770_, new_A9769_, new_A9768_, new_A9767_, new_A9766_, new_A9765_,
    new_A9764_, new_A9763_, new_A9762_, new_A9761_, new_A9760_, new_A9759_,
    new_A9758_, new_A9757_, new_A9756_, new_A9755_, new_A9754_, new_A9753_,
    new_A9752_, new_A9751_, new_A9750_, new_A9749_, new_A9748_, new_A9747_,
    new_A9746_, new_A9745_, new_A9744_, new_A9743_, new_A9742_, new_A9741_,
    new_A9740_, new_A9739_, new_A9738_, new_A9737_, new_A9736_, new_A9735_,
    new_A9734_, new_A9733_, new_A9732_, new_A9731_, new_A9730_, new_A9729_,
    new_A9728_, new_A9721_, new_A9720_, new_A9719_, new_A9718_, new_A9717_,
    new_A9716_, new_A9715_, new_A9714_, new_A9713_, new_A9712_, new_A9711_,
    new_A9710_, new_A9709_, new_A9708_, new_A9707_, new_A9706_, new_A9705_,
    new_A9704_, new_A9703_, new_A9702_, new_A9701_, new_A9700_, new_A9699_,
    new_A9698_, new_A9697_, new_A9696_, new_A9695_, new_A9694_, new_A9693_,
    new_A9692_, new_A9691_, new_A9690_, new_A9689_, new_A9688_, new_A9687_,
    new_A9686_, new_A9685_, new_A9684_, new_A9683_, new_A9682_, new_A9681_,
    new_A9680_, new_A9679_, new_A9678_, new_A9677_, new_A9676_, new_A9675_,
    new_A9674_, new_A9673_, new_A9672_, new_A9671_, new_A9670_, new_A9669_,
    new_A9668_, new_A9667_, new_A9666_, new_A9665_, new_A9664_, new_A9663_,
    new_A9662_, new_A9661_, new_A9654_, new_A9653_, new_A9652_, new_A9651_,
    new_A9650_, new_A9649_, new_A9648_, new_A9647_, new_A9646_, new_A9645_,
    new_A9644_, new_A9643_, new_A9642_, new_A9641_, new_A9640_, new_A9639_,
    new_A9638_, new_A9637_, new_A9636_, new_A9635_, new_A9634_, new_A9633_,
    new_A9632_, new_A9631_, new_A9630_, new_A9629_, new_A9628_, new_A9627_,
    new_A9626_, new_A9625_, new_A9624_, new_A9623_, new_A9622_, new_A9621_,
    new_A9620_, new_A9619_, new_A9618_, new_A9617_, new_A9616_, new_A9615_,
    new_A9614_, new_A9613_, new_A9612_, new_A9611_, new_A9610_, new_A9609_,
    new_A9608_, new_A9607_, new_A9606_, new_A9605_, new_A9604_, new_A9603_,
    new_A9602_, new_A9601_, new_A9600_, new_A9599_, new_A9598_, new_A9597_,
    new_A9596_, new_A9595_, new_A9594_, new_A9587_, new_A9586_, new_A9585_,
    new_A9584_, new_A9583_, new_A9582_, new_A9581_, new_A9580_, new_A9579_,
    new_A9578_, new_A9577_, new_A9576_, new_A9575_, new_A9574_, new_A9573_,
    new_A9572_, new_A9571_, new_A9570_, new_A9569_, new_A9568_, new_A9567_,
    new_A9566_, new_A9565_, new_A9564_, new_A9563_, new_A9562_, new_A9561_,
    new_A9560_, new_A9559_, new_A9558_, new_A9557_, new_A9556_, new_A9555_,
    new_A9554_, new_A9553_, new_A9552_, new_A9551_, new_A9550_, new_A9549_,
    new_A9548_, new_A9547_, new_A9546_, new_A9545_, new_A9544_, new_A9543_,
    new_A9542_, new_A9541_, new_A9540_, new_A9539_, new_A9538_, new_A9537_,
    new_A9536_, new_A9535_, new_A9534_, new_A9533_, new_A9532_, new_A9531_,
    new_A9530_, new_A9529_, new_A9528_, new_A9527_, new_A9520_, new_A9519_,
    new_A9518_, new_A9517_, new_A9516_, new_A9515_, new_A9514_, new_A9513_,
    new_A9512_, new_A9511_, new_A9510_, new_A9509_, new_A9508_, new_A9507_,
    new_A9506_, new_A9505_, new_A9504_, new_A9503_, new_A9502_, new_A9501_,
    new_A9500_, new_A9499_, new_A9498_, new_A9497_, new_A9496_, new_A9495_,
    new_A9494_, new_A9493_, new_A9492_, new_A9491_, new_A9490_, new_A9489_,
    new_A9488_, new_A9487_, new_A9486_, new_A9485_, new_A9484_, new_A9483_,
    new_A9482_, new_A9481_, new_A9480_, new_A9479_, new_A9478_, new_A9477_,
    new_A9476_, new_A9475_, new_A9474_, new_A9473_, new_A9472_, new_A9471_,
    new_A9470_, new_A9469_, new_A9468_, new_A9467_, new_A9466_, new_A9465_,
    new_A9464_, new_A9463_, new_A9462_, new_A9461_, new_A9460_, new_A9453_,
    new_A9452_, new_A9451_, new_A9450_, new_A9449_, new_A9448_, new_A9447_,
    new_A9446_, new_A9445_, new_A9444_, new_A9443_, new_A9442_, new_A9441_,
    new_A9440_, new_A9439_, new_A9438_, new_A9437_, new_A9436_, new_A9435_,
    new_A9434_, new_A9433_, new_A9432_, new_A9431_, new_A9430_, new_A9429_,
    new_A9428_, new_A9427_, new_A9426_, new_A9425_, new_A9424_, new_A9423_,
    new_A9422_, new_A9421_, new_A9420_, new_A9419_, new_A9418_, new_A9417_,
    new_A9416_, new_A9415_, new_A9414_, new_A9413_, new_A9412_, new_A9411_,
    new_A9410_, new_A9409_, new_A9408_, new_A9407_, new_A9406_, new_A9405_,
    new_A9404_, new_A9403_, new_A9402_, new_A9401_, new_A9400_, new_A9399_,
    new_A9398_, new_A9397_, new_A9396_, new_A9395_, new_A9394_, new_A9393_,
    new_A9386_, new_A9385_, new_A9384_, new_A9383_, new_A9382_, new_A9381_,
    new_A9380_, new_A9379_, new_A9378_, new_A9377_, new_A9376_, new_A9375_,
    new_A9374_, new_A9373_, new_A9372_, new_A9371_, new_A9370_, new_A9369_,
    new_A9368_, new_A9367_, new_A9366_, new_A9365_, new_A9364_, new_A9363_,
    new_A9362_, new_A9361_, new_A9360_, new_A9359_, new_A9358_, new_A9357_,
    new_A9356_, new_A9355_, new_A9354_, new_A9353_, new_A9352_, new_A9351_,
    new_A9350_, new_A9349_, new_A9348_, new_A9347_, new_A9346_, new_A9345_,
    new_A9344_, new_A9343_, new_A9342_, new_A9341_, new_A9340_, new_A9339_,
    new_A9338_, new_A9337_, new_A9336_, new_A9335_, new_A9334_, new_A9333_,
    new_A9332_, new_A9331_, new_A9330_, new_A9329_, new_A9328_, new_A9327_,
    new_A9326_, new_A9319_, new_A9318_, new_A9317_, new_A9316_, new_A9315_,
    new_A9314_, new_A9313_, new_A9312_, new_A9311_, new_A9310_, new_A9309_,
    new_A9308_, new_A9307_, new_A9306_, new_A9305_, new_A9304_, new_A9303_,
    new_A9302_, new_A9301_, new_A9300_, new_A9299_, new_A9298_, new_A9297_,
    new_A9296_, new_A9295_, new_A9294_, new_A9293_, new_A9292_, new_A9291_,
    new_A9290_, new_A9289_, new_A9288_, new_A9287_, new_A9286_, new_A9285_,
    new_A9284_, new_A9283_, new_A9282_, new_A9281_, new_A9280_, new_A9279_,
    new_A9278_, new_A9277_, new_A9276_, new_A9275_, new_A9274_, new_A9273_,
    new_A9272_, new_A9271_, new_A9270_, new_A9269_, new_A9268_, new_A9267_,
    new_A9266_, new_A9265_, new_A9264_, new_A9263_, new_A9262_, new_A9261_,
    new_A9260_, new_A9259_, new_A9252_, new_A9251_, new_A9250_, new_A9249_,
    new_A9248_, new_A9247_, new_A9246_, new_A9245_, new_A9244_, new_A9243_,
    new_A9242_, new_A9241_, new_A9240_, new_A9239_, new_A9238_, new_A9237_,
    new_A9236_, new_A9235_, new_A9234_, new_A9233_, new_A9232_, new_A9231_,
    new_A9230_, new_A9229_, new_A9228_, new_A9227_, new_A9226_, new_A9225_,
    new_A9224_, new_A9223_, new_A9222_, new_A9221_, new_A9220_, new_A9219_,
    new_A9218_, new_A9217_, new_A9216_, new_A9215_, new_A9214_, new_A9213_,
    new_A9212_, new_A9211_, new_A9210_, new_A9209_, new_A9208_, new_A9207_,
    new_A9206_, new_A9205_, new_A9204_, new_A9203_, new_A9202_, new_A9201_,
    new_A9200_, new_A9199_, new_A9198_, new_A9197_, new_A9196_, new_A9195_,
    new_A9194_, new_A9193_, new_A9192_, new_A9185_, new_A9184_, new_A9183_,
    new_A9182_, new_A9181_, new_A9180_, new_A9179_, new_A9178_, new_A9177_,
    new_A9176_, new_A9175_, new_A9174_, new_A9173_, new_A9172_, new_A9171_,
    new_A9170_, new_A9169_, new_A9168_, new_A9167_, new_A9166_, new_A9165_,
    new_A9164_, new_A9163_, new_A9162_, new_A9161_, new_A9160_, new_A9159_,
    new_A9158_, new_A9157_, new_A9156_, new_A9155_, new_A9154_, new_A9153_,
    new_A9152_, new_A9151_, new_A9150_, new_A9149_, new_A9148_, new_A9147_,
    new_A9146_, new_A9145_, new_A9144_, new_A9143_, new_A9142_, new_A9141_,
    new_A9140_, new_A9139_, new_A9138_, new_A9137_, new_A9136_, new_A9135_,
    new_A9134_, new_A9133_, new_A9132_, new_A9131_, new_A9130_, new_A9129_,
    new_A9128_, new_A9127_, new_A9126_, new_A9125_, new_A9118_, new_A9117_,
    new_A9116_, new_A9115_, new_A9114_, new_A9113_, new_A9112_, new_A9111_,
    new_A9110_, new_A9109_, new_A9108_, new_A9107_, new_A9106_, new_A9105_,
    new_A9104_, new_A9103_, new_A9102_, new_A9101_, new_A9100_, new_A9099_,
    new_A9098_, new_A9097_, new_A9096_, new_A9095_, new_A9094_, new_A9093_,
    new_A9092_, new_A9091_, new_A9090_, new_A9089_, new_A9088_, new_A9087_,
    new_A9086_, new_A9085_, new_A9084_, new_A9083_, new_A9082_, new_A9081_,
    new_A9080_, new_A9079_, new_A9078_, new_A9077_, new_A9076_, new_A9075_,
    new_A9074_, new_A9073_, new_A9072_, new_A9071_, new_A9070_, new_A9069_,
    new_A9068_, new_A9067_, new_A9066_, new_A9065_, new_A9064_, new_A9063_,
    new_A9062_, new_A9061_, new_A9060_, new_A9059_, new_A9058_, new_A9051_,
    new_A9050_, new_A9049_, new_A9048_, new_A9047_, new_A9046_, new_A9045_,
    new_A9044_, new_A9043_, new_A9042_, new_A9041_, new_A9040_, new_A9039_,
    new_A9038_, new_A9037_, new_A9036_, new_A9035_, new_A9034_, new_A9033_,
    new_A9032_, new_A9031_, new_A9030_, new_A9029_, new_A9028_, new_A9027_,
    new_A9026_, new_A9025_, new_A9024_, new_A9023_, new_A9022_, new_A9021_,
    new_A9020_, new_A9019_, new_A9018_, new_A9017_, new_A9016_, new_A9015_,
    new_A9014_, new_A9013_, new_A9012_, new_A9011_, new_A9010_, new_A9009_,
    new_A9008_, new_A9007_, new_A9006_, new_A9005_, new_A9004_, new_A9003_,
    new_A9002_, new_A9001_, new_A9000_, new_A8999_, new_A8998_, new_A8997_,
    new_A8996_, new_A8995_, new_A8994_, new_A8993_, new_A8992_, new_A8991_,
    new_A8984_, new_A8983_, new_A8982_, new_A8981_, new_A8980_, new_A8979_,
    new_A8978_, new_A8977_, new_A8976_, new_A8975_, new_A8974_, new_A8973_,
    new_A8972_, new_A8971_, new_A8970_, new_A8969_, new_A8968_, new_A8967_,
    new_A8966_, new_A8965_, new_A8964_, new_A8963_, new_A8962_, new_A8961_,
    new_A8960_, new_A8959_, new_A8958_, new_A8957_, new_A8956_, new_A8955_,
    new_A8954_, new_A8953_, new_A8952_, new_A8951_, new_A8950_, new_A8949_,
    new_A8948_, new_A8947_, new_A8946_, new_A8945_, new_A8944_, new_A8943_,
    new_A8942_, new_A8941_, new_A8940_, new_A8939_, new_A8938_, new_A8937_,
    new_A8936_, new_A8935_, new_A8934_, new_A8933_, new_A8932_, new_A8931_,
    new_A8930_, new_A8929_, new_A8928_, new_A8927_, new_A8926_, new_A8925_,
    new_A8924_, new_A8917_, new_A8916_, new_A8915_, new_A8914_, new_A8913_,
    new_A8912_, new_A8911_, new_A8910_, new_A8909_, new_A8908_, new_A8907_,
    new_A8906_, new_A8905_, new_A8904_, new_A8903_, new_A8902_, new_A8901_,
    new_A8900_, new_A8899_, new_A8898_, new_A8897_, new_A8896_, new_A8895_,
    new_A8894_, new_A8893_, new_A8892_, new_A8891_, new_A8890_, new_A8889_,
    new_A8888_, new_A8887_, new_A8886_, new_A8885_, new_A8884_, new_A8883_,
    new_A8882_, new_A8881_, new_A8880_, new_A8879_, new_A8878_, new_A8877_,
    new_A8876_, new_A8875_, new_A8874_, new_A8873_, new_A8872_, new_A8871_,
    new_A8870_, new_A8869_, new_A8868_, new_A8867_, new_A8866_, new_A8865_,
    new_A8864_, new_A8863_, new_A8862_, new_A8861_, new_A8860_, new_A8859_,
    new_A8858_, new_A8857_, new_A8850_, new_A8849_, new_A8848_, new_A8847_,
    new_A8846_, new_A8845_, new_A8844_, new_A8843_, new_A8842_, new_A8841_,
    new_A8840_, new_A8839_, new_A8838_, new_A8837_, new_A8836_, new_A8835_,
    new_A8834_, new_A8833_, new_A8832_, new_A8831_, new_A8830_, new_A8829_,
    new_A8828_, new_A8827_, new_A8826_, new_A8825_, new_A8824_, new_A8823_,
    new_A8822_, new_A8821_, new_A8820_, new_A8819_, new_A8818_, new_A8817_,
    new_A8816_, new_A8815_, new_A8814_, new_A8813_, new_A8812_, new_A8811_,
    new_A8810_, new_A8809_, new_A8808_, new_A8807_, new_A8806_, new_A8805_,
    new_A8804_, new_A8803_, new_A8802_, new_A8801_, new_A8800_, new_A8799_,
    new_A8798_, new_A8797_, new_A8796_, new_A8795_, new_A8794_, new_A8793_,
    new_A8792_, new_A8791_, new_A8790_, new_A8783_, new_A8782_, new_A8781_,
    new_A8780_, new_A8779_, new_A8778_, new_A8777_, new_A8776_, new_A8775_,
    new_A8774_, new_A8773_, new_A8772_, new_A8771_, new_A8770_, new_A8769_,
    new_A8768_, new_A8767_, new_A8766_, new_A8765_, new_A8764_, new_A8763_,
    new_A8762_, new_A8761_, new_A8760_, new_A8759_, new_A8758_, new_A8757_,
    new_A8756_, new_A8755_, new_A8754_, new_A8753_, new_A8752_, new_A8751_,
    new_A8750_, new_A8749_, new_A8748_, new_A8747_, new_A8746_, new_A8745_,
    new_A8744_, new_A8743_, new_A8742_, new_A8741_, new_A8740_, new_A8739_,
    new_A8738_, new_A8737_, new_A8736_, new_A8735_, new_A8734_, new_A8733_,
    new_A8732_, new_A8731_, new_A8730_, new_A8729_, new_A8728_, new_A8727_,
    new_A8726_, new_A8725_, new_A8724_, new_A8723_, new_A8716_, new_A8715_,
    new_A8714_, new_A8713_, new_A8712_, new_A8711_, new_A8710_, new_A8709_,
    new_A8708_, new_A8707_, new_A8706_, new_A8705_, new_A8704_, new_A8703_,
    new_A8702_, new_A8701_, new_A8700_, new_A8699_, new_A8698_, new_A8697_,
    new_A8696_, new_A8695_, new_A8694_, new_A8693_, new_A8692_, new_A8691_,
    new_A8690_, new_A8689_, new_A8688_, new_A8687_, new_A8686_, new_A8685_,
    new_A8684_, new_A8683_, new_A8682_, new_A8681_, new_A8680_, new_A8679_,
    new_A8678_, new_A8677_, new_A8676_, new_A8675_, new_A8674_, new_A8673_,
    new_A8672_, new_A8671_, new_A8670_, new_A8669_, new_A8668_, new_A8667_,
    new_A8666_, new_A8665_, new_A8664_, new_A8663_, new_A8662_, new_A8661_,
    new_A8660_, new_A8659_, new_A8658_, new_A8657_, new_A8656_, new_A8649_,
    new_A8648_, new_A8647_, new_A8646_, new_A8645_, new_A8644_, new_A8643_,
    new_A8642_, new_A8641_, new_A8640_, new_A8639_, new_A8638_, new_A8637_,
    new_A8636_, new_A8635_, new_A8634_, new_A8633_, new_A8632_, new_A8631_,
    new_A8630_, new_A8629_, new_A8628_, new_A8627_, new_A8626_, new_A8625_,
    new_A8624_, new_A8623_, new_A8622_, new_A8621_, new_A8620_, new_A8619_,
    new_A8618_, new_A8617_, new_A8616_, new_A8615_, new_A8614_, new_A8613_,
    new_A8612_, new_A8611_, new_A8610_, new_A8609_, new_A8608_, new_A8607_,
    new_A8606_, new_A8605_, new_A8604_, new_A8603_, new_A8602_, new_A8601_,
    new_A8600_, new_A8599_, new_A8598_, new_A8597_, new_A8596_, new_A8595_,
    new_A8594_, new_A8593_, new_A8592_, new_A8591_, new_A8590_, new_A8589_,
    new_A8582_, new_A8581_, new_A8580_, new_A8579_, new_A8578_, new_A8577_,
    new_A8576_, new_A8575_, new_A8574_, new_A8573_, new_A8572_, new_A8571_,
    new_A8570_, new_A8569_, new_A8568_, new_A8567_, new_A8566_, new_A8565_,
    new_A8564_, new_A8563_, new_A8562_, new_A8561_, new_A8560_, new_A8559_,
    new_A8558_, new_A8557_, new_A8556_, new_A8555_, new_A8554_, new_A8553_,
    new_A8552_, new_A8551_, new_A8550_, new_A8549_, new_A8548_, new_A8547_,
    new_A8546_, new_A8545_, new_A8544_, new_A8543_, new_A8542_, new_A8541_,
    new_A8540_, new_A8539_, new_A8538_, new_A8537_, new_A8536_, new_A8535_,
    new_A8534_, new_A8533_, new_A8532_, new_A8531_, new_A8530_, new_A8529_,
    new_A8528_, new_A8527_, new_A8526_, new_A8525_, new_A8524_, new_A8523_,
    new_A8522_, new_A8515_, new_A8514_, new_A8513_, new_A8512_, new_A8511_,
    new_A8510_, new_A8509_, new_A8508_, new_A8507_, new_A8506_, new_A8505_,
    new_A8504_, new_A8503_, new_A8502_, new_A8501_, new_A8500_, new_A8499_,
    new_A8498_, new_A8497_, new_A8496_, new_A8495_, new_A8494_, new_A8493_,
    new_A8492_, new_A8491_, new_A8490_, new_A8489_, new_A8488_, new_A8487_,
    new_A8486_, new_A8485_, new_A8484_, new_A8483_, new_A8482_, new_A8481_,
    new_A8480_, new_A8479_, new_A8478_, new_A8477_, new_A8476_, new_A8475_,
    new_A8474_, new_A8473_, new_A8472_, new_A8471_, new_A8470_, new_A8469_,
    new_A8468_, new_A8467_, new_A8466_, new_A8465_, new_A8464_, new_A8463_,
    new_A8462_, new_A8461_, new_A8460_, new_A8459_, new_A8458_, new_A8457_,
    new_A8456_, new_A8455_, new_A8448_, new_A8447_, new_A8446_, new_A8445_,
    new_A8444_, new_A8443_, new_A8442_, new_A8441_, new_A8440_, new_A8439_,
    new_A8438_, new_A8437_, new_A8436_, new_A8435_, new_A8434_, new_A8433_,
    new_A8432_, new_A8431_, new_A8430_, new_A8429_, new_A8428_, new_A8427_,
    new_A8426_, new_A8425_, new_A8424_, new_A8423_, new_A8422_, new_A8421_,
    new_A8420_, new_A8419_, new_A8418_, new_A8417_, new_A8416_, new_A8415_,
    new_A8414_, new_A8413_, new_A8412_, new_A8411_, new_A8410_, new_A8409_,
    new_A8408_, new_A8407_, new_A8406_, new_A8405_, new_A8404_, new_A8403_,
    new_A8402_, new_A8401_, new_A8400_, new_A8399_, new_A8398_, new_A8397_,
    new_A8396_, new_A8395_, new_A8394_, new_A8393_, new_A8392_, new_A8391_,
    new_A8390_, new_A8389_, new_A8388_, new_A8381_, new_A8380_, new_A8379_,
    new_A8378_, new_A8377_, new_A8376_, new_A8375_, new_A8374_, new_A8373_,
    new_A8372_, new_A8371_, new_A8370_, new_A8369_, new_A8368_, new_A8367_,
    new_A8366_, new_A8365_, new_A8364_, new_A8363_, new_A8362_, new_A8361_,
    new_A8360_, new_A8359_, new_A8358_, new_A8357_, new_A8356_, new_A8355_,
    new_A8354_, new_A8353_, new_A8352_, new_A8351_, new_A8350_, new_A8349_,
    new_A8348_, new_A8347_, new_A8346_, new_A8345_, new_A8344_, new_A8343_,
    new_A8342_, new_A8341_, new_A8340_, new_A8339_, new_A8338_, new_A8337_,
    new_A8336_, new_A8335_, new_A8334_, new_A8333_, new_A8332_, new_A8331_,
    new_A8330_, new_A8329_, new_A8328_, new_A8327_, new_A8326_, new_A8325_,
    new_A8324_, new_A8323_, new_A8322_, new_A8321_, new_A8314_, new_A8313_,
    new_A8312_, new_A8311_, new_A8310_, new_A8309_, new_A8308_, new_A8307_,
    new_A8306_, new_A8305_, new_A8304_, new_A8303_, new_A8302_, new_A8301_,
    new_A8300_, new_A8299_, new_A8298_, new_A8297_, new_A8296_, new_A8295_,
    new_A8294_, new_A8293_, new_A8292_, new_A8291_, new_A8290_, new_A8289_,
    new_A8288_, new_A8287_, new_A8286_, new_A8285_, new_A8284_, new_A8283_,
    new_A8282_, new_A8281_, new_A8280_, new_A8279_, new_A8278_, new_A8277_,
    new_A8276_, new_A8275_, new_A8274_, new_A8273_, new_A8272_, new_A8271_,
    new_A8270_, new_A8269_, new_A8268_, new_A8267_, new_A8266_, new_A8265_,
    new_A8264_, new_A8263_, new_A8262_, new_A8261_, new_A8260_, new_A8259_,
    new_A8258_, new_A8257_, new_A8256_, new_A8255_, new_A8254_, new_A8247_,
    new_A8246_, new_A8245_, new_A8244_, new_A8243_, new_A8242_, new_A8241_,
    new_A8240_, new_A8239_, new_A8238_, new_A8237_, new_A8236_, new_A8235_,
    new_A8234_, new_A8233_, new_A8232_, new_A8231_, new_A8230_, new_A8229_,
    new_A8228_, new_A8227_, new_A8226_, new_A8225_, new_A8224_, new_A8223_,
    new_A8222_, new_A8221_, new_A8220_, new_A8219_, new_A8218_, new_A8217_,
    new_A8216_, new_A8215_, new_A8214_, new_A8213_, new_A8212_, new_A8211_,
    new_A8210_, new_A8209_, new_A8208_, new_A8207_, new_A8206_, new_A8205_,
    new_A8204_, new_A8203_, new_A8202_, new_A8201_, new_A8200_, new_A8199_,
    new_A8198_, new_A8197_, new_A8196_, new_A8195_, new_A8194_, new_A8193_,
    new_A8192_, new_A8191_, new_A8190_, new_A8189_, new_A8188_, new_A8187_,
    new_A8180_, new_A8179_, new_A8178_, new_A8177_, new_A8176_, new_A8175_,
    new_A8174_, new_A8173_, new_A8172_, new_A8171_, new_A8170_, new_A8169_,
    new_A8168_, new_A8167_, new_A8166_, new_A8165_, new_A8164_, new_A8163_,
    new_A8162_, new_A8161_, new_A8160_, new_A8159_, new_A8158_, new_A8157_,
    new_A8156_, new_A8155_, new_A8154_, new_A8153_, new_A8152_, new_A8151_,
    new_A8150_, new_A8149_, new_A8148_, new_A8147_, new_A8146_, new_A8145_,
    new_A8144_, new_A8143_, new_A8142_, new_A8141_, new_A8140_, new_A8139_,
    new_A8138_, new_A8137_, new_A8136_, new_A8135_, new_A8134_, new_A8133_,
    new_A8132_, new_A8131_, new_A8130_, new_A8129_, new_A8128_, new_A8127_,
    new_A8126_, new_A8125_, new_A8124_, new_A8123_, new_A8122_, new_A8121_,
    new_A8120_, new_A8113_, new_A8112_, new_A8111_, new_A8110_, new_A8109_,
    new_A8108_, new_A8041_, new_A8042_, new_A8043_, new_A8044_, new_A8045_,
    new_A8046_, new_A8053_, new_A8054_, new_A8055_, new_A8056_, new_A8057_,
    new_A8058_, new_A8059_, new_A8060_, new_A8061_, new_A8062_, new_A8063_,
    new_A8064_, new_A8065_, new_A8066_, new_A8067_, new_A8068_, new_A8069_,
    new_A8070_, new_A8071_, new_A8072_, new_A8073_, new_A8074_, new_A8075_,
    new_A8076_, new_A8077_, new_A8078_, new_A8079_, new_A8080_, new_A8081_,
    new_A8082_, new_A8083_, new_A8084_, new_A8085_, new_A8086_, new_A8087_,
    new_A8088_, new_A8089_, new_A8090_, new_A8091_, new_A8092_, new_A8093_,
    new_A8094_, new_A8095_, new_A8096_, new_A8097_, new_A8098_, new_A8099_,
    new_A8100_, new_A8101_, new_A8102_, new_A8103_, new_A8104_, new_A8105_,
    new_A8106_, new_A8107_;
  assign new_F1528_ = ~F1467 & new_F1481_;
  assign new_F1527_ = F1467 & ~new_F1481_;
  assign new_F1526_ = F1467 & ~new_F1481_;
  assign new_F1525_ = ~F1467 & ~new_F1481_;
  assign new_F1524_ = F1467 & new_F1481_;
  assign new_F1523_ = new_F1527_ | new_F1528_;
  assign new_F1522_ = ~F1467 & new_F1481_;
  assign new_F1521_ = new_F1525_ | new_F1526_;
  assign new_F1520_ = ~new_F1496_ & ~new_F1516_;
  assign new_F1519_ = new_F1496_ & new_F1516_;
  assign new_F1518_ = ~F1463 | ~new_F1488_;
  assign new_F1517_ = new_F1481_ & new_F1518_;
  assign new_F1516_ = F1464 | F1465;
  assign new_F1515_ = F1464 | new_F1481_;
  assign new_F1514_ = ~new_F1481_ & ~new_F1517_;
  assign new_F1513_ = new_F1481_ | new_F1518_;
  assign new_F1512_ = F1464 & ~F1465;
  assign new_F1511_ = ~F1464 & F1465;
  assign new_F1510_ = new_F1474_ | new_F1507_;
  assign new_F1509_ = ~new_F1474_ & ~new_F1508_;
  assign new_F1508_ = new_F1474_ & new_F1507_;
  assign new_F1507_ = ~F1463 | ~new_F1488_;
  assign new_F1506_ = ~F1464 & new_F1474_;
  assign new_F1505_ = F1464 & ~new_F1474_;
  assign new_F1504_ = F1466 & new_F1503_;
  assign new_F1503_ = new_F1522_ | new_F1521_;
  assign new_F1502_ = ~F1466 & new_F1501_;
  assign new_F1501_ = new_F1524_ | new_F1523_;
  assign new_F1500_ = F1466 | new_F1499_;
  assign new_F1499_ = new_F1520_ | new_F1519_;
  assign new_F1498_ = ~new_F1478_ & ~new_F1488_;
  assign new_F1497_ = new_F1478_ & new_F1488_;
  assign new_F1496_ = ~new_F1478_ | new_F1488_;
  assign new_F1495_ = F1462 & ~F1463;
  assign new_F1494_ = ~F1462 & F1463;
  assign new_F1493_ = new_F1515_ & ~new_F1516_;
  assign new_F1492_ = ~new_F1515_ & new_F1516_;
  assign new_F1491_ = ~new_F1514_ | ~new_F1513_;
  assign new_F1490_ = new_F1506_ | new_F1505_;
  assign new_F1489_ = new_F1512_ | new_F1511_;
  assign new_F1488_ = new_F1502_ | new_F1504_;
  assign new_F1487_ = ~new_F1509_ | ~new_F1510_;
  assign new_F1486_ = F1462 & ~F1463;
  assign new_F1485_ = new_F1476_ & ~new_F1488_;
  assign new_F1484_ = ~new_F1476_ & new_F1488_;
  assign new_F1483_ = ~new_F1474_ & new_F1500_;
  assign new_F1482_ = new_F1498_ | new_F1497_;
  assign new_F1481_ = new_F1495_ | new_F1494_;
  assign new_F1480_ = F1463 | new_F1496_;
  assign new_F1479_ = new_F1488_ & new_F1491_;
  assign new_F1478_ = new_F1493_ | new_F1492_;
  assign new_F1477_ = new_F1488_ & new_F1487_;
  assign new_F1476_ = new_F1490_ & new_F1489_;
  assign new_F1475_ = new_F1485_ | new_F1484_;
  assign new_F1474_ = F1463 | new_F1486_;
  assign new_F1473_ = new_F1474_ | new_F1483_;
  assign new_F1472_ = new_F1481_ & new_F1482_;
  assign new_F1471_ = new_F1481_ & new_F1480_;
  assign new_F1470_ = new_F1479_ | new_F1478_;
  assign new_F1469_ = new_F1477_ | new_F1476_;
  assign new_F1468_ = new_F1475_ & new_F1474_;
  assign new_F1535_ = new_F1542_ & new_F1541_;
  assign new_F1536_ = new_F1544_ | new_F1543_;
  assign new_F1537_ = new_F1546_ | new_F1545_;
  assign new_F1538_ = new_F1548_ & new_F1547_;
  assign new_F1539_ = new_F1548_ & new_F1549_;
  assign new_F1540_ = new_F1541_ | new_F1550_;
  assign new_F1541_ = F1530 | new_F1553_;
  assign new_F1542_ = new_F1552_ | new_F1551_;
  assign new_F1543_ = new_F1557_ & new_F1556_;
  assign new_F1544_ = new_F1555_ & new_F1554_;
  assign new_F1545_ = new_F1560_ | new_F1559_;
  assign new_F1546_ = new_F1555_ & new_F1558_;
  assign new_F1547_ = F1530 | new_F1563_;
  assign new_F1548_ = new_F1562_ | new_F1561_;
  assign new_F1549_ = new_F1565_ | new_F1564_;
  assign new_F1550_ = ~new_F1541_ & new_F1567_;
  assign new_F1551_ = ~new_F1543_ & new_F1555_;
  assign new_F1552_ = new_F1543_ & ~new_F1555_;
  assign new_F1553_ = F1529 & ~F1530;
  assign new_F1554_ = ~new_F1576_ | ~new_F1577_;
  assign new_F1555_ = new_F1569_ | new_F1571_;
  assign new_F1556_ = new_F1579_ | new_F1578_;
  assign new_F1557_ = new_F1573_ | new_F1572_;
  assign new_F1558_ = ~new_F1581_ | ~new_F1580_;
  assign new_F1559_ = ~new_F1582_ & new_F1583_;
  assign new_F1560_ = new_F1582_ & ~new_F1583_;
  assign new_F1561_ = ~F1529 & F1530;
  assign new_F1562_ = F1529 & ~F1530;
  assign new_F1563_ = ~new_F1545_ | new_F1555_;
  assign new_F1564_ = new_F1545_ & new_F1555_;
  assign new_F1565_ = ~new_F1545_ & ~new_F1555_;
  assign new_F1566_ = new_F1587_ | new_F1586_;
  assign new_F1567_ = F1533 | new_F1566_;
  assign new_F1568_ = new_F1591_ | new_F1590_;
  assign new_F1569_ = ~F1533 & new_F1568_;
  assign new_F1570_ = new_F1589_ | new_F1588_;
  assign new_F1571_ = F1533 & new_F1570_;
  assign new_F1572_ = F1531 & ~new_F1541_;
  assign new_F1573_ = ~F1531 & new_F1541_;
  assign new_F1574_ = ~F1530 | ~new_F1555_;
  assign new_F1575_ = new_F1541_ & new_F1574_;
  assign new_F1576_ = ~new_F1541_ & ~new_F1575_;
  assign new_F1577_ = new_F1541_ | new_F1574_;
  assign new_F1578_ = ~F1531 & F1532;
  assign new_F1579_ = F1531 & ~F1532;
  assign new_F1580_ = new_F1548_ | new_F1585_;
  assign new_F1581_ = ~new_F1548_ & ~new_F1584_;
  assign new_F1582_ = F1531 | new_F1548_;
  assign new_F1583_ = F1531 | F1532;
  assign new_F1584_ = new_F1548_ & new_F1585_;
  assign new_F1585_ = ~F1530 | ~new_F1555_;
  assign new_F1586_ = new_F1563_ & new_F1583_;
  assign new_F1587_ = ~new_F1563_ & ~new_F1583_;
  assign new_F1588_ = new_F1592_ | new_F1593_;
  assign new_F1589_ = ~F1534 & new_F1548_;
  assign new_F1590_ = new_F1594_ | new_F1595_;
  assign new_F1591_ = F1534 & new_F1548_;
  assign new_F1592_ = ~F1534 & ~new_F1548_;
  assign new_F1593_ = F1534 & ~new_F1548_;
  assign new_F1594_ = F1534 & ~new_F1548_;
  assign new_F1595_ = ~F1534 & new_F1548_;
  assign new_F1602_ = new_F1609_ & new_F1608_;
  assign new_F1603_ = new_F1611_ | new_F1610_;
  assign new_F1604_ = new_F1613_ | new_F1612_;
  assign new_F1605_ = new_F1615_ & new_F1614_;
  assign new_F1606_ = new_F1615_ & new_F1616_;
  assign new_F1607_ = new_F1608_ | new_F1617_;
  assign new_F1608_ = F1597 | new_F1620_;
  assign new_F1609_ = new_F1619_ | new_F1618_;
  assign new_F1610_ = new_F1624_ & new_F1623_;
  assign new_F1611_ = new_F1622_ & new_F1621_;
  assign new_F1612_ = new_F1627_ | new_F1626_;
  assign new_F1613_ = new_F1622_ & new_F1625_;
  assign new_F1614_ = F1597 | new_F1630_;
  assign new_F1615_ = new_F1629_ | new_F1628_;
  assign new_F1616_ = new_F1632_ | new_F1631_;
  assign new_F1617_ = ~new_F1608_ & new_F1634_;
  assign new_F1618_ = ~new_F1610_ & new_F1622_;
  assign new_F1619_ = new_F1610_ & ~new_F1622_;
  assign new_F1620_ = F1596 & ~F1597;
  assign new_F1621_ = ~new_F1643_ | ~new_F1644_;
  assign new_F1622_ = new_F1636_ | new_F1638_;
  assign new_F1623_ = new_F1646_ | new_F1645_;
  assign new_F1624_ = new_F1640_ | new_F1639_;
  assign new_F1625_ = ~new_F1648_ | ~new_F1647_;
  assign new_F1626_ = ~new_F1649_ & new_F1650_;
  assign new_F1627_ = new_F1649_ & ~new_F1650_;
  assign new_F1628_ = ~F1596 & F1597;
  assign new_F1629_ = F1596 & ~F1597;
  assign new_F1630_ = ~new_F1612_ | new_F1622_;
  assign new_F1631_ = new_F1612_ & new_F1622_;
  assign new_F1632_ = ~new_F1612_ & ~new_F1622_;
  assign new_F1633_ = new_F1654_ | new_F1653_;
  assign new_F1634_ = F1600 | new_F1633_;
  assign new_F1635_ = new_F1658_ | new_F1657_;
  assign new_F1636_ = ~F1600 & new_F1635_;
  assign new_F1637_ = new_F1656_ | new_F1655_;
  assign new_F1638_ = F1600 & new_F1637_;
  assign new_F1639_ = F1598 & ~new_F1608_;
  assign new_F1640_ = ~F1598 & new_F1608_;
  assign new_F1641_ = ~F1597 | ~new_F1622_;
  assign new_F1642_ = new_F1608_ & new_F1641_;
  assign new_F1643_ = ~new_F1608_ & ~new_F1642_;
  assign new_F1644_ = new_F1608_ | new_F1641_;
  assign new_F1645_ = ~F1598 & F1599;
  assign new_F1646_ = F1598 & ~F1599;
  assign new_F1647_ = new_F1615_ | new_F1652_;
  assign new_F1648_ = ~new_F1615_ & ~new_F1651_;
  assign new_F1649_ = F1598 | new_F1615_;
  assign new_F1650_ = F1598 | F1599;
  assign new_F1651_ = new_F1615_ & new_F1652_;
  assign new_F1652_ = ~F1597 | ~new_F1622_;
  assign new_F1653_ = new_F1630_ & new_F1650_;
  assign new_F1654_ = ~new_F1630_ & ~new_F1650_;
  assign new_F1655_ = new_F1659_ | new_F1660_;
  assign new_F1656_ = ~F1601 & new_F1615_;
  assign new_F1657_ = new_F1661_ | new_F1662_;
  assign new_F1658_ = F1601 & new_F1615_;
  assign new_F1659_ = ~F1601 & ~new_F1615_;
  assign new_F1660_ = F1601 & ~new_F1615_;
  assign new_F1661_ = F1601 & ~new_F1615_;
  assign new_F1662_ = ~F1601 & new_F1615_;
  assign new_F1669_ = new_F1676_ & new_F1675_;
  assign new_F1670_ = new_F1678_ | new_F1677_;
  assign new_F1671_ = new_F1680_ | new_F1679_;
  assign new_F1672_ = new_F1682_ & new_F1681_;
  assign new_F1673_ = new_F1682_ & new_F1683_;
  assign new_F1674_ = new_F1675_ | new_F1684_;
  assign new_F1675_ = F1664 | new_F1687_;
  assign new_F1676_ = new_F1686_ | new_F1685_;
  assign new_F1677_ = new_F1691_ & new_F1690_;
  assign new_F1678_ = new_F1689_ & new_F1688_;
  assign new_F1679_ = new_F1694_ | new_F1693_;
  assign new_F1680_ = new_F1689_ & new_F1692_;
  assign new_F1681_ = F1664 | new_F1697_;
  assign new_F1682_ = new_F1696_ | new_F1695_;
  assign new_F1683_ = new_F1699_ | new_F1698_;
  assign new_F1684_ = ~new_F1675_ & new_F1701_;
  assign new_F1685_ = ~new_F1677_ & new_F1689_;
  assign new_F1686_ = new_F1677_ & ~new_F1689_;
  assign new_F1687_ = F1663 & ~F1664;
  assign new_F1688_ = ~new_F1710_ | ~new_F1711_;
  assign new_F1689_ = new_F1703_ | new_F1705_;
  assign new_F1690_ = new_F1713_ | new_F1712_;
  assign new_F1691_ = new_F1707_ | new_F1706_;
  assign new_F1692_ = ~new_F1715_ | ~new_F1714_;
  assign new_F1693_ = ~new_F1716_ & new_F1717_;
  assign new_F1694_ = new_F1716_ & ~new_F1717_;
  assign new_F1695_ = ~F1663 & F1664;
  assign new_F1696_ = F1663 & ~F1664;
  assign new_F1697_ = ~new_F1679_ | new_F1689_;
  assign new_F1698_ = new_F1679_ & new_F1689_;
  assign new_F1699_ = ~new_F1679_ & ~new_F1689_;
  assign new_F1700_ = new_F1721_ | new_F1720_;
  assign new_F1701_ = F1667 | new_F1700_;
  assign new_F1702_ = new_F1725_ | new_F1724_;
  assign new_F1703_ = ~F1667 & new_F1702_;
  assign new_F1704_ = new_F1723_ | new_F1722_;
  assign new_F1705_ = F1667 & new_F1704_;
  assign new_F1706_ = F1665 & ~new_F1675_;
  assign new_F1707_ = ~F1665 & new_F1675_;
  assign new_F1708_ = ~F1664 | ~new_F1689_;
  assign new_F1709_ = new_F1675_ & new_F1708_;
  assign new_F1710_ = ~new_F1675_ & ~new_F1709_;
  assign new_F1711_ = new_F1675_ | new_F1708_;
  assign new_F1712_ = ~F1665 & F1666;
  assign new_F1713_ = F1665 & ~F1666;
  assign new_F1714_ = new_F1682_ | new_F1719_;
  assign new_F1715_ = ~new_F1682_ & ~new_F1718_;
  assign new_F1716_ = F1665 | new_F1682_;
  assign new_F1717_ = F1665 | F1666;
  assign new_F1718_ = new_F1682_ & new_F1719_;
  assign new_F1719_ = ~F1664 | ~new_F1689_;
  assign new_F1720_ = new_F1697_ & new_F1717_;
  assign new_F1721_ = ~new_F1697_ & ~new_F1717_;
  assign new_F1722_ = new_F1726_ | new_F1727_;
  assign new_F1723_ = ~F1668 & new_F1682_;
  assign new_F1724_ = new_F1728_ | new_F1729_;
  assign new_F1725_ = F1668 & new_F1682_;
  assign new_F1726_ = ~F1668 & ~new_F1682_;
  assign new_F1727_ = F1668 & ~new_F1682_;
  assign new_F1728_ = F1668 & ~new_F1682_;
  assign new_F1729_ = ~F1668 & new_F1682_;
  assign new_F1736_ = new_F1743_ & new_F1742_;
  assign new_F1737_ = new_F1745_ | new_F1744_;
  assign new_F1738_ = new_F1747_ | new_F1746_;
  assign new_F1739_ = new_F1749_ & new_F1748_;
  assign new_F1740_ = new_F1749_ & new_F1750_;
  assign new_F1741_ = new_F1742_ | new_F1751_;
  assign new_F1742_ = F1731 | new_F1754_;
  assign new_F1743_ = new_F1753_ | new_F1752_;
  assign new_F1744_ = new_F1758_ & new_F1757_;
  assign new_F1745_ = new_F1756_ & new_F1755_;
  assign new_F1746_ = new_F1761_ | new_F1760_;
  assign new_F1747_ = new_F1756_ & new_F1759_;
  assign new_F1748_ = F1731 | new_F1764_;
  assign new_F1749_ = new_F1763_ | new_F1762_;
  assign new_F1750_ = new_F1766_ | new_F1765_;
  assign new_F1751_ = ~new_F1742_ & new_F1768_;
  assign new_F1752_ = ~new_F1744_ & new_F1756_;
  assign new_F1753_ = new_F1744_ & ~new_F1756_;
  assign new_F1754_ = F1730 & ~F1731;
  assign new_F1755_ = ~new_F1777_ | ~new_F1778_;
  assign new_F1756_ = new_F1770_ | new_F1772_;
  assign new_F1757_ = new_F1780_ | new_F1779_;
  assign new_F1758_ = new_F1774_ | new_F1773_;
  assign new_F1759_ = ~new_F1782_ | ~new_F1781_;
  assign new_F1760_ = ~new_F1783_ & new_F1784_;
  assign new_F1761_ = new_F1783_ & ~new_F1784_;
  assign new_F1762_ = ~F1730 & F1731;
  assign new_F1763_ = F1730 & ~F1731;
  assign new_F1764_ = ~new_F1746_ | new_F1756_;
  assign new_F1765_ = new_F1746_ & new_F1756_;
  assign new_F1766_ = ~new_F1746_ & ~new_F1756_;
  assign new_F1767_ = new_F1788_ | new_F1787_;
  assign new_F1768_ = F1734 | new_F1767_;
  assign new_F1769_ = new_F1792_ | new_F1791_;
  assign new_F1770_ = ~F1734 & new_F1769_;
  assign new_F1771_ = new_F1790_ | new_F1789_;
  assign new_F1772_ = F1734 & new_F1771_;
  assign new_F1773_ = F1732 & ~new_F1742_;
  assign new_F1774_ = ~F1732 & new_F1742_;
  assign new_F1775_ = ~F1731 | ~new_F1756_;
  assign new_F1776_ = new_F1742_ & new_F1775_;
  assign new_F1777_ = ~new_F1742_ & ~new_F1776_;
  assign new_F1778_ = new_F1742_ | new_F1775_;
  assign new_F1779_ = ~F1732 & F1733;
  assign new_F1780_ = F1732 & ~F1733;
  assign new_F1781_ = new_F1749_ | new_F1786_;
  assign new_F1782_ = ~new_F1749_ & ~new_F1785_;
  assign new_F1783_ = F1732 | new_F1749_;
  assign new_F1784_ = F1732 | F1733;
  assign new_F1785_ = new_F1749_ & new_F1786_;
  assign new_F1786_ = ~F1731 | ~new_F1756_;
  assign new_F1787_ = new_F1764_ & new_F1784_;
  assign new_F1788_ = ~new_F1764_ & ~new_F1784_;
  assign new_F1789_ = new_F1793_ | new_F1794_;
  assign new_F1790_ = ~F1735 & new_F1749_;
  assign new_F1791_ = new_F1795_ | new_F1796_;
  assign new_F1792_ = F1735 & new_F1749_;
  assign new_F1793_ = ~F1735 & ~new_F1749_;
  assign new_F1794_ = F1735 & ~new_F1749_;
  assign new_F1795_ = F1735 & ~new_F1749_;
  assign new_F1796_ = ~F1735 & new_F1749_;
  assign new_F1803_ = new_F1810_ & new_F1809_;
  assign new_F1804_ = new_F1812_ | new_F1811_;
  assign new_F1805_ = new_F1814_ | new_F1813_;
  assign new_F1806_ = new_F1816_ & new_F1815_;
  assign new_F1807_ = new_F1816_ & new_F1817_;
  assign new_F1808_ = new_F1809_ | new_F1818_;
  assign new_F1809_ = F1798 | new_F1821_;
  assign new_F1810_ = new_F1820_ | new_F1819_;
  assign new_F1811_ = new_F1825_ & new_F1824_;
  assign new_F1812_ = new_F1823_ & new_F1822_;
  assign new_F1813_ = new_F1828_ | new_F1827_;
  assign new_F1814_ = new_F1823_ & new_F1826_;
  assign new_F1815_ = F1798 | new_F1831_;
  assign new_F1816_ = new_F1830_ | new_F1829_;
  assign new_F1817_ = new_F1833_ | new_F1832_;
  assign new_F1818_ = ~new_F1809_ & new_F1835_;
  assign new_F1819_ = ~new_F1811_ & new_F1823_;
  assign new_F1820_ = new_F1811_ & ~new_F1823_;
  assign new_F1821_ = F1797 & ~F1798;
  assign new_F1822_ = ~new_F1844_ | ~new_F1845_;
  assign new_F1823_ = new_F1837_ | new_F1839_;
  assign new_F1824_ = new_F1847_ | new_F1846_;
  assign new_F1825_ = new_F1841_ | new_F1840_;
  assign new_F1826_ = ~new_F1849_ | ~new_F1848_;
  assign new_F1827_ = ~new_F1850_ & new_F1851_;
  assign new_F1828_ = new_F1850_ & ~new_F1851_;
  assign new_F1829_ = ~F1797 & F1798;
  assign new_F1830_ = F1797 & ~F1798;
  assign new_F1831_ = ~new_F1813_ | new_F1823_;
  assign new_F1832_ = new_F1813_ & new_F1823_;
  assign new_F1833_ = ~new_F1813_ & ~new_F1823_;
  assign new_F1834_ = new_F1855_ | new_F1854_;
  assign new_F1835_ = F1801 | new_F1834_;
  assign new_F1836_ = new_F1859_ | new_F1858_;
  assign new_F1837_ = ~F1801 & new_F1836_;
  assign new_F1838_ = new_F1857_ | new_F1856_;
  assign new_F1839_ = F1801 & new_F1838_;
  assign new_F1840_ = F1799 & ~new_F1809_;
  assign new_F1841_ = ~F1799 & new_F1809_;
  assign new_F1842_ = ~F1798 | ~new_F1823_;
  assign new_F1843_ = new_F1809_ & new_F1842_;
  assign new_F1844_ = ~new_F1809_ & ~new_F1843_;
  assign new_F1845_ = new_F1809_ | new_F1842_;
  assign new_F1846_ = ~F1799 & F1800;
  assign new_F1847_ = F1799 & ~F1800;
  assign new_F1848_ = new_F1816_ | new_F1853_;
  assign new_F1849_ = ~new_F1816_ & ~new_F1852_;
  assign new_F1850_ = F1799 | new_F1816_;
  assign new_F1851_ = F1799 | F1800;
  assign new_F1852_ = new_F1816_ & new_F1853_;
  assign new_F1853_ = ~F1798 | ~new_F1823_;
  assign new_F1854_ = new_F1831_ & new_F1851_;
  assign new_F1855_ = ~new_F1831_ & ~new_F1851_;
  assign new_F1856_ = new_F1860_ | new_F1861_;
  assign new_F1857_ = ~F1802 & new_F1816_;
  assign new_F1858_ = new_F1862_ | new_F1863_;
  assign new_F1859_ = F1802 & new_F1816_;
  assign new_F1860_ = ~F1802 & ~new_F1816_;
  assign new_F1861_ = F1802 & ~new_F1816_;
  assign new_F1862_ = F1802 & ~new_F1816_;
  assign new_F1863_ = ~F1802 & new_F1816_;
  assign new_F1870_ = new_F1877_ & new_F1876_;
  assign new_F1871_ = new_F1879_ | new_F1878_;
  assign new_F1872_ = new_F1881_ | new_F1880_;
  assign new_F1873_ = new_F1883_ & new_F1882_;
  assign new_F1874_ = new_F1883_ & new_F1884_;
  assign new_F1875_ = new_F1876_ | new_F1885_;
  assign new_F1876_ = F1865 | new_F1888_;
  assign new_F1877_ = new_F1887_ | new_F1886_;
  assign new_F1878_ = new_F1892_ & new_F1891_;
  assign new_F1879_ = new_F1890_ & new_F1889_;
  assign new_F1880_ = new_F1895_ | new_F1894_;
  assign new_F1881_ = new_F1890_ & new_F1893_;
  assign new_F1882_ = F1865 | new_F1898_;
  assign new_F1883_ = new_F1897_ | new_F1896_;
  assign new_F1884_ = new_F1900_ | new_F1899_;
  assign new_F1885_ = ~new_F1876_ & new_F1902_;
  assign new_F1886_ = ~new_F1878_ & new_F1890_;
  assign new_F1887_ = new_F1878_ & ~new_F1890_;
  assign new_F1888_ = F1864 & ~F1865;
  assign new_F1889_ = ~new_F1911_ | ~new_F1912_;
  assign new_F1890_ = new_F1904_ | new_F1906_;
  assign new_F1891_ = new_F1914_ | new_F1913_;
  assign new_F1892_ = new_F1908_ | new_F1907_;
  assign new_F1893_ = ~new_F1916_ | ~new_F1915_;
  assign new_F1894_ = ~new_F1917_ & new_F1918_;
  assign new_F1895_ = new_F1917_ & ~new_F1918_;
  assign new_F1896_ = ~F1864 & F1865;
  assign new_F1897_ = F1864 & ~F1865;
  assign new_F1898_ = ~new_F1880_ | new_F1890_;
  assign new_F1899_ = new_F1880_ & new_F1890_;
  assign new_F1900_ = ~new_F1880_ & ~new_F1890_;
  assign new_F1901_ = new_F1922_ | new_F1921_;
  assign new_F1902_ = F1868 | new_F1901_;
  assign new_F1903_ = new_F1926_ | new_F1925_;
  assign new_F1904_ = ~F1868 & new_F1903_;
  assign new_F1905_ = new_F1924_ | new_F1923_;
  assign new_F1906_ = F1868 & new_F1905_;
  assign new_F1907_ = F1866 & ~new_F1876_;
  assign new_F1908_ = ~F1866 & new_F1876_;
  assign new_F1909_ = ~F1865 | ~new_F1890_;
  assign new_F1910_ = new_F1876_ & new_F1909_;
  assign new_F1911_ = ~new_F1876_ & ~new_F1910_;
  assign new_F1912_ = new_F1876_ | new_F1909_;
  assign new_F1913_ = ~F1866 & F1867;
  assign new_F1914_ = F1866 & ~F1867;
  assign new_F1915_ = new_F1883_ | new_F1920_;
  assign new_F1916_ = ~new_F1883_ & ~new_F1919_;
  assign new_F1917_ = F1866 | new_F1883_;
  assign new_F1918_ = F1866 | F1867;
  assign new_F1919_ = new_F1883_ & new_F1920_;
  assign new_F1920_ = ~F1865 | ~new_F1890_;
  assign new_F1921_ = new_F1898_ & new_F1918_;
  assign new_F1922_ = ~new_F1898_ & ~new_F1918_;
  assign new_F1923_ = new_F1927_ | new_F1928_;
  assign new_F1924_ = ~F1869 & new_F1883_;
  assign new_F1925_ = new_F1929_ | new_F1930_;
  assign new_F1926_ = F1869 & new_F1883_;
  assign new_F1927_ = ~F1869 & ~new_F1883_;
  assign new_F1928_ = F1869 & ~new_F1883_;
  assign new_F1929_ = F1869 & ~new_F1883_;
  assign new_F1930_ = ~F1869 & new_F1883_;
  assign new_F1937_ = new_F1944_ & new_F1943_;
  assign new_F1938_ = new_F1946_ | new_F1945_;
  assign new_F1939_ = new_F1948_ | new_F1947_;
  assign new_F1940_ = new_F1950_ & new_F1949_;
  assign new_F1941_ = new_F1950_ & new_F1951_;
  assign new_F1942_ = new_F1943_ | new_F1952_;
  assign new_F1943_ = F1932 | new_F1955_;
  assign new_F1944_ = new_F1954_ | new_F1953_;
  assign new_F1945_ = new_F1959_ & new_F1958_;
  assign new_F1946_ = new_F1957_ & new_F1956_;
  assign new_F1947_ = new_F1962_ | new_F1961_;
  assign new_F1948_ = new_F1957_ & new_F1960_;
  assign new_F1949_ = F1932 | new_F1965_;
  assign new_F1950_ = new_F1964_ | new_F1963_;
  assign new_F1951_ = new_F1967_ | new_F1966_;
  assign new_F1952_ = ~new_F1943_ & new_F1969_;
  assign new_F1953_ = ~new_F1945_ & new_F1957_;
  assign new_F1954_ = new_F1945_ & ~new_F1957_;
  assign new_F1955_ = F1931 & ~F1932;
  assign new_F1956_ = ~new_F1978_ | ~new_F1979_;
  assign new_F1957_ = new_F1971_ | new_F1973_;
  assign new_F1958_ = new_F1981_ | new_F1980_;
  assign new_F1959_ = new_F1975_ | new_F1974_;
  assign new_F1960_ = ~new_F1983_ | ~new_F1982_;
  assign new_F1961_ = ~new_F1984_ & new_F1985_;
  assign new_F1962_ = new_F1984_ & ~new_F1985_;
  assign new_F1963_ = ~F1931 & F1932;
  assign new_F1964_ = F1931 & ~F1932;
  assign new_F1965_ = ~new_F1947_ | new_F1957_;
  assign new_F1966_ = new_F1947_ & new_F1957_;
  assign new_F1967_ = ~new_F1947_ & ~new_F1957_;
  assign new_F1968_ = new_F1989_ | new_F1988_;
  assign new_F1969_ = F1935 | new_F1968_;
  assign new_F1970_ = new_F1993_ | new_F1992_;
  assign new_F1971_ = ~F1935 & new_F1970_;
  assign new_F1972_ = new_F1991_ | new_F1990_;
  assign new_F1973_ = F1935 & new_F1972_;
  assign new_F1974_ = F1933 & ~new_F1943_;
  assign new_F1975_ = ~F1933 & new_F1943_;
  assign new_F1976_ = ~F1932 | ~new_F1957_;
  assign new_F1977_ = new_F1943_ & new_F1976_;
  assign new_F1978_ = ~new_F1943_ & ~new_F1977_;
  assign new_F1979_ = new_F1943_ | new_F1976_;
  assign new_F1980_ = ~F1933 & F1934;
  assign new_F1981_ = F1933 & ~F1934;
  assign new_F1982_ = new_F1950_ | new_F1987_;
  assign new_F1983_ = ~new_F1950_ & ~new_F1986_;
  assign new_F1984_ = F1933 | new_F1950_;
  assign new_F1985_ = F1933 | F1934;
  assign new_F1986_ = new_F1950_ & new_F1987_;
  assign new_F1987_ = ~F1932 | ~new_F1957_;
  assign new_F1988_ = new_F1965_ & new_F1985_;
  assign new_F1989_ = ~new_F1965_ & ~new_F1985_;
  assign new_F1990_ = new_F1994_ | new_F1995_;
  assign new_F1991_ = ~F1936 & new_F1950_;
  assign new_F1992_ = new_F1996_ | new_F1997_;
  assign new_F1993_ = F1936 & new_F1950_;
  assign new_F1994_ = ~F1936 & ~new_F1950_;
  assign new_F1995_ = F1936 & ~new_F1950_;
  assign new_F1996_ = F1936 & ~new_F1950_;
  assign new_F1997_ = ~F1936 & new_F1950_;
  assign new_F2004_ = new_F2011_ & new_F2010_;
  assign new_F2005_ = new_F2013_ | new_F2012_;
  assign new_F2006_ = new_F2015_ | new_F2014_;
  assign new_F2007_ = new_F2017_ & new_F2016_;
  assign new_F2008_ = new_F2017_ & new_F2018_;
  assign new_F2009_ = new_F2010_ | new_F2019_;
  assign new_F2010_ = F1999 | new_F2022_;
  assign new_F2011_ = new_F2021_ | new_F2020_;
  assign new_F2012_ = new_F2026_ & new_F2025_;
  assign new_F2013_ = new_F2024_ & new_F2023_;
  assign new_F2014_ = new_F2029_ | new_F2028_;
  assign new_F2015_ = new_F2024_ & new_F2027_;
  assign new_F2016_ = F1999 | new_F2032_;
  assign new_F2017_ = new_F2031_ | new_F2030_;
  assign new_F2018_ = new_F2034_ | new_F2033_;
  assign new_F2019_ = ~new_F2010_ & new_F2036_;
  assign new_F2020_ = ~new_F2012_ & new_F2024_;
  assign new_F2021_ = new_F2012_ & ~new_F2024_;
  assign new_F2022_ = F1998 & ~F1999;
  assign new_F2023_ = ~new_F2045_ | ~new_F2046_;
  assign new_F2024_ = new_F2038_ | new_F2040_;
  assign new_F2025_ = new_F2048_ | new_F2047_;
  assign new_F2026_ = new_F2042_ | new_F2041_;
  assign new_F2027_ = ~new_F2050_ | ~new_F2049_;
  assign new_F2028_ = ~new_F2051_ & new_F2052_;
  assign new_F2029_ = new_F2051_ & ~new_F2052_;
  assign new_F2030_ = ~F1998 & F1999;
  assign new_F2031_ = F1998 & ~F1999;
  assign new_F2032_ = ~new_F2014_ | new_F2024_;
  assign new_F2033_ = new_F2014_ & new_F2024_;
  assign new_F2034_ = ~new_F2014_ & ~new_F2024_;
  assign new_F2035_ = new_F2056_ | new_F2055_;
  assign new_F2036_ = F2002 | new_F2035_;
  assign new_F2037_ = new_F2060_ | new_F2059_;
  assign new_F2038_ = ~F2002 & new_F2037_;
  assign new_F2039_ = new_F2058_ | new_F2057_;
  assign new_F2040_ = F2002 & new_F2039_;
  assign new_F2041_ = F2000 & ~new_F2010_;
  assign new_F2042_ = ~F2000 & new_F2010_;
  assign new_F2043_ = ~F1999 | ~new_F2024_;
  assign new_F2044_ = new_F2010_ & new_F2043_;
  assign new_F2045_ = ~new_F2010_ & ~new_F2044_;
  assign new_F2046_ = new_F2010_ | new_F2043_;
  assign new_F2047_ = ~F2000 & F2001;
  assign new_F2048_ = F2000 & ~F2001;
  assign new_F2049_ = new_F2017_ | new_F2054_;
  assign new_F2050_ = ~new_F2017_ & ~new_F2053_;
  assign new_F2051_ = F2000 | new_F2017_;
  assign new_F2052_ = F2000 | F2001;
  assign new_F2053_ = new_F2017_ & new_F2054_;
  assign new_F2054_ = ~F1999 | ~new_F2024_;
  assign new_F2055_ = new_F2032_ & new_F2052_;
  assign new_F2056_ = ~new_F2032_ & ~new_F2052_;
  assign new_F2057_ = new_F2061_ | new_F2062_;
  assign new_F2058_ = ~F2003 & new_F2017_;
  assign new_F2059_ = new_F2063_ | new_F2064_;
  assign new_F2060_ = F2003 & new_F2017_;
  assign new_F2061_ = ~F2003 & ~new_F2017_;
  assign new_F2062_ = F2003 & ~new_F2017_;
  assign new_F2063_ = F2003 & ~new_F2017_;
  assign new_F2064_ = ~F2003 & new_F2017_;
  assign new_F2071_ = new_F2078_ & new_F2077_;
  assign new_F2072_ = new_F2080_ | new_F2079_;
  assign new_F2073_ = new_F2082_ | new_F2081_;
  assign new_F2074_ = new_F2084_ & new_F2083_;
  assign new_F2075_ = new_F2084_ & new_F2085_;
  assign new_F2076_ = new_F2077_ | new_F2086_;
  assign new_F2077_ = F2066 | new_F2089_;
  assign new_F2078_ = new_F2088_ | new_F2087_;
  assign new_F2079_ = new_F2093_ & new_F2092_;
  assign new_F2080_ = new_F2091_ & new_F2090_;
  assign new_F2081_ = new_F2096_ | new_F2095_;
  assign new_F2082_ = new_F2091_ & new_F2094_;
  assign new_F2083_ = F2066 | new_F2099_;
  assign new_F2084_ = new_F2098_ | new_F2097_;
  assign new_F2085_ = new_F2101_ | new_F2100_;
  assign new_F2086_ = ~new_F2077_ & new_F2103_;
  assign new_F2087_ = ~new_F2079_ & new_F2091_;
  assign new_F2088_ = new_F2079_ & ~new_F2091_;
  assign new_F2089_ = F2065 & ~F2066;
  assign new_F2090_ = ~new_F2112_ | ~new_F2113_;
  assign new_F2091_ = new_F2105_ | new_F2107_;
  assign new_F2092_ = new_F2115_ | new_F2114_;
  assign new_F2093_ = new_F2109_ | new_F2108_;
  assign new_F2094_ = ~new_F2117_ | ~new_F2116_;
  assign new_F2095_ = ~new_F2118_ & new_F2119_;
  assign new_F2096_ = new_F2118_ & ~new_F2119_;
  assign new_F2097_ = ~F2065 & F2066;
  assign new_F2098_ = F2065 & ~F2066;
  assign new_F2099_ = ~new_F2081_ | new_F2091_;
  assign new_F2100_ = new_F2081_ & new_F2091_;
  assign new_F2101_ = ~new_F2081_ & ~new_F2091_;
  assign new_F2102_ = new_F2123_ | new_F2122_;
  assign new_F2103_ = F2069 | new_F2102_;
  assign new_F2104_ = new_F2127_ | new_F2126_;
  assign new_F2105_ = ~F2069 & new_F2104_;
  assign new_F2106_ = new_F2125_ | new_F2124_;
  assign new_F2107_ = F2069 & new_F2106_;
  assign new_F2108_ = F2067 & ~new_F2077_;
  assign new_F2109_ = ~F2067 & new_F2077_;
  assign new_F2110_ = ~F2066 | ~new_F2091_;
  assign new_F2111_ = new_F2077_ & new_F2110_;
  assign new_F2112_ = ~new_F2077_ & ~new_F2111_;
  assign new_F2113_ = new_F2077_ | new_F2110_;
  assign new_F2114_ = ~F2067 & F2068;
  assign new_F2115_ = F2067 & ~F2068;
  assign new_F2116_ = new_F2084_ | new_F2121_;
  assign new_F2117_ = ~new_F2084_ & ~new_F2120_;
  assign new_F2118_ = F2067 | new_F2084_;
  assign new_F2119_ = F2067 | F2068;
  assign new_F2120_ = new_F2084_ & new_F2121_;
  assign new_F2121_ = ~F2066 | ~new_F2091_;
  assign new_F2122_ = new_F2099_ & new_F2119_;
  assign new_F2123_ = ~new_F2099_ & ~new_F2119_;
  assign new_F2124_ = new_F2128_ | new_F2129_;
  assign new_F2125_ = ~F2070 & new_F2084_;
  assign new_F2126_ = new_F2130_ | new_F2131_;
  assign new_F2127_ = F2070 & new_F2084_;
  assign new_F2128_ = ~F2070 & ~new_F2084_;
  assign new_F2129_ = F2070 & ~new_F2084_;
  assign new_F2130_ = F2070 & ~new_F2084_;
  assign new_F2131_ = ~F2070 & new_F2084_;
  assign new_F2138_ = new_F2145_ & new_F2144_;
  assign new_F2139_ = new_F2147_ | new_F2146_;
  assign new_F2140_ = new_F2149_ | new_F2148_;
  assign new_F2141_ = new_F2151_ & new_F2150_;
  assign new_F2142_ = new_F2151_ & new_F2152_;
  assign new_F2143_ = new_F2144_ | new_F2153_;
  assign new_F2144_ = F2133 | new_F2156_;
  assign new_F2145_ = new_F2155_ | new_F2154_;
  assign new_F2146_ = new_F2160_ & new_F2159_;
  assign new_F2147_ = new_F2158_ & new_F2157_;
  assign new_F2148_ = new_F2163_ | new_F2162_;
  assign new_F2149_ = new_F2158_ & new_F2161_;
  assign new_F2150_ = F2133 | new_F2166_;
  assign new_F2151_ = new_F2165_ | new_F2164_;
  assign new_F2152_ = new_F2168_ | new_F2167_;
  assign new_F2153_ = ~new_F2144_ & new_F2170_;
  assign new_F2154_ = ~new_F2146_ & new_F2158_;
  assign new_F2155_ = new_F2146_ & ~new_F2158_;
  assign new_F2156_ = F2132 & ~F2133;
  assign new_F2157_ = ~new_F2179_ | ~new_F2180_;
  assign new_F2158_ = new_F2172_ | new_F2174_;
  assign new_F2159_ = new_F2182_ | new_F2181_;
  assign new_F2160_ = new_F2176_ | new_F2175_;
  assign new_F2161_ = ~new_F2184_ | ~new_F2183_;
  assign new_F2162_ = ~new_F2185_ & new_F2186_;
  assign new_F2163_ = new_F2185_ & ~new_F2186_;
  assign new_F2164_ = ~F2132 & F2133;
  assign new_F2165_ = F2132 & ~F2133;
  assign new_F2166_ = ~new_F2148_ | new_F2158_;
  assign new_F2167_ = new_F2148_ & new_F2158_;
  assign new_F2168_ = ~new_F2148_ & ~new_F2158_;
  assign new_F2169_ = new_F2190_ | new_F2189_;
  assign new_F2170_ = F2136 | new_F2169_;
  assign new_F2171_ = new_F2194_ | new_F2193_;
  assign new_F2172_ = ~F2136 & new_F2171_;
  assign new_F2173_ = new_F2192_ | new_F2191_;
  assign new_F2174_ = F2136 & new_F2173_;
  assign new_F2175_ = F2134 & ~new_F2144_;
  assign new_F2176_ = ~F2134 & new_F2144_;
  assign new_F2177_ = ~F2133 | ~new_F2158_;
  assign new_F2178_ = new_F2144_ & new_F2177_;
  assign new_F2179_ = ~new_F2144_ & ~new_F2178_;
  assign new_F2180_ = new_F2144_ | new_F2177_;
  assign new_F2181_ = ~F2134 & F2135;
  assign new_F2182_ = F2134 & ~F2135;
  assign new_F2183_ = new_F2151_ | new_F2188_;
  assign new_F2184_ = ~new_F2151_ & ~new_F2187_;
  assign new_F2185_ = F2134 | new_F2151_;
  assign new_F2186_ = F2134 | F2135;
  assign new_F2187_ = new_F2151_ & new_F2188_;
  assign new_F2188_ = ~F2133 | ~new_F2158_;
  assign new_F2189_ = new_F2166_ & new_F2186_;
  assign new_F2190_ = ~new_F2166_ & ~new_F2186_;
  assign new_F2191_ = new_F2195_ | new_F2196_;
  assign new_F2192_ = ~F2137 & new_F2151_;
  assign new_F2193_ = new_F2197_ | new_F2198_;
  assign new_F2194_ = F2137 & new_F2151_;
  assign new_F2195_ = ~F2137 & ~new_F2151_;
  assign new_F2196_ = F2137 & ~new_F2151_;
  assign new_F2197_ = F2137 & ~new_F2151_;
  assign new_F2198_ = ~F2137 & new_F2151_;
  assign new_F2205_ = new_F2212_ & new_F2211_;
  assign new_F2206_ = new_F2214_ | new_F2213_;
  assign new_F2207_ = new_F2216_ | new_F2215_;
  assign new_F2208_ = new_F2218_ & new_F2217_;
  assign new_F2209_ = new_F2218_ & new_F2219_;
  assign new_F2210_ = new_F2211_ | new_F2220_;
  assign new_F2211_ = F2200 | new_F2223_;
  assign new_F2212_ = new_F2222_ | new_F2221_;
  assign new_F2213_ = new_F2227_ & new_F2226_;
  assign new_F2214_ = new_F2225_ & new_F2224_;
  assign new_F2215_ = new_F2230_ | new_F2229_;
  assign new_F2216_ = new_F2225_ & new_F2228_;
  assign new_F2217_ = F2200 | new_F2233_;
  assign new_F2218_ = new_F2232_ | new_F2231_;
  assign new_F2219_ = new_F2235_ | new_F2234_;
  assign new_F2220_ = ~new_F2211_ & new_F2237_;
  assign new_F2221_ = ~new_F2213_ & new_F2225_;
  assign new_F2222_ = new_F2213_ & ~new_F2225_;
  assign new_F2223_ = F2199 & ~F2200;
  assign new_F2224_ = ~new_F2246_ | ~new_F2247_;
  assign new_F2225_ = new_F2239_ | new_F2241_;
  assign new_F2226_ = new_F2249_ | new_F2248_;
  assign new_F2227_ = new_F2243_ | new_F2242_;
  assign new_F2228_ = ~new_F2251_ | ~new_F2250_;
  assign new_F2229_ = ~new_F2252_ & new_F2253_;
  assign new_F2230_ = new_F2252_ & ~new_F2253_;
  assign new_F2231_ = ~F2199 & F2200;
  assign new_F2232_ = F2199 & ~F2200;
  assign new_F2233_ = ~new_F2215_ | new_F2225_;
  assign new_F2234_ = new_F2215_ & new_F2225_;
  assign new_F2235_ = ~new_F2215_ & ~new_F2225_;
  assign new_F2236_ = new_F2257_ | new_F2256_;
  assign new_F2237_ = F2203 | new_F2236_;
  assign new_F2238_ = new_F2261_ | new_F2260_;
  assign new_F2239_ = ~F2203 & new_F2238_;
  assign new_F2240_ = new_F2259_ | new_F2258_;
  assign new_F2241_ = F2203 & new_F2240_;
  assign new_F2242_ = F2201 & ~new_F2211_;
  assign new_F2243_ = ~F2201 & new_F2211_;
  assign new_F2244_ = ~F2200 | ~new_F2225_;
  assign new_F2245_ = new_F2211_ & new_F2244_;
  assign new_F2246_ = ~new_F2211_ & ~new_F2245_;
  assign new_F2247_ = new_F2211_ | new_F2244_;
  assign new_F2248_ = ~F2201 & F2202;
  assign new_F2249_ = F2201 & ~F2202;
  assign new_F2250_ = new_F2218_ | new_F2255_;
  assign new_F2251_ = ~new_F2218_ & ~new_F2254_;
  assign new_F2252_ = F2201 | new_F2218_;
  assign new_F2253_ = F2201 | F2202;
  assign new_F2254_ = new_F2218_ & new_F2255_;
  assign new_F2255_ = ~F2200 | ~new_F2225_;
  assign new_F2256_ = new_F2233_ & new_F2253_;
  assign new_F2257_ = ~new_F2233_ & ~new_F2253_;
  assign new_F2258_ = new_F2262_ | new_F2263_;
  assign new_F2259_ = ~F2204 & new_F2218_;
  assign new_F2260_ = new_F2264_ | new_F2265_;
  assign new_F2261_ = F2204 & new_F2218_;
  assign new_F2262_ = ~F2204 & ~new_F2218_;
  assign new_F2263_ = F2204 & ~new_F2218_;
  assign new_F2264_ = F2204 & ~new_F2218_;
  assign new_F2265_ = ~F2204 & new_F2218_;
  assign new_F2272_ = new_F2279_ & new_F2278_;
  assign new_F2273_ = new_F2281_ | new_F2280_;
  assign new_F2274_ = new_F2283_ | new_F2282_;
  assign new_F2275_ = new_F2285_ & new_F2284_;
  assign new_F2276_ = new_F2285_ & new_F2286_;
  assign new_F2277_ = new_F2278_ | new_F2287_;
  assign new_F2278_ = F2267 | new_F2290_;
  assign new_F2279_ = new_F2289_ | new_F2288_;
  assign new_F2280_ = new_F2294_ & new_F2293_;
  assign new_F2281_ = new_F2292_ & new_F2291_;
  assign new_F2282_ = new_F2297_ | new_F2296_;
  assign new_F2283_ = new_F2292_ & new_F2295_;
  assign new_F2284_ = F2267 | new_F2300_;
  assign new_F2285_ = new_F2299_ | new_F2298_;
  assign new_F2286_ = new_F2302_ | new_F2301_;
  assign new_F2287_ = ~new_F2278_ & new_F2304_;
  assign new_F2288_ = ~new_F2280_ & new_F2292_;
  assign new_F2289_ = new_F2280_ & ~new_F2292_;
  assign new_F2290_ = F2266 & ~F2267;
  assign new_F2291_ = ~new_F2313_ | ~new_F2314_;
  assign new_F2292_ = new_F2306_ | new_F2308_;
  assign new_F2293_ = new_F2316_ | new_F2315_;
  assign new_F2294_ = new_F2310_ | new_F2309_;
  assign new_F2295_ = ~new_F2318_ | ~new_F2317_;
  assign new_F2296_ = ~new_F2319_ & new_F2320_;
  assign new_F2297_ = new_F2319_ & ~new_F2320_;
  assign new_F2298_ = ~F2266 & F2267;
  assign new_F2299_ = F2266 & ~F2267;
  assign new_F2300_ = ~new_F2282_ | new_F2292_;
  assign new_F2301_ = new_F2282_ & new_F2292_;
  assign new_F2302_ = ~new_F2282_ & ~new_F2292_;
  assign new_F2303_ = new_F2324_ | new_F2323_;
  assign new_F2304_ = F2270 | new_F2303_;
  assign new_F2305_ = new_F2328_ | new_F2327_;
  assign new_F2306_ = ~F2270 & new_F2305_;
  assign new_F2307_ = new_F2326_ | new_F2325_;
  assign new_F2308_ = F2270 & new_F2307_;
  assign new_F2309_ = F2268 & ~new_F2278_;
  assign new_F2310_ = ~F2268 & new_F2278_;
  assign new_F2311_ = ~F2267 | ~new_F2292_;
  assign new_F2312_ = new_F2278_ & new_F2311_;
  assign new_F2313_ = ~new_F2278_ & ~new_F2312_;
  assign new_F2314_ = new_F2278_ | new_F2311_;
  assign new_F2315_ = ~F2268 & F2269;
  assign new_F2316_ = F2268 & ~F2269;
  assign new_F2317_ = new_F2285_ | new_F2322_;
  assign new_F2318_ = ~new_F2285_ & ~new_F2321_;
  assign new_F2319_ = F2268 | new_F2285_;
  assign new_F2320_ = F2268 | F2269;
  assign new_F2321_ = new_F2285_ & new_F2322_;
  assign new_F2322_ = ~F2267 | ~new_F2292_;
  assign new_F2323_ = new_F2300_ & new_F2320_;
  assign new_F2324_ = ~new_F2300_ & ~new_F2320_;
  assign new_F2325_ = new_F2329_ | new_F2330_;
  assign new_F2326_ = ~F2271 & new_F2285_;
  assign new_F2327_ = new_F2331_ | new_F2332_;
  assign new_F2328_ = F2271 & new_F2285_;
  assign new_F2329_ = ~F2271 & ~new_F2285_;
  assign new_F2330_ = F2271 & ~new_F2285_;
  assign new_F2331_ = F2271 & ~new_F2285_;
  assign new_F2332_ = ~F2271 & new_F2285_;
  assign new_F2339_ = new_F2346_ & new_F2345_;
  assign new_F2340_ = new_F2348_ | new_F2347_;
  assign new_F2341_ = new_F2350_ | new_F2349_;
  assign new_F2342_ = new_F2352_ & new_F2351_;
  assign new_F2343_ = new_F2352_ & new_F2353_;
  assign new_F2344_ = new_F2345_ | new_F2354_;
  assign new_F2345_ = F2334 | new_F2357_;
  assign new_F2346_ = new_F2356_ | new_F2355_;
  assign new_F2347_ = new_F2361_ & new_F2360_;
  assign new_F2348_ = new_F2359_ & new_F2358_;
  assign new_F2349_ = new_F2364_ | new_F2363_;
  assign new_F2350_ = new_F2359_ & new_F2362_;
  assign new_F2351_ = F2334 | new_F2367_;
  assign new_F2352_ = new_F2366_ | new_F2365_;
  assign new_F2353_ = new_F2369_ | new_F2368_;
  assign new_F2354_ = ~new_F2345_ & new_F2371_;
  assign new_F2355_ = ~new_F2347_ & new_F2359_;
  assign new_F2356_ = new_F2347_ & ~new_F2359_;
  assign new_F2357_ = F2333 & ~F2334;
  assign new_F2358_ = ~new_F2380_ | ~new_F2381_;
  assign new_F2359_ = new_F2373_ | new_F2375_;
  assign new_F2360_ = new_F2383_ | new_F2382_;
  assign new_F2361_ = new_F2377_ | new_F2376_;
  assign new_F2362_ = ~new_F2385_ | ~new_F2384_;
  assign new_F2363_ = ~new_F2386_ & new_F2387_;
  assign new_F2364_ = new_F2386_ & ~new_F2387_;
  assign new_F2365_ = ~F2333 & F2334;
  assign new_F2366_ = F2333 & ~F2334;
  assign new_F2367_ = ~new_F2349_ | new_F2359_;
  assign new_F2368_ = new_F2349_ & new_F2359_;
  assign new_F2369_ = ~new_F2349_ & ~new_F2359_;
  assign new_F2370_ = new_F2391_ | new_F2390_;
  assign new_F2371_ = F2337 | new_F2370_;
  assign new_F2372_ = new_F2395_ | new_F2394_;
  assign new_F2373_ = ~F2337 & new_F2372_;
  assign new_F2374_ = new_F2393_ | new_F2392_;
  assign new_F2375_ = F2337 & new_F2374_;
  assign new_F2376_ = F2335 & ~new_F2345_;
  assign new_F2377_ = ~F2335 & new_F2345_;
  assign new_F2378_ = ~F2334 | ~new_F2359_;
  assign new_F2379_ = new_F2345_ & new_F2378_;
  assign new_F2380_ = ~new_F2345_ & ~new_F2379_;
  assign new_F2381_ = new_F2345_ | new_F2378_;
  assign new_F2382_ = ~F2335 & F2336;
  assign new_F2383_ = F2335 & ~F2336;
  assign new_F2384_ = new_F2352_ | new_F2389_;
  assign new_F2385_ = ~new_F2352_ & ~new_F2388_;
  assign new_F2386_ = F2335 | new_F2352_;
  assign new_F2387_ = F2335 | F2336;
  assign new_F2388_ = new_F2352_ & new_F2389_;
  assign new_F2389_ = ~F2334 | ~new_F2359_;
  assign new_F2390_ = new_F2367_ & new_F2387_;
  assign new_F2391_ = ~new_F2367_ & ~new_F2387_;
  assign new_F2392_ = new_F2396_ | new_F2397_;
  assign new_F2393_ = ~F2338 & new_F2352_;
  assign new_F2394_ = new_F2398_ | new_F2399_;
  assign new_F2395_ = F2338 & new_F2352_;
  assign new_F2396_ = ~F2338 & ~new_F2352_;
  assign new_F2397_ = F2338 & ~new_F2352_;
  assign new_F2398_ = F2338 & ~new_F2352_;
  assign new_F2399_ = ~F2338 & new_F2352_;
  assign new_F2406_ = new_F2413_ & new_F2412_;
  assign new_F2407_ = new_F2415_ | new_F2414_;
  assign new_F2408_ = new_F2417_ | new_F2416_;
  assign new_F2409_ = new_F2419_ & new_F2418_;
  assign new_F2410_ = new_F2419_ & new_F2420_;
  assign new_F2411_ = new_F2412_ | new_F2421_;
  assign new_F2412_ = F2401 | new_F2424_;
  assign new_F2413_ = new_F2423_ | new_F2422_;
  assign new_F2414_ = new_F2428_ & new_F2427_;
  assign new_F2415_ = new_F2426_ & new_F2425_;
  assign new_F2416_ = new_F2431_ | new_F2430_;
  assign new_F2417_ = new_F2426_ & new_F2429_;
  assign new_F2418_ = F2401 | new_F2434_;
  assign new_F2419_ = new_F2433_ | new_F2432_;
  assign new_F2420_ = new_F2436_ | new_F2435_;
  assign new_F2421_ = ~new_F2412_ & new_F2438_;
  assign new_F2422_ = ~new_F2414_ & new_F2426_;
  assign new_F2423_ = new_F2414_ & ~new_F2426_;
  assign new_F2424_ = F2400 & ~F2401;
  assign new_F2425_ = ~new_F2447_ | ~new_F2448_;
  assign new_F2426_ = new_F2440_ | new_F2442_;
  assign new_F2427_ = new_F2450_ | new_F2449_;
  assign new_F2428_ = new_F2444_ | new_F2443_;
  assign new_F2429_ = ~new_F2452_ | ~new_F2451_;
  assign new_F2430_ = ~new_F2453_ & new_F2454_;
  assign new_F2431_ = new_F2453_ & ~new_F2454_;
  assign new_F2432_ = ~F2400 & F2401;
  assign new_F2433_ = F2400 & ~F2401;
  assign new_F2434_ = ~new_F2416_ | new_F2426_;
  assign new_F2435_ = new_F2416_ & new_F2426_;
  assign new_F2436_ = ~new_F2416_ & ~new_F2426_;
  assign new_F2437_ = new_F2458_ | new_F2457_;
  assign new_F2438_ = F2404 | new_F2437_;
  assign new_F2439_ = new_F2462_ | new_F2461_;
  assign new_F2440_ = ~F2404 & new_F2439_;
  assign new_F2441_ = new_F2460_ | new_F2459_;
  assign new_F2442_ = F2404 & new_F2441_;
  assign new_F2443_ = F2402 & ~new_F2412_;
  assign new_F2444_ = ~F2402 & new_F2412_;
  assign new_F2445_ = ~F2401 | ~new_F2426_;
  assign new_F2446_ = new_F2412_ & new_F2445_;
  assign new_F2447_ = ~new_F2412_ & ~new_F2446_;
  assign new_F2448_ = new_F2412_ | new_F2445_;
  assign new_F2449_ = ~F2402 & F2403;
  assign new_F2450_ = F2402 & ~F2403;
  assign new_F2451_ = new_F2419_ | new_F2456_;
  assign new_F2452_ = ~new_F2419_ & ~new_F2455_;
  assign new_F2453_ = F2402 | new_F2419_;
  assign new_F2454_ = F2402 | F2403;
  assign new_F2455_ = new_F2419_ & new_F2456_;
  assign new_F2456_ = ~F2401 | ~new_F2426_;
  assign new_F2457_ = new_F2434_ & new_F2454_;
  assign new_F2458_ = ~new_F2434_ & ~new_F2454_;
  assign new_F2459_ = new_F2463_ | new_F2464_;
  assign new_F2460_ = ~F2405 & new_F2419_;
  assign new_F2461_ = new_F2465_ | new_F2466_;
  assign new_F2462_ = F2405 & new_F2419_;
  assign new_F2463_ = ~F2405 & ~new_F2419_;
  assign new_F2464_ = F2405 & ~new_F2419_;
  assign new_F2465_ = F2405 & ~new_F2419_;
  assign new_F2466_ = ~F2405 & new_F2419_;
  assign new_F2473_ = new_F2480_ & new_F2479_;
  assign new_F2474_ = new_F2482_ | new_F2481_;
  assign new_F2475_ = new_F2484_ | new_F2483_;
  assign new_F2476_ = new_F2486_ & new_F2485_;
  assign new_F2477_ = new_F2486_ & new_F2487_;
  assign new_F2478_ = new_F2479_ | new_F2488_;
  assign new_F2479_ = F2468 | new_F2491_;
  assign new_F2480_ = new_F2490_ | new_F2489_;
  assign new_F2481_ = new_F2495_ & new_F2494_;
  assign new_F2482_ = new_F2493_ & new_F2492_;
  assign new_F2483_ = new_F2498_ | new_F2497_;
  assign new_F2484_ = new_F2493_ & new_F2496_;
  assign new_F2485_ = F2468 | new_F2501_;
  assign new_F2486_ = new_F2500_ | new_F2499_;
  assign new_F2487_ = new_F2503_ | new_F2502_;
  assign new_F2488_ = ~new_F2479_ & new_F2505_;
  assign new_F2489_ = ~new_F2481_ & new_F2493_;
  assign new_F2490_ = new_F2481_ & ~new_F2493_;
  assign new_F2491_ = F2467 & ~F2468;
  assign new_F2492_ = ~new_F2514_ | ~new_F2515_;
  assign new_F2493_ = new_F2507_ | new_F2509_;
  assign new_F2494_ = new_F2517_ | new_F2516_;
  assign new_F2495_ = new_F2511_ | new_F2510_;
  assign new_F2496_ = ~new_F2519_ | ~new_F2518_;
  assign new_F2497_ = ~new_F2520_ & new_F2521_;
  assign new_F2498_ = new_F2520_ & ~new_F2521_;
  assign new_F2499_ = ~F2467 & F2468;
  assign new_F2500_ = F2467 & ~F2468;
  assign new_F2501_ = ~new_F2483_ | new_F2493_;
  assign new_F2502_ = new_F2483_ & new_F2493_;
  assign new_F2503_ = ~new_F2483_ & ~new_F2493_;
  assign new_F2504_ = new_F2525_ | new_F2524_;
  assign new_F2505_ = F2471 | new_F2504_;
  assign new_F2506_ = new_F2529_ | new_F2528_;
  assign new_F2507_ = ~F2471 & new_F2506_;
  assign new_F2508_ = new_F2527_ | new_F2526_;
  assign new_F2509_ = F2471 & new_F2508_;
  assign new_F2510_ = F2469 & ~new_F2479_;
  assign new_F2511_ = ~F2469 & new_F2479_;
  assign new_F2512_ = ~F2468 | ~new_F2493_;
  assign new_F2513_ = new_F2479_ & new_F2512_;
  assign new_F2514_ = ~new_F2479_ & ~new_F2513_;
  assign new_F2515_ = new_F2479_ | new_F2512_;
  assign new_F2516_ = ~F2469 & F2470;
  assign new_F2517_ = F2469 & ~F2470;
  assign new_F2518_ = new_F2486_ | new_F2523_;
  assign new_F2519_ = ~new_F2486_ & ~new_F2522_;
  assign new_F2520_ = F2469 | new_F2486_;
  assign new_F2521_ = F2469 | F2470;
  assign new_F2522_ = new_F2486_ & new_F2523_;
  assign new_F2523_ = ~F2468 | ~new_F2493_;
  assign new_F2524_ = new_F2501_ & new_F2521_;
  assign new_F2525_ = ~new_F2501_ & ~new_F2521_;
  assign new_F2526_ = new_F2530_ | new_F2531_;
  assign new_F2527_ = ~F2472 & new_F2486_;
  assign new_F2528_ = new_F2532_ | new_F2533_;
  assign new_F2529_ = F2472 & new_F2486_;
  assign new_F2530_ = ~F2472 & ~new_F2486_;
  assign new_F2531_ = F2472 & ~new_F2486_;
  assign new_F2532_ = F2472 & ~new_F2486_;
  assign new_F2533_ = ~F2472 & new_F2486_;
  assign new_F2540_ = new_F2547_ & new_F2546_;
  assign new_F2541_ = new_F2549_ | new_F2548_;
  assign new_F2542_ = new_F2551_ | new_F2550_;
  assign new_F2543_ = new_F2553_ & new_F2552_;
  assign new_F2544_ = new_F2553_ & new_F2554_;
  assign new_F2545_ = new_F2546_ | new_F2555_;
  assign new_F2546_ = F2535 | new_F2558_;
  assign new_F2547_ = new_F2557_ | new_F2556_;
  assign new_F2548_ = new_F2562_ & new_F2561_;
  assign new_F2549_ = new_F2560_ & new_F2559_;
  assign new_F2550_ = new_F2565_ | new_F2564_;
  assign new_F2551_ = new_F2560_ & new_F2563_;
  assign new_F2552_ = F2535 | new_F2568_;
  assign new_F2553_ = new_F2567_ | new_F2566_;
  assign new_F2554_ = new_F2570_ | new_F2569_;
  assign new_F2555_ = ~new_F2546_ & new_F2572_;
  assign new_F2556_ = ~new_F2548_ & new_F2560_;
  assign new_F2557_ = new_F2548_ & ~new_F2560_;
  assign new_F2558_ = F2534 & ~F2535;
  assign new_F2559_ = ~new_F2581_ | ~new_F2582_;
  assign new_F2560_ = new_F2574_ | new_F2576_;
  assign new_F2561_ = new_F2584_ | new_F2583_;
  assign new_F2562_ = new_F2578_ | new_F2577_;
  assign new_F2563_ = ~new_F2586_ | ~new_F2585_;
  assign new_F2564_ = ~new_F2587_ & new_F2588_;
  assign new_F2565_ = new_F2587_ & ~new_F2588_;
  assign new_F2566_ = ~F2534 & F2535;
  assign new_F2567_ = F2534 & ~F2535;
  assign new_F2568_ = ~new_F2550_ | new_F2560_;
  assign new_F2569_ = new_F2550_ & new_F2560_;
  assign new_F2570_ = ~new_F2550_ & ~new_F2560_;
  assign new_F2571_ = new_F2592_ | new_F2591_;
  assign new_F2572_ = F2538 | new_F2571_;
  assign new_F2573_ = new_F2596_ | new_F2595_;
  assign new_F2574_ = ~F2538 & new_F2573_;
  assign new_F2575_ = new_F2594_ | new_F2593_;
  assign new_F2576_ = F2538 & new_F2575_;
  assign new_F2577_ = F2536 & ~new_F2546_;
  assign new_F2578_ = ~F2536 & new_F2546_;
  assign new_F2579_ = ~F2535 | ~new_F2560_;
  assign new_F2580_ = new_F2546_ & new_F2579_;
  assign new_F2581_ = ~new_F2546_ & ~new_F2580_;
  assign new_F2582_ = new_F2546_ | new_F2579_;
  assign new_F2583_ = ~F2536 & F2537;
  assign new_F2584_ = F2536 & ~F2537;
  assign new_F2585_ = new_F2553_ | new_F2590_;
  assign new_F2586_ = ~new_F2553_ & ~new_F2589_;
  assign new_F2587_ = F2536 | new_F2553_;
  assign new_F2588_ = F2536 | F2537;
  assign new_F2589_ = new_F2553_ & new_F2590_;
  assign new_F2590_ = ~F2535 | ~new_F2560_;
  assign new_F2591_ = new_F2568_ & new_F2588_;
  assign new_F2592_ = ~new_F2568_ & ~new_F2588_;
  assign new_F2593_ = new_F2597_ | new_F2598_;
  assign new_F2594_ = ~F2539 & new_F2553_;
  assign new_F2595_ = new_F2599_ | new_F2600_;
  assign new_F2596_ = F2539 & new_F2553_;
  assign new_F2597_ = ~F2539 & ~new_F2553_;
  assign new_F2598_ = F2539 & ~new_F2553_;
  assign new_F2599_ = F2539 & ~new_F2553_;
  assign new_F2600_ = ~F2539 & new_F2553_;
  assign new_F2607_ = new_F2614_ & new_F2613_;
  assign new_F2608_ = new_F2616_ | new_F2615_;
  assign new_F2609_ = new_F2618_ | new_F2617_;
  assign new_F2610_ = new_F2620_ & new_F2619_;
  assign new_F2611_ = new_F2620_ & new_F2621_;
  assign new_F2612_ = new_F2613_ | new_F2622_;
  assign new_F2613_ = F2602 | new_F2625_;
  assign new_F2614_ = new_F2624_ | new_F2623_;
  assign new_F2615_ = new_F2629_ & new_F2628_;
  assign new_F2616_ = new_F2627_ & new_F2626_;
  assign new_F2617_ = new_F2632_ | new_F2631_;
  assign new_F2618_ = new_F2627_ & new_F2630_;
  assign new_F2619_ = F2602 | new_F2635_;
  assign new_F2620_ = new_F2634_ | new_F2633_;
  assign new_F2621_ = new_F2637_ | new_F2636_;
  assign new_F2622_ = ~new_F2613_ & new_F2639_;
  assign new_F2623_ = ~new_F2615_ & new_F2627_;
  assign new_F2624_ = new_F2615_ & ~new_F2627_;
  assign new_F2625_ = F2601 & ~F2602;
  assign new_F2626_ = ~new_F2648_ | ~new_F2649_;
  assign new_F2627_ = new_F2641_ | new_F2643_;
  assign new_F2628_ = new_F2651_ | new_F2650_;
  assign new_F2629_ = new_F2645_ | new_F2644_;
  assign new_F2630_ = ~new_F2653_ | ~new_F2652_;
  assign new_F2631_ = ~new_F2654_ & new_F2655_;
  assign new_F2632_ = new_F2654_ & ~new_F2655_;
  assign new_F2633_ = ~F2601 & F2602;
  assign new_F2634_ = F2601 & ~F2602;
  assign new_F2635_ = ~new_F2617_ | new_F2627_;
  assign new_F2636_ = new_F2617_ & new_F2627_;
  assign new_F2637_ = ~new_F2617_ & ~new_F2627_;
  assign new_F2638_ = new_F2659_ | new_F2658_;
  assign new_F2639_ = F2605 | new_F2638_;
  assign new_F2640_ = new_F2663_ | new_F2662_;
  assign new_F2641_ = ~F2605 & new_F2640_;
  assign new_F2642_ = new_F2661_ | new_F2660_;
  assign new_F2643_ = F2605 & new_F2642_;
  assign new_F2644_ = F2603 & ~new_F2613_;
  assign new_F2645_ = ~F2603 & new_F2613_;
  assign new_F2646_ = ~F2602 | ~new_F2627_;
  assign new_F2647_ = new_F2613_ & new_F2646_;
  assign new_F2648_ = ~new_F2613_ & ~new_F2647_;
  assign new_F2649_ = new_F2613_ | new_F2646_;
  assign new_F2650_ = ~F2603 & F2604;
  assign new_F2651_ = F2603 & ~F2604;
  assign new_F2652_ = new_F2620_ | new_F2657_;
  assign new_F2653_ = ~new_F2620_ & ~new_F2656_;
  assign new_F2654_ = F2603 | new_F2620_;
  assign new_F2655_ = F2603 | F2604;
  assign new_F2656_ = new_F2620_ & new_F2657_;
  assign new_F2657_ = ~F2602 | ~new_F2627_;
  assign new_F2658_ = new_F2635_ & new_F2655_;
  assign new_F2659_ = ~new_F2635_ & ~new_F2655_;
  assign new_F2660_ = new_F2664_ | new_F2665_;
  assign new_F2661_ = ~F2606 & new_F2620_;
  assign new_F2662_ = new_F2666_ | new_F2667_;
  assign new_F2663_ = F2606 & new_F2620_;
  assign new_F2664_ = ~F2606 & ~new_F2620_;
  assign new_F2665_ = F2606 & ~new_F2620_;
  assign new_F2666_ = F2606 & ~new_F2620_;
  assign new_F2667_ = ~F2606 & new_F2620_;
  assign new_F2674_ = new_F2681_ & new_F2680_;
  assign new_F2675_ = new_F2683_ | new_F2682_;
  assign new_F2676_ = new_F2685_ | new_F2684_;
  assign new_F2677_ = new_F2687_ & new_F2686_;
  assign new_F2678_ = new_F2687_ & new_F2688_;
  assign new_F2679_ = new_F2680_ | new_F2689_;
  assign new_F2680_ = F2669 | new_F2692_;
  assign new_F2681_ = new_F2691_ | new_F2690_;
  assign new_F2682_ = new_F2696_ & new_F2695_;
  assign new_F2683_ = new_F2694_ & new_F2693_;
  assign new_F2684_ = new_F2699_ | new_F2698_;
  assign new_F2685_ = new_F2694_ & new_F2697_;
  assign new_F2686_ = F2669 | new_F2702_;
  assign new_F2687_ = new_F2701_ | new_F2700_;
  assign new_F2688_ = new_F2704_ | new_F2703_;
  assign new_F2689_ = ~new_F2680_ & new_F2706_;
  assign new_F2690_ = ~new_F2682_ & new_F2694_;
  assign new_F2691_ = new_F2682_ & ~new_F2694_;
  assign new_F2692_ = F2668 & ~F2669;
  assign new_F2693_ = ~new_F2715_ | ~new_F2716_;
  assign new_F2694_ = new_F2708_ | new_F2710_;
  assign new_F2695_ = new_F2718_ | new_F2717_;
  assign new_F2696_ = new_F2712_ | new_F2711_;
  assign new_F2697_ = ~new_F2720_ | ~new_F2719_;
  assign new_F2698_ = ~new_F2721_ & new_F2722_;
  assign new_F2699_ = new_F2721_ & ~new_F2722_;
  assign new_F2700_ = ~F2668 & F2669;
  assign new_F2701_ = F2668 & ~F2669;
  assign new_F2702_ = ~new_F2684_ | new_F2694_;
  assign new_F2703_ = new_F2684_ & new_F2694_;
  assign new_F2704_ = ~new_F2684_ & ~new_F2694_;
  assign new_F2705_ = new_F2726_ | new_F2725_;
  assign new_F2706_ = F2672 | new_F2705_;
  assign new_F2707_ = new_F2730_ | new_F2729_;
  assign new_F2708_ = ~F2672 & new_F2707_;
  assign new_F2709_ = new_F2728_ | new_F2727_;
  assign new_F2710_ = F2672 & new_F2709_;
  assign new_F2711_ = F2670 & ~new_F2680_;
  assign new_F2712_ = ~F2670 & new_F2680_;
  assign new_F2713_ = ~F2669 | ~new_F2694_;
  assign new_F2714_ = new_F2680_ & new_F2713_;
  assign new_F2715_ = ~new_F2680_ & ~new_F2714_;
  assign new_F2716_ = new_F2680_ | new_F2713_;
  assign new_F2717_ = ~F2670 & F2671;
  assign new_F2718_ = F2670 & ~F2671;
  assign new_F2719_ = new_F2687_ | new_F2724_;
  assign new_F2720_ = ~new_F2687_ & ~new_F2723_;
  assign new_F2721_ = F2670 | new_F2687_;
  assign new_F2722_ = F2670 | F2671;
  assign new_F2723_ = new_F2687_ & new_F2724_;
  assign new_F2724_ = ~F2669 | ~new_F2694_;
  assign new_F2725_ = new_F2702_ & new_F2722_;
  assign new_F2726_ = ~new_F2702_ & ~new_F2722_;
  assign new_F2727_ = new_F2731_ | new_F2732_;
  assign new_F2728_ = ~F2673 & new_F2687_;
  assign new_F2729_ = new_F2733_ | new_F2734_;
  assign new_F2730_ = F2673 & new_F2687_;
  assign new_F2731_ = ~F2673 & ~new_F2687_;
  assign new_F2732_ = F2673 & ~new_F2687_;
  assign new_F2733_ = F2673 & ~new_F2687_;
  assign new_F2734_ = ~F2673 & new_F2687_;
  assign new_F2741_ = new_F2748_ & new_F2747_;
  assign new_F2742_ = new_F2750_ | new_F2749_;
  assign new_F2743_ = new_F2752_ | new_F2751_;
  assign new_F2744_ = new_F2754_ & new_F2753_;
  assign new_F2745_ = new_F2754_ & new_F2755_;
  assign new_F2746_ = new_F2747_ | new_F2756_;
  assign new_F2747_ = F2736 | new_F2759_;
  assign new_F2748_ = new_F2758_ | new_F2757_;
  assign new_F2749_ = new_F2763_ & new_F2762_;
  assign new_F2750_ = new_F2761_ & new_F2760_;
  assign new_F2751_ = new_F2766_ | new_F2765_;
  assign new_F2752_ = new_F2761_ & new_F2764_;
  assign new_F2753_ = F2736 | new_F2769_;
  assign new_F2754_ = new_F2768_ | new_F2767_;
  assign new_F2755_ = new_F2771_ | new_F2770_;
  assign new_F2756_ = ~new_F2747_ & new_F2773_;
  assign new_F2757_ = ~new_F2749_ & new_F2761_;
  assign new_F2758_ = new_F2749_ & ~new_F2761_;
  assign new_F2759_ = F2735 & ~F2736;
  assign new_F2760_ = ~new_F2782_ | ~new_F2783_;
  assign new_F2761_ = new_F2775_ | new_F2777_;
  assign new_F2762_ = new_F2785_ | new_F2784_;
  assign new_F2763_ = new_F2779_ | new_F2778_;
  assign new_F2764_ = ~new_F2787_ | ~new_F2786_;
  assign new_F2765_ = ~new_F2788_ & new_F2789_;
  assign new_F2766_ = new_F2788_ & ~new_F2789_;
  assign new_F2767_ = ~F2735 & F2736;
  assign new_F2768_ = F2735 & ~F2736;
  assign new_F2769_ = ~new_F2751_ | new_F2761_;
  assign new_F2770_ = new_F2751_ & new_F2761_;
  assign new_F2771_ = ~new_F2751_ & ~new_F2761_;
  assign new_F2772_ = new_F2793_ | new_F2792_;
  assign new_F2773_ = F2739 | new_F2772_;
  assign new_F2774_ = new_F2797_ | new_F2796_;
  assign new_F2775_ = ~F2739 & new_F2774_;
  assign new_F2776_ = new_F2795_ | new_F2794_;
  assign new_F2777_ = F2739 & new_F2776_;
  assign new_F2778_ = F2737 & ~new_F2747_;
  assign new_F2779_ = ~F2737 & new_F2747_;
  assign new_F2780_ = ~F2736 | ~new_F2761_;
  assign new_F2781_ = new_F2747_ & new_F2780_;
  assign new_F2782_ = ~new_F2747_ & ~new_F2781_;
  assign new_F2783_ = new_F2747_ | new_F2780_;
  assign new_F2784_ = ~F2737 & F2738;
  assign new_F2785_ = F2737 & ~F2738;
  assign new_F2786_ = new_F2754_ | new_F2791_;
  assign new_F2787_ = ~new_F2754_ & ~new_F2790_;
  assign new_F2788_ = F2737 | new_F2754_;
  assign new_F2789_ = F2737 | F2738;
  assign new_F2790_ = new_F2754_ & new_F2791_;
  assign new_F2791_ = ~F2736 | ~new_F2761_;
  assign new_F2792_ = new_F2769_ & new_F2789_;
  assign new_F2793_ = ~new_F2769_ & ~new_F2789_;
  assign new_F2794_ = new_F2798_ | new_F2799_;
  assign new_F2795_ = ~F2740 & new_F2754_;
  assign new_F2796_ = new_F2800_ | new_F2801_;
  assign new_F2797_ = F2740 & new_F2754_;
  assign new_F2798_ = ~F2740 & ~new_F2754_;
  assign new_F2799_ = F2740 & ~new_F2754_;
  assign new_F2800_ = F2740 & ~new_F2754_;
  assign new_F2801_ = ~F2740 & new_F2754_;
  assign new_F2808_ = new_F2815_ & new_F2814_;
  assign new_F2809_ = new_F2817_ | new_F2816_;
  assign new_F2810_ = new_F2819_ | new_F2818_;
  assign new_F2811_ = new_F2821_ & new_F2820_;
  assign new_F2812_ = new_F2821_ & new_F2822_;
  assign new_F2813_ = new_F2814_ | new_F2823_;
  assign new_F2814_ = F2803 | new_F2826_;
  assign new_F2815_ = new_F2825_ | new_F2824_;
  assign new_F2816_ = new_F2830_ & new_F2829_;
  assign new_F2817_ = new_F2828_ & new_F2827_;
  assign new_F2818_ = new_F2833_ | new_F2832_;
  assign new_F2819_ = new_F2828_ & new_F2831_;
  assign new_F2820_ = F2803 | new_F2836_;
  assign new_F2821_ = new_F2835_ | new_F2834_;
  assign new_F2822_ = new_F2838_ | new_F2837_;
  assign new_F2823_ = ~new_F2814_ & new_F2840_;
  assign new_F2824_ = ~new_F2816_ & new_F2828_;
  assign new_F2825_ = new_F2816_ & ~new_F2828_;
  assign new_F2826_ = F2802 & ~F2803;
  assign new_F2827_ = ~new_F2849_ | ~new_F2850_;
  assign new_F2828_ = new_F2842_ | new_F2844_;
  assign new_F2829_ = new_F2852_ | new_F2851_;
  assign new_F2830_ = new_F2846_ | new_F2845_;
  assign new_F2831_ = ~new_F2854_ | ~new_F2853_;
  assign new_F2832_ = ~new_F2855_ & new_F2856_;
  assign new_F2833_ = new_F2855_ & ~new_F2856_;
  assign new_F2834_ = ~F2802 & F2803;
  assign new_F2835_ = F2802 & ~F2803;
  assign new_F2836_ = ~new_F2818_ | new_F2828_;
  assign new_F2837_ = new_F2818_ & new_F2828_;
  assign new_F2838_ = ~new_F2818_ & ~new_F2828_;
  assign new_F2839_ = new_F2860_ | new_F2859_;
  assign new_F2840_ = F2806 | new_F2839_;
  assign new_F2841_ = new_F2864_ | new_F2863_;
  assign new_F2842_ = ~F2806 & new_F2841_;
  assign new_F2843_ = new_F2862_ | new_F2861_;
  assign new_F2844_ = F2806 & new_F2843_;
  assign new_F2845_ = F2804 & ~new_F2814_;
  assign new_F2846_ = ~F2804 & new_F2814_;
  assign new_F2847_ = ~F2803 | ~new_F2828_;
  assign new_F2848_ = new_F2814_ & new_F2847_;
  assign new_F2849_ = ~new_F2814_ & ~new_F2848_;
  assign new_F2850_ = new_F2814_ | new_F2847_;
  assign new_F2851_ = ~F2804 & F2805;
  assign new_F2852_ = F2804 & ~F2805;
  assign new_F2853_ = new_F2821_ | new_F2858_;
  assign new_F2854_ = ~new_F2821_ & ~new_F2857_;
  assign new_F2855_ = F2804 | new_F2821_;
  assign new_F2856_ = F2804 | F2805;
  assign new_F2857_ = new_F2821_ & new_F2858_;
  assign new_F2858_ = ~F2803 | ~new_F2828_;
  assign new_F2859_ = new_F2836_ & new_F2856_;
  assign new_F2860_ = ~new_F2836_ & ~new_F2856_;
  assign new_F2861_ = new_F2865_ | new_F2866_;
  assign new_F2862_ = ~F2807 & new_F2821_;
  assign new_F2863_ = new_F2867_ | new_F2868_;
  assign new_F2864_ = F2807 & new_F2821_;
  assign new_F2865_ = ~F2807 & ~new_F2821_;
  assign new_F2866_ = F2807 & ~new_F2821_;
  assign new_F2867_ = F2807 & ~new_F2821_;
  assign new_F2868_ = ~F2807 & new_F2821_;
  assign new_F2875_ = new_F2882_ & new_F2881_;
  assign new_F2876_ = new_F2884_ | new_F2883_;
  assign new_F2877_ = new_F2886_ | new_F2885_;
  assign new_F2878_ = new_F2888_ & new_F2887_;
  assign new_F2879_ = new_F2888_ & new_F2889_;
  assign new_F2880_ = new_F2881_ | new_F2890_;
  assign new_F2881_ = F2870 | new_F2893_;
  assign new_F2882_ = new_F2892_ | new_F2891_;
  assign new_F2883_ = new_F2897_ & new_F2896_;
  assign new_F2884_ = new_F2895_ & new_F2894_;
  assign new_F2885_ = new_F2900_ | new_F2899_;
  assign new_F2886_ = new_F2895_ & new_F2898_;
  assign new_F2887_ = F2870 | new_F2903_;
  assign new_F2888_ = new_F2902_ | new_F2901_;
  assign new_F2889_ = new_F2905_ | new_F2904_;
  assign new_F2890_ = ~new_F2881_ & new_F2907_;
  assign new_F2891_ = ~new_F2883_ & new_F2895_;
  assign new_F2892_ = new_F2883_ & ~new_F2895_;
  assign new_F2893_ = F2869 & ~F2870;
  assign new_F2894_ = ~new_F2916_ | ~new_F2917_;
  assign new_F2895_ = new_F2909_ | new_F2911_;
  assign new_F2896_ = new_F2919_ | new_F2918_;
  assign new_F2897_ = new_F2913_ | new_F2912_;
  assign new_F2898_ = ~new_F2921_ | ~new_F2920_;
  assign new_F2899_ = ~new_F2922_ & new_F2923_;
  assign new_F2900_ = new_F2922_ & ~new_F2923_;
  assign new_F2901_ = ~F2869 & F2870;
  assign new_F2902_ = F2869 & ~F2870;
  assign new_F2903_ = ~new_F2885_ | new_F2895_;
  assign new_F2904_ = new_F2885_ & new_F2895_;
  assign new_F2905_ = ~new_F2885_ & ~new_F2895_;
  assign new_F2906_ = new_F2927_ | new_F2926_;
  assign new_F2907_ = F2873 | new_F2906_;
  assign new_F2908_ = new_F2931_ | new_F2930_;
  assign new_F2909_ = ~F2873 & new_F2908_;
  assign new_F2910_ = new_F2929_ | new_F2928_;
  assign new_F2911_ = F2873 & new_F2910_;
  assign new_F2912_ = F2871 & ~new_F2881_;
  assign new_F2913_ = ~F2871 & new_F2881_;
  assign new_F2914_ = ~F2870 | ~new_F2895_;
  assign new_F2915_ = new_F2881_ & new_F2914_;
  assign new_F2916_ = ~new_F2881_ & ~new_F2915_;
  assign new_F2917_ = new_F2881_ | new_F2914_;
  assign new_F2918_ = ~F2871 & F2872;
  assign new_F2919_ = F2871 & ~F2872;
  assign new_F2920_ = new_F2888_ | new_F2925_;
  assign new_F2921_ = ~new_F2888_ & ~new_F2924_;
  assign new_F2922_ = F2871 | new_F2888_;
  assign new_F2923_ = F2871 | F2872;
  assign new_F2924_ = new_F2888_ & new_F2925_;
  assign new_F2925_ = ~F2870 | ~new_F2895_;
  assign new_F2926_ = new_F2903_ & new_F2923_;
  assign new_F2927_ = ~new_F2903_ & ~new_F2923_;
  assign new_F2928_ = new_F2932_ | new_F2933_;
  assign new_F2929_ = ~F2874 & new_F2888_;
  assign new_F2930_ = new_F2934_ | new_F2935_;
  assign new_F2931_ = F2874 & new_F2888_;
  assign new_F2932_ = ~F2874 & ~new_F2888_;
  assign new_F2933_ = F2874 & ~new_F2888_;
  assign new_F2934_ = F2874 & ~new_F2888_;
  assign new_F2935_ = ~F2874 & new_F2888_;
  assign new_F2942_ = new_F2949_ & new_F2948_;
  assign new_F2943_ = new_F2951_ | new_F2950_;
  assign new_F2944_ = new_F2953_ | new_F2952_;
  assign new_F2945_ = new_F2955_ & new_F2954_;
  assign new_F2946_ = new_F2955_ & new_F2956_;
  assign new_F2947_ = new_F2948_ | new_F2957_;
  assign new_F2948_ = F2937 | new_F2960_;
  assign new_F2949_ = new_F2959_ | new_F2958_;
  assign new_F2950_ = new_F2964_ & new_F2963_;
  assign new_F2951_ = new_F2962_ & new_F2961_;
  assign new_F2952_ = new_F2967_ | new_F2966_;
  assign new_F2953_ = new_F2962_ & new_F2965_;
  assign new_F2954_ = F2937 | new_F2970_;
  assign new_F2955_ = new_F2969_ | new_F2968_;
  assign new_F2956_ = new_F2972_ | new_F2971_;
  assign new_F2957_ = ~new_F2948_ & new_F2974_;
  assign new_F2958_ = ~new_F2950_ & new_F2962_;
  assign new_F2959_ = new_F2950_ & ~new_F2962_;
  assign new_F2960_ = F2936 & ~F2937;
  assign new_F2961_ = ~new_F2983_ | ~new_F2984_;
  assign new_F2962_ = new_F2976_ | new_F2978_;
  assign new_F2963_ = new_F2986_ | new_F2985_;
  assign new_F2964_ = new_F2980_ | new_F2979_;
  assign new_F2965_ = ~new_F2988_ | ~new_F2987_;
  assign new_F2966_ = ~new_F2989_ & new_F2990_;
  assign new_F2967_ = new_F2989_ & ~new_F2990_;
  assign new_F2968_ = ~F2936 & F2937;
  assign new_F2969_ = F2936 & ~F2937;
  assign new_F2970_ = ~new_F2952_ | new_F2962_;
  assign new_F2971_ = new_F2952_ & new_F2962_;
  assign new_F2972_ = ~new_F2952_ & ~new_F2962_;
  assign new_F2973_ = new_F2994_ | new_F2993_;
  assign new_F2974_ = F2940 | new_F2973_;
  assign new_F2975_ = new_F2998_ | new_F2997_;
  assign new_F2976_ = ~F2940 & new_F2975_;
  assign new_F2977_ = new_F2996_ | new_F2995_;
  assign new_F2978_ = F2940 & new_F2977_;
  assign new_F2979_ = F2938 & ~new_F2948_;
  assign new_F2980_ = ~F2938 & new_F2948_;
  assign new_F2981_ = ~F2937 | ~new_F2962_;
  assign new_F2982_ = new_F2948_ & new_F2981_;
  assign new_F2983_ = ~new_F2948_ & ~new_F2982_;
  assign new_F2984_ = new_F2948_ | new_F2981_;
  assign new_F2985_ = ~F2938 & F2939;
  assign new_F2986_ = F2938 & ~F2939;
  assign new_F2987_ = new_F2955_ | new_F2992_;
  assign new_F2988_ = ~new_F2955_ & ~new_F2991_;
  assign new_F2989_ = F2938 | new_F2955_;
  assign new_F2990_ = F2938 | F2939;
  assign new_F2991_ = new_F2955_ & new_F2992_;
  assign new_F2992_ = ~F2937 | ~new_F2962_;
  assign new_F2993_ = new_F2970_ & new_F2990_;
  assign new_F2994_ = ~new_F2970_ & ~new_F2990_;
  assign new_F2995_ = new_F2999_ | new_F3000_;
  assign new_F2996_ = ~F2941 & new_F2955_;
  assign new_F2997_ = new_F3001_ | new_F3002_;
  assign new_F2998_ = F2941 & new_F2955_;
  assign new_F2999_ = ~F2941 & ~new_F2955_;
  assign new_F3000_ = F2941 & ~new_F2955_;
  assign new_F3001_ = F2941 & ~new_F2955_;
  assign new_F3002_ = ~F2941 & new_F2955_;
  assign new_F3009_ = new_F3016_ & new_F3015_;
  assign new_F3010_ = new_F3018_ | new_F3017_;
  assign new_F3011_ = new_F3020_ | new_F3019_;
  assign new_F3012_ = new_F3022_ & new_F3021_;
  assign new_F3013_ = new_F3022_ & new_F3023_;
  assign new_F3014_ = new_F3015_ | new_F3024_;
  assign new_F3015_ = F3004 | new_F3027_;
  assign new_F3016_ = new_F3026_ | new_F3025_;
  assign new_F3017_ = new_F3031_ & new_F3030_;
  assign new_F3018_ = new_F3029_ & new_F3028_;
  assign new_F3019_ = new_F3034_ | new_F3033_;
  assign new_F3020_ = new_F3029_ & new_F3032_;
  assign new_F3021_ = F3004 | new_F3037_;
  assign new_F3022_ = new_F3036_ | new_F3035_;
  assign new_F3023_ = new_F3039_ | new_F3038_;
  assign new_F3024_ = ~new_F3015_ & new_F3041_;
  assign new_F3025_ = ~new_F3017_ & new_F3029_;
  assign new_F3026_ = new_F3017_ & ~new_F3029_;
  assign new_F3027_ = F3003 & ~F3004;
  assign new_F3028_ = ~new_F3050_ | ~new_F3051_;
  assign new_F3029_ = new_F3043_ | new_F3045_;
  assign new_F3030_ = new_F3053_ | new_F3052_;
  assign new_F3031_ = new_F3047_ | new_F3046_;
  assign new_F3032_ = ~new_F3055_ | ~new_F3054_;
  assign new_F3033_ = ~new_F3056_ & new_F3057_;
  assign new_F3034_ = new_F3056_ & ~new_F3057_;
  assign new_F3035_ = ~F3003 & F3004;
  assign new_F3036_ = F3003 & ~F3004;
  assign new_F3037_ = ~new_F3019_ | new_F3029_;
  assign new_F3038_ = new_F3019_ & new_F3029_;
  assign new_F3039_ = ~new_F3019_ & ~new_F3029_;
  assign new_F3040_ = new_F3061_ | new_F3060_;
  assign new_F3041_ = F3007 | new_F3040_;
  assign new_F3042_ = new_F3065_ | new_F3064_;
  assign new_F3043_ = ~F3007 & new_F3042_;
  assign new_F3044_ = new_F3063_ | new_F3062_;
  assign new_F3045_ = F3007 & new_F3044_;
  assign new_F3046_ = F3005 & ~new_F3015_;
  assign new_F3047_ = ~F3005 & new_F3015_;
  assign new_F3048_ = ~F3004 | ~new_F3029_;
  assign new_F3049_ = new_F3015_ & new_F3048_;
  assign new_F3050_ = ~new_F3015_ & ~new_F3049_;
  assign new_F3051_ = new_F3015_ | new_F3048_;
  assign new_F3052_ = ~F3005 & F3006;
  assign new_F3053_ = F3005 & ~F3006;
  assign new_F3054_ = new_F3022_ | new_F3059_;
  assign new_F3055_ = ~new_F3022_ & ~new_F3058_;
  assign new_F3056_ = F3005 | new_F3022_;
  assign new_F3057_ = F3005 | F3006;
  assign new_F3058_ = new_F3022_ & new_F3059_;
  assign new_F3059_ = ~F3004 | ~new_F3029_;
  assign new_F3060_ = new_F3037_ & new_F3057_;
  assign new_F3061_ = ~new_F3037_ & ~new_F3057_;
  assign new_F3062_ = new_F3066_ | new_F3067_;
  assign new_F3063_ = ~F3008 & new_F3022_;
  assign new_F3064_ = new_F3068_ | new_F3069_;
  assign new_F3065_ = F3008 & new_F3022_;
  assign new_F3066_ = ~F3008 & ~new_F3022_;
  assign new_F3067_ = F3008 & ~new_F3022_;
  assign new_F3068_ = F3008 & ~new_F3022_;
  assign new_F3069_ = ~F3008 & new_F3022_;
  assign new_F3076_ = new_F3083_ & new_F3082_;
  assign new_F3077_ = new_F3085_ | new_F3084_;
  assign new_F3078_ = new_F3087_ | new_F3086_;
  assign new_F3079_ = new_F3089_ & new_F3088_;
  assign new_F3080_ = new_F3089_ & new_F3090_;
  assign new_F3081_ = new_F3082_ | new_F3091_;
  assign new_F3082_ = F3071 | new_F3094_;
  assign new_F3083_ = new_F3093_ | new_F3092_;
  assign new_F3084_ = new_F3098_ & new_F3097_;
  assign new_F3085_ = new_F3096_ & new_F3095_;
  assign new_F3086_ = new_F3101_ | new_F3100_;
  assign new_F3087_ = new_F3096_ & new_F3099_;
  assign new_F3088_ = F3071 | new_F3104_;
  assign new_F3089_ = new_F3103_ | new_F3102_;
  assign new_F3090_ = new_F3106_ | new_F3105_;
  assign new_F3091_ = ~new_F3082_ & new_F3108_;
  assign new_F3092_ = ~new_F3084_ & new_F3096_;
  assign new_F3093_ = new_F3084_ & ~new_F3096_;
  assign new_F3094_ = F3070 & ~F3071;
  assign new_F3095_ = ~new_F3117_ | ~new_F3118_;
  assign new_F3096_ = new_F3110_ | new_F3112_;
  assign new_F3097_ = new_F3120_ | new_F3119_;
  assign new_F3098_ = new_F3114_ | new_F3113_;
  assign new_F3099_ = ~new_F3122_ | ~new_F3121_;
  assign new_F3100_ = ~new_F3123_ & new_F3124_;
  assign new_F3101_ = new_F3123_ & ~new_F3124_;
  assign new_F3102_ = ~F3070 & F3071;
  assign new_F3103_ = F3070 & ~F3071;
  assign new_F3104_ = ~new_F3086_ | new_F3096_;
  assign new_F3105_ = new_F3086_ & new_F3096_;
  assign new_F3106_ = ~new_F3086_ & ~new_F3096_;
  assign new_F3107_ = new_F3128_ | new_F3127_;
  assign new_F3108_ = F3074 | new_F3107_;
  assign new_F3109_ = new_F3132_ | new_F3131_;
  assign new_F3110_ = ~F3074 & new_F3109_;
  assign new_F3111_ = new_F3130_ | new_F3129_;
  assign new_F3112_ = F3074 & new_F3111_;
  assign new_F3113_ = F3072 & ~new_F3082_;
  assign new_F3114_ = ~F3072 & new_F3082_;
  assign new_F3115_ = ~F3071 | ~new_F3096_;
  assign new_F3116_ = new_F3082_ & new_F3115_;
  assign new_F3117_ = ~new_F3082_ & ~new_F3116_;
  assign new_F3118_ = new_F3082_ | new_F3115_;
  assign new_F3119_ = ~F3072 & F3073;
  assign new_F3120_ = F3072 & ~F3073;
  assign new_F3121_ = new_F3089_ | new_F3126_;
  assign new_F3122_ = ~new_F3089_ & ~new_F3125_;
  assign new_F3123_ = F3072 | new_F3089_;
  assign new_F3124_ = F3072 | F3073;
  assign new_F3125_ = new_F3089_ & new_F3126_;
  assign new_F3126_ = ~F3071 | ~new_F3096_;
  assign new_F3127_ = new_F3104_ & new_F3124_;
  assign new_F3128_ = ~new_F3104_ & ~new_F3124_;
  assign new_F3129_ = new_F3133_ | new_F3134_;
  assign new_F3130_ = ~F3075 & new_F3089_;
  assign new_F3131_ = new_F3135_ | new_F3136_;
  assign new_F3132_ = F3075 & new_F3089_;
  assign new_F3133_ = ~F3075 & ~new_F3089_;
  assign new_F3134_ = F3075 & ~new_F3089_;
  assign new_F3135_ = F3075 & ~new_F3089_;
  assign new_F3136_ = ~F3075 & new_F3089_;
  assign new_F3143_ = new_F3150_ & new_F3149_;
  assign new_F3144_ = new_F3152_ | new_F3151_;
  assign new_F3145_ = new_F3154_ | new_F3153_;
  assign new_F3146_ = new_F3156_ & new_F3155_;
  assign new_F3147_ = new_F3156_ & new_F3157_;
  assign new_F3148_ = new_F3149_ | new_F3158_;
  assign new_F3149_ = F3138 | new_F3161_;
  assign new_F3150_ = new_F3160_ | new_F3159_;
  assign new_F3151_ = new_F3165_ & new_F3164_;
  assign new_F3152_ = new_F3163_ & new_F3162_;
  assign new_F3153_ = new_F3168_ | new_F3167_;
  assign new_F3154_ = new_F3163_ & new_F3166_;
  assign new_F3155_ = F3138 | new_F3171_;
  assign new_F3156_ = new_F3170_ | new_F3169_;
  assign new_F3157_ = new_F3173_ | new_F3172_;
  assign new_F3158_ = ~new_F3149_ & new_F3175_;
  assign new_F3159_ = ~new_F3151_ & new_F3163_;
  assign new_F3160_ = new_F3151_ & ~new_F3163_;
  assign new_F3161_ = F3137 & ~F3138;
  assign new_F3162_ = ~new_F3184_ | ~new_F3185_;
  assign new_F3163_ = new_F3177_ | new_F3179_;
  assign new_F3164_ = new_F3187_ | new_F3186_;
  assign new_F3165_ = new_F3181_ | new_F3180_;
  assign new_F3166_ = ~new_F3189_ | ~new_F3188_;
  assign new_F3167_ = ~new_F3190_ & new_F3191_;
  assign new_F3168_ = new_F3190_ & ~new_F3191_;
  assign new_F3169_ = ~F3137 & F3138;
  assign new_F3170_ = F3137 & ~F3138;
  assign new_F3171_ = ~new_F3153_ | new_F3163_;
  assign new_F3172_ = new_F3153_ & new_F3163_;
  assign new_F3173_ = ~new_F3153_ & ~new_F3163_;
  assign new_F3174_ = new_F3195_ | new_F3194_;
  assign new_F3175_ = F3141 | new_F3174_;
  assign new_F3176_ = new_F3199_ | new_F3198_;
  assign new_F3177_ = ~F3141 & new_F3176_;
  assign new_F3178_ = new_F3197_ | new_F3196_;
  assign new_F3179_ = F3141 & new_F3178_;
  assign new_F3180_ = F3139 & ~new_F3149_;
  assign new_F3181_ = ~F3139 & new_F3149_;
  assign new_F3182_ = ~F3138 | ~new_F3163_;
  assign new_F3183_ = new_F3149_ & new_F3182_;
  assign new_F3184_ = ~new_F3149_ & ~new_F3183_;
  assign new_F3185_ = new_F3149_ | new_F3182_;
  assign new_F3186_ = ~F3139 & F3140;
  assign new_F3187_ = F3139 & ~F3140;
  assign new_F3188_ = new_F3156_ | new_F3193_;
  assign new_F3189_ = ~new_F3156_ & ~new_F3192_;
  assign new_F3190_ = F3139 | new_F3156_;
  assign new_F3191_ = F3139 | F3140;
  assign new_F3192_ = new_F3156_ & new_F3193_;
  assign new_F3193_ = ~F3138 | ~new_F3163_;
  assign new_F3194_ = new_F3171_ & new_F3191_;
  assign new_F3195_ = ~new_F3171_ & ~new_F3191_;
  assign new_F3196_ = new_F3200_ | new_F3201_;
  assign new_F3197_ = ~F3142 & new_F3156_;
  assign new_F3198_ = new_F3202_ | new_F3203_;
  assign new_F3199_ = F3142 & new_F3156_;
  assign new_F3200_ = ~F3142 & ~new_F3156_;
  assign new_F3201_ = F3142 & ~new_F3156_;
  assign new_F3202_ = F3142 & ~new_F3156_;
  assign new_F3203_ = ~F3142 & new_F3156_;
  assign new_F3210_ = new_F3217_ & new_F3216_;
  assign new_F3211_ = new_F3219_ | new_F3218_;
  assign new_F3212_ = new_F3221_ | new_F3220_;
  assign new_F3213_ = new_F3223_ & new_F3222_;
  assign new_F3214_ = new_F3223_ & new_F3224_;
  assign new_F3215_ = new_F3216_ | new_F3225_;
  assign new_F3216_ = F3205 | new_F3228_;
  assign new_F3217_ = new_F3227_ | new_F3226_;
  assign new_F3218_ = new_F3232_ & new_F3231_;
  assign new_F3219_ = new_F3230_ & new_F3229_;
  assign new_F3220_ = new_F3235_ | new_F3234_;
  assign new_F3221_ = new_F3230_ & new_F3233_;
  assign new_F3222_ = F3205 | new_F3238_;
  assign new_F3223_ = new_F3237_ | new_F3236_;
  assign new_F3224_ = new_F3240_ | new_F3239_;
  assign new_F3225_ = ~new_F3216_ & new_F3242_;
  assign new_F3226_ = ~new_F3218_ & new_F3230_;
  assign new_F3227_ = new_F3218_ & ~new_F3230_;
  assign new_F3228_ = F3204 & ~F3205;
  assign new_F3229_ = ~new_F3251_ | ~new_F3252_;
  assign new_F3230_ = new_F3244_ | new_F3246_;
  assign new_F3231_ = new_F3254_ | new_F3253_;
  assign new_F3232_ = new_F3248_ | new_F3247_;
  assign new_F3233_ = ~new_F3256_ | ~new_F3255_;
  assign new_F3234_ = ~new_F3257_ & new_F3258_;
  assign new_F3235_ = new_F3257_ & ~new_F3258_;
  assign new_F3236_ = ~F3204 & F3205;
  assign new_F3237_ = F3204 & ~F3205;
  assign new_F3238_ = ~new_F3220_ | new_F3230_;
  assign new_F3239_ = new_F3220_ & new_F3230_;
  assign new_F3240_ = ~new_F3220_ & ~new_F3230_;
  assign new_F3241_ = new_F3262_ | new_F3261_;
  assign new_F3242_ = F3208 | new_F3241_;
  assign new_F3243_ = new_F3266_ | new_F3265_;
  assign new_F3244_ = ~F3208 & new_F3243_;
  assign new_F3245_ = new_F3264_ | new_F3263_;
  assign new_F3246_ = F3208 & new_F3245_;
  assign new_F3247_ = F3206 & ~new_F3216_;
  assign new_F3248_ = ~F3206 & new_F3216_;
  assign new_F3249_ = ~F3205 | ~new_F3230_;
  assign new_F3250_ = new_F3216_ & new_F3249_;
  assign new_F3251_ = ~new_F3216_ & ~new_F3250_;
  assign new_F3252_ = new_F3216_ | new_F3249_;
  assign new_F3253_ = ~F3206 & F3207;
  assign new_F3254_ = F3206 & ~F3207;
  assign new_F3255_ = new_F3223_ | new_F3260_;
  assign new_F3256_ = ~new_F3223_ & ~new_F3259_;
  assign new_F3257_ = F3206 | new_F3223_;
  assign new_F3258_ = F3206 | F3207;
  assign new_F3259_ = new_F3223_ & new_F3260_;
  assign new_F3260_ = ~F3205 | ~new_F3230_;
  assign new_F3261_ = new_F3238_ & new_F3258_;
  assign new_F3262_ = ~new_F3238_ & ~new_F3258_;
  assign new_F3263_ = new_F3267_ | new_F3268_;
  assign new_F3264_ = ~F3209 & new_F3223_;
  assign new_F3265_ = new_F3269_ | new_F3270_;
  assign new_F3266_ = F3209 & new_F3223_;
  assign new_F3267_ = ~F3209 & ~new_F3223_;
  assign new_F3268_ = F3209 & ~new_F3223_;
  assign new_F3269_ = F3209 & ~new_F3223_;
  assign new_F3270_ = ~F3209 & new_F3223_;
  assign new_F3277_ = new_F3284_ & new_F3283_;
  assign new_F3278_ = new_F3286_ | new_F3285_;
  assign new_F3279_ = new_F3288_ | new_F3287_;
  assign new_F3280_ = new_F3290_ & new_F3289_;
  assign new_F3281_ = new_F3290_ & new_F3291_;
  assign new_F3282_ = new_F3283_ | new_F3292_;
  assign new_F3283_ = F3272 | new_F3295_;
  assign new_F3284_ = new_F3294_ | new_F3293_;
  assign new_F3285_ = new_F3299_ & new_F3298_;
  assign new_F3286_ = new_F3297_ & new_F3296_;
  assign new_F3287_ = new_F3302_ | new_F3301_;
  assign new_F3288_ = new_F3297_ & new_F3300_;
  assign new_F3289_ = F3272 | new_F3305_;
  assign new_F3290_ = new_F3304_ | new_F3303_;
  assign new_F3291_ = new_F3307_ | new_F3306_;
  assign new_F3292_ = ~new_F3283_ & new_F3309_;
  assign new_F3293_ = ~new_F3285_ & new_F3297_;
  assign new_F3294_ = new_F3285_ & ~new_F3297_;
  assign new_F3295_ = F3271 & ~F3272;
  assign new_F3296_ = ~new_F3318_ | ~new_F3319_;
  assign new_F3297_ = new_F3311_ | new_F3313_;
  assign new_F3298_ = new_F3321_ | new_F3320_;
  assign new_F3299_ = new_F3315_ | new_F3314_;
  assign new_F3300_ = ~new_F3323_ | ~new_F3322_;
  assign new_F3301_ = ~new_F3324_ & new_F3325_;
  assign new_F3302_ = new_F3324_ & ~new_F3325_;
  assign new_F3303_ = ~F3271 & F3272;
  assign new_F3304_ = F3271 & ~F3272;
  assign new_F3305_ = ~new_F3287_ | new_F3297_;
  assign new_F3306_ = new_F3287_ & new_F3297_;
  assign new_F3307_ = ~new_F3287_ & ~new_F3297_;
  assign new_F3308_ = new_F3329_ | new_F3328_;
  assign new_F3309_ = F3275 | new_F3308_;
  assign new_F3310_ = new_F3333_ | new_F3332_;
  assign new_F3311_ = ~F3275 & new_F3310_;
  assign new_F3312_ = new_F3331_ | new_F3330_;
  assign new_F3313_ = F3275 & new_F3312_;
  assign new_F3314_ = F3273 & ~new_F3283_;
  assign new_F3315_ = ~F3273 & new_F3283_;
  assign new_F3316_ = ~F3272 | ~new_F3297_;
  assign new_F3317_ = new_F3283_ & new_F3316_;
  assign new_F3318_ = ~new_F3283_ & ~new_F3317_;
  assign new_F3319_ = new_F3283_ | new_F3316_;
  assign new_F3320_ = ~F3273 & F3274;
  assign new_F3321_ = F3273 & ~F3274;
  assign new_F3322_ = new_F3290_ | new_F3327_;
  assign new_F3323_ = ~new_F3290_ & ~new_F3326_;
  assign new_F3324_ = F3273 | new_F3290_;
  assign new_F3325_ = F3273 | F3274;
  assign new_F3326_ = new_F3290_ & new_F3327_;
  assign new_F3327_ = ~F3272 | ~new_F3297_;
  assign new_F3328_ = new_F3305_ & new_F3325_;
  assign new_F3329_ = ~new_F3305_ & ~new_F3325_;
  assign new_F3330_ = new_F3334_ | new_F3335_;
  assign new_F3331_ = ~F3276 & new_F3290_;
  assign new_F3332_ = new_F3336_ | new_F3337_;
  assign new_F3333_ = F3276 & new_F3290_;
  assign new_F3334_ = ~F3276 & ~new_F3290_;
  assign new_F3335_ = F3276 & ~new_F3290_;
  assign new_F3336_ = F3276 & ~new_F3290_;
  assign new_F3337_ = ~F3276 & new_F3290_;
  assign new_F3344_ = new_F3351_ & new_F3350_;
  assign new_F3345_ = new_F3353_ | new_F3352_;
  assign new_F3346_ = new_F3355_ | new_F3354_;
  assign new_F3347_ = new_F3357_ & new_F3356_;
  assign new_F3348_ = new_F3357_ & new_F3358_;
  assign new_F3349_ = new_F3350_ | new_F3359_;
  assign new_F3350_ = F3339 | new_F3362_;
  assign new_F3351_ = new_F3361_ | new_F3360_;
  assign new_F3352_ = new_F3366_ & new_F3365_;
  assign new_F3353_ = new_F3364_ & new_F3363_;
  assign new_F3354_ = new_F3369_ | new_F3368_;
  assign new_F3355_ = new_F3364_ & new_F3367_;
  assign new_F3356_ = F3339 | new_F3372_;
  assign new_F3357_ = new_F3371_ | new_F3370_;
  assign new_F3358_ = new_F3374_ | new_F3373_;
  assign new_F3359_ = ~new_F3350_ & new_F3376_;
  assign new_F3360_ = ~new_F3352_ & new_F3364_;
  assign new_F3361_ = new_F3352_ & ~new_F3364_;
  assign new_F3362_ = F3338 & ~F3339;
  assign new_F3363_ = ~new_F3385_ | ~new_F3386_;
  assign new_F3364_ = new_F3378_ | new_F3380_;
  assign new_F3365_ = new_F3388_ | new_F3387_;
  assign new_F3366_ = new_F3382_ | new_F3381_;
  assign new_F3367_ = ~new_F3390_ | ~new_F3389_;
  assign new_F3368_ = ~new_F3391_ & new_F3392_;
  assign new_F3369_ = new_F3391_ & ~new_F3392_;
  assign new_F3370_ = ~F3338 & F3339;
  assign new_F3371_ = F3338 & ~F3339;
  assign new_F3372_ = ~new_F3354_ | new_F3364_;
  assign new_F3373_ = new_F3354_ & new_F3364_;
  assign new_F3374_ = ~new_F3354_ & ~new_F3364_;
  assign new_F3375_ = new_F3396_ | new_F3395_;
  assign new_F3376_ = F3342 | new_F3375_;
  assign new_F3377_ = new_F3400_ | new_F3399_;
  assign new_F3378_ = ~F3342 & new_F3377_;
  assign new_F3379_ = new_F3398_ | new_F3397_;
  assign new_F3380_ = F3342 & new_F3379_;
  assign new_F3381_ = F3340 & ~new_F3350_;
  assign new_F3382_ = ~F3340 & new_F3350_;
  assign new_F3383_ = ~F3339 | ~new_F3364_;
  assign new_F3384_ = new_F3350_ & new_F3383_;
  assign new_F3385_ = ~new_F3350_ & ~new_F3384_;
  assign new_F3386_ = new_F3350_ | new_F3383_;
  assign new_F3387_ = ~F3340 & F3341;
  assign new_F3388_ = F3340 & ~F3341;
  assign new_F3389_ = new_F3357_ | new_F3394_;
  assign new_F3390_ = ~new_F3357_ & ~new_F3393_;
  assign new_F3391_ = F3340 | new_F3357_;
  assign new_F3392_ = F3340 | F3341;
  assign new_F3393_ = new_F3357_ & new_F3394_;
  assign new_F3394_ = ~F3339 | ~new_F3364_;
  assign new_F3395_ = new_F3372_ & new_F3392_;
  assign new_F3396_ = ~new_F3372_ & ~new_F3392_;
  assign new_F3397_ = new_F3401_ | new_F3402_;
  assign new_F3398_ = ~F3343 & new_F3357_;
  assign new_F3399_ = new_F3403_ | new_F3404_;
  assign new_F3400_ = F3343 & new_F3357_;
  assign new_F3401_ = ~F3343 & ~new_F3357_;
  assign new_F3402_ = F3343 & ~new_F3357_;
  assign new_F3403_ = F3343 & ~new_F3357_;
  assign new_F3404_ = ~F3343 & new_F3357_;
  assign new_F3411_ = new_F3418_ & new_F3417_;
  assign new_F3412_ = new_F3420_ | new_F3419_;
  assign new_F3413_ = new_F3422_ | new_F3421_;
  assign new_F3414_ = new_F3424_ & new_F3423_;
  assign new_F3415_ = new_F3424_ & new_F3425_;
  assign new_F3416_ = new_F3417_ | new_F3426_;
  assign new_F3417_ = F3406 | new_F3429_;
  assign new_F3418_ = new_F3428_ | new_F3427_;
  assign new_F3419_ = new_F3433_ & new_F3432_;
  assign new_F3420_ = new_F3431_ & new_F3430_;
  assign new_F3421_ = new_F3436_ | new_F3435_;
  assign new_F3422_ = new_F3431_ & new_F3434_;
  assign new_F3423_ = F3406 | new_F3439_;
  assign new_F3424_ = new_F3438_ | new_F3437_;
  assign new_F3425_ = new_F3441_ | new_F3440_;
  assign new_F3426_ = ~new_F3417_ & new_F3443_;
  assign new_F3427_ = ~new_F3419_ & new_F3431_;
  assign new_F3428_ = new_F3419_ & ~new_F3431_;
  assign new_F3429_ = F3405 & ~F3406;
  assign new_F3430_ = ~new_F3452_ | ~new_F3453_;
  assign new_F3431_ = new_F3445_ | new_F3447_;
  assign new_F3432_ = new_F3455_ | new_F3454_;
  assign new_F3433_ = new_F3449_ | new_F3448_;
  assign new_F3434_ = ~new_F3457_ | ~new_F3456_;
  assign new_F3435_ = ~new_F3458_ & new_F3459_;
  assign new_F3436_ = new_F3458_ & ~new_F3459_;
  assign new_F3437_ = ~F3405 & F3406;
  assign new_F3438_ = F3405 & ~F3406;
  assign new_F3439_ = ~new_F3421_ | new_F3431_;
  assign new_F3440_ = new_F3421_ & new_F3431_;
  assign new_F3441_ = ~new_F3421_ & ~new_F3431_;
  assign new_F3442_ = new_F3463_ | new_F3462_;
  assign new_F3443_ = F3409 | new_F3442_;
  assign new_F3444_ = new_F3467_ | new_F3466_;
  assign new_F3445_ = ~F3409 & new_F3444_;
  assign new_F3446_ = new_F3465_ | new_F3464_;
  assign new_F3447_ = F3409 & new_F3446_;
  assign new_F3448_ = F3407 & ~new_F3417_;
  assign new_F3449_ = ~F3407 & new_F3417_;
  assign new_F3450_ = ~F3406 | ~new_F3431_;
  assign new_F3451_ = new_F3417_ & new_F3450_;
  assign new_F3452_ = ~new_F3417_ & ~new_F3451_;
  assign new_F3453_ = new_F3417_ | new_F3450_;
  assign new_F3454_ = ~F3407 & F3408;
  assign new_F3455_ = F3407 & ~F3408;
  assign new_F3456_ = new_F3424_ | new_F3461_;
  assign new_F3457_ = ~new_F3424_ & ~new_F3460_;
  assign new_F3458_ = F3407 | new_F3424_;
  assign new_F3459_ = F3407 | F3408;
  assign new_F3460_ = new_F3424_ & new_F3461_;
  assign new_F3461_ = ~F3406 | ~new_F3431_;
  assign new_F3462_ = new_F3439_ & new_F3459_;
  assign new_F3463_ = ~new_F3439_ & ~new_F3459_;
  assign new_F3464_ = new_F3468_ | new_F3469_;
  assign new_F3465_ = ~F3410 & new_F3424_;
  assign new_F3466_ = new_F3470_ | new_F3471_;
  assign new_F3467_ = F3410 & new_F3424_;
  assign new_F3468_ = ~F3410 & ~new_F3424_;
  assign new_F3469_ = F3410 & ~new_F3424_;
  assign new_F3470_ = F3410 & ~new_F3424_;
  assign new_F3471_ = ~F3410 & new_F3424_;
  assign new_F3478_ = new_F3485_ & new_F3484_;
  assign new_F3479_ = new_F3487_ | new_F3486_;
  assign new_F3480_ = new_F3489_ | new_F3488_;
  assign new_F3481_ = new_F3491_ & new_F3490_;
  assign new_F3482_ = new_F3491_ & new_F3492_;
  assign new_F3483_ = new_F3484_ | new_F3493_;
  assign new_F3484_ = F3473 | new_F3496_;
  assign new_F3485_ = new_F3495_ | new_F3494_;
  assign new_F3486_ = new_F3500_ & new_F3499_;
  assign new_F3487_ = new_F3498_ & new_F3497_;
  assign new_F3488_ = new_F3503_ | new_F3502_;
  assign new_F3489_ = new_F3498_ & new_F3501_;
  assign new_F3490_ = F3473 | new_F3506_;
  assign new_F3491_ = new_F3505_ | new_F3504_;
  assign new_F3492_ = new_F3508_ | new_F3507_;
  assign new_F3493_ = ~new_F3484_ & new_F3510_;
  assign new_F3494_ = ~new_F3486_ & new_F3498_;
  assign new_F3495_ = new_F3486_ & ~new_F3498_;
  assign new_F3496_ = F3472 & ~F3473;
  assign new_F3497_ = ~new_F3519_ | ~new_F3520_;
  assign new_F3498_ = new_F3512_ | new_F3514_;
  assign new_F3499_ = new_F3522_ | new_F3521_;
  assign new_F3500_ = new_F3516_ | new_F3515_;
  assign new_F3501_ = ~new_F3524_ | ~new_F3523_;
  assign new_F3502_ = ~new_F3525_ & new_F3526_;
  assign new_F3503_ = new_F3525_ & ~new_F3526_;
  assign new_F3504_ = ~F3472 & F3473;
  assign new_F3505_ = F3472 & ~F3473;
  assign new_F3506_ = ~new_F3488_ | new_F3498_;
  assign new_F3507_ = new_F3488_ & new_F3498_;
  assign new_F3508_ = ~new_F3488_ & ~new_F3498_;
  assign new_F3509_ = new_F3530_ | new_F3529_;
  assign new_F3510_ = F3476 | new_F3509_;
  assign new_F3511_ = new_F3534_ | new_F3533_;
  assign new_F3512_ = ~F3476 & new_F3511_;
  assign new_F3513_ = new_F3532_ | new_F3531_;
  assign new_F3514_ = F3476 & new_F3513_;
  assign new_F3515_ = F3474 & ~new_F3484_;
  assign new_F3516_ = ~F3474 & new_F3484_;
  assign new_F3517_ = ~F3473 | ~new_F3498_;
  assign new_F3518_ = new_F3484_ & new_F3517_;
  assign new_F3519_ = ~new_F3484_ & ~new_F3518_;
  assign new_F3520_ = new_F3484_ | new_F3517_;
  assign new_F3521_ = ~F3474 & F3475;
  assign new_F3522_ = F3474 & ~F3475;
  assign new_F3523_ = new_F3491_ | new_F3528_;
  assign new_F3524_ = ~new_F3491_ & ~new_F3527_;
  assign new_F3525_ = F3474 | new_F3491_;
  assign new_F3526_ = F3474 | F3475;
  assign new_F3527_ = new_F3491_ & new_F3528_;
  assign new_F3528_ = ~F3473 | ~new_F3498_;
  assign new_F3529_ = new_F3506_ & new_F3526_;
  assign new_F3530_ = ~new_F3506_ & ~new_F3526_;
  assign new_F3531_ = new_F3535_ | new_F3536_;
  assign new_F3532_ = ~F3477 & new_F3491_;
  assign new_F3533_ = new_F3537_ | new_F3538_;
  assign new_F3534_ = F3477 & new_F3491_;
  assign new_F3535_ = ~F3477 & ~new_F3491_;
  assign new_F3536_ = F3477 & ~new_F3491_;
  assign new_F3537_ = F3477 & ~new_F3491_;
  assign new_F3538_ = ~F3477 & new_F3491_;
  assign new_F3545_ = new_F3552_ & new_F3551_;
  assign new_F3546_ = new_F3554_ | new_F3553_;
  assign new_F3547_ = new_F3556_ | new_F3555_;
  assign new_F3548_ = new_F3558_ & new_F3557_;
  assign new_F3549_ = new_F3558_ & new_F3559_;
  assign new_F3550_ = new_F3551_ | new_F3560_;
  assign new_F3551_ = F3540 | new_F3563_;
  assign new_F3552_ = new_F3562_ | new_F3561_;
  assign new_F3553_ = new_F3567_ & new_F3566_;
  assign new_F3554_ = new_F3565_ & new_F3564_;
  assign new_F3555_ = new_F3570_ | new_F3569_;
  assign new_F3556_ = new_F3565_ & new_F3568_;
  assign new_F3557_ = F3540 | new_F3573_;
  assign new_F3558_ = new_F3572_ | new_F3571_;
  assign new_F3559_ = new_F3575_ | new_F3574_;
  assign new_F3560_ = ~new_F3551_ & new_F3577_;
  assign new_F3561_ = ~new_F3553_ & new_F3565_;
  assign new_F3562_ = new_F3553_ & ~new_F3565_;
  assign new_F3563_ = F3539 & ~F3540;
  assign new_F3564_ = ~new_F3586_ | ~new_F3587_;
  assign new_F3565_ = new_F3579_ | new_F3581_;
  assign new_F3566_ = new_F3589_ | new_F3588_;
  assign new_F3567_ = new_F3583_ | new_F3582_;
  assign new_F3568_ = ~new_F3591_ | ~new_F3590_;
  assign new_F3569_ = ~new_F3592_ & new_F3593_;
  assign new_F3570_ = new_F3592_ & ~new_F3593_;
  assign new_F3571_ = ~F3539 & F3540;
  assign new_F3572_ = F3539 & ~F3540;
  assign new_F3573_ = ~new_F3555_ | new_F3565_;
  assign new_F3574_ = new_F3555_ & new_F3565_;
  assign new_F3575_ = ~new_F3555_ & ~new_F3565_;
  assign new_F3576_ = new_F3597_ | new_F3596_;
  assign new_F3577_ = F3543 | new_F3576_;
  assign new_F3578_ = new_F3601_ | new_F3600_;
  assign new_F3579_ = ~F3543 & new_F3578_;
  assign new_F3580_ = new_F3599_ | new_F3598_;
  assign new_F3581_ = F3543 & new_F3580_;
  assign new_F3582_ = F3541 & ~new_F3551_;
  assign new_F3583_ = ~F3541 & new_F3551_;
  assign new_F3584_ = ~F3540 | ~new_F3565_;
  assign new_F3585_ = new_F3551_ & new_F3584_;
  assign new_F3586_ = ~new_F3551_ & ~new_F3585_;
  assign new_F3587_ = new_F3551_ | new_F3584_;
  assign new_F3588_ = ~F3541 & F3542;
  assign new_F3589_ = F3541 & ~F3542;
  assign new_F3590_ = new_F3558_ | new_F3595_;
  assign new_F3591_ = ~new_F3558_ & ~new_F3594_;
  assign new_F3592_ = F3541 | new_F3558_;
  assign new_F3593_ = F3541 | F3542;
  assign new_F3594_ = new_F3558_ & new_F3595_;
  assign new_F3595_ = ~F3540 | ~new_F3565_;
  assign new_F3596_ = new_F3573_ & new_F3593_;
  assign new_F3597_ = ~new_F3573_ & ~new_F3593_;
  assign new_F3598_ = new_F3602_ | new_F3603_;
  assign new_F3599_ = ~F3544 & new_F3558_;
  assign new_F3600_ = new_F3604_ | new_F3605_;
  assign new_F3601_ = F3544 & new_F3558_;
  assign new_F3602_ = ~F3544 & ~new_F3558_;
  assign new_F3603_ = F3544 & ~new_F3558_;
  assign new_F3604_ = F3544 & ~new_F3558_;
  assign new_F3605_ = ~F3544 & new_F3558_;
  assign new_F3612_ = new_F3619_ & new_F3618_;
  assign new_F3613_ = new_F3621_ | new_F3620_;
  assign new_F3614_ = new_F3623_ | new_F3622_;
  assign new_F3615_ = new_F3625_ & new_F3624_;
  assign new_F3616_ = new_F3625_ & new_F3626_;
  assign new_F3617_ = new_F3618_ | new_F3627_;
  assign new_F3618_ = F3607 | new_F3630_;
  assign new_F3619_ = new_F3629_ | new_F3628_;
  assign new_F3620_ = new_F3634_ & new_F3633_;
  assign new_F3621_ = new_F3632_ & new_F3631_;
  assign new_F3622_ = new_F3637_ | new_F3636_;
  assign new_F3623_ = new_F3632_ & new_F3635_;
  assign new_F3624_ = F3607 | new_F3640_;
  assign new_F3625_ = new_F3639_ | new_F3638_;
  assign new_F3626_ = new_F3642_ | new_F3641_;
  assign new_F3627_ = ~new_F3618_ & new_F3644_;
  assign new_F3628_ = ~new_F3620_ & new_F3632_;
  assign new_F3629_ = new_F3620_ & ~new_F3632_;
  assign new_F3630_ = F3606 & ~F3607;
  assign new_F3631_ = ~new_F3653_ | ~new_F3654_;
  assign new_F3632_ = new_F3646_ | new_F3648_;
  assign new_F3633_ = new_F3656_ | new_F3655_;
  assign new_F3634_ = new_F3650_ | new_F3649_;
  assign new_F3635_ = ~new_F3658_ | ~new_F3657_;
  assign new_F3636_ = ~new_F3659_ & new_F3660_;
  assign new_F3637_ = new_F3659_ & ~new_F3660_;
  assign new_F3638_ = ~F3606 & F3607;
  assign new_F3639_ = F3606 & ~F3607;
  assign new_F3640_ = ~new_F3622_ | new_F3632_;
  assign new_F3641_ = new_F3622_ & new_F3632_;
  assign new_F3642_ = ~new_F3622_ & ~new_F3632_;
  assign new_F3643_ = new_F3664_ | new_F3663_;
  assign new_F3644_ = F3610 | new_F3643_;
  assign new_F3645_ = new_F3668_ | new_F3667_;
  assign new_F3646_ = ~F3610 & new_F3645_;
  assign new_F3647_ = new_F3666_ | new_F3665_;
  assign new_F3648_ = F3610 & new_F3647_;
  assign new_F3649_ = F3608 & ~new_F3618_;
  assign new_F3650_ = ~F3608 & new_F3618_;
  assign new_F3651_ = ~F3607 | ~new_F3632_;
  assign new_F3652_ = new_F3618_ & new_F3651_;
  assign new_F3653_ = ~new_F3618_ & ~new_F3652_;
  assign new_F3654_ = new_F3618_ | new_F3651_;
  assign new_F3655_ = ~F3608 & F3609;
  assign new_F3656_ = F3608 & ~F3609;
  assign new_F3657_ = new_F3625_ | new_F3662_;
  assign new_F3658_ = ~new_F3625_ & ~new_F3661_;
  assign new_F3659_ = F3608 | new_F3625_;
  assign new_F3660_ = F3608 | F3609;
  assign new_F3661_ = new_F3625_ & new_F3662_;
  assign new_F3662_ = ~F3607 | ~new_F3632_;
  assign new_F3663_ = new_F3640_ & new_F3660_;
  assign new_F3664_ = ~new_F3640_ & ~new_F3660_;
  assign new_F3665_ = new_F3669_ | new_F3670_;
  assign new_F3666_ = ~F3611 & new_F3625_;
  assign new_F3667_ = new_F3671_ | new_F3672_;
  assign new_F3668_ = F3611 & new_F3625_;
  assign new_F3669_ = ~F3611 & ~new_F3625_;
  assign new_F3670_ = F3611 & ~new_F3625_;
  assign new_F3671_ = F3611 & ~new_F3625_;
  assign new_F3672_ = ~F3611 & new_F3625_;
  assign new_F3679_ = new_F3686_ & new_F3685_;
  assign new_F3680_ = new_F3688_ | new_F3687_;
  assign new_F3681_ = new_F3690_ | new_F3689_;
  assign new_F3682_ = new_F3692_ & new_F3691_;
  assign new_F3683_ = new_F3692_ & new_F3693_;
  assign new_F3684_ = new_F3685_ | new_F3694_;
  assign new_F3685_ = F3674 | new_F3697_;
  assign new_F3686_ = new_F3696_ | new_F3695_;
  assign new_F3687_ = new_F3701_ & new_F3700_;
  assign new_F3688_ = new_F3699_ & new_F3698_;
  assign new_F3689_ = new_F3704_ | new_F3703_;
  assign new_F3690_ = new_F3699_ & new_F3702_;
  assign new_F3691_ = F3674 | new_F3707_;
  assign new_F3692_ = new_F3706_ | new_F3705_;
  assign new_F3693_ = new_F3709_ | new_F3708_;
  assign new_F3694_ = ~new_F3685_ & new_F3711_;
  assign new_F3695_ = ~new_F3687_ & new_F3699_;
  assign new_F3696_ = new_F3687_ & ~new_F3699_;
  assign new_F3697_ = F3673 & ~F3674;
  assign new_F3698_ = ~new_F3720_ | ~new_F3721_;
  assign new_F3699_ = new_F3713_ | new_F3715_;
  assign new_F3700_ = new_F3723_ | new_F3722_;
  assign new_F3701_ = new_F3717_ | new_F3716_;
  assign new_F3702_ = ~new_F3725_ | ~new_F3724_;
  assign new_F3703_ = ~new_F3726_ & new_F3727_;
  assign new_F3704_ = new_F3726_ & ~new_F3727_;
  assign new_F3705_ = ~F3673 & F3674;
  assign new_F3706_ = F3673 & ~F3674;
  assign new_F3707_ = ~new_F3689_ | new_F3699_;
  assign new_F3708_ = new_F3689_ & new_F3699_;
  assign new_F3709_ = ~new_F3689_ & ~new_F3699_;
  assign new_F3710_ = new_F3731_ | new_F3730_;
  assign new_F3711_ = F3677 | new_F3710_;
  assign new_F3712_ = new_F3735_ | new_F3734_;
  assign new_F3713_ = ~F3677 & new_F3712_;
  assign new_F3714_ = new_F3733_ | new_F3732_;
  assign new_F3715_ = F3677 & new_F3714_;
  assign new_F3716_ = F3675 & ~new_F3685_;
  assign new_F3717_ = ~F3675 & new_F3685_;
  assign new_F3718_ = ~F3674 | ~new_F3699_;
  assign new_F3719_ = new_F3685_ & new_F3718_;
  assign new_F3720_ = ~new_F3685_ & ~new_F3719_;
  assign new_F3721_ = new_F3685_ | new_F3718_;
  assign new_F3722_ = ~F3675 & F3676;
  assign new_F3723_ = F3675 & ~F3676;
  assign new_F3724_ = new_F3692_ | new_F3729_;
  assign new_F3725_ = ~new_F3692_ & ~new_F3728_;
  assign new_F3726_ = F3675 | new_F3692_;
  assign new_F3727_ = F3675 | F3676;
  assign new_F3728_ = new_F3692_ & new_F3729_;
  assign new_F3729_ = ~F3674 | ~new_F3699_;
  assign new_F3730_ = new_F3707_ & new_F3727_;
  assign new_F3731_ = ~new_F3707_ & ~new_F3727_;
  assign new_F3732_ = new_F3736_ | new_F3737_;
  assign new_F3733_ = ~F3678 & new_F3692_;
  assign new_F3734_ = new_F3738_ | new_F3739_;
  assign new_F3735_ = F3678 & new_F3692_;
  assign new_F3736_ = ~F3678 & ~new_F3692_;
  assign new_F3737_ = F3678 & ~new_F3692_;
  assign new_F3738_ = F3678 & ~new_F3692_;
  assign new_F3739_ = ~F3678 & new_F3692_;
  assign new_F3746_ = new_F3753_ & new_F3752_;
  assign new_F3747_ = new_F3755_ | new_F3754_;
  assign new_F3748_ = new_F3757_ | new_F3756_;
  assign new_F3749_ = new_F3759_ & new_F3758_;
  assign new_F3750_ = new_F3759_ & new_F3760_;
  assign new_F3751_ = new_F3752_ | new_F3761_;
  assign new_F3752_ = F3741 | new_F3764_;
  assign new_F3753_ = new_F3763_ | new_F3762_;
  assign new_F3754_ = new_F3768_ & new_F3767_;
  assign new_F3755_ = new_F3766_ & new_F3765_;
  assign new_F3756_ = new_F3771_ | new_F3770_;
  assign new_F3757_ = new_F3766_ & new_F3769_;
  assign new_F3758_ = F3741 | new_F3774_;
  assign new_F3759_ = new_F3773_ | new_F3772_;
  assign new_F3760_ = new_F3776_ | new_F3775_;
  assign new_F3761_ = ~new_F3752_ & new_F3778_;
  assign new_F3762_ = ~new_F3754_ & new_F3766_;
  assign new_F3763_ = new_F3754_ & ~new_F3766_;
  assign new_F3764_ = F3740 & ~F3741;
  assign new_F3765_ = ~new_F3787_ | ~new_F3788_;
  assign new_F3766_ = new_F3780_ | new_F3782_;
  assign new_F3767_ = new_F3790_ | new_F3789_;
  assign new_F3768_ = new_F3784_ | new_F3783_;
  assign new_F3769_ = ~new_F3792_ | ~new_F3791_;
  assign new_F3770_ = ~new_F3793_ & new_F3794_;
  assign new_F3771_ = new_F3793_ & ~new_F3794_;
  assign new_F3772_ = ~F3740 & F3741;
  assign new_F3773_ = F3740 & ~F3741;
  assign new_F3774_ = ~new_F3756_ | new_F3766_;
  assign new_F3775_ = new_F3756_ & new_F3766_;
  assign new_F3776_ = ~new_F3756_ & ~new_F3766_;
  assign new_F3777_ = new_F3798_ | new_F3797_;
  assign new_F3778_ = F3744 | new_F3777_;
  assign new_F3779_ = new_F3802_ | new_F3801_;
  assign new_F3780_ = ~F3744 & new_F3779_;
  assign new_F3781_ = new_F3800_ | new_F3799_;
  assign new_F3782_ = F3744 & new_F3781_;
  assign new_F3783_ = F3742 & ~new_F3752_;
  assign new_F3784_ = ~F3742 & new_F3752_;
  assign new_F3785_ = ~F3741 | ~new_F3766_;
  assign new_F3786_ = new_F3752_ & new_F3785_;
  assign new_F3787_ = ~new_F3752_ & ~new_F3786_;
  assign new_F3788_ = new_F3752_ | new_F3785_;
  assign new_F3789_ = ~F3742 & F3743;
  assign new_F3790_ = F3742 & ~F3743;
  assign new_F3791_ = new_F3759_ | new_F3796_;
  assign new_F3792_ = ~new_F3759_ & ~new_F3795_;
  assign new_F3793_ = F3742 | new_F3759_;
  assign new_F3794_ = F3742 | F3743;
  assign new_F3795_ = new_F3759_ & new_F3796_;
  assign new_F3796_ = ~F3741 | ~new_F3766_;
  assign new_F3797_ = new_F3774_ & new_F3794_;
  assign new_F3798_ = ~new_F3774_ & ~new_F3794_;
  assign new_F3799_ = new_F3803_ | new_F3804_;
  assign new_F3800_ = ~F3745 & new_F3759_;
  assign new_F3801_ = new_F3805_ | new_F3806_;
  assign new_F3802_ = F3745 & new_F3759_;
  assign new_F3803_ = ~F3745 & ~new_F3759_;
  assign new_F3804_ = F3745 & ~new_F3759_;
  assign new_F3805_ = F3745 & ~new_F3759_;
  assign new_F3806_ = ~F3745 & new_F3759_;
  assign new_F3813_ = new_F3820_ & new_F3819_;
  assign new_F3814_ = new_F3822_ | new_F3821_;
  assign new_F3815_ = new_F3824_ | new_F3823_;
  assign new_F3816_ = new_F3826_ & new_F3825_;
  assign new_F3817_ = new_F3826_ & new_F3827_;
  assign new_F3818_ = new_F3819_ | new_F3828_;
  assign new_F3819_ = F3808 | new_F3831_;
  assign new_F3820_ = new_F3830_ | new_F3829_;
  assign new_F3821_ = new_F3835_ & new_F3834_;
  assign new_F3822_ = new_F3833_ & new_F3832_;
  assign new_F3823_ = new_F3838_ | new_F3837_;
  assign new_F3824_ = new_F3833_ & new_F3836_;
  assign new_F3825_ = F3808 | new_F3841_;
  assign new_F3826_ = new_F3840_ | new_F3839_;
  assign new_F3827_ = new_F3843_ | new_F3842_;
  assign new_F3828_ = ~new_F3819_ & new_F3845_;
  assign new_F3829_ = ~new_F3821_ & new_F3833_;
  assign new_F3830_ = new_F3821_ & ~new_F3833_;
  assign new_F3831_ = F3807 & ~F3808;
  assign new_F3832_ = ~new_F3854_ | ~new_F3855_;
  assign new_F3833_ = new_F3847_ | new_F3849_;
  assign new_F3834_ = new_F3857_ | new_F3856_;
  assign new_F3835_ = new_F3851_ | new_F3850_;
  assign new_F3836_ = ~new_F3859_ | ~new_F3858_;
  assign new_F3837_ = ~new_F3860_ & new_F3861_;
  assign new_F3838_ = new_F3860_ & ~new_F3861_;
  assign new_F3839_ = ~F3807 & F3808;
  assign new_F3840_ = F3807 & ~F3808;
  assign new_F3841_ = ~new_F3823_ | new_F3833_;
  assign new_F3842_ = new_F3823_ & new_F3833_;
  assign new_F3843_ = ~new_F3823_ & ~new_F3833_;
  assign new_F3844_ = new_F3865_ | new_F3864_;
  assign new_F3845_ = F3811 | new_F3844_;
  assign new_F3846_ = new_F3869_ | new_F3868_;
  assign new_F3847_ = ~F3811 & new_F3846_;
  assign new_F3848_ = new_F3867_ | new_F3866_;
  assign new_F3849_ = F3811 & new_F3848_;
  assign new_F3850_ = F3809 & ~new_F3819_;
  assign new_F3851_ = ~F3809 & new_F3819_;
  assign new_F3852_ = ~F3808 | ~new_F3833_;
  assign new_F3853_ = new_F3819_ & new_F3852_;
  assign new_F3854_ = ~new_F3819_ & ~new_F3853_;
  assign new_F3855_ = new_F3819_ | new_F3852_;
  assign new_F3856_ = ~F3809 & F3810;
  assign new_F3857_ = F3809 & ~F3810;
  assign new_F3858_ = new_F3826_ | new_F3863_;
  assign new_F3859_ = ~new_F3826_ & ~new_F3862_;
  assign new_F3860_ = F3809 | new_F3826_;
  assign new_F3861_ = F3809 | F3810;
  assign new_F3862_ = new_F3826_ & new_F3863_;
  assign new_F3863_ = ~F3808 | ~new_F3833_;
  assign new_F3864_ = new_F3841_ & new_F3861_;
  assign new_F3865_ = ~new_F3841_ & ~new_F3861_;
  assign new_F3866_ = new_F3870_ | new_F3871_;
  assign new_F3867_ = ~F3812 & new_F3826_;
  assign new_F3868_ = new_F3872_ | new_F3873_;
  assign new_F3869_ = F3812 & new_F3826_;
  assign new_F3870_ = ~F3812 & ~new_F3826_;
  assign new_F3871_ = F3812 & ~new_F3826_;
  assign new_F3872_ = F3812 & ~new_F3826_;
  assign new_F3873_ = ~F3812 & new_F3826_;
  assign new_F3880_ = new_F3887_ & new_F3886_;
  assign new_F3881_ = new_F3889_ | new_F3888_;
  assign new_F3882_ = new_F3891_ | new_F3890_;
  assign new_F3883_ = new_F3893_ & new_F3892_;
  assign new_F3884_ = new_F3893_ & new_F3894_;
  assign new_F3885_ = new_F3886_ | new_F3895_;
  assign new_F3886_ = F3875 | new_F3898_;
  assign new_F3887_ = new_F3897_ | new_F3896_;
  assign new_F3888_ = new_F3902_ & new_F3901_;
  assign new_F3889_ = new_F3900_ & new_F3899_;
  assign new_F3890_ = new_F3905_ | new_F3904_;
  assign new_F3891_ = new_F3900_ & new_F3903_;
  assign new_F3892_ = F3875 | new_F3908_;
  assign new_F3893_ = new_F3907_ | new_F3906_;
  assign new_F3894_ = new_F3910_ | new_F3909_;
  assign new_F3895_ = ~new_F3886_ & new_F3912_;
  assign new_F3896_ = ~new_F3888_ & new_F3900_;
  assign new_F3897_ = new_F3888_ & ~new_F3900_;
  assign new_F3898_ = F3874 & ~F3875;
  assign new_F3899_ = ~new_F3921_ | ~new_F3922_;
  assign new_F3900_ = new_F3914_ | new_F3916_;
  assign new_F3901_ = new_F3924_ | new_F3923_;
  assign new_F3902_ = new_F3918_ | new_F3917_;
  assign new_F3903_ = ~new_F3926_ | ~new_F3925_;
  assign new_F3904_ = ~new_F3927_ & new_F3928_;
  assign new_F3905_ = new_F3927_ & ~new_F3928_;
  assign new_F3906_ = ~F3874 & F3875;
  assign new_F3907_ = F3874 & ~F3875;
  assign new_F3908_ = ~new_F3890_ | new_F3900_;
  assign new_F3909_ = new_F3890_ & new_F3900_;
  assign new_F3910_ = ~new_F3890_ & ~new_F3900_;
  assign new_F3911_ = new_F3932_ | new_F3931_;
  assign new_F3912_ = F3878 | new_F3911_;
  assign new_F3913_ = new_F3936_ | new_F3935_;
  assign new_F3914_ = ~F3878 & new_F3913_;
  assign new_F3915_ = new_F3934_ | new_F3933_;
  assign new_F3916_ = F3878 & new_F3915_;
  assign new_F3917_ = F3876 & ~new_F3886_;
  assign new_F3918_ = ~F3876 & new_F3886_;
  assign new_F3919_ = ~F3875 | ~new_F3900_;
  assign new_F3920_ = new_F3886_ & new_F3919_;
  assign new_F3921_ = ~new_F3886_ & ~new_F3920_;
  assign new_F3922_ = new_F3886_ | new_F3919_;
  assign new_F3923_ = ~F3876 & F3877;
  assign new_F3924_ = F3876 & ~F3877;
  assign new_F3925_ = new_F3893_ | new_F3930_;
  assign new_F3926_ = ~new_F3893_ & ~new_F3929_;
  assign new_F3927_ = F3876 | new_F3893_;
  assign new_F3928_ = F3876 | F3877;
  assign new_F3929_ = new_F3893_ & new_F3930_;
  assign new_F3930_ = ~F3875 | ~new_F3900_;
  assign new_F3931_ = new_F3908_ & new_F3928_;
  assign new_F3932_ = ~new_F3908_ & ~new_F3928_;
  assign new_F3933_ = new_F3937_ | new_F3938_;
  assign new_F3934_ = ~F3879 & new_F3893_;
  assign new_F3935_ = new_F3939_ | new_F3940_;
  assign new_F3936_ = F3879 & new_F3893_;
  assign new_F3937_ = ~F3879 & ~new_F3893_;
  assign new_F3938_ = F3879 & ~new_F3893_;
  assign new_F3939_ = F3879 & ~new_F3893_;
  assign new_F3940_ = ~F3879 & new_F3893_;
  assign new_F3947_ = new_F3954_ & new_F3953_;
  assign new_F3948_ = new_F3956_ | new_F3955_;
  assign new_F3949_ = new_F3958_ | new_F3957_;
  assign new_F3950_ = new_F3960_ & new_F3959_;
  assign new_F3951_ = new_F3960_ & new_F3961_;
  assign new_F3952_ = new_F3953_ | new_F3962_;
  assign new_F3953_ = F3942 | new_F3965_;
  assign new_F3954_ = new_F3964_ | new_F3963_;
  assign new_F3955_ = new_F3969_ & new_F3968_;
  assign new_F3956_ = new_F3967_ & new_F3966_;
  assign new_F3957_ = new_F3972_ | new_F3971_;
  assign new_F3958_ = new_F3967_ & new_F3970_;
  assign new_F3959_ = F3942 | new_F3975_;
  assign new_F3960_ = new_F3974_ | new_F3973_;
  assign new_F3961_ = new_F3977_ | new_F3976_;
  assign new_F3962_ = ~new_F3953_ & new_F3979_;
  assign new_F3963_ = ~new_F3955_ & new_F3967_;
  assign new_F3964_ = new_F3955_ & ~new_F3967_;
  assign new_F3965_ = F3941 & ~F3942;
  assign new_F3966_ = ~new_F3988_ | ~new_F3989_;
  assign new_F3967_ = new_F3981_ | new_F3983_;
  assign new_F3968_ = new_F3991_ | new_F3990_;
  assign new_F3969_ = new_F3985_ | new_F3984_;
  assign new_F3970_ = ~new_F3993_ | ~new_F3992_;
  assign new_F3971_ = ~new_F3994_ & new_F3995_;
  assign new_F3972_ = new_F3994_ & ~new_F3995_;
  assign new_F3973_ = ~F3941 & F3942;
  assign new_F3974_ = F3941 & ~F3942;
  assign new_F3975_ = ~new_F3957_ | new_F3967_;
  assign new_F3976_ = new_F3957_ & new_F3967_;
  assign new_F3977_ = ~new_F3957_ & ~new_F3967_;
  assign new_F3978_ = new_F3999_ | new_F3998_;
  assign new_F3979_ = F3945 | new_F3978_;
  assign new_F3980_ = new_F4003_ | new_F4002_;
  assign new_F3981_ = ~F3945 & new_F3980_;
  assign new_F3982_ = new_F4001_ | new_F4000_;
  assign new_F3983_ = F3945 & new_F3982_;
  assign new_F3984_ = F3943 & ~new_F3953_;
  assign new_F3985_ = ~F3943 & new_F3953_;
  assign new_F3986_ = ~F3942 | ~new_F3967_;
  assign new_F3987_ = new_F3953_ & new_F3986_;
  assign new_F3988_ = ~new_F3953_ & ~new_F3987_;
  assign new_F3989_ = new_F3953_ | new_F3986_;
  assign new_F3990_ = ~F3943 & F3944;
  assign new_F3991_ = F3943 & ~F3944;
  assign new_F3992_ = new_F3960_ | new_F3997_;
  assign new_F3993_ = ~new_F3960_ & ~new_F3996_;
  assign new_F3994_ = F3943 | new_F3960_;
  assign new_F3995_ = F3943 | F3944;
  assign new_F3996_ = new_F3960_ & new_F3997_;
  assign new_F3997_ = ~F3942 | ~new_F3967_;
  assign new_F3998_ = new_F3975_ & new_F3995_;
  assign new_F3999_ = ~new_F3975_ & ~new_F3995_;
  assign new_F4000_ = new_F4004_ | new_F4005_;
  assign new_F4001_ = ~F3946 & new_F3960_;
  assign new_F4002_ = new_F4006_ | new_F4007_;
  assign new_F4003_ = F3946 & new_F3960_;
  assign new_F4004_ = ~F3946 & ~new_F3960_;
  assign new_F4005_ = F3946 & ~new_F3960_;
  assign new_F4006_ = F3946 & ~new_F3960_;
  assign new_F4007_ = ~F3946 & new_F3960_;
  assign new_F4014_ = new_F4021_ & new_F4020_;
  assign new_F4015_ = new_F4023_ | new_F4022_;
  assign new_F4016_ = new_F4025_ | new_F4024_;
  assign new_F4017_ = new_F4027_ & new_F4026_;
  assign new_F4018_ = new_F4027_ & new_F4028_;
  assign new_F4019_ = new_F4020_ | new_F4029_;
  assign new_F4020_ = F4009 | new_F4032_;
  assign new_F4021_ = new_F4031_ | new_F4030_;
  assign new_F4022_ = new_F4036_ & new_F4035_;
  assign new_F4023_ = new_F4034_ & new_F4033_;
  assign new_F4024_ = new_F4039_ | new_F4038_;
  assign new_F4025_ = new_F4034_ & new_F4037_;
  assign new_F4026_ = F4009 | new_F4042_;
  assign new_F4027_ = new_F4041_ | new_F4040_;
  assign new_F4028_ = new_F4044_ | new_F4043_;
  assign new_F4029_ = ~new_F4020_ & new_F4046_;
  assign new_F4030_ = ~new_F4022_ & new_F4034_;
  assign new_F4031_ = new_F4022_ & ~new_F4034_;
  assign new_F4032_ = F4008 & ~F4009;
  assign new_F4033_ = ~new_F4055_ | ~new_F4056_;
  assign new_F4034_ = new_F4048_ | new_F4050_;
  assign new_F4035_ = new_F4058_ | new_F4057_;
  assign new_F4036_ = new_F4052_ | new_F4051_;
  assign new_F4037_ = ~new_F4060_ | ~new_F4059_;
  assign new_F4038_ = ~new_F4061_ & new_F4062_;
  assign new_F4039_ = new_F4061_ & ~new_F4062_;
  assign new_F4040_ = ~F4008 & F4009;
  assign new_F4041_ = F4008 & ~F4009;
  assign new_F4042_ = ~new_F4024_ | new_F4034_;
  assign new_F4043_ = new_F4024_ & new_F4034_;
  assign new_F4044_ = ~new_F4024_ & ~new_F4034_;
  assign new_F4045_ = new_F4066_ | new_F4065_;
  assign new_F4046_ = F4012 | new_F4045_;
  assign new_F4047_ = new_F4070_ | new_F4069_;
  assign new_F4048_ = ~F4012 & new_F4047_;
  assign new_F4049_ = new_F4068_ | new_F4067_;
  assign new_F4050_ = F4012 & new_F4049_;
  assign new_F4051_ = F4010 & ~new_F4020_;
  assign new_F4052_ = ~F4010 & new_F4020_;
  assign new_F4053_ = ~F4009 | ~new_F4034_;
  assign new_F4054_ = new_F4020_ & new_F4053_;
  assign new_F4055_ = ~new_F4020_ & ~new_F4054_;
  assign new_F4056_ = new_F4020_ | new_F4053_;
  assign new_F4057_ = ~F4010 & F4011;
  assign new_F4058_ = F4010 & ~F4011;
  assign new_F4059_ = new_F4027_ | new_F4064_;
  assign new_F4060_ = ~new_F4027_ & ~new_F4063_;
  assign new_F4061_ = F4010 | new_F4027_;
  assign new_F4062_ = F4010 | F4011;
  assign new_F4063_ = new_F4027_ & new_F4064_;
  assign new_F4064_ = ~F4009 | ~new_F4034_;
  assign new_F4065_ = new_F4042_ & new_F4062_;
  assign new_F4066_ = ~new_F4042_ & ~new_F4062_;
  assign new_F4067_ = new_F4071_ | new_F4072_;
  assign new_F4068_ = ~F4013 & new_F4027_;
  assign new_F4069_ = new_F4073_ | new_F4074_;
  assign new_F4070_ = F4013 & new_F4027_;
  assign new_F4071_ = ~F4013 & ~new_F4027_;
  assign new_F4072_ = F4013 & ~new_F4027_;
  assign new_F4073_ = F4013 & ~new_F4027_;
  assign new_F4074_ = ~F4013 & new_F4027_;
  assign new_F4081_ = new_F4088_ & new_F4087_;
  assign new_F4082_ = new_F4090_ | new_F4089_;
  assign new_F4083_ = new_F4092_ | new_F4091_;
  assign new_F4084_ = new_F4094_ & new_F4093_;
  assign new_F4085_ = new_F4094_ & new_F4095_;
  assign new_F4086_ = new_F4087_ | new_F4096_;
  assign new_F4087_ = F4076 | new_F4099_;
  assign new_F4088_ = new_F4098_ | new_F4097_;
  assign new_F4089_ = new_F4103_ & new_F4102_;
  assign new_F4090_ = new_F4101_ & new_F4100_;
  assign new_F4091_ = new_F4106_ | new_F4105_;
  assign new_F4092_ = new_F4101_ & new_F4104_;
  assign new_F4093_ = F4076 | new_F4109_;
  assign new_F4094_ = new_F4108_ | new_F4107_;
  assign new_F4095_ = new_F4111_ | new_F4110_;
  assign new_F4096_ = ~new_F4087_ & new_F4113_;
  assign new_F4097_ = ~new_F4089_ & new_F4101_;
  assign new_F4098_ = new_F4089_ & ~new_F4101_;
  assign new_F4099_ = F4075 & ~F4076;
  assign new_F4100_ = ~new_F4122_ | ~new_F4123_;
  assign new_F4101_ = new_F4115_ | new_F4117_;
  assign new_F4102_ = new_F4125_ | new_F4124_;
  assign new_F4103_ = new_F4119_ | new_F4118_;
  assign new_F4104_ = ~new_F4127_ | ~new_F4126_;
  assign new_F4105_ = ~new_F4128_ & new_F4129_;
  assign new_F4106_ = new_F4128_ & ~new_F4129_;
  assign new_F4107_ = ~F4075 & F4076;
  assign new_F4108_ = F4075 & ~F4076;
  assign new_F4109_ = ~new_F4091_ | new_F4101_;
  assign new_F4110_ = new_F4091_ & new_F4101_;
  assign new_F4111_ = ~new_F4091_ & ~new_F4101_;
  assign new_F4112_ = new_F4133_ | new_F4132_;
  assign new_F4113_ = F4079 | new_F4112_;
  assign new_F4114_ = new_F4137_ | new_F4136_;
  assign new_F4115_ = ~F4079 & new_F4114_;
  assign new_F4116_ = new_F4135_ | new_F4134_;
  assign new_F4117_ = F4079 & new_F4116_;
  assign new_F4118_ = F4077 & ~new_F4087_;
  assign new_F4119_ = ~F4077 & new_F4087_;
  assign new_F4120_ = ~F4076 | ~new_F4101_;
  assign new_F4121_ = new_F4087_ & new_F4120_;
  assign new_F4122_ = ~new_F4087_ & ~new_F4121_;
  assign new_F4123_ = new_F4087_ | new_F4120_;
  assign new_F4124_ = ~F4077 & F4078;
  assign new_F4125_ = F4077 & ~F4078;
  assign new_F4126_ = new_F4094_ | new_F4131_;
  assign new_F4127_ = ~new_F4094_ & ~new_F4130_;
  assign new_F4128_ = F4077 | new_F4094_;
  assign new_F4129_ = F4077 | F4078;
  assign new_F4130_ = new_F4094_ & new_F4131_;
  assign new_F4131_ = ~F4076 | ~new_F4101_;
  assign new_F4132_ = new_F4109_ & new_F4129_;
  assign new_F4133_ = ~new_F4109_ & ~new_F4129_;
  assign new_F4134_ = new_F4138_ | new_F4139_;
  assign new_F4135_ = ~F4080 & new_F4094_;
  assign new_F4136_ = new_F4140_ | new_F4141_;
  assign new_F4137_ = F4080 & new_F4094_;
  assign new_F4138_ = ~F4080 & ~new_F4094_;
  assign new_F4139_ = F4080 & ~new_F4094_;
  assign new_F4140_ = F4080 & ~new_F4094_;
  assign new_F4141_ = ~F4080 & new_F4094_;
  assign new_F4148_ = new_F4155_ & new_F4154_;
  assign new_F4149_ = new_F4157_ | new_F4156_;
  assign new_F4150_ = new_F4159_ | new_F4158_;
  assign new_F4151_ = new_F4161_ & new_F4160_;
  assign new_F4152_ = new_F4161_ & new_F4162_;
  assign new_F4153_ = new_F4154_ | new_F4163_;
  assign new_F4154_ = F4143 | new_F4166_;
  assign new_F4155_ = new_F4165_ | new_F4164_;
  assign new_F4156_ = new_F4170_ & new_F4169_;
  assign new_F4157_ = new_F4168_ & new_F4167_;
  assign new_F4158_ = new_F4173_ | new_F4172_;
  assign new_F4159_ = new_F4168_ & new_F4171_;
  assign new_F4160_ = F4143 | new_F4176_;
  assign new_F4161_ = new_F4175_ | new_F4174_;
  assign new_F4162_ = new_F4178_ | new_F4177_;
  assign new_F4163_ = ~new_F4154_ & new_F4180_;
  assign new_F4164_ = ~new_F4156_ & new_F4168_;
  assign new_F4165_ = new_F4156_ & ~new_F4168_;
  assign new_F4166_ = F4142 & ~F4143;
  assign new_F4167_ = ~new_F4189_ | ~new_F4190_;
  assign new_F4168_ = new_F4182_ | new_F4184_;
  assign new_F4169_ = new_F4192_ | new_F4191_;
  assign new_F4170_ = new_F4186_ | new_F4185_;
  assign new_F4171_ = ~new_F4194_ | ~new_F4193_;
  assign new_F4172_ = ~new_F4195_ & new_F4196_;
  assign new_F4173_ = new_F4195_ & ~new_F4196_;
  assign new_F4174_ = ~F4142 & F4143;
  assign new_F4175_ = F4142 & ~F4143;
  assign new_F4176_ = ~new_F4158_ | new_F4168_;
  assign new_F4177_ = new_F4158_ & new_F4168_;
  assign new_F4178_ = ~new_F4158_ & ~new_F4168_;
  assign new_F4179_ = new_F4200_ | new_F4199_;
  assign new_F4180_ = F4146 | new_F4179_;
  assign new_F4181_ = new_F4204_ | new_F4203_;
  assign new_F4182_ = ~F4146 & new_F4181_;
  assign new_F4183_ = new_F4202_ | new_F4201_;
  assign new_F4184_ = F4146 & new_F4183_;
  assign new_F4185_ = F4144 & ~new_F4154_;
  assign new_F4186_ = ~F4144 & new_F4154_;
  assign new_F4187_ = ~F4143 | ~new_F4168_;
  assign new_F4188_ = new_F4154_ & new_F4187_;
  assign new_F4189_ = ~new_F4154_ & ~new_F4188_;
  assign new_F4190_ = new_F4154_ | new_F4187_;
  assign new_F4191_ = ~F4144 & F4145;
  assign new_F4192_ = F4144 & ~F4145;
  assign new_F4193_ = new_F4161_ | new_F4198_;
  assign new_F4194_ = ~new_F4161_ & ~new_F4197_;
  assign new_F4195_ = F4144 | new_F4161_;
  assign new_F4196_ = F4144 | F4145;
  assign new_F4197_ = new_F4161_ & new_F4198_;
  assign new_F4198_ = ~F4143 | ~new_F4168_;
  assign new_F4199_ = new_F4176_ & new_F4196_;
  assign new_F4200_ = ~new_F4176_ & ~new_F4196_;
  assign new_F4201_ = new_F4205_ | new_F4206_;
  assign new_F4202_ = ~F4147 & new_F4161_;
  assign new_F4203_ = new_F4207_ | new_F4208_;
  assign new_F4204_ = F4147 & new_F4161_;
  assign new_F4205_ = ~F4147 & ~new_F4161_;
  assign new_F4206_ = F4147 & ~new_F4161_;
  assign new_F4207_ = F4147 & ~new_F4161_;
  assign new_F4208_ = ~F4147 & new_F4161_;
  assign new_F4215_ = new_F4222_ & new_F4221_;
  assign new_F4216_ = new_F4224_ | new_F4223_;
  assign new_F4217_ = new_F4226_ | new_F4225_;
  assign new_F4218_ = new_F4228_ & new_F4227_;
  assign new_F4219_ = new_F4228_ & new_F4229_;
  assign new_F4220_ = new_F4221_ | new_F4230_;
  assign new_F4221_ = F4210 | new_F4233_;
  assign new_F4222_ = new_F4232_ | new_F4231_;
  assign new_F4223_ = new_F4237_ & new_F4236_;
  assign new_F4224_ = new_F4235_ & new_F4234_;
  assign new_F4225_ = new_F4240_ | new_F4239_;
  assign new_F4226_ = new_F4235_ & new_F4238_;
  assign new_F4227_ = F4210 | new_F4243_;
  assign new_F4228_ = new_F4242_ | new_F4241_;
  assign new_F4229_ = new_F4245_ | new_F4244_;
  assign new_F4230_ = ~new_F4221_ & new_F4247_;
  assign new_F4231_ = ~new_F4223_ & new_F4235_;
  assign new_F4232_ = new_F4223_ & ~new_F4235_;
  assign new_F4233_ = F4209 & ~F4210;
  assign new_F4234_ = ~new_F4256_ | ~new_F4257_;
  assign new_F4235_ = new_F4249_ | new_F4251_;
  assign new_F4236_ = new_F4259_ | new_F4258_;
  assign new_F4237_ = new_F4253_ | new_F4252_;
  assign new_F4238_ = ~new_F4261_ | ~new_F4260_;
  assign new_F4239_ = ~new_F4262_ & new_F4263_;
  assign new_F4240_ = new_F4262_ & ~new_F4263_;
  assign new_F4241_ = ~F4209 & F4210;
  assign new_F4242_ = F4209 & ~F4210;
  assign new_F4243_ = ~new_F4225_ | new_F4235_;
  assign new_F4244_ = new_F4225_ & new_F4235_;
  assign new_F4245_ = ~new_F4225_ & ~new_F4235_;
  assign new_F4246_ = new_F4267_ | new_F4266_;
  assign new_F4247_ = F4213 | new_F4246_;
  assign new_F4248_ = new_F4271_ | new_F4270_;
  assign new_F4249_ = ~F4213 & new_F4248_;
  assign new_F4250_ = new_F4269_ | new_F4268_;
  assign new_F4251_ = F4213 & new_F4250_;
  assign new_F4252_ = F4211 & ~new_F4221_;
  assign new_F4253_ = ~F4211 & new_F4221_;
  assign new_F4254_ = ~F4210 | ~new_F4235_;
  assign new_F4255_ = new_F4221_ & new_F4254_;
  assign new_F4256_ = ~new_F4221_ & ~new_F4255_;
  assign new_F4257_ = new_F4221_ | new_F4254_;
  assign new_F4258_ = ~F4211 & F4212;
  assign new_F4259_ = F4211 & ~F4212;
  assign new_F4260_ = new_F4228_ | new_F4265_;
  assign new_F4261_ = ~new_F4228_ & ~new_F4264_;
  assign new_F4262_ = F4211 | new_F4228_;
  assign new_F4263_ = F4211 | F4212;
  assign new_F4264_ = new_F4228_ & new_F4265_;
  assign new_F4265_ = ~F4210 | ~new_F4235_;
  assign new_F4266_ = new_F4243_ & new_F4263_;
  assign new_F4267_ = ~new_F4243_ & ~new_F4263_;
  assign new_F4268_ = new_F4272_ | new_F4273_;
  assign new_F4269_ = ~F4214 & new_F4228_;
  assign new_F4270_ = new_F4274_ | new_F4275_;
  assign new_F4271_ = F4214 & new_F4228_;
  assign new_F4272_ = ~F4214 & ~new_F4228_;
  assign new_F4273_ = F4214 & ~new_F4228_;
  assign new_F4274_ = F4214 & ~new_F4228_;
  assign new_F4275_ = ~F4214 & new_F4228_;
  assign new_F4282_ = new_F4289_ & new_F4288_;
  assign new_F4283_ = new_F4291_ | new_F4290_;
  assign new_F4284_ = new_F4293_ | new_F4292_;
  assign new_F4285_ = new_F4295_ & new_F4294_;
  assign new_F4286_ = new_F4295_ & new_F4296_;
  assign new_F4287_ = new_F4288_ | new_F4297_;
  assign new_F4288_ = F4277 | new_F4300_;
  assign new_F4289_ = new_F4299_ | new_F4298_;
  assign new_F4290_ = new_F4304_ & new_F4303_;
  assign new_F4291_ = new_F4302_ & new_F4301_;
  assign new_F4292_ = new_F4307_ | new_F4306_;
  assign new_F4293_ = new_F4302_ & new_F4305_;
  assign new_F4294_ = F4277 | new_F4310_;
  assign new_F4295_ = new_F4309_ | new_F4308_;
  assign new_F4296_ = new_F4312_ | new_F4311_;
  assign new_F4297_ = ~new_F4288_ & new_F4314_;
  assign new_F4298_ = ~new_F4290_ & new_F4302_;
  assign new_F4299_ = new_F4290_ & ~new_F4302_;
  assign new_F4300_ = F4276 & ~F4277;
  assign new_F4301_ = ~new_F4323_ | ~new_F4324_;
  assign new_F4302_ = new_F4316_ | new_F4318_;
  assign new_F4303_ = new_F4326_ | new_F4325_;
  assign new_F4304_ = new_F4320_ | new_F4319_;
  assign new_F4305_ = ~new_F4328_ | ~new_F4327_;
  assign new_F4306_ = ~new_F4329_ & new_F4330_;
  assign new_F4307_ = new_F4329_ & ~new_F4330_;
  assign new_F4308_ = ~F4276 & F4277;
  assign new_F4309_ = F4276 & ~F4277;
  assign new_F4310_ = ~new_F4292_ | new_F4302_;
  assign new_F4311_ = new_F4292_ & new_F4302_;
  assign new_F4312_ = ~new_F4292_ & ~new_F4302_;
  assign new_F4313_ = new_F4334_ | new_F4333_;
  assign new_F4314_ = F4280 | new_F4313_;
  assign new_F4315_ = new_F4338_ | new_F4337_;
  assign new_F4316_ = ~F4280 & new_F4315_;
  assign new_F4317_ = new_F4336_ | new_F4335_;
  assign new_F4318_ = F4280 & new_F4317_;
  assign new_F4319_ = F4278 & ~new_F4288_;
  assign new_F4320_ = ~F4278 & new_F4288_;
  assign new_F4321_ = ~F4277 | ~new_F4302_;
  assign new_F4322_ = new_F4288_ & new_F4321_;
  assign new_F4323_ = ~new_F4288_ & ~new_F4322_;
  assign new_F4324_ = new_F4288_ | new_F4321_;
  assign new_F4325_ = ~F4278 & F4279;
  assign new_F4326_ = F4278 & ~F4279;
  assign new_F4327_ = new_F4295_ | new_F4332_;
  assign new_F4328_ = ~new_F4295_ & ~new_F4331_;
  assign new_F4329_ = F4278 | new_F4295_;
  assign new_F4330_ = F4278 | F4279;
  assign new_F4331_ = new_F4295_ & new_F4332_;
  assign new_F4332_ = ~F4277 | ~new_F4302_;
  assign new_F4333_ = new_F4310_ & new_F4330_;
  assign new_F4334_ = ~new_F4310_ & ~new_F4330_;
  assign new_F4335_ = new_F4339_ | new_F4340_;
  assign new_F4336_ = ~F4281 & new_F4295_;
  assign new_F4337_ = new_F4341_ | new_F4342_;
  assign new_F4338_ = F4281 & new_F4295_;
  assign new_F4339_ = ~F4281 & ~new_F4295_;
  assign new_F4340_ = F4281 & ~new_F4295_;
  assign new_F4341_ = F4281 & ~new_F4295_;
  assign new_F4342_ = ~F4281 & new_F4295_;
  assign new_F4349_ = new_F4356_ & new_F4355_;
  assign new_F4350_ = new_F4358_ | new_F4357_;
  assign new_F4351_ = new_F4360_ | new_F4359_;
  assign new_F4352_ = new_F4362_ & new_F4361_;
  assign new_F4353_ = new_F4362_ & new_F4363_;
  assign new_F4354_ = new_F4355_ | new_F4364_;
  assign new_F4355_ = F4344 | new_F4367_;
  assign new_F4356_ = new_F4366_ | new_F4365_;
  assign new_F4357_ = new_F4371_ & new_F4370_;
  assign new_F4358_ = new_F4369_ & new_F4368_;
  assign new_F4359_ = new_F4374_ | new_F4373_;
  assign new_F4360_ = new_F4369_ & new_F4372_;
  assign new_F4361_ = F4344 | new_F4377_;
  assign new_F4362_ = new_F4376_ | new_F4375_;
  assign new_F4363_ = new_F4379_ | new_F4378_;
  assign new_F4364_ = ~new_F4355_ & new_F4381_;
  assign new_F4365_ = ~new_F4357_ & new_F4369_;
  assign new_F4366_ = new_F4357_ & ~new_F4369_;
  assign new_F4367_ = F4343 & ~F4344;
  assign new_F4368_ = ~new_F4390_ | ~new_F4391_;
  assign new_F4369_ = new_F4383_ | new_F4385_;
  assign new_F4370_ = new_F4393_ | new_F4392_;
  assign new_F4371_ = new_F4387_ | new_F4386_;
  assign new_F4372_ = ~new_F4395_ | ~new_F4394_;
  assign new_F4373_ = ~new_F4396_ & new_F4397_;
  assign new_F4374_ = new_F4396_ & ~new_F4397_;
  assign new_F4375_ = ~F4343 & F4344;
  assign new_F4376_ = F4343 & ~F4344;
  assign new_F4377_ = ~new_F4359_ | new_F4369_;
  assign new_F4378_ = new_F4359_ & new_F4369_;
  assign new_F4379_ = ~new_F4359_ & ~new_F4369_;
  assign new_F4380_ = new_F4401_ | new_F4400_;
  assign new_F4381_ = F4347 | new_F4380_;
  assign new_F4382_ = new_F4405_ | new_F4404_;
  assign new_F4383_ = ~F4347 & new_F4382_;
  assign new_F4384_ = new_F4403_ | new_F4402_;
  assign new_F4385_ = F4347 & new_F4384_;
  assign new_F4386_ = F4345 & ~new_F4355_;
  assign new_F4387_ = ~F4345 & new_F4355_;
  assign new_F4388_ = ~F4344 | ~new_F4369_;
  assign new_F4389_ = new_F4355_ & new_F4388_;
  assign new_F4390_ = ~new_F4355_ & ~new_F4389_;
  assign new_F4391_ = new_F4355_ | new_F4388_;
  assign new_F4392_ = ~F4345 & F4346;
  assign new_F4393_ = F4345 & ~F4346;
  assign new_F4394_ = new_F4362_ | new_F4399_;
  assign new_F4395_ = ~new_F4362_ & ~new_F4398_;
  assign new_F4396_ = F4345 | new_F4362_;
  assign new_F4397_ = F4345 | F4346;
  assign new_F4398_ = new_F4362_ & new_F4399_;
  assign new_F4399_ = ~F4344 | ~new_F4369_;
  assign new_F4400_ = new_F4377_ & new_F4397_;
  assign new_F4401_ = ~new_F4377_ & ~new_F4397_;
  assign new_F4402_ = new_F4406_ | new_F4407_;
  assign new_F4403_ = ~F4348 & new_F4362_;
  assign new_F4404_ = new_F4408_ | new_F4409_;
  assign new_F4405_ = F4348 & new_F4362_;
  assign new_F4406_ = ~F4348 & ~new_F4362_;
  assign new_F4407_ = F4348 & ~new_F4362_;
  assign new_F4408_ = F4348 & ~new_F4362_;
  assign new_F4409_ = ~F4348 & new_F4362_;
  assign new_F4416_ = new_F4423_ & new_F4422_;
  assign new_F4417_ = new_F4425_ | new_F4424_;
  assign new_F4418_ = new_F4427_ | new_F4426_;
  assign new_F4419_ = new_F4429_ & new_F4428_;
  assign new_F4420_ = new_F4429_ & new_F4430_;
  assign new_F4421_ = new_F4422_ | new_F4431_;
  assign new_F4422_ = F4411 | new_F4434_;
  assign new_F4423_ = new_F4433_ | new_F4432_;
  assign new_F4424_ = new_F4438_ & new_F4437_;
  assign new_F4425_ = new_F4436_ & new_F4435_;
  assign new_F4426_ = new_F4441_ | new_F4440_;
  assign new_F4427_ = new_F4436_ & new_F4439_;
  assign new_F4428_ = F4411 | new_F4444_;
  assign new_F4429_ = new_F4443_ | new_F4442_;
  assign new_F4430_ = new_F4446_ | new_F4445_;
  assign new_F4431_ = ~new_F4422_ & new_F4448_;
  assign new_F4432_ = ~new_F4424_ & new_F4436_;
  assign new_F4433_ = new_F4424_ & ~new_F4436_;
  assign new_F4434_ = F4410 & ~F4411;
  assign new_F4435_ = ~new_F4457_ | ~new_F4458_;
  assign new_F4436_ = new_F4450_ | new_F4452_;
  assign new_F4437_ = new_F4460_ | new_F4459_;
  assign new_F4438_ = new_F4454_ | new_F4453_;
  assign new_F4439_ = ~new_F4462_ | ~new_F4461_;
  assign new_F4440_ = ~new_F4463_ & new_F4464_;
  assign new_F4441_ = new_F4463_ & ~new_F4464_;
  assign new_F4442_ = ~F4410 & F4411;
  assign new_F4443_ = F4410 & ~F4411;
  assign new_F4444_ = ~new_F4426_ | new_F4436_;
  assign new_F4445_ = new_F4426_ & new_F4436_;
  assign new_F4446_ = ~new_F4426_ & ~new_F4436_;
  assign new_F4447_ = new_F4468_ | new_F4467_;
  assign new_F4448_ = F4414 | new_F4447_;
  assign new_F4449_ = new_F4472_ | new_F4471_;
  assign new_F4450_ = ~F4414 & new_F4449_;
  assign new_F4451_ = new_F4470_ | new_F4469_;
  assign new_F4452_ = F4414 & new_F4451_;
  assign new_F4453_ = F4412 & ~new_F4422_;
  assign new_F4454_ = ~F4412 & new_F4422_;
  assign new_F4455_ = ~F4411 | ~new_F4436_;
  assign new_F4456_ = new_F4422_ & new_F4455_;
  assign new_F4457_ = ~new_F4422_ & ~new_F4456_;
  assign new_F4458_ = new_F4422_ | new_F4455_;
  assign new_F4459_ = ~F4412 & F4413;
  assign new_F4460_ = F4412 & ~F4413;
  assign new_F4461_ = new_F4429_ | new_F4466_;
  assign new_F4462_ = ~new_F4429_ & ~new_F4465_;
  assign new_F4463_ = F4412 | new_F4429_;
  assign new_F4464_ = F4412 | F4413;
  assign new_F4465_ = new_F4429_ & new_F4466_;
  assign new_F4466_ = ~F4411 | ~new_F4436_;
  assign new_F4467_ = new_F4444_ & new_F4464_;
  assign new_F4468_ = ~new_F4444_ & ~new_F4464_;
  assign new_F4469_ = new_F4473_ | new_F4474_;
  assign new_F4470_ = ~F4415 & new_F4429_;
  assign new_F4471_ = new_F4475_ | new_F4476_;
  assign new_F4472_ = F4415 & new_F4429_;
  assign new_F4473_ = ~F4415 & ~new_F4429_;
  assign new_F4474_ = F4415 & ~new_F4429_;
  assign new_F4475_ = F4415 & ~new_F4429_;
  assign new_F4476_ = ~F4415 & new_F4429_;
  assign new_F4483_ = new_F4490_ & new_F4489_;
  assign new_F4484_ = new_F4492_ | new_F4491_;
  assign new_F4485_ = new_F4494_ | new_F4493_;
  assign new_F4486_ = new_F4496_ & new_F4495_;
  assign new_F4487_ = new_F4496_ & new_F4497_;
  assign new_F4488_ = new_F4489_ | new_F4498_;
  assign new_F4489_ = F4478 | new_F4501_;
  assign new_F4490_ = new_F4500_ | new_F4499_;
  assign new_F4491_ = new_F4505_ & new_F4504_;
  assign new_F4492_ = new_F4503_ & new_F4502_;
  assign new_F4493_ = new_F4508_ | new_F4507_;
  assign new_F4494_ = new_F4503_ & new_F4506_;
  assign new_F4495_ = F4478 | new_F4511_;
  assign new_F4496_ = new_F4510_ | new_F4509_;
  assign new_F4497_ = new_F4513_ | new_F4512_;
  assign new_F4498_ = ~new_F4489_ & new_F4515_;
  assign new_F4499_ = ~new_F4491_ & new_F4503_;
  assign new_F4500_ = new_F4491_ & ~new_F4503_;
  assign new_F4501_ = F4477 & ~F4478;
  assign new_F4502_ = ~new_F4524_ | ~new_F4525_;
  assign new_F4503_ = new_F4517_ | new_F4519_;
  assign new_F4504_ = new_F4527_ | new_F4526_;
  assign new_F4505_ = new_F4521_ | new_F4520_;
  assign new_F4506_ = ~new_F4529_ | ~new_F4528_;
  assign new_F4507_ = ~new_F4530_ & new_F4531_;
  assign new_F4508_ = new_F4530_ & ~new_F4531_;
  assign new_F4509_ = ~F4477 & F4478;
  assign new_F4510_ = F4477 & ~F4478;
  assign new_F4511_ = ~new_F4493_ | new_F4503_;
  assign new_F4512_ = new_F4493_ & new_F4503_;
  assign new_F4513_ = ~new_F4493_ & ~new_F4503_;
  assign new_F4514_ = new_F4535_ | new_F4534_;
  assign new_F4515_ = F4481 | new_F4514_;
  assign new_F4516_ = new_F4539_ | new_F4538_;
  assign new_F4517_ = ~F4481 & new_F4516_;
  assign new_F4518_ = new_F4537_ | new_F4536_;
  assign new_F4519_ = F4481 & new_F4518_;
  assign new_F4520_ = F4479 & ~new_F4489_;
  assign new_F4521_ = ~F4479 & new_F4489_;
  assign new_F4522_ = ~F4478 | ~new_F4503_;
  assign new_F4523_ = new_F4489_ & new_F4522_;
  assign new_F4524_ = ~new_F4489_ & ~new_F4523_;
  assign new_F4525_ = new_F4489_ | new_F4522_;
  assign new_F4526_ = ~F4479 & F4480;
  assign new_F4527_ = F4479 & ~F4480;
  assign new_F4528_ = new_F4496_ | new_F4533_;
  assign new_F4529_ = ~new_F4496_ & ~new_F4532_;
  assign new_F4530_ = F4479 | new_F4496_;
  assign new_F4531_ = F4479 | F4480;
  assign new_F4532_ = new_F4496_ & new_F4533_;
  assign new_F4533_ = ~F4478 | ~new_F4503_;
  assign new_F4534_ = new_F4511_ & new_F4531_;
  assign new_F4535_ = ~new_F4511_ & ~new_F4531_;
  assign new_F4536_ = new_F4540_ | new_F4541_;
  assign new_F4537_ = ~F4482 & new_F4496_;
  assign new_F4538_ = new_F4542_ | new_F4543_;
  assign new_F4539_ = F4482 & new_F4496_;
  assign new_F4540_ = ~F4482 & ~new_F4496_;
  assign new_F4541_ = F4482 & ~new_F4496_;
  assign new_F4542_ = F4482 & ~new_F4496_;
  assign new_F4543_ = ~F4482 & new_F4496_;
  assign new_F4550_ = new_F4557_ & new_F4556_;
  assign new_F4551_ = new_F4559_ | new_F4558_;
  assign new_F4552_ = new_F4561_ | new_F4560_;
  assign new_F4553_ = new_F4563_ & new_F4562_;
  assign new_F4554_ = new_F4563_ & new_F4564_;
  assign new_F4555_ = new_F4556_ | new_F4565_;
  assign new_F4556_ = F4545 | new_F4568_;
  assign new_F4557_ = new_F4567_ | new_F4566_;
  assign new_F4558_ = new_F4572_ & new_F4571_;
  assign new_F4559_ = new_F4570_ & new_F4569_;
  assign new_F4560_ = new_F4575_ | new_F4574_;
  assign new_F4561_ = new_F4570_ & new_F4573_;
  assign new_F4562_ = F4545 | new_F4578_;
  assign new_F4563_ = new_F4577_ | new_F4576_;
  assign new_F4564_ = new_F4580_ | new_F4579_;
  assign new_F4565_ = ~new_F4556_ & new_F4582_;
  assign new_F4566_ = ~new_F4558_ & new_F4570_;
  assign new_F4567_ = new_F4558_ & ~new_F4570_;
  assign new_F4568_ = F4544 & ~F4545;
  assign new_F4569_ = ~new_F4591_ | ~new_F4592_;
  assign new_F4570_ = new_F4584_ | new_F4586_;
  assign new_F4571_ = new_F4594_ | new_F4593_;
  assign new_F4572_ = new_F4588_ | new_F4587_;
  assign new_F4573_ = ~new_F4596_ | ~new_F4595_;
  assign new_F4574_ = ~new_F4597_ & new_F4598_;
  assign new_F4575_ = new_F4597_ & ~new_F4598_;
  assign new_F4576_ = ~F4544 & F4545;
  assign new_F4577_ = F4544 & ~F4545;
  assign new_F4578_ = ~new_F4560_ | new_F4570_;
  assign new_F4579_ = new_F4560_ & new_F4570_;
  assign new_F4580_ = ~new_F4560_ & ~new_F4570_;
  assign new_F4581_ = new_F4602_ | new_F4601_;
  assign new_F4582_ = F4548 | new_F4581_;
  assign new_F4583_ = new_F4606_ | new_F4605_;
  assign new_F4584_ = ~F4548 & new_F4583_;
  assign new_F4585_ = new_F4604_ | new_F4603_;
  assign new_F4586_ = F4548 & new_F4585_;
  assign new_F4587_ = F4546 & ~new_F4556_;
  assign new_F4588_ = ~F4546 & new_F4556_;
  assign new_F4589_ = ~F4545 | ~new_F4570_;
  assign new_F4590_ = new_F4556_ & new_F4589_;
  assign new_F4591_ = ~new_F4556_ & ~new_F4590_;
  assign new_F4592_ = new_F4556_ | new_F4589_;
  assign new_F4593_ = ~F4546 & F4547;
  assign new_F4594_ = F4546 & ~F4547;
  assign new_F4595_ = new_F4563_ | new_F4600_;
  assign new_F4596_ = ~new_F4563_ & ~new_F4599_;
  assign new_F4597_ = F4546 | new_F4563_;
  assign new_F4598_ = F4546 | F4547;
  assign new_F4599_ = new_F4563_ & new_F4600_;
  assign new_F4600_ = ~F4545 | ~new_F4570_;
  assign new_F4601_ = new_F4578_ & new_F4598_;
  assign new_F4602_ = ~new_F4578_ & ~new_F4598_;
  assign new_F4603_ = new_F4607_ | new_F4608_;
  assign new_F4604_ = ~F4549 & new_F4563_;
  assign new_F4605_ = new_F4609_ | new_F4610_;
  assign new_F4606_ = F4549 & new_F4563_;
  assign new_F4607_ = ~F4549 & ~new_F4563_;
  assign new_F4608_ = F4549 & ~new_F4563_;
  assign new_F4609_ = F4549 & ~new_F4563_;
  assign new_F4610_ = ~F4549 & new_F4563_;
  assign new_F4617_ = new_F4624_ & new_F4623_;
  assign new_F4618_ = new_F4626_ | new_F4625_;
  assign new_F4619_ = new_F4628_ | new_F4627_;
  assign new_F4620_ = new_F4630_ & new_F4629_;
  assign new_F4621_ = new_F4630_ & new_F4631_;
  assign new_F4622_ = new_F4623_ | new_F4632_;
  assign new_F4623_ = F4612 | new_F4635_;
  assign new_F4624_ = new_F4634_ | new_F4633_;
  assign new_F4625_ = new_F4639_ & new_F4638_;
  assign new_F4626_ = new_F4637_ & new_F4636_;
  assign new_F4627_ = new_F4642_ | new_F4641_;
  assign new_F4628_ = new_F4637_ & new_F4640_;
  assign new_F4629_ = F4612 | new_F4645_;
  assign new_F4630_ = new_F4644_ | new_F4643_;
  assign new_F4631_ = new_F4647_ | new_F4646_;
  assign new_F4632_ = ~new_F4623_ & new_F4649_;
  assign new_F4633_ = ~new_F4625_ & new_F4637_;
  assign new_F4634_ = new_F4625_ & ~new_F4637_;
  assign new_F4635_ = F4611 & ~F4612;
  assign new_F4636_ = ~new_F4658_ | ~new_F4659_;
  assign new_F4637_ = new_F4651_ | new_F4653_;
  assign new_F4638_ = new_F4661_ | new_F4660_;
  assign new_F4639_ = new_F4655_ | new_F4654_;
  assign new_F4640_ = ~new_F4663_ | ~new_F4662_;
  assign new_F4641_ = ~new_F4664_ & new_F4665_;
  assign new_F4642_ = new_F4664_ & ~new_F4665_;
  assign new_F4643_ = ~F4611 & F4612;
  assign new_F4644_ = F4611 & ~F4612;
  assign new_F4645_ = ~new_F4627_ | new_F4637_;
  assign new_F4646_ = new_F4627_ & new_F4637_;
  assign new_F4647_ = ~new_F4627_ & ~new_F4637_;
  assign new_F4648_ = new_F4669_ | new_F4668_;
  assign new_F4649_ = F4615 | new_F4648_;
  assign new_F4650_ = new_F4673_ | new_F4672_;
  assign new_F4651_ = ~F4615 & new_F4650_;
  assign new_F4652_ = new_F4671_ | new_F4670_;
  assign new_F4653_ = F4615 & new_F4652_;
  assign new_F4654_ = F4613 & ~new_F4623_;
  assign new_F4655_ = ~F4613 & new_F4623_;
  assign new_F4656_ = ~F4612 | ~new_F4637_;
  assign new_F4657_ = new_F4623_ & new_F4656_;
  assign new_F4658_ = ~new_F4623_ & ~new_F4657_;
  assign new_F4659_ = new_F4623_ | new_F4656_;
  assign new_F4660_ = ~F4613 & F4614;
  assign new_F4661_ = F4613 & ~F4614;
  assign new_F4662_ = new_F4630_ | new_F4667_;
  assign new_F4663_ = ~new_F4630_ & ~new_F4666_;
  assign new_F4664_ = F4613 | new_F4630_;
  assign new_F4665_ = F4613 | F4614;
  assign new_F4666_ = new_F4630_ & new_F4667_;
  assign new_F4667_ = ~F4612 | ~new_F4637_;
  assign new_F4668_ = new_F4645_ & new_F4665_;
  assign new_F4669_ = ~new_F4645_ & ~new_F4665_;
  assign new_F4670_ = new_F4674_ | new_F4675_;
  assign new_F4671_ = ~F4616 & new_F4630_;
  assign new_F4672_ = new_F4676_ | new_F4677_;
  assign new_F4673_ = F4616 & new_F4630_;
  assign new_F4674_ = ~F4616 & ~new_F4630_;
  assign new_F4675_ = F4616 & ~new_F4630_;
  assign new_F4676_ = F4616 & ~new_F4630_;
  assign new_F4677_ = ~F4616 & new_F4630_;
  assign new_F4684_ = new_F4691_ & new_F4690_;
  assign new_F4685_ = new_F4693_ | new_F4692_;
  assign new_F4686_ = new_F4695_ | new_F4694_;
  assign new_F4687_ = new_F4697_ & new_F4696_;
  assign new_F4688_ = new_F4697_ & new_F4698_;
  assign new_F4689_ = new_F4690_ | new_F4699_;
  assign new_F4690_ = F4679 | new_F4702_;
  assign new_F4691_ = new_F4701_ | new_F4700_;
  assign new_F4692_ = new_F4706_ & new_F4705_;
  assign new_F4693_ = new_F4704_ & new_F4703_;
  assign new_F4694_ = new_F4709_ | new_F4708_;
  assign new_F4695_ = new_F4704_ & new_F4707_;
  assign new_F4696_ = F4679 | new_F4712_;
  assign new_F4697_ = new_F4711_ | new_F4710_;
  assign new_F4698_ = new_F4714_ | new_F4713_;
  assign new_F4699_ = ~new_F4690_ & new_F4716_;
  assign new_F4700_ = ~new_F4692_ & new_F4704_;
  assign new_F4701_ = new_F4692_ & ~new_F4704_;
  assign new_F4702_ = F4678 & ~F4679;
  assign new_F4703_ = ~new_F4725_ | ~new_F4726_;
  assign new_F4704_ = new_F4718_ | new_F4720_;
  assign new_F4705_ = new_F4728_ | new_F4727_;
  assign new_F4706_ = new_F4722_ | new_F4721_;
  assign new_F4707_ = ~new_F4730_ | ~new_F4729_;
  assign new_F4708_ = ~new_F4731_ & new_F4732_;
  assign new_F4709_ = new_F4731_ & ~new_F4732_;
  assign new_F4710_ = ~F4678 & F4679;
  assign new_F4711_ = F4678 & ~F4679;
  assign new_F4712_ = ~new_F4694_ | new_F4704_;
  assign new_F4713_ = new_F4694_ & new_F4704_;
  assign new_F4714_ = ~new_F4694_ & ~new_F4704_;
  assign new_F4715_ = new_F4736_ | new_F4735_;
  assign new_F4716_ = F4682 | new_F4715_;
  assign new_F4717_ = new_F4740_ | new_F4739_;
  assign new_F4718_ = ~F4682 & new_F4717_;
  assign new_F4719_ = new_F4738_ | new_F4737_;
  assign new_F4720_ = F4682 & new_F4719_;
  assign new_F4721_ = F4680 & ~new_F4690_;
  assign new_F4722_ = ~F4680 & new_F4690_;
  assign new_F4723_ = ~F4679 | ~new_F4704_;
  assign new_F4724_ = new_F4690_ & new_F4723_;
  assign new_F4725_ = ~new_F4690_ & ~new_F4724_;
  assign new_F4726_ = new_F4690_ | new_F4723_;
  assign new_F4727_ = ~F4680 & F4681;
  assign new_F4728_ = F4680 & ~F4681;
  assign new_F4729_ = new_F4697_ | new_F4734_;
  assign new_F4730_ = ~new_F4697_ & ~new_F4733_;
  assign new_F4731_ = F4680 | new_F4697_;
  assign new_F4732_ = F4680 | F4681;
  assign new_F4733_ = new_F4697_ & new_F4734_;
  assign new_F4734_ = ~F4679 | ~new_F4704_;
  assign new_F4735_ = new_F4712_ & new_F4732_;
  assign new_F4736_ = ~new_F4712_ & ~new_F4732_;
  assign new_F4737_ = new_F4741_ | new_F4742_;
  assign new_F4738_ = ~F4683 & new_F4697_;
  assign new_F4739_ = new_F4743_ | new_F4744_;
  assign new_F4740_ = F4683 & new_F4697_;
  assign new_F4741_ = ~F4683 & ~new_F4697_;
  assign new_F4742_ = F4683 & ~new_F4697_;
  assign new_F4743_ = F4683 & ~new_F4697_;
  assign new_F4744_ = ~F4683 & new_F4697_;
  assign new_F4751_ = new_F4758_ & new_F4757_;
  assign new_F4752_ = new_F4760_ | new_F4759_;
  assign new_F4753_ = new_F4762_ | new_F4761_;
  assign new_F4754_ = new_F4764_ & new_F4763_;
  assign new_F4755_ = new_F4764_ & new_F4765_;
  assign new_F4756_ = new_F4757_ | new_F4766_;
  assign new_F4757_ = F4746 | new_F4769_;
  assign new_F4758_ = new_F4768_ | new_F4767_;
  assign new_F4759_ = new_F4773_ & new_F4772_;
  assign new_F4760_ = new_F4771_ & new_F4770_;
  assign new_F4761_ = new_F4776_ | new_F4775_;
  assign new_F4762_ = new_F4771_ & new_F4774_;
  assign new_F4763_ = F4746 | new_F4779_;
  assign new_F4764_ = new_F4778_ | new_F4777_;
  assign new_F4765_ = new_F4781_ | new_F4780_;
  assign new_F4766_ = ~new_F4757_ & new_F4783_;
  assign new_F4767_ = ~new_F4759_ & new_F4771_;
  assign new_F4768_ = new_F4759_ & ~new_F4771_;
  assign new_F4769_ = F4745 & ~F4746;
  assign new_F4770_ = ~new_F4792_ | ~new_F4793_;
  assign new_F4771_ = new_F4785_ | new_F4787_;
  assign new_F4772_ = new_F4795_ | new_F4794_;
  assign new_F4773_ = new_F4789_ | new_F4788_;
  assign new_F4774_ = ~new_F4797_ | ~new_F4796_;
  assign new_F4775_ = ~new_F4798_ & new_F4799_;
  assign new_F4776_ = new_F4798_ & ~new_F4799_;
  assign new_F4777_ = ~F4745 & F4746;
  assign new_F4778_ = F4745 & ~F4746;
  assign new_F4779_ = ~new_F4761_ | new_F4771_;
  assign new_F4780_ = new_F4761_ & new_F4771_;
  assign new_F4781_ = ~new_F4761_ & ~new_F4771_;
  assign new_F4782_ = new_F4803_ | new_F4802_;
  assign new_F4783_ = F4749 | new_F4782_;
  assign new_F4784_ = new_F4807_ | new_F4806_;
  assign new_F4785_ = ~F4749 & new_F4784_;
  assign new_F4786_ = new_F4805_ | new_F4804_;
  assign new_F4787_ = F4749 & new_F4786_;
  assign new_F4788_ = F4747 & ~new_F4757_;
  assign new_F4789_ = ~F4747 & new_F4757_;
  assign new_F4790_ = ~F4746 | ~new_F4771_;
  assign new_F4791_ = new_F4757_ & new_F4790_;
  assign new_F4792_ = ~new_F4757_ & ~new_F4791_;
  assign new_F4793_ = new_F4757_ | new_F4790_;
  assign new_F4794_ = ~F4747 & F4748;
  assign new_F4795_ = F4747 & ~F4748;
  assign new_F4796_ = new_F4764_ | new_F4801_;
  assign new_F4797_ = ~new_F4764_ & ~new_F4800_;
  assign new_F4798_ = F4747 | new_F4764_;
  assign new_F4799_ = F4747 | F4748;
  assign new_F4800_ = new_F4764_ & new_F4801_;
  assign new_F4801_ = ~F4746 | ~new_F4771_;
  assign new_F4802_ = new_F4779_ & new_F4799_;
  assign new_F4803_ = ~new_F4779_ & ~new_F4799_;
  assign new_F4804_ = new_F4808_ | new_F4809_;
  assign new_F4805_ = ~F4750 & new_F4764_;
  assign new_F4806_ = new_F4810_ | new_F4811_;
  assign new_F4807_ = F4750 & new_F4764_;
  assign new_F4808_ = ~F4750 & ~new_F4764_;
  assign new_F4809_ = F4750 & ~new_F4764_;
  assign new_F4810_ = F4750 & ~new_F4764_;
  assign new_F4811_ = ~F4750 & new_F4764_;
  assign new_F4818_ = new_F4825_ & new_F4824_;
  assign new_F4819_ = new_F4827_ | new_F4826_;
  assign new_F4820_ = new_F4829_ | new_F4828_;
  assign new_F4821_ = new_F4831_ & new_F4830_;
  assign new_F4822_ = new_F4831_ & new_F4832_;
  assign new_F4823_ = new_F4824_ | new_F4833_;
  assign new_F4824_ = F4813 | new_F4836_;
  assign new_F4825_ = new_F4835_ | new_F4834_;
  assign new_F4826_ = new_F4840_ & new_F4839_;
  assign new_F4827_ = new_F4838_ & new_F4837_;
  assign new_F4828_ = new_F4843_ | new_F4842_;
  assign new_F4829_ = new_F4838_ & new_F4841_;
  assign new_F4830_ = F4813 | new_F4846_;
  assign new_F4831_ = new_F4845_ | new_F4844_;
  assign new_F4832_ = new_F4848_ | new_F4847_;
  assign new_F4833_ = ~new_F4824_ & new_F4850_;
  assign new_F4834_ = ~new_F4826_ & new_F4838_;
  assign new_F4835_ = new_F4826_ & ~new_F4838_;
  assign new_F4836_ = F4812 & ~F4813;
  assign new_F4837_ = ~new_F4859_ | ~new_F4860_;
  assign new_F4838_ = new_F4852_ | new_F4854_;
  assign new_F4839_ = new_F4862_ | new_F4861_;
  assign new_F4840_ = new_F4856_ | new_F4855_;
  assign new_F4841_ = ~new_F4864_ | ~new_F4863_;
  assign new_F4842_ = ~new_F4865_ & new_F4866_;
  assign new_F4843_ = new_F4865_ & ~new_F4866_;
  assign new_F4844_ = ~F4812 & F4813;
  assign new_F4845_ = F4812 & ~F4813;
  assign new_F4846_ = ~new_F4828_ | new_F4838_;
  assign new_F4847_ = new_F4828_ & new_F4838_;
  assign new_F4848_ = ~new_F4828_ & ~new_F4838_;
  assign new_F4849_ = new_F4870_ | new_F4869_;
  assign new_F4850_ = F4816 | new_F4849_;
  assign new_F4851_ = new_F4874_ | new_F4873_;
  assign new_F4852_ = ~F4816 & new_F4851_;
  assign new_F4853_ = new_F4872_ | new_F4871_;
  assign new_F4854_ = F4816 & new_F4853_;
  assign new_F4855_ = F4814 & ~new_F4824_;
  assign new_F4856_ = ~F4814 & new_F4824_;
  assign new_F4857_ = ~F4813 | ~new_F4838_;
  assign new_F4858_ = new_F4824_ & new_F4857_;
  assign new_F4859_ = ~new_F4824_ & ~new_F4858_;
  assign new_F4860_ = new_F4824_ | new_F4857_;
  assign new_F4861_ = ~F4814 & F4815;
  assign new_F4862_ = F4814 & ~F4815;
  assign new_F4863_ = new_F4831_ | new_F4868_;
  assign new_F4864_ = ~new_F4831_ & ~new_F4867_;
  assign new_F4865_ = F4814 | new_F4831_;
  assign new_F4866_ = F4814 | F4815;
  assign new_F4867_ = new_F4831_ & new_F4868_;
  assign new_F4868_ = ~F4813 | ~new_F4838_;
  assign new_F4869_ = new_F4846_ & new_F4866_;
  assign new_F4870_ = ~new_F4846_ & ~new_F4866_;
  assign new_F4871_ = new_F4875_ | new_F4876_;
  assign new_F4872_ = ~F4817 & new_F4831_;
  assign new_F4873_ = new_F4877_ | new_F4878_;
  assign new_F4874_ = F4817 & new_F4831_;
  assign new_F4875_ = ~F4817 & ~new_F4831_;
  assign new_F4876_ = F4817 & ~new_F4831_;
  assign new_F4877_ = F4817 & ~new_F4831_;
  assign new_F4878_ = ~F4817 & new_F4831_;
  assign new_F4885_ = new_F4892_ & new_F4891_;
  assign new_F4886_ = new_F4894_ | new_F4893_;
  assign new_F4887_ = new_F4896_ | new_F4895_;
  assign new_F4888_ = new_F4898_ & new_F4897_;
  assign new_F4889_ = new_F4898_ & new_F4899_;
  assign new_F4890_ = new_F4891_ | new_F4900_;
  assign new_F4891_ = F4880 | new_F4903_;
  assign new_F4892_ = new_F4902_ | new_F4901_;
  assign new_F4893_ = new_F4907_ & new_F4906_;
  assign new_F4894_ = new_F4905_ & new_F4904_;
  assign new_F4895_ = new_F4910_ | new_F4909_;
  assign new_F4896_ = new_F4905_ & new_F4908_;
  assign new_F4897_ = F4880 | new_F4913_;
  assign new_F4898_ = new_F4912_ | new_F4911_;
  assign new_F4899_ = new_F4915_ | new_F4914_;
  assign new_F4900_ = ~new_F4891_ & new_F4917_;
  assign new_F4901_ = ~new_F4893_ & new_F4905_;
  assign new_F4902_ = new_F4893_ & ~new_F4905_;
  assign new_F4903_ = F4879 & ~F4880;
  assign new_F4904_ = ~new_F4926_ | ~new_F4927_;
  assign new_F4905_ = new_F4919_ | new_F4921_;
  assign new_F4906_ = new_F4929_ | new_F4928_;
  assign new_F4907_ = new_F4923_ | new_F4922_;
  assign new_F4908_ = ~new_F4931_ | ~new_F4930_;
  assign new_F4909_ = ~new_F4932_ & new_F4933_;
  assign new_F4910_ = new_F4932_ & ~new_F4933_;
  assign new_F4911_ = ~F4879 & F4880;
  assign new_F4912_ = F4879 & ~F4880;
  assign new_F4913_ = ~new_F4895_ | new_F4905_;
  assign new_F4914_ = new_F4895_ & new_F4905_;
  assign new_F4915_ = ~new_F4895_ & ~new_F4905_;
  assign new_F4916_ = new_F4937_ | new_F4936_;
  assign new_F4917_ = F4883 | new_F4916_;
  assign new_F4918_ = new_F4941_ | new_F4940_;
  assign new_F4919_ = ~F4883 & new_F4918_;
  assign new_F4920_ = new_F4939_ | new_F4938_;
  assign new_F4921_ = F4883 & new_F4920_;
  assign new_F4922_ = F4881 & ~new_F4891_;
  assign new_F4923_ = ~F4881 & new_F4891_;
  assign new_F4924_ = ~F4880 | ~new_F4905_;
  assign new_F4925_ = new_F4891_ & new_F4924_;
  assign new_F4926_ = ~new_F4891_ & ~new_F4925_;
  assign new_F4927_ = new_F4891_ | new_F4924_;
  assign new_F4928_ = ~F4881 & F4882;
  assign new_F4929_ = F4881 & ~F4882;
  assign new_F4930_ = new_F4898_ | new_F4935_;
  assign new_F4931_ = ~new_F4898_ & ~new_F4934_;
  assign new_F4932_ = F4881 | new_F4898_;
  assign new_F4933_ = F4881 | F4882;
  assign new_F4934_ = new_F4898_ & new_F4935_;
  assign new_F4935_ = ~F4880 | ~new_F4905_;
  assign new_F4936_ = new_F4913_ & new_F4933_;
  assign new_F4937_ = ~new_F4913_ & ~new_F4933_;
  assign new_F4938_ = new_F4942_ | new_F4943_;
  assign new_F4939_ = ~F4884 & new_F4898_;
  assign new_F4940_ = new_F4944_ | new_F4945_;
  assign new_F4941_ = F4884 & new_F4898_;
  assign new_F4942_ = ~F4884 & ~new_F4898_;
  assign new_F4943_ = F4884 & ~new_F4898_;
  assign new_F4944_ = F4884 & ~new_F4898_;
  assign new_F4945_ = ~F4884 & new_F4898_;
  assign new_F4952_ = new_F4959_ & new_F4958_;
  assign new_F4953_ = new_F4961_ | new_F4960_;
  assign new_F4954_ = new_F4963_ | new_F4962_;
  assign new_F4955_ = new_F4965_ & new_F4964_;
  assign new_F4956_ = new_F4965_ & new_F4966_;
  assign new_F4957_ = new_F4958_ | new_F4967_;
  assign new_F4958_ = F4947 | new_F4970_;
  assign new_F4959_ = new_F4969_ | new_F4968_;
  assign new_F4960_ = new_F4974_ & new_F4973_;
  assign new_F4961_ = new_F4972_ & new_F4971_;
  assign new_F4962_ = new_F4977_ | new_F4976_;
  assign new_F4963_ = new_F4972_ & new_F4975_;
  assign new_F4964_ = F4947 | new_F4980_;
  assign new_F4965_ = new_F4979_ | new_F4978_;
  assign new_F4966_ = new_F4982_ | new_F4981_;
  assign new_F4967_ = ~new_F4958_ & new_F4984_;
  assign new_F4968_ = ~new_F4960_ & new_F4972_;
  assign new_F4969_ = new_F4960_ & ~new_F4972_;
  assign new_F4970_ = F4946 & ~F4947;
  assign new_F4971_ = ~new_F4993_ | ~new_F4994_;
  assign new_F4972_ = new_F4986_ | new_F4988_;
  assign new_F4973_ = new_F4996_ | new_F4995_;
  assign new_F4974_ = new_F4990_ | new_F4989_;
  assign new_F4975_ = ~new_F4998_ | ~new_F4997_;
  assign new_F4976_ = ~new_F4999_ & new_F5000_;
  assign new_F4977_ = new_F4999_ & ~new_F5000_;
  assign new_F4978_ = ~F4946 & F4947;
  assign new_F4979_ = F4946 & ~F4947;
  assign new_F4980_ = ~new_F4962_ | new_F4972_;
  assign new_F4981_ = new_F4962_ & new_F4972_;
  assign new_F4982_ = ~new_F4962_ & ~new_F4972_;
  assign new_F4983_ = new_F5004_ | new_F5003_;
  assign new_F4984_ = F4950 | new_F4983_;
  assign new_F4985_ = new_F5008_ | new_F5007_;
  assign new_F4986_ = ~F4950 & new_F4985_;
  assign new_F4987_ = new_F5006_ | new_F5005_;
  assign new_F4988_ = F4950 & new_F4987_;
  assign new_F4989_ = F4948 & ~new_F4958_;
  assign new_F4990_ = ~F4948 & new_F4958_;
  assign new_F4991_ = ~F4947 | ~new_F4972_;
  assign new_F4992_ = new_F4958_ & new_F4991_;
  assign new_F4993_ = ~new_F4958_ & ~new_F4992_;
  assign new_F4994_ = new_F4958_ | new_F4991_;
  assign new_F4995_ = ~F4948 & F4949;
  assign new_F4996_ = F4948 & ~F4949;
  assign new_F4997_ = new_F4965_ | new_F5002_;
  assign new_F4998_ = ~new_F4965_ & ~new_F5001_;
  assign new_F4999_ = F4948 | new_F4965_;
  assign new_F5000_ = F4948 | F4949;
  assign new_F5001_ = new_F4965_ & new_F5002_;
  assign new_F5002_ = ~F4947 | ~new_F4972_;
  assign new_F5003_ = new_F4980_ & new_F5000_;
  assign new_F5004_ = ~new_F4980_ & ~new_F5000_;
  assign new_F5005_ = new_F5009_ | new_F5010_;
  assign new_F5006_ = ~F4951 & new_F4965_;
  assign new_F5007_ = new_F5011_ | new_F5012_;
  assign new_F5008_ = F4951 & new_F4965_;
  assign new_F5009_ = ~F4951 & ~new_F4965_;
  assign new_F5010_ = F4951 & ~new_F4965_;
  assign new_F5011_ = F4951 & ~new_F4965_;
  assign new_F5012_ = ~F4951 & new_F4965_;
  assign new_F5019_ = new_F5026_ & new_F5025_;
  assign new_F5020_ = new_F5028_ | new_F5027_;
  assign new_F5021_ = new_F5030_ | new_F5029_;
  assign new_F5022_ = new_F5032_ & new_F5031_;
  assign new_F5023_ = new_F5032_ & new_F5033_;
  assign new_F5024_ = new_F5025_ | new_F5034_;
  assign new_F5025_ = F5014 | new_F5037_;
  assign new_F5026_ = new_F5036_ | new_F5035_;
  assign new_F5027_ = new_F5041_ & new_F5040_;
  assign new_F5028_ = new_F5039_ & new_F5038_;
  assign new_F5029_ = new_F5044_ | new_F5043_;
  assign new_F5030_ = new_F5039_ & new_F5042_;
  assign new_F5031_ = F5014 | new_F5047_;
  assign new_F5032_ = new_F5046_ | new_F5045_;
  assign new_F5033_ = new_F5049_ | new_F5048_;
  assign new_F5034_ = ~new_F5025_ & new_F5051_;
  assign new_F5035_ = ~new_F5027_ & new_F5039_;
  assign new_F5036_ = new_F5027_ & ~new_F5039_;
  assign new_F5037_ = F5013 & ~F5014;
  assign new_F5038_ = ~new_F5060_ | ~new_F5061_;
  assign new_F5039_ = new_F5053_ | new_F5055_;
  assign new_F5040_ = new_F5063_ | new_F5062_;
  assign new_F5041_ = new_F5057_ | new_F5056_;
  assign new_F5042_ = ~new_F5065_ | ~new_F5064_;
  assign new_F5043_ = ~new_F5066_ & new_F5067_;
  assign new_F5044_ = new_F5066_ & ~new_F5067_;
  assign new_F5045_ = ~F5013 & F5014;
  assign new_F5046_ = F5013 & ~F5014;
  assign new_F5047_ = ~new_F5029_ | new_F5039_;
  assign new_F5048_ = new_F5029_ & new_F5039_;
  assign new_F5049_ = ~new_F5029_ & ~new_F5039_;
  assign new_F5050_ = new_F5071_ | new_F5070_;
  assign new_F5051_ = F5017 | new_F5050_;
  assign new_F5052_ = new_F5075_ | new_F5074_;
  assign new_F5053_ = ~F5017 & new_F5052_;
  assign new_F5054_ = new_F5073_ | new_F5072_;
  assign new_F5055_ = F5017 & new_F5054_;
  assign new_F5056_ = F5015 & ~new_F5025_;
  assign new_F5057_ = ~F5015 & new_F5025_;
  assign new_F5058_ = ~F5014 | ~new_F5039_;
  assign new_F5059_ = new_F5025_ & new_F5058_;
  assign new_F5060_ = ~new_F5025_ & ~new_F5059_;
  assign new_F5061_ = new_F5025_ | new_F5058_;
  assign new_F5062_ = ~F5015 & F5016;
  assign new_F5063_ = F5015 & ~F5016;
  assign new_F5064_ = new_F5032_ | new_F5069_;
  assign new_F5065_ = ~new_F5032_ & ~new_F5068_;
  assign new_F5066_ = F5015 | new_F5032_;
  assign new_F5067_ = F5015 | F5016;
  assign new_F5068_ = new_F5032_ & new_F5069_;
  assign new_F5069_ = ~F5014 | ~new_F5039_;
  assign new_F5070_ = new_F5047_ & new_F5067_;
  assign new_F5071_ = ~new_F5047_ & ~new_F5067_;
  assign new_F5072_ = new_F5076_ | new_F5077_;
  assign new_F5073_ = ~F5018 & new_F5032_;
  assign new_F5074_ = new_F5078_ | new_F5079_;
  assign new_F5075_ = F5018 & new_F5032_;
  assign new_F5076_ = ~F5018 & ~new_F5032_;
  assign new_F5077_ = F5018 & ~new_F5032_;
  assign new_F5078_ = F5018 & ~new_F5032_;
  assign new_F5079_ = ~F5018 & new_F5032_;
  assign new_F5086_ = new_F5093_ & new_F5092_;
  assign new_F5087_ = new_F5095_ | new_F5094_;
  assign new_F5088_ = new_F5097_ | new_F5096_;
  assign new_F5089_ = new_F5099_ & new_F5098_;
  assign new_F5090_ = new_F5099_ & new_F5100_;
  assign new_F5091_ = new_F5092_ | new_F5101_;
  assign new_F5092_ = F5081 | new_F5104_;
  assign new_F5093_ = new_F5103_ | new_F5102_;
  assign new_F5094_ = new_F5108_ & new_F5107_;
  assign new_F5095_ = new_F5106_ & new_F5105_;
  assign new_F5096_ = new_F5111_ | new_F5110_;
  assign new_F5097_ = new_F5106_ & new_F5109_;
  assign new_F5098_ = F5081 | new_F5114_;
  assign new_F5099_ = new_F5113_ | new_F5112_;
  assign new_F5100_ = new_F5116_ | new_F5115_;
  assign new_F5101_ = ~new_F5092_ & new_F5118_;
  assign new_F5102_ = ~new_F5094_ & new_F5106_;
  assign new_F5103_ = new_F5094_ & ~new_F5106_;
  assign new_F5104_ = F5080 & ~F5081;
  assign new_F5105_ = ~new_F5127_ | ~new_F5128_;
  assign new_F5106_ = new_F5120_ | new_F5122_;
  assign new_F5107_ = new_F5130_ | new_F5129_;
  assign new_F5108_ = new_F5124_ | new_F5123_;
  assign new_F5109_ = ~new_F5132_ | ~new_F5131_;
  assign new_F5110_ = ~new_F5133_ & new_F5134_;
  assign new_F5111_ = new_F5133_ & ~new_F5134_;
  assign new_F5112_ = ~F5080 & F5081;
  assign new_F5113_ = F5080 & ~F5081;
  assign new_F5114_ = ~new_F5096_ | new_F5106_;
  assign new_F5115_ = new_F5096_ & new_F5106_;
  assign new_F5116_ = ~new_F5096_ & ~new_F5106_;
  assign new_F5117_ = new_F5138_ | new_F5137_;
  assign new_F5118_ = F5084 | new_F5117_;
  assign new_F5119_ = new_F5142_ | new_F5141_;
  assign new_F5120_ = ~F5084 & new_F5119_;
  assign new_F5121_ = new_F5140_ | new_F5139_;
  assign new_F5122_ = F5084 & new_F5121_;
  assign new_F5123_ = F5082 & ~new_F5092_;
  assign new_F5124_ = ~F5082 & new_F5092_;
  assign new_F5125_ = ~F5081 | ~new_F5106_;
  assign new_F5126_ = new_F5092_ & new_F5125_;
  assign new_F5127_ = ~new_F5092_ & ~new_F5126_;
  assign new_F5128_ = new_F5092_ | new_F5125_;
  assign new_F5129_ = ~F5082 & F5083;
  assign new_F5130_ = F5082 & ~F5083;
  assign new_F5131_ = new_F5099_ | new_F5136_;
  assign new_F5132_ = ~new_F5099_ & ~new_F5135_;
  assign new_F5133_ = F5082 | new_F5099_;
  assign new_F5134_ = F5082 | F5083;
  assign new_F5135_ = new_F5099_ & new_F5136_;
  assign new_F5136_ = ~F5081 | ~new_F5106_;
  assign new_F5137_ = new_F5114_ & new_F5134_;
  assign new_F5138_ = ~new_F5114_ & ~new_F5134_;
  assign new_F5139_ = new_F5143_ | new_F5144_;
  assign new_F5140_ = ~F5085 & new_F5099_;
  assign new_F5141_ = new_F5145_ | new_F5146_;
  assign new_F5142_ = F5085 & new_F5099_;
  assign new_F5143_ = ~F5085 & ~new_F5099_;
  assign new_F5144_ = F5085 & ~new_F5099_;
  assign new_F5145_ = F5085 & ~new_F5099_;
  assign new_F5146_ = ~F5085 & new_F5099_;
  assign new_F5153_ = new_F5160_ & new_F5159_;
  assign new_F5154_ = new_F5162_ | new_F5161_;
  assign new_F5155_ = new_F5164_ | new_F5163_;
  assign new_F5156_ = new_F5166_ & new_F5165_;
  assign new_F5157_ = new_F5166_ & new_F5167_;
  assign new_F5158_ = new_F5159_ | new_F5168_;
  assign new_F5159_ = F5148 | new_F5171_;
  assign new_F5160_ = new_F5170_ | new_F5169_;
  assign new_F5161_ = new_F5175_ & new_F5174_;
  assign new_F5162_ = new_F5173_ & new_F5172_;
  assign new_F5163_ = new_F5178_ | new_F5177_;
  assign new_F5164_ = new_F5173_ & new_F5176_;
  assign new_F5165_ = F5148 | new_F5181_;
  assign new_F5166_ = new_F5180_ | new_F5179_;
  assign new_F5167_ = new_F5183_ | new_F5182_;
  assign new_F5168_ = ~new_F5159_ & new_F5185_;
  assign new_F5169_ = ~new_F5161_ & new_F5173_;
  assign new_F5170_ = new_F5161_ & ~new_F5173_;
  assign new_F5171_ = F5147 & ~F5148;
  assign new_F5172_ = ~new_F5194_ | ~new_F5195_;
  assign new_F5173_ = new_F5187_ | new_F5189_;
  assign new_F5174_ = new_F5197_ | new_F5196_;
  assign new_F5175_ = new_F5191_ | new_F5190_;
  assign new_F5176_ = ~new_F5199_ | ~new_F5198_;
  assign new_F5177_ = ~new_F5200_ & new_F5201_;
  assign new_F5178_ = new_F5200_ & ~new_F5201_;
  assign new_F5179_ = ~F5147 & F5148;
  assign new_F5180_ = F5147 & ~F5148;
  assign new_F5181_ = ~new_F5163_ | new_F5173_;
  assign new_F5182_ = new_F5163_ & new_F5173_;
  assign new_F5183_ = ~new_F5163_ & ~new_F5173_;
  assign new_F5184_ = new_F5205_ | new_F5204_;
  assign new_F5185_ = F5151 | new_F5184_;
  assign new_F5186_ = new_F5209_ | new_F5208_;
  assign new_F5187_ = ~F5151 & new_F5186_;
  assign new_F5188_ = new_F5207_ | new_F5206_;
  assign new_F5189_ = F5151 & new_F5188_;
  assign new_F5190_ = F5149 & ~new_F5159_;
  assign new_F5191_ = ~F5149 & new_F5159_;
  assign new_F5192_ = ~F5148 | ~new_F5173_;
  assign new_F5193_ = new_F5159_ & new_F5192_;
  assign new_F5194_ = ~new_F5159_ & ~new_F5193_;
  assign new_F5195_ = new_F5159_ | new_F5192_;
  assign new_F5196_ = ~F5149 & F5150;
  assign new_F5197_ = F5149 & ~F5150;
  assign new_F5198_ = new_F5166_ | new_F5203_;
  assign new_F5199_ = ~new_F5166_ & ~new_F5202_;
  assign new_F5200_ = F5149 | new_F5166_;
  assign new_F5201_ = F5149 | F5150;
  assign new_F5202_ = new_F5166_ & new_F5203_;
  assign new_F5203_ = ~F5148 | ~new_F5173_;
  assign new_F5204_ = new_F5181_ & new_F5201_;
  assign new_F5205_ = ~new_F5181_ & ~new_F5201_;
  assign new_F5206_ = new_F5210_ | new_F5211_;
  assign new_F5207_ = ~F5152 & new_F5166_;
  assign new_F5208_ = new_F5212_ | new_F5213_;
  assign new_F5209_ = F5152 & new_F5166_;
  assign new_F5210_ = ~F5152 & ~new_F5166_;
  assign new_F5211_ = F5152 & ~new_F5166_;
  assign new_F5212_ = F5152 & ~new_F5166_;
  assign new_F5213_ = ~F5152 & new_F5166_;
  assign new_F5220_ = new_F5227_ & new_F5226_;
  assign new_F5221_ = new_F5229_ | new_F5228_;
  assign new_F5222_ = new_F5231_ | new_F5230_;
  assign new_F5223_ = new_F5233_ & new_F5232_;
  assign new_F5224_ = new_F5233_ & new_F5234_;
  assign new_F5225_ = new_F5226_ | new_F5235_;
  assign new_F5226_ = F5215 | new_F5238_;
  assign new_F5227_ = new_F5237_ | new_F5236_;
  assign new_F5228_ = new_F5242_ & new_F5241_;
  assign new_F5229_ = new_F5240_ & new_F5239_;
  assign new_F5230_ = new_F5245_ | new_F5244_;
  assign new_F5231_ = new_F5240_ & new_F5243_;
  assign new_F5232_ = F5215 | new_F5248_;
  assign new_F5233_ = new_F5247_ | new_F5246_;
  assign new_F5234_ = new_F5250_ | new_F5249_;
  assign new_F5235_ = ~new_F5226_ & new_F5252_;
  assign new_F5236_ = ~new_F5228_ & new_F5240_;
  assign new_F5237_ = new_F5228_ & ~new_F5240_;
  assign new_F5238_ = F5214 & ~F5215;
  assign new_F5239_ = ~new_F5261_ | ~new_F5262_;
  assign new_F5240_ = new_F5254_ | new_F5256_;
  assign new_F5241_ = new_F5264_ | new_F5263_;
  assign new_F5242_ = new_F5258_ | new_F5257_;
  assign new_F5243_ = ~new_F5266_ | ~new_F5265_;
  assign new_F5244_ = ~new_F5267_ & new_F5268_;
  assign new_F5245_ = new_F5267_ & ~new_F5268_;
  assign new_F5246_ = ~F5214 & F5215;
  assign new_F5247_ = F5214 & ~F5215;
  assign new_F5248_ = ~new_F5230_ | new_F5240_;
  assign new_F5249_ = new_F5230_ & new_F5240_;
  assign new_F5250_ = ~new_F5230_ & ~new_F5240_;
  assign new_F5251_ = new_F5272_ | new_F5271_;
  assign new_F5252_ = F5218 | new_F5251_;
  assign new_F5253_ = new_F5276_ | new_F5275_;
  assign new_F5254_ = ~F5218 & new_F5253_;
  assign new_F5255_ = new_F5274_ | new_F5273_;
  assign new_F5256_ = F5218 & new_F5255_;
  assign new_F5257_ = F5216 & ~new_F5226_;
  assign new_F5258_ = ~F5216 & new_F5226_;
  assign new_F5259_ = ~F5215 | ~new_F5240_;
  assign new_F5260_ = new_F5226_ & new_F5259_;
  assign new_F5261_ = ~new_F5226_ & ~new_F5260_;
  assign new_F5262_ = new_F5226_ | new_F5259_;
  assign new_F5263_ = ~F5216 & F5217;
  assign new_F5264_ = F5216 & ~F5217;
  assign new_F5265_ = new_F5233_ | new_F5270_;
  assign new_F5266_ = ~new_F5233_ & ~new_F5269_;
  assign new_F5267_ = F5216 | new_F5233_;
  assign new_F5268_ = F5216 | F5217;
  assign new_F5269_ = new_F5233_ & new_F5270_;
  assign new_F5270_ = ~F5215 | ~new_F5240_;
  assign new_F5271_ = new_F5248_ & new_F5268_;
  assign new_F5272_ = ~new_F5248_ & ~new_F5268_;
  assign new_F5273_ = new_F5277_ | new_F5278_;
  assign new_F5274_ = ~F5219 & new_F5233_;
  assign new_F5275_ = new_F5279_ | new_F5280_;
  assign new_F5276_ = F5219 & new_F5233_;
  assign new_F5277_ = ~F5219 & ~new_F5233_;
  assign new_F5278_ = F5219 & ~new_F5233_;
  assign new_F5279_ = F5219 & ~new_F5233_;
  assign new_F5280_ = ~F5219 & new_F5233_;
  assign new_F5287_ = new_F5294_ & new_F5293_;
  assign new_F5288_ = new_F5296_ | new_F5295_;
  assign new_F5289_ = new_F5298_ | new_F5297_;
  assign new_F5290_ = new_F5300_ & new_F5299_;
  assign new_F5291_ = new_F5300_ & new_F5301_;
  assign new_F5292_ = new_F5293_ | new_F5302_;
  assign new_F5293_ = F5282 | new_F5305_;
  assign new_F5294_ = new_F5304_ | new_F5303_;
  assign new_F5295_ = new_F5309_ & new_F5308_;
  assign new_F5296_ = new_F5307_ & new_F5306_;
  assign new_F5297_ = new_F5312_ | new_F5311_;
  assign new_F5298_ = new_F5307_ & new_F5310_;
  assign new_F5299_ = F5282 | new_F5315_;
  assign new_F5300_ = new_F5314_ | new_F5313_;
  assign new_F5301_ = new_F5317_ | new_F5316_;
  assign new_F5302_ = ~new_F5293_ & new_F5319_;
  assign new_F5303_ = ~new_F5295_ & new_F5307_;
  assign new_F5304_ = new_F5295_ & ~new_F5307_;
  assign new_F5305_ = F5281 & ~F5282;
  assign new_F5306_ = ~new_F5328_ | ~new_F5329_;
  assign new_F5307_ = new_F5321_ | new_F5323_;
  assign new_F5308_ = new_F5331_ | new_F5330_;
  assign new_F5309_ = new_F5325_ | new_F5324_;
  assign new_F5310_ = ~new_F5333_ | ~new_F5332_;
  assign new_F5311_ = ~new_F5334_ & new_F5335_;
  assign new_F5312_ = new_F5334_ & ~new_F5335_;
  assign new_F5313_ = ~F5281 & F5282;
  assign new_F5314_ = F5281 & ~F5282;
  assign new_F5315_ = ~new_F5297_ | new_F5307_;
  assign new_F5316_ = new_F5297_ & new_F5307_;
  assign new_F5317_ = ~new_F5297_ & ~new_F5307_;
  assign new_F5318_ = new_F5339_ | new_F5338_;
  assign new_F5319_ = F5285 | new_F5318_;
  assign new_F5320_ = new_F5343_ | new_F5342_;
  assign new_F5321_ = ~F5285 & new_F5320_;
  assign new_F5322_ = new_F5341_ | new_F5340_;
  assign new_F5323_ = F5285 & new_F5322_;
  assign new_F5324_ = F5283 & ~new_F5293_;
  assign new_F5325_ = ~F5283 & new_F5293_;
  assign new_F5326_ = ~F5282 | ~new_F5307_;
  assign new_F5327_ = new_F5293_ & new_F5326_;
  assign new_F5328_ = ~new_F5293_ & ~new_F5327_;
  assign new_F5329_ = new_F5293_ | new_F5326_;
  assign new_F5330_ = ~F5283 & F5284;
  assign new_F5331_ = F5283 & ~F5284;
  assign new_F5332_ = new_F5300_ | new_F5337_;
  assign new_F5333_ = ~new_F5300_ & ~new_F5336_;
  assign new_F5334_ = F5283 | new_F5300_;
  assign new_F5335_ = F5283 | F5284;
  assign new_F5336_ = new_F5300_ & new_F5337_;
  assign new_F5337_ = ~F5282 | ~new_F5307_;
  assign new_F5338_ = new_F5315_ & new_F5335_;
  assign new_F5339_ = ~new_F5315_ & ~new_F5335_;
  assign new_F5340_ = new_F5344_ | new_F5345_;
  assign new_F5341_ = ~F5286 & new_F5300_;
  assign new_F5342_ = new_F5346_ | new_F5347_;
  assign new_F5343_ = F5286 & new_F5300_;
  assign new_F5344_ = ~F5286 & ~new_F5300_;
  assign new_F5345_ = F5286 & ~new_F5300_;
  assign new_F5346_ = F5286 & ~new_F5300_;
  assign new_F5347_ = ~F5286 & new_F5300_;
  assign new_F5354_ = new_F5361_ & new_F5360_;
  assign new_F5355_ = new_F5363_ | new_F5362_;
  assign new_F5356_ = new_F5365_ | new_F5364_;
  assign new_F5357_ = new_F5367_ & new_F5366_;
  assign new_F5358_ = new_F5367_ & new_F5368_;
  assign new_F5359_ = new_F5360_ | new_F5369_;
  assign new_F5360_ = F5349 | new_F5372_;
  assign new_F5361_ = new_F5371_ | new_F5370_;
  assign new_F5362_ = new_F5376_ & new_F5375_;
  assign new_F5363_ = new_F5374_ & new_F5373_;
  assign new_F5364_ = new_F5379_ | new_F5378_;
  assign new_F5365_ = new_F5374_ & new_F5377_;
  assign new_F5366_ = F5349 | new_F5382_;
  assign new_F5367_ = new_F5381_ | new_F5380_;
  assign new_F5368_ = new_F5384_ | new_F5383_;
  assign new_F5369_ = ~new_F5360_ & new_F5386_;
  assign new_F5370_ = ~new_F5362_ & new_F5374_;
  assign new_F5371_ = new_F5362_ & ~new_F5374_;
  assign new_F5372_ = F5348 & ~F5349;
  assign new_F5373_ = ~new_F5395_ | ~new_F5396_;
  assign new_F5374_ = new_F5388_ | new_F5390_;
  assign new_F5375_ = new_F5398_ | new_F5397_;
  assign new_F5376_ = new_F5392_ | new_F5391_;
  assign new_F5377_ = ~new_F5400_ | ~new_F5399_;
  assign new_F5378_ = ~new_F5401_ & new_F5402_;
  assign new_F5379_ = new_F5401_ & ~new_F5402_;
  assign new_F5380_ = ~F5348 & F5349;
  assign new_F5381_ = F5348 & ~F5349;
  assign new_F5382_ = ~new_F5364_ | new_F5374_;
  assign new_F5383_ = new_F5364_ & new_F5374_;
  assign new_F5384_ = ~new_F5364_ & ~new_F5374_;
  assign new_F5385_ = new_F5406_ | new_F5405_;
  assign new_F5386_ = F5352 | new_F5385_;
  assign new_F5387_ = new_F5410_ | new_F5409_;
  assign new_F5388_ = ~F5352 & new_F5387_;
  assign new_F5389_ = new_F5408_ | new_F5407_;
  assign new_F5390_ = F5352 & new_F5389_;
  assign new_F5391_ = F5350 & ~new_F5360_;
  assign new_F5392_ = ~F5350 & new_F5360_;
  assign new_F5393_ = ~F5349 | ~new_F5374_;
  assign new_F5394_ = new_F5360_ & new_F5393_;
  assign new_F5395_ = ~new_F5360_ & ~new_F5394_;
  assign new_F5396_ = new_F5360_ | new_F5393_;
  assign new_F5397_ = ~F5350 & F5351;
  assign new_F5398_ = F5350 & ~F5351;
  assign new_F5399_ = new_F5367_ | new_F5404_;
  assign new_F5400_ = ~new_F5367_ & ~new_F5403_;
  assign new_F5401_ = F5350 | new_F5367_;
  assign new_F5402_ = F5350 | F5351;
  assign new_F5403_ = new_F5367_ & new_F5404_;
  assign new_F5404_ = ~F5349 | ~new_F5374_;
  assign new_F5405_ = new_F5382_ & new_F5402_;
  assign new_F5406_ = ~new_F5382_ & ~new_F5402_;
  assign new_F5407_ = new_F5411_ | new_F5412_;
  assign new_F5408_ = ~F5353 & new_F5367_;
  assign new_F5409_ = new_F5413_ | new_F5414_;
  assign new_F5410_ = F5353 & new_F5367_;
  assign new_F5411_ = ~F5353 & ~new_F5367_;
  assign new_F5412_ = F5353 & ~new_F5367_;
  assign new_F5413_ = F5353 & ~new_F5367_;
  assign new_F5414_ = ~F5353 & new_F5367_;
  assign new_F5421_ = new_F5428_ & new_F5427_;
  assign new_F5422_ = new_F5430_ | new_F5429_;
  assign new_F5423_ = new_F5432_ | new_F5431_;
  assign new_F5424_ = new_F5434_ & new_F5433_;
  assign new_F5425_ = new_F5434_ & new_F5435_;
  assign new_F5426_ = new_F5427_ | new_F5436_;
  assign new_F5427_ = F5416 | new_F5439_;
  assign new_F5428_ = new_F5438_ | new_F5437_;
  assign new_F5429_ = new_F5443_ & new_F5442_;
  assign new_F5430_ = new_F5441_ & new_F5440_;
  assign new_F5431_ = new_F5446_ | new_F5445_;
  assign new_F5432_ = new_F5441_ & new_F5444_;
  assign new_F5433_ = F5416 | new_F5449_;
  assign new_F5434_ = new_F5448_ | new_F5447_;
  assign new_F5435_ = new_F5451_ | new_F5450_;
  assign new_F5436_ = ~new_F5427_ & new_F5453_;
  assign new_F5437_ = ~new_F5429_ & new_F5441_;
  assign new_F5438_ = new_F5429_ & ~new_F5441_;
  assign new_F5439_ = F5415 & ~F5416;
  assign new_F5440_ = ~new_F5462_ | ~new_F5463_;
  assign new_F5441_ = new_F5455_ | new_F5457_;
  assign new_F5442_ = new_F5465_ | new_F5464_;
  assign new_F5443_ = new_F5459_ | new_F5458_;
  assign new_F5444_ = ~new_F5467_ | ~new_F5466_;
  assign new_F5445_ = ~new_F5468_ & new_F5469_;
  assign new_F5446_ = new_F5468_ & ~new_F5469_;
  assign new_F5447_ = ~F5415 & F5416;
  assign new_F5448_ = F5415 & ~F5416;
  assign new_F5449_ = ~new_F5431_ | new_F5441_;
  assign new_F5450_ = new_F5431_ & new_F5441_;
  assign new_F5451_ = ~new_F5431_ & ~new_F5441_;
  assign new_F5452_ = new_F5473_ | new_F5472_;
  assign new_F5453_ = F5419 | new_F5452_;
  assign new_F5454_ = new_F5477_ | new_F5476_;
  assign new_F5455_ = ~F5419 & new_F5454_;
  assign new_F5456_ = new_F5475_ | new_F5474_;
  assign new_F5457_ = F5419 & new_F5456_;
  assign new_F5458_ = F5417 & ~new_F5427_;
  assign new_F5459_ = ~F5417 & new_F5427_;
  assign new_F5460_ = ~F5416 | ~new_F5441_;
  assign new_F5461_ = new_F5427_ & new_F5460_;
  assign new_F5462_ = ~new_F5427_ & ~new_F5461_;
  assign new_F5463_ = new_F5427_ | new_F5460_;
  assign new_F5464_ = ~F5417 & F5418;
  assign new_F5465_ = F5417 & ~F5418;
  assign new_F5466_ = new_F5434_ | new_F5471_;
  assign new_F5467_ = ~new_F5434_ & ~new_F5470_;
  assign new_F5468_ = F5417 | new_F5434_;
  assign new_F5469_ = F5417 | F5418;
  assign new_F5470_ = new_F5434_ & new_F5471_;
  assign new_F5471_ = ~F5416 | ~new_F5441_;
  assign new_F5472_ = new_F5449_ & new_F5469_;
  assign new_F5473_ = ~new_F5449_ & ~new_F5469_;
  assign new_F5474_ = new_F5478_ | new_F5479_;
  assign new_F5475_ = ~F5420 & new_F5434_;
  assign new_F5476_ = new_F5480_ | new_F5481_;
  assign new_F5477_ = F5420 & new_F5434_;
  assign new_F5478_ = ~F5420 & ~new_F5434_;
  assign new_F5479_ = F5420 & ~new_F5434_;
  assign new_F5480_ = F5420 & ~new_F5434_;
  assign new_F5481_ = ~F5420 & new_F5434_;
  assign new_F5488_ = new_F5495_ & new_F5494_;
  assign new_F5489_ = new_F5497_ | new_F5496_;
  assign new_F5490_ = new_F5499_ | new_F5498_;
  assign new_F5491_ = new_F5501_ & new_F5500_;
  assign new_F5492_ = new_F5501_ & new_F5502_;
  assign new_F5493_ = new_F5494_ | new_F5503_;
  assign new_F5494_ = F5483 | new_F5506_;
  assign new_F5495_ = new_F5505_ | new_F5504_;
  assign new_F5496_ = new_F5510_ & new_F5509_;
  assign new_F5497_ = new_F5508_ & new_F5507_;
  assign new_F5498_ = new_F5513_ | new_F5512_;
  assign new_F5499_ = new_F5508_ & new_F5511_;
  assign new_F5500_ = F5483 | new_F5516_;
  assign new_F5501_ = new_F5515_ | new_F5514_;
  assign new_F5502_ = new_F5518_ | new_F5517_;
  assign new_F5503_ = ~new_F5494_ & new_F5520_;
  assign new_F5504_ = ~new_F5496_ & new_F5508_;
  assign new_F5505_ = new_F5496_ & ~new_F5508_;
  assign new_F5506_ = F5482 & ~F5483;
  assign new_F5507_ = ~new_F5529_ | ~new_F5530_;
  assign new_F5508_ = new_F5522_ | new_F5524_;
  assign new_F5509_ = new_F5532_ | new_F5531_;
  assign new_F5510_ = new_F5526_ | new_F5525_;
  assign new_F5511_ = ~new_F5534_ | ~new_F5533_;
  assign new_F5512_ = ~new_F5535_ & new_F5536_;
  assign new_F5513_ = new_F5535_ & ~new_F5536_;
  assign new_F5514_ = ~F5482 & F5483;
  assign new_F5515_ = F5482 & ~F5483;
  assign new_F5516_ = ~new_F5498_ | new_F5508_;
  assign new_F5517_ = new_F5498_ & new_F5508_;
  assign new_F5518_ = ~new_F5498_ & ~new_F5508_;
  assign new_F5519_ = new_F5540_ | new_F5539_;
  assign new_F5520_ = F5486 | new_F5519_;
  assign new_F5521_ = new_F5544_ | new_F5543_;
  assign new_F5522_ = ~F5486 & new_F5521_;
  assign new_F5523_ = new_F5542_ | new_F5541_;
  assign new_F5524_ = F5486 & new_F5523_;
  assign new_F5525_ = F5484 & ~new_F5494_;
  assign new_F5526_ = ~F5484 & new_F5494_;
  assign new_F5527_ = ~F5483 | ~new_F5508_;
  assign new_F5528_ = new_F5494_ & new_F5527_;
  assign new_F5529_ = ~new_F5494_ & ~new_F5528_;
  assign new_F5530_ = new_F5494_ | new_F5527_;
  assign new_F5531_ = ~F5484 & F5485;
  assign new_F5532_ = F5484 & ~F5485;
  assign new_F5533_ = new_F5501_ | new_F5538_;
  assign new_F5534_ = ~new_F5501_ & ~new_F5537_;
  assign new_F5535_ = F5484 | new_F5501_;
  assign new_F5536_ = F5484 | F5485;
  assign new_F5537_ = new_F5501_ & new_F5538_;
  assign new_F5538_ = ~F5483 | ~new_F5508_;
  assign new_F5539_ = new_F5516_ & new_F5536_;
  assign new_F5540_ = ~new_F5516_ & ~new_F5536_;
  assign new_F5541_ = new_F5545_ | new_F5546_;
  assign new_F5542_ = ~F5487 & new_F5501_;
  assign new_F5543_ = new_F5547_ | new_F5548_;
  assign new_F5544_ = F5487 & new_F5501_;
  assign new_F5545_ = ~F5487 & ~new_F5501_;
  assign new_F5546_ = F5487 & ~new_F5501_;
  assign new_F5547_ = F5487 & ~new_F5501_;
  assign new_F5548_ = ~F5487 & new_F5501_;
  assign new_F5555_ = new_F5562_ & new_F5561_;
  assign new_F5556_ = new_F5564_ | new_F5563_;
  assign new_F5557_ = new_F5566_ | new_F5565_;
  assign new_F5558_ = new_F5568_ & new_F5567_;
  assign new_F5559_ = new_F5568_ & new_F5569_;
  assign new_F5560_ = new_F5561_ | new_F5570_;
  assign new_F5561_ = F5550 | new_F5573_;
  assign new_F5562_ = new_F5572_ | new_F5571_;
  assign new_F5563_ = new_F5577_ & new_F5576_;
  assign new_F5564_ = new_F5575_ & new_F5574_;
  assign new_F5565_ = new_F5580_ | new_F5579_;
  assign new_F5566_ = new_F5575_ & new_F5578_;
  assign new_F5567_ = F5550 | new_F5583_;
  assign new_F5568_ = new_F5582_ | new_F5581_;
  assign new_F5569_ = new_F5585_ | new_F5584_;
  assign new_F5570_ = ~new_F5561_ & new_F5587_;
  assign new_F5571_ = ~new_F5563_ & new_F5575_;
  assign new_F5572_ = new_F5563_ & ~new_F5575_;
  assign new_F5573_ = F5549 & ~F5550;
  assign new_F5574_ = ~new_F5596_ | ~new_F5597_;
  assign new_F5575_ = new_F5589_ | new_F5591_;
  assign new_F5576_ = new_F5599_ | new_F5598_;
  assign new_F5577_ = new_F5593_ | new_F5592_;
  assign new_F5578_ = ~new_F5601_ | ~new_F5600_;
  assign new_F5579_ = ~new_F5602_ & new_F5603_;
  assign new_F5580_ = new_F5602_ & ~new_F5603_;
  assign new_F5581_ = ~F5549 & F5550;
  assign new_F5582_ = F5549 & ~F5550;
  assign new_F5583_ = ~new_F5565_ | new_F5575_;
  assign new_F5584_ = new_F5565_ & new_F5575_;
  assign new_F5585_ = ~new_F5565_ & ~new_F5575_;
  assign new_F5586_ = new_F5607_ | new_F5606_;
  assign new_F5587_ = F5553 | new_F5586_;
  assign new_F5588_ = new_F5611_ | new_F5610_;
  assign new_F5589_ = ~F5553 & new_F5588_;
  assign new_F5590_ = new_F5609_ | new_F5608_;
  assign new_F5591_ = F5553 & new_F5590_;
  assign new_F5592_ = F5551 & ~new_F5561_;
  assign new_F5593_ = ~F5551 & new_F5561_;
  assign new_F5594_ = ~F5550 | ~new_F5575_;
  assign new_F5595_ = new_F5561_ & new_F5594_;
  assign new_F5596_ = ~new_F5561_ & ~new_F5595_;
  assign new_F5597_ = new_F5561_ | new_F5594_;
  assign new_F5598_ = ~F5551 & F5552;
  assign new_F5599_ = F5551 & ~F5552;
  assign new_F5600_ = new_F5568_ | new_F5605_;
  assign new_F5601_ = ~new_F5568_ & ~new_F5604_;
  assign new_F5602_ = F5551 | new_F5568_;
  assign new_F5603_ = F5551 | F5552;
  assign new_F5604_ = new_F5568_ & new_F5605_;
  assign new_F5605_ = ~F5550 | ~new_F5575_;
  assign new_F5606_ = new_F5583_ & new_F5603_;
  assign new_F5607_ = ~new_F5583_ & ~new_F5603_;
  assign new_F5608_ = new_F5612_ | new_F5613_;
  assign new_F5609_ = ~F5554 & new_F5568_;
  assign new_F5610_ = new_F5614_ | new_F5615_;
  assign new_F5611_ = F5554 & new_F5568_;
  assign new_F5612_ = ~F5554 & ~new_F5568_;
  assign new_F5613_ = F5554 & ~new_F5568_;
  assign new_F5614_ = F5554 & ~new_F5568_;
  assign new_F5615_ = ~F5554 & new_F5568_;
  assign new_F5622_ = new_F5629_ & new_F5628_;
  assign new_F5623_ = new_F5631_ | new_F5630_;
  assign new_F5624_ = new_F5633_ | new_F5632_;
  assign new_F5625_ = new_F5635_ & new_F5634_;
  assign new_F5626_ = new_F5635_ & new_F5636_;
  assign new_F5627_ = new_F5628_ | new_F5637_;
  assign new_F5628_ = F5617 | new_F5640_;
  assign new_F5629_ = new_F5639_ | new_F5638_;
  assign new_F5630_ = new_F5644_ & new_F5643_;
  assign new_F5631_ = new_F5642_ & new_F5641_;
  assign new_F5632_ = new_F5647_ | new_F5646_;
  assign new_F5633_ = new_F5642_ & new_F5645_;
  assign new_F5634_ = F5617 | new_F5650_;
  assign new_F5635_ = new_F5649_ | new_F5648_;
  assign new_F5636_ = new_F5652_ | new_F5651_;
  assign new_F5637_ = ~new_F5628_ & new_F5654_;
  assign new_F5638_ = ~new_F5630_ & new_F5642_;
  assign new_F5639_ = new_F5630_ & ~new_F5642_;
  assign new_F5640_ = F5616 & ~F5617;
  assign new_F5641_ = ~new_F5663_ | ~new_F5664_;
  assign new_F5642_ = new_F5656_ | new_F5658_;
  assign new_F5643_ = new_F5666_ | new_F5665_;
  assign new_F5644_ = new_F5660_ | new_F5659_;
  assign new_F5645_ = ~new_F5668_ | ~new_F5667_;
  assign new_F5646_ = ~new_F5669_ & new_F5670_;
  assign new_F5647_ = new_F5669_ & ~new_F5670_;
  assign new_F5648_ = ~F5616 & F5617;
  assign new_F5649_ = F5616 & ~F5617;
  assign new_F5650_ = ~new_F5632_ | new_F5642_;
  assign new_F5651_ = new_F5632_ & new_F5642_;
  assign new_F5652_ = ~new_F5632_ & ~new_F5642_;
  assign new_F5653_ = new_F5674_ | new_F5673_;
  assign new_F5654_ = F5620 | new_F5653_;
  assign new_F5655_ = new_F5678_ | new_F5677_;
  assign new_F5656_ = ~F5620 & new_F5655_;
  assign new_F5657_ = new_F5676_ | new_F5675_;
  assign new_F5658_ = F5620 & new_F5657_;
  assign new_F5659_ = F5618 & ~new_F5628_;
  assign new_F5660_ = ~F5618 & new_F5628_;
  assign new_F5661_ = ~F5617 | ~new_F5642_;
  assign new_F5662_ = new_F5628_ & new_F5661_;
  assign new_F5663_ = ~new_F5628_ & ~new_F5662_;
  assign new_F5664_ = new_F5628_ | new_F5661_;
  assign new_F5665_ = ~F5618 & F5619;
  assign new_F5666_ = F5618 & ~F5619;
  assign new_F5667_ = new_F5635_ | new_F5672_;
  assign new_F5668_ = ~new_F5635_ & ~new_F5671_;
  assign new_F5669_ = F5618 | new_F5635_;
  assign new_F5670_ = F5618 | F5619;
  assign new_F5671_ = new_F5635_ & new_F5672_;
  assign new_F5672_ = ~F5617 | ~new_F5642_;
  assign new_F5673_ = new_F5650_ & new_F5670_;
  assign new_F5674_ = ~new_F5650_ & ~new_F5670_;
  assign new_F5675_ = new_F5679_ | new_F5680_;
  assign new_F5676_ = ~F5621 & new_F5635_;
  assign new_F5677_ = new_F5681_ | new_F5682_;
  assign new_F5678_ = F5621 & new_F5635_;
  assign new_F5679_ = ~F5621 & ~new_F5635_;
  assign new_F5680_ = F5621 & ~new_F5635_;
  assign new_F5681_ = F5621 & ~new_F5635_;
  assign new_F5682_ = ~F5621 & new_F5635_;
  assign new_F5689_ = new_F5696_ & new_F5695_;
  assign new_F5690_ = new_F5698_ | new_F5697_;
  assign new_F5691_ = new_F5700_ | new_F5699_;
  assign new_F5692_ = new_F5702_ & new_F5701_;
  assign new_F5693_ = new_F5702_ & new_F5703_;
  assign new_F5694_ = new_F5695_ | new_F5704_;
  assign new_F5695_ = F5684 | new_F5707_;
  assign new_F5696_ = new_F5706_ | new_F5705_;
  assign new_F5697_ = new_F5711_ & new_F5710_;
  assign new_F5698_ = new_F5709_ & new_F5708_;
  assign new_F5699_ = new_F5714_ | new_F5713_;
  assign new_F5700_ = new_F5709_ & new_F5712_;
  assign new_F5701_ = F5684 | new_F5717_;
  assign new_F5702_ = new_F5716_ | new_F5715_;
  assign new_F5703_ = new_F5719_ | new_F5718_;
  assign new_F5704_ = ~new_F5695_ & new_F5721_;
  assign new_F5705_ = ~new_F5697_ & new_F5709_;
  assign new_F5706_ = new_F5697_ & ~new_F5709_;
  assign new_F5707_ = F5683 & ~F5684;
  assign new_F5708_ = ~new_F5730_ | ~new_F5731_;
  assign new_F5709_ = new_F5723_ | new_F5725_;
  assign new_F5710_ = new_F5733_ | new_F5732_;
  assign new_F5711_ = new_F5727_ | new_F5726_;
  assign new_F5712_ = ~new_F5735_ | ~new_F5734_;
  assign new_F5713_ = ~new_F5736_ & new_F5737_;
  assign new_F5714_ = new_F5736_ & ~new_F5737_;
  assign new_F5715_ = ~F5683 & F5684;
  assign new_F5716_ = F5683 & ~F5684;
  assign new_F5717_ = ~new_F5699_ | new_F5709_;
  assign new_F5718_ = new_F5699_ & new_F5709_;
  assign new_F5719_ = ~new_F5699_ & ~new_F5709_;
  assign new_F5720_ = new_F5741_ | new_F5740_;
  assign new_F5721_ = F5687 | new_F5720_;
  assign new_F5722_ = new_F5745_ | new_F5744_;
  assign new_F5723_ = ~F5687 & new_F5722_;
  assign new_F5724_ = new_F5743_ | new_F5742_;
  assign new_F5725_ = F5687 & new_F5724_;
  assign new_F5726_ = F5685 & ~new_F5695_;
  assign new_F5727_ = ~F5685 & new_F5695_;
  assign new_F5728_ = ~F5684 | ~new_F5709_;
  assign new_F5729_ = new_F5695_ & new_F5728_;
  assign new_F5730_ = ~new_F5695_ & ~new_F5729_;
  assign new_F5731_ = new_F5695_ | new_F5728_;
  assign new_F5732_ = ~F5685 & F5686;
  assign new_F5733_ = F5685 & ~F5686;
  assign new_F5734_ = new_F5702_ | new_F5739_;
  assign new_F5735_ = ~new_F5702_ & ~new_F5738_;
  assign new_F5736_ = F5685 | new_F5702_;
  assign new_F5737_ = F5685 | F5686;
  assign new_F5738_ = new_F5702_ & new_F5739_;
  assign new_F5739_ = ~F5684 | ~new_F5709_;
  assign new_F5740_ = new_F5717_ & new_F5737_;
  assign new_F5741_ = ~new_F5717_ & ~new_F5737_;
  assign new_F5742_ = new_F5746_ | new_F5747_;
  assign new_F5743_ = ~F5688 & new_F5702_;
  assign new_F5744_ = new_F5748_ | new_F5749_;
  assign new_F5745_ = F5688 & new_F5702_;
  assign new_F5746_ = ~F5688 & ~new_F5702_;
  assign new_F5747_ = F5688 & ~new_F5702_;
  assign new_F5748_ = F5688 & ~new_F5702_;
  assign new_F5749_ = ~F5688 & new_F5702_;
  assign new_F5756_ = new_F5763_ & new_F5762_;
  assign new_F5757_ = new_F5765_ | new_F5764_;
  assign new_F5758_ = new_F5767_ | new_F5766_;
  assign new_F5759_ = new_F5769_ & new_F5768_;
  assign new_F5760_ = new_F5769_ & new_F5770_;
  assign new_F5761_ = new_F5762_ | new_F5771_;
  assign new_F5762_ = F5751 | new_F5774_;
  assign new_F5763_ = new_F5773_ | new_F5772_;
  assign new_F5764_ = new_F5778_ & new_F5777_;
  assign new_F5765_ = new_F5776_ & new_F5775_;
  assign new_F5766_ = new_F5781_ | new_F5780_;
  assign new_F5767_ = new_F5776_ & new_F5779_;
  assign new_F5768_ = F5751 | new_F5784_;
  assign new_F5769_ = new_F5783_ | new_F5782_;
  assign new_F5770_ = new_F5786_ | new_F5785_;
  assign new_F5771_ = ~new_F5762_ & new_F5788_;
  assign new_F5772_ = ~new_F5764_ & new_F5776_;
  assign new_F5773_ = new_F5764_ & ~new_F5776_;
  assign new_F5774_ = F5750 & ~F5751;
  assign new_F5775_ = ~new_F5797_ | ~new_F5798_;
  assign new_F5776_ = new_F5790_ | new_F5792_;
  assign new_F5777_ = new_F5800_ | new_F5799_;
  assign new_F5778_ = new_F5794_ | new_F5793_;
  assign new_F5779_ = ~new_F5802_ | ~new_F5801_;
  assign new_F5780_ = ~new_F5803_ & new_F5804_;
  assign new_F5781_ = new_F5803_ & ~new_F5804_;
  assign new_F5782_ = ~F5750 & F5751;
  assign new_F5783_ = F5750 & ~F5751;
  assign new_F5784_ = ~new_F5766_ | new_F5776_;
  assign new_F5785_ = new_F5766_ & new_F5776_;
  assign new_F5786_ = ~new_F5766_ & ~new_F5776_;
  assign new_F5787_ = new_F5808_ | new_F5807_;
  assign new_F5788_ = F5754 | new_F5787_;
  assign new_F5789_ = new_F5812_ | new_F5811_;
  assign new_F5790_ = ~F5754 & new_F5789_;
  assign new_F5791_ = new_F5810_ | new_F5809_;
  assign new_F5792_ = F5754 & new_F5791_;
  assign new_F5793_ = F5752 & ~new_F5762_;
  assign new_F5794_ = ~F5752 & new_F5762_;
  assign new_F5795_ = ~F5751 | ~new_F5776_;
  assign new_F5796_ = new_F5762_ & new_F5795_;
  assign new_F5797_ = ~new_F5762_ & ~new_F5796_;
  assign new_F5798_ = new_F5762_ | new_F5795_;
  assign new_F5799_ = ~F5752 & F5753;
  assign new_F5800_ = F5752 & ~F5753;
  assign new_F5801_ = new_F5769_ | new_F5806_;
  assign new_F5802_ = ~new_F5769_ & ~new_F5805_;
  assign new_F5803_ = F5752 | new_F5769_;
  assign new_F5804_ = F5752 | F5753;
  assign new_F5805_ = new_F5769_ & new_F5806_;
  assign new_F5806_ = ~F5751 | ~new_F5776_;
  assign new_F5807_ = new_F5784_ & new_F5804_;
  assign new_F5808_ = ~new_F5784_ & ~new_F5804_;
  assign new_F5809_ = new_F5813_ | new_F5814_;
  assign new_F5810_ = ~F5755 & new_F5769_;
  assign new_F5811_ = new_F5815_ | new_F5816_;
  assign new_F5812_ = F5755 & new_F5769_;
  assign new_F5813_ = ~F5755 & ~new_F5769_;
  assign new_F5814_ = F5755 & ~new_F5769_;
  assign new_F5815_ = F5755 & ~new_F5769_;
  assign new_F5816_ = ~F5755 & new_F5769_;
  assign new_F5823_ = new_F5830_ & new_F5829_;
  assign new_F5824_ = new_F5832_ | new_F5831_;
  assign new_F5825_ = new_F5834_ | new_F5833_;
  assign new_F5826_ = new_F5836_ & new_F5835_;
  assign new_F5827_ = new_F5836_ & new_F5837_;
  assign new_F5828_ = new_F5829_ | new_F5838_;
  assign new_F5829_ = F5818 | new_F5841_;
  assign new_F5830_ = new_F5840_ | new_F5839_;
  assign new_F5831_ = new_F5845_ & new_F5844_;
  assign new_F5832_ = new_F5843_ & new_F5842_;
  assign new_F5833_ = new_F5848_ | new_F5847_;
  assign new_F5834_ = new_F5843_ & new_F5846_;
  assign new_F5835_ = F5818 | new_F5851_;
  assign new_F5836_ = new_F5850_ | new_F5849_;
  assign new_F5837_ = new_F5853_ | new_F5852_;
  assign new_F5838_ = ~new_F5829_ & new_F5855_;
  assign new_F5839_ = ~new_F5831_ & new_F5843_;
  assign new_F5840_ = new_F5831_ & ~new_F5843_;
  assign new_F5841_ = F5817 & ~F5818;
  assign new_F5842_ = ~new_F5864_ | ~new_F5865_;
  assign new_F5843_ = new_F5857_ | new_F5859_;
  assign new_F5844_ = new_F5867_ | new_F5866_;
  assign new_F5845_ = new_F5861_ | new_F5860_;
  assign new_F5846_ = ~new_F5869_ | ~new_F5868_;
  assign new_F5847_ = ~new_F5870_ & new_F5871_;
  assign new_F5848_ = new_F5870_ & ~new_F5871_;
  assign new_F5849_ = ~F5817 & F5818;
  assign new_F5850_ = F5817 & ~F5818;
  assign new_F5851_ = ~new_F5833_ | new_F5843_;
  assign new_F5852_ = new_F5833_ & new_F5843_;
  assign new_F5853_ = ~new_F5833_ & ~new_F5843_;
  assign new_F5854_ = new_F5875_ | new_F5874_;
  assign new_F5855_ = F5821 | new_F5854_;
  assign new_F5856_ = new_F5879_ | new_F5878_;
  assign new_F5857_ = ~F5821 & new_F5856_;
  assign new_F5858_ = new_F5877_ | new_F5876_;
  assign new_F5859_ = F5821 & new_F5858_;
  assign new_F5860_ = F5819 & ~new_F5829_;
  assign new_F5861_ = ~F5819 & new_F5829_;
  assign new_F5862_ = ~F5818 | ~new_F5843_;
  assign new_F5863_ = new_F5829_ & new_F5862_;
  assign new_F5864_ = ~new_F5829_ & ~new_F5863_;
  assign new_F5865_ = new_F5829_ | new_F5862_;
  assign new_F5866_ = ~F5819 & F5820;
  assign new_F5867_ = F5819 & ~F5820;
  assign new_F5868_ = new_F5836_ | new_F5873_;
  assign new_F5869_ = ~new_F5836_ & ~new_F5872_;
  assign new_F5870_ = F5819 | new_F5836_;
  assign new_F5871_ = F5819 | F5820;
  assign new_F5872_ = new_F5836_ & new_F5873_;
  assign new_F5873_ = ~F5818 | ~new_F5843_;
  assign new_F5874_ = new_F5851_ & new_F5871_;
  assign new_F5875_ = ~new_F5851_ & ~new_F5871_;
  assign new_F5876_ = new_F5880_ | new_F5881_;
  assign new_F5877_ = ~F5822 & new_F5836_;
  assign new_F5878_ = new_F5882_ | new_F5883_;
  assign new_F5879_ = F5822 & new_F5836_;
  assign new_F5880_ = ~F5822 & ~new_F5836_;
  assign new_F5881_ = F5822 & ~new_F5836_;
  assign new_F5882_ = F5822 & ~new_F5836_;
  assign new_F5883_ = ~F5822 & new_F5836_;
  assign new_F5890_ = new_F5897_ & new_F5896_;
  assign new_F5891_ = new_F5899_ | new_F5898_;
  assign new_F5892_ = new_F5901_ | new_F5900_;
  assign new_F5893_ = new_F5903_ & new_F5902_;
  assign new_F5894_ = new_F5903_ & new_F5904_;
  assign new_F5895_ = new_F5896_ | new_F5905_;
  assign new_F5896_ = F5885 | new_F5908_;
  assign new_F5897_ = new_F5907_ | new_F5906_;
  assign new_F5898_ = new_F5912_ & new_F5911_;
  assign new_F5899_ = new_F5910_ & new_F5909_;
  assign new_F5900_ = new_F5915_ | new_F5914_;
  assign new_F5901_ = new_F5910_ & new_F5913_;
  assign new_F5902_ = F5885 | new_F5918_;
  assign new_F5903_ = new_F5917_ | new_F5916_;
  assign new_F5904_ = new_F5920_ | new_F5919_;
  assign new_F5905_ = ~new_F5896_ & new_F5922_;
  assign new_F5906_ = ~new_F5898_ & new_F5910_;
  assign new_F5907_ = new_F5898_ & ~new_F5910_;
  assign new_F5908_ = F5884 & ~F5885;
  assign new_F5909_ = ~new_F5931_ | ~new_F5932_;
  assign new_F5910_ = new_F5924_ | new_F5926_;
  assign new_F5911_ = new_F5934_ | new_F5933_;
  assign new_F5912_ = new_F5928_ | new_F5927_;
  assign new_F5913_ = ~new_F5936_ | ~new_F5935_;
  assign new_F5914_ = ~new_F5937_ & new_F5938_;
  assign new_F5915_ = new_F5937_ & ~new_F5938_;
  assign new_F5916_ = ~F5884 & F5885;
  assign new_F5917_ = F5884 & ~F5885;
  assign new_F5918_ = ~new_F5900_ | new_F5910_;
  assign new_F5919_ = new_F5900_ & new_F5910_;
  assign new_F5920_ = ~new_F5900_ & ~new_F5910_;
  assign new_F5921_ = new_F5942_ | new_F5941_;
  assign new_F5922_ = F5888 | new_F5921_;
  assign new_F5923_ = new_F5946_ | new_F5945_;
  assign new_F5924_ = ~F5888 & new_F5923_;
  assign new_F5925_ = new_F5944_ | new_F5943_;
  assign new_F5926_ = F5888 & new_F5925_;
  assign new_F5927_ = F5886 & ~new_F5896_;
  assign new_F5928_ = ~F5886 & new_F5896_;
  assign new_F5929_ = ~F5885 | ~new_F5910_;
  assign new_F5930_ = new_F5896_ & new_F5929_;
  assign new_F5931_ = ~new_F5896_ & ~new_F5930_;
  assign new_F5932_ = new_F5896_ | new_F5929_;
  assign new_F5933_ = ~F5886 & F5887;
  assign new_F5934_ = F5886 & ~F5887;
  assign new_F5935_ = new_F5903_ | new_F5940_;
  assign new_F5936_ = ~new_F5903_ & ~new_F5939_;
  assign new_F5937_ = F5886 | new_F5903_;
  assign new_F5938_ = F5886 | F5887;
  assign new_F5939_ = new_F5903_ & new_F5940_;
  assign new_F5940_ = ~F5885 | ~new_F5910_;
  assign new_F5941_ = new_F5918_ & new_F5938_;
  assign new_F5942_ = ~new_F5918_ & ~new_F5938_;
  assign new_F5943_ = new_F5947_ | new_F5948_;
  assign new_F5944_ = ~F5889 & new_F5903_;
  assign new_F5945_ = new_F5949_ | new_F5950_;
  assign new_F5946_ = F5889 & new_F5903_;
  assign new_F5947_ = ~F5889 & ~new_F5903_;
  assign new_F5948_ = F5889 & ~new_F5903_;
  assign new_F5949_ = F5889 & ~new_F5903_;
  assign new_F5950_ = ~F5889 & new_F5903_;
  assign new_F5957_ = new_F5964_ & new_F5963_;
  assign new_F5958_ = new_F5966_ | new_F5965_;
  assign new_F5959_ = new_F5968_ | new_F5967_;
  assign new_F5960_ = new_F5970_ & new_F5969_;
  assign new_F5961_ = new_F5970_ & new_F5971_;
  assign new_F5962_ = new_F5963_ | new_F5972_;
  assign new_F5963_ = F5952 | new_F5975_;
  assign new_F5964_ = new_F5974_ | new_F5973_;
  assign new_F5965_ = new_F5979_ & new_F5978_;
  assign new_F5966_ = new_F5977_ & new_F5976_;
  assign new_F5967_ = new_F5982_ | new_F5981_;
  assign new_F5968_ = new_F5977_ & new_F5980_;
  assign new_F5969_ = F5952 | new_F5985_;
  assign new_F5970_ = new_F5984_ | new_F5983_;
  assign new_F5971_ = new_F5987_ | new_F5986_;
  assign new_F5972_ = ~new_F5963_ & new_F5989_;
  assign new_F5973_ = ~new_F5965_ & new_F5977_;
  assign new_F5974_ = new_F5965_ & ~new_F5977_;
  assign new_F5975_ = F5951 & ~F5952;
  assign new_F5976_ = ~new_F5998_ | ~new_F5999_;
  assign new_F5977_ = new_F5991_ | new_F5993_;
  assign new_F5978_ = new_F6001_ | new_F6000_;
  assign new_F5979_ = new_F5995_ | new_F5994_;
  assign new_F5980_ = ~new_F6003_ | ~new_F6002_;
  assign new_F5981_ = ~new_F6004_ & new_F6005_;
  assign new_F5982_ = new_F6004_ & ~new_F6005_;
  assign new_F5983_ = ~F5951 & F5952;
  assign new_F5984_ = F5951 & ~F5952;
  assign new_F5985_ = ~new_F5967_ | new_F5977_;
  assign new_F5986_ = new_F5967_ & new_F5977_;
  assign new_F5987_ = ~new_F5967_ & ~new_F5977_;
  assign new_F5988_ = new_F6009_ | new_F6008_;
  assign new_F5989_ = F5955 | new_F5988_;
  assign new_F5990_ = new_F6013_ | new_F6012_;
  assign new_F5991_ = ~F5955 & new_F5990_;
  assign new_F5992_ = new_F6011_ | new_F6010_;
  assign new_F5993_ = F5955 & new_F5992_;
  assign new_F5994_ = F5953 & ~new_F5963_;
  assign new_F5995_ = ~F5953 & new_F5963_;
  assign new_F5996_ = ~F5952 | ~new_F5977_;
  assign new_F5997_ = new_F5963_ & new_F5996_;
  assign new_F5998_ = ~new_F5963_ & ~new_F5997_;
  assign new_F5999_ = new_F5963_ | new_F5996_;
  assign new_F6000_ = ~F5953 & F5954;
  assign new_F6001_ = F5953 & ~F5954;
  assign new_F6002_ = new_F5970_ | new_F6007_;
  assign new_F6003_ = ~new_F5970_ & ~new_F6006_;
  assign new_F6004_ = F5953 | new_F5970_;
  assign new_F6005_ = F5953 | F5954;
  assign new_F6006_ = new_F5970_ & new_F6007_;
  assign new_F6007_ = ~F5952 | ~new_F5977_;
  assign new_F6008_ = new_F5985_ & new_F6005_;
  assign new_F6009_ = ~new_F5985_ & ~new_F6005_;
  assign new_F6010_ = new_F6014_ | new_F6015_;
  assign new_F6011_ = ~F5956 & new_F5970_;
  assign new_F6012_ = new_F6016_ | new_F6017_;
  assign new_F6013_ = F5956 & new_F5970_;
  assign new_F6014_ = ~F5956 & ~new_F5970_;
  assign new_F6015_ = F5956 & ~new_F5970_;
  assign new_F6016_ = F5956 & ~new_F5970_;
  assign new_F6017_ = ~F5956 & new_F5970_;
  assign new_F6024_ = new_F6031_ & new_F6030_;
  assign new_F6025_ = new_F6033_ | new_F6032_;
  assign new_F6026_ = new_F6035_ | new_F6034_;
  assign new_F6027_ = new_F6037_ & new_F6036_;
  assign new_F6028_ = new_F6037_ & new_F6038_;
  assign new_F6029_ = new_F6030_ | new_F6039_;
  assign new_F6030_ = F6019 | new_F6042_;
  assign new_F6031_ = new_F6041_ | new_F6040_;
  assign new_F6032_ = new_F6046_ & new_F6045_;
  assign new_F6033_ = new_F6044_ & new_F6043_;
  assign new_F6034_ = new_F6049_ | new_F6048_;
  assign new_F6035_ = new_F6044_ & new_F6047_;
  assign new_F6036_ = F6019 | new_F6052_;
  assign new_F6037_ = new_F6051_ | new_F6050_;
  assign new_F6038_ = new_F6054_ | new_F6053_;
  assign new_F6039_ = ~new_F6030_ & new_F6056_;
  assign new_F6040_ = ~new_F6032_ & new_F6044_;
  assign new_F6041_ = new_F6032_ & ~new_F6044_;
  assign new_F6042_ = F6018 & ~F6019;
  assign new_F6043_ = ~new_F6065_ | ~new_F6066_;
  assign new_F6044_ = new_F6058_ | new_F6060_;
  assign new_F6045_ = new_F6068_ | new_F6067_;
  assign new_F6046_ = new_F6062_ | new_F6061_;
  assign new_F6047_ = ~new_F6070_ | ~new_F6069_;
  assign new_F6048_ = ~new_F6071_ & new_F6072_;
  assign new_F6049_ = new_F6071_ & ~new_F6072_;
  assign new_F6050_ = ~F6018 & F6019;
  assign new_F6051_ = F6018 & ~F6019;
  assign new_F6052_ = ~new_F6034_ | new_F6044_;
  assign new_F6053_ = new_F6034_ & new_F6044_;
  assign new_F6054_ = ~new_F6034_ & ~new_F6044_;
  assign new_F6055_ = new_F6076_ | new_F6075_;
  assign new_F6056_ = F6022 | new_F6055_;
  assign new_F6057_ = new_F6080_ | new_F6079_;
  assign new_F6058_ = ~F6022 & new_F6057_;
  assign new_F6059_ = new_F6078_ | new_F6077_;
  assign new_F6060_ = F6022 & new_F6059_;
  assign new_F6061_ = F6020 & ~new_F6030_;
  assign new_F6062_ = ~F6020 & new_F6030_;
  assign new_F6063_ = ~F6019 | ~new_F6044_;
  assign new_F6064_ = new_F6030_ & new_F6063_;
  assign new_F6065_ = ~new_F6030_ & ~new_F6064_;
  assign new_F6066_ = new_F6030_ | new_F6063_;
  assign new_F6067_ = ~F6020 & F6021;
  assign new_F6068_ = F6020 & ~F6021;
  assign new_F6069_ = new_F6037_ | new_F6074_;
  assign new_F6070_ = ~new_F6037_ & ~new_F6073_;
  assign new_F6071_ = F6020 | new_F6037_;
  assign new_F6072_ = F6020 | F6021;
  assign new_F6073_ = new_F6037_ & new_F6074_;
  assign new_F6074_ = ~F6019 | ~new_F6044_;
  assign new_F6075_ = new_F6052_ & new_F6072_;
  assign new_F6076_ = ~new_F6052_ & ~new_F6072_;
  assign new_F6077_ = new_F6081_ | new_F6082_;
  assign new_F6078_ = ~F6023 & new_F6037_;
  assign new_F6079_ = new_F6083_ | new_F6084_;
  assign new_F6080_ = F6023 & new_F6037_;
  assign new_F6081_ = ~F6023 & ~new_F6037_;
  assign new_F6082_ = F6023 & ~new_F6037_;
  assign new_F6083_ = F6023 & ~new_F6037_;
  assign new_F6084_ = ~F6023 & new_F6037_;
  assign new_F6091_ = new_F6098_ & new_F6097_;
  assign new_F6092_ = new_F6100_ | new_F6099_;
  assign new_F6093_ = new_F6102_ | new_F6101_;
  assign new_F6094_ = new_F6104_ & new_F6103_;
  assign new_F6095_ = new_F6104_ & new_F6105_;
  assign new_F6096_ = new_F6097_ | new_F6106_;
  assign new_F6097_ = F6086 | new_F6109_;
  assign new_F6098_ = new_F6108_ | new_F6107_;
  assign new_F6099_ = new_F6113_ & new_F6112_;
  assign new_F6100_ = new_F6111_ & new_F6110_;
  assign new_F6101_ = new_F6116_ | new_F6115_;
  assign new_F6102_ = new_F6111_ & new_F6114_;
  assign new_F6103_ = F6086 | new_F6119_;
  assign new_F6104_ = new_F6118_ | new_F6117_;
  assign new_F6105_ = new_F6121_ | new_F6120_;
  assign new_F6106_ = ~new_F6097_ & new_F6123_;
  assign new_F6107_ = ~new_F6099_ & new_F6111_;
  assign new_F6108_ = new_F6099_ & ~new_F6111_;
  assign new_F6109_ = F6085 & ~F6086;
  assign new_F6110_ = ~new_F6132_ | ~new_F6133_;
  assign new_F6111_ = new_F6125_ | new_F6127_;
  assign new_F6112_ = new_F6135_ | new_F6134_;
  assign new_F6113_ = new_F6129_ | new_F6128_;
  assign new_F6114_ = ~new_F6137_ | ~new_F6136_;
  assign new_F6115_ = ~new_F6138_ & new_F6139_;
  assign new_F6116_ = new_F6138_ & ~new_F6139_;
  assign new_F6117_ = ~F6085 & F6086;
  assign new_F6118_ = F6085 & ~F6086;
  assign new_F6119_ = ~new_F6101_ | new_F6111_;
  assign new_F6120_ = new_F6101_ & new_F6111_;
  assign new_F6121_ = ~new_F6101_ & ~new_F6111_;
  assign new_F6122_ = new_F6143_ | new_F6142_;
  assign new_F6123_ = F6089 | new_F6122_;
  assign new_F6124_ = new_F6147_ | new_F6146_;
  assign new_F6125_ = ~F6089 & new_F6124_;
  assign new_F6126_ = new_F6145_ | new_F6144_;
  assign new_F6127_ = F6089 & new_F6126_;
  assign new_F6128_ = F6087 & ~new_F6097_;
  assign new_F6129_ = ~F6087 & new_F6097_;
  assign new_F6130_ = ~F6086 | ~new_F6111_;
  assign new_F6131_ = new_F6097_ & new_F6130_;
  assign new_F6132_ = ~new_F6097_ & ~new_F6131_;
  assign new_F6133_ = new_F6097_ | new_F6130_;
  assign new_F6134_ = ~F6087 & F6088;
  assign new_F6135_ = F6087 & ~F6088;
  assign new_F6136_ = new_F6104_ | new_F6141_;
  assign new_F6137_ = ~new_F6104_ & ~new_F6140_;
  assign new_F6138_ = F6087 | new_F6104_;
  assign new_F6139_ = F6087 | F6088;
  assign new_F6140_ = new_F6104_ & new_F6141_;
  assign new_F6141_ = ~F6086 | ~new_F6111_;
  assign new_F6142_ = new_F6119_ & new_F6139_;
  assign new_F6143_ = ~new_F6119_ & ~new_F6139_;
  assign new_F6144_ = new_F6148_ | new_F6149_;
  assign new_F6145_ = ~F6090 & new_F6104_;
  assign new_F6146_ = new_F6150_ | new_F6151_;
  assign new_F6147_ = F6090 & new_F6104_;
  assign new_F6148_ = ~F6090 & ~new_F6104_;
  assign new_F6149_ = F6090 & ~new_F6104_;
  assign new_F6150_ = F6090 & ~new_F6104_;
  assign new_F6151_ = ~F6090 & new_F6104_;
  assign new_F6158_ = new_F6165_ & new_F6164_;
  assign new_F6159_ = new_F6167_ | new_F6166_;
  assign new_F6160_ = new_F6169_ | new_F6168_;
  assign new_F6161_ = new_F6171_ & new_F6170_;
  assign new_F6162_ = new_F6171_ & new_F6172_;
  assign new_F6163_ = new_F6164_ | new_F6173_;
  assign new_F6164_ = F6153 | new_F6176_;
  assign new_F6165_ = new_F6175_ | new_F6174_;
  assign new_F6166_ = new_F6180_ & new_F6179_;
  assign new_F6167_ = new_F6178_ & new_F6177_;
  assign new_F6168_ = new_F6183_ | new_F6182_;
  assign new_F6169_ = new_F6178_ & new_F6181_;
  assign new_F6170_ = F6153 | new_F6186_;
  assign new_F6171_ = new_F6185_ | new_F6184_;
  assign new_F6172_ = new_F6188_ | new_F6187_;
  assign new_F6173_ = ~new_F6164_ & new_F6190_;
  assign new_F6174_ = ~new_F6166_ & new_F6178_;
  assign new_F6175_ = new_F6166_ & ~new_F6178_;
  assign new_F6176_ = F6152 & ~F6153;
  assign new_F6177_ = ~new_F6199_ | ~new_F6200_;
  assign new_F6178_ = new_F6192_ | new_F6194_;
  assign new_F6179_ = new_F6202_ | new_F6201_;
  assign new_F6180_ = new_F6196_ | new_F6195_;
  assign new_F6181_ = ~new_F6204_ | ~new_F6203_;
  assign new_F6182_ = ~new_F6205_ & new_F6206_;
  assign new_F6183_ = new_F6205_ & ~new_F6206_;
  assign new_F6184_ = ~F6152 & F6153;
  assign new_F6185_ = F6152 & ~F6153;
  assign new_F6186_ = ~new_F6168_ | new_F6178_;
  assign new_F6187_ = new_F6168_ & new_F6178_;
  assign new_F6188_ = ~new_F6168_ & ~new_F6178_;
  assign new_F6189_ = new_F6210_ | new_F6209_;
  assign new_F6190_ = F6156 | new_F6189_;
  assign new_F6191_ = new_F6214_ | new_F6213_;
  assign new_F6192_ = ~F6156 & new_F6191_;
  assign new_F6193_ = new_F6212_ | new_F6211_;
  assign new_F6194_ = F6156 & new_F6193_;
  assign new_F6195_ = F6154 & ~new_F6164_;
  assign new_F6196_ = ~F6154 & new_F6164_;
  assign new_F6197_ = ~F6153 | ~new_F6178_;
  assign new_F6198_ = new_F6164_ & new_F6197_;
  assign new_F6199_ = ~new_F6164_ & ~new_F6198_;
  assign new_F6200_ = new_F6164_ | new_F6197_;
  assign new_F6201_ = ~F6154 & F6155;
  assign new_F6202_ = F6154 & ~F6155;
  assign new_F6203_ = new_F6171_ | new_F6208_;
  assign new_F6204_ = ~new_F6171_ & ~new_F6207_;
  assign new_F6205_ = F6154 | new_F6171_;
  assign new_F6206_ = F6154 | F6155;
  assign new_F6207_ = new_F6171_ & new_F6208_;
  assign new_F6208_ = ~F6153 | ~new_F6178_;
  assign new_F6209_ = new_F6186_ & new_F6206_;
  assign new_F6210_ = ~new_F6186_ & ~new_F6206_;
  assign new_F6211_ = new_F6215_ | new_F6216_;
  assign new_F6212_ = ~F6157 & new_F6171_;
  assign new_F6213_ = new_F6217_ | new_F6218_;
  assign new_F6214_ = F6157 & new_F6171_;
  assign new_F6215_ = ~F6157 & ~new_F6171_;
  assign new_F6216_ = F6157 & ~new_F6171_;
  assign new_F6217_ = F6157 & ~new_F6171_;
  assign new_F6218_ = ~F6157 & new_F6171_;
  assign new_F6225_ = new_F6232_ & new_F6231_;
  assign new_F6226_ = new_F6234_ | new_F6233_;
  assign new_F6227_ = new_F6236_ | new_F6235_;
  assign new_F6228_ = new_F6238_ & new_F6237_;
  assign new_F6229_ = new_F6238_ & new_F6239_;
  assign new_F6230_ = new_F6231_ | new_F6240_;
  assign new_F6231_ = F6220 | new_F6243_;
  assign new_F6232_ = new_F6242_ | new_F6241_;
  assign new_F6233_ = new_F6247_ & new_F6246_;
  assign new_F6234_ = new_F6245_ & new_F6244_;
  assign new_F6235_ = new_F6250_ | new_F6249_;
  assign new_F6236_ = new_F6245_ & new_F6248_;
  assign new_F6237_ = F6220 | new_F6253_;
  assign new_F6238_ = new_F6252_ | new_F6251_;
  assign new_F6239_ = new_F6255_ | new_F6254_;
  assign new_F6240_ = ~new_F6231_ & new_F6257_;
  assign new_F6241_ = ~new_F6233_ & new_F6245_;
  assign new_F6242_ = new_F6233_ & ~new_F6245_;
  assign new_F6243_ = F6219 & ~F6220;
  assign new_F6244_ = ~new_F6266_ | ~new_F6267_;
  assign new_F6245_ = new_F6259_ | new_F6261_;
  assign new_F6246_ = new_F6269_ | new_F6268_;
  assign new_F6247_ = new_F6263_ | new_F6262_;
  assign new_F6248_ = ~new_F6271_ | ~new_F6270_;
  assign new_F6249_ = ~new_F6272_ & new_F6273_;
  assign new_F6250_ = new_F6272_ & ~new_F6273_;
  assign new_F6251_ = ~F6219 & F6220;
  assign new_F6252_ = F6219 & ~F6220;
  assign new_F6253_ = ~new_F6235_ | new_F6245_;
  assign new_F6254_ = new_F6235_ & new_F6245_;
  assign new_F6255_ = ~new_F6235_ & ~new_F6245_;
  assign new_F6256_ = new_F6277_ | new_F6276_;
  assign new_F6257_ = F6223 | new_F6256_;
  assign new_F6258_ = new_F6281_ | new_F6280_;
  assign new_F6259_ = ~F6223 & new_F6258_;
  assign new_F6260_ = new_F6279_ | new_F6278_;
  assign new_F6261_ = F6223 & new_F6260_;
  assign new_F6262_ = F6221 & ~new_F6231_;
  assign new_F6263_ = ~F6221 & new_F6231_;
  assign new_F6264_ = ~F6220 | ~new_F6245_;
  assign new_F6265_ = new_F6231_ & new_F6264_;
  assign new_F6266_ = ~new_F6231_ & ~new_F6265_;
  assign new_F6267_ = new_F6231_ | new_F6264_;
  assign new_F6268_ = ~F6221 & F6222;
  assign new_F6269_ = F6221 & ~F6222;
  assign new_F6270_ = new_F6238_ | new_F6275_;
  assign new_F6271_ = ~new_F6238_ & ~new_F6274_;
  assign new_F6272_ = F6221 | new_F6238_;
  assign new_F6273_ = F6221 | F6222;
  assign new_F6274_ = new_F6238_ & new_F6275_;
  assign new_F6275_ = ~F6220 | ~new_F6245_;
  assign new_F6276_ = new_F6253_ & new_F6273_;
  assign new_F6277_ = ~new_F6253_ & ~new_F6273_;
  assign new_F6278_ = new_F6282_ | new_F6283_;
  assign new_F6279_ = ~F6224 & new_F6238_;
  assign new_F6280_ = new_F6284_ | new_F6285_;
  assign new_F6281_ = F6224 & new_F6238_;
  assign new_F6282_ = ~F6224 & ~new_F6238_;
  assign new_F6283_ = F6224 & ~new_F6238_;
  assign new_F6284_ = F6224 & ~new_F6238_;
  assign new_F6285_ = ~F6224 & new_F6238_;
  assign new_F6292_ = new_F6299_ & new_F6298_;
  assign new_F6293_ = new_F6301_ | new_F6300_;
  assign new_F6294_ = new_F6303_ | new_F6302_;
  assign new_F6295_ = new_F6305_ & new_F6304_;
  assign new_F6296_ = new_F6305_ & new_F6306_;
  assign new_F6297_ = new_F6298_ | new_F6307_;
  assign new_F6298_ = F6287 | new_F6310_;
  assign new_F6299_ = new_F6309_ | new_F6308_;
  assign new_F6300_ = new_F6314_ & new_F6313_;
  assign new_F6301_ = new_F6312_ & new_F6311_;
  assign new_F6302_ = new_F6317_ | new_F6316_;
  assign new_F6303_ = new_F6312_ & new_F6315_;
  assign new_F6304_ = F6287 | new_F6320_;
  assign new_F6305_ = new_F6319_ | new_F6318_;
  assign new_F6306_ = new_F6322_ | new_F6321_;
  assign new_F6307_ = ~new_F6298_ & new_F6324_;
  assign new_F6308_ = ~new_F6300_ & new_F6312_;
  assign new_F6309_ = new_F6300_ & ~new_F6312_;
  assign new_F6310_ = F6286 & ~F6287;
  assign new_F6311_ = ~new_F6333_ | ~new_F6334_;
  assign new_F6312_ = new_F6326_ | new_F6328_;
  assign new_F6313_ = new_F6336_ | new_F6335_;
  assign new_F6314_ = new_F6330_ | new_F6329_;
  assign new_F6315_ = ~new_F6338_ | ~new_F6337_;
  assign new_F6316_ = ~new_F6339_ & new_F6340_;
  assign new_F6317_ = new_F6339_ & ~new_F6340_;
  assign new_F6318_ = ~F6286 & F6287;
  assign new_F6319_ = F6286 & ~F6287;
  assign new_F6320_ = ~new_F6302_ | new_F6312_;
  assign new_F6321_ = new_F6302_ & new_F6312_;
  assign new_F6322_ = ~new_F6302_ & ~new_F6312_;
  assign new_F6323_ = new_F6344_ | new_F6343_;
  assign new_F6324_ = F6290 | new_F6323_;
  assign new_F6325_ = new_F6348_ | new_F6347_;
  assign new_F6326_ = ~F6290 & new_F6325_;
  assign new_F6327_ = new_F6346_ | new_F6345_;
  assign new_F6328_ = F6290 & new_F6327_;
  assign new_F6329_ = F6288 & ~new_F6298_;
  assign new_F6330_ = ~F6288 & new_F6298_;
  assign new_F6331_ = ~F6287 | ~new_F6312_;
  assign new_F6332_ = new_F6298_ & new_F6331_;
  assign new_F6333_ = ~new_F6298_ & ~new_F6332_;
  assign new_F6334_ = new_F6298_ | new_F6331_;
  assign new_F6335_ = ~F6288 & F6289;
  assign new_F6336_ = F6288 & ~F6289;
  assign new_F6337_ = new_F6305_ | new_F6342_;
  assign new_F6338_ = ~new_F6305_ & ~new_F6341_;
  assign new_F6339_ = F6288 | new_F6305_;
  assign new_F6340_ = F6288 | F6289;
  assign new_F6341_ = new_F6305_ & new_F6342_;
  assign new_F6342_ = ~F6287 | ~new_F6312_;
  assign new_F6343_ = new_F6320_ & new_F6340_;
  assign new_F6344_ = ~new_F6320_ & ~new_F6340_;
  assign new_F6345_ = new_F6349_ | new_F6350_;
  assign new_F6346_ = ~F6291 & new_F6305_;
  assign new_F6347_ = new_F6351_ | new_F6352_;
  assign new_F6348_ = F6291 & new_F6305_;
  assign new_F6349_ = ~F6291 & ~new_F6305_;
  assign new_F6350_ = F6291 & ~new_F6305_;
  assign new_F6351_ = F6291 & ~new_F6305_;
  assign new_F6352_ = ~F6291 & new_F6305_;
  assign new_F6359_ = new_F6366_ & new_F6365_;
  assign new_F6360_ = new_F6368_ | new_F6367_;
  assign new_F6361_ = new_F6370_ | new_F6369_;
  assign new_F6362_ = new_F6372_ & new_F6371_;
  assign new_F6363_ = new_F6372_ & new_F6373_;
  assign new_F6364_ = new_F6365_ | new_F6374_;
  assign new_F6365_ = F6354 | new_F6377_;
  assign new_F6366_ = new_F6376_ | new_F6375_;
  assign new_F6367_ = new_F6381_ & new_F6380_;
  assign new_F6368_ = new_F6379_ & new_F6378_;
  assign new_F6369_ = new_F6384_ | new_F6383_;
  assign new_F6370_ = new_F6379_ & new_F6382_;
  assign new_F6371_ = F6354 | new_F6387_;
  assign new_F6372_ = new_F6386_ | new_F6385_;
  assign new_F6373_ = new_F6389_ | new_F6388_;
  assign new_F6374_ = ~new_F6365_ & new_F6391_;
  assign new_F6375_ = ~new_F6367_ & new_F6379_;
  assign new_F6376_ = new_F6367_ & ~new_F6379_;
  assign new_F6377_ = F6353 & ~F6354;
  assign new_F6378_ = ~new_F6400_ | ~new_F6401_;
  assign new_F6379_ = new_F6393_ | new_F6395_;
  assign new_F6380_ = new_F6403_ | new_F6402_;
  assign new_F6381_ = new_F6397_ | new_F6396_;
  assign new_F6382_ = ~new_F6405_ | ~new_F6404_;
  assign new_F6383_ = ~new_F6406_ & new_F6407_;
  assign new_F6384_ = new_F6406_ & ~new_F6407_;
  assign new_F6385_ = ~F6353 & F6354;
  assign new_F6386_ = F6353 & ~F6354;
  assign new_F6387_ = ~new_F6369_ | new_F6379_;
  assign new_F6388_ = new_F6369_ & new_F6379_;
  assign new_F6389_ = ~new_F6369_ & ~new_F6379_;
  assign new_F6390_ = new_F6411_ | new_F6410_;
  assign new_F6391_ = F6357 | new_F6390_;
  assign new_F6392_ = new_F6415_ | new_F6414_;
  assign new_F6393_ = ~F6357 & new_F6392_;
  assign new_F6394_ = new_F6413_ | new_F6412_;
  assign new_F6395_ = F6357 & new_F6394_;
  assign new_F6396_ = F6355 & ~new_F6365_;
  assign new_F6397_ = ~F6355 & new_F6365_;
  assign new_F6398_ = ~F6354 | ~new_F6379_;
  assign new_F6399_ = new_F6365_ & new_F6398_;
  assign new_F6400_ = ~new_F6365_ & ~new_F6399_;
  assign new_F6401_ = new_F6365_ | new_F6398_;
  assign new_F6402_ = ~F6355 & F6356;
  assign new_F6403_ = F6355 & ~F6356;
  assign new_F6404_ = new_F6372_ | new_F6409_;
  assign new_F6405_ = ~new_F6372_ & ~new_F6408_;
  assign new_F6406_ = F6355 | new_F6372_;
  assign new_F6407_ = F6355 | F6356;
  assign new_F6408_ = new_F6372_ & new_F6409_;
  assign new_F6409_ = ~F6354 | ~new_F6379_;
  assign new_F6410_ = new_F6387_ & new_F6407_;
  assign new_F6411_ = ~new_F6387_ & ~new_F6407_;
  assign new_F6412_ = new_F6416_ | new_F6417_;
  assign new_F6413_ = ~F6358 & new_F6372_;
  assign new_F6414_ = new_F6418_ | new_F6419_;
  assign new_F6415_ = F6358 & new_F6372_;
  assign new_F6416_ = ~F6358 & ~new_F6372_;
  assign new_F6417_ = F6358 & ~new_F6372_;
  assign new_F6418_ = F6358 & ~new_F6372_;
  assign new_F6419_ = ~F6358 & new_F6372_;
  assign new_F6426_ = new_F6433_ & new_F6432_;
  assign new_F6427_ = new_F6435_ | new_F6434_;
  assign new_F6428_ = new_F6437_ | new_F6436_;
  assign new_F6429_ = new_F6439_ & new_F6438_;
  assign new_F6430_ = new_F6439_ & new_F6440_;
  assign new_F6431_ = new_F6432_ | new_F6441_;
  assign new_F6432_ = F6421 | new_F6444_;
  assign new_F6433_ = new_F6443_ | new_F6442_;
  assign new_F6434_ = new_F6448_ & new_F6447_;
  assign new_F6435_ = new_F6446_ & new_F6445_;
  assign new_F6436_ = new_F6451_ | new_F6450_;
  assign new_F6437_ = new_F6446_ & new_F6449_;
  assign new_F6438_ = F6421 | new_F6454_;
  assign new_F6439_ = new_F6453_ | new_F6452_;
  assign new_F6440_ = new_F6456_ | new_F6455_;
  assign new_F6441_ = ~new_F6432_ & new_F6458_;
  assign new_F6442_ = ~new_F6434_ & new_F6446_;
  assign new_F6443_ = new_F6434_ & ~new_F6446_;
  assign new_F6444_ = F6420 & ~F6421;
  assign new_F6445_ = ~new_F6467_ | ~new_F6468_;
  assign new_F6446_ = new_F6460_ | new_F6462_;
  assign new_F6447_ = new_F6470_ | new_F6469_;
  assign new_F6448_ = new_F6464_ | new_F6463_;
  assign new_F6449_ = ~new_F6472_ | ~new_F6471_;
  assign new_F6450_ = ~new_F6473_ & new_F6474_;
  assign new_F6451_ = new_F6473_ & ~new_F6474_;
  assign new_F6452_ = ~F6420 & F6421;
  assign new_F6453_ = F6420 & ~F6421;
  assign new_F6454_ = ~new_F6436_ | new_F6446_;
  assign new_F6455_ = new_F6436_ & new_F6446_;
  assign new_F6456_ = ~new_F6436_ & ~new_F6446_;
  assign new_F6457_ = new_F6478_ | new_F6477_;
  assign new_F6458_ = F6424 | new_F6457_;
  assign new_F6459_ = new_F6482_ | new_F6481_;
  assign new_F6460_ = ~F6424 & new_F6459_;
  assign new_F6461_ = new_F6480_ | new_F6479_;
  assign new_F6462_ = F6424 & new_F6461_;
  assign new_F6463_ = F6422 & ~new_F6432_;
  assign new_F6464_ = ~F6422 & new_F6432_;
  assign new_F6465_ = ~F6421 | ~new_F6446_;
  assign new_F6466_ = new_F6432_ & new_F6465_;
  assign new_F6467_ = ~new_F6432_ & ~new_F6466_;
  assign new_F6468_ = new_F6432_ | new_F6465_;
  assign new_F6469_ = ~F6422 & F6423;
  assign new_F6470_ = F6422 & ~F6423;
  assign new_F6471_ = new_F6439_ | new_F6476_;
  assign new_F6472_ = ~new_F6439_ & ~new_F6475_;
  assign new_F6473_ = F6422 | new_F6439_;
  assign new_F6474_ = F6422 | F6423;
  assign new_F6475_ = new_F6439_ & new_F6476_;
  assign new_F6476_ = ~F6421 | ~new_F6446_;
  assign new_F6477_ = new_F6454_ & new_F6474_;
  assign new_F6478_ = ~new_F6454_ & ~new_F6474_;
  assign new_F6479_ = new_F6483_ | new_F6484_;
  assign new_F6480_ = ~F6425 & new_F6439_;
  assign new_F6481_ = new_F6485_ | new_F6486_;
  assign new_F6482_ = F6425 & new_F6439_;
  assign new_F6483_ = ~F6425 & ~new_F6439_;
  assign new_F6484_ = F6425 & ~new_F6439_;
  assign new_F6485_ = F6425 & ~new_F6439_;
  assign new_F6486_ = ~F6425 & new_F6439_;
  assign new_F6493_ = new_F6500_ & new_F6499_;
  assign new_F6494_ = new_F6502_ | new_F6501_;
  assign new_F6495_ = new_F6504_ | new_F6503_;
  assign new_F6496_ = new_F6506_ & new_F6505_;
  assign new_F6497_ = new_F6506_ & new_F6507_;
  assign new_F6498_ = new_F6499_ | new_F6508_;
  assign new_F6499_ = F6488 | new_F6511_;
  assign new_F6500_ = new_F6510_ | new_F6509_;
  assign new_F6501_ = new_F6515_ & new_F6514_;
  assign new_F6502_ = new_F6513_ & new_F6512_;
  assign new_F6503_ = new_F6518_ | new_F6517_;
  assign new_F6504_ = new_F6513_ & new_F6516_;
  assign new_F6505_ = F6488 | new_F6521_;
  assign new_F6506_ = new_F6520_ | new_F6519_;
  assign new_F6507_ = new_F6523_ | new_F6522_;
  assign new_F6508_ = ~new_F6499_ & new_F6525_;
  assign new_F6509_ = ~new_F6501_ & new_F6513_;
  assign new_F6510_ = new_F6501_ & ~new_F6513_;
  assign new_F6511_ = F6487 & ~F6488;
  assign new_F6512_ = ~new_F6534_ | ~new_F6535_;
  assign new_F6513_ = new_F6527_ | new_F6529_;
  assign new_F6514_ = new_F6537_ | new_F6536_;
  assign new_F6515_ = new_F6531_ | new_F6530_;
  assign new_F6516_ = ~new_F6539_ | ~new_F6538_;
  assign new_F6517_ = ~new_F6540_ & new_F6541_;
  assign new_F6518_ = new_F6540_ & ~new_F6541_;
  assign new_F6519_ = ~F6487 & F6488;
  assign new_F6520_ = F6487 & ~F6488;
  assign new_F6521_ = ~new_F6503_ | new_F6513_;
  assign new_F6522_ = new_F6503_ & new_F6513_;
  assign new_F6523_ = ~new_F6503_ & ~new_F6513_;
  assign new_F6524_ = new_F6545_ | new_F6544_;
  assign new_F6525_ = F6491 | new_F6524_;
  assign new_F6526_ = new_F6549_ | new_F6548_;
  assign new_F6527_ = ~F6491 & new_F6526_;
  assign new_F6528_ = new_F6547_ | new_F6546_;
  assign new_F6529_ = F6491 & new_F6528_;
  assign new_F6530_ = F6489 & ~new_F6499_;
  assign new_F6531_ = ~F6489 & new_F6499_;
  assign new_F6532_ = ~F6488 | ~new_F6513_;
  assign new_F6533_ = new_F6499_ & new_F6532_;
  assign new_F6534_ = ~new_F6499_ & ~new_F6533_;
  assign new_F6535_ = new_F6499_ | new_F6532_;
  assign new_F6536_ = ~F6489 & F6490;
  assign new_F6537_ = F6489 & ~F6490;
  assign new_F6538_ = new_F6506_ | new_F6543_;
  assign new_F6539_ = ~new_F6506_ & ~new_F6542_;
  assign new_F6540_ = F6489 | new_F6506_;
  assign new_F6541_ = F6489 | F6490;
  assign new_F6542_ = new_F6506_ & new_F6543_;
  assign new_F6543_ = ~F6488 | ~new_F6513_;
  assign new_F6544_ = new_F6521_ & new_F6541_;
  assign new_F6545_ = ~new_F6521_ & ~new_F6541_;
  assign new_F6546_ = new_F6550_ | new_F6551_;
  assign new_F6547_ = ~F6492 & new_F6506_;
  assign new_F6548_ = new_F6552_ | new_F6553_;
  assign new_F6549_ = F6492 & new_F6506_;
  assign new_F6550_ = ~F6492 & ~new_F6506_;
  assign new_F6551_ = F6492 & ~new_F6506_;
  assign new_F6552_ = F6492 & ~new_F6506_;
  assign new_F6553_ = ~F6492 & new_F6506_;
  assign new_F6560_ = new_F6567_ & new_F6566_;
  assign new_F6561_ = new_F6569_ | new_F6568_;
  assign new_F6562_ = new_F6571_ | new_F6570_;
  assign new_F6563_ = new_F6573_ & new_F6572_;
  assign new_F6564_ = new_F6573_ & new_F6574_;
  assign new_F6565_ = new_F6566_ | new_F6575_;
  assign new_F6566_ = F6555 | new_F6578_;
  assign new_F6567_ = new_F6577_ | new_F6576_;
  assign new_F6568_ = new_F6582_ & new_F6581_;
  assign new_F6569_ = new_F6580_ & new_F6579_;
  assign new_F6570_ = new_F6585_ | new_F6584_;
  assign new_F6571_ = new_F6580_ & new_F6583_;
  assign new_F6572_ = F6555 | new_F6588_;
  assign new_F6573_ = new_F6587_ | new_F6586_;
  assign new_F6574_ = new_F6590_ | new_F6589_;
  assign new_F6575_ = ~new_F6566_ & new_F6592_;
  assign new_F6576_ = ~new_F6568_ & new_F6580_;
  assign new_F6577_ = new_F6568_ & ~new_F6580_;
  assign new_F6578_ = F6554 & ~F6555;
  assign new_F6579_ = ~new_F6601_ | ~new_F6602_;
  assign new_F6580_ = new_F6594_ | new_F6596_;
  assign new_F6581_ = new_F6604_ | new_F6603_;
  assign new_F6582_ = new_F6598_ | new_F6597_;
  assign new_F6583_ = ~new_F6606_ | ~new_F6605_;
  assign new_F6584_ = ~new_F6607_ & new_F6608_;
  assign new_F6585_ = new_F6607_ & ~new_F6608_;
  assign new_F6586_ = ~F6554 & F6555;
  assign new_F6587_ = F6554 & ~F6555;
  assign new_F6588_ = ~new_F6570_ | new_F6580_;
  assign new_F6589_ = new_F6570_ & new_F6580_;
  assign new_F6590_ = ~new_F6570_ & ~new_F6580_;
  assign new_F6591_ = new_F6612_ | new_F6611_;
  assign new_F6592_ = F6558 | new_F6591_;
  assign new_F6593_ = new_F6616_ | new_F6615_;
  assign new_F6594_ = ~F6558 & new_F6593_;
  assign new_F6595_ = new_F6614_ | new_F6613_;
  assign new_F6596_ = F6558 & new_F6595_;
  assign new_F6597_ = F6556 & ~new_F6566_;
  assign new_F6598_ = ~F6556 & new_F6566_;
  assign new_F6599_ = ~F6555 | ~new_F6580_;
  assign new_F6600_ = new_F6566_ & new_F6599_;
  assign new_F6601_ = ~new_F6566_ & ~new_F6600_;
  assign new_F6602_ = new_F6566_ | new_F6599_;
  assign new_F6603_ = ~F6556 & F6557;
  assign new_F6604_ = F6556 & ~F6557;
  assign new_F6605_ = new_F6573_ | new_F6610_;
  assign new_F6606_ = ~new_F6573_ & ~new_F6609_;
  assign new_F6607_ = F6556 | new_F6573_;
  assign new_F6608_ = F6556 | F6557;
  assign new_F6609_ = new_F6573_ & new_F6610_;
  assign new_F6610_ = ~F6555 | ~new_F6580_;
  assign new_F6611_ = new_F6588_ & new_F6608_;
  assign new_F6612_ = ~new_F6588_ & ~new_F6608_;
  assign new_F6613_ = new_F6617_ | new_F6618_;
  assign new_F6614_ = ~F6559 & new_F6573_;
  assign new_F6615_ = new_F6619_ | new_F6620_;
  assign new_F6616_ = F6559 & new_F6573_;
  assign new_F6617_ = ~F6559 & ~new_F6573_;
  assign new_F6618_ = F6559 & ~new_F6573_;
  assign new_F6619_ = F6559 & ~new_F6573_;
  assign new_F6620_ = ~F6559 & new_F6573_;
  assign new_F6627_ = new_F6634_ & new_F6633_;
  assign new_F6628_ = new_F6636_ | new_F6635_;
  assign new_F6629_ = new_F6638_ | new_F6637_;
  assign new_F6630_ = new_F6640_ & new_F6639_;
  assign new_F6631_ = new_F6640_ & new_F6641_;
  assign new_F6632_ = new_F6633_ | new_F6642_;
  assign new_F6633_ = F6622 | new_F6645_;
  assign new_F6634_ = new_F6644_ | new_F6643_;
  assign new_F6635_ = new_F6649_ & new_F6648_;
  assign new_F6636_ = new_F6647_ & new_F6646_;
  assign new_F6637_ = new_F6652_ | new_F6651_;
  assign new_F6638_ = new_F6647_ & new_F6650_;
  assign new_F6639_ = F6622 | new_F6655_;
  assign new_F6640_ = new_F6654_ | new_F6653_;
  assign new_F6641_ = new_F6657_ | new_F6656_;
  assign new_F6642_ = ~new_F6633_ & new_F6659_;
  assign new_F6643_ = ~new_F6635_ & new_F6647_;
  assign new_F6644_ = new_F6635_ & ~new_F6647_;
  assign new_F6645_ = F6621 & ~F6622;
  assign new_F6646_ = ~new_F6668_ | ~new_F6669_;
  assign new_F6647_ = new_F6661_ | new_F6663_;
  assign new_F6648_ = new_F6671_ | new_F6670_;
  assign new_F6649_ = new_F6665_ | new_F6664_;
  assign new_F6650_ = ~new_F6673_ | ~new_F6672_;
  assign new_F6651_ = ~new_F6674_ & new_F6675_;
  assign new_F6652_ = new_F6674_ & ~new_F6675_;
  assign new_F6653_ = ~F6621 & F6622;
  assign new_F6654_ = F6621 & ~F6622;
  assign new_F6655_ = ~new_F6637_ | new_F6647_;
  assign new_F6656_ = new_F6637_ & new_F6647_;
  assign new_F6657_ = ~new_F6637_ & ~new_F6647_;
  assign new_F6658_ = new_F6679_ | new_F6678_;
  assign new_F6659_ = F6625 | new_F6658_;
  assign new_F6660_ = new_F6683_ | new_F6682_;
  assign new_F6661_ = ~F6625 & new_F6660_;
  assign new_F6662_ = new_F6681_ | new_F6680_;
  assign new_F6663_ = F6625 & new_F6662_;
  assign new_F6664_ = F6623 & ~new_F6633_;
  assign new_F6665_ = ~F6623 & new_F6633_;
  assign new_F6666_ = ~F6622 | ~new_F6647_;
  assign new_F6667_ = new_F6633_ & new_F6666_;
  assign new_F6668_ = ~new_F6633_ & ~new_F6667_;
  assign new_F6669_ = new_F6633_ | new_F6666_;
  assign new_F6670_ = ~F6623 & F6624;
  assign new_F6671_ = F6623 & ~F6624;
  assign new_F6672_ = new_F6640_ | new_F6677_;
  assign new_F6673_ = ~new_F6640_ & ~new_F6676_;
  assign new_F6674_ = F6623 | new_F6640_;
  assign new_F6675_ = F6623 | F6624;
  assign new_F6676_ = new_F6640_ & new_F6677_;
  assign new_F6677_ = ~F6622 | ~new_F6647_;
  assign new_F6678_ = new_F6655_ & new_F6675_;
  assign new_F6679_ = ~new_F6655_ & ~new_F6675_;
  assign new_F6680_ = new_F6684_ | new_F6685_;
  assign new_F6681_ = ~F6626 & new_F6640_;
  assign new_F6682_ = new_F6686_ | new_F6687_;
  assign new_F6683_ = F6626 & new_F6640_;
  assign new_F6684_ = ~F6626 & ~new_F6640_;
  assign new_F6685_ = F6626 & ~new_F6640_;
  assign new_F6686_ = F6626 & ~new_F6640_;
  assign new_F6687_ = ~F6626 & new_F6640_;
  assign new_F6694_ = new_F6701_ & new_F6700_;
  assign new_F6695_ = new_F6703_ | new_F6702_;
  assign new_F6696_ = new_F6705_ | new_F6704_;
  assign new_F6697_ = new_F6707_ & new_F6706_;
  assign new_F6698_ = new_F6707_ & new_F6708_;
  assign new_F6699_ = new_F6700_ | new_F6709_;
  assign new_F6700_ = F6689 | new_F6712_;
  assign new_F6701_ = new_F6711_ | new_F6710_;
  assign new_F6702_ = new_F6716_ & new_F6715_;
  assign new_F6703_ = new_F6714_ & new_F6713_;
  assign new_F6704_ = new_F6719_ | new_F6718_;
  assign new_F6705_ = new_F6714_ & new_F6717_;
  assign new_F6706_ = F6689 | new_F6722_;
  assign new_F6707_ = new_F6721_ | new_F6720_;
  assign new_F6708_ = new_F6724_ | new_F6723_;
  assign new_F6709_ = ~new_F6700_ & new_F6726_;
  assign new_F6710_ = ~new_F6702_ & new_F6714_;
  assign new_F6711_ = new_F6702_ & ~new_F6714_;
  assign new_F6712_ = F6688 & ~F6689;
  assign new_F6713_ = ~new_F6735_ | ~new_F6736_;
  assign new_F6714_ = new_F6728_ | new_F6730_;
  assign new_F6715_ = new_F6738_ | new_F6737_;
  assign new_F6716_ = new_F6732_ | new_F6731_;
  assign new_F6717_ = ~new_F6740_ | ~new_F6739_;
  assign new_F6718_ = ~new_F6741_ & new_F6742_;
  assign new_F6719_ = new_F6741_ & ~new_F6742_;
  assign new_F6720_ = ~F6688 & F6689;
  assign new_F6721_ = F6688 & ~F6689;
  assign new_F6722_ = ~new_F6704_ | new_F6714_;
  assign new_F6723_ = new_F6704_ & new_F6714_;
  assign new_F6724_ = ~new_F6704_ & ~new_F6714_;
  assign new_F6725_ = new_F6746_ | new_F6745_;
  assign new_F6726_ = F6692 | new_F6725_;
  assign new_F6727_ = new_F6750_ | new_F6749_;
  assign new_F6728_ = ~F6692 & new_F6727_;
  assign new_F6729_ = new_F6748_ | new_F6747_;
  assign new_F6730_ = F6692 & new_F6729_;
  assign new_F6731_ = F6690 & ~new_F6700_;
  assign new_F6732_ = ~F6690 & new_F6700_;
  assign new_F6733_ = ~F6689 | ~new_F6714_;
  assign new_F6734_ = new_F6700_ & new_F6733_;
  assign new_F6735_ = ~new_F6700_ & ~new_F6734_;
  assign new_F6736_ = new_F6700_ | new_F6733_;
  assign new_F6737_ = ~F6690 & F6691;
  assign new_F6738_ = F6690 & ~F6691;
  assign new_F6739_ = new_F6707_ | new_F6744_;
  assign new_F6740_ = ~new_F6707_ & ~new_F6743_;
  assign new_F6741_ = F6690 | new_F6707_;
  assign new_F6742_ = F6690 | F6691;
  assign new_F6743_ = new_F6707_ & new_F6744_;
  assign new_F6744_ = ~F6689 | ~new_F6714_;
  assign new_F6745_ = new_F6722_ & new_F6742_;
  assign new_F6746_ = ~new_F6722_ & ~new_F6742_;
  assign new_F6747_ = new_F6751_ | new_F6752_;
  assign new_F6748_ = ~F6693 & new_F6707_;
  assign new_F6749_ = new_F6753_ | new_F6754_;
  assign new_F6750_ = F6693 & new_F6707_;
  assign new_F6751_ = ~F6693 & ~new_F6707_;
  assign new_F6752_ = F6693 & ~new_F6707_;
  assign new_F6753_ = F6693 & ~new_F6707_;
  assign new_F6754_ = ~F6693 & new_F6707_;
  assign new_F6761_ = new_F6768_ & new_F6767_;
  assign new_F6762_ = new_F6770_ | new_F6769_;
  assign new_F6763_ = new_F6772_ | new_F6771_;
  assign new_F6764_ = new_F6774_ & new_F6773_;
  assign new_F6765_ = new_F6774_ & new_F6775_;
  assign new_F6766_ = new_F6767_ | new_F6776_;
  assign new_F6767_ = F6756 | new_F6779_;
  assign new_F6768_ = new_F6778_ | new_F6777_;
  assign new_F6769_ = new_F6783_ & new_F6782_;
  assign new_F6770_ = new_F6781_ & new_F6780_;
  assign new_F6771_ = new_F6786_ | new_F6785_;
  assign new_F6772_ = new_F6781_ & new_F6784_;
  assign new_F6773_ = F6756 | new_F6789_;
  assign new_F6774_ = new_F6788_ | new_F6787_;
  assign new_F6775_ = new_F6791_ | new_F6790_;
  assign new_F6776_ = ~new_F6767_ & new_F6793_;
  assign new_F6777_ = ~new_F6769_ & new_F6781_;
  assign new_F6778_ = new_F6769_ & ~new_F6781_;
  assign new_F6779_ = F6755 & ~F6756;
  assign new_F6780_ = ~new_F6802_ | ~new_F6803_;
  assign new_F6781_ = new_F6795_ | new_F6797_;
  assign new_F6782_ = new_F6805_ | new_F6804_;
  assign new_F6783_ = new_F6799_ | new_F6798_;
  assign new_F6784_ = ~new_F6807_ | ~new_F6806_;
  assign new_F6785_ = ~new_F6808_ & new_F6809_;
  assign new_F6786_ = new_F6808_ & ~new_F6809_;
  assign new_F6787_ = ~F6755 & F6756;
  assign new_F6788_ = F6755 & ~F6756;
  assign new_F6789_ = ~new_F6771_ | new_F6781_;
  assign new_F6790_ = new_F6771_ & new_F6781_;
  assign new_F6791_ = ~new_F6771_ & ~new_F6781_;
  assign new_F6792_ = new_F6813_ | new_F6812_;
  assign new_F6793_ = F6759 | new_F6792_;
  assign new_F6794_ = new_F6817_ | new_F6816_;
  assign new_F6795_ = ~F6759 & new_F6794_;
  assign new_F6796_ = new_F6815_ | new_F6814_;
  assign new_F6797_ = F6759 & new_F6796_;
  assign new_F6798_ = F6757 & ~new_F6767_;
  assign new_F6799_ = ~F6757 & new_F6767_;
  assign new_F6800_ = ~F6756 | ~new_F6781_;
  assign new_F6801_ = new_F6767_ & new_F6800_;
  assign new_F6802_ = ~new_F6767_ & ~new_F6801_;
  assign new_F6803_ = new_F6767_ | new_F6800_;
  assign new_F6804_ = ~F6757 & F6758;
  assign new_F6805_ = F6757 & ~F6758;
  assign new_F6806_ = new_F6774_ | new_F6811_;
  assign new_F6807_ = ~new_F6774_ & ~new_F6810_;
  assign new_F6808_ = F6757 | new_F6774_;
  assign new_F6809_ = F6757 | F6758;
  assign new_F6810_ = new_F6774_ & new_F6811_;
  assign new_F6811_ = ~F6756 | ~new_F6781_;
  assign new_F6812_ = new_F6789_ & new_F6809_;
  assign new_F6813_ = ~new_F6789_ & ~new_F6809_;
  assign new_F6814_ = new_F6818_ | new_F6819_;
  assign new_F6815_ = ~F6760 & new_F6774_;
  assign new_F6816_ = new_F6820_ | new_F6821_;
  assign new_F6817_ = F6760 & new_F6774_;
  assign new_F6818_ = ~F6760 & ~new_F6774_;
  assign new_F6819_ = F6760 & ~new_F6774_;
  assign new_F6820_ = F6760 & ~new_F6774_;
  assign new_F6821_ = ~F6760 & new_F6774_;
  assign new_F6828_ = new_F6835_ & new_F6834_;
  assign new_F6829_ = new_F6837_ | new_F6836_;
  assign new_F6830_ = new_F6839_ | new_F6838_;
  assign new_F6831_ = new_F6841_ & new_F6840_;
  assign new_F6832_ = new_F6841_ & new_F6842_;
  assign new_F6833_ = new_F6834_ | new_F6843_;
  assign new_F6834_ = F6823 | new_F6846_;
  assign new_F6835_ = new_F6845_ | new_F6844_;
  assign new_F6836_ = new_F6850_ & new_F6849_;
  assign new_F6837_ = new_F6848_ & new_F6847_;
  assign new_F6838_ = new_F6853_ | new_F6852_;
  assign new_F6839_ = new_F6848_ & new_F6851_;
  assign new_F6840_ = F6823 | new_F6856_;
  assign new_F6841_ = new_F6855_ | new_F6854_;
  assign new_F6842_ = new_F6858_ | new_F6857_;
  assign new_F6843_ = ~new_F6834_ & new_F6860_;
  assign new_F6844_ = ~new_F6836_ & new_F6848_;
  assign new_F6845_ = new_F6836_ & ~new_F6848_;
  assign new_F6846_ = F6822 & ~F6823;
  assign new_F6847_ = ~new_F6869_ | ~new_F6870_;
  assign new_F6848_ = new_F6862_ | new_F6864_;
  assign new_F6849_ = new_F6872_ | new_F6871_;
  assign new_F6850_ = new_F6866_ | new_F6865_;
  assign new_F6851_ = ~new_F6874_ | ~new_F6873_;
  assign new_F6852_ = ~new_F6875_ & new_F6876_;
  assign new_F6853_ = new_F6875_ & ~new_F6876_;
  assign new_F6854_ = ~F6822 & F6823;
  assign new_F6855_ = F6822 & ~F6823;
  assign new_F6856_ = ~new_F6838_ | new_F6848_;
  assign new_F6857_ = new_F6838_ & new_F6848_;
  assign new_F6858_ = ~new_F6838_ & ~new_F6848_;
  assign new_F6859_ = new_F6880_ | new_F6879_;
  assign new_F6860_ = F6826 | new_F6859_;
  assign new_F6861_ = new_F6884_ | new_F6883_;
  assign new_F6862_ = ~F6826 & new_F6861_;
  assign new_F6863_ = new_F6882_ | new_F6881_;
  assign new_F6864_ = F6826 & new_F6863_;
  assign new_F6865_ = F6824 & ~new_F6834_;
  assign new_F6866_ = ~F6824 & new_F6834_;
  assign new_F6867_ = ~F6823 | ~new_F6848_;
  assign new_F6868_ = new_F6834_ & new_F6867_;
  assign new_F6869_ = ~new_F6834_ & ~new_F6868_;
  assign new_F6870_ = new_F6834_ | new_F6867_;
  assign new_F6871_ = ~F6824 & F6825;
  assign new_F6872_ = F6824 & ~F6825;
  assign new_F6873_ = new_F6841_ | new_F6878_;
  assign new_F6874_ = ~new_F6841_ & ~new_F6877_;
  assign new_F6875_ = F6824 | new_F6841_;
  assign new_F6876_ = F6824 | F6825;
  assign new_F6877_ = new_F6841_ & new_F6878_;
  assign new_F6878_ = ~F6823 | ~new_F6848_;
  assign new_F6879_ = new_F6856_ & new_F6876_;
  assign new_F6880_ = ~new_F6856_ & ~new_F6876_;
  assign new_F6881_ = new_F6885_ | new_F6886_;
  assign new_F6882_ = ~F6827 & new_F6841_;
  assign new_F6883_ = new_F6887_ | new_F6888_;
  assign new_F6884_ = F6827 & new_F6841_;
  assign new_F6885_ = ~F6827 & ~new_F6841_;
  assign new_F6886_ = F6827 & ~new_F6841_;
  assign new_F6887_ = F6827 & ~new_F6841_;
  assign new_F6888_ = ~F6827 & new_F6841_;
  assign new_F6895_ = new_F6902_ & new_F6901_;
  assign new_F6896_ = new_F6904_ | new_F6903_;
  assign new_F6897_ = new_F6906_ | new_F6905_;
  assign new_F6898_ = new_F6908_ & new_F6907_;
  assign new_F6899_ = new_F6908_ & new_F6909_;
  assign new_F6900_ = new_F6901_ | new_F6910_;
  assign new_F6901_ = F6890 | new_F6913_;
  assign new_F6902_ = new_F6912_ | new_F6911_;
  assign new_F6903_ = new_F6917_ & new_F6916_;
  assign new_F6904_ = new_F6915_ & new_F6914_;
  assign new_F6905_ = new_F6920_ | new_F6919_;
  assign new_F6906_ = new_F6915_ & new_F6918_;
  assign new_F6907_ = F6890 | new_F6923_;
  assign new_F6908_ = new_F6922_ | new_F6921_;
  assign new_F6909_ = new_F6925_ | new_F6924_;
  assign new_F6910_ = ~new_F6901_ & new_F6927_;
  assign new_F6911_ = ~new_F6903_ & new_F6915_;
  assign new_F6912_ = new_F6903_ & ~new_F6915_;
  assign new_F6913_ = F6889 & ~F6890;
  assign new_F6914_ = ~new_F6936_ | ~new_F6937_;
  assign new_F6915_ = new_F6929_ | new_F6931_;
  assign new_F6916_ = new_F6939_ | new_F6938_;
  assign new_F6917_ = new_F6933_ | new_F6932_;
  assign new_F6918_ = ~new_F6941_ | ~new_F6940_;
  assign new_F6919_ = ~new_F6942_ & new_F6943_;
  assign new_F6920_ = new_F6942_ & ~new_F6943_;
  assign new_F6921_ = ~F6889 & F6890;
  assign new_F6922_ = F6889 & ~F6890;
  assign new_F6923_ = ~new_F6905_ | new_F6915_;
  assign new_F6924_ = new_F6905_ & new_F6915_;
  assign new_F6925_ = ~new_F6905_ & ~new_F6915_;
  assign new_F6926_ = new_F6947_ | new_F6946_;
  assign new_F6927_ = F6893 | new_F6926_;
  assign new_F6928_ = new_F6951_ | new_F6950_;
  assign new_F6929_ = ~F6893 & new_F6928_;
  assign new_F6930_ = new_F6949_ | new_F6948_;
  assign new_F6931_ = F6893 & new_F6930_;
  assign new_F6932_ = F6891 & ~new_F6901_;
  assign new_F6933_ = ~F6891 & new_F6901_;
  assign new_F6934_ = ~F6890 | ~new_F6915_;
  assign new_F6935_ = new_F6901_ & new_F6934_;
  assign new_F6936_ = ~new_F6901_ & ~new_F6935_;
  assign new_F6937_ = new_F6901_ | new_F6934_;
  assign new_F6938_ = ~F6891 & F6892;
  assign new_F6939_ = F6891 & ~F6892;
  assign new_F6940_ = new_F6908_ | new_F6945_;
  assign new_F6941_ = ~new_F6908_ & ~new_F6944_;
  assign new_F6942_ = F6891 | new_F6908_;
  assign new_F6943_ = F6891 | F6892;
  assign new_F6944_ = new_F6908_ & new_F6945_;
  assign new_F6945_ = ~F6890 | ~new_F6915_;
  assign new_F6946_ = new_F6923_ & new_F6943_;
  assign new_F6947_ = ~new_F6923_ & ~new_F6943_;
  assign new_F6948_ = new_F6952_ | new_F6953_;
  assign new_F6949_ = ~F6894 & new_F6908_;
  assign new_F6950_ = new_F6954_ | new_F6955_;
  assign new_F6951_ = F6894 & new_F6908_;
  assign new_F6952_ = ~F6894 & ~new_F6908_;
  assign new_F6953_ = F6894 & ~new_F6908_;
  assign new_F6954_ = F6894 & ~new_F6908_;
  assign new_F6955_ = ~F6894 & new_F6908_;
  assign new_F6962_ = new_F6969_ & new_F6968_;
  assign new_F6963_ = new_F6971_ | new_F6970_;
  assign new_F6964_ = new_F6973_ | new_F6972_;
  assign new_F6965_ = new_F6975_ & new_F6974_;
  assign new_F6966_ = new_F6975_ & new_F6976_;
  assign new_F6967_ = new_F6968_ | new_F6977_;
  assign new_F6968_ = F6957 | new_F6980_;
  assign new_F6969_ = new_F6979_ | new_F6978_;
  assign new_F6970_ = new_F6984_ & new_F6983_;
  assign new_F6971_ = new_F6982_ & new_F6981_;
  assign new_F6972_ = new_F6987_ | new_F6986_;
  assign new_F6973_ = new_F6982_ & new_F6985_;
  assign new_F6974_ = F6957 | new_F6990_;
  assign new_F6975_ = new_F6989_ | new_F6988_;
  assign new_F6976_ = new_F6992_ | new_F6991_;
  assign new_F6977_ = ~new_F6968_ & new_F6994_;
  assign new_F6978_ = ~new_F6970_ & new_F6982_;
  assign new_F6979_ = new_F6970_ & ~new_F6982_;
  assign new_F6980_ = F6956 & ~F6957;
  assign new_F6981_ = ~new_F7003_ | ~new_F7004_;
  assign new_F6982_ = new_F6996_ | new_F6998_;
  assign new_F6983_ = new_F7006_ | new_F7005_;
  assign new_F6984_ = new_F7000_ | new_F6999_;
  assign new_F6985_ = ~new_F7008_ | ~new_F7007_;
  assign new_F6986_ = ~new_F7009_ & new_F7010_;
  assign new_F6987_ = new_F7009_ & ~new_F7010_;
  assign new_F6988_ = ~F6956 & F6957;
  assign new_F6989_ = F6956 & ~F6957;
  assign new_F6990_ = ~new_F6972_ | new_F6982_;
  assign new_F6991_ = new_F6972_ & new_F6982_;
  assign new_F6992_ = ~new_F6972_ & ~new_F6982_;
  assign new_F6993_ = new_F7014_ | new_F7013_;
  assign new_F6994_ = F6960 | new_F6993_;
  assign new_F6995_ = new_F7018_ | new_F7017_;
  assign new_F6996_ = ~F6960 & new_F6995_;
  assign new_F6997_ = new_F7016_ | new_F7015_;
  assign new_F6998_ = F6960 & new_F6997_;
  assign new_F6999_ = F6958 & ~new_F6968_;
  assign new_F7000_ = ~F6958 & new_F6968_;
  assign new_F7001_ = ~F6957 | ~new_F6982_;
  assign new_F7002_ = new_F6968_ & new_F7001_;
  assign new_F7003_ = ~new_F6968_ & ~new_F7002_;
  assign new_F7004_ = new_F6968_ | new_F7001_;
  assign new_F7005_ = ~F6958 & F6959;
  assign new_F7006_ = F6958 & ~F6959;
  assign new_F7007_ = new_F6975_ | new_F7012_;
  assign new_F7008_ = ~new_F6975_ & ~new_F7011_;
  assign new_F7009_ = F6958 | new_F6975_;
  assign new_F7010_ = F6958 | F6959;
  assign new_F7011_ = new_F6975_ & new_F7012_;
  assign new_F7012_ = ~F6957 | ~new_F6982_;
  assign new_F7013_ = new_F6990_ & new_F7010_;
  assign new_F7014_ = ~new_F6990_ & ~new_F7010_;
  assign new_F7015_ = new_F7019_ | new_F7020_;
  assign new_F7016_ = ~F6961 & new_F6975_;
  assign new_F7017_ = new_F7021_ | new_F7022_;
  assign new_F7018_ = F6961 & new_F6975_;
  assign new_F7019_ = ~F6961 & ~new_F6975_;
  assign new_F7020_ = F6961 & ~new_F6975_;
  assign new_F7021_ = F6961 & ~new_F6975_;
  assign new_F7022_ = ~F6961 & new_F6975_;
  assign new_F7029_ = new_F7036_ & new_F7035_;
  assign new_F7030_ = new_F7038_ | new_F7037_;
  assign new_F7031_ = new_F7040_ | new_F7039_;
  assign new_F7032_ = new_F7042_ & new_F7041_;
  assign new_F7033_ = new_F7042_ & new_F7043_;
  assign new_F7034_ = new_F7035_ | new_F7044_;
  assign new_F7035_ = F7024 | new_F7047_;
  assign new_F7036_ = new_F7046_ | new_F7045_;
  assign new_F7037_ = new_F7051_ & new_F7050_;
  assign new_F7038_ = new_F7049_ & new_F7048_;
  assign new_F7039_ = new_F7054_ | new_F7053_;
  assign new_F7040_ = new_F7049_ & new_F7052_;
  assign new_F7041_ = F7024 | new_F7057_;
  assign new_F7042_ = new_F7056_ | new_F7055_;
  assign new_F7043_ = new_F7059_ | new_F7058_;
  assign new_F7044_ = ~new_F7035_ & new_F7061_;
  assign new_F7045_ = ~new_F7037_ & new_F7049_;
  assign new_F7046_ = new_F7037_ & ~new_F7049_;
  assign new_F7047_ = F7023 & ~F7024;
  assign new_F7048_ = ~new_F7070_ | ~new_F7071_;
  assign new_F7049_ = new_F7063_ | new_F7065_;
  assign new_F7050_ = new_F7073_ | new_F7072_;
  assign new_F7051_ = new_F7067_ | new_F7066_;
  assign new_F7052_ = ~new_F7075_ | ~new_F7074_;
  assign new_F7053_ = ~new_F7076_ & new_F7077_;
  assign new_F7054_ = new_F7076_ & ~new_F7077_;
  assign new_F7055_ = ~F7023 & F7024;
  assign new_F7056_ = F7023 & ~F7024;
  assign new_F7057_ = ~new_F7039_ | new_F7049_;
  assign new_F7058_ = new_F7039_ & new_F7049_;
  assign new_F7059_ = ~new_F7039_ & ~new_F7049_;
  assign new_F7060_ = new_F7081_ | new_F7080_;
  assign new_F7061_ = F7027 | new_F7060_;
  assign new_F7062_ = new_F7085_ | new_F7084_;
  assign new_F7063_ = ~F7027 & new_F7062_;
  assign new_F7064_ = new_F7083_ | new_F7082_;
  assign new_F7065_ = F7027 & new_F7064_;
  assign new_F7066_ = F7025 & ~new_F7035_;
  assign new_F7067_ = ~F7025 & new_F7035_;
  assign new_F7068_ = ~F7024 | ~new_F7049_;
  assign new_F7069_ = new_F7035_ & new_F7068_;
  assign new_F7070_ = ~new_F7035_ & ~new_F7069_;
  assign new_F7071_ = new_F7035_ | new_F7068_;
  assign new_F7072_ = ~F7025 & F7026;
  assign new_F7073_ = F7025 & ~F7026;
  assign new_F7074_ = new_F7042_ | new_F7079_;
  assign new_F7075_ = ~new_F7042_ & ~new_F7078_;
  assign new_F7076_ = F7025 | new_F7042_;
  assign new_F7077_ = F7025 | F7026;
  assign new_F7078_ = new_F7042_ & new_F7079_;
  assign new_F7079_ = ~F7024 | ~new_F7049_;
  assign new_F7080_ = new_F7057_ & new_F7077_;
  assign new_F7081_ = ~new_F7057_ & ~new_F7077_;
  assign new_F7082_ = new_F7086_ | new_F7087_;
  assign new_F7083_ = ~F7028 & new_F7042_;
  assign new_F7084_ = new_F7088_ | new_F7089_;
  assign new_F7085_ = F7028 & new_F7042_;
  assign new_F7086_ = ~F7028 & ~new_F7042_;
  assign new_F7087_ = F7028 & ~new_F7042_;
  assign new_F7088_ = F7028 & ~new_F7042_;
  assign new_F7089_ = ~F7028 & new_F7042_;
  assign new_F7096_ = new_F7103_ & new_F7102_;
  assign new_F7097_ = new_F7105_ | new_F7104_;
  assign new_F7098_ = new_F7107_ | new_F7106_;
  assign new_F7099_ = new_F7109_ & new_F7108_;
  assign new_F7100_ = new_F7109_ & new_F7110_;
  assign new_F7101_ = new_F7102_ | new_F7111_;
  assign new_F7102_ = F7091 | new_F7114_;
  assign new_F7103_ = new_F7113_ | new_F7112_;
  assign new_F7104_ = new_F7118_ & new_F7117_;
  assign new_F7105_ = new_F7116_ & new_F7115_;
  assign new_F7106_ = new_F7121_ | new_F7120_;
  assign new_F7107_ = new_F7116_ & new_F7119_;
  assign new_F7108_ = F7091 | new_F7124_;
  assign new_F7109_ = new_F7123_ | new_F7122_;
  assign new_F7110_ = new_F7126_ | new_F7125_;
  assign new_F7111_ = ~new_F7102_ & new_F7128_;
  assign new_F7112_ = ~new_F7104_ & new_F7116_;
  assign new_F7113_ = new_F7104_ & ~new_F7116_;
  assign new_F7114_ = F7090 & ~F7091;
  assign new_F7115_ = ~new_F7137_ | ~new_F7138_;
  assign new_F7116_ = new_F7130_ | new_F7132_;
  assign new_F7117_ = new_F7140_ | new_F7139_;
  assign new_F7118_ = new_F7134_ | new_F7133_;
  assign new_F7119_ = ~new_F7142_ | ~new_F7141_;
  assign new_F7120_ = ~new_F7143_ & new_F7144_;
  assign new_F7121_ = new_F7143_ & ~new_F7144_;
  assign new_F7122_ = ~F7090 & F7091;
  assign new_F7123_ = F7090 & ~F7091;
  assign new_F7124_ = ~new_F7106_ | new_F7116_;
  assign new_F7125_ = new_F7106_ & new_F7116_;
  assign new_F7126_ = ~new_F7106_ & ~new_F7116_;
  assign new_F7127_ = new_F7148_ | new_F7147_;
  assign new_F7128_ = F7094 | new_F7127_;
  assign new_F7129_ = new_F7152_ | new_F7151_;
  assign new_F7130_ = ~F7094 & new_F7129_;
  assign new_F7131_ = new_F7150_ | new_F7149_;
  assign new_F7132_ = F7094 & new_F7131_;
  assign new_F7133_ = F7092 & ~new_F7102_;
  assign new_F7134_ = ~F7092 & new_F7102_;
  assign new_F7135_ = ~F7091 | ~new_F7116_;
  assign new_F7136_ = new_F7102_ & new_F7135_;
  assign new_F7137_ = ~new_F7102_ & ~new_F7136_;
  assign new_F7138_ = new_F7102_ | new_F7135_;
  assign new_F7139_ = ~F7092 & F7093;
  assign new_F7140_ = F7092 & ~F7093;
  assign new_F7141_ = new_F7109_ | new_F7146_;
  assign new_F7142_ = ~new_F7109_ & ~new_F7145_;
  assign new_F7143_ = F7092 | new_F7109_;
  assign new_F7144_ = F7092 | F7093;
  assign new_F7145_ = new_F7109_ & new_F7146_;
  assign new_F7146_ = ~F7091 | ~new_F7116_;
  assign new_F7147_ = new_F7124_ & new_F7144_;
  assign new_F7148_ = ~new_F7124_ & ~new_F7144_;
  assign new_F7149_ = new_F7153_ | new_F7154_;
  assign new_F7150_ = ~F7095 & new_F7109_;
  assign new_F7151_ = new_F7155_ | new_F7156_;
  assign new_F7152_ = F7095 & new_F7109_;
  assign new_F7153_ = ~F7095 & ~new_F7109_;
  assign new_F7154_ = F7095 & ~new_F7109_;
  assign new_F7155_ = F7095 & ~new_F7109_;
  assign new_F7156_ = ~F7095 & new_F7109_;
  assign new_F7163_ = new_F7170_ & new_F7169_;
  assign new_F7164_ = new_F7172_ | new_F7171_;
  assign new_F7165_ = new_F7174_ | new_F7173_;
  assign new_F7166_ = new_F7176_ & new_F7175_;
  assign new_F7167_ = new_F7176_ & new_F7177_;
  assign new_F7168_ = new_F7169_ | new_F7178_;
  assign new_F7169_ = F7158 | new_F7181_;
  assign new_F7170_ = new_F7180_ | new_F7179_;
  assign new_F7171_ = new_F7185_ & new_F7184_;
  assign new_F7172_ = new_F7183_ & new_F7182_;
  assign new_F7173_ = new_F7188_ | new_F7187_;
  assign new_F7174_ = new_F7183_ & new_F7186_;
  assign new_F7175_ = F7158 | new_F7191_;
  assign new_F7176_ = new_F7190_ | new_F7189_;
  assign new_F7177_ = new_F7193_ | new_F7192_;
  assign new_F7178_ = ~new_F7169_ & new_F7195_;
  assign new_F7179_ = ~new_F7171_ & new_F7183_;
  assign new_F7180_ = new_F7171_ & ~new_F7183_;
  assign new_F7181_ = F7157 & ~F7158;
  assign new_F7182_ = ~new_F7204_ | ~new_F7205_;
  assign new_F7183_ = new_F7197_ | new_F7199_;
  assign new_F7184_ = new_F7207_ | new_F7206_;
  assign new_F7185_ = new_F7201_ | new_F7200_;
  assign new_F7186_ = ~new_F7209_ | ~new_F7208_;
  assign new_F7187_ = ~new_F7210_ & new_F7211_;
  assign new_F7188_ = new_F7210_ & ~new_F7211_;
  assign new_F7189_ = ~F7157 & F7158;
  assign new_F7190_ = F7157 & ~F7158;
  assign new_F7191_ = ~new_F7173_ | new_F7183_;
  assign new_F7192_ = new_F7173_ & new_F7183_;
  assign new_F7193_ = ~new_F7173_ & ~new_F7183_;
  assign new_F7194_ = new_F7215_ | new_F7214_;
  assign new_F7195_ = F7161 | new_F7194_;
  assign new_F7196_ = new_F7219_ | new_F7218_;
  assign new_F7197_ = ~F7161 & new_F7196_;
  assign new_F7198_ = new_F7217_ | new_F7216_;
  assign new_F7199_ = F7161 & new_F7198_;
  assign new_F7200_ = F7159 & ~new_F7169_;
  assign new_F7201_ = ~F7159 & new_F7169_;
  assign new_F7202_ = ~F7158 | ~new_F7183_;
  assign new_F7203_ = new_F7169_ & new_F7202_;
  assign new_F7204_ = ~new_F7169_ & ~new_F7203_;
  assign new_F7205_ = new_F7169_ | new_F7202_;
  assign new_F7206_ = ~F7159 & F7160;
  assign new_F7207_ = F7159 & ~F7160;
  assign new_F7208_ = new_F7176_ | new_F7213_;
  assign new_F7209_ = ~new_F7176_ & ~new_F7212_;
  assign new_F7210_ = F7159 | new_F7176_;
  assign new_F7211_ = F7159 | F7160;
  assign new_F7212_ = new_F7176_ & new_F7213_;
  assign new_F7213_ = ~F7158 | ~new_F7183_;
  assign new_F7214_ = new_F7191_ & new_F7211_;
  assign new_F7215_ = ~new_F7191_ & ~new_F7211_;
  assign new_F7216_ = new_F7220_ | new_F7221_;
  assign new_F7217_ = ~F7162 & new_F7176_;
  assign new_F7218_ = new_F7222_ | new_F7223_;
  assign new_F7219_ = F7162 & new_F7176_;
  assign new_F7220_ = ~F7162 & ~new_F7176_;
  assign new_F7221_ = F7162 & ~new_F7176_;
  assign new_F7222_ = F7162 & ~new_F7176_;
  assign new_F7223_ = ~F7162 & new_F7176_;
  assign new_F7230_ = new_F7237_ & new_F7236_;
  assign new_F7231_ = new_F7239_ | new_F7238_;
  assign new_F7232_ = new_F7241_ | new_F7240_;
  assign new_F7233_ = new_F7243_ & new_F7242_;
  assign new_F7234_ = new_F7243_ & new_F7244_;
  assign new_F7235_ = new_F7236_ | new_F7245_;
  assign new_F7236_ = F7225 | new_F7248_;
  assign new_F7237_ = new_F7247_ | new_F7246_;
  assign new_F7238_ = new_F7252_ & new_F7251_;
  assign new_F7239_ = new_F7250_ & new_F7249_;
  assign new_F7240_ = new_F7255_ | new_F7254_;
  assign new_F7241_ = new_F7250_ & new_F7253_;
  assign new_F7242_ = F7225 | new_F7258_;
  assign new_F7243_ = new_F7257_ | new_F7256_;
  assign new_F7244_ = new_F7260_ | new_F7259_;
  assign new_F7245_ = ~new_F7236_ & new_F7262_;
  assign new_F7246_ = ~new_F7238_ & new_F7250_;
  assign new_F7247_ = new_F7238_ & ~new_F7250_;
  assign new_F7248_ = F7224 & ~F7225;
  assign new_F7249_ = ~new_F7271_ | ~new_F7272_;
  assign new_F7250_ = new_F7264_ | new_F7266_;
  assign new_F7251_ = new_F7274_ | new_F7273_;
  assign new_F7252_ = new_F7268_ | new_F7267_;
  assign new_F7253_ = ~new_F7276_ | ~new_F7275_;
  assign new_F7254_ = ~new_F7277_ & new_F7278_;
  assign new_F7255_ = new_F7277_ & ~new_F7278_;
  assign new_F7256_ = ~F7224 & F7225;
  assign new_F7257_ = F7224 & ~F7225;
  assign new_F7258_ = ~new_F7240_ | new_F7250_;
  assign new_F7259_ = new_F7240_ & new_F7250_;
  assign new_F7260_ = ~new_F7240_ & ~new_F7250_;
  assign new_F7261_ = new_F7282_ | new_F7281_;
  assign new_F7262_ = F7228 | new_F7261_;
  assign new_F7263_ = new_F7286_ | new_F7285_;
  assign new_F7264_ = ~F7228 & new_F7263_;
  assign new_F7265_ = new_F7284_ | new_F7283_;
  assign new_F7266_ = F7228 & new_F7265_;
  assign new_F7267_ = F7226 & ~new_F7236_;
  assign new_F7268_ = ~F7226 & new_F7236_;
  assign new_F7269_ = ~F7225 | ~new_F7250_;
  assign new_F7270_ = new_F7236_ & new_F7269_;
  assign new_F7271_ = ~new_F7236_ & ~new_F7270_;
  assign new_F7272_ = new_F7236_ | new_F7269_;
  assign new_F7273_ = ~F7226 & F7227;
  assign new_F7274_ = F7226 & ~F7227;
  assign new_F7275_ = new_F7243_ | new_F7280_;
  assign new_F7276_ = ~new_F7243_ & ~new_F7279_;
  assign new_F7277_ = F7226 | new_F7243_;
  assign new_F7278_ = F7226 | F7227;
  assign new_F7279_ = new_F7243_ & new_F7280_;
  assign new_F7280_ = ~F7225 | ~new_F7250_;
  assign new_F7281_ = new_F7258_ & new_F7278_;
  assign new_F7282_ = ~new_F7258_ & ~new_F7278_;
  assign new_F7283_ = new_F7287_ | new_F7288_;
  assign new_F7284_ = ~F7229 & new_F7243_;
  assign new_F7285_ = new_F7289_ | new_F7290_;
  assign new_F7286_ = F7229 & new_F7243_;
  assign new_F7287_ = ~F7229 & ~new_F7243_;
  assign new_F7288_ = F7229 & ~new_F7243_;
  assign new_F7289_ = F7229 & ~new_F7243_;
  assign new_F7290_ = ~F7229 & new_F7243_;
  assign new_F7297_ = new_F7304_ & new_F7303_;
  assign new_F7298_ = new_F7306_ | new_F7305_;
  assign new_F7299_ = new_F7308_ | new_F7307_;
  assign new_F7300_ = new_F7310_ & new_F7309_;
  assign new_F7301_ = new_F7310_ & new_F7311_;
  assign new_F7302_ = new_F7303_ | new_F7312_;
  assign new_F7303_ = F7292 | new_F7315_;
  assign new_F7304_ = new_F7314_ | new_F7313_;
  assign new_F7305_ = new_F7319_ & new_F7318_;
  assign new_F7306_ = new_F7317_ & new_F7316_;
  assign new_F7307_ = new_F7322_ | new_F7321_;
  assign new_F7308_ = new_F7317_ & new_F7320_;
  assign new_F7309_ = F7292 | new_F7325_;
  assign new_F7310_ = new_F7324_ | new_F7323_;
  assign new_F7311_ = new_F7327_ | new_F7326_;
  assign new_F7312_ = ~new_F7303_ & new_F7329_;
  assign new_F7313_ = ~new_F7305_ & new_F7317_;
  assign new_F7314_ = new_F7305_ & ~new_F7317_;
  assign new_F7315_ = F7291 & ~F7292;
  assign new_F7316_ = ~new_F7338_ | ~new_F7339_;
  assign new_F7317_ = new_F7331_ | new_F7333_;
  assign new_F7318_ = new_F7341_ | new_F7340_;
  assign new_F7319_ = new_F7335_ | new_F7334_;
  assign new_F7320_ = ~new_F7343_ | ~new_F7342_;
  assign new_F7321_ = ~new_F7344_ & new_F7345_;
  assign new_F7322_ = new_F7344_ & ~new_F7345_;
  assign new_F7323_ = ~F7291 & F7292;
  assign new_F7324_ = F7291 & ~F7292;
  assign new_F7325_ = ~new_F7307_ | new_F7317_;
  assign new_F7326_ = new_F7307_ & new_F7317_;
  assign new_F7327_ = ~new_F7307_ & ~new_F7317_;
  assign new_F7328_ = new_F7349_ | new_F7348_;
  assign new_F7329_ = F7295 | new_F7328_;
  assign new_F7330_ = new_F7353_ | new_F7352_;
  assign new_F7331_ = ~F7295 & new_F7330_;
  assign new_F7332_ = new_F7351_ | new_F7350_;
  assign new_F7333_ = F7295 & new_F7332_;
  assign new_F7334_ = F7293 & ~new_F7303_;
  assign new_F7335_ = ~F7293 & new_F7303_;
  assign new_F7336_ = ~F7292 | ~new_F7317_;
  assign new_F7337_ = new_F7303_ & new_F7336_;
  assign new_F7338_ = ~new_F7303_ & ~new_F7337_;
  assign new_F7339_ = new_F7303_ | new_F7336_;
  assign new_F7340_ = ~F7293 & F7294;
  assign new_F7341_ = F7293 & ~F7294;
  assign new_F7342_ = new_F7310_ | new_F7347_;
  assign new_F7343_ = ~new_F7310_ & ~new_F7346_;
  assign new_F7344_ = F7293 | new_F7310_;
  assign new_F7345_ = F7293 | F7294;
  assign new_F7346_ = new_F7310_ & new_F7347_;
  assign new_F7347_ = ~F7292 | ~new_F7317_;
  assign new_F7348_ = new_F7325_ & new_F7345_;
  assign new_F7349_ = ~new_F7325_ & ~new_F7345_;
  assign new_F7350_ = new_F7354_ | new_F7355_;
  assign new_F7351_ = ~F7296 & new_F7310_;
  assign new_F7352_ = new_F7356_ | new_F7357_;
  assign new_F7353_ = F7296 & new_F7310_;
  assign new_F7354_ = ~F7296 & ~new_F7310_;
  assign new_F7355_ = F7296 & ~new_F7310_;
  assign new_F7356_ = F7296 & ~new_F7310_;
  assign new_F7357_ = ~F7296 & new_F7310_;
  assign new_F7364_ = new_F7371_ & new_F7370_;
  assign new_F7365_ = new_F7373_ | new_F7372_;
  assign new_F7366_ = new_F7375_ | new_F7374_;
  assign new_F7367_ = new_F7377_ & new_F7376_;
  assign new_F7368_ = new_F7377_ & new_F7378_;
  assign new_F7369_ = new_F7370_ | new_F7379_;
  assign new_F7370_ = F7359 | new_F7382_;
  assign new_F7371_ = new_F7381_ | new_F7380_;
  assign new_F7372_ = new_F7386_ & new_F7385_;
  assign new_F7373_ = new_F7384_ & new_F7383_;
  assign new_F7374_ = new_F7389_ | new_F7388_;
  assign new_F7375_ = new_F7384_ & new_F7387_;
  assign new_F7376_ = F7359 | new_F7392_;
  assign new_F7377_ = new_F7391_ | new_F7390_;
  assign new_F7378_ = new_F7394_ | new_F7393_;
  assign new_F7379_ = ~new_F7370_ & new_F7396_;
  assign new_F7380_ = ~new_F7372_ & new_F7384_;
  assign new_F7381_ = new_F7372_ & ~new_F7384_;
  assign new_F7382_ = F7358 & ~F7359;
  assign new_F7383_ = ~new_F7405_ | ~new_F7406_;
  assign new_F7384_ = new_F7398_ | new_F7400_;
  assign new_F7385_ = new_F7408_ | new_F7407_;
  assign new_F7386_ = new_F7402_ | new_F7401_;
  assign new_F7387_ = ~new_F7410_ | ~new_F7409_;
  assign new_F7388_ = ~new_F7411_ & new_F7412_;
  assign new_F7389_ = new_F7411_ & ~new_F7412_;
  assign new_F7390_ = ~F7358 & F7359;
  assign new_F7391_ = F7358 & ~F7359;
  assign new_F7392_ = ~new_F7374_ | new_F7384_;
  assign new_F7393_ = new_F7374_ & new_F7384_;
  assign new_F7394_ = ~new_F7374_ & ~new_F7384_;
  assign new_F7395_ = new_F7416_ | new_F7415_;
  assign new_F7396_ = F7362 | new_F7395_;
  assign new_F7397_ = new_F7420_ | new_F7419_;
  assign new_F7398_ = ~F7362 & new_F7397_;
  assign new_F7399_ = new_F7418_ | new_F7417_;
  assign new_F7400_ = F7362 & new_F7399_;
  assign new_F7401_ = F7360 & ~new_F7370_;
  assign new_F7402_ = ~F7360 & new_F7370_;
  assign new_F7403_ = ~F7359 | ~new_F7384_;
  assign new_F7404_ = new_F7370_ & new_F7403_;
  assign new_F7405_ = ~new_F7370_ & ~new_F7404_;
  assign new_F7406_ = new_F7370_ | new_F7403_;
  assign new_F7407_ = ~F7360 & F7361;
  assign new_F7408_ = F7360 & ~F7361;
  assign new_F7409_ = new_F7377_ | new_F7414_;
  assign new_F7410_ = ~new_F7377_ & ~new_F7413_;
  assign new_F7411_ = F7360 | new_F7377_;
  assign new_F7412_ = F7360 | F7361;
  assign new_F7413_ = new_F7377_ & new_F7414_;
  assign new_F7414_ = ~F7359 | ~new_F7384_;
  assign new_F7415_ = new_F7392_ & new_F7412_;
  assign new_F7416_ = ~new_F7392_ & ~new_F7412_;
  assign new_F7417_ = new_F7421_ | new_F7422_;
  assign new_F7418_ = ~F7363 & new_F7377_;
  assign new_F7419_ = new_F7423_ | new_F7424_;
  assign new_F7420_ = F7363 & new_F7377_;
  assign new_F7421_ = ~F7363 & ~new_F7377_;
  assign new_F7422_ = F7363 & ~new_F7377_;
  assign new_F7423_ = F7363 & ~new_F7377_;
  assign new_F7424_ = ~F7363 & new_F7377_;
  assign new_F7431_ = new_F7438_ & new_F7437_;
  assign new_F7432_ = new_F7440_ | new_F7439_;
  assign new_F7433_ = new_F7442_ | new_F7441_;
  assign new_F7434_ = new_F7444_ & new_F7443_;
  assign new_F7435_ = new_F7444_ & new_F7445_;
  assign new_F7436_ = new_F7437_ | new_F7446_;
  assign new_F7437_ = F7426 | new_F7449_;
  assign new_F7438_ = new_F7448_ | new_F7447_;
  assign new_F7439_ = new_F7453_ & new_F7452_;
  assign new_F7440_ = new_F7451_ & new_F7450_;
  assign new_F7441_ = new_F7456_ | new_F7455_;
  assign new_F7442_ = new_F7451_ & new_F7454_;
  assign new_F7443_ = F7426 | new_F7459_;
  assign new_F7444_ = new_F7458_ | new_F7457_;
  assign new_F7445_ = new_F7461_ | new_F7460_;
  assign new_F7446_ = ~new_F7437_ & new_F7463_;
  assign new_F7447_ = ~new_F7439_ & new_F7451_;
  assign new_F7448_ = new_F7439_ & ~new_F7451_;
  assign new_F7449_ = F7425 & ~F7426;
  assign new_F7450_ = ~new_F7472_ | ~new_F7473_;
  assign new_F7451_ = new_F7465_ | new_F7467_;
  assign new_F7452_ = new_F7475_ | new_F7474_;
  assign new_F7453_ = new_F7469_ | new_F7468_;
  assign new_F7454_ = ~new_F7477_ | ~new_F7476_;
  assign new_F7455_ = ~new_F7478_ & new_F7479_;
  assign new_F7456_ = new_F7478_ & ~new_F7479_;
  assign new_F7457_ = ~F7425 & F7426;
  assign new_F7458_ = F7425 & ~F7426;
  assign new_F7459_ = ~new_F7441_ | new_F7451_;
  assign new_F7460_ = new_F7441_ & new_F7451_;
  assign new_F7461_ = ~new_F7441_ & ~new_F7451_;
  assign new_F7462_ = new_F7483_ | new_F7482_;
  assign new_F7463_ = F7429 | new_F7462_;
  assign new_F7464_ = new_F7487_ | new_F7486_;
  assign new_F7465_ = ~F7429 & new_F7464_;
  assign new_F7466_ = new_F7485_ | new_F7484_;
  assign new_F7467_ = F7429 & new_F7466_;
  assign new_F7468_ = F7427 & ~new_F7437_;
  assign new_F7469_ = ~F7427 & new_F7437_;
  assign new_F7470_ = ~F7426 | ~new_F7451_;
  assign new_F7471_ = new_F7437_ & new_F7470_;
  assign new_F7472_ = ~new_F7437_ & ~new_F7471_;
  assign new_F7473_ = new_F7437_ | new_F7470_;
  assign new_F7474_ = ~F7427 & F7428;
  assign new_F7475_ = F7427 & ~F7428;
  assign new_F7476_ = new_F7444_ | new_F7481_;
  assign new_F7477_ = ~new_F7444_ & ~new_F7480_;
  assign new_F7478_ = F7427 | new_F7444_;
  assign new_F7479_ = F7427 | F7428;
  assign new_F7480_ = new_F7444_ & new_F7481_;
  assign new_F7481_ = ~F7426 | ~new_F7451_;
  assign new_F7482_ = new_F7459_ & new_F7479_;
  assign new_F7483_ = ~new_F7459_ & ~new_F7479_;
  assign new_F7484_ = new_F7488_ | new_F7489_;
  assign new_F7485_ = ~F7430 & new_F7444_;
  assign new_F7486_ = new_F7490_ | new_F7491_;
  assign new_F7487_ = F7430 & new_F7444_;
  assign new_F7488_ = ~F7430 & ~new_F7444_;
  assign new_F7489_ = F7430 & ~new_F7444_;
  assign new_F7490_ = F7430 & ~new_F7444_;
  assign new_F7491_ = ~F7430 & new_F7444_;
  assign new_F7498_ = new_F7505_ & new_F7504_;
  assign new_F7499_ = new_F7507_ | new_F7506_;
  assign new_F7500_ = new_F7509_ | new_F7508_;
  assign new_F7501_ = new_F7511_ & new_F7510_;
  assign new_F7502_ = new_F7511_ & new_F7512_;
  assign new_F7503_ = new_F7504_ | new_F7513_;
  assign new_F7504_ = F7493 | new_F7516_;
  assign new_F7505_ = new_F7515_ | new_F7514_;
  assign new_F7506_ = new_F7520_ & new_F7519_;
  assign new_F7507_ = new_F7518_ & new_F7517_;
  assign new_F7508_ = new_F7523_ | new_F7522_;
  assign new_F7509_ = new_F7518_ & new_F7521_;
  assign new_F7510_ = F7493 | new_F7526_;
  assign new_F7511_ = new_F7525_ | new_F7524_;
  assign new_F7512_ = new_F7528_ | new_F7527_;
  assign new_F7513_ = ~new_F7504_ & new_F7530_;
  assign new_F7514_ = ~new_F7506_ & new_F7518_;
  assign new_F7515_ = new_F7506_ & ~new_F7518_;
  assign new_F7516_ = F7492 & ~F7493;
  assign new_F7517_ = ~new_F7539_ | ~new_F7540_;
  assign new_F7518_ = new_F7532_ | new_F7534_;
  assign new_F7519_ = new_F7542_ | new_F7541_;
  assign new_F7520_ = new_F7536_ | new_F7535_;
  assign new_F7521_ = ~new_F7544_ | ~new_F7543_;
  assign new_F7522_ = ~new_F7545_ & new_F7546_;
  assign new_F7523_ = new_F7545_ & ~new_F7546_;
  assign new_F7524_ = ~F7492 & F7493;
  assign new_F7525_ = F7492 & ~F7493;
  assign new_F7526_ = ~new_F7508_ | new_F7518_;
  assign new_F7527_ = new_F7508_ & new_F7518_;
  assign new_F7528_ = ~new_F7508_ & ~new_F7518_;
  assign new_F7529_ = new_F7550_ | new_F7549_;
  assign new_F7530_ = F7496 | new_F7529_;
  assign new_F7531_ = new_F7554_ | new_F7553_;
  assign new_F7532_ = ~F7496 & new_F7531_;
  assign new_F7533_ = new_F7552_ | new_F7551_;
  assign new_F7534_ = F7496 & new_F7533_;
  assign new_F7535_ = F7494 & ~new_F7504_;
  assign new_F7536_ = ~F7494 & new_F7504_;
  assign new_F7537_ = ~F7493 | ~new_F7518_;
  assign new_F7538_ = new_F7504_ & new_F7537_;
  assign new_F7539_ = ~new_F7504_ & ~new_F7538_;
  assign new_F7540_ = new_F7504_ | new_F7537_;
  assign new_F7541_ = ~F7494 & F7495;
  assign new_F7542_ = F7494 & ~F7495;
  assign new_F7543_ = new_F7511_ | new_F7548_;
  assign new_F7544_ = ~new_F7511_ & ~new_F7547_;
  assign new_F7545_ = F7494 | new_F7511_;
  assign new_F7546_ = F7494 | F7495;
  assign new_F7547_ = new_F7511_ & new_F7548_;
  assign new_F7548_ = ~F7493 | ~new_F7518_;
  assign new_F7549_ = new_F7526_ & new_F7546_;
  assign new_F7550_ = ~new_F7526_ & ~new_F7546_;
  assign new_F7551_ = new_F7555_ | new_F7556_;
  assign new_F7552_ = ~F7497 & new_F7511_;
  assign new_F7553_ = new_F7557_ | new_F7558_;
  assign new_F7554_ = F7497 & new_F7511_;
  assign new_F7555_ = ~F7497 & ~new_F7511_;
  assign new_F7556_ = F7497 & ~new_F7511_;
  assign new_F7557_ = F7497 & ~new_F7511_;
  assign new_F7558_ = ~F7497 & new_F7511_;
  assign new_F7565_ = new_F7572_ & new_F7571_;
  assign new_F7566_ = new_F7574_ | new_F7573_;
  assign new_F7567_ = new_F7576_ | new_F7575_;
  assign new_F7568_ = new_F7578_ & new_F7577_;
  assign new_F7569_ = new_F7578_ & new_F7579_;
  assign new_F7570_ = new_F7571_ | new_F7580_;
  assign new_F7571_ = F7560 | new_F7583_;
  assign new_F7572_ = new_F7582_ | new_F7581_;
  assign new_F7573_ = new_F7587_ & new_F7586_;
  assign new_F7574_ = new_F7585_ & new_F7584_;
  assign new_F7575_ = new_F7590_ | new_F7589_;
  assign new_F7576_ = new_F7585_ & new_F7588_;
  assign new_F7577_ = F7560 | new_F7593_;
  assign new_F7578_ = new_F7592_ | new_F7591_;
  assign new_F7579_ = new_F7595_ | new_F7594_;
  assign new_F7580_ = ~new_F7571_ & new_F7597_;
  assign new_F7581_ = ~new_F7573_ & new_F7585_;
  assign new_F7582_ = new_F7573_ & ~new_F7585_;
  assign new_F7583_ = F7559 & ~F7560;
  assign new_F7584_ = ~new_F7606_ | ~new_F7607_;
  assign new_F7585_ = new_F7599_ | new_F7601_;
  assign new_F7586_ = new_F7609_ | new_F7608_;
  assign new_F7587_ = new_F7603_ | new_F7602_;
  assign new_F7588_ = ~new_F7611_ | ~new_F7610_;
  assign new_F7589_ = ~new_F7612_ & new_F7613_;
  assign new_F7590_ = new_F7612_ & ~new_F7613_;
  assign new_F7591_ = ~F7559 & F7560;
  assign new_F7592_ = F7559 & ~F7560;
  assign new_F7593_ = ~new_F7575_ | new_F7585_;
  assign new_F7594_ = new_F7575_ & new_F7585_;
  assign new_F7595_ = ~new_F7575_ & ~new_F7585_;
  assign new_F7596_ = new_F7617_ | new_F7616_;
  assign new_F7597_ = F7563 | new_F7596_;
  assign new_F7598_ = new_F7621_ | new_F7620_;
  assign new_F7599_ = ~F7563 & new_F7598_;
  assign new_F7600_ = new_F7619_ | new_F7618_;
  assign new_F7601_ = F7563 & new_F7600_;
  assign new_F7602_ = F7561 & ~new_F7571_;
  assign new_F7603_ = ~F7561 & new_F7571_;
  assign new_F7604_ = ~F7560 | ~new_F7585_;
  assign new_F7605_ = new_F7571_ & new_F7604_;
  assign new_F7606_ = ~new_F7571_ & ~new_F7605_;
  assign new_F7607_ = new_F7571_ | new_F7604_;
  assign new_F7608_ = ~F7561 & F7562;
  assign new_F7609_ = F7561 & ~F7562;
  assign new_F7610_ = new_F7578_ | new_F7615_;
  assign new_F7611_ = ~new_F7578_ & ~new_F7614_;
  assign new_F7612_ = F7561 | new_F7578_;
  assign new_F7613_ = F7561 | F7562;
  assign new_F7614_ = new_F7578_ & new_F7615_;
  assign new_F7615_ = ~F7560 | ~new_F7585_;
  assign new_F7616_ = new_F7593_ & new_F7613_;
  assign new_F7617_ = ~new_F7593_ & ~new_F7613_;
  assign new_F7618_ = new_F7622_ | new_F7623_;
  assign new_F7619_ = ~F7564 & new_F7578_;
  assign new_F7620_ = new_F7624_ | new_F7625_;
  assign new_F7621_ = F7564 & new_F7578_;
  assign new_F7622_ = ~F7564 & ~new_F7578_;
  assign new_F7623_ = F7564 & ~new_F7578_;
  assign new_F7624_ = F7564 & ~new_F7578_;
  assign new_F7625_ = ~F7564 & new_F7578_;
  assign new_F7632_ = new_F7639_ & new_F7638_;
  assign new_F7633_ = new_F7641_ | new_F7640_;
  assign new_F7634_ = new_F7643_ | new_F7642_;
  assign new_F7635_ = new_F7645_ & new_F7644_;
  assign new_F7636_ = new_F7645_ & new_F7646_;
  assign new_F7637_ = new_F7638_ | new_F7647_;
  assign new_F7638_ = F7627 | new_F7650_;
  assign new_F7639_ = new_F7649_ | new_F7648_;
  assign new_F7640_ = new_F7654_ & new_F7653_;
  assign new_F7641_ = new_F7652_ & new_F7651_;
  assign new_F7642_ = new_F7657_ | new_F7656_;
  assign new_F7643_ = new_F7652_ & new_F7655_;
  assign new_F7644_ = F7627 | new_F7660_;
  assign new_F7645_ = new_F7659_ | new_F7658_;
  assign new_F7646_ = new_F7662_ | new_F7661_;
  assign new_F7647_ = ~new_F7638_ & new_F7664_;
  assign new_F7648_ = ~new_F7640_ & new_F7652_;
  assign new_F7649_ = new_F7640_ & ~new_F7652_;
  assign new_F7650_ = F7626 & ~F7627;
  assign new_F7651_ = ~new_F7673_ | ~new_F7674_;
  assign new_F7652_ = new_F7666_ | new_F7668_;
  assign new_F7653_ = new_F7676_ | new_F7675_;
  assign new_F7654_ = new_F7670_ | new_F7669_;
  assign new_F7655_ = ~new_F7678_ | ~new_F7677_;
  assign new_F7656_ = ~new_F7679_ & new_F7680_;
  assign new_F7657_ = new_F7679_ & ~new_F7680_;
  assign new_F7658_ = ~F7626 & F7627;
  assign new_F7659_ = F7626 & ~F7627;
  assign new_F7660_ = ~new_F7642_ | new_F7652_;
  assign new_F7661_ = new_F7642_ & new_F7652_;
  assign new_F7662_ = ~new_F7642_ & ~new_F7652_;
  assign new_F7663_ = new_F7684_ | new_F7683_;
  assign new_F7664_ = F7630 | new_F7663_;
  assign new_F7665_ = new_F7688_ | new_F7687_;
  assign new_F7666_ = ~F7630 & new_F7665_;
  assign new_F7667_ = new_F7686_ | new_F7685_;
  assign new_F7668_ = F7630 & new_F7667_;
  assign new_F7669_ = F7628 & ~new_F7638_;
  assign new_F7670_ = ~F7628 & new_F7638_;
  assign new_F7671_ = ~F7627 | ~new_F7652_;
  assign new_F7672_ = new_F7638_ & new_F7671_;
  assign new_F7673_ = ~new_F7638_ & ~new_F7672_;
  assign new_F7674_ = new_F7638_ | new_F7671_;
  assign new_F7675_ = ~F7628 & F7629;
  assign new_F7676_ = F7628 & ~F7629;
  assign new_F7677_ = new_F7645_ | new_F7682_;
  assign new_F7678_ = ~new_F7645_ & ~new_F7681_;
  assign new_F7679_ = F7628 | new_F7645_;
  assign new_F7680_ = F7628 | F7629;
  assign new_F7681_ = new_F7645_ & new_F7682_;
  assign new_F7682_ = ~F7627 | ~new_F7652_;
  assign new_F7683_ = new_F7660_ & new_F7680_;
  assign new_F7684_ = ~new_F7660_ & ~new_F7680_;
  assign new_F7685_ = new_F7689_ | new_F7690_;
  assign new_F7686_ = ~F7631 & new_F7645_;
  assign new_F7687_ = new_F7691_ | new_F7692_;
  assign new_F7688_ = F7631 & new_F7645_;
  assign new_F7689_ = ~F7631 & ~new_F7645_;
  assign new_F7690_ = F7631 & ~new_F7645_;
  assign new_F7691_ = F7631 & ~new_F7645_;
  assign new_F7692_ = ~F7631 & new_F7645_;
  assign new_F7699_ = new_F7706_ & new_F7705_;
  assign new_F7700_ = new_F7708_ | new_F7707_;
  assign new_F7701_ = new_F7710_ | new_F7709_;
  assign new_F7702_ = new_F7712_ & new_F7711_;
  assign new_F7703_ = new_F7712_ & new_F7713_;
  assign new_F7704_ = new_F7705_ | new_F7714_;
  assign new_F7705_ = F7694 | new_F7717_;
  assign new_F7706_ = new_F7716_ | new_F7715_;
  assign new_F7707_ = new_F7721_ & new_F7720_;
  assign new_F7708_ = new_F7719_ & new_F7718_;
  assign new_F7709_ = new_F7724_ | new_F7723_;
  assign new_F7710_ = new_F7719_ & new_F7722_;
  assign new_F7711_ = F7694 | new_F7727_;
  assign new_F7712_ = new_F7726_ | new_F7725_;
  assign new_F7713_ = new_F7729_ | new_F7728_;
  assign new_F7714_ = ~new_F7705_ & new_F7731_;
  assign new_F7715_ = ~new_F7707_ & new_F7719_;
  assign new_F7716_ = new_F7707_ & ~new_F7719_;
  assign new_F7717_ = F7693 & ~F7694;
  assign new_F7718_ = ~new_F7740_ | ~new_F7741_;
  assign new_F7719_ = new_F7733_ | new_F7735_;
  assign new_F7720_ = new_F7743_ | new_F7742_;
  assign new_F7721_ = new_F7737_ | new_F7736_;
  assign new_F7722_ = ~new_F7745_ | ~new_F7744_;
  assign new_F7723_ = ~new_F7746_ & new_F7747_;
  assign new_F7724_ = new_F7746_ & ~new_F7747_;
  assign new_F7725_ = ~F7693 & F7694;
  assign new_F7726_ = F7693 & ~F7694;
  assign new_F7727_ = ~new_F7709_ | new_F7719_;
  assign new_F7728_ = new_F7709_ & new_F7719_;
  assign new_F7729_ = ~new_F7709_ & ~new_F7719_;
  assign new_F7730_ = new_F7751_ | new_F7750_;
  assign new_F7731_ = F7697 | new_F7730_;
  assign new_F7732_ = new_F7755_ | new_F7754_;
  assign new_F7733_ = ~F7697 & new_F7732_;
  assign new_F7734_ = new_F7753_ | new_F7752_;
  assign new_F7735_ = F7697 & new_F7734_;
  assign new_F7736_ = F7695 & ~new_F7705_;
  assign new_F7737_ = ~F7695 & new_F7705_;
  assign new_F7738_ = ~F7694 | ~new_F7719_;
  assign new_F7739_ = new_F7705_ & new_F7738_;
  assign new_F7740_ = ~new_F7705_ & ~new_F7739_;
  assign new_F7741_ = new_F7705_ | new_F7738_;
  assign new_F7742_ = ~F7695 & F7696;
  assign new_F7743_ = F7695 & ~F7696;
  assign new_F7744_ = new_F7712_ | new_F7749_;
  assign new_F7745_ = ~new_F7712_ & ~new_F7748_;
  assign new_F7746_ = F7695 | new_F7712_;
  assign new_F7747_ = F7695 | F7696;
  assign new_F7748_ = new_F7712_ & new_F7749_;
  assign new_F7749_ = ~F7694 | ~new_F7719_;
  assign new_F7750_ = new_F7727_ & new_F7747_;
  assign new_F7751_ = ~new_F7727_ & ~new_F7747_;
  assign new_F7752_ = new_F7756_ | new_F7757_;
  assign new_F7753_ = ~F7698 & new_F7712_;
  assign new_F7754_ = new_F7758_ | new_F7759_;
  assign new_F7755_ = F7698 & new_F7712_;
  assign new_F7756_ = ~F7698 & ~new_F7712_;
  assign new_F7757_ = F7698 & ~new_F7712_;
  assign new_F7758_ = F7698 & ~new_F7712_;
  assign new_F7759_ = ~F7698 & new_F7712_;
  assign new_F7766_ = new_F7773_ & new_F7772_;
  assign new_F7767_ = new_F7775_ | new_F7774_;
  assign new_F7768_ = new_F7777_ | new_F7776_;
  assign new_F7769_ = new_F7779_ & new_F7778_;
  assign new_F7770_ = new_F7779_ & new_F7780_;
  assign new_F7771_ = new_F7772_ | new_F7781_;
  assign new_F7772_ = F7761 | new_F7784_;
  assign new_F7773_ = new_F7783_ | new_F7782_;
  assign new_F7774_ = new_F7788_ & new_F7787_;
  assign new_F7775_ = new_F7786_ & new_F7785_;
  assign new_F7776_ = new_F7791_ | new_F7790_;
  assign new_F7777_ = new_F7786_ & new_F7789_;
  assign new_F7778_ = F7761 | new_F7794_;
  assign new_F7779_ = new_F7793_ | new_F7792_;
  assign new_F7780_ = new_F7796_ | new_F7795_;
  assign new_F7781_ = ~new_F7772_ & new_F7798_;
  assign new_F7782_ = ~new_F7774_ & new_F7786_;
  assign new_F7783_ = new_F7774_ & ~new_F7786_;
  assign new_F7784_ = F7760 & ~F7761;
  assign new_F7785_ = ~new_F7807_ | ~new_F7808_;
  assign new_F7786_ = new_F7800_ | new_F7802_;
  assign new_F7787_ = new_F7810_ | new_F7809_;
  assign new_F7788_ = new_F7804_ | new_F7803_;
  assign new_F7789_ = ~new_F7812_ | ~new_F7811_;
  assign new_F7790_ = ~new_F7813_ & new_F7814_;
  assign new_F7791_ = new_F7813_ & ~new_F7814_;
  assign new_F7792_ = ~F7760 & F7761;
  assign new_F7793_ = F7760 & ~F7761;
  assign new_F7794_ = ~new_F7776_ | new_F7786_;
  assign new_F7795_ = new_F7776_ & new_F7786_;
  assign new_F7796_ = ~new_F7776_ & ~new_F7786_;
  assign new_F7797_ = new_F7818_ | new_F7817_;
  assign new_F7798_ = F7764 | new_F7797_;
  assign new_F7799_ = new_F7822_ | new_F7821_;
  assign new_F7800_ = ~F7764 & new_F7799_;
  assign new_F7801_ = new_F7820_ | new_F7819_;
  assign new_F7802_ = F7764 & new_F7801_;
  assign new_F7803_ = F7762 & ~new_F7772_;
  assign new_F7804_ = ~F7762 & new_F7772_;
  assign new_F7805_ = ~F7761 | ~new_F7786_;
  assign new_F7806_ = new_F7772_ & new_F7805_;
  assign new_F7807_ = ~new_F7772_ & ~new_F7806_;
  assign new_F7808_ = new_F7772_ | new_F7805_;
  assign new_F7809_ = ~F7762 & F7763;
  assign new_F7810_ = F7762 & ~F7763;
  assign new_F7811_ = new_F7779_ | new_F7816_;
  assign new_F7812_ = ~new_F7779_ & ~new_F7815_;
  assign new_F7813_ = F7762 | new_F7779_;
  assign new_F7814_ = F7762 | F7763;
  assign new_F7815_ = new_F7779_ & new_F7816_;
  assign new_F7816_ = ~F7761 | ~new_F7786_;
  assign new_F7817_ = new_F7794_ & new_F7814_;
  assign new_F7818_ = ~new_F7794_ & ~new_F7814_;
  assign new_F7819_ = new_F7823_ | new_F7824_;
  assign new_F7820_ = ~F7765 & new_F7779_;
  assign new_F7821_ = new_F7825_ | new_F7826_;
  assign new_F7822_ = F7765 & new_F7779_;
  assign new_F7823_ = ~F7765 & ~new_F7779_;
  assign new_F7824_ = F7765 & ~new_F7779_;
  assign new_F7825_ = F7765 & ~new_F7779_;
  assign new_F7826_ = ~F7765 & new_F7779_;
  assign new_F7833_ = new_F7840_ & new_F7839_;
  assign new_F7834_ = new_F7842_ | new_F7841_;
  assign new_F7835_ = new_F7844_ | new_F7843_;
  assign new_F7836_ = new_F7846_ & new_F7845_;
  assign new_F7837_ = new_F7846_ & new_F7847_;
  assign new_F7838_ = new_F7839_ | new_F7848_;
  assign new_F7839_ = F7828 | new_F7851_;
  assign new_F7840_ = new_F7850_ | new_F7849_;
  assign new_F7841_ = new_F7855_ & new_F7854_;
  assign new_F7842_ = new_F7853_ & new_F7852_;
  assign new_F7843_ = new_F7858_ | new_F7857_;
  assign new_F7844_ = new_F7853_ & new_F7856_;
  assign new_F7845_ = F7828 | new_F7861_;
  assign new_F7846_ = new_F7860_ | new_F7859_;
  assign new_F7847_ = new_F7863_ | new_F7862_;
  assign new_F7848_ = ~new_F7839_ & new_F7865_;
  assign new_F7849_ = ~new_F7841_ & new_F7853_;
  assign new_F7850_ = new_F7841_ & ~new_F7853_;
  assign new_F7851_ = F7827 & ~F7828;
  assign new_F7852_ = ~new_F7874_ | ~new_F7875_;
  assign new_F7853_ = new_F7867_ | new_F7869_;
  assign new_F7854_ = new_F7877_ | new_F7876_;
  assign new_F7855_ = new_F7871_ | new_F7870_;
  assign new_F7856_ = ~new_F7879_ | ~new_F7878_;
  assign new_F7857_ = ~new_F7880_ & new_F7881_;
  assign new_F7858_ = new_F7880_ & ~new_F7881_;
  assign new_F7859_ = ~F7827 & F7828;
  assign new_F7860_ = F7827 & ~F7828;
  assign new_F7861_ = ~new_F7843_ | new_F7853_;
  assign new_F7862_ = new_F7843_ & new_F7853_;
  assign new_F7863_ = ~new_F7843_ & ~new_F7853_;
  assign new_F7864_ = new_F7885_ | new_F7884_;
  assign new_F7865_ = F7831 | new_F7864_;
  assign new_F7866_ = new_F7889_ | new_F7888_;
  assign new_F7867_ = ~F7831 & new_F7866_;
  assign new_F7868_ = new_F7887_ | new_F7886_;
  assign new_F7869_ = F7831 & new_F7868_;
  assign new_F7870_ = F7829 & ~new_F7839_;
  assign new_F7871_ = ~F7829 & new_F7839_;
  assign new_F7872_ = ~F7828 | ~new_F7853_;
  assign new_F7873_ = new_F7839_ & new_F7872_;
  assign new_F7874_ = ~new_F7839_ & ~new_F7873_;
  assign new_F7875_ = new_F7839_ | new_F7872_;
  assign new_F7876_ = ~F7829 & F7830;
  assign new_F7877_ = F7829 & ~F7830;
  assign new_F7878_ = new_F7846_ | new_F7883_;
  assign new_F7879_ = ~new_F7846_ & ~new_F7882_;
  assign new_F7880_ = F7829 | new_F7846_;
  assign new_F7881_ = F7829 | F7830;
  assign new_F7882_ = new_F7846_ & new_F7883_;
  assign new_F7883_ = ~F7828 | ~new_F7853_;
  assign new_F7884_ = new_F7861_ & new_F7881_;
  assign new_F7885_ = ~new_F7861_ & ~new_F7881_;
  assign new_F7886_ = new_F7890_ | new_F7891_;
  assign new_F7887_ = ~F7832 & new_F7846_;
  assign new_F7888_ = new_F7892_ | new_F7893_;
  assign new_F7889_ = F7832 & new_F7846_;
  assign new_F7890_ = ~F7832 & ~new_F7846_;
  assign new_F7891_ = F7832 & ~new_F7846_;
  assign new_F7892_ = F7832 & ~new_F7846_;
  assign new_F7893_ = ~F7832 & new_F7846_;
  assign new_F7900_ = new_F7907_ & new_F7906_;
  assign new_F7901_ = new_F7909_ | new_F7908_;
  assign new_F7902_ = new_F7911_ | new_F7910_;
  assign new_F7903_ = new_F7913_ & new_F7912_;
  assign new_F7904_ = new_F7913_ & new_F7914_;
  assign new_F7905_ = new_F7906_ | new_F7915_;
  assign new_F7906_ = F7895 | new_F7918_;
  assign new_F7907_ = new_F7917_ | new_F7916_;
  assign new_F7908_ = new_F7922_ & new_F7921_;
  assign new_F7909_ = new_F7920_ & new_F7919_;
  assign new_F7910_ = new_F7925_ | new_F7924_;
  assign new_F7911_ = new_F7920_ & new_F7923_;
  assign new_F7912_ = F7895 | new_F7928_;
  assign new_F7913_ = new_F7927_ | new_F7926_;
  assign new_F7914_ = new_F7930_ | new_F7929_;
  assign new_F7915_ = ~new_F7906_ & new_F7932_;
  assign new_F7916_ = ~new_F7908_ & new_F7920_;
  assign new_F7917_ = new_F7908_ & ~new_F7920_;
  assign new_F7918_ = F7894 & ~F7895;
  assign new_F7919_ = ~new_F7941_ | ~new_F7942_;
  assign new_F7920_ = new_F7934_ | new_F7936_;
  assign new_F7921_ = new_F7944_ | new_F7943_;
  assign new_F7922_ = new_F7938_ | new_F7937_;
  assign new_F7923_ = ~new_F7946_ | ~new_F7945_;
  assign new_F7924_ = ~new_F7947_ & new_F7948_;
  assign new_F7925_ = new_F7947_ & ~new_F7948_;
  assign new_F7926_ = ~F7894 & F7895;
  assign new_F7927_ = F7894 & ~F7895;
  assign new_F7928_ = ~new_F7910_ | new_F7920_;
  assign new_F7929_ = new_F7910_ & new_F7920_;
  assign new_F7930_ = ~new_F7910_ & ~new_F7920_;
  assign new_F7931_ = new_F7952_ | new_F7951_;
  assign new_F7932_ = F7898 | new_F7931_;
  assign new_F7933_ = new_F7956_ | new_F7955_;
  assign new_F7934_ = ~F7898 & new_F7933_;
  assign new_F7935_ = new_F7954_ | new_F7953_;
  assign new_F7936_ = F7898 & new_F7935_;
  assign new_F7937_ = F7896 & ~new_F7906_;
  assign new_F7938_ = ~F7896 & new_F7906_;
  assign new_F7939_ = ~F7895 | ~new_F7920_;
  assign new_F7940_ = new_F7906_ & new_F7939_;
  assign new_F7941_ = ~new_F7906_ & ~new_F7940_;
  assign new_F7942_ = new_F7906_ | new_F7939_;
  assign new_F7943_ = ~F7896 & F7897;
  assign new_F7944_ = F7896 & ~F7897;
  assign new_F7945_ = new_F7913_ | new_F7950_;
  assign new_F7946_ = ~new_F7913_ & ~new_F7949_;
  assign new_F7947_ = F7896 | new_F7913_;
  assign new_F7948_ = F7896 | F7897;
  assign new_F7949_ = new_F7913_ & new_F7950_;
  assign new_F7950_ = ~F7895 | ~new_F7920_;
  assign new_F7951_ = new_F7928_ & new_F7948_;
  assign new_F7952_ = ~new_F7928_ & ~new_F7948_;
  assign new_F7953_ = new_F7957_ | new_F7958_;
  assign new_F7954_ = ~F7899 & new_F7913_;
  assign new_F7955_ = new_F7959_ | new_F7960_;
  assign new_F7956_ = F7899 & new_F7913_;
  assign new_F7957_ = ~F7899 & ~new_F7913_;
  assign new_F7958_ = F7899 & ~new_F7913_;
  assign new_F7959_ = F7899 & ~new_F7913_;
  assign new_F7960_ = ~F7899 & new_F7913_;
  assign new_F7967_ = new_F7974_ & new_F7973_;
  assign new_F7968_ = new_F7976_ | new_F7975_;
  assign new_F7969_ = new_F7978_ | new_F7977_;
  assign new_F7970_ = new_F7980_ & new_F7979_;
  assign new_F7971_ = new_F7980_ & new_F7981_;
  assign new_F7972_ = new_F7973_ | new_F7982_;
  assign new_F7973_ = F7962 | new_F7985_;
  assign new_F7974_ = new_F7984_ | new_F7983_;
  assign new_F7975_ = new_F7989_ & new_F7988_;
  assign new_F7976_ = new_F7987_ & new_F7986_;
  assign new_F7977_ = new_F7992_ | new_F7991_;
  assign new_F7978_ = new_F7987_ & new_F7990_;
  assign new_F7979_ = F7962 | new_F7995_;
  assign new_F7980_ = new_F7994_ | new_F7993_;
  assign new_F7981_ = new_F7997_ | new_F7996_;
  assign new_F7982_ = ~new_F7973_ & new_F7999_;
  assign new_F7983_ = ~new_F7975_ & new_F7987_;
  assign new_F7984_ = new_F7975_ & ~new_F7987_;
  assign new_F7985_ = F7961 & ~F7962;
  assign new_F7986_ = ~new_F8008_ | ~new_F8009_;
  assign new_F7987_ = new_F8001_ | new_F8003_;
  assign new_F7988_ = new_F8011_ | new_F8010_;
  assign new_F7989_ = new_F8005_ | new_F8004_;
  assign new_F7990_ = ~new_F8013_ | ~new_F8012_;
  assign new_F7991_ = ~new_F8014_ & new_F8015_;
  assign new_F7992_ = new_F8014_ & ~new_F8015_;
  assign new_F7993_ = ~F7961 & F7962;
  assign new_F7994_ = F7961 & ~F7962;
  assign new_F7995_ = ~new_F7977_ | new_F7987_;
  assign new_F7996_ = new_F7977_ & new_F7987_;
  assign new_F7997_ = ~new_F7977_ & ~new_F7987_;
  assign new_F7998_ = new_F8019_ | new_F8018_;
  assign new_F7999_ = F7965 | new_F7998_;
  assign new_F8000_ = new_F8023_ | new_F8022_;
  assign new_F8001_ = ~F7965 & new_F8000_;
  assign new_F8002_ = new_F8021_ | new_F8020_;
  assign new_F8003_ = F7965 & new_F8002_;
  assign new_F8004_ = F7963 & ~new_F7973_;
  assign new_F8005_ = ~F7963 & new_F7973_;
  assign new_F8006_ = ~F7962 | ~new_F7987_;
  assign new_F8007_ = new_F7973_ & new_F8006_;
  assign new_F8008_ = ~new_F7973_ & ~new_F8007_;
  assign new_F8009_ = new_F7973_ | new_F8006_;
  assign new_F8010_ = ~F7963 & F7964;
  assign new_F8011_ = F7963 & ~F7964;
  assign new_F8012_ = new_F7980_ | new_F8017_;
  assign new_F8013_ = ~new_F7980_ & ~new_F8016_;
  assign new_F8014_ = F7963 | new_F7980_;
  assign new_F8015_ = F7963 | F7964;
  assign new_F8016_ = new_F7980_ & new_F8017_;
  assign new_F8017_ = ~F7962 | ~new_F7987_;
  assign new_F8018_ = new_F7995_ & new_F8015_;
  assign new_F8019_ = ~new_F7995_ & ~new_F8015_;
  assign new_F8020_ = new_F8024_ | new_F8025_;
  assign new_F8021_ = ~F7966 & new_F7980_;
  assign new_F8022_ = new_F8026_ | new_F8027_;
  assign new_F8023_ = F7966 & new_F7980_;
  assign new_F8024_ = ~F7966 & ~new_F7980_;
  assign new_F8025_ = F7966 & ~new_F7980_;
  assign new_F8026_ = F7966 & ~new_F7980_;
  assign new_F8027_ = ~F7966 & new_F7980_;
  assign new_F8034_ = new_F8041_ & new_F8040_;
  assign new_F8035_ = new_F8043_ | new_F8042_;
  assign new_F8036_ = new_F8045_ | new_F8044_;
  assign new_F8037_ = new_F8047_ & new_F8046_;
  assign new_F8038_ = new_F8047_ & new_F8048_;
  assign new_F8039_ = new_F8040_ | new_F8049_;
  assign new_F8040_ = F8029 | new_F8052_;
  assign new_F8041_ = new_F8051_ | new_F8050_;
  assign new_F8042_ = new_F8056_ & new_F8055_;
  assign new_F8043_ = new_F8054_ & new_F8053_;
  assign new_F8044_ = new_F8059_ | new_F8058_;
  assign new_F8045_ = new_F8054_ & new_F8057_;
  assign new_F8046_ = F8029 | new_F8062_;
  assign new_F8047_ = new_F8061_ | new_F8060_;
  assign new_F8048_ = new_F8064_ | new_F8063_;
  assign new_F8049_ = ~new_F8040_ & new_F8066_;
  assign new_F8050_ = ~new_F8042_ & new_F8054_;
  assign new_F8051_ = new_F8042_ & ~new_F8054_;
  assign new_F8052_ = F8028 & ~F8029;
  assign new_F8053_ = ~new_F8075_ | ~new_F8076_;
  assign new_F8054_ = new_F8068_ | new_F8070_;
  assign new_F8055_ = new_F8078_ | new_F8077_;
  assign new_F8056_ = new_F8072_ | new_F8071_;
  assign new_F8057_ = ~new_F8080_ | ~new_F8079_;
  assign new_F8058_ = ~new_F8081_ & new_F8082_;
  assign new_F8059_ = new_F8081_ & ~new_F8082_;
  assign new_F8060_ = ~F8028 & F8029;
  assign new_F8061_ = F8028 & ~F8029;
  assign new_F8062_ = ~new_F8044_ | new_F8054_;
  assign new_F8063_ = new_F8044_ & new_F8054_;
  assign new_F8064_ = ~new_F8044_ & ~new_F8054_;
  assign new_F8065_ = new_F8086_ | new_F8085_;
  assign new_F8066_ = F8032 | new_F8065_;
  assign new_F8067_ = new_F8090_ | new_F8089_;
  assign new_F8068_ = ~F8032 & new_F8067_;
  assign new_F8069_ = new_F8088_ | new_F8087_;
  assign new_F8070_ = F8032 & new_F8069_;
  assign new_F8071_ = F8030 & ~new_F8040_;
  assign new_F8072_ = ~F8030 & new_F8040_;
  assign new_F8073_ = ~F8029 | ~new_F8054_;
  assign new_F8074_ = new_F8040_ & new_F8073_;
  assign new_F8075_ = ~new_F8040_ & ~new_F8074_;
  assign new_F8076_ = new_F8040_ | new_F8073_;
  assign new_F8077_ = ~F8030 & F8031;
  assign new_F8078_ = F8030 & ~F8031;
  assign new_F8079_ = new_F8047_ | new_F8084_;
  assign new_F8080_ = ~new_F8047_ & ~new_F8083_;
  assign new_F8081_ = F8030 | new_F8047_;
  assign new_F8082_ = F8030 | F8031;
  assign new_F8083_ = new_F8047_ & new_F8084_;
  assign new_F8084_ = ~F8029 | ~new_F8054_;
  assign new_F8085_ = new_F8062_ & new_F8082_;
  assign new_F8086_ = ~new_F8062_ & ~new_F8082_;
  assign new_F8087_ = new_F8091_ | new_F8092_;
  assign new_F8088_ = ~F8033 & new_F8047_;
  assign new_F8089_ = new_F8093_ | new_F8094_;
  assign new_F8090_ = F8033 & new_F8047_;
  assign new_F8091_ = ~F8033 & ~new_F8047_;
  assign new_F8092_ = F8033 & ~new_F8047_;
  assign new_F8093_ = F8033 & ~new_F8047_;
  assign new_F8094_ = ~F8033 & new_F8047_;
  assign new_F8101_ = new_F8108_ & new_F8107_;
  assign new_F8102_ = new_F8110_ | new_F8109_;
  assign new_F8103_ = new_F8112_ | new_F8111_;
  assign new_F8104_ = new_F8114_ & new_F8113_;
  assign new_F8105_ = new_F8114_ & new_F8115_;
  assign new_F8106_ = new_F8107_ | new_F8116_;
  assign new_F8107_ = F8096 | new_F8119_;
  assign new_F8108_ = new_F8118_ | new_F8117_;
  assign new_F8109_ = new_F8123_ & new_F8122_;
  assign new_F8110_ = new_F8121_ & new_F8120_;
  assign new_F8111_ = new_F8126_ | new_F8125_;
  assign new_F8112_ = new_F8121_ & new_F8124_;
  assign new_F8113_ = F8096 | new_F8129_;
  assign new_F8114_ = new_F8128_ | new_F8127_;
  assign new_F8115_ = new_F8131_ | new_F8130_;
  assign new_F8116_ = ~new_F8107_ & new_F8133_;
  assign new_F8117_ = ~new_F8109_ & new_F8121_;
  assign new_F8118_ = new_F8109_ & ~new_F8121_;
  assign new_F8119_ = F8095 & ~F8096;
  assign new_F8120_ = ~new_F8142_ | ~new_F8143_;
  assign new_F8121_ = new_F8135_ | new_F8137_;
  assign new_F8122_ = new_F8145_ | new_F8144_;
  assign new_F8123_ = new_F8139_ | new_F8138_;
  assign new_F8124_ = ~new_F8147_ | ~new_F8146_;
  assign new_F8125_ = ~new_F8148_ & new_F8149_;
  assign new_F8126_ = new_F8148_ & ~new_F8149_;
  assign new_F8127_ = ~F8095 & F8096;
  assign new_F8128_ = F8095 & ~F8096;
  assign new_F8129_ = ~new_F8111_ | new_F8121_;
  assign new_F8130_ = new_F8111_ & new_F8121_;
  assign new_F8131_ = ~new_F8111_ & ~new_F8121_;
  assign new_F8132_ = new_F8153_ | new_F8152_;
  assign new_F8133_ = F8099 | new_F8132_;
  assign new_F8134_ = new_F8157_ | new_F8156_;
  assign new_F8135_ = ~F8099 & new_F8134_;
  assign new_F8136_ = new_F8155_ | new_F8154_;
  assign new_F8137_ = F8099 & new_F8136_;
  assign new_F8138_ = F8097 & ~new_F8107_;
  assign new_F8139_ = ~F8097 & new_F8107_;
  assign new_F8140_ = ~F8096 | ~new_F8121_;
  assign new_F8141_ = new_F8107_ & new_F8140_;
  assign new_F8142_ = ~new_F8107_ & ~new_F8141_;
  assign new_F8143_ = new_F8107_ | new_F8140_;
  assign new_F8144_ = ~F8097 & F8098;
  assign new_F8145_ = F8097 & ~F8098;
  assign new_F8146_ = new_F8114_ | new_F8151_;
  assign new_F8147_ = ~new_F8114_ & ~new_F8150_;
  assign new_F8148_ = F8097 | new_F8114_;
  assign new_F8149_ = F8097 | F8098;
  assign new_F8150_ = new_F8114_ & new_F8151_;
  assign new_F8151_ = ~F8096 | ~new_F8121_;
  assign new_F8152_ = new_F8129_ & new_F8149_;
  assign new_F8153_ = ~new_F8129_ & ~new_F8149_;
  assign new_F8154_ = new_F8158_ | new_F8159_;
  assign new_F8155_ = ~F8100 & new_F8114_;
  assign new_F8156_ = new_F8160_ | new_F8161_;
  assign new_F8157_ = F8100 & new_F8114_;
  assign new_F8158_ = ~F8100 & ~new_F8114_;
  assign new_F8159_ = F8100 & ~new_F8114_;
  assign new_F8160_ = F8100 & ~new_F8114_;
  assign new_F8161_ = ~F8100 & new_F8114_;
  assign new_F8168_ = new_F8175_ & new_F8174_;
  assign new_F8169_ = new_F8177_ | new_F8176_;
  assign new_F8170_ = new_F8179_ | new_F8178_;
  assign new_F8171_ = new_F8181_ & new_F8180_;
  assign new_F8172_ = new_F8181_ & new_F8182_;
  assign new_F8173_ = new_F8174_ | new_F8183_;
  assign new_F8174_ = F8163 | new_F8186_;
  assign new_F8175_ = new_F8185_ | new_F8184_;
  assign new_F8176_ = new_F8190_ & new_F8189_;
  assign new_F8177_ = new_F8188_ & new_F8187_;
  assign new_F8178_ = new_F8193_ | new_F8192_;
  assign new_F8179_ = new_F8188_ & new_F8191_;
  assign new_F8180_ = F8163 | new_F8196_;
  assign new_F8181_ = new_F8195_ | new_F8194_;
  assign new_F8182_ = new_F8198_ | new_F8197_;
  assign new_F8183_ = ~new_F8174_ & new_F8200_;
  assign new_F8184_ = ~new_F8176_ & new_F8188_;
  assign new_F8185_ = new_F8176_ & ~new_F8188_;
  assign new_F8186_ = F8162 & ~F8163;
  assign new_F8187_ = ~new_F8209_ | ~new_F8210_;
  assign new_F8188_ = new_F8202_ | new_F8204_;
  assign new_F8189_ = new_F8212_ | new_F8211_;
  assign new_F8190_ = new_F8206_ | new_F8205_;
  assign new_F8191_ = ~new_F8214_ | ~new_F8213_;
  assign new_F8192_ = ~new_F8215_ & new_F8216_;
  assign new_F8193_ = new_F8215_ & ~new_F8216_;
  assign new_F8194_ = ~F8162 & F8163;
  assign new_F8195_ = F8162 & ~F8163;
  assign new_F8196_ = ~new_F8178_ | new_F8188_;
  assign new_F8197_ = new_F8178_ & new_F8188_;
  assign new_F8198_ = ~new_F8178_ & ~new_F8188_;
  assign new_F8199_ = new_F8220_ | new_F8219_;
  assign new_F8200_ = F8166 | new_F8199_;
  assign new_F8201_ = new_F8224_ | new_F8223_;
  assign new_F8202_ = ~F8166 & new_F8201_;
  assign new_F8203_ = new_F8222_ | new_F8221_;
  assign new_F8204_ = F8166 & new_F8203_;
  assign new_F8205_ = F8164 & ~new_F8174_;
  assign new_F8206_ = ~F8164 & new_F8174_;
  assign new_F8207_ = ~F8163 | ~new_F8188_;
  assign new_F8208_ = new_F8174_ & new_F8207_;
  assign new_F8209_ = ~new_F8174_ & ~new_F8208_;
  assign new_F8210_ = new_F8174_ | new_F8207_;
  assign new_F8211_ = ~F8164 & F8165;
  assign new_F8212_ = F8164 & ~F8165;
  assign new_F8213_ = new_F8181_ | new_F8218_;
  assign new_F8214_ = ~new_F8181_ & ~new_F8217_;
  assign new_F8215_ = F8164 | new_F8181_;
  assign new_F8216_ = F8164 | F8165;
  assign new_F8217_ = new_F8181_ & new_F8218_;
  assign new_F8218_ = ~F8163 | ~new_F8188_;
  assign new_F8219_ = new_F8196_ & new_F8216_;
  assign new_F8220_ = ~new_F8196_ & ~new_F8216_;
  assign new_F8221_ = new_F8225_ | new_F8226_;
  assign new_F8222_ = ~F8167 & new_F8181_;
  assign new_F8223_ = new_F8227_ | new_F8228_;
  assign new_F8224_ = F8167 & new_F8181_;
  assign new_F8225_ = ~F8167 & ~new_F8181_;
  assign new_F8226_ = F8167 & ~new_F8181_;
  assign new_F8227_ = F8167 & ~new_F8181_;
  assign new_F8228_ = ~F8167 & new_F8181_;
  assign new_F8235_ = new_F8242_ & new_F8241_;
  assign new_F8236_ = new_F8244_ | new_F8243_;
  assign new_F8237_ = new_F8246_ | new_F8245_;
  assign new_F8238_ = new_F8248_ & new_F8247_;
  assign new_F8239_ = new_F8248_ & new_F8249_;
  assign new_F8240_ = new_F8241_ | new_F8250_;
  assign new_F8241_ = F8230 | new_F8253_;
  assign new_F8242_ = new_F8252_ | new_F8251_;
  assign new_F8243_ = new_F8257_ & new_F8256_;
  assign new_F8244_ = new_F8255_ & new_F8254_;
  assign new_F8245_ = new_F8260_ | new_F8259_;
  assign new_F8246_ = new_F8255_ & new_F8258_;
  assign new_F8247_ = F8230 | new_F8263_;
  assign new_F8248_ = new_F8262_ | new_F8261_;
  assign new_F8249_ = new_F8265_ | new_F8264_;
  assign new_F8250_ = ~new_F8241_ & new_F8267_;
  assign new_F8251_ = ~new_F8243_ & new_F8255_;
  assign new_F8252_ = new_F8243_ & ~new_F8255_;
  assign new_F8253_ = F8229 & ~F8230;
  assign new_F8254_ = ~new_F8276_ | ~new_F8277_;
  assign new_F8255_ = new_F8269_ | new_F8271_;
  assign new_F8256_ = new_F8279_ | new_F8278_;
  assign new_F8257_ = new_F8273_ | new_F8272_;
  assign new_F8258_ = ~new_F8281_ | ~new_F8280_;
  assign new_F8259_ = ~new_F8282_ & new_F8283_;
  assign new_F8260_ = new_F8282_ & ~new_F8283_;
  assign new_F8261_ = ~F8229 & F8230;
  assign new_F8262_ = F8229 & ~F8230;
  assign new_F8263_ = ~new_F8245_ | new_F8255_;
  assign new_F8264_ = new_F8245_ & new_F8255_;
  assign new_F8265_ = ~new_F8245_ & ~new_F8255_;
  assign new_F8266_ = new_F8287_ | new_F8286_;
  assign new_F8267_ = F8233 | new_F8266_;
  assign new_F8268_ = new_F8291_ | new_F8290_;
  assign new_F8269_ = ~F8233 & new_F8268_;
  assign new_F8270_ = new_F8289_ | new_F8288_;
  assign new_F8271_ = F8233 & new_F8270_;
  assign new_F8272_ = F8231 & ~new_F8241_;
  assign new_F8273_ = ~F8231 & new_F8241_;
  assign new_F8274_ = ~F8230 | ~new_F8255_;
  assign new_F8275_ = new_F8241_ & new_F8274_;
  assign new_F8276_ = ~new_F8241_ & ~new_F8275_;
  assign new_F8277_ = new_F8241_ | new_F8274_;
  assign new_F8278_ = ~F8231 & F8232;
  assign new_F8279_ = F8231 & ~F8232;
  assign new_F8280_ = new_F8248_ | new_F8285_;
  assign new_F8281_ = ~new_F8248_ & ~new_F8284_;
  assign new_F8282_ = F8231 | new_F8248_;
  assign new_F8283_ = F8231 | F8232;
  assign new_F8284_ = new_F8248_ & new_F8285_;
  assign new_F8285_ = ~F8230 | ~new_F8255_;
  assign new_F8286_ = new_F8263_ & new_F8283_;
  assign new_F8287_ = ~new_F8263_ & ~new_F8283_;
  assign new_F8288_ = new_F8292_ | new_F8293_;
  assign new_F8289_ = ~F8234 & new_F8248_;
  assign new_F8290_ = new_F8294_ | new_F8295_;
  assign new_F8291_ = F8234 & new_F8248_;
  assign new_F8292_ = ~F8234 & ~new_F8248_;
  assign new_F8293_ = F8234 & ~new_F8248_;
  assign new_F8294_ = F8234 & ~new_F8248_;
  assign new_F8295_ = ~F8234 & new_F8248_;
  assign new_F8302_ = new_F8309_ & new_F8308_;
  assign new_F8303_ = new_F8311_ | new_F8310_;
  assign new_F8304_ = new_F8313_ | new_F8312_;
  assign new_F8305_ = new_F8315_ & new_F8314_;
  assign new_F8306_ = new_F8315_ & new_F8316_;
  assign new_F8307_ = new_F8308_ | new_F8317_;
  assign new_F8308_ = F8297 | new_F8320_;
  assign new_F8309_ = new_F8319_ | new_F8318_;
  assign new_F8310_ = new_F8324_ & new_F8323_;
  assign new_F8311_ = new_F8322_ & new_F8321_;
  assign new_F8312_ = new_F8327_ | new_F8326_;
  assign new_F8313_ = new_F8322_ & new_F8325_;
  assign new_F8314_ = F8297 | new_F8330_;
  assign new_F8315_ = new_F8329_ | new_F8328_;
  assign new_F8316_ = new_F8332_ | new_F8331_;
  assign new_F8317_ = ~new_F8308_ & new_F8334_;
  assign new_F8318_ = ~new_F8310_ & new_F8322_;
  assign new_F8319_ = new_F8310_ & ~new_F8322_;
  assign new_F8320_ = F8296 & ~F8297;
  assign new_F8321_ = ~new_F8343_ | ~new_F8344_;
  assign new_F8322_ = new_F8336_ | new_F8338_;
  assign new_F8323_ = new_F8346_ | new_F8345_;
  assign new_F8324_ = new_F8340_ | new_F8339_;
  assign new_F8325_ = ~new_F8348_ | ~new_F8347_;
  assign new_F8326_ = ~new_F8349_ & new_F8350_;
  assign new_F8327_ = new_F8349_ & ~new_F8350_;
  assign new_F8328_ = ~F8296 & F8297;
  assign new_F8329_ = F8296 & ~F8297;
  assign new_F8330_ = ~new_F8312_ | new_F8322_;
  assign new_F8331_ = new_F8312_ & new_F8322_;
  assign new_F8332_ = ~new_F8312_ & ~new_F8322_;
  assign new_F8333_ = new_F8354_ | new_F8353_;
  assign new_F8334_ = F8300 | new_F8333_;
  assign new_F8335_ = new_F8358_ | new_F8357_;
  assign new_F8336_ = ~F8300 & new_F8335_;
  assign new_F8337_ = new_F8356_ | new_F8355_;
  assign new_F8338_ = F8300 & new_F8337_;
  assign new_F8339_ = F8298 & ~new_F8308_;
  assign new_F8340_ = ~F8298 & new_F8308_;
  assign new_F8341_ = ~F8297 | ~new_F8322_;
  assign new_F8342_ = new_F8308_ & new_F8341_;
  assign new_F8343_ = ~new_F8308_ & ~new_F8342_;
  assign new_F8344_ = new_F8308_ | new_F8341_;
  assign new_F8345_ = ~F8298 & F8299;
  assign new_F8346_ = F8298 & ~F8299;
  assign new_F8347_ = new_F8315_ | new_F8352_;
  assign new_F8348_ = ~new_F8315_ & ~new_F8351_;
  assign new_F8349_ = F8298 | new_F8315_;
  assign new_F8350_ = F8298 | F8299;
  assign new_F8351_ = new_F8315_ & new_F8352_;
  assign new_F8352_ = ~F8297 | ~new_F8322_;
  assign new_F8353_ = new_F8330_ & new_F8350_;
  assign new_F8354_ = ~new_F8330_ & ~new_F8350_;
  assign new_F8355_ = new_F8359_ | new_F8360_;
  assign new_F8356_ = ~F8301 & new_F8315_;
  assign new_F8357_ = new_F8361_ | new_F8362_;
  assign new_F8358_ = F8301 & new_F8315_;
  assign new_F8359_ = ~F8301 & ~new_F8315_;
  assign new_F8360_ = F8301 & ~new_F8315_;
  assign new_F8361_ = F8301 & ~new_F8315_;
  assign new_F8362_ = ~F8301 & new_F8315_;
  assign new_F8369_ = new_F8376_ & new_F8375_;
  assign new_F8370_ = new_F8378_ | new_F8377_;
  assign new_F8371_ = new_F8380_ | new_F8379_;
  assign new_F8372_ = new_F8382_ & new_F8381_;
  assign new_F8373_ = new_F8382_ & new_F8383_;
  assign new_F8374_ = new_F8375_ | new_F8384_;
  assign new_F8375_ = F8364 | new_F8387_;
  assign new_F8376_ = new_F8386_ | new_F8385_;
  assign new_F8377_ = new_F8391_ & new_F8390_;
  assign new_F8378_ = new_F8389_ & new_F8388_;
  assign new_F8379_ = new_F8394_ | new_F8393_;
  assign new_F8380_ = new_F8389_ & new_F8392_;
  assign new_F8381_ = F8364 | new_F8397_;
  assign new_F8382_ = new_F8396_ | new_F8395_;
  assign new_F8383_ = new_F8399_ | new_F8398_;
  assign new_F8384_ = ~new_F8375_ & new_F8401_;
  assign new_F8385_ = ~new_F8377_ & new_F8389_;
  assign new_F8386_ = new_F8377_ & ~new_F8389_;
  assign new_F8387_ = F8363 & ~F8364;
  assign new_F8388_ = ~new_F8410_ | ~new_F8411_;
  assign new_F8389_ = new_F8403_ | new_F8405_;
  assign new_F8390_ = new_F8413_ | new_F8412_;
  assign new_F8391_ = new_F8407_ | new_F8406_;
  assign new_F8392_ = ~new_F8415_ | ~new_F8414_;
  assign new_F8393_ = ~new_F8416_ & new_F8417_;
  assign new_F8394_ = new_F8416_ & ~new_F8417_;
  assign new_F8395_ = ~F8363 & F8364;
  assign new_F8396_ = F8363 & ~F8364;
  assign new_F8397_ = ~new_F8379_ | new_F8389_;
  assign new_F8398_ = new_F8379_ & new_F8389_;
  assign new_F8399_ = ~new_F8379_ & ~new_F8389_;
  assign new_F8400_ = new_F8421_ | new_F8420_;
  assign new_F8401_ = F8367 | new_F8400_;
  assign new_F8402_ = new_F8425_ | new_F8424_;
  assign new_F8403_ = ~F8367 & new_F8402_;
  assign new_F8404_ = new_F8423_ | new_F8422_;
  assign new_F8405_ = F8367 & new_F8404_;
  assign new_F8406_ = F8365 & ~new_F8375_;
  assign new_F8407_ = ~F8365 & new_F8375_;
  assign new_F8408_ = ~F8364 | ~new_F8389_;
  assign new_F8409_ = new_F8375_ & new_F8408_;
  assign new_F8410_ = ~new_F8375_ & ~new_F8409_;
  assign new_F8411_ = new_F8375_ | new_F8408_;
  assign new_F8412_ = ~F8365 & F8366;
  assign new_F8413_ = F8365 & ~F8366;
  assign new_F8414_ = new_F8382_ | new_F8419_;
  assign new_F8415_ = ~new_F8382_ & ~new_F8418_;
  assign new_F8416_ = F8365 | new_F8382_;
  assign new_F8417_ = F8365 | F8366;
  assign new_F8418_ = new_F8382_ & new_F8419_;
  assign new_F8419_ = ~F8364 | ~new_F8389_;
  assign new_F8420_ = new_F8397_ & new_F8417_;
  assign new_F8421_ = ~new_F8397_ & ~new_F8417_;
  assign new_F8422_ = new_F8426_ | new_F8427_;
  assign new_F8423_ = ~F8368 & new_F8382_;
  assign new_F8424_ = new_F8428_ | new_F8429_;
  assign new_F8425_ = F8368 & new_F8382_;
  assign new_F8426_ = ~F8368 & ~new_F8382_;
  assign new_F8427_ = F8368 & ~new_F8382_;
  assign new_F8428_ = F8368 & ~new_F8382_;
  assign new_F8429_ = ~F8368 & new_F8382_;
  assign new_F8436_ = new_F8443_ & new_F8442_;
  assign new_F8437_ = new_F8445_ | new_F8444_;
  assign new_F8438_ = new_F8447_ | new_F8446_;
  assign new_F8439_ = new_F8449_ & new_F8448_;
  assign new_F8440_ = new_F8449_ & new_F8450_;
  assign new_F8441_ = new_F8442_ | new_F8451_;
  assign new_F8442_ = F8431 | new_F8454_;
  assign new_F8443_ = new_F8453_ | new_F8452_;
  assign new_F8444_ = new_F8458_ & new_F8457_;
  assign new_F8445_ = new_F8456_ & new_F8455_;
  assign new_F8446_ = new_F8461_ | new_F8460_;
  assign new_F8447_ = new_F8456_ & new_F8459_;
  assign new_F8448_ = F8431 | new_F8464_;
  assign new_F8449_ = new_F8463_ | new_F8462_;
  assign new_F8450_ = new_F8466_ | new_F8465_;
  assign new_F8451_ = ~new_F8442_ & new_F8468_;
  assign new_F8452_ = ~new_F8444_ & new_F8456_;
  assign new_F8453_ = new_F8444_ & ~new_F8456_;
  assign new_F8454_ = F8430 & ~F8431;
  assign new_F8455_ = ~new_F8477_ | ~new_F8478_;
  assign new_F8456_ = new_F8470_ | new_F8472_;
  assign new_F8457_ = new_F8480_ | new_F8479_;
  assign new_F8458_ = new_F8474_ | new_F8473_;
  assign new_F8459_ = ~new_F8482_ | ~new_F8481_;
  assign new_F8460_ = ~new_F8483_ & new_F8484_;
  assign new_F8461_ = new_F8483_ & ~new_F8484_;
  assign new_F8462_ = ~F8430 & F8431;
  assign new_F8463_ = F8430 & ~F8431;
  assign new_F8464_ = ~new_F8446_ | new_F8456_;
  assign new_F8465_ = new_F8446_ & new_F8456_;
  assign new_F8466_ = ~new_F8446_ & ~new_F8456_;
  assign new_F8467_ = new_F8488_ | new_F8487_;
  assign new_F8468_ = F8434 | new_F8467_;
  assign new_F8469_ = new_F8492_ | new_F8491_;
  assign new_F8470_ = ~F8434 & new_F8469_;
  assign new_F8471_ = new_F8490_ | new_F8489_;
  assign new_F8472_ = F8434 & new_F8471_;
  assign new_F8473_ = F8432 & ~new_F8442_;
  assign new_F8474_ = ~F8432 & new_F8442_;
  assign new_F8475_ = ~F8431 | ~new_F8456_;
  assign new_F8476_ = new_F8442_ & new_F8475_;
  assign new_F8477_ = ~new_F8442_ & ~new_F8476_;
  assign new_F8478_ = new_F8442_ | new_F8475_;
  assign new_F8479_ = ~F8432 & F8433;
  assign new_F8480_ = F8432 & ~F8433;
  assign new_F8481_ = new_F8449_ | new_F8486_;
  assign new_F8482_ = ~new_F8449_ & ~new_F8485_;
  assign new_F8483_ = F8432 | new_F8449_;
  assign new_F8484_ = F8432 | F8433;
  assign new_F8485_ = new_F8449_ & new_F8486_;
  assign new_F8486_ = ~F8431 | ~new_F8456_;
  assign new_F8487_ = new_F8464_ & new_F8484_;
  assign new_F8488_ = ~new_F8464_ & ~new_F8484_;
  assign new_F8489_ = new_F8493_ | new_F8494_;
  assign new_F8490_ = ~F8435 & new_F8449_;
  assign new_F8491_ = new_F8495_ | new_F8496_;
  assign new_F8492_ = F8435 & new_F8449_;
  assign new_F8493_ = ~F8435 & ~new_F8449_;
  assign new_F8494_ = F8435 & ~new_F8449_;
  assign new_F8495_ = F8435 & ~new_F8449_;
  assign new_F8496_ = ~F8435 & new_F8449_;
  assign new_F8503_ = new_F8510_ & new_F8509_;
  assign new_F8504_ = new_F8512_ | new_F8511_;
  assign new_F8505_ = new_F8514_ | new_F8513_;
  assign new_F8506_ = new_F8516_ & new_F8515_;
  assign new_F8507_ = new_F8516_ & new_F8517_;
  assign new_F8508_ = new_F8509_ | new_F8518_;
  assign new_F8509_ = F8498 | new_F8521_;
  assign new_F8510_ = new_F8520_ | new_F8519_;
  assign new_F8511_ = new_F8525_ & new_F8524_;
  assign new_F8512_ = new_F8523_ & new_F8522_;
  assign new_F8513_ = new_F8528_ | new_F8527_;
  assign new_F8514_ = new_F8523_ & new_F8526_;
  assign new_F8515_ = F8498 | new_F8531_;
  assign new_F8516_ = new_F8530_ | new_F8529_;
  assign new_F8517_ = new_F8533_ | new_F8532_;
  assign new_F8518_ = ~new_F8509_ & new_F8535_;
  assign new_F8519_ = ~new_F8511_ & new_F8523_;
  assign new_F8520_ = new_F8511_ & ~new_F8523_;
  assign new_F8521_ = F8497 & ~F8498;
  assign new_F8522_ = ~new_F8544_ | ~new_F8545_;
  assign new_F8523_ = new_F8537_ | new_F8539_;
  assign new_F8524_ = new_F8547_ | new_F8546_;
  assign new_F8525_ = new_F8541_ | new_F8540_;
  assign new_F8526_ = ~new_F8549_ | ~new_F8548_;
  assign new_F8527_ = ~new_F8550_ & new_F8551_;
  assign new_F8528_ = new_F8550_ & ~new_F8551_;
  assign new_F8529_ = ~F8497 & F8498;
  assign new_F8530_ = F8497 & ~F8498;
  assign new_F8531_ = ~new_F8513_ | new_F8523_;
  assign new_F8532_ = new_F8513_ & new_F8523_;
  assign new_F8533_ = ~new_F8513_ & ~new_F8523_;
  assign new_F8534_ = new_F8555_ | new_F8554_;
  assign new_F8535_ = F8501 | new_F8534_;
  assign new_F8536_ = new_F8559_ | new_F8558_;
  assign new_F8537_ = ~F8501 & new_F8536_;
  assign new_F8538_ = new_F8557_ | new_F8556_;
  assign new_F8539_ = F8501 & new_F8538_;
  assign new_F8540_ = F8499 & ~new_F8509_;
  assign new_F8541_ = ~F8499 & new_F8509_;
  assign new_F8542_ = ~F8498 | ~new_F8523_;
  assign new_F8543_ = new_F8509_ & new_F8542_;
  assign new_F8544_ = ~new_F8509_ & ~new_F8543_;
  assign new_F8545_ = new_F8509_ | new_F8542_;
  assign new_F8546_ = ~F8499 & F8500;
  assign new_F8547_ = F8499 & ~F8500;
  assign new_F8548_ = new_F8516_ | new_F8553_;
  assign new_F8549_ = ~new_F8516_ & ~new_F8552_;
  assign new_F8550_ = F8499 | new_F8516_;
  assign new_F8551_ = F8499 | F8500;
  assign new_F8552_ = new_F8516_ & new_F8553_;
  assign new_F8553_ = ~F8498 | ~new_F8523_;
  assign new_F8554_ = new_F8531_ & new_F8551_;
  assign new_F8555_ = ~new_F8531_ & ~new_F8551_;
  assign new_F8556_ = new_F8560_ | new_F8561_;
  assign new_F8557_ = ~F8502 & new_F8516_;
  assign new_F8558_ = new_F8562_ | new_F8563_;
  assign new_F8559_ = F8502 & new_F8516_;
  assign new_F8560_ = ~F8502 & ~new_F8516_;
  assign new_F8561_ = F8502 & ~new_F8516_;
  assign new_F8562_ = F8502 & ~new_F8516_;
  assign new_F8563_ = ~F8502 & new_F8516_;
  assign new_F8570_ = new_F8577_ & new_F8576_;
  assign new_F8571_ = new_F8579_ | new_F8578_;
  assign new_F8572_ = new_F8581_ | new_F8580_;
  assign new_F8573_ = new_F8583_ & new_F8582_;
  assign new_F8574_ = new_F8583_ & new_F8584_;
  assign new_F8575_ = new_F8576_ | new_F8585_;
  assign new_F8576_ = F8565 | new_F8588_;
  assign new_F8577_ = new_F8587_ | new_F8586_;
  assign new_F8578_ = new_F8592_ & new_F8591_;
  assign new_F8579_ = new_F8590_ & new_F8589_;
  assign new_F8580_ = new_F8595_ | new_F8594_;
  assign new_F8581_ = new_F8590_ & new_F8593_;
  assign new_F8582_ = F8565 | new_F8598_;
  assign new_F8583_ = new_F8597_ | new_F8596_;
  assign new_F8584_ = new_F8600_ | new_F8599_;
  assign new_F8585_ = ~new_F8576_ & new_F8602_;
  assign new_F8586_ = ~new_F8578_ & new_F8590_;
  assign new_F8587_ = new_F8578_ & ~new_F8590_;
  assign new_F8588_ = F8564 & ~F8565;
  assign new_F8589_ = ~new_F8611_ | ~new_F8612_;
  assign new_F8590_ = new_F8604_ | new_F8606_;
  assign new_F8591_ = new_F8614_ | new_F8613_;
  assign new_F8592_ = new_F8608_ | new_F8607_;
  assign new_F8593_ = ~new_F8616_ | ~new_F8615_;
  assign new_F8594_ = ~new_F8617_ & new_F8618_;
  assign new_F8595_ = new_F8617_ & ~new_F8618_;
  assign new_F8596_ = ~F8564 & F8565;
  assign new_F8597_ = F8564 & ~F8565;
  assign new_F8598_ = ~new_F8580_ | new_F8590_;
  assign new_F8599_ = new_F8580_ & new_F8590_;
  assign new_F8600_ = ~new_F8580_ & ~new_F8590_;
  assign new_F8601_ = new_F8622_ | new_F8621_;
  assign new_F8602_ = F8568 | new_F8601_;
  assign new_F8603_ = new_F8626_ | new_F8625_;
  assign new_F8604_ = ~F8568 & new_F8603_;
  assign new_F8605_ = new_F8624_ | new_F8623_;
  assign new_F8606_ = F8568 & new_F8605_;
  assign new_F8607_ = F8566 & ~new_F8576_;
  assign new_F8608_ = ~F8566 & new_F8576_;
  assign new_F8609_ = ~F8565 | ~new_F8590_;
  assign new_F8610_ = new_F8576_ & new_F8609_;
  assign new_F8611_ = ~new_F8576_ & ~new_F8610_;
  assign new_F8612_ = new_F8576_ | new_F8609_;
  assign new_F8613_ = ~F8566 & F8567;
  assign new_F8614_ = F8566 & ~F8567;
  assign new_F8615_ = new_F8583_ | new_F8620_;
  assign new_F8616_ = ~new_F8583_ & ~new_F8619_;
  assign new_F8617_ = F8566 | new_F8583_;
  assign new_F8618_ = F8566 | F8567;
  assign new_F8619_ = new_F8583_ & new_F8620_;
  assign new_F8620_ = ~F8565 | ~new_F8590_;
  assign new_F8621_ = new_F8598_ & new_F8618_;
  assign new_F8622_ = ~new_F8598_ & ~new_F8618_;
  assign new_F8623_ = new_F8627_ | new_F8628_;
  assign new_F8624_ = ~F8569 & new_F8583_;
  assign new_F8625_ = new_F8629_ | new_F8630_;
  assign new_F8626_ = F8569 & new_F8583_;
  assign new_F8627_ = ~F8569 & ~new_F8583_;
  assign new_F8628_ = F8569 & ~new_F8583_;
  assign new_F8629_ = F8569 & ~new_F8583_;
  assign new_F8630_ = ~F8569 & new_F8583_;
  assign new_F8637_ = new_F8644_ & new_F8643_;
  assign new_F8638_ = new_F8646_ | new_F8645_;
  assign new_F8639_ = new_F8648_ | new_F8647_;
  assign new_F8640_ = new_F8650_ & new_F8649_;
  assign new_F8641_ = new_F8650_ & new_F8651_;
  assign new_F8642_ = new_F8643_ | new_F8652_;
  assign new_F8643_ = F8632 | new_F8655_;
  assign new_F8644_ = new_F8654_ | new_F8653_;
  assign new_F8645_ = new_F8659_ & new_F8658_;
  assign new_F8646_ = new_F8657_ & new_F8656_;
  assign new_F8647_ = new_F8662_ | new_F8661_;
  assign new_F8648_ = new_F8657_ & new_F8660_;
  assign new_F8649_ = F8632 | new_F8665_;
  assign new_F8650_ = new_F8664_ | new_F8663_;
  assign new_F8651_ = new_F8667_ | new_F8666_;
  assign new_F8652_ = ~new_F8643_ & new_F8669_;
  assign new_F8653_ = ~new_F8645_ & new_F8657_;
  assign new_F8654_ = new_F8645_ & ~new_F8657_;
  assign new_F8655_ = F8631 & ~F8632;
  assign new_F8656_ = ~new_F8678_ | ~new_F8679_;
  assign new_F8657_ = new_F8671_ | new_F8673_;
  assign new_F8658_ = new_F8681_ | new_F8680_;
  assign new_F8659_ = new_F8675_ | new_F8674_;
  assign new_F8660_ = ~new_F8683_ | ~new_F8682_;
  assign new_F8661_ = ~new_F8684_ & new_F8685_;
  assign new_F8662_ = new_F8684_ & ~new_F8685_;
  assign new_F8663_ = ~F8631 & F8632;
  assign new_F8664_ = F8631 & ~F8632;
  assign new_F8665_ = ~new_F8647_ | new_F8657_;
  assign new_F8666_ = new_F8647_ & new_F8657_;
  assign new_F8667_ = ~new_F8647_ & ~new_F8657_;
  assign new_F8668_ = new_F8689_ | new_F8688_;
  assign new_F8669_ = F8635 | new_F8668_;
  assign new_F8670_ = new_F8693_ | new_F8692_;
  assign new_F8671_ = ~F8635 & new_F8670_;
  assign new_F8672_ = new_F8691_ | new_F8690_;
  assign new_F8673_ = F8635 & new_F8672_;
  assign new_F8674_ = F8633 & ~new_F8643_;
  assign new_F8675_ = ~F8633 & new_F8643_;
  assign new_F8676_ = ~F8632 | ~new_F8657_;
  assign new_F8677_ = new_F8643_ & new_F8676_;
  assign new_F8678_ = ~new_F8643_ & ~new_F8677_;
  assign new_F8679_ = new_F8643_ | new_F8676_;
  assign new_F8680_ = ~F8633 & F8634;
  assign new_F8681_ = F8633 & ~F8634;
  assign new_F8682_ = new_F8650_ | new_F8687_;
  assign new_F8683_ = ~new_F8650_ & ~new_F8686_;
  assign new_F8684_ = F8633 | new_F8650_;
  assign new_F8685_ = F8633 | F8634;
  assign new_F8686_ = new_F8650_ & new_F8687_;
  assign new_F8687_ = ~F8632 | ~new_F8657_;
  assign new_F8688_ = new_F8665_ & new_F8685_;
  assign new_F8689_ = ~new_F8665_ & ~new_F8685_;
  assign new_F8690_ = new_F8694_ | new_F8695_;
  assign new_F8691_ = ~F8636 & new_F8650_;
  assign new_F8692_ = new_F8696_ | new_F8697_;
  assign new_F8693_ = F8636 & new_F8650_;
  assign new_F8694_ = ~F8636 & ~new_F8650_;
  assign new_F8695_ = F8636 & ~new_F8650_;
  assign new_F8696_ = F8636 & ~new_F8650_;
  assign new_F8697_ = ~F8636 & new_F8650_;
  assign new_F8704_ = new_F8711_ & new_F8710_;
  assign new_F8705_ = new_F8713_ | new_F8712_;
  assign new_F8706_ = new_F8715_ | new_F8714_;
  assign new_F8707_ = new_F8717_ & new_F8716_;
  assign new_F8708_ = new_F8717_ & new_F8718_;
  assign new_F8709_ = new_F8710_ | new_F8719_;
  assign new_F8710_ = F8699 | new_F8722_;
  assign new_F8711_ = new_F8721_ | new_F8720_;
  assign new_F8712_ = new_F8726_ & new_F8725_;
  assign new_F8713_ = new_F8724_ & new_F8723_;
  assign new_F8714_ = new_F8729_ | new_F8728_;
  assign new_F8715_ = new_F8724_ & new_F8727_;
  assign new_F8716_ = F8699 | new_F8732_;
  assign new_F8717_ = new_F8731_ | new_F8730_;
  assign new_F8718_ = new_F8734_ | new_F8733_;
  assign new_F8719_ = ~new_F8710_ & new_F8736_;
  assign new_F8720_ = ~new_F8712_ & new_F8724_;
  assign new_F8721_ = new_F8712_ & ~new_F8724_;
  assign new_F8722_ = F8698 & ~F8699;
  assign new_F8723_ = ~new_F8745_ | ~new_F8746_;
  assign new_F8724_ = new_F8738_ | new_F8740_;
  assign new_F8725_ = new_F8748_ | new_F8747_;
  assign new_F8726_ = new_F8742_ | new_F8741_;
  assign new_F8727_ = ~new_F8750_ | ~new_F8749_;
  assign new_F8728_ = ~new_F8751_ & new_F8752_;
  assign new_F8729_ = new_F8751_ & ~new_F8752_;
  assign new_F8730_ = ~F8698 & F8699;
  assign new_F8731_ = F8698 & ~F8699;
  assign new_F8732_ = ~new_F8714_ | new_F8724_;
  assign new_F8733_ = new_F8714_ & new_F8724_;
  assign new_F8734_ = ~new_F8714_ & ~new_F8724_;
  assign new_F8735_ = new_F8756_ | new_F8755_;
  assign new_F8736_ = F8702 | new_F8735_;
  assign new_F8737_ = new_F8760_ | new_F8759_;
  assign new_F8738_ = ~F8702 & new_F8737_;
  assign new_F8739_ = new_F8758_ | new_F8757_;
  assign new_F8740_ = F8702 & new_F8739_;
  assign new_F8741_ = F8700 & ~new_F8710_;
  assign new_F8742_ = ~F8700 & new_F8710_;
  assign new_F8743_ = ~F8699 | ~new_F8724_;
  assign new_F8744_ = new_F8710_ & new_F8743_;
  assign new_F8745_ = ~new_F8710_ & ~new_F8744_;
  assign new_F8746_ = new_F8710_ | new_F8743_;
  assign new_F8747_ = ~F8700 & F8701;
  assign new_F8748_ = F8700 & ~F8701;
  assign new_F8749_ = new_F8717_ | new_F8754_;
  assign new_F8750_ = ~new_F8717_ & ~new_F8753_;
  assign new_F8751_ = F8700 | new_F8717_;
  assign new_F8752_ = F8700 | F8701;
  assign new_F8753_ = new_F8717_ & new_F8754_;
  assign new_F8754_ = ~F8699 | ~new_F8724_;
  assign new_F8755_ = new_F8732_ & new_F8752_;
  assign new_F8756_ = ~new_F8732_ & ~new_F8752_;
  assign new_F8757_ = new_F8761_ | new_F8762_;
  assign new_F8758_ = ~F8703 & new_F8717_;
  assign new_F8759_ = new_F8763_ | new_F8764_;
  assign new_F8760_ = F8703 & new_F8717_;
  assign new_F8761_ = ~F8703 & ~new_F8717_;
  assign new_F8762_ = F8703 & ~new_F8717_;
  assign new_F8763_ = F8703 & ~new_F8717_;
  assign new_F8764_ = ~F8703 & new_F8717_;
  assign new_F8771_ = new_F8778_ & new_F8777_;
  assign new_F8772_ = new_F8780_ | new_F8779_;
  assign new_F8773_ = new_F8782_ | new_F8781_;
  assign new_F8774_ = new_F8784_ & new_F8783_;
  assign new_F8775_ = new_F8784_ & new_F8785_;
  assign new_F8776_ = new_F8777_ | new_F8786_;
  assign new_F8777_ = F8766 | new_F8789_;
  assign new_F8778_ = new_F8788_ | new_F8787_;
  assign new_F8779_ = new_F8793_ & new_F8792_;
  assign new_F8780_ = new_F8791_ & new_F8790_;
  assign new_F8781_ = new_F8796_ | new_F8795_;
  assign new_F8782_ = new_F8791_ & new_F8794_;
  assign new_F8783_ = F8766 | new_F8799_;
  assign new_F8784_ = new_F8798_ | new_F8797_;
  assign new_F8785_ = new_F8801_ | new_F8800_;
  assign new_F8786_ = ~new_F8777_ & new_F8803_;
  assign new_F8787_ = ~new_F8779_ & new_F8791_;
  assign new_F8788_ = new_F8779_ & ~new_F8791_;
  assign new_F8789_ = F8765 & ~F8766;
  assign new_F8790_ = ~new_F8812_ | ~new_F8813_;
  assign new_F8791_ = new_F8805_ | new_F8807_;
  assign new_F8792_ = new_F8815_ | new_F8814_;
  assign new_F8793_ = new_F8809_ | new_F8808_;
  assign new_F8794_ = ~new_F8817_ | ~new_F8816_;
  assign new_F8795_ = ~new_F8818_ & new_F8819_;
  assign new_F8796_ = new_F8818_ & ~new_F8819_;
  assign new_F8797_ = ~F8765 & F8766;
  assign new_F8798_ = F8765 & ~F8766;
  assign new_F8799_ = ~new_F8781_ | new_F8791_;
  assign new_F8800_ = new_F8781_ & new_F8791_;
  assign new_F8801_ = ~new_F8781_ & ~new_F8791_;
  assign new_F8802_ = new_F8823_ | new_F8822_;
  assign new_F8803_ = F8769 | new_F8802_;
  assign new_F8804_ = new_F8827_ | new_F8826_;
  assign new_F8805_ = ~F8769 & new_F8804_;
  assign new_F8806_ = new_F8825_ | new_F8824_;
  assign new_F8807_ = F8769 & new_F8806_;
  assign new_F8808_ = F8767 & ~new_F8777_;
  assign new_F8809_ = ~F8767 & new_F8777_;
  assign new_F8810_ = ~F8766 | ~new_F8791_;
  assign new_F8811_ = new_F8777_ & new_F8810_;
  assign new_F8812_ = ~new_F8777_ & ~new_F8811_;
  assign new_F8813_ = new_F8777_ | new_F8810_;
  assign new_F8814_ = ~F8767 & F8768;
  assign new_F8815_ = F8767 & ~F8768;
  assign new_F8816_ = new_F8784_ | new_F8821_;
  assign new_F8817_ = ~new_F8784_ & ~new_F8820_;
  assign new_F8818_ = F8767 | new_F8784_;
  assign new_F8819_ = F8767 | F8768;
  assign new_F8820_ = new_F8784_ & new_F8821_;
  assign new_F8821_ = ~F8766 | ~new_F8791_;
  assign new_F8822_ = new_F8799_ & new_F8819_;
  assign new_F8823_ = ~new_F8799_ & ~new_F8819_;
  assign new_F8824_ = new_F8828_ | new_F8829_;
  assign new_F8825_ = ~F8770 & new_F8784_;
  assign new_F8826_ = new_F8830_ | new_F8831_;
  assign new_F8827_ = F8770 & new_F8784_;
  assign new_F8828_ = ~F8770 & ~new_F8784_;
  assign new_F8829_ = F8770 & ~new_F8784_;
  assign new_F8830_ = F8770 & ~new_F8784_;
  assign new_F8831_ = ~F8770 & new_F8784_;
  assign new_F8838_ = new_F8845_ & new_F8844_;
  assign new_F8839_ = new_F8847_ | new_F8846_;
  assign new_F8840_ = new_F8849_ | new_F8848_;
  assign new_F8841_ = new_F8851_ & new_F8850_;
  assign new_F8842_ = new_F8851_ & new_F8852_;
  assign new_F8843_ = new_F8844_ | new_F8853_;
  assign new_F8844_ = F8833 | new_F8856_;
  assign new_F8845_ = new_F8855_ | new_F8854_;
  assign new_F8846_ = new_F8860_ & new_F8859_;
  assign new_F8847_ = new_F8858_ & new_F8857_;
  assign new_F8848_ = new_F8863_ | new_F8862_;
  assign new_F8849_ = new_F8858_ & new_F8861_;
  assign new_F8850_ = F8833 | new_F8866_;
  assign new_F8851_ = new_F8865_ | new_F8864_;
  assign new_F8852_ = new_F8868_ | new_F8867_;
  assign new_F8853_ = ~new_F8844_ & new_F8870_;
  assign new_F8854_ = ~new_F8846_ & new_F8858_;
  assign new_F8855_ = new_F8846_ & ~new_F8858_;
  assign new_F8856_ = F8832 & ~F8833;
  assign new_F8857_ = ~new_F8879_ | ~new_F8880_;
  assign new_F8858_ = new_F8872_ | new_F8874_;
  assign new_F8859_ = new_F8882_ | new_F8881_;
  assign new_F8860_ = new_F8876_ | new_F8875_;
  assign new_F8861_ = ~new_F8884_ | ~new_F8883_;
  assign new_F8862_ = ~new_F8885_ & new_F8886_;
  assign new_F8863_ = new_F8885_ & ~new_F8886_;
  assign new_F8864_ = ~F8832 & F8833;
  assign new_F8865_ = F8832 & ~F8833;
  assign new_F8866_ = ~new_F8848_ | new_F8858_;
  assign new_F8867_ = new_F8848_ & new_F8858_;
  assign new_F8868_ = ~new_F8848_ & ~new_F8858_;
  assign new_F8869_ = new_F8890_ | new_F8889_;
  assign new_F8870_ = F8836 | new_F8869_;
  assign new_F8871_ = new_F8894_ | new_F8893_;
  assign new_F8872_ = ~F8836 & new_F8871_;
  assign new_F8873_ = new_F8892_ | new_F8891_;
  assign new_F8874_ = F8836 & new_F8873_;
  assign new_F8875_ = F8834 & ~new_F8844_;
  assign new_F8876_ = ~F8834 & new_F8844_;
  assign new_F8877_ = ~F8833 | ~new_F8858_;
  assign new_F8878_ = new_F8844_ & new_F8877_;
  assign new_F8879_ = ~new_F8844_ & ~new_F8878_;
  assign new_F8880_ = new_F8844_ | new_F8877_;
  assign new_F8881_ = ~F8834 & F8835;
  assign new_F8882_ = F8834 & ~F8835;
  assign new_F8883_ = new_F8851_ | new_F8888_;
  assign new_F8884_ = ~new_F8851_ & ~new_F8887_;
  assign new_F8885_ = F8834 | new_F8851_;
  assign new_F8886_ = F8834 | F8835;
  assign new_F8887_ = new_F8851_ & new_F8888_;
  assign new_F8888_ = ~F8833 | ~new_F8858_;
  assign new_F8889_ = new_F8866_ & new_F8886_;
  assign new_F8890_ = ~new_F8866_ & ~new_F8886_;
  assign new_F8891_ = new_F8895_ | new_F8896_;
  assign new_F8892_ = ~F8837 & new_F8851_;
  assign new_F8893_ = new_F8897_ | new_F8898_;
  assign new_F8894_ = F8837 & new_F8851_;
  assign new_F8895_ = ~F8837 & ~new_F8851_;
  assign new_F8896_ = F8837 & ~new_F8851_;
  assign new_F8897_ = F8837 & ~new_F8851_;
  assign new_F8898_ = ~F8837 & new_F8851_;
  assign new_F8905_ = new_F8912_ & new_F8911_;
  assign new_F8906_ = new_F8914_ | new_F8913_;
  assign new_F8907_ = new_F8916_ | new_F8915_;
  assign new_F8908_ = new_F8918_ & new_F8917_;
  assign new_F8909_ = new_F8918_ & new_F8919_;
  assign new_F8910_ = new_F8911_ | new_F8920_;
  assign new_F8911_ = F8900 | new_F8923_;
  assign new_F8912_ = new_F8922_ | new_F8921_;
  assign new_F8913_ = new_F8927_ & new_F8926_;
  assign new_F8914_ = new_F8925_ & new_F8924_;
  assign new_F8915_ = new_F8930_ | new_F8929_;
  assign new_F8916_ = new_F8925_ & new_F8928_;
  assign new_F8917_ = F8900 | new_F8933_;
  assign new_F8918_ = new_F8932_ | new_F8931_;
  assign new_F8919_ = new_F8935_ | new_F8934_;
  assign new_F8920_ = ~new_F8911_ & new_F8937_;
  assign new_F8921_ = ~new_F8913_ & new_F8925_;
  assign new_F8922_ = new_F8913_ & ~new_F8925_;
  assign new_F8923_ = F8899 & ~F8900;
  assign new_F8924_ = ~new_F8946_ | ~new_F8947_;
  assign new_F8925_ = new_F8939_ | new_F8941_;
  assign new_F8926_ = new_F8949_ | new_F8948_;
  assign new_F8927_ = new_F8943_ | new_F8942_;
  assign new_F8928_ = ~new_F8951_ | ~new_F8950_;
  assign new_F8929_ = ~new_F8952_ & new_F8953_;
  assign new_F8930_ = new_F8952_ & ~new_F8953_;
  assign new_F8931_ = ~F8899 & F8900;
  assign new_F8932_ = F8899 & ~F8900;
  assign new_F8933_ = ~new_F8915_ | new_F8925_;
  assign new_F8934_ = new_F8915_ & new_F8925_;
  assign new_F8935_ = ~new_F8915_ & ~new_F8925_;
  assign new_F8936_ = new_F8957_ | new_F8956_;
  assign new_F8937_ = F8903 | new_F8936_;
  assign new_F8938_ = new_F8961_ | new_F8960_;
  assign new_F8939_ = ~F8903 & new_F8938_;
  assign new_F8940_ = new_F8959_ | new_F8958_;
  assign new_F8941_ = F8903 & new_F8940_;
  assign new_F8942_ = F8901 & ~new_F8911_;
  assign new_F8943_ = ~F8901 & new_F8911_;
  assign new_F8944_ = ~F8900 | ~new_F8925_;
  assign new_F8945_ = new_F8911_ & new_F8944_;
  assign new_F8946_ = ~new_F8911_ & ~new_F8945_;
  assign new_F8947_ = new_F8911_ | new_F8944_;
  assign new_F8948_ = ~F8901 & F8902;
  assign new_F8949_ = F8901 & ~F8902;
  assign new_F8950_ = new_F8918_ | new_F8955_;
  assign new_F8951_ = ~new_F8918_ & ~new_F8954_;
  assign new_F8952_ = F8901 | new_F8918_;
  assign new_F8953_ = F8901 | F8902;
  assign new_F8954_ = new_F8918_ & new_F8955_;
  assign new_F8955_ = ~F8900 | ~new_F8925_;
  assign new_F8956_ = new_F8933_ & new_F8953_;
  assign new_F8957_ = ~new_F8933_ & ~new_F8953_;
  assign new_F8958_ = new_F8962_ | new_F8963_;
  assign new_F8959_ = ~F8904 & new_F8918_;
  assign new_F8960_ = new_F8964_ | new_F8965_;
  assign new_F8961_ = F8904 & new_F8918_;
  assign new_F8962_ = ~F8904 & ~new_F8918_;
  assign new_F8963_ = F8904 & ~new_F8918_;
  assign new_F8964_ = F8904 & ~new_F8918_;
  assign new_F8965_ = ~F8904 & new_F8918_;
  assign new_F8972_ = new_F8979_ & new_F8978_;
  assign new_F8973_ = new_F8981_ | new_F8980_;
  assign new_F8974_ = new_F8983_ | new_F8982_;
  assign new_F8975_ = new_F8985_ & new_F8984_;
  assign new_F8976_ = new_F8985_ & new_F8986_;
  assign new_F8977_ = new_F8978_ | new_F8987_;
  assign new_F8978_ = F8967 | new_F8990_;
  assign new_F8979_ = new_F8989_ | new_F8988_;
  assign new_F8980_ = new_F8994_ & new_F8993_;
  assign new_F8981_ = new_F8992_ & new_F8991_;
  assign new_F8982_ = new_F8997_ | new_F8996_;
  assign new_F8983_ = new_F8992_ & new_F8995_;
  assign new_F8984_ = F8967 | new_F9000_;
  assign new_F8985_ = new_F8999_ | new_F8998_;
  assign new_F8986_ = new_F9002_ | new_F9001_;
  assign new_F8987_ = ~new_F8978_ & new_F9004_;
  assign new_F8988_ = ~new_F8980_ & new_F8992_;
  assign new_F8989_ = new_F8980_ & ~new_F8992_;
  assign new_F8990_ = F8966 & ~F8967;
  assign new_F8991_ = ~new_F9013_ | ~new_F9014_;
  assign new_F8992_ = new_F9006_ | new_F9008_;
  assign new_F8993_ = new_F9016_ | new_F9015_;
  assign new_F8994_ = new_F9010_ | new_F9009_;
  assign new_F8995_ = ~new_F9018_ | ~new_F9017_;
  assign new_F8996_ = ~new_F9019_ & new_F9020_;
  assign new_F8997_ = new_F9019_ & ~new_F9020_;
  assign new_F8998_ = ~F8966 & F8967;
  assign new_F8999_ = F8966 & ~F8967;
  assign new_F9000_ = ~new_F8982_ | new_F8992_;
  assign new_F9001_ = new_F8982_ & new_F8992_;
  assign new_F9002_ = ~new_F8982_ & ~new_F8992_;
  assign new_F9003_ = new_F9024_ | new_F9023_;
  assign new_F9004_ = F8970 | new_F9003_;
  assign new_F9005_ = new_F9028_ | new_F9027_;
  assign new_F9006_ = ~F8970 & new_F9005_;
  assign new_F9007_ = new_F9026_ | new_F9025_;
  assign new_F9008_ = F8970 & new_F9007_;
  assign new_F9009_ = F8968 & ~new_F8978_;
  assign new_F9010_ = ~F8968 & new_F8978_;
  assign new_F9011_ = ~F8967 | ~new_F8992_;
  assign new_F9012_ = new_F8978_ & new_F9011_;
  assign new_F9013_ = ~new_F8978_ & ~new_F9012_;
  assign new_F9014_ = new_F8978_ | new_F9011_;
  assign new_F9015_ = ~F8968 & F8969;
  assign new_F9016_ = F8968 & ~F8969;
  assign new_F9017_ = new_F8985_ | new_F9022_;
  assign new_F9018_ = ~new_F8985_ & ~new_F9021_;
  assign new_F9019_ = F8968 | new_F8985_;
  assign new_F9020_ = F8968 | F8969;
  assign new_F9021_ = new_F8985_ & new_F9022_;
  assign new_F9022_ = ~F8967 | ~new_F8992_;
  assign new_F9023_ = new_F9000_ & new_F9020_;
  assign new_F9024_ = ~new_F9000_ & ~new_F9020_;
  assign new_F9025_ = new_F9029_ | new_F9030_;
  assign new_F9026_ = ~F8971 & new_F8985_;
  assign new_F9027_ = new_F9031_ | new_F9032_;
  assign new_F9028_ = F8971 & new_F8985_;
  assign new_F9029_ = ~F8971 & ~new_F8985_;
  assign new_F9030_ = F8971 & ~new_F8985_;
  assign new_F9031_ = F8971 & ~new_F8985_;
  assign new_F9032_ = ~F8971 & new_F8985_;
  assign new_F9039_ = new_F9046_ & new_F9045_;
  assign new_F9040_ = new_F9048_ | new_F9047_;
  assign new_F9041_ = new_F9050_ | new_F9049_;
  assign new_F9042_ = new_F9052_ & new_F9051_;
  assign new_F9043_ = new_F9052_ & new_F9053_;
  assign new_F9044_ = new_F9045_ | new_F9054_;
  assign new_F9045_ = F9034 | new_F9057_;
  assign new_F9046_ = new_F9056_ | new_F9055_;
  assign new_F9047_ = new_F9061_ & new_F9060_;
  assign new_F9048_ = new_F9059_ & new_F9058_;
  assign new_F9049_ = new_F9064_ | new_F9063_;
  assign new_F9050_ = new_F9059_ & new_F9062_;
  assign new_F9051_ = F9034 | new_F9067_;
  assign new_F9052_ = new_F9066_ | new_F9065_;
  assign new_F9053_ = new_F9069_ | new_F9068_;
  assign new_F9054_ = ~new_F9045_ & new_F9071_;
  assign new_F9055_ = ~new_F9047_ & new_F9059_;
  assign new_F9056_ = new_F9047_ & ~new_F9059_;
  assign new_F9057_ = F9033 & ~F9034;
  assign new_F9058_ = ~new_F9080_ | ~new_F9081_;
  assign new_F9059_ = new_F9073_ | new_F9075_;
  assign new_F9060_ = new_F9083_ | new_F9082_;
  assign new_F9061_ = new_F9077_ | new_F9076_;
  assign new_F9062_ = ~new_F9085_ | ~new_F9084_;
  assign new_F9063_ = ~new_F9086_ & new_F9087_;
  assign new_F9064_ = new_F9086_ & ~new_F9087_;
  assign new_F9065_ = ~F9033 & F9034;
  assign new_F9066_ = F9033 & ~F9034;
  assign new_F9067_ = ~new_F9049_ | new_F9059_;
  assign new_F9068_ = new_F9049_ & new_F9059_;
  assign new_F9069_ = ~new_F9049_ & ~new_F9059_;
  assign new_F9070_ = new_F9091_ | new_F9090_;
  assign new_F9071_ = F9037 | new_F9070_;
  assign new_F9072_ = new_F9095_ | new_F9094_;
  assign new_F9073_ = ~F9037 & new_F9072_;
  assign new_F9074_ = new_F9093_ | new_F9092_;
  assign new_F9075_ = F9037 & new_F9074_;
  assign new_F9076_ = F9035 & ~new_F9045_;
  assign new_F9077_ = ~F9035 & new_F9045_;
  assign new_F9078_ = ~F9034 | ~new_F9059_;
  assign new_F9079_ = new_F9045_ & new_F9078_;
  assign new_F9080_ = ~new_F9045_ & ~new_F9079_;
  assign new_F9081_ = new_F9045_ | new_F9078_;
  assign new_F9082_ = ~F9035 & F9036;
  assign new_F9083_ = F9035 & ~F9036;
  assign new_F9084_ = new_F9052_ | new_F9089_;
  assign new_F9085_ = ~new_F9052_ & ~new_F9088_;
  assign new_F9086_ = F9035 | new_F9052_;
  assign new_F9087_ = F9035 | F9036;
  assign new_F9088_ = new_F9052_ & new_F9089_;
  assign new_F9089_ = ~F9034 | ~new_F9059_;
  assign new_F9090_ = new_F9067_ & new_F9087_;
  assign new_F9091_ = ~new_F9067_ & ~new_F9087_;
  assign new_F9092_ = new_F9096_ | new_F9097_;
  assign new_F9093_ = ~F9038 & new_F9052_;
  assign new_F9094_ = new_F9098_ | new_F9099_;
  assign new_F9095_ = F9038 & new_F9052_;
  assign new_F9096_ = ~F9038 & ~new_F9052_;
  assign new_F9097_ = F9038 & ~new_F9052_;
  assign new_F9098_ = F9038 & ~new_F9052_;
  assign new_F9099_ = ~F9038 & new_F9052_;
  assign new_F9106_ = new_F9113_ & new_F9112_;
  assign new_F9107_ = new_F9115_ | new_F9114_;
  assign new_F9108_ = new_F9117_ | new_F9116_;
  assign new_F9109_ = new_F9119_ & new_F9118_;
  assign new_F9110_ = new_F9119_ & new_F9120_;
  assign new_F9111_ = new_F9112_ | new_F9121_;
  assign new_F9112_ = F9101 | new_F9124_;
  assign new_F9113_ = new_F9123_ | new_F9122_;
  assign new_F9114_ = new_F9128_ & new_F9127_;
  assign new_F9115_ = new_F9126_ & new_F9125_;
  assign new_F9116_ = new_F9131_ | new_F9130_;
  assign new_F9117_ = new_F9126_ & new_F9129_;
  assign new_F9118_ = F9101 | new_F9134_;
  assign new_F9119_ = new_F9133_ | new_F9132_;
  assign new_F9120_ = new_F9136_ | new_F9135_;
  assign new_F9121_ = ~new_F9112_ & new_F9138_;
  assign new_F9122_ = ~new_F9114_ & new_F9126_;
  assign new_F9123_ = new_F9114_ & ~new_F9126_;
  assign new_F9124_ = F9100 & ~F9101;
  assign new_F9125_ = ~new_F9147_ | ~new_F9148_;
  assign new_F9126_ = new_F9140_ | new_F9142_;
  assign new_F9127_ = new_F9150_ | new_F9149_;
  assign new_F9128_ = new_F9144_ | new_F9143_;
  assign new_F9129_ = ~new_F9152_ | ~new_F9151_;
  assign new_F9130_ = ~new_F9153_ & new_F9154_;
  assign new_F9131_ = new_F9153_ & ~new_F9154_;
  assign new_F9132_ = ~F9100 & F9101;
  assign new_F9133_ = F9100 & ~F9101;
  assign new_F9134_ = ~new_F9116_ | new_F9126_;
  assign new_F9135_ = new_F9116_ & new_F9126_;
  assign new_F9136_ = ~new_F9116_ & ~new_F9126_;
  assign new_F9137_ = new_F9158_ | new_F9157_;
  assign new_F9138_ = F9104 | new_F9137_;
  assign new_F9139_ = new_F9162_ | new_F9161_;
  assign new_F9140_ = ~F9104 & new_F9139_;
  assign new_F9141_ = new_F9160_ | new_F9159_;
  assign new_F9142_ = F9104 & new_F9141_;
  assign new_F9143_ = F9102 & ~new_F9112_;
  assign new_F9144_ = ~F9102 & new_F9112_;
  assign new_F9145_ = ~F9101 | ~new_F9126_;
  assign new_F9146_ = new_F9112_ & new_F9145_;
  assign new_F9147_ = ~new_F9112_ & ~new_F9146_;
  assign new_F9148_ = new_F9112_ | new_F9145_;
  assign new_F9149_ = ~F9102 & F9103;
  assign new_F9150_ = F9102 & ~F9103;
  assign new_F9151_ = new_F9119_ | new_F9156_;
  assign new_F9152_ = ~new_F9119_ & ~new_F9155_;
  assign new_F9153_ = F9102 | new_F9119_;
  assign new_F9154_ = F9102 | F9103;
  assign new_F9155_ = new_F9119_ & new_F9156_;
  assign new_F9156_ = ~F9101 | ~new_F9126_;
  assign new_F9157_ = new_F9134_ & new_F9154_;
  assign new_F9158_ = ~new_F9134_ & ~new_F9154_;
  assign new_F9159_ = new_F9163_ | new_F9164_;
  assign new_F9160_ = ~F9105 & new_F9119_;
  assign new_F9161_ = new_F9165_ | new_F9166_;
  assign new_F9162_ = F9105 & new_F9119_;
  assign new_F9163_ = ~F9105 & ~new_F9119_;
  assign new_F9164_ = F9105 & ~new_F9119_;
  assign new_F9165_ = F9105 & ~new_F9119_;
  assign new_F9166_ = ~F9105 & new_F9119_;
  assign new_F9173_ = new_F9180_ & new_F9179_;
  assign new_F9174_ = new_F9182_ | new_F9181_;
  assign new_F9175_ = new_F9184_ | new_F9183_;
  assign new_F9176_ = new_F9186_ & new_F9185_;
  assign new_F9177_ = new_F9186_ & new_F9187_;
  assign new_F9178_ = new_F9179_ | new_F9188_;
  assign new_F9179_ = F9168 | new_F9191_;
  assign new_F9180_ = new_F9190_ | new_F9189_;
  assign new_F9181_ = new_F9195_ & new_F9194_;
  assign new_F9182_ = new_F9193_ & new_F9192_;
  assign new_F9183_ = new_F9198_ | new_F9197_;
  assign new_F9184_ = new_F9193_ & new_F9196_;
  assign new_F9185_ = F9168 | new_F9201_;
  assign new_F9186_ = new_F9200_ | new_F9199_;
  assign new_F9187_ = new_F9203_ | new_F9202_;
  assign new_F9188_ = ~new_F9179_ & new_F9205_;
  assign new_F9189_ = ~new_F9181_ & new_F9193_;
  assign new_F9190_ = new_F9181_ & ~new_F9193_;
  assign new_F9191_ = F9167 & ~F9168;
  assign new_F9192_ = ~new_F9214_ | ~new_F9215_;
  assign new_F9193_ = new_F9207_ | new_F9209_;
  assign new_F9194_ = new_F9217_ | new_F9216_;
  assign new_F9195_ = new_F9211_ | new_F9210_;
  assign new_F9196_ = ~new_F9219_ | ~new_F9218_;
  assign new_F9197_ = ~new_F9220_ & new_F9221_;
  assign new_F9198_ = new_F9220_ & ~new_F9221_;
  assign new_F9199_ = ~F9167 & F9168;
  assign new_F9200_ = F9167 & ~F9168;
  assign new_F9201_ = ~new_F9183_ | new_F9193_;
  assign new_F9202_ = new_F9183_ & new_F9193_;
  assign new_F9203_ = ~new_F9183_ & ~new_F9193_;
  assign new_F9204_ = new_F9225_ | new_F9224_;
  assign new_F9205_ = F9171 | new_F9204_;
  assign new_F9206_ = new_F9229_ | new_F9228_;
  assign new_F9207_ = ~F9171 & new_F9206_;
  assign new_F9208_ = new_F9227_ | new_F9226_;
  assign new_F9209_ = F9171 & new_F9208_;
  assign new_F9210_ = F9169 & ~new_F9179_;
  assign new_F9211_ = ~F9169 & new_F9179_;
  assign new_F9212_ = ~F9168 | ~new_F9193_;
  assign new_F9213_ = new_F9179_ & new_F9212_;
  assign new_F9214_ = ~new_F9179_ & ~new_F9213_;
  assign new_F9215_ = new_F9179_ | new_F9212_;
  assign new_F9216_ = ~F9169 & F9170;
  assign new_F9217_ = F9169 & ~F9170;
  assign new_F9218_ = new_F9186_ | new_F9223_;
  assign new_F9219_ = ~new_F9186_ & ~new_F9222_;
  assign new_F9220_ = F9169 | new_F9186_;
  assign new_F9221_ = F9169 | F9170;
  assign new_F9222_ = new_F9186_ & new_F9223_;
  assign new_F9223_ = ~F9168 | ~new_F9193_;
  assign new_F9224_ = new_F9201_ & new_F9221_;
  assign new_F9225_ = ~new_F9201_ & ~new_F9221_;
  assign new_F9226_ = new_F9230_ | new_F9231_;
  assign new_F9227_ = ~F9172 & new_F9186_;
  assign new_F9228_ = new_F9232_ | new_F9233_;
  assign new_F9229_ = F9172 & new_F9186_;
  assign new_F9230_ = ~F9172 & ~new_F9186_;
  assign new_F9231_ = F9172 & ~new_F9186_;
  assign new_F9232_ = F9172 & ~new_F9186_;
  assign new_F9233_ = ~F9172 & new_F9186_;
  assign new_F9240_ = new_F9247_ & new_F9246_;
  assign new_F9241_ = new_F9249_ | new_F9248_;
  assign new_F9242_ = new_F9251_ | new_F9250_;
  assign new_F9243_ = new_F9253_ & new_F9252_;
  assign new_F9244_ = new_F9253_ & new_F9254_;
  assign new_F9245_ = new_F9246_ | new_F9255_;
  assign new_F9246_ = F9235 | new_F9258_;
  assign new_F9247_ = new_F9257_ | new_F9256_;
  assign new_F9248_ = new_F9262_ & new_F9261_;
  assign new_F9249_ = new_F9260_ & new_F9259_;
  assign new_F9250_ = new_F9265_ | new_F9264_;
  assign new_F9251_ = new_F9260_ & new_F9263_;
  assign new_F9252_ = F9235 | new_F9268_;
  assign new_F9253_ = new_F9267_ | new_F9266_;
  assign new_F9254_ = new_F9270_ | new_F9269_;
  assign new_F9255_ = ~new_F9246_ & new_F9272_;
  assign new_F9256_ = ~new_F9248_ & new_F9260_;
  assign new_F9257_ = new_F9248_ & ~new_F9260_;
  assign new_F9258_ = F9234 & ~F9235;
  assign new_F9259_ = ~new_F9281_ | ~new_F9282_;
  assign new_F9260_ = new_F9274_ | new_F9276_;
  assign new_F9261_ = new_F9284_ | new_F9283_;
  assign new_F9262_ = new_F9278_ | new_F9277_;
  assign new_F9263_ = ~new_F9286_ | ~new_F9285_;
  assign new_F9264_ = ~new_F9287_ & new_F9288_;
  assign new_F9265_ = new_F9287_ & ~new_F9288_;
  assign new_F9266_ = ~F9234 & F9235;
  assign new_F9267_ = F9234 & ~F9235;
  assign new_F9268_ = ~new_F9250_ | new_F9260_;
  assign new_F9269_ = new_F9250_ & new_F9260_;
  assign new_F9270_ = ~new_F9250_ & ~new_F9260_;
  assign new_F9271_ = new_F9292_ | new_F9291_;
  assign new_F9272_ = F9238 | new_F9271_;
  assign new_F9273_ = new_F9296_ | new_F9295_;
  assign new_F9274_ = ~F9238 & new_F9273_;
  assign new_F9275_ = new_F9294_ | new_F9293_;
  assign new_F9276_ = F9238 & new_F9275_;
  assign new_F9277_ = F9236 & ~new_F9246_;
  assign new_F9278_ = ~F9236 & new_F9246_;
  assign new_F9279_ = ~F9235 | ~new_F9260_;
  assign new_F9280_ = new_F9246_ & new_F9279_;
  assign new_F9281_ = ~new_F9246_ & ~new_F9280_;
  assign new_F9282_ = new_F9246_ | new_F9279_;
  assign new_F9283_ = ~F9236 & F9237;
  assign new_F9284_ = F9236 & ~F9237;
  assign new_F9285_ = new_F9253_ | new_F9290_;
  assign new_F9286_ = ~new_F9253_ & ~new_F9289_;
  assign new_F9287_ = F9236 | new_F9253_;
  assign new_F9288_ = F9236 | F9237;
  assign new_F9289_ = new_F9253_ & new_F9290_;
  assign new_F9290_ = ~F9235 | ~new_F9260_;
  assign new_F9291_ = new_F9268_ & new_F9288_;
  assign new_F9292_ = ~new_F9268_ & ~new_F9288_;
  assign new_F9293_ = new_F9297_ | new_F9298_;
  assign new_F9294_ = ~F9239 & new_F9253_;
  assign new_F9295_ = new_F9299_ | new_F9300_;
  assign new_F9296_ = F9239 & new_F9253_;
  assign new_F9297_ = ~F9239 & ~new_F9253_;
  assign new_F9298_ = F9239 & ~new_F9253_;
  assign new_F9299_ = F9239 & ~new_F9253_;
  assign new_F9300_ = ~F9239 & new_F9253_;
  assign new_F9307_ = new_F9314_ & new_F9313_;
  assign new_F9308_ = new_F9316_ | new_F9315_;
  assign new_F9309_ = new_F9318_ | new_F9317_;
  assign new_F9310_ = new_F9320_ & new_F9319_;
  assign new_F9311_ = new_F9320_ & new_F9321_;
  assign new_F9312_ = new_F9313_ | new_F9322_;
  assign new_F9313_ = F9302 | new_F9325_;
  assign new_F9314_ = new_F9324_ | new_F9323_;
  assign new_F9315_ = new_F9329_ & new_F9328_;
  assign new_F9316_ = new_F9327_ & new_F9326_;
  assign new_F9317_ = new_F9332_ | new_F9331_;
  assign new_F9318_ = new_F9327_ & new_F9330_;
  assign new_F9319_ = F9302 | new_F9335_;
  assign new_F9320_ = new_F9334_ | new_F9333_;
  assign new_F9321_ = new_F9337_ | new_F9336_;
  assign new_F9322_ = ~new_F9313_ & new_F9339_;
  assign new_F9323_ = ~new_F9315_ & new_F9327_;
  assign new_F9324_ = new_F9315_ & ~new_F9327_;
  assign new_F9325_ = F9301 & ~F9302;
  assign new_F9326_ = ~new_F9348_ | ~new_F9349_;
  assign new_F9327_ = new_F9341_ | new_F9343_;
  assign new_F9328_ = new_F9351_ | new_F9350_;
  assign new_F9329_ = new_F9345_ | new_F9344_;
  assign new_F9330_ = ~new_F9353_ | ~new_F9352_;
  assign new_F9331_ = ~new_F9354_ & new_F9355_;
  assign new_F9332_ = new_F9354_ & ~new_F9355_;
  assign new_F9333_ = ~F9301 & F9302;
  assign new_F9334_ = F9301 & ~F9302;
  assign new_F9335_ = ~new_F9317_ | new_F9327_;
  assign new_F9336_ = new_F9317_ & new_F9327_;
  assign new_F9337_ = ~new_F9317_ & ~new_F9327_;
  assign new_F9338_ = new_F9359_ | new_F9358_;
  assign new_F9339_ = F9305 | new_F9338_;
  assign new_F9340_ = new_F9363_ | new_F9362_;
  assign new_F9341_ = ~F9305 & new_F9340_;
  assign new_F9342_ = new_F9361_ | new_F9360_;
  assign new_F9343_ = F9305 & new_F9342_;
  assign new_F9344_ = F9303 & ~new_F9313_;
  assign new_F9345_ = ~F9303 & new_F9313_;
  assign new_F9346_ = ~F9302 | ~new_F9327_;
  assign new_F9347_ = new_F9313_ & new_F9346_;
  assign new_F9348_ = ~new_F9313_ & ~new_F9347_;
  assign new_F9349_ = new_F9313_ | new_F9346_;
  assign new_F9350_ = ~F9303 & F9304;
  assign new_F9351_ = F9303 & ~F9304;
  assign new_F9352_ = new_F9320_ | new_F9357_;
  assign new_F9353_ = ~new_F9320_ & ~new_F9356_;
  assign new_F9354_ = F9303 | new_F9320_;
  assign new_F9355_ = F9303 | F9304;
  assign new_F9356_ = new_F9320_ & new_F9357_;
  assign new_F9357_ = ~F9302 | ~new_F9327_;
  assign new_F9358_ = new_F9335_ & new_F9355_;
  assign new_F9359_ = ~new_F9335_ & ~new_F9355_;
  assign new_F9360_ = new_F9364_ | new_F9365_;
  assign new_F9361_ = ~F9306 & new_F9320_;
  assign new_F9362_ = new_F9366_ | new_F9367_;
  assign new_F9363_ = F9306 & new_F9320_;
  assign new_F9364_ = ~F9306 & ~new_F9320_;
  assign new_F9365_ = F9306 & ~new_F9320_;
  assign new_F9366_ = F9306 & ~new_F9320_;
  assign new_F9367_ = ~F9306 & new_F9320_;
  assign new_F9374_ = new_F9381_ & new_F9380_;
  assign new_F9375_ = new_F9383_ | new_F9382_;
  assign new_F9376_ = new_F9385_ | new_F9384_;
  assign new_F9377_ = new_F9387_ & new_F9386_;
  assign new_F9378_ = new_F9387_ & new_F9388_;
  assign new_F9379_ = new_F9380_ | new_F9389_;
  assign new_F9380_ = F9369 | new_F9392_;
  assign new_F9381_ = new_F9391_ | new_F9390_;
  assign new_F9382_ = new_F9396_ & new_F9395_;
  assign new_F9383_ = new_F9394_ & new_F9393_;
  assign new_F9384_ = new_F9399_ | new_F9398_;
  assign new_F9385_ = new_F9394_ & new_F9397_;
  assign new_F9386_ = F9369 | new_F9402_;
  assign new_F9387_ = new_F9401_ | new_F9400_;
  assign new_F9388_ = new_F9404_ | new_F9403_;
  assign new_F9389_ = ~new_F9380_ & new_F9406_;
  assign new_F9390_ = ~new_F9382_ & new_F9394_;
  assign new_F9391_ = new_F9382_ & ~new_F9394_;
  assign new_F9392_ = F9368 & ~F9369;
  assign new_F9393_ = ~new_F9415_ | ~new_F9416_;
  assign new_F9394_ = new_F9408_ | new_F9410_;
  assign new_F9395_ = new_F9418_ | new_F9417_;
  assign new_F9396_ = new_F9412_ | new_F9411_;
  assign new_F9397_ = ~new_F9420_ | ~new_F9419_;
  assign new_F9398_ = ~new_F9421_ & new_F9422_;
  assign new_F9399_ = new_F9421_ & ~new_F9422_;
  assign new_F9400_ = ~F9368 & F9369;
  assign new_F9401_ = F9368 & ~F9369;
  assign new_F9402_ = ~new_F9384_ | new_F9394_;
  assign new_F9403_ = new_F9384_ & new_F9394_;
  assign new_F9404_ = ~new_F9384_ & ~new_F9394_;
  assign new_F9405_ = new_F9426_ | new_F9425_;
  assign new_F9406_ = F9372 | new_F9405_;
  assign new_F9407_ = new_F9430_ | new_F9429_;
  assign new_F9408_ = ~F9372 & new_F9407_;
  assign new_F9409_ = new_F9428_ | new_F9427_;
  assign new_F9410_ = F9372 & new_F9409_;
  assign new_F9411_ = F9370 & ~new_F9380_;
  assign new_F9412_ = ~F9370 & new_F9380_;
  assign new_F9413_ = ~F9369 | ~new_F9394_;
  assign new_F9414_ = new_F9380_ & new_F9413_;
  assign new_F9415_ = ~new_F9380_ & ~new_F9414_;
  assign new_F9416_ = new_F9380_ | new_F9413_;
  assign new_F9417_ = ~F9370 & F9371;
  assign new_F9418_ = F9370 & ~F9371;
  assign new_F9419_ = new_F9387_ | new_F9424_;
  assign new_F9420_ = ~new_F9387_ & ~new_F9423_;
  assign new_F9421_ = F9370 | new_F9387_;
  assign new_F9422_ = F9370 | F9371;
  assign new_F9423_ = new_F9387_ & new_F9424_;
  assign new_F9424_ = ~F9369 | ~new_F9394_;
  assign new_F9425_ = new_F9402_ & new_F9422_;
  assign new_F9426_ = ~new_F9402_ & ~new_F9422_;
  assign new_F9427_ = new_F9431_ | new_F9432_;
  assign new_F9428_ = ~F9373 & new_F9387_;
  assign new_F9429_ = new_F9433_ | new_F9434_;
  assign new_F9430_ = F9373 & new_F9387_;
  assign new_F9431_ = ~F9373 & ~new_F9387_;
  assign new_F9432_ = F9373 & ~new_F9387_;
  assign new_F9433_ = F9373 & ~new_F9387_;
  assign new_F9434_ = ~F9373 & new_F9387_;
  assign new_F9441_ = new_F9448_ & new_F9447_;
  assign new_F9442_ = new_F9450_ | new_F9449_;
  assign new_F9443_ = new_F9452_ | new_F9451_;
  assign new_F9444_ = new_F9454_ & new_F9453_;
  assign new_F9445_ = new_F9454_ & new_F9455_;
  assign new_F9446_ = new_F9447_ | new_F9456_;
  assign new_F9447_ = F9436 | new_F9459_;
  assign new_F9448_ = new_F9458_ | new_F9457_;
  assign new_F9449_ = new_F9463_ & new_F9462_;
  assign new_F9450_ = new_F9461_ & new_F9460_;
  assign new_F9451_ = new_F9466_ | new_F9465_;
  assign new_F9452_ = new_F9461_ & new_F9464_;
  assign new_F9453_ = F9436 | new_F9469_;
  assign new_F9454_ = new_F9468_ | new_F9467_;
  assign new_F9455_ = new_F9471_ | new_F9470_;
  assign new_F9456_ = ~new_F9447_ & new_F9473_;
  assign new_F9457_ = ~new_F9449_ & new_F9461_;
  assign new_F9458_ = new_F9449_ & ~new_F9461_;
  assign new_F9459_ = F9435 & ~F9436;
  assign new_F9460_ = ~new_F9482_ | ~new_F9483_;
  assign new_F9461_ = new_F9475_ | new_F9477_;
  assign new_F9462_ = new_F9485_ | new_F9484_;
  assign new_F9463_ = new_F9479_ | new_F9478_;
  assign new_F9464_ = ~new_F9487_ | ~new_F9486_;
  assign new_F9465_ = ~new_F9488_ & new_F9489_;
  assign new_F9466_ = new_F9488_ & ~new_F9489_;
  assign new_F9467_ = ~F9435 & F9436;
  assign new_F9468_ = F9435 & ~F9436;
  assign new_F9469_ = ~new_F9451_ | new_F9461_;
  assign new_F9470_ = new_F9451_ & new_F9461_;
  assign new_F9471_ = ~new_F9451_ & ~new_F9461_;
  assign new_F9472_ = new_F9493_ | new_F9492_;
  assign new_F9473_ = F9439 | new_F9472_;
  assign new_F9474_ = new_F9497_ | new_F9496_;
  assign new_F9475_ = ~F9439 & new_F9474_;
  assign new_F9476_ = new_F9495_ | new_F9494_;
  assign new_F9477_ = F9439 & new_F9476_;
  assign new_F9478_ = F9437 & ~new_F9447_;
  assign new_F9479_ = ~F9437 & new_F9447_;
  assign new_F9480_ = ~F9436 | ~new_F9461_;
  assign new_F9481_ = new_F9447_ & new_F9480_;
  assign new_F9482_ = ~new_F9447_ & ~new_F9481_;
  assign new_F9483_ = new_F9447_ | new_F9480_;
  assign new_F9484_ = ~F9437 & F9438;
  assign new_F9485_ = F9437 & ~F9438;
  assign new_F9486_ = new_F9454_ | new_F9491_;
  assign new_F9487_ = ~new_F9454_ & ~new_F9490_;
  assign new_F9488_ = F9437 | new_F9454_;
  assign new_F9489_ = F9437 | F9438;
  assign new_F9490_ = new_F9454_ & new_F9491_;
  assign new_F9491_ = ~F9436 | ~new_F9461_;
  assign new_F9492_ = new_F9469_ & new_F9489_;
  assign new_F9493_ = ~new_F9469_ & ~new_F9489_;
  assign new_F9494_ = new_F9498_ | new_F9499_;
  assign new_F9495_ = ~F9440 & new_F9454_;
  assign new_F9496_ = new_F9500_ | new_F9501_;
  assign new_F9497_ = F9440 & new_F9454_;
  assign new_F9498_ = ~F9440 & ~new_F9454_;
  assign new_F9499_ = F9440 & ~new_F9454_;
  assign new_F9500_ = F9440 & ~new_F9454_;
  assign new_F9501_ = ~F9440 & new_F9454_;
  assign new_F9508_ = new_F9515_ & new_F9514_;
  assign new_F9509_ = new_F9517_ | new_F9516_;
  assign new_F9510_ = new_F9519_ | new_F9518_;
  assign new_F9511_ = new_F9521_ & new_F9520_;
  assign new_F9512_ = new_F9521_ & new_F9522_;
  assign new_F9513_ = new_F9514_ | new_F9523_;
  assign new_F9514_ = F9503 | new_F9526_;
  assign new_F9515_ = new_F9525_ | new_F9524_;
  assign new_F9516_ = new_F9530_ & new_F9529_;
  assign new_F9517_ = new_F9528_ & new_F9527_;
  assign new_F9518_ = new_F9533_ | new_F9532_;
  assign new_F9519_ = new_F9528_ & new_F9531_;
  assign new_F9520_ = F9503 | new_F9536_;
  assign new_F9521_ = new_F9535_ | new_F9534_;
  assign new_F9522_ = new_F9538_ | new_F9537_;
  assign new_F9523_ = ~new_F9514_ & new_F9540_;
  assign new_F9524_ = ~new_F9516_ & new_F9528_;
  assign new_F9525_ = new_F9516_ & ~new_F9528_;
  assign new_F9526_ = F9502 & ~F9503;
  assign new_F9527_ = ~new_F9549_ | ~new_F9550_;
  assign new_F9528_ = new_F9542_ | new_F9544_;
  assign new_F9529_ = new_F9552_ | new_F9551_;
  assign new_F9530_ = new_F9546_ | new_F9545_;
  assign new_F9531_ = ~new_F9554_ | ~new_F9553_;
  assign new_F9532_ = ~new_F9555_ & new_F9556_;
  assign new_F9533_ = new_F9555_ & ~new_F9556_;
  assign new_F9534_ = ~F9502 & F9503;
  assign new_F9535_ = F9502 & ~F9503;
  assign new_F9536_ = ~new_F9518_ | new_F9528_;
  assign new_F9537_ = new_F9518_ & new_F9528_;
  assign new_F9538_ = ~new_F9518_ & ~new_F9528_;
  assign new_F9539_ = new_F9560_ | new_F9559_;
  assign new_F9540_ = F9506 | new_F9539_;
  assign new_F9541_ = new_F9564_ | new_F9563_;
  assign new_F9542_ = ~F9506 & new_F9541_;
  assign new_F9543_ = new_F9562_ | new_F9561_;
  assign new_F9544_ = F9506 & new_F9543_;
  assign new_F9545_ = F9504 & ~new_F9514_;
  assign new_F9546_ = ~F9504 & new_F9514_;
  assign new_F9547_ = ~F9503 | ~new_F9528_;
  assign new_F9548_ = new_F9514_ & new_F9547_;
  assign new_F9549_ = ~new_F9514_ & ~new_F9548_;
  assign new_F9550_ = new_F9514_ | new_F9547_;
  assign new_F9551_ = ~F9504 & F9505;
  assign new_F9552_ = F9504 & ~F9505;
  assign new_F9553_ = new_F9521_ | new_F9558_;
  assign new_F9554_ = ~new_F9521_ & ~new_F9557_;
  assign new_F9555_ = F9504 | new_F9521_;
  assign new_F9556_ = F9504 | F9505;
  assign new_F9557_ = new_F9521_ & new_F9558_;
  assign new_F9558_ = ~F9503 | ~new_F9528_;
  assign new_F9559_ = new_F9536_ & new_F9556_;
  assign new_F9560_ = ~new_F9536_ & ~new_F9556_;
  assign new_F9561_ = new_F9565_ | new_F9566_;
  assign new_F9562_ = ~F9507 & new_F9521_;
  assign new_F9563_ = new_F9567_ | new_F9568_;
  assign new_F9564_ = F9507 & new_F9521_;
  assign new_F9565_ = ~F9507 & ~new_F9521_;
  assign new_F9566_ = F9507 & ~new_F9521_;
  assign new_F9567_ = F9507 & ~new_F9521_;
  assign new_F9568_ = ~F9507 & new_F9521_;
  assign new_F9575_ = new_F9582_ & new_F9581_;
  assign new_F9576_ = new_F9584_ | new_F9583_;
  assign new_F9577_ = new_F9586_ | new_F9585_;
  assign new_F9578_ = new_F9588_ & new_F9587_;
  assign new_F9579_ = new_F9588_ & new_F9589_;
  assign new_F9580_ = new_F9581_ | new_F9590_;
  assign new_F9581_ = F9570 | new_F9593_;
  assign new_F9582_ = new_F9592_ | new_F9591_;
  assign new_F9583_ = new_F9597_ & new_F9596_;
  assign new_F9584_ = new_F9595_ & new_F9594_;
  assign new_F9585_ = new_F9600_ | new_F9599_;
  assign new_F9586_ = new_F9595_ & new_F9598_;
  assign new_F9587_ = F9570 | new_F9603_;
  assign new_F9588_ = new_F9602_ | new_F9601_;
  assign new_F9589_ = new_F9605_ | new_F9604_;
  assign new_F9590_ = ~new_F9581_ & new_F9607_;
  assign new_F9591_ = ~new_F9583_ & new_F9595_;
  assign new_F9592_ = new_F9583_ & ~new_F9595_;
  assign new_F9593_ = F9569 & ~F9570;
  assign new_F9594_ = ~new_F9616_ | ~new_F9617_;
  assign new_F9595_ = new_F9609_ | new_F9611_;
  assign new_F9596_ = new_F9619_ | new_F9618_;
  assign new_F9597_ = new_F9613_ | new_F9612_;
  assign new_F9598_ = ~new_F9621_ | ~new_F9620_;
  assign new_F9599_ = ~new_F9622_ & new_F9623_;
  assign new_F9600_ = new_F9622_ & ~new_F9623_;
  assign new_F9601_ = ~F9569 & F9570;
  assign new_F9602_ = F9569 & ~F9570;
  assign new_F9603_ = ~new_F9585_ | new_F9595_;
  assign new_F9604_ = new_F9585_ & new_F9595_;
  assign new_F9605_ = ~new_F9585_ & ~new_F9595_;
  assign new_F9606_ = new_F9627_ | new_F9626_;
  assign new_F9607_ = F9573 | new_F9606_;
  assign new_F9608_ = new_F9631_ | new_F9630_;
  assign new_F9609_ = ~F9573 & new_F9608_;
  assign new_F9610_ = new_F9629_ | new_F9628_;
  assign new_F9611_ = F9573 & new_F9610_;
  assign new_F9612_ = F9571 & ~new_F9581_;
  assign new_F9613_ = ~F9571 & new_F9581_;
  assign new_F9614_ = ~F9570 | ~new_F9595_;
  assign new_F9615_ = new_F9581_ & new_F9614_;
  assign new_F9616_ = ~new_F9581_ & ~new_F9615_;
  assign new_F9617_ = new_F9581_ | new_F9614_;
  assign new_F9618_ = ~F9571 & F9572;
  assign new_F9619_ = F9571 & ~F9572;
  assign new_F9620_ = new_F9588_ | new_F9625_;
  assign new_F9621_ = ~new_F9588_ & ~new_F9624_;
  assign new_F9622_ = F9571 | new_F9588_;
  assign new_F9623_ = F9571 | F9572;
  assign new_F9624_ = new_F9588_ & new_F9625_;
  assign new_F9625_ = ~F9570 | ~new_F9595_;
  assign new_F9626_ = new_F9603_ & new_F9623_;
  assign new_F9627_ = ~new_F9603_ & ~new_F9623_;
  assign new_F9628_ = new_F9632_ | new_F9633_;
  assign new_F9629_ = ~F9574 & new_F9588_;
  assign new_F9630_ = new_F9634_ | new_F9635_;
  assign new_F9631_ = F9574 & new_F9588_;
  assign new_F9632_ = ~F9574 & ~new_F9588_;
  assign new_F9633_ = F9574 & ~new_F9588_;
  assign new_F9634_ = F9574 & ~new_F9588_;
  assign new_F9635_ = ~F9574 & new_F9588_;
  assign new_F9642_ = new_F9649_ & new_F9648_;
  assign new_F9643_ = new_F9651_ | new_F9650_;
  assign new_F9644_ = new_F9653_ | new_F9652_;
  assign new_F9645_ = new_F9655_ & new_F9654_;
  assign new_F9646_ = new_F9655_ & new_F9656_;
  assign new_F9647_ = new_F9648_ | new_F9657_;
  assign new_F9648_ = F9637 | new_F9660_;
  assign new_F9649_ = new_F9659_ | new_F9658_;
  assign new_F9650_ = new_F9664_ & new_F9663_;
  assign new_F9651_ = new_F9662_ & new_F9661_;
  assign new_F9652_ = new_F9667_ | new_F9666_;
  assign new_F9653_ = new_F9662_ & new_F9665_;
  assign new_F9654_ = F9637 | new_F9670_;
  assign new_F9655_ = new_F9669_ | new_F9668_;
  assign new_F9656_ = new_F9672_ | new_F9671_;
  assign new_F9657_ = ~new_F9648_ & new_F9674_;
  assign new_F9658_ = ~new_F9650_ & new_F9662_;
  assign new_F9659_ = new_F9650_ & ~new_F9662_;
  assign new_F9660_ = F9636 & ~F9637;
  assign new_F9661_ = ~new_F9683_ | ~new_F9684_;
  assign new_F9662_ = new_F9676_ | new_F9678_;
  assign new_F9663_ = new_F9686_ | new_F9685_;
  assign new_F9664_ = new_F9680_ | new_F9679_;
  assign new_F9665_ = ~new_F9688_ | ~new_F9687_;
  assign new_F9666_ = ~new_F9689_ & new_F9690_;
  assign new_F9667_ = new_F9689_ & ~new_F9690_;
  assign new_F9668_ = ~F9636 & F9637;
  assign new_F9669_ = F9636 & ~F9637;
  assign new_F9670_ = ~new_F9652_ | new_F9662_;
  assign new_F9671_ = new_F9652_ & new_F9662_;
  assign new_F9672_ = ~new_F9652_ & ~new_F9662_;
  assign new_F9673_ = new_F9694_ | new_F9693_;
  assign new_F9674_ = F9640 | new_F9673_;
  assign new_F9675_ = new_F9698_ | new_F9697_;
  assign new_F9676_ = ~F9640 & new_F9675_;
  assign new_F9677_ = new_F9696_ | new_F9695_;
  assign new_F9678_ = F9640 & new_F9677_;
  assign new_F9679_ = F9638 & ~new_F9648_;
  assign new_F9680_ = ~F9638 & new_F9648_;
  assign new_F9681_ = ~F9637 | ~new_F9662_;
  assign new_F9682_ = new_F9648_ & new_F9681_;
  assign new_F9683_ = ~new_F9648_ & ~new_F9682_;
  assign new_F9684_ = new_F9648_ | new_F9681_;
  assign new_F9685_ = ~F9638 & F9639;
  assign new_F9686_ = F9638 & ~F9639;
  assign new_F9687_ = new_F9655_ | new_F9692_;
  assign new_F9688_ = ~new_F9655_ & ~new_F9691_;
  assign new_F9689_ = F9638 | new_F9655_;
  assign new_F9690_ = F9638 | F9639;
  assign new_F9691_ = new_F9655_ & new_F9692_;
  assign new_F9692_ = ~F9637 | ~new_F9662_;
  assign new_F9693_ = new_F9670_ & new_F9690_;
  assign new_F9694_ = ~new_F9670_ & ~new_F9690_;
  assign new_F9695_ = new_F9699_ | new_F9700_;
  assign new_F9696_ = ~F9641 & new_F9655_;
  assign new_F9697_ = new_F9701_ | new_F9702_;
  assign new_F9698_ = F9641 & new_F9655_;
  assign new_F9699_ = ~F9641 & ~new_F9655_;
  assign new_F9700_ = F9641 & ~new_F9655_;
  assign new_F9701_ = F9641 & ~new_F9655_;
  assign new_F9702_ = ~F9641 & new_F9655_;
  assign new_F9709_ = new_F9716_ & new_F9715_;
  assign new_F9710_ = new_F9718_ | new_F9717_;
  assign new_F9711_ = new_F9720_ | new_F9719_;
  assign new_F9712_ = new_F9722_ & new_F9721_;
  assign new_F9713_ = new_F9722_ & new_F9723_;
  assign new_F9714_ = new_F9715_ | new_F9724_;
  assign new_F9715_ = F9704 | new_F9727_;
  assign new_F9716_ = new_F9726_ | new_F9725_;
  assign new_F9717_ = new_F9731_ & new_F9730_;
  assign new_F9718_ = new_F9729_ & new_F9728_;
  assign new_F9719_ = new_F9734_ | new_F9733_;
  assign new_F9720_ = new_F9729_ & new_F9732_;
  assign new_F9721_ = F9704 | new_F9737_;
  assign new_F9722_ = new_F9736_ | new_F9735_;
  assign new_F9723_ = new_F9739_ | new_F9738_;
  assign new_F9724_ = ~new_F9715_ & new_F9741_;
  assign new_F9725_ = ~new_F9717_ & new_F9729_;
  assign new_F9726_ = new_F9717_ & ~new_F9729_;
  assign new_F9727_ = F9703 & ~F9704;
  assign new_F9728_ = ~new_F9750_ | ~new_F9751_;
  assign new_F9729_ = new_F9743_ | new_F9745_;
  assign new_F9730_ = new_F9753_ | new_F9752_;
  assign new_F9731_ = new_F9747_ | new_F9746_;
  assign new_F9732_ = ~new_F9755_ | ~new_F9754_;
  assign new_F9733_ = ~new_F9756_ & new_F9757_;
  assign new_F9734_ = new_F9756_ & ~new_F9757_;
  assign new_F9735_ = ~F9703 & F9704;
  assign new_F9736_ = F9703 & ~F9704;
  assign new_F9737_ = ~new_F9719_ | new_F9729_;
  assign new_F9738_ = new_F9719_ & new_F9729_;
  assign new_F9739_ = ~new_F9719_ & ~new_F9729_;
  assign new_F9740_ = new_F9761_ | new_F9760_;
  assign new_F9741_ = F9707 | new_F9740_;
  assign new_F9742_ = new_F9765_ | new_F9764_;
  assign new_F9743_ = ~F9707 & new_F9742_;
  assign new_F9744_ = new_F9763_ | new_F9762_;
  assign new_F9745_ = F9707 & new_F9744_;
  assign new_F9746_ = F9705 & ~new_F9715_;
  assign new_F9747_ = ~F9705 & new_F9715_;
  assign new_F9748_ = ~F9704 | ~new_F9729_;
  assign new_F9749_ = new_F9715_ & new_F9748_;
  assign new_F9750_ = ~new_F9715_ & ~new_F9749_;
  assign new_F9751_ = new_F9715_ | new_F9748_;
  assign new_F9752_ = ~F9705 & F9706;
  assign new_F9753_ = F9705 & ~F9706;
  assign new_F9754_ = new_F9722_ | new_F9759_;
  assign new_F9755_ = ~new_F9722_ & ~new_F9758_;
  assign new_F9756_ = F9705 | new_F9722_;
  assign new_F9757_ = F9705 | F9706;
  assign new_F9758_ = new_F9722_ & new_F9759_;
  assign new_F9759_ = ~F9704 | ~new_F9729_;
  assign new_F9760_ = new_F9737_ & new_F9757_;
  assign new_F9761_ = ~new_F9737_ & ~new_F9757_;
  assign new_F9762_ = new_F9766_ | new_F9767_;
  assign new_F9763_ = ~F9708 & new_F9722_;
  assign new_F9764_ = new_F9768_ | new_F9769_;
  assign new_F9765_ = F9708 & new_F9722_;
  assign new_F9766_ = ~F9708 & ~new_F9722_;
  assign new_F9767_ = F9708 & ~new_F9722_;
  assign new_F9768_ = F9708 & ~new_F9722_;
  assign new_F9769_ = ~F9708 & new_F9722_;
  assign new_F9776_ = new_F9783_ & new_F9782_;
  assign new_F9777_ = new_F9785_ | new_F9784_;
  assign new_F9778_ = new_F9787_ | new_F9786_;
  assign new_F9779_ = new_F9789_ & new_F9788_;
  assign new_F9780_ = new_F9789_ & new_F9790_;
  assign new_F9781_ = new_F9782_ | new_F9791_;
  assign new_F9782_ = F9771 | new_F9794_;
  assign new_F9783_ = new_F9793_ | new_F9792_;
  assign new_F9784_ = new_F9798_ & new_F9797_;
  assign new_F9785_ = new_F9796_ & new_F9795_;
  assign new_F9786_ = new_F9801_ | new_F9800_;
  assign new_F9787_ = new_F9796_ & new_F9799_;
  assign new_F9788_ = F9771 | new_F9804_;
  assign new_F9789_ = new_F9803_ | new_F9802_;
  assign new_F9790_ = new_F9806_ | new_F9805_;
  assign new_F9791_ = ~new_F9782_ & new_F9808_;
  assign new_F9792_ = ~new_F9784_ & new_F9796_;
  assign new_F9793_ = new_F9784_ & ~new_F9796_;
  assign new_F9794_ = F9770 & ~F9771;
  assign new_F9795_ = ~new_F9817_ | ~new_F9818_;
  assign new_F9796_ = new_F9810_ | new_F9812_;
  assign new_F9797_ = new_F9820_ | new_F9819_;
  assign new_F9798_ = new_F9814_ | new_F9813_;
  assign new_F9799_ = ~new_F9822_ | ~new_F9821_;
  assign new_F9800_ = ~new_F9823_ & new_F9824_;
  assign new_F9801_ = new_F9823_ & ~new_F9824_;
  assign new_F9802_ = ~F9770 & F9771;
  assign new_F9803_ = F9770 & ~F9771;
  assign new_F9804_ = ~new_F9786_ | new_F9796_;
  assign new_F9805_ = new_F9786_ & new_F9796_;
  assign new_F9806_ = ~new_F9786_ & ~new_F9796_;
  assign new_F9807_ = new_F9828_ | new_F9827_;
  assign new_F9808_ = F9774 | new_F9807_;
  assign new_F9809_ = new_F9832_ | new_F9831_;
  assign new_F9810_ = ~F9774 & new_F9809_;
  assign new_F9811_ = new_F9830_ | new_F9829_;
  assign new_F9812_ = F9774 & new_F9811_;
  assign new_F9813_ = F9772 & ~new_F9782_;
  assign new_F9814_ = ~F9772 & new_F9782_;
  assign new_F9815_ = ~F9771 | ~new_F9796_;
  assign new_F9816_ = new_F9782_ & new_F9815_;
  assign new_F9817_ = ~new_F9782_ & ~new_F9816_;
  assign new_F9818_ = new_F9782_ | new_F9815_;
  assign new_F9819_ = ~F9772 & F9773;
  assign new_F9820_ = F9772 & ~F9773;
  assign new_F9821_ = new_F9789_ | new_F9826_;
  assign new_F9822_ = ~new_F9789_ & ~new_F9825_;
  assign new_F9823_ = F9772 | new_F9789_;
  assign new_F9824_ = F9772 | F9773;
  assign new_F9825_ = new_F9789_ & new_F9826_;
  assign new_F9826_ = ~F9771 | ~new_F9796_;
  assign new_F9827_ = new_F9804_ & new_F9824_;
  assign new_F9828_ = ~new_F9804_ & ~new_F9824_;
  assign new_F9829_ = new_F9833_ | new_F9834_;
  assign new_F9830_ = ~F9775 & new_F9789_;
  assign new_F9831_ = new_F9835_ | new_F9836_;
  assign new_F9832_ = F9775 & new_F9789_;
  assign new_F9833_ = ~F9775 & ~new_F9789_;
  assign new_F9834_ = F9775 & ~new_F9789_;
  assign new_F9835_ = F9775 & ~new_F9789_;
  assign new_F9836_ = ~F9775 & new_F9789_;
  assign new_F9843_ = new_F9850_ & new_F9849_;
  assign new_F9844_ = new_F9852_ | new_F9851_;
  assign new_F9845_ = new_F9854_ | new_F9853_;
  assign new_F9846_ = new_F9856_ & new_F9855_;
  assign new_F9847_ = new_F9856_ & new_F9857_;
  assign new_F9848_ = new_F9849_ | new_F9858_;
  assign new_F9849_ = F9838 | new_F9861_;
  assign new_F9850_ = new_F9860_ | new_F9859_;
  assign new_F9851_ = new_F9865_ & new_F9864_;
  assign new_F9852_ = new_F9863_ & new_F9862_;
  assign new_F9853_ = new_F9868_ | new_F9867_;
  assign new_F9854_ = new_F9863_ & new_F9866_;
  assign new_F9855_ = F9838 | new_F9871_;
  assign new_F9856_ = new_F9870_ | new_F9869_;
  assign new_F9857_ = new_F9873_ | new_F9872_;
  assign new_F9858_ = ~new_F9849_ & new_F9875_;
  assign new_F9859_ = ~new_F9851_ & new_F9863_;
  assign new_F9860_ = new_F9851_ & ~new_F9863_;
  assign new_F9861_ = F9837 & ~F9838;
  assign new_F9862_ = ~new_F9884_ | ~new_F9885_;
  assign new_F9863_ = new_F9877_ | new_F9879_;
  assign new_F9864_ = new_F9887_ | new_F9886_;
  assign new_F9865_ = new_F9881_ | new_F9880_;
  assign new_F9866_ = ~new_F9889_ | ~new_F9888_;
  assign new_F9867_ = ~new_F9890_ & new_F9891_;
  assign new_F9868_ = new_F9890_ & ~new_F9891_;
  assign new_F9869_ = ~F9837 & F9838;
  assign new_F9870_ = F9837 & ~F9838;
  assign new_F9871_ = ~new_F9853_ | new_F9863_;
  assign new_F9872_ = new_F9853_ & new_F9863_;
  assign new_F9873_ = ~new_F9853_ & ~new_F9863_;
  assign new_F9874_ = new_F9895_ | new_F9894_;
  assign new_F9875_ = F9841 | new_F9874_;
  assign new_F9876_ = new_F9899_ | new_F9898_;
  assign new_F9877_ = ~F9841 & new_F9876_;
  assign new_F9878_ = new_F9897_ | new_F9896_;
  assign new_F9879_ = F9841 & new_F9878_;
  assign new_F9880_ = F9839 & ~new_F9849_;
  assign new_F9881_ = ~F9839 & new_F9849_;
  assign new_F9882_ = ~F9838 | ~new_F9863_;
  assign new_F9883_ = new_F9849_ & new_F9882_;
  assign new_F9884_ = ~new_F9849_ & ~new_F9883_;
  assign new_F9885_ = new_F9849_ | new_F9882_;
  assign new_F9886_ = ~F9839 & F9840;
  assign new_F9887_ = F9839 & ~F9840;
  assign new_F9888_ = new_F9856_ | new_F9893_;
  assign new_F9889_ = ~new_F9856_ & ~new_F9892_;
  assign new_F9890_ = F9839 | new_F9856_;
  assign new_F9891_ = F9839 | F9840;
  assign new_F9892_ = new_F9856_ & new_F9893_;
  assign new_F9893_ = ~F9838 | ~new_F9863_;
  assign new_F9894_ = new_F9871_ & new_F9891_;
  assign new_F9895_ = ~new_F9871_ & ~new_F9891_;
  assign new_F9896_ = new_F9900_ | new_F9901_;
  assign new_F9897_ = ~F9842 & new_F9856_;
  assign new_F9898_ = new_F9902_ | new_F9903_;
  assign new_F9899_ = F9842 & new_F9856_;
  assign new_F9900_ = ~F9842 & ~new_F9856_;
  assign new_F9901_ = F9842 & ~new_F9856_;
  assign new_F9902_ = F9842 & ~new_F9856_;
  assign new_F9903_ = ~F9842 & new_F9856_;
  assign new_F9910_ = new_F9917_ & new_F9916_;
  assign new_F9911_ = new_F9919_ | new_F9918_;
  assign new_F9912_ = new_F9921_ | new_F9920_;
  assign new_F9913_ = new_F9923_ & new_F9922_;
  assign new_F9914_ = new_F9923_ & new_F9924_;
  assign new_F9915_ = new_F9916_ | new_F9925_;
  assign new_F9916_ = F9905 | new_F9928_;
  assign new_F9917_ = new_F9927_ | new_F9926_;
  assign new_F9918_ = new_F9932_ & new_F9931_;
  assign new_F9919_ = new_F9930_ & new_F9929_;
  assign new_F9920_ = new_F9935_ | new_F9934_;
  assign new_F9921_ = new_F9930_ & new_F9933_;
  assign new_F9922_ = F9905 | new_F9938_;
  assign new_F9923_ = new_F9937_ | new_F9936_;
  assign new_F9924_ = new_F9940_ | new_F9939_;
  assign new_F9925_ = ~new_F9916_ & new_F9942_;
  assign new_F9926_ = ~new_F9918_ & new_F9930_;
  assign new_F9927_ = new_F9918_ & ~new_F9930_;
  assign new_F9928_ = F9904 & ~F9905;
  assign new_F9929_ = ~new_F9951_ | ~new_F9952_;
  assign new_F9930_ = new_F9944_ | new_F9946_;
  assign new_F9931_ = new_F9954_ | new_F9953_;
  assign new_F9932_ = new_F9948_ | new_F9947_;
  assign new_F9933_ = ~new_F9956_ | ~new_F9955_;
  assign new_F9934_ = ~new_F9957_ & new_F9958_;
  assign new_F9935_ = new_F9957_ & ~new_F9958_;
  assign new_F9936_ = ~F9904 & F9905;
  assign new_F9937_ = F9904 & ~F9905;
  assign new_F9938_ = ~new_F9920_ | new_F9930_;
  assign new_F9939_ = new_F9920_ & new_F9930_;
  assign new_F9940_ = ~new_F9920_ & ~new_F9930_;
  assign new_F9941_ = new_F9962_ | new_F9961_;
  assign new_F9942_ = F9908 | new_F9941_;
  assign new_F9943_ = new_F9966_ | new_F9965_;
  assign new_F9944_ = ~F9908 & new_F9943_;
  assign new_F9945_ = new_F9964_ | new_F9963_;
  assign new_F9946_ = F9908 & new_F9945_;
  assign new_F9947_ = F9906 & ~new_F9916_;
  assign new_F9948_ = ~F9906 & new_F9916_;
  assign new_F9949_ = ~F9905 | ~new_F9930_;
  assign new_F9950_ = new_F9916_ & new_F9949_;
  assign new_F9951_ = ~new_F9916_ & ~new_F9950_;
  assign new_F9952_ = new_F9916_ | new_F9949_;
  assign new_F9953_ = ~F9906 & F9907;
  assign new_F9954_ = F9906 & ~F9907;
  assign new_F9955_ = new_F9923_ | new_F9960_;
  assign new_F9956_ = ~new_F9923_ & ~new_F9959_;
  assign new_F9957_ = F9906 | new_F9923_;
  assign new_F9958_ = F9906 | F9907;
  assign new_F9959_ = new_F9923_ & new_F9960_;
  assign new_F9960_ = ~F9905 | ~new_F9930_;
  assign new_F9961_ = new_F9938_ & new_F9958_;
  assign new_F9962_ = ~new_F9938_ & ~new_F9958_;
  assign new_F9963_ = new_F9967_ | new_F9968_;
  assign new_F9964_ = ~F9909 & new_F9923_;
  assign new_F9965_ = new_F9969_ | new_F9970_;
  assign new_F9966_ = F9909 & new_F9923_;
  assign new_F9967_ = ~F9909 & ~new_F9923_;
  assign new_F9968_ = F9909 & ~new_F9923_;
  assign new_F9969_ = F9909 & ~new_F9923_;
  assign new_F9970_ = ~F9909 & new_F9923_;
  assign new_F9977_ = new_F9984_ & new_F9983_;
  assign new_F9978_ = new_F9986_ | new_F9985_;
  assign new_F9979_ = new_F9988_ | new_F9987_;
  assign new_F9980_ = new_F9990_ & new_F9989_;
  assign new_F9981_ = new_F9990_ & new_F9991_;
  assign new_F9982_ = new_F9983_ | new_F9992_;
  assign new_F9983_ = F9972 | new_F9995_;
  assign new_F9984_ = new_F9994_ | new_F9993_;
  assign new_F9985_ = new_F9999_ & new_F9998_;
  assign new_F9986_ = new_F9997_ & new_F9996_;
  assign new_F9987_ = new_G3_ | new_G2_;
  assign new_F9988_ = new_F9997_ & new_G1_;
  assign new_F9989_ = F9972 | new_G6_;
  assign new_F9990_ = new_G5_ | new_G4_;
  assign new_F9991_ = new_G8_ | new_G7_;
  assign new_F9992_ = ~new_F9983_ & new_G10_;
  assign new_F9993_ = ~new_F9985_ & new_F9997_;
  assign new_F9994_ = new_F9985_ & ~new_F9997_;
  assign new_F9995_ = F9971 & ~F9972;
  assign new_F9996_ = ~new_G19_ | ~new_G20_;
  assign new_F9997_ = new_G12_ | new_G14_;
  assign new_F9998_ = new_G22_ | new_G21_;
  assign new_F9999_ = new_G16_ | new_G15_;
  assign new_G1_ = ~new_G24_ | ~new_G23_;
  assign new_G2_ = ~new_G25_ & new_G26_;
  assign new_G3_ = new_G25_ & ~new_G26_;
  assign new_G4_ = ~F9971 & F9972;
  assign new_G5_ = F9971 & ~F9972;
  assign new_G6_ = ~new_F9987_ | new_F9997_;
  assign new_G7_ = new_F9987_ & new_F9997_;
  assign new_G8_ = ~new_F9987_ & ~new_F9997_;
  assign new_G9_ = new_G30_ | new_G29_;
  assign new_G10_ = F9975 | new_G9_;
  assign new_G11_ = new_G34_ | new_G33_;
  assign new_G12_ = ~F9975 & new_G11_;
  assign new_G13_ = new_G32_ | new_G31_;
  assign new_G14_ = F9975 & new_G13_;
  assign new_G15_ = F9973 & ~new_F9983_;
  assign new_G16_ = ~F9973 & new_F9983_;
  assign new_G17_ = ~F9972 | ~new_F9997_;
  assign new_G18_ = new_F9983_ & new_G17_;
  assign new_G19_ = ~new_F9983_ & ~new_G18_;
  assign new_G20_ = new_F9983_ | new_G17_;
  assign new_G21_ = ~F9973 & F9974;
  assign new_G22_ = F9973 & ~F9974;
  assign new_G23_ = new_F9990_ | new_G28_;
  assign new_G24_ = ~new_F9990_ & ~new_G27_;
  assign new_G25_ = F9973 | new_F9990_;
  assign new_G26_ = F9973 | F9974;
  assign new_G27_ = new_F9990_ & new_G28_;
  assign new_G28_ = ~F9972 | ~new_F9997_;
  assign new_G29_ = new_G6_ & new_G26_;
  assign new_G30_ = ~new_G6_ & ~new_G26_;
  assign new_G31_ = new_G35_ | new_G36_;
  assign new_G32_ = ~F9976 & new_F9990_;
  assign new_G33_ = new_G37_ | new_G38_;
  assign new_G34_ = F9976 & new_F9990_;
  assign new_G35_ = ~F9976 & ~new_F9990_;
  assign new_G36_ = F9976 & ~new_F9990_;
  assign new_G37_ = F9976 & ~new_F9990_;
  assign new_G38_ = ~F9976 & new_F9990_;
  assign new_G45_ = new_G52_ & new_G51_;
  assign new_G46_ = new_G54_ | new_G53_;
  assign new_G47_ = new_G56_ | new_G55_;
  assign new_G48_ = new_G58_ & new_G57_;
  assign new_G49_ = new_G58_ & new_G59_;
  assign new_G50_ = new_G51_ | new_G60_;
  assign new_G51_ = G40 | new_G63_;
  assign new_G52_ = new_G62_ | new_G61_;
  assign new_G53_ = new_G67_ & new_G66_;
  assign new_G54_ = new_G65_ & new_G64_;
  assign new_G55_ = new_G70_ | new_G69_;
  assign new_G56_ = new_G65_ & new_G68_;
  assign new_G57_ = G40 | new_G73_;
  assign new_G58_ = new_G72_ | new_G71_;
  assign new_G59_ = new_G75_ | new_G74_;
  assign new_G60_ = ~new_G51_ & new_G77_;
  assign new_G61_ = ~new_G53_ & new_G65_;
  assign new_G62_ = new_G53_ & ~new_G65_;
  assign new_G63_ = G39 & ~G40;
  assign new_G64_ = ~new_G86_ | ~new_G87_;
  assign new_G65_ = new_G79_ | new_G81_;
  assign new_G66_ = new_G89_ | new_G88_;
  assign new_G67_ = new_G83_ | new_G82_;
  assign new_G68_ = ~new_G91_ | ~new_G90_;
  assign new_G69_ = ~new_G92_ & new_G93_;
  assign new_G70_ = new_G92_ & ~new_G93_;
  assign new_G71_ = ~G39 & G40;
  assign new_G72_ = G39 & ~G40;
  assign new_G73_ = ~new_G55_ | new_G65_;
  assign new_G74_ = new_G55_ & new_G65_;
  assign new_G75_ = ~new_G55_ & ~new_G65_;
  assign new_G76_ = new_G97_ | new_G96_;
  assign new_G77_ = G43 | new_G76_;
  assign new_G78_ = new_G101_ | new_G100_;
  assign new_G79_ = ~G43 & new_G78_;
  assign new_G80_ = new_G99_ | new_G98_;
  assign new_G81_ = G43 & new_G80_;
  assign new_G82_ = G41 & ~new_G51_;
  assign new_G83_ = ~G41 & new_G51_;
  assign new_G84_ = ~G40 | ~new_G65_;
  assign new_G85_ = new_G51_ & new_G84_;
  assign new_G86_ = ~new_G51_ & ~new_G85_;
  assign new_G87_ = new_G51_ | new_G84_;
  assign new_G88_ = ~G41 & G42;
  assign new_G89_ = G41 & ~G42;
  assign new_G90_ = new_G58_ | new_G95_;
  assign new_G91_ = ~new_G58_ & ~new_G94_;
  assign new_G92_ = G41 | new_G58_;
  assign new_G93_ = G41 | G42;
  assign new_G94_ = new_G58_ & new_G95_;
  assign new_G95_ = ~G40 | ~new_G65_;
  assign new_G96_ = new_G73_ & new_G93_;
  assign new_G97_ = ~new_G73_ & ~new_G93_;
  assign new_G98_ = new_G102_ | new_G103_;
  assign new_G99_ = ~G44 & new_G58_;
  assign new_G100_ = new_G104_ | new_G105_;
  assign new_G101_ = G44 & new_G58_;
  assign new_G102_ = ~G44 & ~new_G58_;
  assign new_G103_ = G44 & ~new_G58_;
  assign new_G104_ = G44 & ~new_G58_;
  assign new_G105_ = ~G44 & new_G58_;
  assign new_G112_ = new_G119_ & new_G118_;
  assign new_G113_ = new_G121_ | new_G120_;
  assign new_G114_ = new_G123_ | new_G122_;
  assign new_G115_ = new_G125_ & new_G124_;
  assign new_G116_ = new_G125_ & new_G126_;
  assign new_G117_ = new_G118_ | new_G127_;
  assign new_G118_ = G107 | new_G130_;
  assign new_G119_ = new_G129_ | new_G128_;
  assign new_G120_ = new_G134_ & new_G133_;
  assign new_G121_ = new_G132_ & new_G131_;
  assign new_G122_ = new_G137_ | new_G136_;
  assign new_G123_ = new_G132_ & new_G135_;
  assign new_G124_ = G107 | new_G140_;
  assign new_G125_ = new_G139_ | new_G138_;
  assign new_G126_ = new_G142_ | new_G141_;
  assign new_G127_ = ~new_G118_ & new_G144_;
  assign new_G128_ = ~new_G120_ & new_G132_;
  assign new_G129_ = new_G120_ & ~new_G132_;
  assign new_G130_ = G106 & ~G107;
  assign new_G131_ = ~new_G153_ | ~new_G154_;
  assign new_G132_ = new_G146_ | new_G148_;
  assign new_G133_ = new_G156_ | new_G155_;
  assign new_G134_ = new_G150_ | new_G149_;
  assign new_G135_ = ~new_G158_ | ~new_G157_;
  assign new_G136_ = ~new_G159_ & new_G160_;
  assign new_G137_ = new_G159_ & ~new_G160_;
  assign new_G138_ = ~G106 & G107;
  assign new_G139_ = G106 & ~G107;
  assign new_G140_ = ~new_G122_ | new_G132_;
  assign new_G141_ = new_G122_ & new_G132_;
  assign new_G142_ = ~new_G122_ & ~new_G132_;
  assign new_G143_ = new_G164_ | new_G163_;
  assign new_G144_ = G110 | new_G143_;
  assign new_G145_ = new_G168_ | new_G167_;
  assign new_G146_ = ~G110 & new_G145_;
  assign new_G147_ = new_G166_ | new_G165_;
  assign new_G148_ = G110 & new_G147_;
  assign new_G149_ = G108 & ~new_G118_;
  assign new_G150_ = ~G108 & new_G118_;
  assign new_G151_ = ~G107 | ~new_G132_;
  assign new_G152_ = new_G118_ & new_G151_;
  assign new_G153_ = ~new_G118_ & ~new_G152_;
  assign new_G154_ = new_G118_ | new_G151_;
  assign new_G155_ = ~G108 & G109;
  assign new_G156_ = G108 & ~G109;
  assign new_G157_ = new_G125_ | new_G162_;
  assign new_G158_ = ~new_G125_ & ~new_G161_;
  assign new_G159_ = G108 | new_G125_;
  assign new_G160_ = G108 | G109;
  assign new_G161_ = new_G125_ & new_G162_;
  assign new_G162_ = ~G107 | ~new_G132_;
  assign new_G163_ = new_G140_ & new_G160_;
  assign new_G164_ = ~new_G140_ & ~new_G160_;
  assign new_G165_ = new_G169_ | new_G170_;
  assign new_G166_ = ~G111 & new_G125_;
  assign new_G167_ = new_G171_ | new_G172_;
  assign new_G168_ = G111 & new_G125_;
  assign new_G169_ = ~G111 & ~new_G125_;
  assign new_G170_ = G111 & ~new_G125_;
  assign new_G171_ = G111 & ~new_G125_;
  assign new_G172_ = ~G111 & new_G125_;
  assign new_G179_ = new_G186_ & new_G185_;
  assign new_G180_ = new_G188_ | new_G187_;
  assign new_G181_ = new_G190_ | new_G189_;
  assign new_G182_ = new_G192_ & new_G191_;
  assign new_G183_ = new_G192_ & new_G193_;
  assign new_G184_ = new_G185_ | new_G194_;
  assign new_G185_ = G174 | new_G197_;
  assign new_G186_ = new_G196_ | new_G195_;
  assign new_G187_ = new_G201_ & new_G200_;
  assign new_G188_ = new_G199_ & new_G198_;
  assign new_G189_ = new_G204_ | new_G203_;
  assign new_G190_ = new_G199_ & new_G202_;
  assign new_G191_ = G174 | new_G207_;
  assign new_G192_ = new_G206_ | new_G205_;
  assign new_G193_ = new_G209_ | new_G208_;
  assign new_G194_ = ~new_G185_ & new_G211_;
  assign new_G195_ = ~new_G187_ & new_G199_;
  assign new_G196_ = new_G187_ & ~new_G199_;
  assign new_G197_ = G173 & ~G174;
  assign new_G198_ = ~new_G220_ | ~new_G221_;
  assign new_G199_ = new_G213_ | new_G215_;
  assign new_G200_ = new_G223_ | new_G222_;
  assign new_G201_ = new_G217_ | new_G216_;
  assign new_G202_ = ~new_G225_ | ~new_G224_;
  assign new_G203_ = ~new_G226_ & new_G227_;
  assign new_G204_ = new_G226_ & ~new_G227_;
  assign new_G205_ = ~G173 & G174;
  assign new_G206_ = G173 & ~G174;
  assign new_G207_ = ~new_G189_ | new_G199_;
  assign new_G208_ = new_G189_ & new_G199_;
  assign new_G209_ = ~new_G189_ & ~new_G199_;
  assign new_G210_ = new_G231_ | new_G230_;
  assign new_G211_ = G177 | new_G210_;
  assign new_G212_ = new_G235_ | new_G234_;
  assign new_G213_ = ~G177 & new_G212_;
  assign new_G214_ = new_G233_ | new_G232_;
  assign new_G215_ = G177 & new_G214_;
  assign new_G216_ = G175 & ~new_G185_;
  assign new_G217_ = ~G175 & new_G185_;
  assign new_G218_ = ~G174 | ~new_G199_;
  assign new_G219_ = new_G185_ & new_G218_;
  assign new_G220_ = ~new_G185_ & ~new_G219_;
  assign new_G221_ = new_G185_ | new_G218_;
  assign new_G222_ = ~G175 & G176;
  assign new_G223_ = G175 & ~G176;
  assign new_G224_ = new_G192_ | new_G229_;
  assign new_G225_ = ~new_G192_ & ~new_G228_;
  assign new_G226_ = G175 | new_G192_;
  assign new_G227_ = G175 | G176;
  assign new_G228_ = new_G192_ & new_G229_;
  assign new_G229_ = ~G174 | ~new_G199_;
  assign new_G230_ = new_G207_ & new_G227_;
  assign new_G231_ = ~new_G207_ & ~new_G227_;
  assign new_G232_ = new_G236_ | new_G237_;
  assign new_G233_ = ~G178 & new_G192_;
  assign new_G234_ = new_G238_ | new_G239_;
  assign new_G235_ = G178 & new_G192_;
  assign new_G236_ = ~G178 & ~new_G192_;
  assign new_G237_ = G178 & ~new_G192_;
  assign new_G238_ = G178 & ~new_G192_;
  assign new_G239_ = ~G178 & new_G192_;
  assign new_G246_ = new_G253_ & new_G252_;
  assign new_G247_ = new_G255_ | new_G254_;
  assign new_G248_ = new_G257_ | new_G256_;
  assign new_G249_ = new_G259_ & new_G258_;
  assign new_G250_ = new_G259_ & new_G260_;
  assign new_G251_ = new_G252_ | new_G261_;
  assign new_G252_ = G241 | new_G264_;
  assign new_G253_ = new_G263_ | new_G262_;
  assign new_G254_ = new_G268_ & new_G267_;
  assign new_G255_ = new_G266_ & new_G265_;
  assign new_G256_ = new_G271_ | new_G270_;
  assign new_G257_ = new_G266_ & new_G269_;
  assign new_G258_ = G241 | new_G274_;
  assign new_G259_ = new_G273_ | new_G272_;
  assign new_G260_ = new_G276_ | new_G275_;
  assign new_G261_ = ~new_G252_ & new_G278_;
  assign new_G262_ = ~new_G254_ & new_G266_;
  assign new_G263_ = new_G254_ & ~new_G266_;
  assign new_G264_ = G240 & ~G241;
  assign new_G265_ = ~new_G287_ | ~new_G288_;
  assign new_G266_ = new_G280_ | new_G282_;
  assign new_G267_ = new_G290_ | new_G289_;
  assign new_G268_ = new_G284_ | new_G283_;
  assign new_G269_ = ~new_G292_ | ~new_G291_;
  assign new_G270_ = ~new_G293_ & new_G294_;
  assign new_G271_ = new_G293_ & ~new_G294_;
  assign new_G272_ = ~G240 & G241;
  assign new_G273_ = G240 & ~G241;
  assign new_G274_ = ~new_G256_ | new_G266_;
  assign new_G275_ = new_G256_ & new_G266_;
  assign new_G276_ = ~new_G256_ & ~new_G266_;
  assign new_G277_ = new_G298_ | new_G297_;
  assign new_G278_ = G244 | new_G277_;
  assign new_G279_ = new_G302_ | new_G301_;
  assign new_G280_ = ~G244 & new_G279_;
  assign new_G281_ = new_G300_ | new_G299_;
  assign new_G282_ = G244 & new_G281_;
  assign new_G283_ = G242 & ~new_G252_;
  assign new_G284_ = ~G242 & new_G252_;
  assign new_G285_ = ~G241 | ~new_G266_;
  assign new_G286_ = new_G252_ & new_G285_;
  assign new_G287_ = ~new_G252_ & ~new_G286_;
  assign new_G288_ = new_G252_ | new_G285_;
  assign new_G289_ = ~G242 & G243;
  assign new_G290_ = G242 & ~G243;
  assign new_G291_ = new_G259_ | new_G296_;
  assign new_G292_ = ~new_G259_ & ~new_G295_;
  assign new_G293_ = G242 | new_G259_;
  assign new_G294_ = G242 | G243;
  assign new_G295_ = new_G259_ & new_G296_;
  assign new_G296_ = ~G241 | ~new_G266_;
  assign new_G297_ = new_G274_ & new_G294_;
  assign new_G298_ = ~new_G274_ & ~new_G294_;
  assign new_G299_ = new_G303_ | new_G304_;
  assign new_G300_ = ~G245 & new_G259_;
  assign new_G301_ = new_G305_ | new_G306_;
  assign new_G302_ = G245 & new_G259_;
  assign new_G303_ = ~G245 & ~new_G259_;
  assign new_G304_ = G245 & ~new_G259_;
  assign new_G305_ = G245 & ~new_G259_;
  assign new_G306_ = ~G245 & new_G259_;
  assign new_G313_ = new_G320_ & new_G319_;
  assign new_G314_ = new_G322_ | new_G321_;
  assign new_G315_ = new_G324_ | new_G323_;
  assign new_G316_ = new_G326_ & new_G325_;
  assign new_G317_ = new_G326_ & new_G327_;
  assign new_G318_ = new_G319_ | new_G328_;
  assign new_G319_ = G308 | new_G331_;
  assign new_G320_ = new_G330_ | new_G329_;
  assign new_G321_ = new_G335_ & new_G334_;
  assign new_G322_ = new_G333_ & new_G332_;
  assign new_G323_ = new_G338_ | new_G337_;
  assign new_G324_ = new_G333_ & new_G336_;
  assign new_G325_ = G308 | new_G341_;
  assign new_G326_ = new_G340_ | new_G339_;
  assign new_G327_ = new_G343_ | new_G342_;
  assign new_G328_ = ~new_G319_ & new_G345_;
  assign new_G329_ = ~new_G321_ & new_G333_;
  assign new_G330_ = new_G321_ & ~new_G333_;
  assign new_G331_ = G307 & ~G308;
  assign new_G332_ = ~new_G354_ | ~new_G355_;
  assign new_G333_ = new_G347_ | new_G349_;
  assign new_G334_ = new_G357_ | new_G356_;
  assign new_G335_ = new_G351_ | new_G350_;
  assign new_G336_ = ~new_G359_ | ~new_G358_;
  assign new_G337_ = ~new_G360_ & new_G361_;
  assign new_G338_ = new_G360_ & ~new_G361_;
  assign new_G339_ = ~G307 & G308;
  assign new_G340_ = G307 & ~G308;
  assign new_G341_ = ~new_G323_ | new_G333_;
  assign new_G342_ = new_G323_ & new_G333_;
  assign new_G343_ = ~new_G323_ & ~new_G333_;
  assign new_G344_ = new_G365_ | new_G364_;
  assign new_G345_ = G311 | new_G344_;
  assign new_G346_ = new_G369_ | new_G368_;
  assign new_G347_ = ~G311 & new_G346_;
  assign new_G348_ = new_G367_ | new_G366_;
  assign new_G349_ = G311 & new_G348_;
  assign new_G350_ = G309 & ~new_G319_;
  assign new_G351_ = ~G309 & new_G319_;
  assign new_G352_ = ~G308 | ~new_G333_;
  assign new_G353_ = new_G319_ & new_G352_;
  assign new_G354_ = ~new_G319_ & ~new_G353_;
  assign new_G355_ = new_G319_ | new_G352_;
  assign new_G356_ = ~G309 & G310;
  assign new_G357_ = G309 & ~G310;
  assign new_G358_ = new_G326_ | new_G363_;
  assign new_G359_ = ~new_G326_ & ~new_G362_;
  assign new_G360_ = G309 | new_G326_;
  assign new_G361_ = G309 | G310;
  assign new_G362_ = new_G326_ & new_G363_;
  assign new_G363_ = ~G308 | ~new_G333_;
  assign new_G364_ = new_G341_ & new_G361_;
  assign new_G365_ = ~new_G341_ & ~new_G361_;
  assign new_G366_ = new_G370_ | new_G371_;
  assign new_G367_ = ~G312 & new_G326_;
  assign new_G368_ = new_G372_ | new_G373_;
  assign new_G369_ = G312 & new_G326_;
  assign new_G370_ = ~G312 & ~new_G326_;
  assign new_G371_ = G312 & ~new_G326_;
  assign new_G372_ = G312 & ~new_G326_;
  assign new_G373_ = ~G312 & new_G326_;
  assign new_G380_ = new_G387_ & new_G386_;
  assign new_G381_ = new_G389_ | new_G388_;
  assign new_G382_ = new_G391_ | new_G390_;
  assign new_G383_ = new_G393_ & new_G392_;
  assign new_G384_ = new_G393_ & new_G394_;
  assign new_G385_ = new_G386_ | new_G395_;
  assign new_G386_ = G375 | new_G398_;
  assign new_G387_ = new_G397_ | new_G396_;
  assign new_G388_ = new_G402_ & new_G401_;
  assign new_G389_ = new_G400_ & new_G399_;
  assign new_G390_ = new_G405_ | new_G404_;
  assign new_G391_ = new_G400_ & new_G403_;
  assign new_G392_ = G375 | new_G408_;
  assign new_G393_ = new_G407_ | new_G406_;
  assign new_G394_ = new_G410_ | new_G409_;
  assign new_G395_ = ~new_G386_ & new_G412_;
  assign new_G396_ = ~new_G388_ & new_G400_;
  assign new_G397_ = new_G388_ & ~new_G400_;
  assign new_G398_ = G374 & ~G375;
  assign new_G399_ = ~new_G421_ | ~new_G422_;
  assign new_G400_ = new_G414_ | new_G416_;
  assign new_G401_ = new_G424_ | new_G423_;
  assign new_G402_ = new_G418_ | new_G417_;
  assign new_G403_ = ~new_G426_ | ~new_G425_;
  assign new_G404_ = ~new_G427_ & new_G428_;
  assign new_G405_ = new_G427_ & ~new_G428_;
  assign new_G406_ = ~G374 & G375;
  assign new_G407_ = G374 & ~G375;
  assign new_G408_ = ~new_G390_ | new_G400_;
  assign new_G409_ = new_G390_ & new_G400_;
  assign new_G410_ = ~new_G390_ & ~new_G400_;
  assign new_G411_ = new_G432_ | new_G431_;
  assign new_G412_ = G378 | new_G411_;
  assign new_G413_ = new_G436_ | new_G435_;
  assign new_G414_ = ~G378 & new_G413_;
  assign new_G415_ = new_G434_ | new_G433_;
  assign new_G416_ = G378 & new_G415_;
  assign new_G417_ = G376 & ~new_G386_;
  assign new_G418_ = ~G376 & new_G386_;
  assign new_G419_ = ~G375 | ~new_G400_;
  assign new_G420_ = new_G386_ & new_G419_;
  assign new_G421_ = ~new_G386_ & ~new_G420_;
  assign new_G422_ = new_G386_ | new_G419_;
  assign new_G423_ = ~G376 & G377;
  assign new_G424_ = G376 & ~G377;
  assign new_G425_ = new_G393_ | new_G430_;
  assign new_G426_ = ~new_G393_ & ~new_G429_;
  assign new_G427_ = G376 | new_G393_;
  assign new_G428_ = G376 | G377;
  assign new_G429_ = new_G393_ & new_G430_;
  assign new_G430_ = ~G375 | ~new_G400_;
  assign new_G431_ = new_G408_ & new_G428_;
  assign new_G432_ = ~new_G408_ & ~new_G428_;
  assign new_G433_ = new_G437_ | new_G438_;
  assign new_G434_ = ~G379 & new_G393_;
  assign new_G435_ = new_G439_ | new_G440_;
  assign new_G436_ = G379 & new_G393_;
  assign new_G437_ = ~G379 & ~new_G393_;
  assign new_G438_ = G379 & ~new_G393_;
  assign new_G439_ = G379 & ~new_G393_;
  assign new_G440_ = ~G379 & new_G393_;
  assign new_G447_ = new_G454_ & new_G453_;
  assign new_G448_ = new_G456_ | new_G455_;
  assign new_G449_ = new_G458_ | new_G457_;
  assign new_G450_ = new_G460_ & new_G459_;
  assign new_G451_ = new_G460_ & new_G461_;
  assign new_G452_ = new_G453_ | new_G462_;
  assign new_G453_ = G442 | new_G465_;
  assign new_G454_ = new_G464_ | new_G463_;
  assign new_G455_ = new_G469_ & new_G468_;
  assign new_G456_ = new_G467_ & new_G466_;
  assign new_G457_ = new_G472_ | new_G471_;
  assign new_G458_ = new_G467_ & new_G470_;
  assign new_G459_ = G442 | new_G475_;
  assign new_G460_ = new_G474_ | new_G473_;
  assign new_G461_ = new_G477_ | new_G476_;
  assign new_G462_ = ~new_G453_ & new_G479_;
  assign new_G463_ = ~new_G455_ & new_G467_;
  assign new_G464_ = new_G455_ & ~new_G467_;
  assign new_G465_ = G441 & ~G442;
  assign new_G466_ = ~new_G488_ | ~new_G489_;
  assign new_G467_ = new_G481_ | new_G483_;
  assign new_G468_ = new_G491_ | new_G490_;
  assign new_G469_ = new_G485_ | new_G484_;
  assign new_G470_ = ~new_G493_ | ~new_G492_;
  assign new_G471_ = ~new_G494_ & new_G495_;
  assign new_G472_ = new_G494_ & ~new_G495_;
  assign new_G473_ = ~G441 & G442;
  assign new_G474_ = G441 & ~G442;
  assign new_G475_ = ~new_G457_ | new_G467_;
  assign new_G476_ = new_G457_ & new_G467_;
  assign new_G477_ = ~new_G457_ & ~new_G467_;
  assign new_G478_ = new_G499_ | new_G498_;
  assign new_G479_ = G445 | new_G478_;
  assign new_G480_ = new_G503_ | new_G502_;
  assign new_G481_ = ~G445 & new_G480_;
  assign new_G482_ = new_G501_ | new_G500_;
  assign new_G483_ = G445 & new_G482_;
  assign new_G484_ = G443 & ~new_G453_;
  assign new_G485_ = ~G443 & new_G453_;
  assign new_G486_ = ~G442 | ~new_G467_;
  assign new_G487_ = new_G453_ & new_G486_;
  assign new_G488_ = ~new_G453_ & ~new_G487_;
  assign new_G489_ = new_G453_ | new_G486_;
  assign new_G490_ = ~G443 & G444;
  assign new_G491_ = G443 & ~G444;
  assign new_G492_ = new_G460_ | new_G497_;
  assign new_G493_ = ~new_G460_ & ~new_G496_;
  assign new_G494_ = G443 | new_G460_;
  assign new_G495_ = G443 | G444;
  assign new_G496_ = new_G460_ & new_G497_;
  assign new_G497_ = ~G442 | ~new_G467_;
  assign new_G498_ = new_G475_ & new_G495_;
  assign new_G499_ = ~new_G475_ & ~new_G495_;
  assign new_G500_ = new_G504_ | new_G505_;
  assign new_G501_ = ~G446 & new_G460_;
  assign new_G502_ = new_G506_ | new_G507_;
  assign new_G503_ = G446 & new_G460_;
  assign new_G504_ = ~G446 & ~new_G460_;
  assign new_G505_ = G446 & ~new_G460_;
  assign new_G506_ = G446 & ~new_G460_;
  assign new_G507_ = ~G446 & new_G460_;
  assign new_G514_ = new_G521_ & new_G520_;
  assign new_G515_ = new_G523_ | new_G522_;
  assign new_G516_ = new_G525_ | new_G524_;
  assign new_G517_ = new_G527_ & new_G526_;
  assign new_G518_ = new_G527_ & new_G528_;
  assign new_G519_ = new_G520_ | new_G529_;
  assign new_G520_ = G509 | new_G532_;
  assign new_G521_ = new_G531_ | new_G530_;
  assign new_G522_ = new_G536_ & new_G535_;
  assign new_G523_ = new_G534_ & new_G533_;
  assign new_G524_ = new_G539_ | new_G538_;
  assign new_G525_ = new_G534_ & new_G537_;
  assign new_G526_ = G509 | new_G542_;
  assign new_G527_ = new_G541_ | new_G540_;
  assign new_G528_ = new_G544_ | new_G543_;
  assign new_G529_ = ~new_G520_ & new_G546_;
  assign new_G530_ = ~new_G522_ & new_G534_;
  assign new_G531_ = new_G522_ & ~new_G534_;
  assign new_G532_ = G508 & ~G509;
  assign new_G533_ = ~new_G555_ | ~new_G556_;
  assign new_G534_ = new_G548_ | new_G550_;
  assign new_G535_ = new_G558_ | new_G557_;
  assign new_G536_ = new_G552_ | new_G551_;
  assign new_G537_ = ~new_G560_ | ~new_G559_;
  assign new_G538_ = ~new_G561_ & new_G562_;
  assign new_G539_ = new_G561_ & ~new_G562_;
  assign new_G540_ = ~G508 & G509;
  assign new_G541_ = G508 & ~G509;
  assign new_G542_ = ~new_G524_ | new_G534_;
  assign new_G543_ = new_G524_ & new_G534_;
  assign new_G544_ = ~new_G524_ & ~new_G534_;
  assign new_G545_ = new_G566_ | new_G565_;
  assign new_G546_ = G512 | new_G545_;
  assign new_G547_ = new_G570_ | new_G569_;
  assign new_G548_ = ~G512 & new_G547_;
  assign new_G549_ = new_G568_ | new_G567_;
  assign new_G550_ = G512 & new_G549_;
  assign new_G551_ = G510 & ~new_G520_;
  assign new_G552_ = ~G510 & new_G520_;
  assign new_G553_ = ~G509 | ~new_G534_;
  assign new_G554_ = new_G520_ & new_G553_;
  assign new_G555_ = ~new_G520_ & ~new_G554_;
  assign new_G556_ = new_G520_ | new_G553_;
  assign new_G557_ = ~G510 & G511;
  assign new_G558_ = G510 & ~G511;
  assign new_G559_ = new_G527_ | new_G564_;
  assign new_G560_ = ~new_G527_ & ~new_G563_;
  assign new_G561_ = G510 | new_G527_;
  assign new_G562_ = G510 | G511;
  assign new_G563_ = new_G527_ & new_G564_;
  assign new_G564_ = ~G509 | ~new_G534_;
  assign new_G565_ = new_G542_ & new_G562_;
  assign new_G566_ = ~new_G542_ & ~new_G562_;
  assign new_G567_ = new_G571_ | new_G572_;
  assign new_G568_ = ~G513 & new_G527_;
  assign new_G569_ = new_G573_ | new_G574_;
  assign new_G570_ = G513 & new_G527_;
  assign new_G571_ = ~G513 & ~new_G527_;
  assign new_G572_ = G513 & ~new_G527_;
  assign new_G573_ = G513 & ~new_G527_;
  assign new_G574_ = ~G513 & new_G527_;
  assign new_G581_ = new_G588_ & new_G587_;
  assign new_G582_ = new_G590_ | new_G589_;
  assign new_G583_ = new_G592_ | new_G591_;
  assign new_G584_ = new_G594_ & new_G593_;
  assign new_G585_ = new_G594_ & new_G595_;
  assign new_G586_ = new_G587_ | new_G596_;
  assign new_G587_ = G576 | new_G599_;
  assign new_G588_ = new_G598_ | new_G597_;
  assign new_G589_ = new_G603_ & new_G602_;
  assign new_G590_ = new_G601_ & new_G600_;
  assign new_G591_ = new_G606_ | new_G605_;
  assign new_G592_ = new_G601_ & new_G604_;
  assign new_G593_ = G576 | new_G609_;
  assign new_G594_ = new_G608_ | new_G607_;
  assign new_G595_ = new_G611_ | new_G610_;
  assign new_G596_ = ~new_G587_ & new_G613_;
  assign new_G597_ = ~new_G589_ & new_G601_;
  assign new_G598_ = new_G589_ & ~new_G601_;
  assign new_G599_ = G575 & ~G576;
  assign new_G600_ = ~new_G622_ | ~new_G623_;
  assign new_G601_ = new_G615_ | new_G617_;
  assign new_G602_ = new_G625_ | new_G624_;
  assign new_G603_ = new_G619_ | new_G618_;
  assign new_G604_ = ~new_G627_ | ~new_G626_;
  assign new_G605_ = ~new_G628_ & new_G629_;
  assign new_G606_ = new_G628_ & ~new_G629_;
  assign new_G607_ = ~G575 & G576;
  assign new_G608_ = G575 & ~G576;
  assign new_G609_ = ~new_G591_ | new_G601_;
  assign new_G610_ = new_G591_ & new_G601_;
  assign new_G611_ = ~new_G591_ & ~new_G601_;
  assign new_G612_ = new_G633_ | new_G632_;
  assign new_G613_ = G579 | new_G612_;
  assign new_G614_ = new_G637_ | new_G636_;
  assign new_G615_ = ~G579 & new_G614_;
  assign new_G616_ = new_G635_ | new_G634_;
  assign new_G617_ = G579 & new_G616_;
  assign new_G618_ = G577 & ~new_G587_;
  assign new_G619_ = ~G577 & new_G587_;
  assign new_G620_ = ~G576 | ~new_G601_;
  assign new_G621_ = new_G587_ & new_G620_;
  assign new_G622_ = ~new_G587_ & ~new_G621_;
  assign new_G623_ = new_G587_ | new_G620_;
  assign new_G624_ = ~G577 & G578;
  assign new_G625_ = G577 & ~G578;
  assign new_G626_ = new_G594_ | new_G631_;
  assign new_G627_ = ~new_G594_ & ~new_G630_;
  assign new_G628_ = G577 | new_G594_;
  assign new_G629_ = G577 | G578;
  assign new_G630_ = new_G594_ & new_G631_;
  assign new_G631_ = ~G576 | ~new_G601_;
  assign new_G632_ = new_G609_ & new_G629_;
  assign new_G633_ = ~new_G609_ & ~new_G629_;
  assign new_G634_ = new_G638_ | new_G639_;
  assign new_G635_ = ~G580 & new_G594_;
  assign new_G636_ = new_G640_ | new_G641_;
  assign new_G637_ = G580 & new_G594_;
  assign new_G638_ = ~G580 & ~new_G594_;
  assign new_G639_ = G580 & ~new_G594_;
  assign new_G640_ = G580 & ~new_G594_;
  assign new_G641_ = ~G580 & new_G594_;
  assign new_G648_ = new_G655_ & new_G654_;
  assign new_G649_ = new_G657_ | new_G656_;
  assign new_G650_ = new_G659_ | new_G658_;
  assign new_G651_ = new_G661_ & new_G660_;
  assign new_G652_ = new_G661_ & new_G662_;
  assign new_G653_ = new_G654_ | new_G663_;
  assign new_G654_ = G643 | new_G666_;
  assign new_G655_ = new_G665_ | new_G664_;
  assign new_G656_ = new_G670_ & new_G669_;
  assign new_G657_ = new_G668_ & new_G667_;
  assign new_G658_ = new_G673_ | new_G672_;
  assign new_G659_ = new_G668_ & new_G671_;
  assign new_G660_ = G643 | new_G676_;
  assign new_G661_ = new_G675_ | new_G674_;
  assign new_G662_ = new_G678_ | new_G677_;
  assign new_G663_ = ~new_G654_ & new_G680_;
  assign new_G664_ = ~new_G656_ & new_G668_;
  assign new_G665_ = new_G656_ & ~new_G668_;
  assign new_G666_ = G642 & ~G643;
  assign new_G667_ = ~new_G689_ | ~new_G690_;
  assign new_G668_ = new_G682_ | new_G684_;
  assign new_G669_ = new_G692_ | new_G691_;
  assign new_G670_ = new_G686_ | new_G685_;
  assign new_G671_ = ~new_G694_ | ~new_G693_;
  assign new_G672_ = ~new_G695_ & new_G696_;
  assign new_G673_ = new_G695_ & ~new_G696_;
  assign new_G674_ = ~G642 & G643;
  assign new_G675_ = G642 & ~G643;
  assign new_G676_ = ~new_G658_ | new_G668_;
  assign new_G677_ = new_G658_ & new_G668_;
  assign new_G678_ = ~new_G658_ & ~new_G668_;
  assign new_G679_ = new_G700_ | new_G699_;
  assign new_G680_ = G646 | new_G679_;
  assign new_G681_ = new_G704_ | new_G703_;
  assign new_G682_ = ~G646 & new_G681_;
  assign new_G683_ = new_G702_ | new_G701_;
  assign new_G684_ = G646 & new_G683_;
  assign new_G685_ = G644 & ~new_G654_;
  assign new_G686_ = ~G644 & new_G654_;
  assign new_G687_ = ~G643 | ~new_G668_;
  assign new_G688_ = new_G654_ & new_G687_;
  assign new_G689_ = ~new_G654_ & ~new_G688_;
  assign new_G690_ = new_G654_ | new_G687_;
  assign new_G691_ = ~G644 & G645;
  assign new_G692_ = G644 & ~G645;
  assign new_G693_ = new_G661_ | new_G698_;
  assign new_G694_ = ~new_G661_ & ~new_G697_;
  assign new_G695_ = G644 | new_G661_;
  assign new_G696_ = G644 | G645;
  assign new_G697_ = new_G661_ & new_G698_;
  assign new_G698_ = ~G643 | ~new_G668_;
  assign new_G699_ = new_G676_ & new_G696_;
  assign new_G700_ = ~new_G676_ & ~new_G696_;
  assign new_G701_ = new_G705_ | new_G706_;
  assign new_G702_ = ~G647 & new_G661_;
  assign new_G703_ = new_G707_ | new_G708_;
  assign new_G704_ = G647 & new_G661_;
  assign new_G705_ = ~G647 & ~new_G661_;
  assign new_G706_ = G647 & ~new_G661_;
  assign new_G707_ = G647 & ~new_G661_;
  assign new_G708_ = ~G647 & new_G661_;
  assign new_G715_ = new_G722_ & new_G721_;
  assign new_G716_ = new_G724_ | new_G723_;
  assign new_G717_ = new_G726_ | new_G725_;
  assign new_G718_ = new_G728_ & new_G727_;
  assign new_G719_ = new_G728_ & new_G729_;
  assign new_G720_ = new_G721_ | new_G730_;
  assign new_G721_ = G710 | new_G733_;
  assign new_G722_ = new_G732_ | new_G731_;
  assign new_G723_ = new_G737_ & new_G736_;
  assign new_G724_ = new_G735_ & new_G734_;
  assign new_G725_ = new_G740_ | new_G739_;
  assign new_G726_ = new_G735_ & new_G738_;
  assign new_G727_ = G710 | new_G743_;
  assign new_G728_ = new_G742_ | new_G741_;
  assign new_G729_ = new_G745_ | new_G744_;
  assign new_G730_ = ~new_G721_ & new_G747_;
  assign new_G731_ = ~new_G723_ & new_G735_;
  assign new_G732_ = new_G723_ & ~new_G735_;
  assign new_G733_ = G709 & ~G710;
  assign new_G734_ = ~new_G756_ | ~new_G757_;
  assign new_G735_ = new_G749_ | new_G751_;
  assign new_G736_ = new_G759_ | new_G758_;
  assign new_G737_ = new_G753_ | new_G752_;
  assign new_G738_ = ~new_G761_ | ~new_G760_;
  assign new_G739_ = ~new_G762_ & new_G763_;
  assign new_G740_ = new_G762_ & ~new_G763_;
  assign new_G741_ = ~G709 & G710;
  assign new_G742_ = G709 & ~G710;
  assign new_G743_ = ~new_G725_ | new_G735_;
  assign new_G744_ = new_G725_ & new_G735_;
  assign new_G745_ = ~new_G725_ & ~new_G735_;
  assign new_G746_ = new_G767_ | new_G766_;
  assign new_G747_ = G713 | new_G746_;
  assign new_G748_ = new_G771_ | new_G770_;
  assign new_G749_ = ~G713 & new_G748_;
  assign new_G750_ = new_G769_ | new_G768_;
  assign new_G751_ = G713 & new_G750_;
  assign new_G752_ = G711 & ~new_G721_;
  assign new_G753_ = ~G711 & new_G721_;
  assign new_G754_ = ~G710 | ~new_G735_;
  assign new_G755_ = new_G721_ & new_G754_;
  assign new_G756_ = ~new_G721_ & ~new_G755_;
  assign new_G757_ = new_G721_ | new_G754_;
  assign new_G758_ = ~G711 & G712;
  assign new_G759_ = G711 & ~G712;
  assign new_G760_ = new_G728_ | new_G765_;
  assign new_G761_ = ~new_G728_ & ~new_G764_;
  assign new_G762_ = G711 | new_G728_;
  assign new_G763_ = G711 | G712;
  assign new_G764_ = new_G728_ & new_G765_;
  assign new_G765_ = ~G710 | ~new_G735_;
  assign new_G766_ = new_G743_ & new_G763_;
  assign new_G767_ = ~new_G743_ & ~new_G763_;
  assign new_G768_ = new_G772_ | new_G773_;
  assign new_G769_ = ~G714 & new_G728_;
  assign new_G770_ = new_G774_ | new_G775_;
  assign new_G771_ = G714 & new_G728_;
  assign new_G772_ = ~G714 & ~new_G728_;
  assign new_G773_ = G714 & ~new_G728_;
  assign new_G774_ = G714 & ~new_G728_;
  assign new_G775_ = ~G714 & new_G728_;
  assign new_G782_ = new_G789_ & new_G788_;
  assign new_G783_ = new_G791_ | new_G790_;
  assign new_G784_ = new_G793_ | new_G792_;
  assign new_G785_ = new_G795_ & new_G794_;
  assign new_G786_ = new_G795_ & new_G796_;
  assign new_G787_ = new_G788_ | new_G797_;
  assign new_G788_ = G777 | new_G800_;
  assign new_G789_ = new_G799_ | new_G798_;
  assign new_G790_ = new_G804_ & new_G803_;
  assign new_G791_ = new_G802_ & new_G801_;
  assign new_G792_ = new_G807_ | new_G806_;
  assign new_G793_ = new_G802_ & new_G805_;
  assign new_G794_ = G777 | new_G810_;
  assign new_G795_ = new_G809_ | new_G808_;
  assign new_G796_ = new_G812_ | new_G811_;
  assign new_G797_ = ~new_G788_ & new_G814_;
  assign new_G798_ = ~new_G790_ & new_G802_;
  assign new_G799_ = new_G790_ & ~new_G802_;
  assign new_G800_ = G776 & ~G777;
  assign new_G801_ = ~new_G823_ | ~new_G824_;
  assign new_G802_ = new_G816_ | new_G818_;
  assign new_G803_ = new_G826_ | new_G825_;
  assign new_G804_ = new_G820_ | new_G819_;
  assign new_G805_ = ~new_G828_ | ~new_G827_;
  assign new_G806_ = ~new_G829_ & new_G830_;
  assign new_G807_ = new_G829_ & ~new_G830_;
  assign new_G808_ = ~G776 & G777;
  assign new_G809_ = G776 & ~G777;
  assign new_G810_ = ~new_G792_ | new_G802_;
  assign new_G811_ = new_G792_ & new_G802_;
  assign new_G812_ = ~new_G792_ & ~new_G802_;
  assign new_G813_ = new_G834_ | new_G833_;
  assign new_G814_ = G780 | new_G813_;
  assign new_G815_ = new_G838_ | new_G837_;
  assign new_G816_ = ~G780 & new_G815_;
  assign new_G817_ = new_G836_ | new_G835_;
  assign new_G818_ = G780 & new_G817_;
  assign new_G819_ = G778 & ~new_G788_;
  assign new_G820_ = ~G778 & new_G788_;
  assign new_G821_ = ~G777 | ~new_G802_;
  assign new_G822_ = new_G788_ & new_G821_;
  assign new_G823_ = ~new_G788_ & ~new_G822_;
  assign new_G824_ = new_G788_ | new_G821_;
  assign new_G825_ = ~G778 & G779;
  assign new_G826_ = G778 & ~G779;
  assign new_G827_ = new_G795_ | new_G832_;
  assign new_G828_ = ~new_G795_ & ~new_G831_;
  assign new_G829_ = G778 | new_G795_;
  assign new_G830_ = G778 | G779;
  assign new_G831_ = new_G795_ & new_G832_;
  assign new_G832_ = ~G777 | ~new_G802_;
  assign new_G833_ = new_G810_ & new_G830_;
  assign new_G834_ = ~new_G810_ & ~new_G830_;
  assign new_G835_ = new_G839_ | new_G840_;
  assign new_G836_ = ~G781 & new_G795_;
  assign new_G837_ = new_G841_ | new_G842_;
  assign new_G838_ = G781 & new_G795_;
  assign new_G839_ = ~G781 & ~new_G795_;
  assign new_G840_ = G781 & ~new_G795_;
  assign new_G841_ = G781 & ~new_G795_;
  assign new_G842_ = ~G781 & new_G795_;
  assign new_G849_ = new_G856_ & new_G855_;
  assign new_G850_ = new_G858_ | new_G857_;
  assign new_G851_ = new_G860_ | new_G859_;
  assign new_G852_ = new_G862_ & new_G861_;
  assign new_G853_ = new_G862_ & new_G863_;
  assign new_G854_ = new_G855_ | new_G864_;
  assign new_G855_ = G844 | new_G867_;
  assign new_G856_ = new_G866_ | new_G865_;
  assign new_G857_ = new_G871_ & new_G870_;
  assign new_G858_ = new_G869_ & new_G868_;
  assign new_G859_ = new_G874_ | new_G873_;
  assign new_G860_ = new_G869_ & new_G872_;
  assign new_G861_ = G844 | new_G877_;
  assign new_G862_ = new_G876_ | new_G875_;
  assign new_G863_ = new_G879_ | new_G878_;
  assign new_G864_ = ~new_G855_ & new_G881_;
  assign new_G865_ = ~new_G857_ & new_G869_;
  assign new_G866_ = new_G857_ & ~new_G869_;
  assign new_G867_ = G843 & ~G844;
  assign new_G868_ = ~new_G890_ | ~new_G891_;
  assign new_G869_ = new_G883_ | new_G885_;
  assign new_G870_ = new_G893_ | new_G892_;
  assign new_G871_ = new_G887_ | new_G886_;
  assign new_G872_ = ~new_G895_ | ~new_G894_;
  assign new_G873_ = ~new_G896_ & new_G897_;
  assign new_G874_ = new_G896_ & ~new_G897_;
  assign new_G875_ = ~G843 & G844;
  assign new_G876_ = G843 & ~G844;
  assign new_G877_ = ~new_G859_ | new_G869_;
  assign new_G878_ = new_G859_ & new_G869_;
  assign new_G879_ = ~new_G859_ & ~new_G869_;
  assign new_G880_ = new_G901_ | new_G900_;
  assign new_G881_ = G847 | new_G880_;
  assign new_G882_ = new_G905_ | new_G904_;
  assign new_G883_ = ~G847 & new_G882_;
  assign new_G884_ = new_G903_ | new_G902_;
  assign new_G885_ = G847 & new_G884_;
  assign new_G886_ = G845 & ~new_G855_;
  assign new_G887_ = ~G845 & new_G855_;
  assign new_G888_ = ~G844 | ~new_G869_;
  assign new_G889_ = new_G855_ & new_G888_;
  assign new_G890_ = ~new_G855_ & ~new_G889_;
  assign new_G891_ = new_G855_ | new_G888_;
  assign new_G892_ = ~G845 & G846;
  assign new_G893_ = G845 & ~G846;
  assign new_G894_ = new_G862_ | new_G899_;
  assign new_G895_ = ~new_G862_ & ~new_G898_;
  assign new_G896_ = G845 | new_G862_;
  assign new_G897_ = G845 | G846;
  assign new_G898_ = new_G862_ & new_G899_;
  assign new_G899_ = ~G844 | ~new_G869_;
  assign new_G900_ = new_G877_ & new_G897_;
  assign new_G901_ = ~new_G877_ & ~new_G897_;
  assign new_G902_ = new_G906_ | new_G907_;
  assign new_G903_ = ~G848 & new_G862_;
  assign new_G904_ = new_G908_ | new_G909_;
  assign new_G905_ = G848 & new_G862_;
  assign new_G906_ = ~G848 & ~new_G862_;
  assign new_G907_ = G848 & ~new_G862_;
  assign new_G908_ = G848 & ~new_G862_;
  assign new_G909_ = ~G848 & new_G862_;
  assign new_G916_ = new_G923_ & new_G922_;
  assign new_G917_ = new_G925_ | new_G924_;
  assign new_G918_ = new_G927_ | new_G926_;
  assign new_G919_ = new_G929_ & new_G928_;
  assign new_G920_ = new_G929_ & new_G930_;
  assign new_G921_ = new_G922_ | new_G931_;
  assign new_G922_ = G911 | new_G934_;
  assign new_G923_ = new_G933_ | new_G932_;
  assign new_G924_ = new_G938_ & new_G937_;
  assign new_G925_ = new_G936_ & new_G935_;
  assign new_G926_ = new_G941_ | new_G940_;
  assign new_G927_ = new_G936_ & new_G939_;
  assign new_G928_ = G911 | new_G944_;
  assign new_G929_ = new_G943_ | new_G942_;
  assign new_G930_ = new_G946_ | new_G945_;
  assign new_G931_ = ~new_G922_ & new_G948_;
  assign new_G932_ = ~new_G924_ & new_G936_;
  assign new_G933_ = new_G924_ & ~new_G936_;
  assign new_G934_ = G910 & ~G911;
  assign new_G935_ = ~new_G957_ | ~new_G958_;
  assign new_G936_ = new_G950_ | new_G952_;
  assign new_G937_ = new_G960_ | new_G959_;
  assign new_G938_ = new_G954_ | new_G953_;
  assign new_G939_ = ~new_G962_ | ~new_G961_;
  assign new_G940_ = ~new_G963_ & new_G964_;
  assign new_G941_ = new_G963_ & ~new_G964_;
  assign new_G942_ = ~G910 & G911;
  assign new_G943_ = G910 & ~G911;
  assign new_G944_ = ~new_G926_ | new_G936_;
  assign new_G945_ = new_G926_ & new_G936_;
  assign new_G946_ = ~new_G926_ & ~new_G936_;
  assign new_G947_ = new_G968_ | new_G967_;
  assign new_G948_ = G914 | new_G947_;
  assign new_G949_ = new_G972_ | new_G971_;
  assign new_G950_ = ~G914 & new_G949_;
  assign new_G951_ = new_G970_ | new_G969_;
  assign new_G952_ = G914 & new_G951_;
  assign new_G953_ = G912 & ~new_G922_;
  assign new_G954_ = ~G912 & new_G922_;
  assign new_G955_ = ~G911 | ~new_G936_;
  assign new_G956_ = new_G922_ & new_G955_;
  assign new_G957_ = ~new_G922_ & ~new_G956_;
  assign new_G958_ = new_G922_ | new_G955_;
  assign new_G959_ = ~G912 & G913;
  assign new_G960_ = G912 & ~G913;
  assign new_G961_ = new_G929_ | new_G966_;
  assign new_G962_ = ~new_G929_ & ~new_G965_;
  assign new_G963_ = G912 | new_G929_;
  assign new_G964_ = G912 | G913;
  assign new_G965_ = new_G929_ & new_G966_;
  assign new_G966_ = ~G911 | ~new_G936_;
  assign new_G967_ = new_G944_ & new_G964_;
  assign new_G968_ = ~new_G944_ & ~new_G964_;
  assign new_G969_ = new_G973_ | new_G974_;
  assign new_G970_ = ~G915 & new_G929_;
  assign new_G971_ = new_G975_ | new_G976_;
  assign new_G972_ = G915 & new_G929_;
  assign new_G973_ = ~G915 & ~new_G929_;
  assign new_G974_ = G915 & ~new_G929_;
  assign new_G975_ = G915 & ~new_G929_;
  assign new_G976_ = ~G915 & new_G929_;
  assign new_G983_ = new_G990_ & new_G989_;
  assign new_G984_ = new_G992_ | new_G991_;
  assign new_G985_ = new_G994_ | new_G993_;
  assign new_G986_ = new_G996_ & new_G995_;
  assign new_G987_ = new_G996_ & new_G997_;
  assign new_G988_ = new_G989_ | new_G998_;
  assign new_G989_ = G978 | new_G1001_;
  assign new_G990_ = new_G1000_ | new_G999_;
  assign new_G991_ = new_G1005_ & new_G1004_;
  assign new_G992_ = new_G1003_ & new_G1002_;
  assign new_G993_ = new_G1008_ | new_G1007_;
  assign new_G994_ = new_G1003_ & new_G1006_;
  assign new_G995_ = G978 | new_G1011_;
  assign new_G996_ = new_G1010_ | new_G1009_;
  assign new_G997_ = new_G1013_ | new_G1012_;
  assign new_G998_ = ~new_G989_ & new_G1015_;
  assign new_G999_ = ~new_G991_ & new_G1003_;
  assign new_G1000_ = new_G991_ & ~new_G1003_;
  assign new_G1001_ = G977 & ~G978;
  assign new_G1002_ = ~new_G1024_ | ~new_G1025_;
  assign new_G1003_ = new_G1017_ | new_G1019_;
  assign new_G1004_ = new_G1027_ | new_G1026_;
  assign new_G1005_ = new_G1021_ | new_G1020_;
  assign new_G1006_ = ~new_G1029_ | ~new_G1028_;
  assign new_G1007_ = ~new_G1030_ & new_G1031_;
  assign new_G1008_ = new_G1030_ & ~new_G1031_;
  assign new_G1009_ = ~G977 & G978;
  assign new_G1010_ = G977 & ~G978;
  assign new_G1011_ = ~new_G993_ | new_G1003_;
  assign new_G1012_ = new_G993_ & new_G1003_;
  assign new_G1013_ = ~new_G993_ & ~new_G1003_;
  assign new_G1014_ = new_G1035_ | new_G1034_;
  assign new_G1015_ = G981 | new_G1014_;
  assign new_G1016_ = new_G1039_ | new_G1038_;
  assign new_G1017_ = ~G981 & new_G1016_;
  assign new_G1018_ = new_G1037_ | new_G1036_;
  assign new_G1019_ = G981 & new_G1018_;
  assign new_G1020_ = G979 & ~new_G989_;
  assign new_G1021_ = ~G979 & new_G989_;
  assign new_G1022_ = ~G978 | ~new_G1003_;
  assign new_G1023_ = new_G989_ & new_G1022_;
  assign new_G1024_ = ~new_G989_ & ~new_G1023_;
  assign new_G1025_ = new_G989_ | new_G1022_;
  assign new_G1026_ = ~G979 & G980;
  assign new_G1027_ = G979 & ~G980;
  assign new_G1028_ = new_G996_ | new_G1033_;
  assign new_G1029_ = ~new_G996_ & ~new_G1032_;
  assign new_G1030_ = G979 | new_G996_;
  assign new_G1031_ = G979 | G980;
  assign new_G1032_ = new_G996_ & new_G1033_;
  assign new_G1033_ = ~G978 | ~new_G1003_;
  assign new_G1034_ = new_G1011_ & new_G1031_;
  assign new_G1035_ = ~new_G1011_ & ~new_G1031_;
  assign new_G1036_ = new_G1040_ | new_G1041_;
  assign new_G1037_ = ~G982 & new_G996_;
  assign new_G1038_ = new_G1042_ | new_G1043_;
  assign new_G1039_ = G982 & new_G996_;
  assign new_G1040_ = ~G982 & ~new_G996_;
  assign new_G1041_ = G982 & ~new_G996_;
  assign new_G1042_ = G982 & ~new_G996_;
  assign new_G1043_ = ~G982 & new_G996_;
  assign new_G1050_ = new_G1057_ & new_G1056_;
  assign new_G1051_ = new_G1059_ | new_G1058_;
  assign new_G1052_ = new_G1061_ | new_G1060_;
  assign new_G1053_ = new_G1063_ & new_G1062_;
  assign new_G1054_ = new_G1063_ & new_G1064_;
  assign new_G1055_ = new_G1056_ | new_G1065_;
  assign new_G1056_ = G1045 | new_G1068_;
  assign new_G1057_ = new_G1067_ | new_G1066_;
  assign new_G1058_ = new_G1072_ & new_G1071_;
  assign new_G1059_ = new_G1070_ & new_G1069_;
  assign new_G1060_ = new_G1075_ | new_G1074_;
  assign new_G1061_ = new_G1070_ & new_G1073_;
  assign new_G1062_ = G1045 | new_G1078_;
  assign new_G1063_ = new_G1077_ | new_G1076_;
  assign new_G1064_ = new_G1080_ | new_G1079_;
  assign new_G1065_ = ~new_G1056_ & new_G1082_;
  assign new_G1066_ = ~new_G1058_ & new_G1070_;
  assign new_G1067_ = new_G1058_ & ~new_G1070_;
  assign new_G1068_ = G1044 & ~G1045;
  assign new_G1069_ = ~new_G1091_ | ~new_G1092_;
  assign new_G1070_ = new_G1084_ | new_G1086_;
  assign new_G1071_ = new_G1094_ | new_G1093_;
  assign new_G1072_ = new_G1088_ | new_G1087_;
  assign new_G1073_ = ~new_G1096_ | ~new_G1095_;
  assign new_G1074_ = ~new_G1097_ & new_G1098_;
  assign new_G1075_ = new_G1097_ & ~new_G1098_;
  assign new_G1076_ = ~G1044 & G1045;
  assign new_G1077_ = G1044 & ~G1045;
  assign new_G1078_ = ~new_G1060_ | new_G1070_;
  assign new_G1079_ = new_G1060_ & new_G1070_;
  assign new_G1080_ = ~new_G1060_ & ~new_G1070_;
  assign new_G1081_ = new_G1102_ | new_G1101_;
  assign new_G1082_ = G1048 | new_G1081_;
  assign new_G1083_ = new_G1106_ | new_G1105_;
  assign new_G1084_ = ~G1048 & new_G1083_;
  assign new_G1085_ = new_G1104_ | new_G1103_;
  assign new_G1086_ = G1048 & new_G1085_;
  assign new_G1087_ = G1046 & ~new_G1056_;
  assign new_G1088_ = ~G1046 & new_G1056_;
  assign new_G1089_ = ~G1045 | ~new_G1070_;
  assign new_G1090_ = new_G1056_ & new_G1089_;
  assign new_G1091_ = ~new_G1056_ & ~new_G1090_;
  assign new_G1092_ = new_G1056_ | new_G1089_;
  assign new_G1093_ = ~G1046 & G1047;
  assign new_G1094_ = G1046 & ~G1047;
  assign new_G1095_ = new_G1063_ | new_G1100_;
  assign new_G1096_ = ~new_G1063_ & ~new_G1099_;
  assign new_G1097_ = G1046 | new_G1063_;
  assign new_G1098_ = G1046 | G1047;
  assign new_G1099_ = new_G1063_ & new_G1100_;
  assign new_G1100_ = ~G1045 | ~new_G1070_;
  assign new_G1101_ = new_G1078_ & new_G1098_;
  assign new_G1102_ = ~new_G1078_ & ~new_G1098_;
  assign new_G1103_ = new_G1107_ | new_G1108_;
  assign new_G1104_ = ~G1049 & new_G1063_;
  assign new_G1105_ = new_G1109_ | new_G1110_;
  assign new_G1106_ = G1049 & new_G1063_;
  assign new_G1107_ = ~G1049 & ~new_G1063_;
  assign new_G1108_ = G1049 & ~new_G1063_;
  assign new_G1109_ = G1049 & ~new_G1063_;
  assign new_G1110_ = ~G1049 & new_G1063_;
  assign new_G1117_ = new_G1124_ & new_G1123_;
  assign new_G1118_ = new_G1126_ | new_G1125_;
  assign new_G1119_ = new_G1128_ | new_G1127_;
  assign new_G1120_ = new_G1130_ & new_G1129_;
  assign new_G1121_ = new_G1130_ & new_G1131_;
  assign new_G1122_ = new_G1123_ | new_G1132_;
  assign new_G1123_ = G1112 | new_G1135_;
  assign new_G1124_ = new_G1134_ | new_G1133_;
  assign new_G1125_ = new_G1139_ & new_G1138_;
  assign new_G1126_ = new_G1137_ & new_G1136_;
  assign new_G1127_ = new_G1142_ | new_G1141_;
  assign new_G1128_ = new_G1137_ & new_G1140_;
  assign new_G1129_ = G1112 | new_G1145_;
  assign new_G1130_ = new_G1144_ | new_G1143_;
  assign new_G1131_ = new_G1147_ | new_G1146_;
  assign new_G1132_ = ~new_G1123_ & new_G1149_;
  assign new_G1133_ = ~new_G1125_ & new_G1137_;
  assign new_G1134_ = new_G1125_ & ~new_G1137_;
  assign new_G1135_ = G1111 & ~G1112;
  assign new_G1136_ = ~new_G1158_ | ~new_G1159_;
  assign new_G1137_ = new_G1151_ | new_G1153_;
  assign new_G1138_ = new_G1161_ | new_G1160_;
  assign new_G1139_ = new_G1155_ | new_G1154_;
  assign new_G1140_ = ~new_G1163_ | ~new_G1162_;
  assign new_G1141_ = ~new_G1164_ & new_G1165_;
  assign new_G1142_ = new_G1164_ & ~new_G1165_;
  assign new_G1143_ = ~G1111 & G1112;
  assign new_G1144_ = G1111 & ~G1112;
  assign new_G1145_ = ~new_G1127_ | new_G1137_;
  assign new_G1146_ = new_G1127_ & new_G1137_;
  assign new_G1147_ = ~new_G1127_ & ~new_G1137_;
  assign new_G1148_ = new_G1169_ | new_G1168_;
  assign new_G1149_ = G1115 | new_G1148_;
  assign new_G1150_ = new_G1173_ | new_G1172_;
  assign new_G1151_ = ~G1115 & new_G1150_;
  assign new_G1152_ = new_G1171_ | new_G1170_;
  assign new_G1153_ = G1115 & new_G1152_;
  assign new_G1154_ = G1113 & ~new_G1123_;
  assign new_G1155_ = ~G1113 & new_G1123_;
  assign new_G1156_ = ~G1112 | ~new_G1137_;
  assign new_G1157_ = new_G1123_ & new_G1156_;
  assign new_G1158_ = ~new_G1123_ & ~new_G1157_;
  assign new_G1159_ = new_G1123_ | new_G1156_;
  assign new_G1160_ = ~G1113 & G1114;
  assign new_G1161_ = G1113 & ~G1114;
  assign new_G1162_ = new_G1130_ | new_G1167_;
  assign new_G1163_ = ~new_G1130_ & ~new_G1166_;
  assign new_G1164_ = G1113 | new_G1130_;
  assign new_G1165_ = G1113 | G1114;
  assign new_G1166_ = new_G1130_ & new_G1167_;
  assign new_G1167_ = ~G1112 | ~new_G1137_;
  assign new_G1168_ = new_G1145_ & new_G1165_;
  assign new_G1169_ = ~new_G1145_ & ~new_G1165_;
  assign new_G1170_ = new_G1174_ | new_G1175_;
  assign new_G1171_ = ~G1116 & new_G1130_;
  assign new_G1172_ = new_G1176_ | new_G1177_;
  assign new_G1173_ = G1116 & new_G1130_;
  assign new_G1174_ = ~G1116 & ~new_G1130_;
  assign new_G1175_ = G1116 & ~new_G1130_;
  assign new_G1176_ = G1116 & ~new_G1130_;
  assign new_G1177_ = ~G1116 & new_G1130_;
  assign new_G1184_ = new_G1191_ & new_G1190_;
  assign new_G1185_ = new_G1193_ | new_G1192_;
  assign new_G1186_ = new_G1195_ | new_G1194_;
  assign new_G1187_ = new_G1197_ & new_G1196_;
  assign new_G1188_ = new_G1197_ & new_G1198_;
  assign new_G1189_ = new_G1190_ | new_G1199_;
  assign new_G1190_ = G1179 | new_G1202_;
  assign new_G1191_ = new_G1201_ | new_G1200_;
  assign new_G1192_ = new_G1206_ & new_G1205_;
  assign new_G1193_ = new_G1204_ & new_G1203_;
  assign new_G1194_ = new_G1209_ | new_G1208_;
  assign new_G1195_ = new_G1204_ & new_G1207_;
  assign new_G1196_ = G1179 | new_G1212_;
  assign new_G1197_ = new_G1211_ | new_G1210_;
  assign new_G1198_ = new_G1214_ | new_G1213_;
  assign new_G1199_ = ~new_G1190_ & new_G1216_;
  assign new_G1200_ = ~new_G1192_ & new_G1204_;
  assign new_G1201_ = new_G1192_ & ~new_G1204_;
  assign new_G1202_ = G1178 & ~G1179;
  assign new_G1203_ = ~new_G1225_ | ~new_G1226_;
  assign new_G1204_ = new_G1218_ | new_G1220_;
  assign new_G1205_ = new_G1228_ | new_G1227_;
  assign new_G1206_ = new_G1222_ | new_G1221_;
  assign new_G1207_ = ~new_G1230_ | ~new_G1229_;
  assign new_G1208_ = ~new_G1231_ & new_G1232_;
  assign new_G1209_ = new_G1231_ & ~new_G1232_;
  assign new_G1210_ = ~G1178 & G1179;
  assign new_G1211_ = G1178 & ~G1179;
  assign new_G1212_ = ~new_G1194_ | new_G1204_;
  assign new_G1213_ = new_G1194_ & new_G1204_;
  assign new_G1214_ = ~new_G1194_ & ~new_G1204_;
  assign new_G1215_ = new_G1236_ | new_G1235_;
  assign new_G1216_ = G1182 | new_G1215_;
  assign new_G1217_ = new_G1240_ | new_G1239_;
  assign new_G1218_ = ~G1182 & new_G1217_;
  assign new_G1219_ = new_G1238_ | new_G1237_;
  assign new_G1220_ = G1182 & new_G1219_;
  assign new_G1221_ = G1180 & ~new_G1190_;
  assign new_G1222_ = ~G1180 & new_G1190_;
  assign new_G1223_ = ~G1179 | ~new_G1204_;
  assign new_G1224_ = new_G1190_ & new_G1223_;
  assign new_G1225_ = ~new_G1190_ & ~new_G1224_;
  assign new_G1226_ = new_G1190_ | new_G1223_;
  assign new_G1227_ = ~G1180 & G1181;
  assign new_G1228_ = G1180 & ~G1181;
  assign new_G1229_ = new_G1197_ | new_G1234_;
  assign new_G1230_ = ~new_G1197_ & ~new_G1233_;
  assign new_G1231_ = G1180 | new_G1197_;
  assign new_G1232_ = G1180 | G1181;
  assign new_G1233_ = new_G1197_ & new_G1234_;
  assign new_G1234_ = ~G1179 | ~new_G1204_;
  assign new_G1235_ = new_G1212_ & new_G1232_;
  assign new_G1236_ = ~new_G1212_ & ~new_G1232_;
  assign new_G1237_ = new_G1241_ | new_G1242_;
  assign new_G1238_ = ~G1183 & new_G1197_;
  assign new_G1239_ = new_G1243_ | new_G1244_;
  assign new_G1240_ = G1183 & new_G1197_;
  assign new_G1241_ = ~G1183 & ~new_G1197_;
  assign new_G1242_ = G1183 & ~new_G1197_;
  assign new_G1243_ = G1183 & ~new_G1197_;
  assign new_G1244_ = ~G1183 & new_G1197_;
  assign new_G1251_ = new_G1258_ & new_G1257_;
  assign new_G1252_ = new_G1260_ | new_G1259_;
  assign new_G1253_ = new_G1262_ | new_G1261_;
  assign new_G1254_ = new_G1264_ & new_G1263_;
  assign new_G1255_ = new_G1264_ & new_G1265_;
  assign new_G1256_ = new_G1257_ | new_G1266_;
  assign new_G1257_ = G1246 | new_G1269_;
  assign new_G1258_ = new_G1268_ | new_G1267_;
  assign new_G1259_ = new_G1273_ & new_G1272_;
  assign new_G1260_ = new_G1271_ & new_G1270_;
  assign new_G1261_ = new_G1276_ | new_G1275_;
  assign new_G1262_ = new_G1271_ & new_G1274_;
  assign new_G1263_ = G1246 | new_G1279_;
  assign new_G1264_ = new_G1278_ | new_G1277_;
  assign new_G1265_ = new_G1281_ | new_G1280_;
  assign new_G1266_ = ~new_G1257_ & new_G1283_;
  assign new_G1267_ = ~new_G1259_ & new_G1271_;
  assign new_G1268_ = new_G1259_ & ~new_G1271_;
  assign new_G1269_ = G1245 & ~G1246;
  assign new_G1270_ = ~new_G1292_ | ~new_G1293_;
  assign new_G1271_ = new_G1285_ | new_G1287_;
  assign new_G1272_ = new_G1295_ | new_G1294_;
  assign new_G1273_ = new_G1289_ | new_G1288_;
  assign new_G1274_ = ~new_G1297_ | ~new_G1296_;
  assign new_G1275_ = ~new_G1298_ & new_G1299_;
  assign new_G1276_ = new_G1298_ & ~new_G1299_;
  assign new_G1277_ = ~G1245 & G1246;
  assign new_G1278_ = G1245 & ~G1246;
  assign new_G1279_ = ~new_G1261_ | new_G1271_;
  assign new_G1280_ = new_G1261_ & new_G1271_;
  assign new_G1281_ = ~new_G1261_ & ~new_G1271_;
  assign new_G1282_ = new_G1303_ | new_G1302_;
  assign new_G1283_ = G1249 | new_G1282_;
  assign new_G1284_ = new_G1307_ | new_G1306_;
  assign new_G1285_ = ~G1249 & new_G1284_;
  assign new_G1286_ = new_G1305_ | new_G1304_;
  assign new_G1287_ = G1249 & new_G1286_;
  assign new_G1288_ = G1247 & ~new_G1257_;
  assign new_G1289_ = ~G1247 & new_G1257_;
  assign new_G1290_ = ~G1246 | ~new_G1271_;
  assign new_G1291_ = new_G1257_ & new_G1290_;
  assign new_G1292_ = ~new_G1257_ & ~new_G1291_;
  assign new_G1293_ = new_G1257_ | new_G1290_;
  assign new_G1294_ = ~G1247 & G1248;
  assign new_G1295_ = G1247 & ~G1248;
  assign new_G1296_ = new_G1264_ | new_G1301_;
  assign new_G1297_ = ~new_G1264_ & ~new_G1300_;
  assign new_G1298_ = G1247 | new_G1264_;
  assign new_G1299_ = G1247 | G1248;
  assign new_G1300_ = new_G1264_ & new_G1301_;
  assign new_G1301_ = ~G1246 | ~new_G1271_;
  assign new_G1302_ = new_G1279_ & new_G1299_;
  assign new_G1303_ = ~new_G1279_ & ~new_G1299_;
  assign new_G1304_ = new_G1308_ | new_G1309_;
  assign new_G1305_ = ~G1250 & new_G1264_;
  assign new_G1306_ = new_G1310_ | new_G1311_;
  assign new_G1307_ = G1250 & new_G1264_;
  assign new_G1308_ = ~G1250 & ~new_G1264_;
  assign new_G1309_ = G1250 & ~new_G1264_;
  assign new_G1310_ = G1250 & ~new_G1264_;
  assign new_G1311_ = ~G1250 & new_G1264_;
  assign new_G1318_ = new_G1325_ & new_G1324_;
  assign new_G1319_ = new_G1327_ | new_G1326_;
  assign new_G1320_ = new_G1329_ | new_G1328_;
  assign new_G1321_ = new_G1331_ & new_G1330_;
  assign new_G1322_ = new_G1331_ & new_G1332_;
  assign new_G1323_ = new_G1324_ | new_G1333_;
  assign new_G1324_ = G1313 | new_G1336_;
  assign new_G1325_ = new_G1335_ | new_G1334_;
  assign new_G1326_ = new_G1340_ & new_G1339_;
  assign new_G1327_ = new_G1338_ & new_G1337_;
  assign new_G1328_ = new_G1343_ | new_G1342_;
  assign new_G1329_ = new_G1338_ & new_G1341_;
  assign new_G1330_ = G1313 | new_G1346_;
  assign new_G1331_ = new_G1345_ | new_G1344_;
  assign new_G1332_ = new_G1348_ | new_G1347_;
  assign new_G1333_ = ~new_G1324_ & new_G1350_;
  assign new_G1334_ = ~new_G1326_ & new_G1338_;
  assign new_G1335_ = new_G1326_ & ~new_G1338_;
  assign new_G1336_ = G1312 & ~G1313;
  assign new_G1337_ = ~new_G1359_ | ~new_G1360_;
  assign new_G1338_ = new_G1352_ | new_G1354_;
  assign new_G1339_ = new_G1362_ | new_G1361_;
  assign new_G1340_ = new_G1356_ | new_G1355_;
  assign new_G1341_ = ~new_G1364_ | ~new_G1363_;
  assign new_G1342_ = ~new_G1365_ & new_G1366_;
  assign new_G1343_ = new_G1365_ & ~new_G1366_;
  assign new_G1344_ = ~G1312 & G1313;
  assign new_G1345_ = G1312 & ~G1313;
  assign new_G1346_ = ~new_G1328_ | new_G1338_;
  assign new_G1347_ = new_G1328_ & new_G1338_;
  assign new_G1348_ = ~new_G1328_ & ~new_G1338_;
  assign new_G1349_ = new_G1370_ | new_G1369_;
  assign new_G1350_ = G1316 | new_G1349_;
  assign new_G1351_ = new_G1374_ | new_G1373_;
  assign new_G1352_ = ~G1316 & new_G1351_;
  assign new_G1353_ = new_G1372_ | new_G1371_;
  assign new_G1354_ = G1316 & new_G1353_;
  assign new_G1355_ = G1314 & ~new_G1324_;
  assign new_G1356_ = ~G1314 & new_G1324_;
  assign new_G1357_ = ~G1313 | ~new_G1338_;
  assign new_G1358_ = new_G1324_ & new_G1357_;
  assign new_G1359_ = ~new_G1324_ & ~new_G1358_;
  assign new_G1360_ = new_G1324_ | new_G1357_;
  assign new_G1361_ = ~G1314 & G1315;
  assign new_G1362_ = G1314 & ~G1315;
  assign new_G1363_ = new_G1331_ | new_G1368_;
  assign new_G1364_ = ~new_G1331_ & ~new_G1367_;
  assign new_G1365_ = G1314 | new_G1331_;
  assign new_G1366_ = G1314 | G1315;
  assign new_G1367_ = new_G1331_ & new_G1368_;
  assign new_G1368_ = ~G1313 | ~new_G1338_;
  assign new_G1369_ = new_G1346_ & new_G1366_;
  assign new_G1370_ = ~new_G1346_ & ~new_G1366_;
  assign new_G1371_ = new_G1375_ | new_G1376_;
  assign new_G1372_ = ~G1317 & new_G1331_;
  assign new_G1373_ = new_G1377_ | new_G1378_;
  assign new_G1374_ = G1317 & new_G1331_;
  assign new_G1375_ = ~G1317 & ~new_G1331_;
  assign new_G1376_ = G1317 & ~new_G1331_;
  assign new_G1377_ = G1317 & ~new_G1331_;
  assign new_G1378_ = ~G1317 & new_G1331_;
  assign new_G1385_ = new_G1392_ & new_G1391_;
  assign new_G1386_ = new_G1394_ | new_G1393_;
  assign new_G1387_ = new_G1396_ | new_G1395_;
  assign new_G1388_ = new_G1398_ & new_G1397_;
  assign new_G1389_ = new_G1398_ & new_G1399_;
  assign new_G1390_ = new_G1391_ | new_G1400_;
  assign new_G1391_ = G1380 | new_G1403_;
  assign new_G1392_ = new_G1402_ | new_G1401_;
  assign new_G1393_ = new_G1407_ & new_G1406_;
  assign new_G1394_ = new_G1405_ & new_G1404_;
  assign new_G1395_ = new_G1410_ | new_G1409_;
  assign new_G1396_ = new_G1405_ & new_G1408_;
  assign new_G1397_ = G1380 | new_G1413_;
  assign new_G1398_ = new_G1412_ | new_G1411_;
  assign new_G1399_ = new_G1415_ | new_G1414_;
  assign new_G1400_ = ~new_G1391_ & new_G1417_;
  assign new_G1401_ = ~new_G1393_ & new_G1405_;
  assign new_G1402_ = new_G1393_ & ~new_G1405_;
  assign new_G1403_ = G1379 & ~G1380;
  assign new_G1404_ = ~new_G1426_ | ~new_G1427_;
  assign new_G1405_ = new_G1419_ | new_G1421_;
  assign new_G1406_ = new_G1429_ | new_G1428_;
  assign new_G1407_ = new_G1423_ | new_G1422_;
  assign new_G1408_ = ~new_G1431_ | ~new_G1430_;
  assign new_G1409_ = ~new_G1432_ & new_G1433_;
  assign new_G1410_ = new_G1432_ & ~new_G1433_;
  assign new_G1411_ = ~G1379 & G1380;
  assign new_G1412_ = G1379 & ~G1380;
  assign new_G1413_ = ~new_G1395_ | new_G1405_;
  assign new_G1414_ = new_G1395_ & new_G1405_;
  assign new_G1415_ = ~new_G1395_ & ~new_G1405_;
  assign new_G1416_ = new_G1437_ | new_G1436_;
  assign new_G1417_ = G1383 | new_G1416_;
  assign new_G1418_ = new_G1441_ | new_G1440_;
  assign new_G1419_ = ~G1383 & new_G1418_;
  assign new_G1420_ = new_G1439_ | new_G1438_;
  assign new_G1421_ = G1383 & new_G1420_;
  assign new_G1422_ = G1381 & ~new_G1391_;
  assign new_G1423_ = ~G1381 & new_G1391_;
  assign new_G1424_ = ~G1380 | ~new_G1405_;
  assign new_G1425_ = new_G1391_ & new_G1424_;
  assign new_G1426_ = ~new_G1391_ & ~new_G1425_;
  assign new_G1427_ = new_G1391_ | new_G1424_;
  assign new_G1428_ = ~G1381 & G1382;
  assign new_G1429_ = G1381 & ~G1382;
  assign new_G1430_ = new_G1398_ | new_G1435_;
  assign new_G1431_ = ~new_G1398_ & ~new_G1434_;
  assign new_G1432_ = G1381 | new_G1398_;
  assign new_G1433_ = G1381 | G1382;
  assign new_G1434_ = new_G1398_ & new_G1435_;
  assign new_G1435_ = ~G1380 | ~new_G1405_;
  assign new_G1436_ = new_G1413_ & new_G1433_;
  assign new_G1437_ = ~new_G1413_ & ~new_G1433_;
  assign new_G1438_ = new_G1442_ | new_G1443_;
  assign new_G1439_ = ~G1384 & new_G1398_;
  assign new_G1440_ = new_G1444_ | new_G1445_;
  assign new_G1441_ = G1384 & new_G1398_;
  assign new_G1442_ = ~G1384 & ~new_G1398_;
  assign new_G1443_ = G1384 & ~new_G1398_;
  assign new_G1444_ = G1384 & ~new_G1398_;
  assign new_G1445_ = ~G1384 & new_G1398_;
  assign new_G1452_ = new_G1459_ & new_G1458_;
  assign new_G1453_ = new_G1461_ | new_G1460_;
  assign new_G1454_ = new_G1463_ | new_G1462_;
  assign new_G1455_ = new_G1465_ & new_G1464_;
  assign new_G1456_ = new_G1465_ & new_G1466_;
  assign new_G1457_ = new_G1458_ | new_G1467_;
  assign new_G1458_ = G1447 | new_G1470_;
  assign new_G1459_ = new_G1469_ | new_G1468_;
  assign new_G1460_ = new_G1474_ & new_G1473_;
  assign new_G1461_ = new_G1472_ & new_G1471_;
  assign new_G1462_ = new_G1477_ | new_G1476_;
  assign new_G1463_ = new_G1472_ & new_G1475_;
  assign new_G1464_ = G1447 | new_G1480_;
  assign new_G1465_ = new_G1479_ | new_G1478_;
  assign new_G1466_ = new_G1482_ | new_G1481_;
  assign new_G1467_ = ~new_G1458_ & new_G1484_;
  assign new_G1468_ = ~new_G1460_ & new_G1472_;
  assign new_G1469_ = new_G1460_ & ~new_G1472_;
  assign new_G1470_ = G1446 & ~G1447;
  assign new_G1471_ = ~new_G1493_ | ~new_G1494_;
  assign new_G1472_ = new_G1486_ | new_G1488_;
  assign new_G1473_ = new_G1496_ | new_G1495_;
  assign new_G1474_ = new_G1490_ | new_G1489_;
  assign new_G1475_ = ~new_G1498_ | ~new_G1497_;
  assign new_G1476_ = ~new_G1499_ & new_G1500_;
  assign new_G1477_ = new_G1499_ & ~new_G1500_;
  assign new_G1478_ = ~G1446 & G1447;
  assign new_G1479_ = G1446 & ~G1447;
  assign new_G1480_ = ~new_G1462_ | new_G1472_;
  assign new_G1481_ = new_G1462_ & new_G1472_;
  assign new_G1482_ = ~new_G1462_ & ~new_G1472_;
  assign new_G1483_ = new_G1504_ | new_G1503_;
  assign new_G1484_ = G1450 | new_G1483_;
  assign new_G1485_ = new_G1508_ | new_G1507_;
  assign new_G1486_ = ~G1450 & new_G1485_;
  assign new_G1487_ = new_G1506_ | new_G1505_;
  assign new_G1488_ = G1450 & new_G1487_;
  assign new_G1489_ = G1448 & ~new_G1458_;
  assign new_G1490_ = ~G1448 & new_G1458_;
  assign new_G1491_ = ~G1447 | ~new_G1472_;
  assign new_G1492_ = new_G1458_ & new_G1491_;
  assign new_G1493_ = ~new_G1458_ & ~new_G1492_;
  assign new_G1494_ = new_G1458_ | new_G1491_;
  assign new_G1495_ = ~G1448 & G1449;
  assign new_G1496_ = G1448 & ~G1449;
  assign new_G1497_ = new_G1465_ | new_G1502_;
  assign new_G1498_ = ~new_G1465_ & ~new_G1501_;
  assign new_G1499_ = G1448 | new_G1465_;
  assign new_G1500_ = G1448 | G1449;
  assign new_G1501_ = new_G1465_ & new_G1502_;
  assign new_G1502_ = ~G1447 | ~new_G1472_;
  assign new_G1503_ = new_G1480_ & new_G1500_;
  assign new_G1504_ = ~new_G1480_ & ~new_G1500_;
  assign new_G1505_ = new_G1509_ | new_G1510_;
  assign new_G1506_ = ~G1451 & new_G1465_;
  assign new_G1507_ = new_G1511_ | new_G1512_;
  assign new_G1508_ = G1451 & new_G1465_;
  assign new_G1509_ = ~G1451 & ~new_G1465_;
  assign new_G1510_ = G1451 & ~new_G1465_;
  assign new_G1511_ = G1451 & ~new_G1465_;
  assign new_G1512_ = ~G1451 & new_G1465_;
  assign new_G1519_ = new_G1526_ & new_G1525_;
  assign new_G1520_ = new_G1528_ | new_G1527_;
  assign new_G1521_ = new_G1530_ | new_G1529_;
  assign new_G1522_ = new_G1532_ & new_G1531_;
  assign new_G1523_ = new_G1532_ & new_G1533_;
  assign new_G1524_ = new_G1525_ | new_G1534_;
  assign new_G1525_ = G1514 | new_G1537_;
  assign new_G1526_ = new_G1536_ | new_G1535_;
  assign new_G1527_ = new_G1541_ & new_G1540_;
  assign new_G1528_ = new_G1539_ & new_G1538_;
  assign new_G1529_ = new_G1544_ | new_G1543_;
  assign new_G1530_ = new_G1539_ & new_G1542_;
  assign new_G1531_ = G1514 | new_G1547_;
  assign new_G1532_ = new_G1546_ | new_G1545_;
  assign new_G1533_ = new_G1549_ | new_G1548_;
  assign new_G1534_ = ~new_G1525_ & new_G1551_;
  assign new_G1535_ = ~new_G1527_ & new_G1539_;
  assign new_G1536_ = new_G1527_ & ~new_G1539_;
  assign new_G1537_ = G1513 & ~G1514;
  assign new_G1538_ = ~new_G1560_ | ~new_G1561_;
  assign new_G1539_ = new_G1553_ | new_G1555_;
  assign new_G1540_ = new_G1563_ | new_G1562_;
  assign new_G1541_ = new_G1557_ | new_G1556_;
  assign new_G1542_ = ~new_G1565_ | ~new_G1564_;
  assign new_G1543_ = ~new_G1566_ & new_G1567_;
  assign new_G1544_ = new_G1566_ & ~new_G1567_;
  assign new_G1545_ = ~G1513 & G1514;
  assign new_G1546_ = G1513 & ~G1514;
  assign new_G1547_ = ~new_G1529_ | new_G1539_;
  assign new_G1548_ = new_G1529_ & new_G1539_;
  assign new_G1549_ = ~new_G1529_ & ~new_G1539_;
  assign new_G1550_ = new_G1571_ | new_G1570_;
  assign new_G1551_ = G1517 | new_G1550_;
  assign new_G1552_ = new_G1575_ | new_G1574_;
  assign new_G1553_ = ~G1517 & new_G1552_;
  assign new_G1554_ = new_G1573_ | new_G1572_;
  assign new_G1555_ = G1517 & new_G1554_;
  assign new_G1556_ = G1515 & ~new_G1525_;
  assign new_G1557_ = ~G1515 & new_G1525_;
  assign new_G1558_ = ~G1514 | ~new_G1539_;
  assign new_G1559_ = new_G1525_ & new_G1558_;
  assign new_G1560_ = ~new_G1525_ & ~new_G1559_;
  assign new_G1561_ = new_G1525_ | new_G1558_;
  assign new_G1562_ = ~G1515 & G1516;
  assign new_G1563_ = G1515 & ~G1516;
  assign new_G1564_ = new_G1532_ | new_G1569_;
  assign new_G1565_ = ~new_G1532_ & ~new_G1568_;
  assign new_G1566_ = G1515 | new_G1532_;
  assign new_G1567_ = G1515 | G1516;
  assign new_G1568_ = new_G1532_ & new_G1569_;
  assign new_G1569_ = ~G1514 | ~new_G1539_;
  assign new_G1570_ = new_G1547_ & new_G1567_;
  assign new_G1571_ = ~new_G1547_ & ~new_G1567_;
  assign new_G1572_ = new_G1576_ | new_G1577_;
  assign new_G1573_ = ~G1518 & new_G1532_;
  assign new_G1574_ = new_G1578_ | new_G1579_;
  assign new_G1575_ = G1518 & new_G1532_;
  assign new_G1576_ = ~G1518 & ~new_G1532_;
  assign new_G1577_ = G1518 & ~new_G1532_;
  assign new_G1578_ = G1518 & ~new_G1532_;
  assign new_G1579_ = ~G1518 & new_G1532_;
  assign new_G1586_ = new_G1593_ & new_G1592_;
  assign new_G1587_ = new_G1595_ | new_G1594_;
  assign new_G1588_ = new_G1597_ | new_G1596_;
  assign new_G1589_ = new_G1599_ & new_G1598_;
  assign new_G1590_ = new_G1599_ & new_G1600_;
  assign new_G1591_ = new_G1592_ | new_G1601_;
  assign new_G1592_ = G1581 | new_G1604_;
  assign new_G1593_ = new_G1603_ | new_G1602_;
  assign new_G1594_ = new_G1608_ & new_G1607_;
  assign new_G1595_ = new_G1606_ & new_G1605_;
  assign new_G1596_ = new_G1611_ | new_G1610_;
  assign new_G1597_ = new_G1606_ & new_G1609_;
  assign new_G1598_ = G1581 | new_G1614_;
  assign new_G1599_ = new_G1613_ | new_G1612_;
  assign new_G1600_ = new_G1616_ | new_G1615_;
  assign new_G1601_ = ~new_G1592_ & new_G1618_;
  assign new_G1602_ = ~new_G1594_ & new_G1606_;
  assign new_G1603_ = new_G1594_ & ~new_G1606_;
  assign new_G1604_ = G1580 & ~G1581;
  assign new_G1605_ = ~new_G1627_ | ~new_G1628_;
  assign new_G1606_ = new_G1620_ | new_G1622_;
  assign new_G1607_ = new_G1630_ | new_G1629_;
  assign new_G1608_ = new_G1624_ | new_G1623_;
  assign new_G1609_ = ~new_G1632_ | ~new_G1631_;
  assign new_G1610_ = ~new_G1633_ & new_G1634_;
  assign new_G1611_ = new_G1633_ & ~new_G1634_;
  assign new_G1612_ = ~G1580 & G1581;
  assign new_G1613_ = G1580 & ~G1581;
  assign new_G1614_ = ~new_G1596_ | new_G1606_;
  assign new_G1615_ = new_G1596_ & new_G1606_;
  assign new_G1616_ = ~new_G1596_ & ~new_G1606_;
  assign new_G1617_ = new_G1638_ | new_G1637_;
  assign new_G1618_ = G1584 | new_G1617_;
  assign new_G1619_ = new_G1642_ | new_G1641_;
  assign new_G1620_ = ~G1584 & new_G1619_;
  assign new_G1621_ = new_G1640_ | new_G1639_;
  assign new_G1622_ = G1584 & new_G1621_;
  assign new_G1623_ = G1582 & ~new_G1592_;
  assign new_G1624_ = ~G1582 & new_G1592_;
  assign new_G1625_ = ~G1581 | ~new_G1606_;
  assign new_G1626_ = new_G1592_ & new_G1625_;
  assign new_G1627_ = ~new_G1592_ & ~new_G1626_;
  assign new_G1628_ = new_G1592_ | new_G1625_;
  assign new_G1629_ = ~G1582 & G1583;
  assign new_G1630_ = G1582 & ~G1583;
  assign new_G1631_ = new_G1599_ | new_G1636_;
  assign new_G1632_ = ~new_G1599_ & ~new_G1635_;
  assign new_G1633_ = G1582 | new_G1599_;
  assign new_G1634_ = G1582 | G1583;
  assign new_G1635_ = new_G1599_ & new_G1636_;
  assign new_G1636_ = ~G1581 | ~new_G1606_;
  assign new_G1637_ = new_G1614_ & new_G1634_;
  assign new_G1638_ = ~new_G1614_ & ~new_G1634_;
  assign new_G1639_ = new_G1643_ | new_G1644_;
  assign new_G1640_ = ~G1585 & new_G1599_;
  assign new_G1641_ = new_G1645_ | new_G1646_;
  assign new_G1642_ = G1585 & new_G1599_;
  assign new_G1643_ = ~G1585 & ~new_G1599_;
  assign new_G1644_ = G1585 & ~new_G1599_;
  assign new_G1645_ = G1585 & ~new_G1599_;
  assign new_G1646_ = ~G1585 & new_G1599_;
  assign new_G1653_ = new_G1660_ & new_G1659_;
  assign new_G1654_ = new_G1662_ | new_G1661_;
  assign new_G1655_ = new_G1664_ | new_G1663_;
  assign new_G1656_ = new_G1666_ & new_G1665_;
  assign new_G1657_ = new_G1666_ & new_G1667_;
  assign new_G1658_ = new_G1659_ | new_G1668_;
  assign new_G1659_ = G1648 | new_G1671_;
  assign new_G1660_ = new_G1670_ | new_G1669_;
  assign new_G1661_ = new_G1675_ & new_G1674_;
  assign new_G1662_ = new_G1673_ & new_G1672_;
  assign new_G1663_ = new_G1678_ | new_G1677_;
  assign new_G1664_ = new_G1673_ & new_G1676_;
  assign new_G1665_ = G1648 | new_G1681_;
  assign new_G1666_ = new_G1680_ | new_G1679_;
  assign new_G1667_ = new_G1683_ | new_G1682_;
  assign new_G1668_ = ~new_G1659_ & new_G1685_;
  assign new_G1669_ = ~new_G1661_ & new_G1673_;
  assign new_G1670_ = new_G1661_ & ~new_G1673_;
  assign new_G1671_ = G1647 & ~G1648;
  assign new_G1672_ = ~new_G1694_ | ~new_G1695_;
  assign new_G1673_ = new_G1687_ | new_G1689_;
  assign new_G1674_ = new_G1697_ | new_G1696_;
  assign new_G1675_ = new_G1691_ | new_G1690_;
  assign new_G1676_ = ~new_G1699_ | ~new_G1698_;
  assign new_G1677_ = ~new_G1700_ & new_G1701_;
  assign new_G1678_ = new_G1700_ & ~new_G1701_;
  assign new_G1679_ = ~G1647 & G1648;
  assign new_G1680_ = G1647 & ~G1648;
  assign new_G1681_ = ~new_G1663_ | new_G1673_;
  assign new_G1682_ = new_G1663_ & new_G1673_;
  assign new_G1683_ = ~new_G1663_ & ~new_G1673_;
  assign new_G1684_ = new_G1705_ | new_G1704_;
  assign new_G1685_ = G1651 | new_G1684_;
  assign new_G1686_ = new_G1709_ | new_G1708_;
  assign new_G1687_ = ~G1651 & new_G1686_;
  assign new_G1688_ = new_G1707_ | new_G1706_;
  assign new_G1689_ = G1651 & new_G1688_;
  assign new_G1690_ = G1649 & ~new_G1659_;
  assign new_G1691_ = ~G1649 & new_G1659_;
  assign new_G1692_ = ~G1648 | ~new_G1673_;
  assign new_G1693_ = new_G1659_ & new_G1692_;
  assign new_G1694_ = ~new_G1659_ & ~new_G1693_;
  assign new_G1695_ = new_G1659_ | new_G1692_;
  assign new_G1696_ = ~G1649 & G1650;
  assign new_G1697_ = G1649 & ~G1650;
  assign new_G1698_ = new_G1666_ | new_G1703_;
  assign new_G1699_ = ~new_G1666_ & ~new_G1702_;
  assign new_G1700_ = G1649 | new_G1666_;
  assign new_G1701_ = G1649 | G1650;
  assign new_G1702_ = new_G1666_ & new_G1703_;
  assign new_G1703_ = ~G1648 | ~new_G1673_;
  assign new_G1704_ = new_G1681_ & new_G1701_;
  assign new_G1705_ = ~new_G1681_ & ~new_G1701_;
  assign new_G1706_ = new_G1710_ | new_G1711_;
  assign new_G1707_ = ~G1652 & new_G1666_;
  assign new_G1708_ = new_G1712_ | new_G1713_;
  assign new_G1709_ = G1652 & new_G1666_;
  assign new_G1710_ = ~G1652 & ~new_G1666_;
  assign new_G1711_ = G1652 & ~new_G1666_;
  assign new_G1712_ = G1652 & ~new_G1666_;
  assign new_G1713_ = ~G1652 & new_G1666_;
  assign new_G1720_ = new_G1727_ & new_G1726_;
  assign new_G1721_ = new_G1729_ | new_G1728_;
  assign new_G1722_ = new_G1731_ | new_G1730_;
  assign new_G1723_ = new_G1733_ & new_G1732_;
  assign new_G1724_ = new_G1733_ & new_G1734_;
  assign new_G1725_ = new_G1726_ | new_G1735_;
  assign new_G1726_ = G1715 | new_G1738_;
  assign new_G1727_ = new_G1737_ | new_G1736_;
  assign new_G1728_ = new_G1742_ & new_G1741_;
  assign new_G1729_ = new_G1740_ & new_G1739_;
  assign new_G1730_ = new_G1745_ | new_G1744_;
  assign new_G1731_ = new_G1740_ & new_G1743_;
  assign new_G1732_ = G1715 | new_G1748_;
  assign new_G1733_ = new_G1747_ | new_G1746_;
  assign new_G1734_ = new_G1750_ | new_G1749_;
  assign new_G1735_ = ~new_G1726_ & new_G1752_;
  assign new_G1736_ = ~new_G1728_ & new_G1740_;
  assign new_G1737_ = new_G1728_ & ~new_G1740_;
  assign new_G1738_ = G1714 & ~G1715;
  assign new_G1739_ = ~new_G1761_ | ~new_G1762_;
  assign new_G1740_ = new_G1754_ | new_G1756_;
  assign new_G1741_ = new_G1764_ | new_G1763_;
  assign new_G1742_ = new_G1758_ | new_G1757_;
  assign new_G1743_ = ~new_G1766_ | ~new_G1765_;
  assign new_G1744_ = ~new_G1767_ & new_G1768_;
  assign new_G1745_ = new_G1767_ & ~new_G1768_;
  assign new_G1746_ = ~G1714 & G1715;
  assign new_G1747_ = G1714 & ~G1715;
  assign new_G1748_ = ~new_G1730_ | new_G1740_;
  assign new_G1749_ = new_G1730_ & new_G1740_;
  assign new_G1750_ = ~new_G1730_ & ~new_G1740_;
  assign new_G1751_ = new_G1772_ | new_G1771_;
  assign new_G1752_ = G1718 | new_G1751_;
  assign new_G1753_ = new_G1776_ | new_G1775_;
  assign new_G1754_ = ~G1718 & new_G1753_;
  assign new_G1755_ = new_G1774_ | new_G1773_;
  assign new_G1756_ = G1718 & new_G1755_;
  assign new_G1757_ = G1716 & ~new_G1726_;
  assign new_G1758_ = ~G1716 & new_G1726_;
  assign new_G1759_ = ~G1715 | ~new_G1740_;
  assign new_G1760_ = new_G1726_ & new_G1759_;
  assign new_G1761_ = ~new_G1726_ & ~new_G1760_;
  assign new_G1762_ = new_G1726_ | new_G1759_;
  assign new_G1763_ = ~G1716 & G1717;
  assign new_G1764_ = G1716 & ~G1717;
  assign new_G1765_ = new_G1733_ | new_G1770_;
  assign new_G1766_ = ~new_G1733_ & ~new_G1769_;
  assign new_G1767_ = G1716 | new_G1733_;
  assign new_G1768_ = G1716 | G1717;
  assign new_G1769_ = new_G1733_ & new_G1770_;
  assign new_G1770_ = ~G1715 | ~new_G1740_;
  assign new_G1771_ = new_G1748_ & new_G1768_;
  assign new_G1772_ = ~new_G1748_ & ~new_G1768_;
  assign new_G1773_ = new_G1777_ | new_G1778_;
  assign new_G1774_ = ~G1719 & new_G1733_;
  assign new_G1775_ = new_G1779_ | new_G1780_;
  assign new_G1776_ = G1719 & new_G1733_;
  assign new_G1777_ = ~G1719 & ~new_G1733_;
  assign new_G1778_ = G1719 & ~new_G1733_;
  assign new_G1779_ = G1719 & ~new_G1733_;
  assign new_G1780_ = ~G1719 & new_G1733_;
  assign new_G1787_ = new_G1794_ & new_G1793_;
  assign new_G1788_ = new_G1796_ | new_G1795_;
  assign new_G1789_ = new_G1798_ | new_G1797_;
  assign new_G1790_ = new_G1800_ & new_G1799_;
  assign new_G1791_ = new_G1800_ & new_G1801_;
  assign new_G1792_ = new_G1793_ | new_G1802_;
  assign new_G1793_ = G1782 | new_G1805_;
  assign new_G1794_ = new_G1804_ | new_G1803_;
  assign new_G1795_ = new_G1809_ & new_G1808_;
  assign new_G1796_ = new_G1807_ & new_G1806_;
  assign new_G1797_ = new_G1812_ | new_G1811_;
  assign new_G1798_ = new_G1807_ & new_G1810_;
  assign new_G1799_ = G1782 | new_G1815_;
  assign new_G1800_ = new_G1814_ | new_G1813_;
  assign new_G1801_ = new_G1817_ | new_G1816_;
  assign new_G1802_ = ~new_G1793_ & new_G1819_;
  assign new_G1803_ = ~new_G1795_ & new_G1807_;
  assign new_G1804_ = new_G1795_ & ~new_G1807_;
  assign new_G1805_ = G1781 & ~G1782;
  assign new_G1806_ = ~new_G1828_ | ~new_G1829_;
  assign new_G1807_ = new_G1821_ | new_G1823_;
  assign new_G1808_ = new_G1831_ | new_G1830_;
  assign new_G1809_ = new_G1825_ | new_G1824_;
  assign new_G1810_ = ~new_G1833_ | ~new_G1832_;
  assign new_G1811_ = ~new_G1834_ & new_G1835_;
  assign new_G1812_ = new_G1834_ & ~new_G1835_;
  assign new_G1813_ = ~G1781 & G1782;
  assign new_G1814_ = G1781 & ~G1782;
  assign new_G1815_ = ~new_G1797_ | new_G1807_;
  assign new_G1816_ = new_G1797_ & new_G1807_;
  assign new_G1817_ = ~new_G1797_ & ~new_G1807_;
  assign new_G1818_ = new_G1839_ | new_G1838_;
  assign new_G1819_ = G1785 | new_G1818_;
  assign new_G1820_ = new_G1843_ | new_G1842_;
  assign new_G1821_ = ~G1785 & new_G1820_;
  assign new_G1822_ = new_G1841_ | new_G1840_;
  assign new_G1823_ = G1785 & new_G1822_;
  assign new_G1824_ = G1783 & ~new_G1793_;
  assign new_G1825_ = ~G1783 & new_G1793_;
  assign new_G1826_ = ~G1782 | ~new_G1807_;
  assign new_G1827_ = new_G1793_ & new_G1826_;
  assign new_G1828_ = ~new_G1793_ & ~new_G1827_;
  assign new_G1829_ = new_G1793_ | new_G1826_;
  assign new_G1830_ = ~G1783 & G1784;
  assign new_G1831_ = G1783 & ~G1784;
  assign new_G1832_ = new_G1800_ | new_G1837_;
  assign new_G1833_ = ~new_G1800_ & ~new_G1836_;
  assign new_G1834_ = G1783 | new_G1800_;
  assign new_G1835_ = G1783 | G1784;
  assign new_G1836_ = new_G1800_ & new_G1837_;
  assign new_G1837_ = ~G1782 | ~new_G1807_;
  assign new_G1838_ = new_G1815_ & new_G1835_;
  assign new_G1839_ = ~new_G1815_ & ~new_G1835_;
  assign new_G1840_ = new_G1844_ | new_G1845_;
  assign new_G1841_ = ~G1786 & new_G1800_;
  assign new_G1842_ = new_G1846_ | new_G1847_;
  assign new_G1843_ = G1786 & new_G1800_;
  assign new_G1844_ = ~G1786 & ~new_G1800_;
  assign new_G1845_ = G1786 & ~new_G1800_;
  assign new_G1846_ = G1786 & ~new_G1800_;
  assign new_G1847_ = ~G1786 & new_G1800_;
  assign new_G1854_ = new_G1861_ & new_G1860_;
  assign new_G1855_ = new_G1863_ | new_G1862_;
  assign new_G1856_ = new_G1865_ | new_G1864_;
  assign new_G1857_ = new_G1867_ & new_G1866_;
  assign new_G1858_ = new_G1867_ & new_G1868_;
  assign new_G1859_ = new_G1860_ | new_G1869_;
  assign new_G1860_ = G1849 | new_G1872_;
  assign new_G1861_ = new_G1871_ | new_G1870_;
  assign new_G1862_ = new_G1876_ & new_G1875_;
  assign new_G1863_ = new_G1874_ & new_G1873_;
  assign new_G1864_ = new_G1879_ | new_G1878_;
  assign new_G1865_ = new_G1874_ & new_G1877_;
  assign new_G1866_ = G1849 | new_G1882_;
  assign new_G1867_ = new_G1881_ | new_G1880_;
  assign new_G1868_ = new_G1884_ | new_G1883_;
  assign new_G1869_ = ~new_G1860_ & new_G1886_;
  assign new_G1870_ = ~new_G1862_ & new_G1874_;
  assign new_G1871_ = new_G1862_ & ~new_G1874_;
  assign new_G1872_ = G1848 & ~G1849;
  assign new_G1873_ = ~new_G1895_ | ~new_G1896_;
  assign new_G1874_ = new_G1888_ | new_G1890_;
  assign new_G1875_ = new_G1898_ | new_G1897_;
  assign new_G1876_ = new_G1892_ | new_G1891_;
  assign new_G1877_ = ~new_G1900_ | ~new_G1899_;
  assign new_G1878_ = ~new_G1901_ & new_G1902_;
  assign new_G1879_ = new_G1901_ & ~new_G1902_;
  assign new_G1880_ = ~G1848 & G1849;
  assign new_G1881_ = G1848 & ~G1849;
  assign new_G1882_ = ~new_G1864_ | new_G1874_;
  assign new_G1883_ = new_G1864_ & new_G1874_;
  assign new_G1884_ = ~new_G1864_ & ~new_G1874_;
  assign new_G1885_ = new_G1906_ | new_G1905_;
  assign new_G1886_ = G1852 | new_G1885_;
  assign new_G1887_ = new_G1910_ | new_G1909_;
  assign new_G1888_ = ~G1852 & new_G1887_;
  assign new_G1889_ = new_G1908_ | new_G1907_;
  assign new_G1890_ = G1852 & new_G1889_;
  assign new_G1891_ = G1850 & ~new_G1860_;
  assign new_G1892_ = ~G1850 & new_G1860_;
  assign new_G1893_ = ~G1849 | ~new_G1874_;
  assign new_G1894_ = new_G1860_ & new_G1893_;
  assign new_G1895_ = ~new_G1860_ & ~new_G1894_;
  assign new_G1896_ = new_G1860_ | new_G1893_;
  assign new_G1897_ = ~G1850 & G1851;
  assign new_G1898_ = G1850 & ~G1851;
  assign new_G1899_ = new_G1867_ | new_G1904_;
  assign new_G1900_ = ~new_G1867_ & ~new_G1903_;
  assign new_G1901_ = G1850 | new_G1867_;
  assign new_G1902_ = G1850 | G1851;
  assign new_G1903_ = new_G1867_ & new_G1904_;
  assign new_G1904_ = ~G1849 | ~new_G1874_;
  assign new_G1905_ = new_G1882_ & new_G1902_;
  assign new_G1906_ = ~new_G1882_ & ~new_G1902_;
  assign new_G1907_ = new_G1911_ | new_G1912_;
  assign new_G1908_ = ~G1853 & new_G1867_;
  assign new_G1909_ = new_G1913_ | new_G1914_;
  assign new_G1910_ = G1853 & new_G1867_;
  assign new_G1911_ = ~G1853 & ~new_G1867_;
  assign new_G1912_ = G1853 & ~new_G1867_;
  assign new_G1913_ = G1853 & ~new_G1867_;
  assign new_G1914_ = ~G1853 & new_G1867_;
  assign new_G1921_ = new_G1928_ & new_G1927_;
  assign new_G1922_ = new_G1930_ | new_G1929_;
  assign new_G1923_ = new_G1932_ | new_G1931_;
  assign new_G1924_ = new_G1934_ & new_G1933_;
  assign new_G1925_ = new_G1934_ & new_G1935_;
  assign new_G1926_ = new_G1927_ | new_G1936_;
  assign new_G1927_ = G1916 | new_G1939_;
  assign new_G1928_ = new_G1938_ | new_G1937_;
  assign new_G1929_ = new_G1943_ & new_G1942_;
  assign new_G1930_ = new_G1941_ & new_G1940_;
  assign new_G1931_ = new_G1946_ | new_G1945_;
  assign new_G1932_ = new_G1941_ & new_G1944_;
  assign new_G1933_ = G1916 | new_G1949_;
  assign new_G1934_ = new_G1948_ | new_G1947_;
  assign new_G1935_ = new_G1951_ | new_G1950_;
  assign new_G1936_ = ~new_G1927_ & new_G1953_;
  assign new_G1937_ = ~new_G1929_ & new_G1941_;
  assign new_G1938_ = new_G1929_ & ~new_G1941_;
  assign new_G1939_ = G1915 & ~G1916;
  assign new_G1940_ = ~new_G1962_ | ~new_G1963_;
  assign new_G1941_ = new_G1955_ | new_G1957_;
  assign new_G1942_ = new_G1965_ | new_G1964_;
  assign new_G1943_ = new_G1959_ | new_G1958_;
  assign new_G1944_ = ~new_G1967_ | ~new_G1966_;
  assign new_G1945_ = ~new_G1968_ & new_G1969_;
  assign new_G1946_ = new_G1968_ & ~new_G1969_;
  assign new_G1947_ = ~G1915 & G1916;
  assign new_G1948_ = G1915 & ~G1916;
  assign new_G1949_ = ~new_G1931_ | new_G1941_;
  assign new_G1950_ = new_G1931_ & new_G1941_;
  assign new_G1951_ = ~new_G1931_ & ~new_G1941_;
  assign new_G1952_ = new_G1973_ | new_G1972_;
  assign new_G1953_ = G1919 | new_G1952_;
  assign new_G1954_ = new_G1977_ | new_G1976_;
  assign new_G1955_ = ~G1919 & new_G1954_;
  assign new_G1956_ = new_G1975_ | new_G1974_;
  assign new_G1957_ = G1919 & new_G1956_;
  assign new_G1958_ = G1917 & ~new_G1927_;
  assign new_G1959_ = ~G1917 & new_G1927_;
  assign new_G1960_ = ~G1916 | ~new_G1941_;
  assign new_G1961_ = new_G1927_ & new_G1960_;
  assign new_G1962_ = ~new_G1927_ & ~new_G1961_;
  assign new_G1963_ = new_G1927_ | new_G1960_;
  assign new_G1964_ = ~G1917 & G1918;
  assign new_G1965_ = G1917 & ~G1918;
  assign new_G1966_ = new_G1934_ | new_G1971_;
  assign new_G1967_ = ~new_G1934_ & ~new_G1970_;
  assign new_G1968_ = G1917 | new_G1934_;
  assign new_G1969_ = G1917 | G1918;
  assign new_G1970_ = new_G1934_ & new_G1971_;
  assign new_G1971_ = ~G1916 | ~new_G1941_;
  assign new_G1972_ = new_G1949_ & new_G1969_;
  assign new_G1973_ = ~new_G1949_ & ~new_G1969_;
  assign new_G1974_ = new_G1978_ | new_G1979_;
  assign new_G1975_ = ~G1920 & new_G1934_;
  assign new_G1976_ = new_G1980_ | new_G1981_;
  assign new_G1977_ = G1920 & new_G1934_;
  assign new_G1978_ = ~G1920 & ~new_G1934_;
  assign new_G1979_ = G1920 & ~new_G1934_;
  assign new_G1980_ = G1920 & ~new_G1934_;
  assign new_G1981_ = ~G1920 & new_G1934_;
  assign new_G1988_ = new_G1995_ & new_G1994_;
  assign new_G1989_ = new_G1997_ | new_G1996_;
  assign new_G1990_ = new_G1999_ | new_G1998_;
  assign new_G1991_ = new_G2001_ & new_G2000_;
  assign new_G1992_ = new_G2001_ & new_G2002_;
  assign new_G1993_ = new_G1994_ | new_G2003_;
  assign new_G1994_ = G1983 | new_G2006_;
  assign new_G1995_ = new_G2005_ | new_G2004_;
  assign new_G1996_ = new_G2010_ & new_G2009_;
  assign new_G1997_ = new_G2008_ & new_G2007_;
  assign new_G1998_ = new_G2013_ | new_G2012_;
  assign new_G1999_ = new_G2008_ & new_G2011_;
  assign new_G2000_ = G1983 | new_G2016_;
  assign new_G2001_ = new_G2015_ | new_G2014_;
  assign new_G2002_ = new_G2018_ | new_G2017_;
  assign new_G2003_ = ~new_G1994_ & new_G2020_;
  assign new_G2004_ = ~new_G1996_ & new_G2008_;
  assign new_G2005_ = new_G1996_ & ~new_G2008_;
  assign new_G2006_ = G1982 & ~G1983;
  assign new_G2007_ = ~new_G2029_ | ~new_G2030_;
  assign new_G2008_ = new_G2022_ | new_G2024_;
  assign new_G2009_ = new_G2032_ | new_G2031_;
  assign new_G2010_ = new_G2026_ | new_G2025_;
  assign new_G2011_ = ~new_G2034_ | ~new_G2033_;
  assign new_G2012_ = ~new_G2035_ & new_G2036_;
  assign new_G2013_ = new_G2035_ & ~new_G2036_;
  assign new_G2014_ = ~G1982 & G1983;
  assign new_G2015_ = G1982 & ~G1983;
  assign new_G2016_ = ~new_G1998_ | new_G2008_;
  assign new_G2017_ = new_G1998_ & new_G2008_;
  assign new_G2018_ = ~new_G1998_ & ~new_G2008_;
  assign new_G2019_ = new_G2040_ | new_G2039_;
  assign new_G2020_ = G1986 | new_G2019_;
  assign new_G2021_ = new_G2044_ | new_G2043_;
  assign new_G2022_ = ~G1986 & new_G2021_;
  assign new_G2023_ = new_G2042_ | new_G2041_;
  assign new_G2024_ = G1986 & new_G2023_;
  assign new_G2025_ = G1984 & ~new_G1994_;
  assign new_G2026_ = ~G1984 & new_G1994_;
  assign new_G2027_ = ~G1983 | ~new_G2008_;
  assign new_G2028_ = new_G1994_ & new_G2027_;
  assign new_G2029_ = ~new_G1994_ & ~new_G2028_;
  assign new_G2030_ = new_G1994_ | new_G2027_;
  assign new_G2031_ = ~G1984 & G1985;
  assign new_G2032_ = G1984 & ~G1985;
  assign new_G2033_ = new_G2001_ | new_G2038_;
  assign new_G2034_ = ~new_G2001_ & ~new_G2037_;
  assign new_G2035_ = G1984 | new_G2001_;
  assign new_G2036_ = G1984 | G1985;
  assign new_G2037_ = new_G2001_ & new_G2038_;
  assign new_G2038_ = ~G1983 | ~new_G2008_;
  assign new_G2039_ = new_G2016_ & new_G2036_;
  assign new_G2040_ = ~new_G2016_ & ~new_G2036_;
  assign new_G2041_ = new_G2045_ | new_G2046_;
  assign new_G2042_ = ~G1987 & new_G2001_;
  assign new_G2043_ = new_G2047_ | new_G2048_;
  assign new_G2044_ = G1987 & new_G2001_;
  assign new_G2045_ = ~G1987 & ~new_G2001_;
  assign new_G2046_ = G1987 & ~new_G2001_;
  assign new_G2047_ = G1987 & ~new_G2001_;
  assign new_G2048_ = ~G1987 & new_G2001_;
  assign new_G2055_ = new_G2062_ & new_G2061_;
  assign new_G2056_ = new_G2064_ | new_G2063_;
  assign new_G2057_ = new_G2066_ | new_G2065_;
  assign new_G2058_ = new_G2068_ & new_G2067_;
  assign new_G2059_ = new_G2068_ & new_G2069_;
  assign new_G2060_ = new_G2061_ | new_G2070_;
  assign new_G2061_ = G2050 | new_G2073_;
  assign new_G2062_ = new_G2072_ | new_G2071_;
  assign new_G2063_ = new_G2077_ & new_G2076_;
  assign new_G2064_ = new_G2075_ & new_G2074_;
  assign new_G2065_ = new_G2080_ | new_G2079_;
  assign new_G2066_ = new_G2075_ & new_G2078_;
  assign new_G2067_ = G2050 | new_G2083_;
  assign new_G2068_ = new_G2082_ | new_G2081_;
  assign new_G2069_ = new_G2085_ | new_G2084_;
  assign new_G2070_ = ~new_G2061_ & new_G2087_;
  assign new_G2071_ = ~new_G2063_ & new_G2075_;
  assign new_G2072_ = new_G2063_ & ~new_G2075_;
  assign new_G2073_ = G2049 & ~G2050;
  assign new_G2074_ = ~new_G2096_ | ~new_G2097_;
  assign new_G2075_ = new_G2089_ | new_G2091_;
  assign new_G2076_ = new_G2099_ | new_G2098_;
  assign new_G2077_ = new_G2093_ | new_G2092_;
  assign new_G2078_ = ~new_G2101_ | ~new_G2100_;
  assign new_G2079_ = ~new_G2102_ & new_G2103_;
  assign new_G2080_ = new_G2102_ & ~new_G2103_;
  assign new_G2081_ = ~G2049 & G2050;
  assign new_G2082_ = G2049 & ~G2050;
  assign new_G2083_ = ~new_G2065_ | new_G2075_;
  assign new_G2084_ = new_G2065_ & new_G2075_;
  assign new_G2085_ = ~new_G2065_ & ~new_G2075_;
  assign new_G2086_ = new_G2107_ | new_G2106_;
  assign new_G2087_ = G2053 | new_G2086_;
  assign new_G2088_ = new_G2111_ | new_G2110_;
  assign new_G2089_ = ~G2053 & new_G2088_;
  assign new_G2090_ = new_G2109_ | new_G2108_;
  assign new_G2091_ = G2053 & new_G2090_;
  assign new_G2092_ = G2051 & ~new_G2061_;
  assign new_G2093_ = ~G2051 & new_G2061_;
  assign new_G2094_ = ~G2050 | ~new_G2075_;
  assign new_G2095_ = new_G2061_ & new_G2094_;
  assign new_G2096_ = ~new_G2061_ & ~new_G2095_;
  assign new_G2097_ = new_G2061_ | new_G2094_;
  assign new_G2098_ = ~G2051 & G2052;
  assign new_G2099_ = G2051 & ~G2052;
  assign new_G2100_ = new_G2068_ | new_G2105_;
  assign new_G2101_ = ~new_G2068_ & ~new_G2104_;
  assign new_G2102_ = G2051 | new_G2068_;
  assign new_G2103_ = G2051 | G2052;
  assign new_G2104_ = new_G2068_ & new_G2105_;
  assign new_G2105_ = ~G2050 | ~new_G2075_;
  assign new_G2106_ = new_G2083_ & new_G2103_;
  assign new_G2107_ = ~new_G2083_ & ~new_G2103_;
  assign new_G2108_ = new_G2112_ | new_G2113_;
  assign new_G2109_ = ~G2054 & new_G2068_;
  assign new_G2110_ = new_G2114_ | new_G2115_;
  assign new_G2111_ = G2054 & new_G2068_;
  assign new_G2112_ = ~G2054 & ~new_G2068_;
  assign new_G2113_ = G2054 & ~new_G2068_;
  assign new_G2114_ = G2054 & ~new_G2068_;
  assign new_G2115_ = ~G2054 & new_G2068_;
  assign new_G2122_ = new_G2129_ & new_G2128_;
  assign new_G2123_ = new_G2131_ | new_G2130_;
  assign new_G2124_ = new_G2133_ | new_G2132_;
  assign new_G2125_ = new_G2135_ & new_G2134_;
  assign new_G2126_ = new_G2135_ & new_G2136_;
  assign new_G2127_ = new_G2128_ | new_G2137_;
  assign new_G2128_ = G2117 | new_G2140_;
  assign new_G2129_ = new_G2139_ | new_G2138_;
  assign new_G2130_ = new_G2144_ & new_G2143_;
  assign new_G2131_ = new_G2142_ & new_G2141_;
  assign new_G2132_ = new_G2147_ | new_G2146_;
  assign new_G2133_ = new_G2142_ & new_G2145_;
  assign new_G2134_ = G2117 | new_G2150_;
  assign new_G2135_ = new_G2149_ | new_G2148_;
  assign new_G2136_ = new_G2152_ | new_G2151_;
  assign new_G2137_ = ~new_G2128_ & new_G2154_;
  assign new_G2138_ = ~new_G2130_ & new_G2142_;
  assign new_G2139_ = new_G2130_ & ~new_G2142_;
  assign new_G2140_ = G2116 & ~G2117;
  assign new_G2141_ = ~new_G2163_ | ~new_G2164_;
  assign new_G2142_ = new_G2156_ | new_G2158_;
  assign new_G2143_ = new_G2166_ | new_G2165_;
  assign new_G2144_ = new_G2160_ | new_G2159_;
  assign new_G2145_ = ~new_G2168_ | ~new_G2167_;
  assign new_G2146_ = ~new_G2169_ & new_G2170_;
  assign new_G2147_ = new_G2169_ & ~new_G2170_;
  assign new_G2148_ = ~G2116 & G2117;
  assign new_G2149_ = G2116 & ~G2117;
  assign new_G2150_ = ~new_G2132_ | new_G2142_;
  assign new_G2151_ = new_G2132_ & new_G2142_;
  assign new_G2152_ = ~new_G2132_ & ~new_G2142_;
  assign new_G2153_ = new_G2174_ | new_G2173_;
  assign new_G2154_ = G2120 | new_G2153_;
  assign new_G2155_ = new_G2178_ | new_G2177_;
  assign new_G2156_ = ~G2120 & new_G2155_;
  assign new_G2157_ = new_G2176_ | new_G2175_;
  assign new_G2158_ = G2120 & new_G2157_;
  assign new_G2159_ = G2118 & ~new_G2128_;
  assign new_G2160_ = ~G2118 & new_G2128_;
  assign new_G2161_ = ~G2117 | ~new_G2142_;
  assign new_G2162_ = new_G2128_ & new_G2161_;
  assign new_G2163_ = ~new_G2128_ & ~new_G2162_;
  assign new_G2164_ = new_G2128_ | new_G2161_;
  assign new_G2165_ = ~G2118 & G2119;
  assign new_G2166_ = G2118 & ~G2119;
  assign new_G2167_ = new_G2135_ | new_G2172_;
  assign new_G2168_ = ~new_G2135_ & ~new_G2171_;
  assign new_G2169_ = G2118 | new_G2135_;
  assign new_G2170_ = G2118 | G2119;
  assign new_G2171_ = new_G2135_ & new_G2172_;
  assign new_G2172_ = ~G2117 | ~new_G2142_;
  assign new_G2173_ = new_G2150_ & new_G2170_;
  assign new_G2174_ = ~new_G2150_ & ~new_G2170_;
  assign new_G2175_ = new_G2179_ | new_G2180_;
  assign new_G2176_ = ~G2121 & new_G2135_;
  assign new_G2177_ = new_G2181_ | new_G2182_;
  assign new_G2178_ = G2121 & new_G2135_;
  assign new_G2179_ = ~G2121 & ~new_G2135_;
  assign new_G2180_ = G2121 & ~new_G2135_;
  assign new_G2181_ = G2121 & ~new_G2135_;
  assign new_G2182_ = ~G2121 & new_G2135_;
  assign new_G2189_ = new_G2196_ & new_G2195_;
  assign new_G2190_ = new_G2198_ | new_G2197_;
  assign new_G2191_ = new_G2200_ | new_G2199_;
  assign new_G2192_ = new_G2202_ & new_G2201_;
  assign new_G2193_ = new_G2202_ & new_G2203_;
  assign new_G2194_ = new_G2195_ | new_G2204_;
  assign new_G2195_ = G2184 | new_G2207_;
  assign new_G2196_ = new_G2206_ | new_G2205_;
  assign new_G2197_ = new_G2211_ & new_G2210_;
  assign new_G2198_ = new_G2209_ & new_G2208_;
  assign new_G2199_ = new_G2214_ | new_G2213_;
  assign new_G2200_ = new_G2209_ & new_G2212_;
  assign new_G2201_ = G2184 | new_G2217_;
  assign new_G2202_ = new_G2216_ | new_G2215_;
  assign new_G2203_ = new_G2219_ | new_G2218_;
  assign new_G2204_ = ~new_G2195_ & new_G2221_;
  assign new_G2205_ = ~new_G2197_ & new_G2209_;
  assign new_G2206_ = new_G2197_ & ~new_G2209_;
  assign new_G2207_ = G2183 & ~G2184;
  assign new_G2208_ = ~new_G2230_ | ~new_G2231_;
  assign new_G2209_ = new_G2223_ | new_G2225_;
  assign new_G2210_ = new_G2233_ | new_G2232_;
  assign new_G2211_ = new_G2227_ | new_G2226_;
  assign new_G2212_ = ~new_G2235_ | ~new_G2234_;
  assign new_G2213_ = ~new_G2236_ & new_G2237_;
  assign new_G2214_ = new_G2236_ & ~new_G2237_;
  assign new_G2215_ = ~G2183 & G2184;
  assign new_G2216_ = G2183 & ~G2184;
  assign new_G2217_ = ~new_G2199_ | new_G2209_;
  assign new_G2218_ = new_G2199_ & new_G2209_;
  assign new_G2219_ = ~new_G2199_ & ~new_G2209_;
  assign new_G2220_ = new_G2241_ | new_G2240_;
  assign new_G2221_ = G2187 | new_G2220_;
  assign new_G2222_ = new_G2245_ | new_G2244_;
  assign new_G2223_ = ~G2187 & new_G2222_;
  assign new_G2224_ = new_G2243_ | new_G2242_;
  assign new_G2225_ = G2187 & new_G2224_;
  assign new_G2226_ = G2185 & ~new_G2195_;
  assign new_G2227_ = ~G2185 & new_G2195_;
  assign new_G2228_ = ~G2184 | ~new_G2209_;
  assign new_G2229_ = new_G2195_ & new_G2228_;
  assign new_G2230_ = ~new_G2195_ & ~new_G2229_;
  assign new_G2231_ = new_G2195_ | new_G2228_;
  assign new_G2232_ = ~G2185 & G2186;
  assign new_G2233_ = G2185 & ~G2186;
  assign new_G2234_ = new_G2202_ | new_G2239_;
  assign new_G2235_ = ~new_G2202_ & ~new_G2238_;
  assign new_G2236_ = G2185 | new_G2202_;
  assign new_G2237_ = G2185 | G2186;
  assign new_G2238_ = new_G2202_ & new_G2239_;
  assign new_G2239_ = ~G2184 | ~new_G2209_;
  assign new_G2240_ = new_G2217_ & new_G2237_;
  assign new_G2241_ = ~new_G2217_ & ~new_G2237_;
  assign new_G2242_ = new_G2246_ | new_G2247_;
  assign new_G2243_ = ~G2188 & new_G2202_;
  assign new_G2244_ = new_G2248_ | new_G2249_;
  assign new_G2245_ = G2188 & new_G2202_;
  assign new_G2246_ = ~G2188 & ~new_G2202_;
  assign new_G2247_ = G2188 & ~new_G2202_;
  assign new_G2248_ = G2188 & ~new_G2202_;
  assign new_G2249_ = ~G2188 & new_G2202_;
  assign new_G2256_ = new_G2263_ & new_G2262_;
  assign new_G2257_ = new_G2265_ | new_G2264_;
  assign new_G2258_ = new_G2267_ | new_G2266_;
  assign new_G2259_ = new_G2269_ & new_G2268_;
  assign new_G2260_ = new_G2269_ & new_G2270_;
  assign new_G2261_ = new_G2262_ | new_G2271_;
  assign new_G2262_ = G2251 | new_G2274_;
  assign new_G2263_ = new_G2273_ | new_G2272_;
  assign new_G2264_ = new_G2278_ & new_G2277_;
  assign new_G2265_ = new_G2276_ & new_G2275_;
  assign new_G2266_ = new_G2281_ | new_G2280_;
  assign new_G2267_ = new_G2276_ & new_G2279_;
  assign new_G2268_ = G2251 | new_G2284_;
  assign new_G2269_ = new_G2283_ | new_G2282_;
  assign new_G2270_ = new_G2286_ | new_G2285_;
  assign new_G2271_ = ~new_G2262_ & new_G2288_;
  assign new_G2272_ = ~new_G2264_ & new_G2276_;
  assign new_G2273_ = new_G2264_ & ~new_G2276_;
  assign new_G2274_ = G2250 & ~G2251;
  assign new_G2275_ = ~new_G2297_ | ~new_G2298_;
  assign new_G2276_ = new_G2290_ | new_G2292_;
  assign new_G2277_ = new_G2300_ | new_G2299_;
  assign new_G2278_ = new_G2294_ | new_G2293_;
  assign new_G2279_ = ~new_G2302_ | ~new_G2301_;
  assign new_G2280_ = ~new_G2303_ & new_G2304_;
  assign new_G2281_ = new_G2303_ & ~new_G2304_;
  assign new_G2282_ = ~G2250 & G2251;
  assign new_G2283_ = G2250 & ~G2251;
  assign new_G2284_ = ~new_G2266_ | new_G2276_;
  assign new_G2285_ = new_G2266_ & new_G2276_;
  assign new_G2286_ = ~new_G2266_ & ~new_G2276_;
  assign new_G2287_ = new_G2308_ | new_G2307_;
  assign new_G2288_ = G2254 | new_G2287_;
  assign new_G2289_ = new_G2312_ | new_G2311_;
  assign new_G2290_ = ~G2254 & new_G2289_;
  assign new_G2291_ = new_G2310_ | new_G2309_;
  assign new_G2292_ = G2254 & new_G2291_;
  assign new_G2293_ = G2252 & ~new_G2262_;
  assign new_G2294_ = ~G2252 & new_G2262_;
  assign new_G2295_ = ~G2251 | ~new_G2276_;
  assign new_G2296_ = new_G2262_ & new_G2295_;
  assign new_G2297_ = ~new_G2262_ & ~new_G2296_;
  assign new_G2298_ = new_G2262_ | new_G2295_;
  assign new_G2299_ = ~G2252 & G2253;
  assign new_G2300_ = G2252 & ~G2253;
  assign new_G2301_ = new_G2269_ | new_G2306_;
  assign new_G2302_ = ~new_G2269_ & ~new_G2305_;
  assign new_G2303_ = G2252 | new_G2269_;
  assign new_G2304_ = G2252 | G2253;
  assign new_G2305_ = new_G2269_ & new_G2306_;
  assign new_G2306_ = ~G2251 | ~new_G2276_;
  assign new_G2307_ = new_G2284_ & new_G2304_;
  assign new_G2308_ = ~new_G2284_ & ~new_G2304_;
  assign new_G2309_ = new_G2313_ | new_G2314_;
  assign new_G2310_ = ~G2255 & new_G2269_;
  assign new_G2311_ = new_G2315_ | new_G2316_;
  assign new_G2312_ = G2255 & new_G2269_;
  assign new_G2313_ = ~G2255 & ~new_G2269_;
  assign new_G2314_ = G2255 & ~new_G2269_;
  assign new_G2315_ = G2255 & ~new_G2269_;
  assign new_G2316_ = ~G2255 & new_G2269_;
  assign new_G2323_ = new_G2330_ & new_G2329_;
  assign new_G2324_ = new_G2332_ | new_G2331_;
  assign new_G2325_ = new_G2334_ | new_G2333_;
  assign new_G2326_ = new_G2336_ & new_G2335_;
  assign new_G2327_ = new_G2336_ & new_G2337_;
  assign new_G2328_ = new_G2329_ | new_G2338_;
  assign new_G2329_ = G2318 | new_G2341_;
  assign new_G2330_ = new_G2340_ | new_G2339_;
  assign new_G2331_ = new_G2345_ & new_G2344_;
  assign new_G2332_ = new_G2343_ & new_G2342_;
  assign new_G2333_ = new_G2348_ | new_G2347_;
  assign new_G2334_ = new_G2343_ & new_G2346_;
  assign new_G2335_ = G2318 | new_G2351_;
  assign new_G2336_ = new_G2350_ | new_G2349_;
  assign new_G2337_ = new_G2353_ | new_G2352_;
  assign new_G2338_ = ~new_G2329_ & new_G2355_;
  assign new_G2339_ = ~new_G2331_ & new_G2343_;
  assign new_G2340_ = new_G2331_ & ~new_G2343_;
  assign new_G2341_ = G2317 & ~G2318;
  assign new_G2342_ = ~new_G2364_ | ~new_G2365_;
  assign new_G2343_ = new_G2357_ | new_G2359_;
  assign new_G2344_ = new_G2367_ | new_G2366_;
  assign new_G2345_ = new_G2361_ | new_G2360_;
  assign new_G2346_ = ~new_G2369_ | ~new_G2368_;
  assign new_G2347_ = ~new_G2370_ & new_G2371_;
  assign new_G2348_ = new_G2370_ & ~new_G2371_;
  assign new_G2349_ = ~G2317 & G2318;
  assign new_G2350_ = G2317 & ~G2318;
  assign new_G2351_ = ~new_G2333_ | new_G2343_;
  assign new_G2352_ = new_G2333_ & new_G2343_;
  assign new_G2353_ = ~new_G2333_ & ~new_G2343_;
  assign new_G2354_ = new_G2375_ | new_G2374_;
  assign new_G2355_ = G2321 | new_G2354_;
  assign new_G2356_ = new_G2379_ | new_G2378_;
  assign new_G2357_ = ~G2321 & new_G2356_;
  assign new_G2358_ = new_G2377_ | new_G2376_;
  assign new_G2359_ = G2321 & new_G2358_;
  assign new_G2360_ = G2319 & ~new_G2329_;
  assign new_G2361_ = ~G2319 & new_G2329_;
  assign new_G2362_ = ~G2318 | ~new_G2343_;
  assign new_G2363_ = new_G2329_ & new_G2362_;
  assign new_G2364_ = ~new_G2329_ & ~new_G2363_;
  assign new_G2365_ = new_G2329_ | new_G2362_;
  assign new_G2366_ = ~G2319 & G2320;
  assign new_G2367_ = G2319 & ~G2320;
  assign new_G2368_ = new_G2336_ | new_G2373_;
  assign new_G2369_ = ~new_G2336_ & ~new_G2372_;
  assign new_G2370_ = G2319 | new_G2336_;
  assign new_G2371_ = G2319 | G2320;
  assign new_G2372_ = new_G2336_ & new_G2373_;
  assign new_G2373_ = ~G2318 | ~new_G2343_;
  assign new_G2374_ = new_G2351_ & new_G2371_;
  assign new_G2375_ = ~new_G2351_ & ~new_G2371_;
  assign new_G2376_ = new_G2380_ | new_G2381_;
  assign new_G2377_ = ~G2322 & new_G2336_;
  assign new_G2378_ = new_G2382_ | new_G2383_;
  assign new_G2379_ = G2322 & new_G2336_;
  assign new_G2380_ = ~G2322 & ~new_G2336_;
  assign new_G2381_ = G2322 & ~new_G2336_;
  assign new_G2382_ = G2322 & ~new_G2336_;
  assign new_G2383_ = ~G2322 & new_G2336_;
  assign new_G2390_ = new_G2397_ & new_G2396_;
  assign new_G2391_ = new_G2399_ | new_G2398_;
  assign new_G2392_ = new_G2401_ | new_G2400_;
  assign new_G2393_ = new_G2403_ & new_G2402_;
  assign new_G2394_ = new_G2403_ & new_G2404_;
  assign new_G2395_ = new_G2396_ | new_G2405_;
  assign new_G2396_ = G2385 | new_G2408_;
  assign new_G2397_ = new_G2407_ | new_G2406_;
  assign new_G2398_ = new_G2412_ & new_G2411_;
  assign new_G2399_ = new_G2410_ & new_G2409_;
  assign new_G2400_ = new_G2415_ | new_G2414_;
  assign new_G2401_ = new_G2410_ & new_G2413_;
  assign new_G2402_ = G2385 | new_G2418_;
  assign new_G2403_ = new_G2417_ | new_G2416_;
  assign new_G2404_ = new_G2420_ | new_G2419_;
  assign new_G2405_ = ~new_G2396_ & new_G2422_;
  assign new_G2406_ = ~new_G2398_ & new_G2410_;
  assign new_G2407_ = new_G2398_ & ~new_G2410_;
  assign new_G2408_ = G2384 & ~G2385;
  assign new_G2409_ = ~new_G2431_ | ~new_G2432_;
  assign new_G2410_ = new_G2424_ | new_G2426_;
  assign new_G2411_ = new_G2434_ | new_G2433_;
  assign new_G2412_ = new_G2428_ | new_G2427_;
  assign new_G2413_ = ~new_G2436_ | ~new_G2435_;
  assign new_G2414_ = ~new_G2437_ & new_G2438_;
  assign new_G2415_ = new_G2437_ & ~new_G2438_;
  assign new_G2416_ = ~G2384 & G2385;
  assign new_G2417_ = G2384 & ~G2385;
  assign new_G2418_ = ~new_G2400_ | new_G2410_;
  assign new_G2419_ = new_G2400_ & new_G2410_;
  assign new_G2420_ = ~new_G2400_ & ~new_G2410_;
  assign new_G2421_ = new_G2442_ | new_G2441_;
  assign new_G2422_ = G2388 | new_G2421_;
  assign new_G2423_ = new_G2446_ | new_G2445_;
  assign new_G2424_ = ~G2388 & new_G2423_;
  assign new_G2425_ = new_G2444_ | new_G2443_;
  assign new_G2426_ = G2388 & new_G2425_;
  assign new_G2427_ = G2386 & ~new_G2396_;
  assign new_G2428_ = ~G2386 & new_G2396_;
  assign new_G2429_ = ~G2385 | ~new_G2410_;
  assign new_G2430_ = new_G2396_ & new_G2429_;
  assign new_G2431_ = ~new_G2396_ & ~new_G2430_;
  assign new_G2432_ = new_G2396_ | new_G2429_;
  assign new_G2433_ = ~G2386 & G2387;
  assign new_G2434_ = G2386 & ~G2387;
  assign new_G2435_ = new_G2403_ | new_G2440_;
  assign new_G2436_ = ~new_G2403_ & ~new_G2439_;
  assign new_G2437_ = G2386 | new_G2403_;
  assign new_G2438_ = G2386 | G2387;
  assign new_G2439_ = new_G2403_ & new_G2440_;
  assign new_G2440_ = ~G2385 | ~new_G2410_;
  assign new_G2441_ = new_G2418_ & new_G2438_;
  assign new_G2442_ = ~new_G2418_ & ~new_G2438_;
  assign new_G2443_ = new_G2447_ | new_G2448_;
  assign new_G2444_ = ~G2389 & new_G2403_;
  assign new_G2445_ = new_G2449_ | new_G2450_;
  assign new_G2446_ = G2389 & new_G2403_;
  assign new_G2447_ = ~G2389 & ~new_G2403_;
  assign new_G2448_ = G2389 & ~new_G2403_;
  assign new_G2449_ = G2389 & ~new_G2403_;
  assign new_G2450_ = ~G2389 & new_G2403_;
  assign new_G2457_ = new_G2464_ & new_G2463_;
  assign new_G2458_ = new_G2466_ | new_G2465_;
  assign new_G2459_ = new_G2468_ | new_G2467_;
  assign new_G2460_ = new_G2470_ & new_G2469_;
  assign new_G2461_ = new_G2470_ & new_G2471_;
  assign new_G2462_ = new_G2463_ | new_G2472_;
  assign new_G2463_ = G2452 | new_G2475_;
  assign new_G2464_ = new_G2474_ | new_G2473_;
  assign new_G2465_ = new_G2479_ & new_G2478_;
  assign new_G2466_ = new_G2477_ & new_G2476_;
  assign new_G2467_ = new_G2482_ | new_G2481_;
  assign new_G2468_ = new_G2477_ & new_G2480_;
  assign new_G2469_ = G2452 | new_G2485_;
  assign new_G2470_ = new_G2484_ | new_G2483_;
  assign new_G2471_ = new_G2487_ | new_G2486_;
  assign new_G2472_ = ~new_G2463_ & new_G2489_;
  assign new_G2473_ = ~new_G2465_ & new_G2477_;
  assign new_G2474_ = new_G2465_ & ~new_G2477_;
  assign new_G2475_ = G2451 & ~G2452;
  assign new_G2476_ = ~new_G2498_ | ~new_G2499_;
  assign new_G2477_ = new_G2491_ | new_G2493_;
  assign new_G2478_ = new_G2501_ | new_G2500_;
  assign new_G2479_ = new_G2495_ | new_G2494_;
  assign new_G2480_ = ~new_G2503_ | ~new_G2502_;
  assign new_G2481_ = ~new_G2504_ & new_G2505_;
  assign new_G2482_ = new_G2504_ & ~new_G2505_;
  assign new_G2483_ = ~G2451 & G2452;
  assign new_G2484_ = G2451 & ~G2452;
  assign new_G2485_ = ~new_G2467_ | new_G2477_;
  assign new_G2486_ = new_G2467_ & new_G2477_;
  assign new_G2487_ = ~new_G2467_ & ~new_G2477_;
  assign new_G2488_ = new_G2509_ | new_G2508_;
  assign new_G2489_ = G2455 | new_G2488_;
  assign new_G2490_ = new_G2513_ | new_G2512_;
  assign new_G2491_ = ~G2455 & new_G2490_;
  assign new_G2492_ = new_G2511_ | new_G2510_;
  assign new_G2493_ = G2455 & new_G2492_;
  assign new_G2494_ = G2453 & ~new_G2463_;
  assign new_G2495_ = ~G2453 & new_G2463_;
  assign new_G2496_ = ~G2452 | ~new_G2477_;
  assign new_G2497_ = new_G2463_ & new_G2496_;
  assign new_G2498_ = ~new_G2463_ & ~new_G2497_;
  assign new_G2499_ = new_G2463_ | new_G2496_;
  assign new_G2500_ = ~G2453 & G2454;
  assign new_G2501_ = G2453 & ~G2454;
  assign new_G2502_ = new_G2470_ | new_G2507_;
  assign new_G2503_ = ~new_G2470_ & ~new_G2506_;
  assign new_G2504_ = G2453 | new_G2470_;
  assign new_G2505_ = G2453 | G2454;
  assign new_G2506_ = new_G2470_ & new_G2507_;
  assign new_G2507_ = ~G2452 | ~new_G2477_;
  assign new_G2508_ = new_G2485_ & new_G2505_;
  assign new_G2509_ = ~new_G2485_ & ~new_G2505_;
  assign new_G2510_ = new_G2514_ | new_G2515_;
  assign new_G2511_ = ~G2456 & new_G2470_;
  assign new_G2512_ = new_G2516_ | new_G2517_;
  assign new_G2513_ = G2456 & new_G2470_;
  assign new_G2514_ = ~G2456 & ~new_G2470_;
  assign new_G2515_ = G2456 & ~new_G2470_;
  assign new_G2516_ = G2456 & ~new_G2470_;
  assign new_G2517_ = ~G2456 & new_G2470_;
  assign new_G2524_ = new_G2531_ & new_G2530_;
  assign new_G2525_ = new_G2533_ | new_G2532_;
  assign new_G2526_ = new_G2535_ | new_G2534_;
  assign new_G2527_ = new_G2537_ & new_G2536_;
  assign new_G2528_ = new_G2537_ & new_G2538_;
  assign new_G2529_ = new_G2530_ | new_G2539_;
  assign new_G2530_ = G2519 | new_G2542_;
  assign new_G2531_ = new_G2541_ | new_G2540_;
  assign new_G2532_ = new_G2546_ & new_G2545_;
  assign new_G2533_ = new_G2544_ & new_G2543_;
  assign new_G2534_ = new_G2549_ | new_G2548_;
  assign new_G2535_ = new_G2544_ & new_G2547_;
  assign new_G2536_ = G2519 | new_G2552_;
  assign new_G2537_ = new_G2551_ | new_G2550_;
  assign new_G2538_ = new_G2554_ | new_G2553_;
  assign new_G2539_ = ~new_G2530_ & new_G2556_;
  assign new_G2540_ = ~new_G2532_ & new_G2544_;
  assign new_G2541_ = new_G2532_ & ~new_G2544_;
  assign new_G2542_ = G2518 & ~G2519;
  assign new_G2543_ = ~new_G2565_ | ~new_G2566_;
  assign new_G2544_ = new_G2558_ | new_G2560_;
  assign new_G2545_ = new_G2568_ | new_G2567_;
  assign new_G2546_ = new_G2562_ | new_G2561_;
  assign new_G2547_ = ~new_G2570_ | ~new_G2569_;
  assign new_G2548_ = ~new_G2571_ & new_G2572_;
  assign new_G2549_ = new_G2571_ & ~new_G2572_;
  assign new_G2550_ = ~G2518 & G2519;
  assign new_G2551_ = G2518 & ~G2519;
  assign new_G2552_ = ~new_G2534_ | new_G2544_;
  assign new_G2553_ = new_G2534_ & new_G2544_;
  assign new_G2554_ = ~new_G2534_ & ~new_G2544_;
  assign new_G2555_ = new_G2576_ | new_G2575_;
  assign new_G2556_ = G2522 | new_G2555_;
  assign new_G2557_ = new_G2580_ | new_G2579_;
  assign new_G2558_ = ~G2522 & new_G2557_;
  assign new_G2559_ = new_G2578_ | new_G2577_;
  assign new_G2560_ = G2522 & new_G2559_;
  assign new_G2561_ = G2520 & ~new_G2530_;
  assign new_G2562_ = ~G2520 & new_G2530_;
  assign new_G2563_ = ~G2519 | ~new_G2544_;
  assign new_G2564_ = new_G2530_ & new_G2563_;
  assign new_G2565_ = ~new_G2530_ & ~new_G2564_;
  assign new_G2566_ = new_G2530_ | new_G2563_;
  assign new_G2567_ = ~G2520 & G2521;
  assign new_G2568_ = G2520 & ~G2521;
  assign new_G2569_ = new_G2537_ | new_G2574_;
  assign new_G2570_ = ~new_G2537_ & ~new_G2573_;
  assign new_G2571_ = G2520 | new_G2537_;
  assign new_G2572_ = G2520 | G2521;
  assign new_G2573_ = new_G2537_ & new_G2574_;
  assign new_G2574_ = ~G2519 | ~new_G2544_;
  assign new_G2575_ = new_G2552_ & new_G2572_;
  assign new_G2576_ = ~new_G2552_ & ~new_G2572_;
  assign new_G2577_ = new_G2581_ | new_G2582_;
  assign new_G2578_ = ~G2523 & new_G2537_;
  assign new_G2579_ = new_G2583_ | new_G2584_;
  assign new_G2580_ = G2523 & new_G2537_;
  assign new_G2581_ = ~G2523 & ~new_G2537_;
  assign new_G2582_ = G2523 & ~new_G2537_;
  assign new_G2583_ = G2523 & ~new_G2537_;
  assign new_G2584_ = ~G2523 & new_G2537_;
  assign new_G2591_ = new_G2598_ & new_G2597_;
  assign new_G2592_ = new_G2600_ | new_G2599_;
  assign new_G2593_ = new_G2602_ | new_G2601_;
  assign new_G2594_ = new_G2604_ & new_G2603_;
  assign new_G2595_ = new_G2604_ & new_G2605_;
  assign new_G2596_ = new_G2597_ | new_G2606_;
  assign new_G2597_ = G2586 | new_G2609_;
  assign new_G2598_ = new_G2608_ | new_G2607_;
  assign new_G2599_ = new_G2613_ & new_G2612_;
  assign new_G2600_ = new_G2611_ & new_G2610_;
  assign new_G2601_ = new_G2616_ | new_G2615_;
  assign new_G2602_ = new_G2611_ & new_G2614_;
  assign new_G2603_ = G2586 | new_G2619_;
  assign new_G2604_ = new_G2618_ | new_G2617_;
  assign new_G2605_ = new_G2621_ | new_G2620_;
  assign new_G2606_ = ~new_G2597_ & new_G2623_;
  assign new_G2607_ = ~new_G2599_ & new_G2611_;
  assign new_G2608_ = new_G2599_ & ~new_G2611_;
  assign new_G2609_ = G2585 & ~G2586;
  assign new_G2610_ = ~new_G2632_ | ~new_G2633_;
  assign new_G2611_ = new_G2625_ | new_G2627_;
  assign new_G2612_ = new_G2635_ | new_G2634_;
  assign new_G2613_ = new_G2629_ | new_G2628_;
  assign new_G2614_ = ~new_G2637_ | ~new_G2636_;
  assign new_G2615_ = ~new_G2638_ & new_G2639_;
  assign new_G2616_ = new_G2638_ & ~new_G2639_;
  assign new_G2617_ = ~G2585 & G2586;
  assign new_G2618_ = G2585 & ~G2586;
  assign new_G2619_ = ~new_G2601_ | new_G2611_;
  assign new_G2620_ = new_G2601_ & new_G2611_;
  assign new_G2621_ = ~new_G2601_ & ~new_G2611_;
  assign new_G2622_ = new_G2643_ | new_G2642_;
  assign new_G2623_ = G2589 | new_G2622_;
  assign new_G2624_ = new_G2647_ | new_G2646_;
  assign new_G2625_ = ~G2589 & new_G2624_;
  assign new_G2626_ = new_G2645_ | new_G2644_;
  assign new_G2627_ = G2589 & new_G2626_;
  assign new_G2628_ = G2587 & ~new_G2597_;
  assign new_G2629_ = ~G2587 & new_G2597_;
  assign new_G2630_ = ~G2586 | ~new_G2611_;
  assign new_G2631_ = new_G2597_ & new_G2630_;
  assign new_G2632_ = ~new_G2597_ & ~new_G2631_;
  assign new_G2633_ = new_G2597_ | new_G2630_;
  assign new_G2634_ = ~G2587 & G2588;
  assign new_G2635_ = G2587 & ~G2588;
  assign new_G2636_ = new_G2604_ | new_G2641_;
  assign new_G2637_ = ~new_G2604_ & ~new_G2640_;
  assign new_G2638_ = G2587 | new_G2604_;
  assign new_G2639_ = G2587 | G2588;
  assign new_G2640_ = new_G2604_ & new_G2641_;
  assign new_G2641_ = ~G2586 | ~new_G2611_;
  assign new_G2642_ = new_G2619_ & new_G2639_;
  assign new_G2643_ = ~new_G2619_ & ~new_G2639_;
  assign new_G2644_ = new_G2648_ | new_G2649_;
  assign new_G2645_ = ~G2590 & new_G2604_;
  assign new_G2646_ = new_G2650_ | new_G2651_;
  assign new_G2647_ = G2590 & new_G2604_;
  assign new_G2648_ = ~G2590 & ~new_G2604_;
  assign new_G2649_ = G2590 & ~new_G2604_;
  assign new_G2650_ = G2590 & ~new_G2604_;
  assign new_G2651_ = ~G2590 & new_G2604_;
  assign new_G2658_ = new_G2665_ & new_G2664_;
  assign new_G2659_ = new_G2667_ | new_G2666_;
  assign new_G2660_ = new_G2669_ | new_G2668_;
  assign new_G2661_ = new_G2671_ & new_G2670_;
  assign new_G2662_ = new_G2671_ & new_G2672_;
  assign new_G2663_ = new_G2664_ | new_G2673_;
  assign new_G2664_ = G2653 | new_G2676_;
  assign new_G2665_ = new_G2675_ | new_G2674_;
  assign new_G2666_ = new_G2680_ & new_G2679_;
  assign new_G2667_ = new_G2678_ & new_G2677_;
  assign new_G2668_ = new_G2683_ | new_G2682_;
  assign new_G2669_ = new_G2678_ & new_G2681_;
  assign new_G2670_ = G2653 | new_G2686_;
  assign new_G2671_ = new_G2685_ | new_G2684_;
  assign new_G2672_ = new_G2688_ | new_G2687_;
  assign new_G2673_ = ~new_G2664_ & new_G2690_;
  assign new_G2674_ = ~new_G2666_ & new_G2678_;
  assign new_G2675_ = new_G2666_ & ~new_G2678_;
  assign new_G2676_ = G2652 & ~G2653;
  assign new_G2677_ = ~new_G2699_ | ~new_G2700_;
  assign new_G2678_ = new_G2692_ | new_G2694_;
  assign new_G2679_ = new_G2702_ | new_G2701_;
  assign new_G2680_ = new_G2696_ | new_G2695_;
  assign new_G2681_ = ~new_G2704_ | ~new_G2703_;
  assign new_G2682_ = ~new_G2705_ & new_G2706_;
  assign new_G2683_ = new_G2705_ & ~new_G2706_;
  assign new_G2684_ = ~G2652 & G2653;
  assign new_G2685_ = G2652 & ~G2653;
  assign new_G2686_ = ~new_G2668_ | new_G2678_;
  assign new_G2687_ = new_G2668_ & new_G2678_;
  assign new_G2688_ = ~new_G2668_ & ~new_G2678_;
  assign new_G2689_ = new_G2710_ | new_G2709_;
  assign new_G2690_ = G2656 | new_G2689_;
  assign new_G2691_ = new_G2714_ | new_G2713_;
  assign new_G2692_ = ~G2656 & new_G2691_;
  assign new_G2693_ = new_G2712_ | new_G2711_;
  assign new_G2694_ = G2656 & new_G2693_;
  assign new_G2695_ = G2654 & ~new_G2664_;
  assign new_G2696_ = ~G2654 & new_G2664_;
  assign new_G2697_ = ~G2653 | ~new_G2678_;
  assign new_G2698_ = new_G2664_ & new_G2697_;
  assign new_G2699_ = ~new_G2664_ & ~new_G2698_;
  assign new_G2700_ = new_G2664_ | new_G2697_;
  assign new_G2701_ = ~G2654 & G2655;
  assign new_G2702_ = G2654 & ~G2655;
  assign new_G2703_ = new_G2671_ | new_G2708_;
  assign new_G2704_ = ~new_G2671_ & ~new_G2707_;
  assign new_G2705_ = G2654 | new_G2671_;
  assign new_G2706_ = G2654 | G2655;
  assign new_G2707_ = new_G2671_ & new_G2708_;
  assign new_G2708_ = ~G2653 | ~new_G2678_;
  assign new_G2709_ = new_G2686_ & new_G2706_;
  assign new_G2710_ = ~new_G2686_ & ~new_G2706_;
  assign new_G2711_ = new_G2715_ | new_G2716_;
  assign new_G2712_ = ~G2657 & new_G2671_;
  assign new_G2713_ = new_G2717_ | new_G2718_;
  assign new_G2714_ = G2657 & new_G2671_;
  assign new_G2715_ = ~G2657 & ~new_G2671_;
  assign new_G2716_ = G2657 & ~new_G2671_;
  assign new_G2717_ = G2657 & ~new_G2671_;
  assign new_G2718_ = ~G2657 & new_G2671_;
  assign new_G2725_ = new_G2732_ & new_G2731_;
  assign new_G2726_ = new_G2734_ | new_G2733_;
  assign new_G2727_ = new_G2736_ | new_G2735_;
  assign new_G2728_ = new_G2738_ & new_G2737_;
  assign new_G2729_ = new_G2738_ & new_G2739_;
  assign new_G2730_ = new_G2731_ | new_G2740_;
  assign new_G2731_ = G2720 | new_G2743_;
  assign new_G2732_ = new_G2742_ | new_G2741_;
  assign new_G2733_ = new_G2747_ & new_G2746_;
  assign new_G2734_ = new_G2745_ & new_G2744_;
  assign new_G2735_ = new_G2750_ | new_G2749_;
  assign new_G2736_ = new_G2745_ & new_G2748_;
  assign new_G2737_ = G2720 | new_G2753_;
  assign new_G2738_ = new_G2752_ | new_G2751_;
  assign new_G2739_ = new_G2755_ | new_G2754_;
  assign new_G2740_ = ~new_G2731_ & new_G2757_;
  assign new_G2741_ = ~new_G2733_ & new_G2745_;
  assign new_G2742_ = new_G2733_ & ~new_G2745_;
  assign new_G2743_ = G2719 & ~G2720;
  assign new_G2744_ = ~new_G2766_ | ~new_G2767_;
  assign new_G2745_ = new_G2759_ | new_G2761_;
  assign new_G2746_ = new_G2769_ | new_G2768_;
  assign new_G2747_ = new_G2763_ | new_G2762_;
  assign new_G2748_ = ~new_G2771_ | ~new_G2770_;
  assign new_G2749_ = ~new_G2772_ & new_G2773_;
  assign new_G2750_ = new_G2772_ & ~new_G2773_;
  assign new_G2751_ = ~G2719 & G2720;
  assign new_G2752_ = G2719 & ~G2720;
  assign new_G2753_ = ~new_G2735_ | new_G2745_;
  assign new_G2754_ = new_G2735_ & new_G2745_;
  assign new_G2755_ = ~new_G2735_ & ~new_G2745_;
  assign new_G2756_ = new_G2777_ | new_G2776_;
  assign new_G2757_ = G2723 | new_G2756_;
  assign new_G2758_ = new_G2781_ | new_G2780_;
  assign new_G2759_ = ~G2723 & new_G2758_;
  assign new_G2760_ = new_G2779_ | new_G2778_;
  assign new_G2761_ = G2723 & new_G2760_;
  assign new_G2762_ = G2721 & ~new_G2731_;
  assign new_G2763_ = ~G2721 & new_G2731_;
  assign new_G2764_ = ~G2720 | ~new_G2745_;
  assign new_G2765_ = new_G2731_ & new_G2764_;
  assign new_G2766_ = ~new_G2731_ & ~new_G2765_;
  assign new_G2767_ = new_G2731_ | new_G2764_;
  assign new_G2768_ = ~G2721 & G2722;
  assign new_G2769_ = G2721 & ~G2722;
  assign new_G2770_ = new_G2738_ | new_G2775_;
  assign new_G2771_ = ~new_G2738_ & ~new_G2774_;
  assign new_G2772_ = G2721 | new_G2738_;
  assign new_G2773_ = G2721 | G2722;
  assign new_G2774_ = new_G2738_ & new_G2775_;
  assign new_G2775_ = ~G2720 | ~new_G2745_;
  assign new_G2776_ = new_G2753_ & new_G2773_;
  assign new_G2777_ = ~new_G2753_ & ~new_G2773_;
  assign new_G2778_ = new_G2782_ | new_G2783_;
  assign new_G2779_ = ~G2724 & new_G2738_;
  assign new_G2780_ = new_G2784_ | new_G2785_;
  assign new_G2781_ = G2724 & new_G2738_;
  assign new_G2782_ = ~G2724 & ~new_G2738_;
  assign new_G2783_ = G2724 & ~new_G2738_;
  assign new_G2784_ = G2724 & ~new_G2738_;
  assign new_G2785_ = ~G2724 & new_G2738_;
  assign new_G2792_ = new_G2799_ & new_G2798_;
  assign new_G2793_ = new_G2801_ | new_G2800_;
  assign new_G2794_ = new_G2803_ | new_G2802_;
  assign new_G2795_ = new_G2805_ & new_G2804_;
  assign new_G2796_ = new_G2805_ & new_G2806_;
  assign new_G2797_ = new_G2798_ | new_G2807_;
  assign new_G2798_ = G2787 | new_G2810_;
  assign new_G2799_ = new_G2809_ | new_G2808_;
  assign new_G2800_ = new_G2814_ & new_G2813_;
  assign new_G2801_ = new_G2812_ & new_G2811_;
  assign new_G2802_ = new_G2817_ | new_G2816_;
  assign new_G2803_ = new_G2812_ & new_G2815_;
  assign new_G2804_ = G2787 | new_G2820_;
  assign new_G2805_ = new_G2819_ | new_G2818_;
  assign new_G2806_ = new_G2822_ | new_G2821_;
  assign new_G2807_ = ~new_G2798_ & new_G2824_;
  assign new_G2808_ = ~new_G2800_ & new_G2812_;
  assign new_G2809_ = new_G2800_ & ~new_G2812_;
  assign new_G2810_ = G2786 & ~G2787;
  assign new_G2811_ = ~new_G2833_ | ~new_G2834_;
  assign new_G2812_ = new_G2826_ | new_G2828_;
  assign new_G2813_ = new_G2836_ | new_G2835_;
  assign new_G2814_ = new_G2830_ | new_G2829_;
  assign new_G2815_ = ~new_G2838_ | ~new_G2837_;
  assign new_G2816_ = ~new_G2839_ & new_G2840_;
  assign new_G2817_ = new_G2839_ & ~new_G2840_;
  assign new_G2818_ = ~G2786 & G2787;
  assign new_G2819_ = G2786 & ~G2787;
  assign new_G2820_ = ~new_G2802_ | new_G2812_;
  assign new_G2821_ = new_G2802_ & new_G2812_;
  assign new_G2822_ = ~new_G2802_ & ~new_G2812_;
  assign new_G2823_ = new_G2844_ | new_G2843_;
  assign new_G2824_ = G2790 | new_G2823_;
  assign new_G2825_ = new_G2848_ | new_G2847_;
  assign new_G2826_ = ~G2790 & new_G2825_;
  assign new_G2827_ = new_G2846_ | new_G2845_;
  assign new_G2828_ = G2790 & new_G2827_;
  assign new_G2829_ = G2788 & ~new_G2798_;
  assign new_G2830_ = ~G2788 & new_G2798_;
  assign new_G2831_ = ~G2787 | ~new_G2812_;
  assign new_G2832_ = new_G2798_ & new_G2831_;
  assign new_G2833_ = ~new_G2798_ & ~new_G2832_;
  assign new_G2834_ = new_G2798_ | new_G2831_;
  assign new_G2835_ = ~G2788 & G2789;
  assign new_G2836_ = G2788 & ~G2789;
  assign new_G2837_ = new_G2805_ | new_G2842_;
  assign new_G2838_ = ~new_G2805_ & ~new_G2841_;
  assign new_G2839_ = G2788 | new_G2805_;
  assign new_G2840_ = G2788 | G2789;
  assign new_G2841_ = new_G2805_ & new_G2842_;
  assign new_G2842_ = ~G2787 | ~new_G2812_;
  assign new_G2843_ = new_G2820_ & new_G2840_;
  assign new_G2844_ = ~new_G2820_ & ~new_G2840_;
  assign new_G2845_ = new_G2849_ | new_G2850_;
  assign new_G2846_ = ~G2791 & new_G2805_;
  assign new_G2847_ = new_G2851_ | new_G2852_;
  assign new_G2848_ = G2791 & new_G2805_;
  assign new_G2849_ = ~G2791 & ~new_G2805_;
  assign new_G2850_ = G2791 & ~new_G2805_;
  assign new_G2851_ = G2791 & ~new_G2805_;
  assign new_G2852_ = ~G2791 & new_G2805_;
  assign new_G2859_ = new_G2866_ & new_G2865_;
  assign new_G2860_ = new_G2868_ | new_G2867_;
  assign new_G2861_ = new_G2870_ | new_G2869_;
  assign new_G2862_ = new_G2872_ & new_G2871_;
  assign new_G2863_ = new_G2872_ & new_G2873_;
  assign new_G2864_ = new_G2865_ | new_G2874_;
  assign new_G2865_ = G2854 | new_G2877_;
  assign new_G2866_ = new_G2876_ | new_G2875_;
  assign new_G2867_ = new_G2881_ & new_G2880_;
  assign new_G2868_ = new_G2879_ & new_G2878_;
  assign new_G2869_ = new_G2884_ | new_G2883_;
  assign new_G2870_ = new_G2879_ & new_G2882_;
  assign new_G2871_ = G2854 | new_G2887_;
  assign new_G2872_ = new_G2886_ | new_G2885_;
  assign new_G2873_ = new_G2889_ | new_G2888_;
  assign new_G2874_ = ~new_G2865_ & new_G2891_;
  assign new_G2875_ = ~new_G2867_ & new_G2879_;
  assign new_G2876_ = new_G2867_ & ~new_G2879_;
  assign new_G2877_ = G2853 & ~G2854;
  assign new_G2878_ = ~new_G2900_ | ~new_G2901_;
  assign new_G2879_ = new_G2893_ | new_G2895_;
  assign new_G2880_ = new_G2903_ | new_G2902_;
  assign new_G2881_ = new_G2897_ | new_G2896_;
  assign new_G2882_ = ~new_G2905_ | ~new_G2904_;
  assign new_G2883_ = ~new_G2906_ & new_G2907_;
  assign new_G2884_ = new_G2906_ & ~new_G2907_;
  assign new_G2885_ = ~G2853 & G2854;
  assign new_G2886_ = G2853 & ~G2854;
  assign new_G2887_ = ~new_G2869_ | new_G2879_;
  assign new_G2888_ = new_G2869_ & new_G2879_;
  assign new_G2889_ = ~new_G2869_ & ~new_G2879_;
  assign new_G2890_ = new_G2911_ | new_G2910_;
  assign new_G2891_ = G2857 | new_G2890_;
  assign new_G2892_ = new_G2915_ | new_G2914_;
  assign new_G2893_ = ~G2857 & new_G2892_;
  assign new_G2894_ = new_G2913_ | new_G2912_;
  assign new_G2895_ = G2857 & new_G2894_;
  assign new_G2896_ = G2855 & ~new_G2865_;
  assign new_G2897_ = ~G2855 & new_G2865_;
  assign new_G2898_ = ~G2854 | ~new_G2879_;
  assign new_G2899_ = new_G2865_ & new_G2898_;
  assign new_G2900_ = ~new_G2865_ & ~new_G2899_;
  assign new_G2901_ = new_G2865_ | new_G2898_;
  assign new_G2902_ = ~G2855 & G2856;
  assign new_G2903_ = G2855 & ~G2856;
  assign new_G2904_ = new_G2872_ | new_G2909_;
  assign new_G2905_ = ~new_G2872_ & ~new_G2908_;
  assign new_G2906_ = G2855 | new_G2872_;
  assign new_G2907_ = G2855 | G2856;
  assign new_G2908_ = new_G2872_ & new_G2909_;
  assign new_G2909_ = ~G2854 | ~new_G2879_;
  assign new_G2910_ = new_G2887_ & new_G2907_;
  assign new_G2911_ = ~new_G2887_ & ~new_G2907_;
  assign new_G2912_ = new_G2916_ | new_G2917_;
  assign new_G2913_ = ~G2858 & new_G2872_;
  assign new_G2914_ = new_G2918_ | new_G2919_;
  assign new_G2915_ = G2858 & new_G2872_;
  assign new_G2916_ = ~G2858 & ~new_G2872_;
  assign new_G2917_ = G2858 & ~new_G2872_;
  assign new_G2918_ = G2858 & ~new_G2872_;
  assign new_G2919_ = ~G2858 & new_G2872_;
  assign new_G2926_ = new_G2933_ & new_G2932_;
  assign new_G2927_ = new_G2935_ | new_G2934_;
  assign new_G2928_ = new_G2937_ | new_G2936_;
  assign new_G2929_ = new_G2939_ & new_G2938_;
  assign new_G2930_ = new_G2939_ & new_G2940_;
  assign new_G2931_ = new_G2932_ | new_G2941_;
  assign new_G2932_ = G2921 | new_G2944_;
  assign new_G2933_ = new_G2943_ | new_G2942_;
  assign new_G2934_ = new_G2948_ & new_G2947_;
  assign new_G2935_ = new_G2946_ & new_G2945_;
  assign new_G2936_ = new_G2951_ | new_G2950_;
  assign new_G2937_ = new_G2946_ & new_G2949_;
  assign new_G2938_ = G2921 | new_G2954_;
  assign new_G2939_ = new_G2953_ | new_G2952_;
  assign new_G2940_ = new_G2956_ | new_G2955_;
  assign new_G2941_ = ~new_G2932_ & new_G2958_;
  assign new_G2942_ = ~new_G2934_ & new_G2946_;
  assign new_G2943_ = new_G2934_ & ~new_G2946_;
  assign new_G2944_ = G2920 & ~G2921;
  assign new_G2945_ = ~new_G2967_ | ~new_G2968_;
  assign new_G2946_ = new_G2960_ | new_G2962_;
  assign new_G2947_ = new_G2970_ | new_G2969_;
  assign new_G2948_ = new_G2964_ | new_G2963_;
  assign new_G2949_ = ~new_G2972_ | ~new_G2971_;
  assign new_G2950_ = ~new_G2973_ & new_G2974_;
  assign new_G2951_ = new_G2973_ & ~new_G2974_;
  assign new_G2952_ = ~G2920 & G2921;
  assign new_G2953_ = G2920 & ~G2921;
  assign new_G2954_ = ~new_G2936_ | new_G2946_;
  assign new_G2955_ = new_G2936_ & new_G2946_;
  assign new_G2956_ = ~new_G2936_ & ~new_G2946_;
  assign new_G2957_ = new_G2978_ | new_G2977_;
  assign new_G2958_ = G2924 | new_G2957_;
  assign new_G2959_ = new_G2982_ | new_G2981_;
  assign new_G2960_ = ~G2924 & new_G2959_;
  assign new_G2961_ = new_G2980_ | new_G2979_;
  assign new_G2962_ = G2924 & new_G2961_;
  assign new_G2963_ = G2922 & ~new_G2932_;
  assign new_G2964_ = ~G2922 & new_G2932_;
  assign new_G2965_ = ~G2921 | ~new_G2946_;
  assign new_G2966_ = new_G2932_ & new_G2965_;
  assign new_G2967_ = ~new_G2932_ & ~new_G2966_;
  assign new_G2968_ = new_G2932_ | new_G2965_;
  assign new_G2969_ = ~G2922 & G2923;
  assign new_G2970_ = G2922 & ~G2923;
  assign new_G2971_ = new_G2939_ | new_G2976_;
  assign new_G2972_ = ~new_G2939_ & ~new_G2975_;
  assign new_G2973_ = G2922 | new_G2939_;
  assign new_G2974_ = G2922 | G2923;
  assign new_G2975_ = new_G2939_ & new_G2976_;
  assign new_G2976_ = ~G2921 | ~new_G2946_;
  assign new_G2977_ = new_G2954_ & new_G2974_;
  assign new_G2978_ = ~new_G2954_ & ~new_G2974_;
  assign new_G2979_ = new_G2983_ | new_G2984_;
  assign new_G2980_ = ~G2925 & new_G2939_;
  assign new_G2981_ = new_G2985_ | new_G2986_;
  assign new_G2982_ = G2925 & new_G2939_;
  assign new_G2983_ = ~G2925 & ~new_G2939_;
  assign new_G2984_ = G2925 & ~new_G2939_;
  assign new_G2985_ = G2925 & ~new_G2939_;
  assign new_G2986_ = ~G2925 & new_G2939_;
  assign new_G2993_ = new_G3000_ & new_G2999_;
  assign new_G2994_ = new_G3002_ | new_G3001_;
  assign new_G2995_ = new_G3004_ | new_G3003_;
  assign new_G2996_ = new_G3006_ & new_G3005_;
  assign new_G2997_ = new_G3006_ & new_G3007_;
  assign new_G2998_ = new_G2999_ | new_G3008_;
  assign new_G2999_ = G2988 | new_G3011_;
  assign new_G3000_ = new_G3010_ | new_G3009_;
  assign new_G3001_ = new_G3015_ & new_G3014_;
  assign new_G3002_ = new_G3013_ & new_G3012_;
  assign new_G3003_ = new_G3018_ | new_G3017_;
  assign new_G3004_ = new_G3013_ & new_G3016_;
  assign new_G3005_ = G2988 | new_G3021_;
  assign new_G3006_ = new_G3020_ | new_G3019_;
  assign new_G3007_ = new_G3023_ | new_G3022_;
  assign new_G3008_ = ~new_G2999_ & new_G3025_;
  assign new_G3009_ = ~new_G3001_ & new_G3013_;
  assign new_G3010_ = new_G3001_ & ~new_G3013_;
  assign new_G3011_ = G2987 & ~G2988;
  assign new_G3012_ = ~new_G3034_ | ~new_G3035_;
  assign new_G3013_ = new_G3027_ | new_G3029_;
  assign new_G3014_ = new_G3037_ | new_G3036_;
  assign new_G3015_ = new_G3031_ | new_G3030_;
  assign new_G3016_ = ~new_G3039_ | ~new_G3038_;
  assign new_G3017_ = ~new_G3040_ & new_G3041_;
  assign new_G3018_ = new_G3040_ & ~new_G3041_;
  assign new_G3019_ = ~G2987 & G2988;
  assign new_G3020_ = G2987 & ~G2988;
  assign new_G3021_ = ~new_G3003_ | new_G3013_;
  assign new_G3022_ = new_G3003_ & new_G3013_;
  assign new_G3023_ = ~new_G3003_ & ~new_G3013_;
  assign new_G3024_ = new_G3045_ | new_G3044_;
  assign new_G3025_ = G2991 | new_G3024_;
  assign new_G3026_ = new_G3049_ | new_G3048_;
  assign new_G3027_ = ~G2991 & new_G3026_;
  assign new_G3028_ = new_G3047_ | new_G3046_;
  assign new_G3029_ = G2991 & new_G3028_;
  assign new_G3030_ = G2989 & ~new_G2999_;
  assign new_G3031_ = ~G2989 & new_G2999_;
  assign new_G3032_ = ~G2988 | ~new_G3013_;
  assign new_G3033_ = new_G2999_ & new_G3032_;
  assign new_G3034_ = ~new_G2999_ & ~new_G3033_;
  assign new_G3035_ = new_G2999_ | new_G3032_;
  assign new_G3036_ = ~G2989 & G2990;
  assign new_G3037_ = G2989 & ~G2990;
  assign new_G3038_ = new_G3006_ | new_G3043_;
  assign new_G3039_ = ~new_G3006_ & ~new_G3042_;
  assign new_G3040_ = G2989 | new_G3006_;
  assign new_G3041_ = G2989 | G2990;
  assign new_G3042_ = new_G3006_ & new_G3043_;
  assign new_G3043_ = ~G2988 | ~new_G3013_;
  assign new_G3044_ = new_G3021_ & new_G3041_;
  assign new_G3045_ = ~new_G3021_ & ~new_G3041_;
  assign new_G3046_ = new_G3050_ | new_G3051_;
  assign new_G3047_ = ~G2992 & new_G3006_;
  assign new_G3048_ = new_G3052_ | new_G3053_;
  assign new_G3049_ = G2992 & new_G3006_;
  assign new_G3050_ = ~G2992 & ~new_G3006_;
  assign new_G3051_ = G2992 & ~new_G3006_;
  assign new_G3052_ = G2992 & ~new_G3006_;
  assign new_G3053_ = ~G2992 & new_G3006_;
  assign new_G3060_ = new_G3067_ & new_G3066_;
  assign new_G3061_ = new_G3069_ | new_G3068_;
  assign new_G3062_ = new_G3071_ | new_G3070_;
  assign new_G3063_ = new_G3073_ & new_G3072_;
  assign new_G3064_ = new_G3073_ & new_G3074_;
  assign new_G3065_ = new_G3066_ | new_G3075_;
  assign new_G3066_ = G3055 | new_G3078_;
  assign new_G3067_ = new_G3077_ | new_G3076_;
  assign new_G3068_ = new_G3082_ & new_G3081_;
  assign new_G3069_ = new_G3080_ & new_G3079_;
  assign new_G3070_ = new_G3085_ | new_G3084_;
  assign new_G3071_ = new_G3080_ & new_G3083_;
  assign new_G3072_ = G3055 | new_G3088_;
  assign new_G3073_ = new_G3087_ | new_G3086_;
  assign new_G3074_ = new_G3090_ | new_G3089_;
  assign new_G3075_ = ~new_G3066_ & new_G3092_;
  assign new_G3076_ = ~new_G3068_ & new_G3080_;
  assign new_G3077_ = new_G3068_ & ~new_G3080_;
  assign new_G3078_ = G3054 & ~G3055;
  assign new_G3079_ = ~new_G3101_ | ~new_G3102_;
  assign new_G3080_ = new_G3094_ | new_G3096_;
  assign new_G3081_ = new_G3104_ | new_G3103_;
  assign new_G3082_ = new_G3098_ | new_G3097_;
  assign new_G3083_ = ~new_G3106_ | ~new_G3105_;
  assign new_G3084_ = ~new_G3107_ & new_G3108_;
  assign new_G3085_ = new_G3107_ & ~new_G3108_;
  assign new_G3086_ = ~G3054 & G3055;
  assign new_G3087_ = G3054 & ~G3055;
  assign new_G3088_ = ~new_G3070_ | new_G3080_;
  assign new_G3089_ = new_G3070_ & new_G3080_;
  assign new_G3090_ = ~new_G3070_ & ~new_G3080_;
  assign new_G3091_ = new_G3112_ | new_G3111_;
  assign new_G3092_ = G3058 | new_G3091_;
  assign new_G3093_ = new_G3116_ | new_G3115_;
  assign new_G3094_ = ~G3058 & new_G3093_;
  assign new_G3095_ = new_G3114_ | new_G3113_;
  assign new_G3096_ = G3058 & new_G3095_;
  assign new_G3097_ = G3056 & ~new_G3066_;
  assign new_G3098_ = ~G3056 & new_G3066_;
  assign new_G3099_ = ~G3055 | ~new_G3080_;
  assign new_G3100_ = new_G3066_ & new_G3099_;
  assign new_G3101_ = ~new_G3066_ & ~new_G3100_;
  assign new_G3102_ = new_G3066_ | new_G3099_;
  assign new_G3103_ = ~G3056 & G3057;
  assign new_G3104_ = G3056 & ~G3057;
  assign new_G3105_ = new_G3073_ | new_G3110_;
  assign new_G3106_ = ~new_G3073_ & ~new_G3109_;
  assign new_G3107_ = G3056 | new_G3073_;
  assign new_G3108_ = G3056 | G3057;
  assign new_G3109_ = new_G3073_ & new_G3110_;
  assign new_G3110_ = ~G3055 | ~new_G3080_;
  assign new_G3111_ = new_G3088_ & new_G3108_;
  assign new_G3112_ = ~new_G3088_ & ~new_G3108_;
  assign new_G3113_ = new_G3117_ | new_G3118_;
  assign new_G3114_ = ~G3059 & new_G3073_;
  assign new_G3115_ = new_G3119_ | new_G3120_;
  assign new_G3116_ = G3059 & new_G3073_;
  assign new_G3117_ = ~G3059 & ~new_G3073_;
  assign new_G3118_ = G3059 & ~new_G3073_;
  assign new_G3119_ = G3059 & ~new_G3073_;
  assign new_G3120_ = ~G3059 & new_G3073_;
  assign new_G3127_ = new_G3134_ & new_G3133_;
  assign new_G3128_ = new_G3136_ | new_G3135_;
  assign new_G3129_ = new_G3138_ | new_G3137_;
  assign new_G3130_ = new_G3140_ & new_G3139_;
  assign new_G3131_ = new_G3140_ & new_G3141_;
  assign new_G3132_ = new_G3133_ | new_G3142_;
  assign new_G3133_ = G3122 | new_G3145_;
  assign new_G3134_ = new_G3144_ | new_G3143_;
  assign new_G3135_ = new_G3149_ & new_G3148_;
  assign new_G3136_ = new_G3147_ & new_G3146_;
  assign new_G3137_ = new_G3152_ | new_G3151_;
  assign new_G3138_ = new_G3147_ & new_G3150_;
  assign new_G3139_ = G3122 | new_G3155_;
  assign new_G3140_ = new_G3154_ | new_G3153_;
  assign new_G3141_ = new_G3157_ | new_G3156_;
  assign new_G3142_ = ~new_G3133_ & new_G3159_;
  assign new_G3143_ = ~new_G3135_ & new_G3147_;
  assign new_G3144_ = new_G3135_ & ~new_G3147_;
  assign new_G3145_ = G3121 & ~G3122;
  assign new_G3146_ = ~new_G3168_ | ~new_G3169_;
  assign new_G3147_ = new_G3161_ | new_G3163_;
  assign new_G3148_ = new_G3171_ | new_G3170_;
  assign new_G3149_ = new_G3165_ | new_G3164_;
  assign new_G3150_ = ~new_G3173_ | ~new_G3172_;
  assign new_G3151_ = ~new_G3174_ & new_G3175_;
  assign new_G3152_ = new_G3174_ & ~new_G3175_;
  assign new_G3153_ = ~G3121 & G3122;
  assign new_G3154_ = G3121 & ~G3122;
  assign new_G3155_ = ~new_G3137_ | new_G3147_;
  assign new_G3156_ = new_G3137_ & new_G3147_;
  assign new_G3157_ = ~new_G3137_ & ~new_G3147_;
  assign new_G3158_ = new_G3179_ | new_G3178_;
  assign new_G3159_ = G3125 | new_G3158_;
  assign new_G3160_ = new_G3183_ | new_G3182_;
  assign new_G3161_ = ~G3125 & new_G3160_;
  assign new_G3162_ = new_G3181_ | new_G3180_;
  assign new_G3163_ = G3125 & new_G3162_;
  assign new_G3164_ = G3123 & ~new_G3133_;
  assign new_G3165_ = ~G3123 & new_G3133_;
  assign new_G3166_ = ~G3122 | ~new_G3147_;
  assign new_G3167_ = new_G3133_ & new_G3166_;
  assign new_G3168_ = ~new_G3133_ & ~new_G3167_;
  assign new_G3169_ = new_G3133_ | new_G3166_;
  assign new_G3170_ = ~G3123 & G3124;
  assign new_G3171_ = G3123 & ~G3124;
  assign new_G3172_ = new_G3140_ | new_G3177_;
  assign new_G3173_ = ~new_G3140_ & ~new_G3176_;
  assign new_G3174_ = G3123 | new_G3140_;
  assign new_G3175_ = G3123 | G3124;
  assign new_G3176_ = new_G3140_ & new_G3177_;
  assign new_G3177_ = ~G3122 | ~new_G3147_;
  assign new_G3178_ = new_G3155_ & new_G3175_;
  assign new_G3179_ = ~new_G3155_ & ~new_G3175_;
  assign new_G3180_ = new_G3184_ | new_G3185_;
  assign new_G3181_ = ~G3126 & new_G3140_;
  assign new_G3182_ = new_G3186_ | new_G3187_;
  assign new_G3183_ = G3126 & new_G3140_;
  assign new_G3184_ = ~G3126 & ~new_G3140_;
  assign new_G3185_ = G3126 & ~new_G3140_;
  assign new_G3186_ = G3126 & ~new_G3140_;
  assign new_G3187_ = ~G3126 & new_G3140_;
  assign new_G3194_ = new_G3201_ & new_G3200_;
  assign new_G3195_ = new_G3203_ | new_G3202_;
  assign new_G3196_ = new_G3205_ | new_G3204_;
  assign new_G3197_ = new_G3207_ & new_G3206_;
  assign new_G3198_ = new_G3207_ & new_G3208_;
  assign new_G3199_ = new_G3200_ | new_G3209_;
  assign new_G3200_ = G3189 | new_G3212_;
  assign new_G3201_ = new_G3211_ | new_G3210_;
  assign new_G3202_ = new_G3216_ & new_G3215_;
  assign new_G3203_ = new_G3214_ & new_G3213_;
  assign new_G3204_ = new_G3219_ | new_G3218_;
  assign new_G3205_ = new_G3214_ & new_G3217_;
  assign new_G3206_ = G3189 | new_G3222_;
  assign new_G3207_ = new_G3221_ | new_G3220_;
  assign new_G3208_ = new_G3224_ | new_G3223_;
  assign new_G3209_ = ~new_G3200_ & new_G3226_;
  assign new_G3210_ = ~new_G3202_ & new_G3214_;
  assign new_G3211_ = new_G3202_ & ~new_G3214_;
  assign new_G3212_ = G3188 & ~G3189;
  assign new_G3213_ = ~new_G3235_ | ~new_G3236_;
  assign new_G3214_ = new_G3228_ | new_G3230_;
  assign new_G3215_ = new_G3238_ | new_G3237_;
  assign new_G3216_ = new_G3232_ | new_G3231_;
  assign new_G3217_ = ~new_G3240_ | ~new_G3239_;
  assign new_G3218_ = ~new_G3241_ & new_G3242_;
  assign new_G3219_ = new_G3241_ & ~new_G3242_;
  assign new_G3220_ = ~G3188 & G3189;
  assign new_G3221_ = G3188 & ~G3189;
  assign new_G3222_ = ~new_G3204_ | new_G3214_;
  assign new_G3223_ = new_G3204_ & new_G3214_;
  assign new_G3224_ = ~new_G3204_ & ~new_G3214_;
  assign new_G3225_ = new_G3246_ | new_G3245_;
  assign new_G3226_ = G3192 | new_G3225_;
  assign new_G3227_ = new_G3250_ | new_G3249_;
  assign new_G3228_ = ~G3192 & new_G3227_;
  assign new_G3229_ = new_G3248_ | new_G3247_;
  assign new_G3230_ = G3192 & new_G3229_;
  assign new_G3231_ = G3190 & ~new_G3200_;
  assign new_G3232_ = ~G3190 & new_G3200_;
  assign new_G3233_ = ~G3189 | ~new_G3214_;
  assign new_G3234_ = new_G3200_ & new_G3233_;
  assign new_G3235_ = ~new_G3200_ & ~new_G3234_;
  assign new_G3236_ = new_G3200_ | new_G3233_;
  assign new_G3237_ = ~G3190 & G3191;
  assign new_G3238_ = G3190 & ~G3191;
  assign new_G3239_ = new_G3207_ | new_G3244_;
  assign new_G3240_ = ~new_G3207_ & ~new_G3243_;
  assign new_G3241_ = G3190 | new_G3207_;
  assign new_G3242_ = G3190 | G3191;
  assign new_G3243_ = new_G3207_ & new_G3244_;
  assign new_G3244_ = ~G3189 | ~new_G3214_;
  assign new_G3245_ = new_G3222_ & new_G3242_;
  assign new_G3246_ = ~new_G3222_ & ~new_G3242_;
  assign new_G3247_ = new_G3251_ | new_G3252_;
  assign new_G3248_ = ~G3193 & new_G3207_;
  assign new_G3249_ = new_G3253_ | new_G3254_;
  assign new_G3250_ = G3193 & new_G3207_;
  assign new_G3251_ = ~G3193 & ~new_G3207_;
  assign new_G3252_ = G3193 & ~new_G3207_;
  assign new_G3253_ = G3193 & ~new_G3207_;
  assign new_G3254_ = ~G3193 & new_G3207_;
  assign new_G3261_ = new_G3268_ & new_G3267_;
  assign new_G3262_ = new_G3270_ | new_G3269_;
  assign new_G3263_ = new_G3272_ | new_G3271_;
  assign new_G3264_ = new_G3274_ & new_G3273_;
  assign new_G3265_ = new_G3274_ & new_G3275_;
  assign new_G3266_ = new_G3267_ | new_G3276_;
  assign new_G3267_ = G3256 | new_G3279_;
  assign new_G3268_ = new_G3278_ | new_G3277_;
  assign new_G3269_ = new_G3283_ & new_G3282_;
  assign new_G3270_ = new_G3281_ & new_G3280_;
  assign new_G3271_ = new_G3286_ | new_G3285_;
  assign new_G3272_ = new_G3281_ & new_G3284_;
  assign new_G3273_ = G3256 | new_G3289_;
  assign new_G3274_ = new_G3288_ | new_G3287_;
  assign new_G3275_ = new_G3291_ | new_G3290_;
  assign new_G3276_ = ~new_G3267_ & new_G3293_;
  assign new_G3277_ = ~new_G3269_ & new_G3281_;
  assign new_G3278_ = new_G3269_ & ~new_G3281_;
  assign new_G3279_ = G3255 & ~G3256;
  assign new_G3280_ = ~new_G3302_ | ~new_G3303_;
  assign new_G3281_ = new_G3295_ | new_G3297_;
  assign new_G3282_ = new_G3305_ | new_G3304_;
  assign new_G3283_ = new_G3299_ | new_G3298_;
  assign new_G3284_ = ~new_G3307_ | ~new_G3306_;
  assign new_G3285_ = ~new_G3308_ & new_G3309_;
  assign new_G3286_ = new_G3308_ & ~new_G3309_;
  assign new_G3287_ = ~G3255 & G3256;
  assign new_G3288_ = G3255 & ~G3256;
  assign new_G3289_ = ~new_G3271_ | new_G3281_;
  assign new_G3290_ = new_G3271_ & new_G3281_;
  assign new_G3291_ = ~new_G3271_ & ~new_G3281_;
  assign new_G3292_ = new_G3313_ | new_G3312_;
  assign new_G3293_ = G3259 | new_G3292_;
  assign new_G3294_ = new_G3317_ | new_G3316_;
  assign new_G3295_ = ~G3259 & new_G3294_;
  assign new_G3296_ = new_G3315_ | new_G3314_;
  assign new_G3297_ = G3259 & new_G3296_;
  assign new_G3298_ = G3257 & ~new_G3267_;
  assign new_G3299_ = ~G3257 & new_G3267_;
  assign new_G3300_ = ~G3256 | ~new_G3281_;
  assign new_G3301_ = new_G3267_ & new_G3300_;
  assign new_G3302_ = ~new_G3267_ & ~new_G3301_;
  assign new_G3303_ = new_G3267_ | new_G3300_;
  assign new_G3304_ = ~G3257 & G3258;
  assign new_G3305_ = G3257 & ~G3258;
  assign new_G3306_ = new_G3274_ | new_G3311_;
  assign new_G3307_ = ~new_G3274_ & ~new_G3310_;
  assign new_G3308_ = G3257 | new_G3274_;
  assign new_G3309_ = G3257 | G3258;
  assign new_G3310_ = new_G3274_ & new_G3311_;
  assign new_G3311_ = ~G3256 | ~new_G3281_;
  assign new_G3312_ = new_G3289_ & new_G3309_;
  assign new_G3313_ = ~new_G3289_ & ~new_G3309_;
  assign new_G3314_ = new_G3318_ | new_G3319_;
  assign new_G3315_ = ~G3260 & new_G3274_;
  assign new_G3316_ = new_G3320_ | new_G3321_;
  assign new_G3317_ = G3260 & new_G3274_;
  assign new_G3318_ = ~G3260 & ~new_G3274_;
  assign new_G3319_ = G3260 & ~new_G3274_;
  assign new_G3320_ = G3260 & ~new_G3274_;
  assign new_G3321_ = ~G3260 & new_G3274_;
  assign new_G3328_ = new_G3335_ & new_G3334_;
  assign new_G3329_ = new_G3337_ | new_G3336_;
  assign new_G3330_ = new_G3339_ | new_G3338_;
  assign new_G3331_ = new_G3341_ & new_G3340_;
  assign new_G3332_ = new_G3341_ & new_G3342_;
  assign new_G3333_ = new_G3334_ | new_G3343_;
  assign new_G3334_ = G3323 | new_G3346_;
  assign new_G3335_ = new_G3345_ | new_G3344_;
  assign new_G3336_ = new_G3350_ & new_G3349_;
  assign new_G3337_ = new_G3348_ & new_G3347_;
  assign new_G3338_ = new_G3353_ | new_G3352_;
  assign new_G3339_ = new_G3348_ & new_G3351_;
  assign new_G3340_ = G3323 | new_G3356_;
  assign new_G3341_ = new_G3355_ | new_G3354_;
  assign new_G3342_ = new_G3358_ | new_G3357_;
  assign new_G3343_ = ~new_G3334_ & new_G3360_;
  assign new_G3344_ = ~new_G3336_ & new_G3348_;
  assign new_G3345_ = new_G3336_ & ~new_G3348_;
  assign new_G3346_ = G3322 & ~G3323;
  assign new_G3347_ = ~new_G3369_ | ~new_G3370_;
  assign new_G3348_ = new_G3362_ | new_G3364_;
  assign new_G3349_ = new_G3372_ | new_G3371_;
  assign new_G3350_ = new_G3366_ | new_G3365_;
  assign new_G3351_ = ~new_G3374_ | ~new_G3373_;
  assign new_G3352_ = ~new_G3375_ & new_G3376_;
  assign new_G3353_ = new_G3375_ & ~new_G3376_;
  assign new_G3354_ = ~G3322 & G3323;
  assign new_G3355_ = G3322 & ~G3323;
  assign new_G3356_ = ~new_G3338_ | new_G3348_;
  assign new_G3357_ = new_G3338_ & new_G3348_;
  assign new_G3358_ = ~new_G3338_ & ~new_G3348_;
  assign new_G3359_ = new_G3380_ | new_G3379_;
  assign new_G3360_ = G3326 | new_G3359_;
  assign new_G3361_ = new_G3384_ | new_G3383_;
  assign new_G3362_ = ~G3326 & new_G3361_;
  assign new_G3363_ = new_G3382_ | new_G3381_;
  assign new_G3364_ = G3326 & new_G3363_;
  assign new_G3365_ = G3324 & ~new_G3334_;
  assign new_G3366_ = ~G3324 & new_G3334_;
  assign new_G3367_ = ~G3323 | ~new_G3348_;
  assign new_G3368_ = new_G3334_ & new_G3367_;
  assign new_G3369_ = ~new_G3334_ & ~new_G3368_;
  assign new_G3370_ = new_G3334_ | new_G3367_;
  assign new_G3371_ = ~G3324 & G3325;
  assign new_G3372_ = G3324 & ~G3325;
  assign new_G3373_ = new_G3341_ | new_G3378_;
  assign new_G3374_ = ~new_G3341_ & ~new_G3377_;
  assign new_G3375_ = G3324 | new_G3341_;
  assign new_G3376_ = G3324 | G3325;
  assign new_G3377_ = new_G3341_ & new_G3378_;
  assign new_G3378_ = ~G3323 | ~new_G3348_;
  assign new_G3379_ = new_G3356_ & new_G3376_;
  assign new_G3380_ = ~new_G3356_ & ~new_G3376_;
  assign new_G3381_ = new_G3385_ | new_G3386_;
  assign new_G3382_ = ~G3327 & new_G3341_;
  assign new_G3383_ = new_G3387_ | new_G3388_;
  assign new_G3384_ = G3327 & new_G3341_;
  assign new_G3385_ = ~G3327 & ~new_G3341_;
  assign new_G3386_ = G3327 & ~new_G3341_;
  assign new_G3387_ = G3327 & ~new_G3341_;
  assign new_G3388_ = ~G3327 & new_G3341_;
  assign new_G3395_ = new_G3402_ & new_G3401_;
  assign new_G3396_ = new_G3404_ | new_G3403_;
  assign new_G3397_ = new_G3406_ | new_G3405_;
  assign new_G3398_ = new_G3408_ & new_G3407_;
  assign new_G3399_ = new_G3408_ & new_G3409_;
  assign new_G3400_ = new_G3401_ | new_G3410_;
  assign new_G3401_ = G3390 | new_G3413_;
  assign new_G3402_ = new_G3412_ | new_G3411_;
  assign new_G3403_ = new_G3417_ & new_G3416_;
  assign new_G3404_ = new_G3415_ & new_G3414_;
  assign new_G3405_ = new_G3420_ | new_G3419_;
  assign new_G3406_ = new_G3415_ & new_G3418_;
  assign new_G3407_ = G3390 | new_G3423_;
  assign new_G3408_ = new_G3422_ | new_G3421_;
  assign new_G3409_ = new_G3425_ | new_G3424_;
  assign new_G3410_ = ~new_G3401_ & new_G3427_;
  assign new_G3411_ = ~new_G3403_ & new_G3415_;
  assign new_G3412_ = new_G3403_ & ~new_G3415_;
  assign new_G3413_ = G3389 & ~G3390;
  assign new_G3414_ = ~new_G3436_ | ~new_G3437_;
  assign new_G3415_ = new_G3429_ | new_G3431_;
  assign new_G3416_ = new_G3439_ | new_G3438_;
  assign new_G3417_ = new_G3433_ | new_G3432_;
  assign new_G3418_ = ~new_G3441_ | ~new_G3440_;
  assign new_G3419_ = ~new_G3442_ & new_G3443_;
  assign new_G3420_ = new_G3442_ & ~new_G3443_;
  assign new_G3421_ = ~G3389 & G3390;
  assign new_G3422_ = G3389 & ~G3390;
  assign new_G3423_ = ~new_G3405_ | new_G3415_;
  assign new_G3424_ = new_G3405_ & new_G3415_;
  assign new_G3425_ = ~new_G3405_ & ~new_G3415_;
  assign new_G3426_ = new_G3447_ | new_G3446_;
  assign new_G3427_ = G3393 | new_G3426_;
  assign new_G3428_ = new_G3451_ | new_G3450_;
  assign new_G3429_ = ~G3393 & new_G3428_;
  assign new_G3430_ = new_G3449_ | new_G3448_;
  assign new_G3431_ = G3393 & new_G3430_;
  assign new_G3432_ = G3391 & ~new_G3401_;
  assign new_G3433_ = ~G3391 & new_G3401_;
  assign new_G3434_ = ~G3390 | ~new_G3415_;
  assign new_G3435_ = new_G3401_ & new_G3434_;
  assign new_G3436_ = ~new_G3401_ & ~new_G3435_;
  assign new_G3437_ = new_G3401_ | new_G3434_;
  assign new_G3438_ = ~G3391 & G3392;
  assign new_G3439_ = G3391 & ~G3392;
  assign new_G3440_ = new_G3408_ | new_G3445_;
  assign new_G3441_ = ~new_G3408_ & ~new_G3444_;
  assign new_G3442_ = G3391 | new_G3408_;
  assign new_G3443_ = G3391 | G3392;
  assign new_G3444_ = new_G3408_ & new_G3445_;
  assign new_G3445_ = ~G3390 | ~new_G3415_;
  assign new_G3446_ = new_G3423_ & new_G3443_;
  assign new_G3447_ = ~new_G3423_ & ~new_G3443_;
  assign new_G3448_ = new_G3452_ | new_G3453_;
  assign new_G3449_ = ~G3394 & new_G3408_;
  assign new_G3450_ = new_G3454_ | new_G3455_;
  assign new_G3451_ = G3394 & new_G3408_;
  assign new_G3452_ = ~G3394 & ~new_G3408_;
  assign new_G3453_ = G3394 & ~new_G3408_;
  assign new_G3454_ = G3394 & ~new_G3408_;
  assign new_G3455_ = ~G3394 & new_G3408_;
  assign new_G3462_ = new_G3469_ & new_G3468_;
  assign new_G3463_ = new_G3471_ | new_G3470_;
  assign new_G3464_ = new_G3473_ | new_G3472_;
  assign new_G3465_ = new_G3475_ & new_G3474_;
  assign new_G3466_ = new_G3475_ & new_G3476_;
  assign new_G3467_ = new_G3468_ | new_G3477_;
  assign new_G3468_ = G3457 | new_G3480_;
  assign new_G3469_ = new_G3479_ | new_G3478_;
  assign new_G3470_ = new_G3484_ & new_G3483_;
  assign new_G3471_ = new_G3482_ & new_G3481_;
  assign new_G3472_ = new_G3487_ | new_G3486_;
  assign new_G3473_ = new_G3482_ & new_G3485_;
  assign new_G3474_ = G3457 | new_G3490_;
  assign new_G3475_ = new_G3489_ | new_G3488_;
  assign new_G3476_ = new_G3492_ | new_G3491_;
  assign new_G3477_ = ~new_G3468_ & new_G3494_;
  assign new_G3478_ = ~new_G3470_ & new_G3482_;
  assign new_G3479_ = new_G3470_ & ~new_G3482_;
  assign new_G3480_ = G3456 & ~G3457;
  assign new_G3481_ = ~new_G3503_ | ~new_G3504_;
  assign new_G3482_ = new_G3496_ | new_G3498_;
  assign new_G3483_ = new_G3506_ | new_G3505_;
  assign new_G3484_ = new_G3500_ | new_G3499_;
  assign new_G3485_ = ~new_G3508_ | ~new_G3507_;
  assign new_G3486_ = ~new_G3509_ & new_G3510_;
  assign new_G3487_ = new_G3509_ & ~new_G3510_;
  assign new_G3488_ = ~G3456 & G3457;
  assign new_G3489_ = G3456 & ~G3457;
  assign new_G3490_ = ~new_G3472_ | new_G3482_;
  assign new_G3491_ = new_G3472_ & new_G3482_;
  assign new_G3492_ = ~new_G3472_ & ~new_G3482_;
  assign new_G3493_ = new_G3514_ | new_G3513_;
  assign new_G3494_ = G3460 | new_G3493_;
  assign new_G3495_ = new_G3518_ | new_G3517_;
  assign new_G3496_ = ~G3460 & new_G3495_;
  assign new_G3497_ = new_G3516_ | new_G3515_;
  assign new_G3498_ = G3460 & new_G3497_;
  assign new_G3499_ = G3458 & ~new_G3468_;
  assign new_G3500_ = ~G3458 & new_G3468_;
  assign new_G3501_ = ~G3457 | ~new_G3482_;
  assign new_G3502_ = new_G3468_ & new_G3501_;
  assign new_G3503_ = ~new_G3468_ & ~new_G3502_;
  assign new_G3504_ = new_G3468_ | new_G3501_;
  assign new_G3505_ = ~G3458 & G3459;
  assign new_G3506_ = G3458 & ~G3459;
  assign new_G3507_ = new_G3475_ | new_G3512_;
  assign new_G3508_ = ~new_G3475_ & ~new_G3511_;
  assign new_G3509_ = G3458 | new_G3475_;
  assign new_G3510_ = G3458 | G3459;
  assign new_G3511_ = new_G3475_ & new_G3512_;
  assign new_G3512_ = ~G3457 | ~new_G3482_;
  assign new_G3513_ = new_G3490_ & new_G3510_;
  assign new_G3514_ = ~new_G3490_ & ~new_G3510_;
  assign new_G3515_ = new_G3519_ | new_G3520_;
  assign new_G3516_ = ~G3461 & new_G3475_;
  assign new_G3517_ = new_G3521_ | new_G3522_;
  assign new_G3518_ = G3461 & new_G3475_;
  assign new_G3519_ = ~G3461 & ~new_G3475_;
  assign new_G3520_ = G3461 & ~new_G3475_;
  assign new_G3521_ = G3461 & ~new_G3475_;
  assign new_G3522_ = ~G3461 & new_G3475_;
  assign new_G3529_ = new_G3536_ & new_G3535_;
  assign new_G3530_ = new_G3538_ | new_G3537_;
  assign new_G3531_ = new_G3540_ | new_G3539_;
  assign new_G3532_ = new_G3542_ & new_G3541_;
  assign new_G3533_ = new_G3542_ & new_G3543_;
  assign new_G3534_ = new_G3535_ | new_G3544_;
  assign new_G3535_ = G3524 | new_G3547_;
  assign new_G3536_ = new_G3546_ | new_G3545_;
  assign new_G3537_ = new_G3551_ & new_G3550_;
  assign new_G3538_ = new_G3549_ & new_G3548_;
  assign new_G3539_ = new_G3554_ | new_G3553_;
  assign new_G3540_ = new_G3549_ & new_G3552_;
  assign new_G3541_ = G3524 | new_G3557_;
  assign new_G3542_ = new_G3556_ | new_G3555_;
  assign new_G3543_ = new_G3559_ | new_G3558_;
  assign new_G3544_ = ~new_G3535_ & new_G3561_;
  assign new_G3545_ = ~new_G3537_ & new_G3549_;
  assign new_G3546_ = new_G3537_ & ~new_G3549_;
  assign new_G3547_ = G3523 & ~G3524;
  assign new_G3548_ = ~new_G3570_ | ~new_G3571_;
  assign new_G3549_ = new_G3563_ | new_G3565_;
  assign new_G3550_ = new_G3573_ | new_G3572_;
  assign new_G3551_ = new_G3567_ | new_G3566_;
  assign new_G3552_ = ~new_G3575_ | ~new_G3574_;
  assign new_G3553_ = ~new_G3576_ & new_G3577_;
  assign new_G3554_ = new_G3576_ & ~new_G3577_;
  assign new_G3555_ = ~G3523 & G3524;
  assign new_G3556_ = G3523 & ~G3524;
  assign new_G3557_ = ~new_G3539_ | new_G3549_;
  assign new_G3558_ = new_G3539_ & new_G3549_;
  assign new_G3559_ = ~new_G3539_ & ~new_G3549_;
  assign new_G3560_ = new_G3581_ | new_G3580_;
  assign new_G3561_ = G3527 | new_G3560_;
  assign new_G3562_ = new_G3585_ | new_G3584_;
  assign new_G3563_ = ~G3527 & new_G3562_;
  assign new_G3564_ = new_G3583_ | new_G3582_;
  assign new_G3565_ = G3527 & new_G3564_;
  assign new_G3566_ = G3525 & ~new_G3535_;
  assign new_G3567_ = ~G3525 & new_G3535_;
  assign new_G3568_ = ~G3524 | ~new_G3549_;
  assign new_G3569_ = new_G3535_ & new_G3568_;
  assign new_G3570_ = ~new_G3535_ & ~new_G3569_;
  assign new_G3571_ = new_G3535_ | new_G3568_;
  assign new_G3572_ = ~G3525 & G3526;
  assign new_G3573_ = G3525 & ~G3526;
  assign new_G3574_ = new_G3542_ | new_G3579_;
  assign new_G3575_ = ~new_G3542_ & ~new_G3578_;
  assign new_G3576_ = G3525 | new_G3542_;
  assign new_G3577_ = G3525 | G3526;
  assign new_G3578_ = new_G3542_ & new_G3579_;
  assign new_G3579_ = ~G3524 | ~new_G3549_;
  assign new_G3580_ = new_G3557_ & new_G3577_;
  assign new_G3581_ = ~new_G3557_ & ~new_G3577_;
  assign new_G3582_ = new_G3586_ | new_G3587_;
  assign new_G3583_ = ~G3528 & new_G3542_;
  assign new_G3584_ = new_G3588_ | new_G3589_;
  assign new_G3585_ = G3528 & new_G3542_;
  assign new_G3586_ = ~G3528 & ~new_G3542_;
  assign new_G3587_ = G3528 & ~new_G3542_;
  assign new_G3588_ = G3528 & ~new_G3542_;
  assign new_G3589_ = ~G3528 & new_G3542_;
  assign new_G3596_ = new_G3603_ & new_G3602_;
  assign new_G3597_ = new_G3605_ | new_G3604_;
  assign new_G3598_ = new_G3607_ | new_G3606_;
  assign new_G3599_ = new_G3609_ & new_G3608_;
  assign new_G3600_ = new_G3609_ & new_G3610_;
  assign new_G3601_ = new_G3602_ | new_G3611_;
  assign new_G3602_ = G3591 | new_G3614_;
  assign new_G3603_ = new_G3613_ | new_G3612_;
  assign new_G3604_ = new_G3618_ & new_G3617_;
  assign new_G3605_ = new_G3616_ & new_G3615_;
  assign new_G3606_ = new_G3621_ | new_G3620_;
  assign new_G3607_ = new_G3616_ & new_G3619_;
  assign new_G3608_ = G3591 | new_G3624_;
  assign new_G3609_ = new_G3623_ | new_G3622_;
  assign new_G3610_ = new_G3626_ | new_G3625_;
  assign new_G3611_ = ~new_G3602_ & new_G3628_;
  assign new_G3612_ = ~new_G3604_ & new_G3616_;
  assign new_G3613_ = new_G3604_ & ~new_G3616_;
  assign new_G3614_ = G3590 & ~G3591;
  assign new_G3615_ = ~new_G3637_ | ~new_G3638_;
  assign new_G3616_ = new_G3630_ | new_G3632_;
  assign new_G3617_ = new_G3640_ | new_G3639_;
  assign new_G3618_ = new_G3634_ | new_G3633_;
  assign new_G3619_ = ~new_G3642_ | ~new_G3641_;
  assign new_G3620_ = ~new_G3643_ & new_G3644_;
  assign new_G3621_ = new_G3643_ & ~new_G3644_;
  assign new_G3622_ = ~G3590 & G3591;
  assign new_G3623_ = G3590 & ~G3591;
  assign new_G3624_ = ~new_G3606_ | new_G3616_;
  assign new_G3625_ = new_G3606_ & new_G3616_;
  assign new_G3626_ = ~new_G3606_ & ~new_G3616_;
  assign new_G3627_ = new_G3648_ | new_G3647_;
  assign new_G3628_ = G3594 | new_G3627_;
  assign new_G3629_ = new_G3652_ | new_G3651_;
  assign new_G3630_ = ~G3594 & new_G3629_;
  assign new_G3631_ = new_G3650_ | new_G3649_;
  assign new_G3632_ = G3594 & new_G3631_;
  assign new_G3633_ = G3592 & ~new_G3602_;
  assign new_G3634_ = ~G3592 & new_G3602_;
  assign new_G3635_ = ~G3591 | ~new_G3616_;
  assign new_G3636_ = new_G3602_ & new_G3635_;
  assign new_G3637_ = ~new_G3602_ & ~new_G3636_;
  assign new_G3638_ = new_G3602_ | new_G3635_;
  assign new_G3639_ = ~G3592 & G3593;
  assign new_G3640_ = G3592 & ~G3593;
  assign new_G3641_ = new_G3609_ | new_G3646_;
  assign new_G3642_ = ~new_G3609_ & ~new_G3645_;
  assign new_G3643_ = G3592 | new_G3609_;
  assign new_G3644_ = G3592 | G3593;
  assign new_G3645_ = new_G3609_ & new_G3646_;
  assign new_G3646_ = ~G3591 | ~new_G3616_;
  assign new_G3647_ = new_G3624_ & new_G3644_;
  assign new_G3648_ = ~new_G3624_ & ~new_G3644_;
  assign new_G3649_ = new_G3653_ | new_G3654_;
  assign new_G3650_ = ~G3595 & new_G3609_;
  assign new_G3651_ = new_G3655_ | new_G3656_;
  assign new_G3652_ = G3595 & new_G3609_;
  assign new_G3653_ = ~G3595 & ~new_G3609_;
  assign new_G3654_ = G3595 & ~new_G3609_;
  assign new_G3655_ = G3595 & ~new_G3609_;
  assign new_G3656_ = ~G3595 & new_G3609_;
  assign new_G3663_ = new_G3670_ & new_G3669_;
  assign new_G3664_ = new_G3672_ | new_G3671_;
  assign new_G3665_ = new_G3674_ | new_G3673_;
  assign new_G3666_ = new_G3676_ & new_G3675_;
  assign new_G3667_ = new_G3676_ & new_G3677_;
  assign new_G3668_ = new_G3669_ | new_G3678_;
  assign new_G3669_ = G3658 | new_G3681_;
  assign new_G3670_ = new_G3680_ | new_G3679_;
  assign new_G3671_ = new_G3685_ & new_G3684_;
  assign new_G3672_ = new_G3683_ & new_G3682_;
  assign new_G3673_ = new_G3688_ | new_G3687_;
  assign new_G3674_ = new_G3683_ & new_G3686_;
  assign new_G3675_ = G3658 | new_G3691_;
  assign new_G3676_ = new_G3690_ | new_G3689_;
  assign new_G3677_ = new_G3693_ | new_G3692_;
  assign new_G3678_ = ~new_G3669_ & new_G3695_;
  assign new_G3679_ = ~new_G3671_ & new_G3683_;
  assign new_G3680_ = new_G3671_ & ~new_G3683_;
  assign new_G3681_ = G3657 & ~G3658;
  assign new_G3682_ = ~new_G3704_ | ~new_G3705_;
  assign new_G3683_ = new_G3697_ | new_G3699_;
  assign new_G3684_ = new_G3707_ | new_G3706_;
  assign new_G3685_ = new_G3701_ | new_G3700_;
  assign new_G3686_ = ~new_G3709_ | ~new_G3708_;
  assign new_G3687_ = ~new_G3710_ & new_G3711_;
  assign new_G3688_ = new_G3710_ & ~new_G3711_;
  assign new_G3689_ = ~G3657 & G3658;
  assign new_G3690_ = G3657 & ~G3658;
  assign new_G3691_ = ~new_G3673_ | new_G3683_;
  assign new_G3692_ = new_G3673_ & new_G3683_;
  assign new_G3693_ = ~new_G3673_ & ~new_G3683_;
  assign new_G3694_ = new_G3715_ | new_G3714_;
  assign new_G3695_ = G3661 | new_G3694_;
  assign new_G3696_ = new_G3719_ | new_G3718_;
  assign new_G3697_ = ~G3661 & new_G3696_;
  assign new_G3698_ = new_G3717_ | new_G3716_;
  assign new_G3699_ = G3661 & new_G3698_;
  assign new_G3700_ = G3659 & ~new_G3669_;
  assign new_G3701_ = ~G3659 & new_G3669_;
  assign new_G3702_ = ~G3658 | ~new_G3683_;
  assign new_G3703_ = new_G3669_ & new_G3702_;
  assign new_G3704_ = ~new_G3669_ & ~new_G3703_;
  assign new_G3705_ = new_G3669_ | new_G3702_;
  assign new_G3706_ = ~G3659 & G3660;
  assign new_G3707_ = G3659 & ~G3660;
  assign new_G3708_ = new_G3676_ | new_G3713_;
  assign new_G3709_ = ~new_G3676_ & ~new_G3712_;
  assign new_G3710_ = G3659 | new_G3676_;
  assign new_G3711_ = G3659 | G3660;
  assign new_G3712_ = new_G3676_ & new_G3713_;
  assign new_G3713_ = ~G3658 | ~new_G3683_;
  assign new_G3714_ = new_G3691_ & new_G3711_;
  assign new_G3715_ = ~new_G3691_ & ~new_G3711_;
  assign new_G3716_ = new_G3720_ | new_G3721_;
  assign new_G3717_ = ~G3662 & new_G3676_;
  assign new_G3718_ = new_G3722_ | new_G3723_;
  assign new_G3719_ = G3662 & new_G3676_;
  assign new_G3720_ = ~G3662 & ~new_G3676_;
  assign new_G3721_ = G3662 & ~new_G3676_;
  assign new_G3722_ = G3662 & ~new_G3676_;
  assign new_G3723_ = ~G3662 & new_G3676_;
  assign new_G3730_ = new_G3737_ & new_G3736_;
  assign new_G3731_ = new_G3739_ | new_G3738_;
  assign new_G3732_ = new_G3741_ | new_G3740_;
  assign new_G3733_ = new_G3743_ & new_G3742_;
  assign new_G3734_ = new_G3743_ & new_G3744_;
  assign new_G3735_ = new_G3736_ | new_G3745_;
  assign new_G3736_ = G3725 | new_G3748_;
  assign new_G3737_ = new_G3747_ | new_G3746_;
  assign new_G3738_ = new_G3752_ & new_G3751_;
  assign new_G3739_ = new_G3750_ & new_G3749_;
  assign new_G3740_ = new_G3755_ | new_G3754_;
  assign new_G3741_ = new_G3750_ & new_G3753_;
  assign new_G3742_ = G3725 | new_G3758_;
  assign new_G3743_ = new_G3757_ | new_G3756_;
  assign new_G3744_ = new_G3760_ | new_G3759_;
  assign new_G3745_ = ~new_G3736_ & new_G3762_;
  assign new_G3746_ = ~new_G3738_ & new_G3750_;
  assign new_G3747_ = new_G3738_ & ~new_G3750_;
  assign new_G3748_ = G3724 & ~G3725;
  assign new_G3749_ = ~new_G3771_ | ~new_G3772_;
  assign new_G3750_ = new_G3764_ | new_G3766_;
  assign new_G3751_ = new_G3774_ | new_G3773_;
  assign new_G3752_ = new_G3768_ | new_G3767_;
  assign new_G3753_ = ~new_G3776_ | ~new_G3775_;
  assign new_G3754_ = ~new_G3777_ & new_G3778_;
  assign new_G3755_ = new_G3777_ & ~new_G3778_;
  assign new_G3756_ = ~G3724 & G3725;
  assign new_G3757_ = G3724 & ~G3725;
  assign new_G3758_ = ~new_G3740_ | new_G3750_;
  assign new_G3759_ = new_G3740_ & new_G3750_;
  assign new_G3760_ = ~new_G3740_ & ~new_G3750_;
  assign new_G3761_ = new_G3782_ | new_G3781_;
  assign new_G3762_ = G3728 | new_G3761_;
  assign new_G3763_ = new_G3786_ | new_G3785_;
  assign new_G3764_ = ~G3728 & new_G3763_;
  assign new_G3765_ = new_G3784_ | new_G3783_;
  assign new_G3766_ = G3728 & new_G3765_;
  assign new_G3767_ = G3726 & ~new_G3736_;
  assign new_G3768_ = ~G3726 & new_G3736_;
  assign new_G3769_ = ~G3725 | ~new_G3750_;
  assign new_G3770_ = new_G3736_ & new_G3769_;
  assign new_G3771_ = ~new_G3736_ & ~new_G3770_;
  assign new_G3772_ = new_G3736_ | new_G3769_;
  assign new_G3773_ = ~G3726 & G3727;
  assign new_G3774_ = G3726 & ~G3727;
  assign new_G3775_ = new_G3743_ | new_G3780_;
  assign new_G3776_ = ~new_G3743_ & ~new_G3779_;
  assign new_G3777_ = G3726 | new_G3743_;
  assign new_G3778_ = G3726 | G3727;
  assign new_G3779_ = new_G3743_ & new_G3780_;
  assign new_G3780_ = ~G3725 | ~new_G3750_;
  assign new_G3781_ = new_G3758_ & new_G3778_;
  assign new_G3782_ = ~new_G3758_ & ~new_G3778_;
  assign new_G3783_ = new_G3787_ | new_G3788_;
  assign new_G3784_ = ~G3729 & new_G3743_;
  assign new_G3785_ = new_G3789_ | new_G3790_;
  assign new_G3786_ = G3729 & new_G3743_;
  assign new_G3787_ = ~G3729 & ~new_G3743_;
  assign new_G3788_ = G3729 & ~new_G3743_;
  assign new_G3789_ = G3729 & ~new_G3743_;
  assign new_G3790_ = ~G3729 & new_G3743_;
  assign new_G3797_ = new_G3804_ & new_G3803_;
  assign new_G3798_ = new_G3806_ | new_G3805_;
  assign new_G3799_ = new_G3808_ | new_G3807_;
  assign new_G3800_ = new_G3810_ & new_G3809_;
  assign new_G3801_ = new_G3810_ & new_G3811_;
  assign new_G3802_ = new_G3803_ | new_G3812_;
  assign new_G3803_ = G3792 | new_G3815_;
  assign new_G3804_ = new_G3814_ | new_G3813_;
  assign new_G3805_ = new_G3819_ & new_G3818_;
  assign new_G3806_ = new_G3817_ & new_G3816_;
  assign new_G3807_ = new_G3822_ | new_G3821_;
  assign new_G3808_ = new_G3817_ & new_G3820_;
  assign new_G3809_ = G3792 | new_G3825_;
  assign new_G3810_ = new_G3824_ | new_G3823_;
  assign new_G3811_ = new_G3827_ | new_G3826_;
  assign new_G3812_ = ~new_G3803_ & new_G3829_;
  assign new_G3813_ = ~new_G3805_ & new_G3817_;
  assign new_G3814_ = new_G3805_ & ~new_G3817_;
  assign new_G3815_ = G3791 & ~G3792;
  assign new_G3816_ = ~new_G3838_ | ~new_G3839_;
  assign new_G3817_ = new_G3831_ | new_G3833_;
  assign new_G3818_ = new_G3841_ | new_G3840_;
  assign new_G3819_ = new_G3835_ | new_G3834_;
  assign new_G3820_ = ~new_G3843_ | ~new_G3842_;
  assign new_G3821_ = ~new_G3844_ & new_G3845_;
  assign new_G3822_ = new_G3844_ & ~new_G3845_;
  assign new_G3823_ = ~G3791 & G3792;
  assign new_G3824_ = G3791 & ~G3792;
  assign new_G3825_ = ~new_G3807_ | new_G3817_;
  assign new_G3826_ = new_G3807_ & new_G3817_;
  assign new_G3827_ = ~new_G3807_ & ~new_G3817_;
  assign new_G3828_ = new_G3849_ | new_G3848_;
  assign new_G3829_ = G3795 | new_G3828_;
  assign new_G3830_ = new_G3853_ | new_G3852_;
  assign new_G3831_ = ~G3795 & new_G3830_;
  assign new_G3832_ = new_G3851_ | new_G3850_;
  assign new_G3833_ = G3795 & new_G3832_;
  assign new_G3834_ = G3793 & ~new_G3803_;
  assign new_G3835_ = ~G3793 & new_G3803_;
  assign new_G3836_ = ~G3792 | ~new_G3817_;
  assign new_G3837_ = new_G3803_ & new_G3836_;
  assign new_G3838_ = ~new_G3803_ & ~new_G3837_;
  assign new_G3839_ = new_G3803_ | new_G3836_;
  assign new_G3840_ = ~G3793 & G3794;
  assign new_G3841_ = G3793 & ~G3794;
  assign new_G3842_ = new_G3810_ | new_G3847_;
  assign new_G3843_ = ~new_G3810_ & ~new_G3846_;
  assign new_G3844_ = G3793 | new_G3810_;
  assign new_G3845_ = G3793 | G3794;
  assign new_G3846_ = new_G3810_ & new_G3847_;
  assign new_G3847_ = ~G3792 | ~new_G3817_;
  assign new_G3848_ = new_G3825_ & new_G3845_;
  assign new_G3849_ = ~new_G3825_ & ~new_G3845_;
  assign new_G3850_ = new_G3854_ | new_G3855_;
  assign new_G3851_ = ~G3796 & new_G3810_;
  assign new_G3852_ = new_G3856_ | new_G3857_;
  assign new_G3853_ = G3796 & new_G3810_;
  assign new_G3854_ = ~G3796 & ~new_G3810_;
  assign new_G3855_ = G3796 & ~new_G3810_;
  assign new_G3856_ = G3796 & ~new_G3810_;
  assign new_G3857_ = ~G3796 & new_G3810_;
  assign new_G3864_ = new_G3871_ & new_G3870_;
  assign new_G3865_ = new_G3873_ | new_G3872_;
  assign new_G3866_ = new_G3875_ | new_G3874_;
  assign new_G3867_ = new_G3877_ & new_G3876_;
  assign new_G3868_ = new_G3877_ & new_G3878_;
  assign new_G3869_ = new_G3870_ | new_G3879_;
  assign new_G3870_ = G3859 | new_G3882_;
  assign new_G3871_ = new_G3881_ | new_G3880_;
  assign new_G3872_ = new_G3886_ & new_G3885_;
  assign new_G3873_ = new_G3884_ & new_G3883_;
  assign new_G3874_ = new_G3889_ | new_G3888_;
  assign new_G3875_ = new_G3884_ & new_G3887_;
  assign new_G3876_ = G3859 | new_G3892_;
  assign new_G3877_ = new_G3891_ | new_G3890_;
  assign new_G3878_ = new_G3894_ | new_G3893_;
  assign new_G3879_ = ~new_G3870_ & new_G3896_;
  assign new_G3880_ = ~new_G3872_ & new_G3884_;
  assign new_G3881_ = new_G3872_ & ~new_G3884_;
  assign new_G3882_ = G3858 & ~G3859;
  assign new_G3883_ = ~new_G3905_ | ~new_G3906_;
  assign new_G3884_ = new_G3898_ | new_G3900_;
  assign new_G3885_ = new_G3908_ | new_G3907_;
  assign new_G3886_ = new_G3902_ | new_G3901_;
  assign new_G3887_ = ~new_G3910_ | ~new_G3909_;
  assign new_G3888_ = ~new_G3911_ & new_G3912_;
  assign new_G3889_ = new_G3911_ & ~new_G3912_;
  assign new_G3890_ = ~G3858 & G3859;
  assign new_G3891_ = G3858 & ~G3859;
  assign new_G3892_ = ~new_G3874_ | new_G3884_;
  assign new_G3893_ = new_G3874_ & new_G3884_;
  assign new_G3894_ = ~new_G3874_ & ~new_G3884_;
  assign new_G3895_ = new_G3916_ | new_G3915_;
  assign new_G3896_ = G3862 | new_G3895_;
  assign new_G3897_ = new_G3920_ | new_G3919_;
  assign new_G3898_ = ~G3862 & new_G3897_;
  assign new_G3899_ = new_G3918_ | new_G3917_;
  assign new_G3900_ = G3862 & new_G3899_;
  assign new_G3901_ = G3860 & ~new_G3870_;
  assign new_G3902_ = ~G3860 & new_G3870_;
  assign new_G3903_ = ~G3859 | ~new_G3884_;
  assign new_G3904_ = new_G3870_ & new_G3903_;
  assign new_G3905_ = ~new_G3870_ & ~new_G3904_;
  assign new_G3906_ = new_G3870_ | new_G3903_;
  assign new_G3907_ = ~G3860 & G3861;
  assign new_G3908_ = G3860 & ~G3861;
  assign new_G3909_ = new_G3877_ | new_G3914_;
  assign new_G3910_ = ~new_G3877_ & ~new_G3913_;
  assign new_G3911_ = G3860 | new_G3877_;
  assign new_G3912_ = G3860 | G3861;
  assign new_G3913_ = new_G3877_ & new_G3914_;
  assign new_G3914_ = ~G3859 | ~new_G3884_;
  assign new_G3915_ = new_G3892_ & new_G3912_;
  assign new_G3916_ = ~new_G3892_ & ~new_G3912_;
  assign new_G3917_ = new_G3921_ | new_G3922_;
  assign new_G3918_ = ~G3863 & new_G3877_;
  assign new_G3919_ = new_G3923_ | new_G3924_;
  assign new_G3920_ = G3863 & new_G3877_;
  assign new_G3921_ = ~G3863 & ~new_G3877_;
  assign new_G3922_ = G3863 & ~new_G3877_;
  assign new_G3923_ = G3863 & ~new_G3877_;
  assign new_G3924_ = ~G3863 & new_G3877_;
  assign new_G3931_ = new_G3938_ & new_G3937_;
  assign new_G3932_ = new_G3940_ | new_G3939_;
  assign new_G3933_ = new_G3942_ | new_G3941_;
  assign new_G3934_ = new_G3944_ & new_G3943_;
  assign new_G3935_ = new_G3944_ & new_G3945_;
  assign new_G3936_ = new_G3937_ | new_G3946_;
  assign new_G3937_ = G3926 | new_G3949_;
  assign new_G3938_ = new_G3948_ | new_G3947_;
  assign new_G3939_ = new_G3953_ & new_G3952_;
  assign new_G3940_ = new_G3951_ & new_G3950_;
  assign new_G3941_ = new_G3956_ | new_G3955_;
  assign new_G3942_ = new_G3951_ & new_G3954_;
  assign new_G3943_ = G3926 | new_G3959_;
  assign new_G3944_ = new_G3958_ | new_G3957_;
  assign new_G3945_ = new_G3961_ | new_G3960_;
  assign new_G3946_ = ~new_G3937_ & new_G3963_;
  assign new_G3947_ = ~new_G3939_ & new_G3951_;
  assign new_G3948_ = new_G3939_ & ~new_G3951_;
  assign new_G3949_ = G3925 & ~G3926;
  assign new_G3950_ = ~new_G3972_ | ~new_G3973_;
  assign new_G3951_ = new_G3965_ | new_G3967_;
  assign new_G3952_ = new_G3975_ | new_G3974_;
  assign new_G3953_ = new_G3969_ | new_G3968_;
  assign new_G3954_ = ~new_G3977_ | ~new_G3976_;
  assign new_G3955_ = ~new_G3978_ & new_G3979_;
  assign new_G3956_ = new_G3978_ & ~new_G3979_;
  assign new_G3957_ = ~G3925 & G3926;
  assign new_G3958_ = G3925 & ~G3926;
  assign new_G3959_ = ~new_G3941_ | new_G3951_;
  assign new_G3960_ = new_G3941_ & new_G3951_;
  assign new_G3961_ = ~new_G3941_ & ~new_G3951_;
  assign new_G3962_ = new_G3983_ | new_G3982_;
  assign new_G3963_ = G3929 | new_G3962_;
  assign new_G3964_ = new_G3987_ | new_G3986_;
  assign new_G3965_ = ~G3929 & new_G3964_;
  assign new_G3966_ = new_G3985_ | new_G3984_;
  assign new_G3967_ = G3929 & new_G3966_;
  assign new_G3968_ = G3927 & ~new_G3937_;
  assign new_G3969_ = ~G3927 & new_G3937_;
  assign new_G3970_ = ~G3926 | ~new_G3951_;
  assign new_G3971_ = new_G3937_ & new_G3970_;
  assign new_G3972_ = ~new_G3937_ & ~new_G3971_;
  assign new_G3973_ = new_G3937_ | new_G3970_;
  assign new_G3974_ = ~G3927 & G3928;
  assign new_G3975_ = G3927 & ~G3928;
  assign new_G3976_ = new_G3944_ | new_G3981_;
  assign new_G3977_ = ~new_G3944_ & ~new_G3980_;
  assign new_G3978_ = G3927 | new_G3944_;
  assign new_G3979_ = G3927 | G3928;
  assign new_G3980_ = new_G3944_ & new_G3981_;
  assign new_G3981_ = ~G3926 | ~new_G3951_;
  assign new_G3982_ = new_G3959_ & new_G3979_;
  assign new_G3983_ = ~new_G3959_ & ~new_G3979_;
  assign new_G3984_ = new_G3988_ | new_G3989_;
  assign new_G3985_ = ~G3930 & new_G3944_;
  assign new_G3986_ = new_G3990_ | new_G3991_;
  assign new_G3987_ = G3930 & new_G3944_;
  assign new_G3988_ = ~G3930 & ~new_G3944_;
  assign new_G3989_ = G3930 & ~new_G3944_;
  assign new_G3990_ = G3930 & ~new_G3944_;
  assign new_G3991_ = ~G3930 & new_G3944_;
  assign new_G3998_ = new_G4005_ & new_G4004_;
  assign new_G3999_ = new_G4007_ | new_G4006_;
  assign new_G4000_ = new_G4009_ | new_G4008_;
  assign new_G4001_ = new_G4011_ & new_G4010_;
  assign new_G4002_ = new_G4011_ & new_G4012_;
  assign new_G4003_ = new_G4004_ | new_G4013_;
  assign new_G4004_ = G3993 | new_G4016_;
  assign new_G4005_ = new_G4015_ | new_G4014_;
  assign new_G4006_ = new_G4020_ & new_G4019_;
  assign new_G4007_ = new_G4018_ & new_G4017_;
  assign new_G4008_ = new_G4023_ | new_G4022_;
  assign new_G4009_ = new_G4018_ & new_G4021_;
  assign new_G4010_ = G3993 | new_G4026_;
  assign new_G4011_ = new_G4025_ | new_G4024_;
  assign new_G4012_ = new_G4028_ | new_G4027_;
  assign new_G4013_ = ~new_G4004_ & new_G4030_;
  assign new_G4014_ = ~new_G4006_ & new_G4018_;
  assign new_G4015_ = new_G4006_ & ~new_G4018_;
  assign new_G4016_ = G3992 & ~G3993;
  assign new_G4017_ = ~new_G4039_ | ~new_G4040_;
  assign new_G4018_ = new_G4032_ | new_G4034_;
  assign new_G4019_ = new_G4042_ | new_G4041_;
  assign new_G4020_ = new_G4036_ | new_G4035_;
  assign new_G4021_ = ~new_G4044_ | ~new_G4043_;
  assign new_G4022_ = ~new_G4045_ & new_G4046_;
  assign new_G4023_ = new_G4045_ & ~new_G4046_;
  assign new_G4024_ = ~G3992 & G3993;
  assign new_G4025_ = G3992 & ~G3993;
  assign new_G4026_ = ~new_G4008_ | new_G4018_;
  assign new_G4027_ = new_G4008_ & new_G4018_;
  assign new_G4028_ = ~new_G4008_ & ~new_G4018_;
  assign new_G4029_ = new_G4050_ | new_G4049_;
  assign new_G4030_ = G3996 | new_G4029_;
  assign new_G4031_ = new_G4054_ | new_G4053_;
  assign new_G4032_ = ~G3996 & new_G4031_;
  assign new_G4033_ = new_G4052_ | new_G4051_;
  assign new_G4034_ = G3996 & new_G4033_;
  assign new_G4035_ = G3994 & ~new_G4004_;
  assign new_G4036_ = ~G3994 & new_G4004_;
  assign new_G4037_ = ~G3993 | ~new_G4018_;
  assign new_G4038_ = new_G4004_ & new_G4037_;
  assign new_G4039_ = ~new_G4004_ & ~new_G4038_;
  assign new_G4040_ = new_G4004_ | new_G4037_;
  assign new_G4041_ = ~G3994 & G3995;
  assign new_G4042_ = G3994 & ~G3995;
  assign new_G4043_ = new_G4011_ | new_G4048_;
  assign new_G4044_ = ~new_G4011_ & ~new_G4047_;
  assign new_G4045_ = G3994 | new_G4011_;
  assign new_G4046_ = G3994 | G3995;
  assign new_G4047_ = new_G4011_ & new_G4048_;
  assign new_G4048_ = ~G3993 | ~new_G4018_;
  assign new_G4049_ = new_G4026_ & new_G4046_;
  assign new_G4050_ = ~new_G4026_ & ~new_G4046_;
  assign new_G4051_ = new_G4055_ | new_G4056_;
  assign new_G4052_ = ~G3997 & new_G4011_;
  assign new_G4053_ = new_G4057_ | new_G4058_;
  assign new_G4054_ = G3997 & new_G4011_;
  assign new_G4055_ = ~G3997 & ~new_G4011_;
  assign new_G4056_ = G3997 & ~new_G4011_;
  assign new_G4057_ = G3997 & ~new_G4011_;
  assign new_G4058_ = ~G3997 & new_G4011_;
  assign new_G4065_ = new_G4072_ & new_G4071_;
  assign new_G4066_ = new_G4074_ | new_G4073_;
  assign new_G4067_ = new_G4076_ | new_G4075_;
  assign new_G4068_ = new_G4078_ & new_G4077_;
  assign new_G4069_ = new_G4078_ & new_G4079_;
  assign new_G4070_ = new_G4071_ | new_G4080_;
  assign new_G4071_ = G4060 | new_G4083_;
  assign new_G4072_ = new_G4082_ | new_G4081_;
  assign new_G4073_ = new_G4087_ & new_G4086_;
  assign new_G4074_ = new_G4085_ & new_G4084_;
  assign new_G4075_ = new_G4090_ | new_G4089_;
  assign new_G4076_ = new_G4085_ & new_G4088_;
  assign new_G4077_ = G4060 | new_G4093_;
  assign new_G4078_ = new_G4092_ | new_G4091_;
  assign new_G4079_ = new_G4095_ | new_G4094_;
  assign new_G4080_ = ~new_G4071_ & new_G4097_;
  assign new_G4081_ = ~new_G4073_ & new_G4085_;
  assign new_G4082_ = new_G4073_ & ~new_G4085_;
  assign new_G4083_ = G4059 & ~G4060;
  assign new_G4084_ = ~new_G4106_ | ~new_G4107_;
  assign new_G4085_ = new_G4099_ | new_G4101_;
  assign new_G4086_ = new_G4109_ | new_G4108_;
  assign new_G4087_ = new_G4103_ | new_G4102_;
  assign new_G4088_ = ~new_G4111_ | ~new_G4110_;
  assign new_G4089_ = ~new_G4112_ & new_G4113_;
  assign new_G4090_ = new_G4112_ & ~new_G4113_;
  assign new_G4091_ = ~G4059 & G4060;
  assign new_G4092_ = G4059 & ~G4060;
  assign new_G4093_ = ~new_G4075_ | new_G4085_;
  assign new_G4094_ = new_G4075_ & new_G4085_;
  assign new_G4095_ = ~new_G4075_ & ~new_G4085_;
  assign new_G4096_ = new_G4117_ | new_G4116_;
  assign new_G4097_ = G4063 | new_G4096_;
  assign new_G4098_ = new_G4121_ | new_G4120_;
  assign new_G4099_ = ~G4063 & new_G4098_;
  assign new_G4100_ = new_G4119_ | new_G4118_;
  assign new_G4101_ = G4063 & new_G4100_;
  assign new_G4102_ = G4061 & ~new_G4071_;
  assign new_G4103_ = ~G4061 & new_G4071_;
  assign new_G4104_ = ~G4060 | ~new_G4085_;
  assign new_G4105_ = new_G4071_ & new_G4104_;
  assign new_G4106_ = ~new_G4071_ & ~new_G4105_;
  assign new_G4107_ = new_G4071_ | new_G4104_;
  assign new_G4108_ = ~G4061 & G4062;
  assign new_G4109_ = G4061 & ~G4062;
  assign new_G4110_ = new_G4078_ | new_G4115_;
  assign new_G4111_ = ~new_G4078_ & ~new_G4114_;
  assign new_G4112_ = G4061 | new_G4078_;
  assign new_G4113_ = G4061 | G4062;
  assign new_G4114_ = new_G4078_ & new_G4115_;
  assign new_G4115_ = ~G4060 | ~new_G4085_;
  assign new_G4116_ = new_G4093_ & new_G4113_;
  assign new_G4117_ = ~new_G4093_ & ~new_G4113_;
  assign new_G4118_ = new_G4122_ | new_G4123_;
  assign new_G4119_ = ~G4064 & new_G4078_;
  assign new_G4120_ = new_G4124_ | new_G4125_;
  assign new_G4121_ = G4064 & new_G4078_;
  assign new_G4122_ = ~G4064 & ~new_G4078_;
  assign new_G4123_ = G4064 & ~new_G4078_;
  assign new_G4124_ = G4064 & ~new_G4078_;
  assign new_G4125_ = ~G4064 & new_G4078_;
  assign new_G4132_ = new_G4139_ & new_G4138_;
  assign new_G4133_ = new_G4141_ | new_G4140_;
  assign new_G4134_ = new_G4143_ | new_G4142_;
  assign new_G4135_ = new_G4145_ & new_G4144_;
  assign new_G4136_ = new_G4145_ & new_G4146_;
  assign new_G4137_ = new_G4138_ | new_G4147_;
  assign new_G4138_ = G4127 | new_G4150_;
  assign new_G4139_ = new_G4149_ | new_G4148_;
  assign new_G4140_ = new_G4154_ & new_G4153_;
  assign new_G4141_ = new_G4152_ & new_G4151_;
  assign new_G4142_ = new_G4157_ | new_G4156_;
  assign new_G4143_ = new_G4152_ & new_G4155_;
  assign new_G4144_ = G4127 | new_G4160_;
  assign new_G4145_ = new_G4159_ | new_G4158_;
  assign new_G4146_ = new_G4162_ | new_G4161_;
  assign new_G4147_ = ~new_G4138_ & new_G4164_;
  assign new_G4148_ = ~new_G4140_ & new_G4152_;
  assign new_G4149_ = new_G4140_ & ~new_G4152_;
  assign new_G4150_ = G4126 & ~G4127;
  assign new_G4151_ = ~new_G4173_ | ~new_G4174_;
  assign new_G4152_ = new_G4166_ | new_G4168_;
  assign new_G4153_ = new_G4176_ | new_G4175_;
  assign new_G4154_ = new_G4170_ | new_G4169_;
  assign new_G4155_ = ~new_G4178_ | ~new_G4177_;
  assign new_G4156_ = ~new_G4179_ & new_G4180_;
  assign new_G4157_ = new_G4179_ & ~new_G4180_;
  assign new_G4158_ = ~G4126 & G4127;
  assign new_G4159_ = G4126 & ~G4127;
  assign new_G4160_ = ~new_G4142_ | new_G4152_;
  assign new_G4161_ = new_G4142_ & new_G4152_;
  assign new_G4162_ = ~new_G4142_ & ~new_G4152_;
  assign new_G4163_ = new_G4184_ | new_G4183_;
  assign new_G4164_ = G4130 | new_G4163_;
  assign new_G4165_ = new_G4188_ | new_G4187_;
  assign new_G4166_ = ~G4130 & new_G4165_;
  assign new_G4167_ = new_G4186_ | new_G4185_;
  assign new_G4168_ = G4130 & new_G4167_;
  assign new_G4169_ = G4128 & ~new_G4138_;
  assign new_G4170_ = ~G4128 & new_G4138_;
  assign new_G4171_ = ~G4127 | ~new_G4152_;
  assign new_G4172_ = new_G4138_ & new_G4171_;
  assign new_G4173_ = ~new_G4138_ & ~new_G4172_;
  assign new_G4174_ = new_G4138_ | new_G4171_;
  assign new_G4175_ = ~G4128 & G4129;
  assign new_G4176_ = G4128 & ~G4129;
  assign new_G4177_ = new_G4145_ | new_G4182_;
  assign new_G4178_ = ~new_G4145_ & ~new_G4181_;
  assign new_G4179_ = G4128 | new_G4145_;
  assign new_G4180_ = G4128 | G4129;
  assign new_G4181_ = new_G4145_ & new_G4182_;
  assign new_G4182_ = ~G4127 | ~new_G4152_;
  assign new_G4183_ = new_G4160_ & new_G4180_;
  assign new_G4184_ = ~new_G4160_ & ~new_G4180_;
  assign new_G4185_ = new_G4189_ | new_G4190_;
  assign new_G4186_ = ~G4131 & new_G4145_;
  assign new_G4187_ = new_G4191_ | new_G4192_;
  assign new_G4188_ = G4131 & new_G4145_;
  assign new_G4189_ = ~G4131 & ~new_G4145_;
  assign new_G4190_ = G4131 & ~new_G4145_;
  assign new_G4191_ = G4131 & ~new_G4145_;
  assign new_G4192_ = ~G4131 & new_G4145_;
  assign new_G4199_ = new_G4206_ & new_G4205_;
  assign new_G4200_ = new_G4208_ | new_G4207_;
  assign new_G4201_ = new_G4210_ | new_G4209_;
  assign new_G4202_ = new_G4212_ & new_G4211_;
  assign new_G4203_ = new_G4212_ & new_G4213_;
  assign new_G4204_ = new_G4205_ | new_G4214_;
  assign new_G4205_ = G4194 | new_G4217_;
  assign new_G4206_ = new_G4216_ | new_G4215_;
  assign new_G4207_ = new_G4221_ & new_G4220_;
  assign new_G4208_ = new_G4219_ & new_G4218_;
  assign new_G4209_ = new_G4224_ | new_G4223_;
  assign new_G4210_ = new_G4219_ & new_G4222_;
  assign new_G4211_ = G4194 | new_G4227_;
  assign new_G4212_ = new_G4226_ | new_G4225_;
  assign new_G4213_ = new_G4229_ | new_G4228_;
  assign new_G4214_ = ~new_G4205_ & new_G4231_;
  assign new_G4215_ = ~new_G4207_ & new_G4219_;
  assign new_G4216_ = new_G4207_ & ~new_G4219_;
  assign new_G4217_ = G4193 & ~G4194;
  assign new_G4218_ = ~new_G4240_ | ~new_G4241_;
  assign new_G4219_ = new_G4233_ | new_G4235_;
  assign new_G4220_ = new_G4243_ | new_G4242_;
  assign new_G4221_ = new_G4237_ | new_G4236_;
  assign new_G4222_ = ~new_G4245_ | ~new_G4244_;
  assign new_G4223_ = ~new_G4246_ & new_G4247_;
  assign new_G4224_ = new_G4246_ & ~new_G4247_;
  assign new_G4225_ = ~G4193 & G4194;
  assign new_G4226_ = G4193 & ~G4194;
  assign new_G4227_ = ~new_G4209_ | new_G4219_;
  assign new_G4228_ = new_G4209_ & new_G4219_;
  assign new_G4229_ = ~new_G4209_ & ~new_G4219_;
  assign new_G4230_ = new_G4251_ | new_G4250_;
  assign new_G4231_ = G4197 | new_G4230_;
  assign new_G4232_ = new_G4255_ | new_G4254_;
  assign new_G4233_ = ~G4197 & new_G4232_;
  assign new_G4234_ = new_G4253_ | new_G4252_;
  assign new_G4235_ = G4197 & new_G4234_;
  assign new_G4236_ = G4195 & ~new_G4205_;
  assign new_G4237_ = ~G4195 & new_G4205_;
  assign new_G4238_ = ~G4194 | ~new_G4219_;
  assign new_G4239_ = new_G4205_ & new_G4238_;
  assign new_G4240_ = ~new_G4205_ & ~new_G4239_;
  assign new_G4241_ = new_G4205_ | new_G4238_;
  assign new_G4242_ = ~G4195 & G4196;
  assign new_G4243_ = G4195 & ~G4196;
  assign new_G4244_ = new_G4212_ | new_G4249_;
  assign new_G4245_ = ~new_G4212_ & ~new_G4248_;
  assign new_G4246_ = G4195 | new_G4212_;
  assign new_G4247_ = G4195 | G4196;
  assign new_G4248_ = new_G4212_ & new_G4249_;
  assign new_G4249_ = ~G4194 | ~new_G4219_;
  assign new_G4250_ = new_G4227_ & new_G4247_;
  assign new_G4251_ = ~new_G4227_ & ~new_G4247_;
  assign new_G4252_ = new_G4256_ | new_G4257_;
  assign new_G4253_ = ~G4198 & new_G4212_;
  assign new_G4254_ = new_G4258_ | new_G4259_;
  assign new_G4255_ = G4198 & new_G4212_;
  assign new_G4256_ = ~G4198 & ~new_G4212_;
  assign new_G4257_ = G4198 & ~new_G4212_;
  assign new_G4258_ = G4198 & ~new_G4212_;
  assign new_G4259_ = ~G4198 & new_G4212_;
  assign new_G4266_ = new_G4273_ & new_G4272_;
  assign new_G4267_ = new_G4275_ | new_G4274_;
  assign new_G4268_ = new_G4277_ | new_G4276_;
  assign new_G4269_ = new_G4279_ & new_G4278_;
  assign new_G4270_ = new_G4279_ & new_G4280_;
  assign new_G4271_ = new_G4272_ | new_G4281_;
  assign new_G4272_ = G4261 | new_G4284_;
  assign new_G4273_ = new_G4283_ | new_G4282_;
  assign new_G4274_ = new_G4288_ & new_G4287_;
  assign new_G4275_ = new_G4286_ & new_G4285_;
  assign new_G4276_ = new_G4291_ | new_G4290_;
  assign new_G4277_ = new_G4286_ & new_G4289_;
  assign new_G4278_ = G4261 | new_G4294_;
  assign new_G4279_ = new_G4293_ | new_G4292_;
  assign new_G4280_ = new_G4296_ | new_G4295_;
  assign new_G4281_ = ~new_G4272_ & new_G4298_;
  assign new_G4282_ = ~new_G4274_ & new_G4286_;
  assign new_G4283_ = new_G4274_ & ~new_G4286_;
  assign new_G4284_ = G4260 & ~G4261;
  assign new_G4285_ = ~new_G4307_ | ~new_G4308_;
  assign new_G4286_ = new_G4300_ | new_G4302_;
  assign new_G4287_ = new_G4310_ | new_G4309_;
  assign new_G4288_ = new_G4304_ | new_G4303_;
  assign new_G4289_ = ~new_G4312_ | ~new_G4311_;
  assign new_G4290_ = ~new_G4313_ & new_G4314_;
  assign new_G4291_ = new_G4313_ & ~new_G4314_;
  assign new_G4292_ = ~G4260 & G4261;
  assign new_G4293_ = G4260 & ~G4261;
  assign new_G4294_ = ~new_G4276_ | new_G4286_;
  assign new_G4295_ = new_G4276_ & new_G4286_;
  assign new_G4296_ = ~new_G4276_ & ~new_G4286_;
  assign new_G4297_ = new_G4318_ | new_G4317_;
  assign new_G4298_ = G4264 | new_G4297_;
  assign new_G4299_ = new_G4322_ | new_G4321_;
  assign new_G4300_ = ~G4264 & new_G4299_;
  assign new_G4301_ = new_G4320_ | new_G4319_;
  assign new_G4302_ = G4264 & new_G4301_;
  assign new_G4303_ = G4262 & ~new_G4272_;
  assign new_G4304_ = ~G4262 & new_G4272_;
  assign new_G4305_ = ~G4261 | ~new_G4286_;
  assign new_G4306_ = new_G4272_ & new_G4305_;
  assign new_G4307_ = ~new_G4272_ & ~new_G4306_;
  assign new_G4308_ = new_G4272_ | new_G4305_;
  assign new_G4309_ = ~G4262 & G4263;
  assign new_G4310_ = G4262 & ~G4263;
  assign new_G4311_ = new_G4279_ | new_G4316_;
  assign new_G4312_ = ~new_G4279_ & ~new_G4315_;
  assign new_G4313_ = G4262 | new_G4279_;
  assign new_G4314_ = G4262 | G4263;
  assign new_G4315_ = new_G4279_ & new_G4316_;
  assign new_G4316_ = ~G4261 | ~new_G4286_;
  assign new_G4317_ = new_G4294_ & new_G4314_;
  assign new_G4318_ = ~new_G4294_ & ~new_G4314_;
  assign new_G4319_ = new_G4323_ | new_G4324_;
  assign new_G4320_ = ~G4265 & new_G4279_;
  assign new_G4321_ = new_G4325_ | new_G4326_;
  assign new_G4322_ = G4265 & new_G4279_;
  assign new_G4323_ = ~G4265 & ~new_G4279_;
  assign new_G4324_ = G4265 & ~new_G4279_;
  assign new_G4325_ = G4265 & ~new_G4279_;
  assign new_G4326_ = ~G4265 & new_G4279_;
  assign new_G4333_ = new_G4340_ & new_G4339_;
  assign new_G4334_ = new_G4342_ | new_G4341_;
  assign new_G4335_ = new_G4344_ | new_G4343_;
  assign new_G4336_ = new_G4346_ & new_G4345_;
  assign new_G4337_ = new_G4346_ & new_G4347_;
  assign new_G4338_ = new_G4339_ | new_G4348_;
  assign new_G4339_ = G4328 | new_G4351_;
  assign new_G4340_ = new_G4350_ | new_G4349_;
  assign new_G4341_ = new_G4355_ & new_G4354_;
  assign new_G4342_ = new_G4353_ & new_G4352_;
  assign new_G4343_ = new_G4358_ | new_G4357_;
  assign new_G4344_ = new_G4353_ & new_G4356_;
  assign new_G4345_ = G4328 | new_G4361_;
  assign new_G4346_ = new_G4360_ | new_G4359_;
  assign new_G4347_ = new_G4363_ | new_G4362_;
  assign new_G4348_ = ~new_G4339_ & new_G4365_;
  assign new_G4349_ = ~new_G4341_ & new_G4353_;
  assign new_G4350_ = new_G4341_ & ~new_G4353_;
  assign new_G4351_ = G4327 & ~G4328;
  assign new_G4352_ = ~new_G4374_ | ~new_G4375_;
  assign new_G4353_ = new_G4367_ | new_G4369_;
  assign new_G4354_ = new_G4377_ | new_G4376_;
  assign new_G4355_ = new_G4371_ | new_G4370_;
  assign new_G4356_ = ~new_G4379_ | ~new_G4378_;
  assign new_G4357_ = ~new_G4380_ & new_G4381_;
  assign new_G4358_ = new_G4380_ & ~new_G4381_;
  assign new_G4359_ = ~G4327 & G4328;
  assign new_G4360_ = G4327 & ~G4328;
  assign new_G4361_ = ~new_G4343_ | new_G4353_;
  assign new_G4362_ = new_G4343_ & new_G4353_;
  assign new_G4363_ = ~new_G4343_ & ~new_G4353_;
  assign new_G4364_ = new_G4385_ | new_G4384_;
  assign new_G4365_ = G4331 | new_G4364_;
  assign new_G4366_ = new_G4389_ | new_G4388_;
  assign new_G4367_ = ~G4331 & new_G4366_;
  assign new_G4368_ = new_G4387_ | new_G4386_;
  assign new_G4369_ = G4331 & new_G4368_;
  assign new_G4370_ = G4329 & ~new_G4339_;
  assign new_G4371_ = ~G4329 & new_G4339_;
  assign new_G4372_ = ~G4328 | ~new_G4353_;
  assign new_G4373_ = new_G4339_ & new_G4372_;
  assign new_G4374_ = ~new_G4339_ & ~new_G4373_;
  assign new_G4375_ = new_G4339_ | new_G4372_;
  assign new_G4376_ = ~G4329 & G4330;
  assign new_G4377_ = G4329 & ~G4330;
  assign new_G4378_ = new_G4346_ | new_G4383_;
  assign new_G4379_ = ~new_G4346_ & ~new_G4382_;
  assign new_G4380_ = G4329 | new_G4346_;
  assign new_G4381_ = G4329 | G4330;
  assign new_G4382_ = new_G4346_ & new_G4383_;
  assign new_G4383_ = ~G4328 | ~new_G4353_;
  assign new_G4384_ = new_G4361_ & new_G4381_;
  assign new_G4385_ = ~new_G4361_ & ~new_G4381_;
  assign new_G4386_ = new_G4390_ | new_G4391_;
  assign new_G4387_ = ~G4332 & new_G4346_;
  assign new_G4388_ = new_G4392_ | new_G4393_;
  assign new_G4389_ = G4332 & new_G4346_;
  assign new_G4390_ = ~G4332 & ~new_G4346_;
  assign new_G4391_ = G4332 & ~new_G4346_;
  assign new_G4392_ = G4332 & ~new_G4346_;
  assign new_G4393_ = ~G4332 & new_G4346_;
  assign new_G4400_ = new_G4407_ & new_G4406_;
  assign new_G4401_ = new_G4409_ | new_G4408_;
  assign new_G4402_ = new_G4411_ | new_G4410_;
  assign new_G4403_ = new_G4413_ & new_G4412_;
  assign new_G4404_ = new_G4413_ & new_G4414_;
  assign new_G4405_ = new_G4406_ | new_G4415_;
  assign new_G4406_ = G4395 | new_G4418_;
  assign new_G4407_ = new_G4417_ | new_G4416_;
  assign new_G4408_ = new_G4422_ & new_G4421_;
  assign new_G4409_ = new_G4420_ & new_G4419_;
  assign new_G4410_ = new_G4425_ | new_G4424_;
  assign new_G4411_ = new_G4420_ & new_G4423_;
  assign new_G4412_ = G4395 | new_G4428_;
  assign new_G4413_ = new_G4427_ | new_G4426_;
  assign new_G4414_ = new_G4430_ | new_G4429_;
  assign new_G4415_ = ~new_G4406_ & new_G4432_;
  assign new_G4416_ = ~new_G4408_ & new_G4420_;
  assign new_G4417_ = new_G4408_ & ~new_G4420_;
  assign new_G4418_ = G4394 & ~G4395;
  assign new_G4419_ = ~new_G4441_ | ~new_G4442_;
  assign new_G4420_ = new_G4434_ | new_G4436_;
  assign new_G4421_ = new_G4444_ | new_G4443_;
  assign new_G4422_ = new_G4438_ | new_G4437_;
  assign new_G4423_ = ~new_G4446_ | ~new_G4445_;
  assign new_G4424_ = ~new_G4447_ & new_G4448_;
  assign new_G4425_ = new_G4447_ & ~new_G4448_;
  assign new_G4426_ = ~G4394 & G4395;
  assign new_G4427_ = G4394 & ~G4395;
  assign new_G4428_ = ~new_G4410_ | new_G4420_;
  assign new_G4429_ = new_G4410_ & new_G4420_;
  assign new_G4430_ = ~new_G4410_ & ~new_G4420_;
  assign new_G4431_ = new_G4452_ | new_G4451_;
  assign new_G4432_ = G4398 | new_G4431_;
  assign new_G4433_ = new_G4456_ | new_G4455_;
  assign new_G4434_ = ~G4398 & new_G4433_;
  assign new_G4435_ = new_G4454_ | new_G4453_;
  assign new_G4436_ = G4398 & new_G4435_;
  assign new_G4437_ = G4396 & ~new_G4406_;
  assign new_G4438_ = ~G4396 & new_G4406_;
  assign new_G4439_ = ~G4395 | ~new_G4420_;
  assign new_G4440_ = new_G4406_ & new_G4439_;
  assign new_G4441_ = ~new_G4406_ & ~new_G4440_;
  assign new_G4442_ = new_G4406_ | new_G4439_;
  assign new_G4443_ = ~G4396 & G4397;
  assign new_G4444_ = G4396 & ~G4397;
  assign new_G4445_ = new_G4413_ | new_G4450_;
  assign new_G4446_ = ~new_G4413_ & ~new_G4449_;
  assign new_G4447_ = G4396 | new_G4413_;
  assign new_G4448_ = G4396 | G4397;
  assign new_G4449_ = new_G4413_ & new_G4450_;
  assign new_G4450_ = ~G4395 | ~new_G4420_;
  assign new_G4451_ = new_G4428_ & new_G4448_;
  assign new_G4452_ = ~new_G4428_ & ~new_G4448_;
  assign new_G4453_ = new_G4457_ | new_G4458_;
  assign new_G4454_ = ~G4399 & new_G4413_;
  assign new_G4455_ = new_G4459_ | new_G4460_;
  assign new_G4456_ = G4399 & new_G4413_;
  assign new_G4457_ = ~G4399 & ~new_G4413_;
  assign new_G4458_ = G4399 & ~new_G4413_;
  assign new_G4459_ = G4399 & ~new_G4413_;
  assign new_G4460_ = ~G4399 & new_G4413_;
  assign new_G4467_ = new_G4474_ & new_G4473_;
  assign new_G4468_ = new_G4476_ | new_G4475_;
  assign new_G4469_ = new_G4478_ | new_G4477_;
  assign new_G4470_ = new_G4480_ & new_G4479_;
  assign new_G4471_ = new_G4480_ & new_G4481_;
  assign new_G4472_ = new_G4473_ | new_G4482_;
  assign new_G4473_ = G4462 | new_G4485_;
  assign new_G4474_ = new_G4484_ | new_G4483_;
  assign new_G4475_ = new_G4489_ & new_G4488_;
  assign new_G4476_ = new_G4487_ & new_G4486_;
  assign new_G4477_ = new_G4492_ | new_G4491_;
  assign new_G4478_ = new_G4487_ & new_G4490_;
  assign new_G4479_ = G4462 | new_G4495_;
  assign new_G4480_ = new_G4494_ | new_G4493_;
  assign new_G4481_ = new_G4497_ | new_G4496_;
  assign new_G4482_ = ~new_G4473_ & new_G4499_;
  assign new_G4483_ = ~new_G4475_ & new_G4487_;
  assign new_G4484_ = new_G4475_ & ~new_G4487_;
  assign new_G4485_ = G4461 & ~G4462;
  assign new_G4486_ = ~new_G4508_ | ~new_G4509_;
  assign new_G4487_ = new_G4501_ | new_G4503_;
  assign new_G4488_ = new_G4511_ | new_G4510_;
  assign new_G4489_ = new_G4505_ | new_G4504_;
  assign new_G4490_ = ~new_G4513_ | ~new_G4512_;
  assign new_G4491_ = ~new_G4514_ & new_G4515_;
  assign new_G4492_ = new_G4514_ & ~new_G4515_;
  assign new_G4493_ = ~G4461 & G4462;
  assign new_G4494_ = G4461 & ~G4462;
  assign new_G4495_ = ~new_G4477_ | new_G4487_;
  assign new_G4496_ = new_G4477_ & new_G4487_;
  assign new_G4497_ = ~new_G4477_ & ~new_G4487_;
  assign new_G4498_ = new_G4519_ | new_G4518_;
  assign new_G4499_ = G4465 | new_G4498_;
  assign new_G4500_ = new_G4523_ | new_G4522_;
  assign new_G4501_ = ~G4465 & new_G4500_;
  assign new_G4502_ = new_G4521_ | new_G4520_;
  assign new_G4503_ = G4465 & new_G4502_;
  assign new_G4504_ = G4463 & ~new_G4473_;
  assign new_G4505_ = ~G4463 & new_G4473_;
  assign new_G4506_ = ~G4462 | ~new_G4487_;
  assign new_G4507_ = new_G4473_ & new_G4506_;
  assign new_G4508_ = ~new_G4473_ & ~new_G4507_;
  assign new_G4509_ = new_G4473_ | new_G4506_;
  assign new_G4510_ = ~G4463 & G4464;
  assign new_G4511_ = G4463 & ~G4464;
  assign new_G4512_ = new_G4480_ | new_G4517_;
  assign new_G4513_ = ~new_G4480_ & ~new_G4516_;
  assign new_G4514_ = G4463 | new_G4480_;
  assign new_G4515_ = G4463 | G4464;
  assign new_G4516_ = new_G4480_ & new_G4517_;
  assign new_G4517_ = ~G4462 | ~new_G4487_;
  assign new_G4518_ = new_G4495_ & new_G4515_;
  assign new_G4519_ = ~new_G4495_ & ~new_G4515_;
  assign new_G4520_ = new_G4524_ | new_G4525_;
  assign new_G4521_ = ~G4466 & new_G4480_;
  assign new_G4522_ = new_G4526_ | new_G4527_;
  assign new_G4523_ = G4466 & new_G4480_;
  assign new_G4524_ = ~G4466 & ~new_G4480_;
  assign new_G4525_ = G4466 & ~new_G4480_;
  assign new_G4526_ = G4466 & ~new_G4480_;
  assign new_G4527_ = ~G4466 & new_G4480_;
  assign new_G4534_ = new_G4541_ & new_G4540_;
  assign new_G4535_ = new_G4543_ | new_G4542_;
  assign new_G4536_ = new_G4545_ | new_G4544_;
  assign new_G4537_ = new_G4547_ & new_G4546_;
  assign new_G4538_ = new_G4547_ & new_G4548_;
  assign new_G4539_ = new_G4540_ | new_G4549_;
  assign new_G4540_ = G4529 | new_G4552_;
  assign new_G4541_ = new_G4551_ | new_G4550_;
  assign new_G4542_ = new_G4556_ & new_G4555_;
  assign new_G4543_ = new_G4554_ & new_G4553_;
  assign new_G4544_ = new_G4559_ | new_G4558_;
  assign new_G4545_ = new_G4554_ & new_G4557_;
  assign new_G4546_ = G4529 | new_G4562_;
  assign new_G4547_ = new_G4561_ | new_G4560_;
  assign new_G4548_ = new_G4564_ | new_G4563_;
  assign new_G4549_ = ~new_G4540_ & new_G4566_;
  assign new_G4550_ = ~new_G4542_ & new_G4554_;
  assign new_G4551_ = new_G4542_ & ~new_G4554_;
  assign new_G4552_ = G4528 & ~G4529;
  assign new_G4553_ = ~new_G4575_ | ~new_G4576_;
  assign new_G4554_ = new_G4568_ | new_G4570_;
  assign new_G4555_ = new_G4578_ | new_G4577_;
  assign new_G4556_ = new_G4572_ | new_G4571_;
  assign new_G4557_ = ~new_G4580_ | ~new_G4579_;
  assign new_G4558_ = ~new_G4581_ & new_G4582_;
  assign new_G4559_ = new_G4581_ & ~new_G4582_;
  assign new_G4560_ = ~G4528 & G4529;
  assign new_G4561_ = G4528 & ~G4529;
  assign new_G4562_ = ~new_G4544_ | new_G4554_;
  assign new_G4563_ = new_G4544_ & new_G4554_;
  assign new_G4564_ = ~new_G4544_ & ~new_G4554_;
  assign new_G4565_ = new_G4586_ | new_G4585_;
  assign new_G4566_ = G4532 | new_G4565_;
  assign new_G4567_ = new_G4590_ | new_G4589_;
  assign new_G4568_ = ~G4532 & new_G4567_;
  assign new_G4569_ = new_G4588_ | new_G4587_;
  assign new_G4570_ = G4532 & new_G4569_;
  assign new_G4571_ = G4530 & ~new_G4540_;
  assign new_G4572_ = ~G4530 & new_G4540_;
  assign new_G4573_ = ~G4529 | ~new_G4554_;
  assign new_G4574_ = new_G4540_ & new_G4573_;
  assign new_G4575_ = ~new_G4540_ & ~new_G4574_;
  assign new_G4576_ = new_G4540_ | new_G4573_;
  assign new_G4577_ = ~G4530 & G4531;
  assign new_G4578_ = G4530 & ~G4531;
  assign new_G4579_ = new_G4547_ | new_G4584_;
  assign new_G4580_ = ~new_G4547_ & ~new_G4583_;
  assign new_G4581_ = G4530 | new_G4547_;
  assign new_G4582_ = G4530 | G4531;
  assign new_G4583_ = new_G4547_ & new_G4584_;
  assign new_G4584_ = ~G4529 | ~new_G4554_;
  assign new_G4585_ = new_G4562_ & new_G4582_;
  assign new_G4586_ = ~new_G4562_ & ~new_G4582_;
  assign new_G4587_ = new_G4591_ | new_G4592_;
  assign new_G4588_ = ~G4533 & new_G4547_;
  assign new_G4589_ = new_G4593_ | new_G4594_;
  assign new_G4590_ = G4533 & new_G4547_;
  assign new_G4591_ = ~G4533 & ~new_G4547_;
  assign new_G4592_ = G4533 & ~new_G4547_;
  assign new_G4593_ = G4533 & ~new_G4547_;
  assign new_G4594_ = ~G4533 & new_G4547_;
  assign new_G4601_ = new_G4608_ & new_G4607_;
  assign new_G4602_ = new_G4610_ | new_G4609_;
  assign new_G4603_ = new_G4612_ | new_G4611_;
  assign new_G4604_ = new_G4614_ & new_G4613_;
  assign new_G4605_ = new_G4614_ & new_G4615_;
  assign new_G4606_ = new_G4607_ | new_G4616_;
  assign new_G4607_ = G4596 | new_G4619_;
  assign new_G4608_ = new_G4618_ | new_G4617_;
  assign new_G4609_ = new_G4623_ & new_G4622_;
  assign new_G4610_ = new_G4621_ & new_G4620_;
  assign new_G4611_ = new_G4626_ | new_G4625_;
  assign new_G4612_ = new_G4621_ & new_G4624_;
  assign new_G4613_ = G4596 | new_G4629_;
  assign new_G4614_ = new_G4628_ | new_G4627_;
  assign new_G4615_ = new_G4631_ | new_G4630_;
  assign new_G4616_ = ~new_G4607_ & new_G4633_;
  assign new_G4617_ = ~new_G4609_ & new_G4621_;
  assign new_G4618_ = new_G4609_ & ~new_G4621_;
  assign new_G4619_ = G4595 & ~G4596;
  assign new_G4620_ = ~new_G4642_ | ~new_G4643_;
  assign new_G4621_ = new_G4635_ | new_G4637_;
  assign new_G4622_ = new_G4645_ | new_G4644_;
  assign new_G4623_ = new_G4639_ | new_G4638_;
  assign new_G4624_ = ~new_G4647_ | ~new_G4646_;
  assign new_G4625_ = ~new_G4648_ & new_G4649_;
  assign new_G4626_ = new_G4648_ & ~new_G4649_;
  assign new_G4627_ = ~G4595 & G4596;
  assign new_G4628_ = G4595 & ~G4596;
  assign new_G4629_ = ~new_G4611_ | new_G4621_;
  assign new_G4630_ = new_G4611_ & new_G4621_;
  assign new_G4631_ = ~new_G4611_ & ~new_G4621_;
  assign new_G4632_ = new_G4653_ | new_G4652_;
  assign new_G4633_ = G4599 | new_G4632_;
  assign new_G4634_ = new_G4657_ | new_G4656_;
  assign new_G4635_ = ~G4599 & new_G4634_;
  assign new_G4636_ = new_G4655_ | new_G4654_;
  assign new_G4637_ = G4599 & new_G4636_;
  assign new_G4638_ = G4597 & ~new_G4607_;
  assign new_G4639_ = ~G4597 & new_G4607_;
  assign new_G4640_ = ~G4596 | ~new_G4621_;
  assign new_G4641_ = new_G4607_ & new_G4640_;
  assign new_G4642_ = ~new_G4607_ & ~new_G4641_;
  assign new_G4643_ = new_G4607_ | new_G4640_;
  assign new_G4644_ = ~G4597 & G4598;
  assign new_G4645_ = G4597 & ~G4598;
  assign new_G4646_ = new_G4614_ | new_G4651_;
  assign new_G4647_ = ~new_G4614_ & ~new_G4650_;
  assign new_G4648_ = G4597 | new_G4614_;
  assign new_G4649_ = G4597 | G4598;
  assign new_G4650_ = new_G4614_ & new_G4651_;
  assign new_G4651_ = ~G4596 | ~new_G4621_;
  assign new_G4652_ = new_G4629_ & new_G4649_;
  assign new_G4653_ = ~new_G4629_ & ~new_G4649_;
  assign new_G4654_ = new_G4658_ | new_G4659_;
  assign new_G4655_ = ~G4600 & new_G4614_;
  assign new_G4656_ = new_G4660_ | new_G4661_;
  assign new_G4657_ = G4600 & new_G4614_;
  assign new_G4658_ = ~G4600 & ~new_G4614_;
  assign new_G4659_ = G4600 & ~new_G4614_;
  assign new_G4660_ = G4600 & ~new_G4614_;
  assign new_G4661_ = ~G4600 & new_G4614_;
  assign new_G4668_ = new_G4675_ & new_G4674_;
  assign new_G4669_ = new_G4677_ | new_G4676_;
  assign new_G4670_ = new_G4679_ | new_G4678_;
  assign new_G4671_ = new_G4681_ & new_G4680_;
  assign new_G4672_ = new_G4681_ & new_G4682_;
  assign new_G4673_ = new_G4674_ | new_G4683_;
  assign new_G4674_ = G4663 | new_G4686_;
  assign new_G4675_ = new_G4685_ | new_G4684_;
  assign new_G4676_ = new_G4690_ & new_G4689_;
  assign new_G4677_ = new_G4688_ & new_G4687_;
  assign new_G4678_ = new_G4693_ | new_G4692_;
  assign new_G4679_ = new_G4688_ & new_G4691_;
  assign new_G4680_ = G4663 | new_G4696_;
  assign new_G4681_ = new_G4695_ | new_G4694_;
  assign new_G4682_ = new_G4698_ | new_G4697_;
  assign new_G4683_ = ~new_G4674_ & new_G4700_;
  assign new_G4684_ = ~new_G4676_ & new_G4688_;
  assign new_G4685_ = new_G4676_ & ~new_G4688_;
  assign new_G4686_ = G4662 & ~G4663;
  assign new_G4687_ = ~new_G4709_ | ~new_G4710_;
  assign new_G4688_ = new_G4702_ | new_G4704_;
  assign new_G4689_ = new_G4712_ | new_G4711_;
  assign new_G4690_ = new_G4706_ | new_G4705_;
  assign new_G4691_ = ~new_G4714_ | ~new_G4713_;
  assign new_G4692_ = ~new_G4715_ & new_G4716_;
  assign new_G4693_ = new_G4715_ & ~new_G4716_;
  assign new_G4694_ = ~G4662 & G4663;
  assign new_G4695_ = G4662 & ~G4663;
  assign new_G4696_ = ~new_G4678_ | new_G4688_;
  assign new_G4697_ = new_G4678_ & new_G4688_;
  assign new_G4698_ = ~new_G4678_ & ~new_G4688_;
  assign new_G4699_ = new_G4720_ | new_G4719_;
  assign new_G4700_ = G4666 | new_G4699_;
  assign new_G4701_ = new_G4724_ | new_G4723_;
  assign new_G4702_ = ~G4666 & new_G4701_;
  assign new_G4703_ = new_G4722_ | new_G4721_;
  assign new_G4704_ = G4666 & new_G4703_;
  assign new_G4705_ = G4664 & ~new_G4674_;
  assign new_G4706_ = ~G4664 & new_G4674_;
  assign new_G4707_ = ~G4663 | ~new_G4688_;
  assign new_G4708_ = new_G4674_ & new_G4707_;
  assign new_G4709_ = ~new_G4674_ & ~new_G4708_;
  assign new_G4710_ = new_G4674_ | new_G4707_;
  assign new_G4711_ = ~G4664 & G4665;
  assign new_G4712_ = G4664 & ~G4665;
  assign new_G4713_ = new_G4681_ | new_G4718_;
  assign new_G4714_ = ~new_G4681_ & ~new_G4717_;
  assign new_G4715_ = G4664 | new_G4681_;
  assign new_G4716_ = G4664 | G4665;
  assign new_G4717_ = new_G4681_ & new_G4718_;
  assign new_G4718_ = ~G4663 | ~new_G4688_;
  assign new_G4719_ = new_G4696_ & new_G4716_;
  assign new_G4720_ = ~new_G4696_ & ~new_G4716_;
  assign new_G4721_ = new_G4725_ | new_G4726_;
  assign new_G4722_ = ~G4667 & new_G4681_;
  assign new_G4723_ = new_G4727_ | new_G4728_;
  assign new_G4724_ = G4667 & new_G4681_;
  assign new_G4725_ = ~G4667 & ~new_G4681_;
  assign new_G4726_ = G4667 & ~new_G4681_;
  assign new_G4727_ = G4667 & ~new_G4681_;
  assign new_G4728_ = ~G4667 & new_G4681_;
  assign new_G4735_ = new_G4742_ & new_G4741_;
  assign new_G4736_ = new_G4744_ | new_G4743_;
  assign new_G4737_ = new_G4746_ | new_G4745_;
  assign new_G4738_ = new_G4748_ & new_G4747_;
  assign new_G4739_ = new_G4748_ & new_G4749_;
  assign new_G4740_ = new_G4741_ | new_G4750_;
  assign new_G4741_ = G4730 | new_G4753_;
  assign new_G4742_ = new_G4752_ | new_G4751_;
  assign new_G4743_ = new_G4757_ & new_G4756_;
  assign new_G4744_ = new_G4755_ & new_G4754_;
  assign new_G4745_ = new_G4760_ | new_G4759_;
  assign new_G4746_ = new_G4755_ & new_G4758_;
  assign new_G4747_ = G4730 | new_G4763_;
  assign new_G4748_ = new_G4762_ | new_G4761_;
  assign new_G4749_ = new_G4765_ | new_G4764_;
  assign new_G4750_ = ~new_G4741_ & new_G4767_;
  assign new_G4751_ = ~new_G4743_ & new_G4755_;
  assign new_G4752_ = new_G4743_ & ~new_G4755_;
  assign new_G4753_ = G4729 & ~G4730;
  assign new_G4754_ = ~new_G4776_ | ~new_G4777_;
  assign new_G4755_ = new_G4769_ | new_G4771_;
  assign new_G4756_ = new_G4779_ | new_G4778_;
  assign new_G4757_ = new_G4773_ | new_G4772_;
  assign new_G4758_ = ~new_G4781_ | ~new_G4780_;
  assign new_G4759_ = ~new_G4782_ & new_G4783_;
  assign new_G4760_ = new_G4782_ & ~new_G4783_;
  assign new_G4761_ = ~G4729 & G4730;
  assign new_G4762_ = G4729 & ~G4730;
  assign new_G4763_ = ~new_G4745_ | new_G4755_;
  assign new_G4764_ = new_G4745_ & new_G4755_;
  assign new_G4765_ = ~new_G4745_ & ~new_G4755_;
  assign new_G4766_ = new_G4787_ | new_G4786_;
  assign new_G4767_ = G4733 | new_G4766_;
  assign new_G4768_ = new_G4791_ | new_G4790_;
  assign new_G4769_ = ~G4733 & new_G4768_;
  assign new_G4770_ = new_G4789_ | new_G4788_;
  assign new_G4771_ = G4733 & new_G4770_;
  assign new_G4772_ = G4731 & ~new_G4741_;
  assign new_G4773_ = ~G4731 & new_G4741_;
  assign new_G4774_ = ~G4730 | ~new_G4755_;
  assign new_G4775_ = new_G4741_ & new_G4774_;
  assign new_G4776_ = ~new_G4741_ & ~new_G4775_;
  assign new_G4777_ = new_G4741_ | new_G4774_;
  assign new_G4778_ = ~G4731 & G4732;
  assign new_G4779_ = G4731 & ~G4732;
  assign new_G4780_ = new_G4748_ | new_G4785_;
  assign new_G4781_ = ~new_G4748_ & ~new_G4784_;
  assign new_G4782_ = G4731 | new_G4748_;
  assign new_G4783_ = G4731 | G4732;
  assign new_G4784_ = new_G4748_ & new_G4785_;
  assign new_G4785_ = ~G4730 | ~new_G4755_;
  assign new_G4786_ = new_G4763_ & new_G4783_;
  assign new_G4787_ = ~new_G4763_ & ~new_G4783_;
  assign new_G4788_ = new_G4792_ | new_G4793_;
  assign new_G4789_ = ~G4734 & new_G4748_;
  assign new_G4790_ = new_G4794_ | new_G4795_;
  assign new_G4791_ = G4734 & new_G4748_;
  assign new_G4792_ = ~G4734 & ~new_G4748_;
  assign new_G4793_ = G4734 & ~new_G4748_;
  assign new_G4794_ = G4734 & ~new_G4748_;
  assign new_G4795_ = ~G4734 & new_G4748_;
  assign new_G4802_ = new_G4809_ & new_G4808_;
  assign new_G4803_ = new_G4811_ | new_G4810_;
  assign new_G4804_ = new_G4813_ | new_G4812_;
  assign new_G4805_ = new_G4815_ & new_G4814_;
  assign new_G4806_ = new_G4815_ & new_G4816_;
  assign new_G4807_ = new_G4808_ | new_G4817_;
  assign new_G4808_ = G4797 | new_G4820_;
  assign new_G4809_ = new_G4819_ | new_G4818_;
  assign new_G4810_ = new_G4824_ & new_G4823_;
  assign new_G4811_ = new_G4822_ & new_G4821_;
  assign new_G4812_ = new_G4827_ | new_G4826_;
  assign new_G4813_ = new_G4822_ & new_G4825_;
  assign new_G4814_ = G4797 | new_G4830_;
  assign new_G4815_ = new_G4829_ | new_G4828_;
  assign new_G4816_ = new_G4832_ | new_G4831_;
  assign new_G4817_ = ~new_G4808_ & new_G4834_;
  assign new_G4818_ = ~new_G4810_ & new_G4822_;
  assign new_G4819_ = new_G4810_ & ~new_G4822_;
  assign new_G4820_ = G4796 & ~G4797;
  assign new_G4821_ = ~new_G4843_ | ~new_G4844_;
  assign new_G4822_ = new_G4836_ | new_G4838_;
  assign new_G4823_ = new_G4846_ | new_G4845_;
  assign new_G4824_ = new_G4840_ | new_G4839_;
  assign new_G4825_ = ~new_G4848_ | ~new_G4847_;
  assign new_G4826_ = ~new_G4849_ & new_G4850_;
  assign new_G4827_ = new_G4849_ & ~new_G4850_;
  assign new_G4828_ = ~G4796 & G4797;
  assign new_G4829_ = G4796 & ~G4797;
  assign new_G4830_ = ~new_G4812_ | new_G4822_;
  assign new_G4831_ = new_G4812_ & new_G4822_;
  assign new_G4832_ = ~new_G4812_ & ~new_G4822_;
  assign new_G4833_ = new_G4854_ | new_G4853_;
  assign new_G4834_ = G4800 | new_G4833_;
  assign new_G4835_ = new_G4858_ | new_G4857_;
  assign new_G4836_ = ~G4800 & new_G4835_;
  assign new_G4837_ = new_G4856_ | new_G4855_;
  assign new_G4838_ = G4800 & new_G4837_;
  assign new_G4839_ = G4798 & ~new_G4808_;
  assign new_G4840_ = ~G4798 & new_G4808_;
  assign new_G4841_ = ~G4797 | ~new_G4822_;
  assign new_G4842_ = new_G4808_ & new_G4841_;
  assign new_G4843_ = ~new_G4808_ & ~new_G4842_;
  assign new_G4844_ = new_G4808_ | new_G4841_;
  assign new_G4845_ = ~G4798 & G4799;
  assign new_G4846_ = G4798 & ~G4799;
  assign new_G4847_ = new_G4815_ | new_G4852_;
  assign new_G4848_ = ~new_G4815_ & ~new_G4851_;
  assign new_G4849_ = G4798 | new_G4815_;
  assign new_G4850_ = G4798 | G4799;
  assign new_G4851_ = new_G4815_ & new_G4852_;
  assign new_G4852_ = ~G4797 | ~new_G4822_;
  assign new_G4853_ = new_G4830_ & new_G4850_;
  assign new_G4854_ = ~new_G4830_ & ~new_G4850_;
  assign new_G4855_ = new_G4859_ | new_G4860_;
  assign new_G4856_ = ~G4801 & new_G4815_;
  assign new_G4857_ = new_G4861_ | new_G4862_;
  assign new_G4858_ = G4801 & new_G4815_;
  assign new_G4859_ = ~G4801 & ~new_G4815_;
  assign new_G4860_ = G4801 & ~new_G4815_;
  assign new_G4861_ = G4801 & ~new_G4815_;
  assign new_G4862_ = ~G4801 & new_G4815_;
  assign new_G4869_ = new_G4876_ & new_G4875_;
  assign new_G4870_ = new_G4878_ | new_G4877_;
  assign new_G4871_ = new_G4880_ | new_G4879_;
  assign new_G4872_ = new_G4882_ & new_G4881_;
  assign new_G4873_ = new_G4882_ & new_G4883_;
  assign new_G4874_ = new_G4875_ | new_G4884_;
  assign new_G4875_ = G4864 | new_G4887_;
  assign new_G4876_ = new_G4886_ | new_G4885_;
  assign new_G4877_ = new_G4891_ & new_G4890_;
  assign new_G4878_ = new_G4889_ & new_G4888_;
  assign new_G4879_ = new_G4894_ | new_G4893_;
  assign new_G4880_ = new_G4889_ & new_G4892_;
  assign new_G4881_ = G4864 | new_G4897_;
  assign new_G4882_ = new_G4896_ | new_G4895_;
  assign new_G4883_ = new_G4899_ | new_G4898_;
  assign new_G4884_ = ~new_G4875_ & new_G4901_;
  assign new_G4885_ = ~new_G4877_ & new_G4889_;
  assign new_G4886_ = new_G4877_ & ~new_G4889_;
  assign new_G4887_ = G4863 & ~G4864;
  assign new_G4888_ = ~new_G4910_ | ~new_G4911_;
  assign new_G4889_ = new_G4903_ | new_G4905_;
  assign new_G4890_ = new_G4913_ | new_G4912_;
  assign new_G4891_ = new_G4907_ | new_G4906_;
  assign new_G4892_ = ~new_G4915_ | ~new_G4914_;
  assign new_G4893_ = ~new_G4916_ & new_G4917_;
  assign new_G4894_ = new_G4916_ & ~new_G4917_;
  assign new_G4895_ = ~G4863 & G4864;
  assign new_G4896_ = G4863 & ~G4864;
  assign new_G4897_ = ~new_G4879_ | new_G4889_;
  assign new_G4898_ = new_G4879_ & new_G4889_;
  assign new_G4899_ = ~new_G4879_ & ~new_G4889_;
  assign new_G4900_ = new_G4921_ | new_G4920_;
  assign new_G4901_ = G4867 | new_G4900_;
  assign new_G4902_ = new_G4925_ | new_G4924_;
  assign new_G4903_ = ~G4867 & new_G4902_;
  assign new_G4904_ = new_G4923_ | new_G4922_;
  assign new_G4905_ = G4867 & new_G4904_;
  assign new_G4906_ = G4865 & ~new_G4875_;
  assign new_G4907_ = ~G4865 & new_G4875_;
  assign new_G4908_ = ~G4864 | ~new_G4889_;
  assign new_G4909_ = new_G4875_ & new_G4908_;
  assign new_G4910_ = ~new_G4875_ & ~new_G4909_;
  assign new_G4911_ = new_G4875_ | new_G4908_;
  assign new_G4912_ = ~G4865 & G4866;
  assign new_G4913_ = G4865 & ~G4866;
  assign new_G4914_ = new_G4882_ | new_G4919_;
  assign new_G4915_ = ~new_G4882_ & ~new_G4918_;
  assign new_G4916_ = G4865 | new_G4882_;
  assign new_G4917_ = G4865 | G4866;
  assign new_G4918_ = new_G4882_ & new_G4919_;
  assign new_G4919_ = ~G4864 | ~new_G4889_;
  assign new_G4920_ = new_G4897_ & new_G4917_;
  assign new_G4921_ = ~new_G4897_ & ~new_G4917_;
  assign new_G4922_ = new_G4926_ | new_G4927_;
  assign new_G4923_ = ~G4868 & new_G4882_;
  assign new_G4924_ = new_G4928_ | new_G4929_;
  assign new_G4925_ = G4868 & new_G4882_;
  assign new_G4926_ = ~G4868 & ~new_G4882_;
  assign new_G4927_ = G4868 & ~new_G4882_;
  assign new_G4928_ = G4868 & ~new_G4882_;
  assign new_G4929_ = ~G4868 & new_G4882_;
  assign new_G4936_ = new_G4943_ & new_G4942_;
  assign new_G4937_ = new_G4945_ | new_G4944_;
  assign new_G4938_ = new_G4947_ | new_G4946_;
  assign new_G4939_ = new_G4949_ & new_G4948_;
  assign new_G4940_ = new_G4949_ & new_G4950_;
  assign new_G4941_ = new_G4942_ | new_G4951_;
  assign new_G4942_ = G4931 | new_G4954_;
  assign new_G4943_ = new_G4953_ | new_G4952_;
  assign new_G4944_ = new_G4958_ & new_G4957_;
  assign new_G4945_ = new_G4956_ & new_G4955_;
  assign new_G4946_ = new_G4961_ | new_G4960_;
  assign new_G4947_ = new_G4956_ & new_G4959_;
  assign new_G4948_ = G4931 | new_G4964_;
  assign new_G4949_ = new_G4963_ | new_G4962_;
  assign new_G4950_ = new_G4966_ | new_G4965_;
  assign new_G4951_ = ~new_G4942_ & new_G4968_;
  assign new_G4952_ = ~new_G4944_ & new_G4956_;
  assign new_G4953_ = new_G4944_ & ~new_G4956_;
  assign new_G4954_ = G4930 & ~G4931;
  assign new_G4955_ = ~new_G4977_ | ~new_G4978_;
  assign new_G4956_ = new_G4970_ | new_G4972_;
  assign new_G4957_ = new_G4980_ | new_G4979_;
  assign new_G4958_ = new_G4974_ | new_G4973_;
  assign new_G4959_ = ~new_G4982_ | ~new_G4981_;
  assign new_G4960_ = ~new_G4983_ & new_G4984_;
  assign new_G4961_ = new_G4983_ & ~new_G4984_;
  assign new_G4962_ = ~G4930 & G4931;
  assign new_G4963_ = G4930 & ~G4931;
  assign new_G4964_ = ~new_G4946_ | new_G4956_;
  assign new_G4965_ = new_G4946_ & new_G4956_;
  assign new_G4966_ = ~new_G4946_ & ~new_G4956_;
  assign new_G4967_ = new_G4988_ | new_G4987_;
  assign new_G4968_ = G4934 | new_G4967_;
  assign new_G4969_ = new_G4992_ | new_G4991_;
  assign new_G4970_ = ~G4934 & new_G4969_;
  assign new_G4971_ = new_G4990_ | new_G4989_;
  assign new_G4972_ = G4934 & new_G4971_;
  assign new_G4973_ = G4932 & ~new_G4942_;
  assign new_G4974_ = ~G4932 & new_G4942_;
  assign new_G4975_ = ~G4931 | ~new_G4956_;
  assign new_G4976_ = new_G4942_ & new_G4975_;
  assign new_G4977_ = ~new_G4942_ & ~new_G4976_;
  assign new_G4978_ = new_G4942_ | new_G4975_;
  assign new_G4979_ = ~G4932 & G4933;
  assign new_G4980_ = G4932 & ~G4933;
  assign new_G4981_ = new_G4949_ | new_G4986_;
  assign new_G4982_ = ~new_G4949_ & ~new_G4985_;
  assign new_G4983_ = G4932 | new_G4949_;
  assign new_G4984_ = G4932 | G4933;
  assign new_G4985_ = new_G4949_ & new_G4986_;
  assign new_G4986_ = ~G4931 | ~new_G4956_;
  assign new_G4987_ = new_G4964_ & new_G4984_;
  assign new_G4988_ = ~new_G4964_ & ~new_G4984_;
  assign new_G4989_ = new_G4993_ | new_G4994_;
  assign new_G4990_ = ~G4935 & new_G4949_;
  assign new_G4991_ = new_G4995_ | new_G4996_;
  assign new_G4992_ = G4935 & new_G4949_;
  assign new_G4993_ = ~G4935 & ~new_G4949_;
  assign new_G4994_ = G4935 & ~new_G4949_;
  assign new_G4995_ = G4935 & ~new_G4949_;
  assign new_G4996_ = ~G4935 & new_G4949_;
  assign new_G5003_ = new_G5010_ & new_G5009_;
  assign new_G5004_ = new_G5012_ | new_G5011_;
  assign new_G5005_ = new_G5014_ | new_G5013_;
  assign new_G5006_ = new_G5016_ & new_G5015_;
  assign new_G5007_ = new_G5016_ & new_G5017_;
  assign new_G5008_ = new_G5009_ | new_G5018_;
  assign new_G5009_ = G4998 | new_G5021_;
  assign new_G5010_ = new_G5020_ | new_G5019_;
  assign new_G5011_ = new_G5025_ & new_G5024_;
  assign new_G5012_ = new_G5023_ & new_G5022_;
  assign new_G5013_ = new_G5028_ | new_G5027_;
  assign new_G5014_ = new_G5023_ & new_G5026_;
  assign new_G5015_ = G4998 | new_G5031_;
  assign new_G5016_ = new_G5030_ | new_G5029_;
  assign new_G5017_ = new_G5033_ | new_G5032_;
  assign new_G5018_ = ~new_G5009_ & new_G5035_;
  assign new_G5019_ = ~new_G5011_ & new_G5023_;
  assign new_G5020_ = new_G5011_ & ~new_G5023_;
  assign new_G5021_ = G4997 & ~G4998;
  assign new_G5022_ = ~new_G5044_ | ~new_G5045_;
  assign new_G5023_ = new_G5037_ | new_G5039_;
  assign new_G5024_ = new_G5047_ | new_G5046_;
  assign new_G5025_ = new_G5041_ | new_G5040_;
  assign new_G5026_ = ~new_G5049_ | ~new_G5048_;
  assign new_G5027_ = ~new_G5050_ & new_G5051_;
  assign new_G5028_ = new_G5050_ & ~new_G5051_;
  assign new_G5029_ = ~G4997 & G4998;
  assign new_G5030_ = G4997 & ~G4998;
  assign new_G5031_ = ~new_G5013_ | new_G5023_;
  assign new_G5032_ = new_G5013_ & new_G5023_;
  assign new_G5033_ = ~new_G5013_ & ~new_G5023_;
  assign new_G5034_ = new_G5055_ | new_G5054_;
  assign new_G5035_ = G5001 | new_G5034_;
  assign new_G5036_ = new_G5059_ | new_G5058_;
  assign new_G5037_ = ~G5001 & new_G5036_;
  assign new_G5038_ = new_G5057_ | new_G5056_;
  assign new_G5039_ = G5001 & new_G5038_;
  assign new_G5040_ = G4999 & ~new_G5009_;
  assign new_G5041_ = ~G4999 & new_G5009_;
  assign new_G5042_ = ~G4998 | ~new_G5023_;
  assign new_G5043_ = new_G5009_ & new_G5042_;
  assign new_G5044_ = ~new_G5009_ & ~new_G5043_;
  assign new_G5045_ = new_G5009_ | new_G5042_;
  assign new_G5046_ = ~G4999 & G5000;
  assign new_G5047_ = G4999 & ~G5000;
  assign new_G5048_ = new_G5016_ | new_G5053_;
  assign new_G5049_ = ~new_G5016_ & ~new_G5052_;
  assign new_G5050_ = G4999 | new_G5016_;
  assign new_G5051_ = G4999 | G5000;
  assign new_G5052_ = new_G5016_ & new_G5053_;
  assign new_G5053_ = ~G4998 | ~new_G5023_;
  assign new_G5054_ = new_G5031_ & new_G5051_;
  assign new_G5055_ = ~new_G5031_ & ~new_G5051_;
  assign new_G5056_ = new_G5060_ | new_G5061_;
  assign new_G5057_ = ~G5002 & new_G5016_;
  assign new_G5058_ = new_G5062_ | new_G5063_;
  assign new_G5059_ = G5002 & new_G5016_;
  assign new_G5060_ = ~G5002 & ~new_G5016_;
  assign new_G5061_ = G5002 & ~new_G5016_;
  assign new_G5062_ = G5002 & ~new_G5016_;
  assign new_G5063_ = ~G5002 & new_G5016_;
  assign new_G5070_ = new_G5077_ & new_G5076_;
  assign new_G5071_ = new_G5079_ | new_G5078_;
  assign new_G5072_ = new_G5081_ | new_G5080_;
  assign new_G5073_ = new_G5083_ & new_G5082_;
  assign new_G5074_ = new_G5083_ & new_G5084_;
  assign new_G5075_ = new_G5076_ | new_G5085_;
  assign new_G5076_ = G5065 | new_G5088_;
  assign new_G5077_ = new_G5087_ | new_G5086_;
  assign new_G5078_ = new_G5092_ & new_G5091_;
  assign new_G5079_ = new_G5090_ & new_G5089_;
  assign new_G5080_ = new_G5095_ | new_G5094_;
  assign new_G5081_ = new_G5090_ & new_G5093_;
  assign new_G5082_ = G5065 | new_G5098_;
  assign new_G5083_ = new_G5097_ | new_G5096_;
  assign new_G5084_ = new_G5100_ | new_G5099_;
  assign new_G5085_ = ~new_G5076_ & new_G5102_;
  assign new_G5086_ = ~new_G5078_ & new_G5090_;
  assign new_G5087_ = new_G5078_ & ~new_G5090_;
  assign new_G5088_ = G5064 & ~G5065;
  assign new_G5089_ = ~new_G5111_ | ~new_G5112_;
  assign new_G5090_ = new_G5104_ | new_G5106_;
  assign new_G5091_ = new_G5114_ | new_G5113_;
  assign new_G5092_ = new_G5108_ | new_G5107_;
  assign new_G5093_ = ~new_G5116_ | ~new_G5115_;
  assign new_G5094_ = ~new_G5117_ & new_G5118_;
  assign new_G5095_ = new_G5117_ & ~new_G5118_;
  assign new_G5096_ = ~G5064 & G5065;
  assign new_G5097_ = G5064 & ~G5065;
  assign new_G5098_ = ~new_G5080_ | new_G5090_;
  assign new_G5099_ = new_G5080_ & new_G5090_;
  assign new_G5100_ = ~new_G5080_ & ~new_G5090_;
  assign new_G5101_ = new_G5122_ | new_G5121_;
  assign new_G5102_ = G5068 | new_G5101_;
  assign new_G5103_ = new_G5126_ | new_G5125_;
  assign new_G5104_ = ~G5068 & new_G5103_;
  assign new_G5105_ = new_G5124_ | new_G5123_;
  assign new_G5106_ = G5068 & new_G5105_;
  assign new_G5107_ = G5066 & ~new_G5076_;
  assign new_G5108_ = ~G5066 & new_G5076_;
  assign new_G5109_ = ~G5065 | ~new_G5090_;
  assign new_G5110_ = new_G5076_ & new_G5109_;
  assign new_G5111_ = ~new_G5076_ & ~new_G5110_;
  assign new_G5112_ = new_G5076_ | new_G5109_;
  assign new_G5113_ = ~G5066 & G5067;
  assign new_G5114_ = G5066 & ~G5067;
  assign new_G5115_ = new_G5083_ | new_G5120_;
  assign new_G5116_ = ~new_G5083_ & ~new_G5119_;
  assign new_G5117_ = G5066 | new_G5083_;
  assign new_G5118_ = G5066 | G5067;
  assign new_G5119_ = new_G5083_ & new_G5120_;
  assign new_G5120_ = ~G5065 | ~new_G5090_;
  assign new_G5121_ = new_G5098_ & new_G5118_;
  assign new_G5122_ = ~new_G5098_ & ~new_G5118_;
  assign new_G5123_ = new_G5127_ | new_G5128_;
  assign new_G5124_ = ~G5069 & new_G5083_;
  assign new_G5125_ = new_G5129_ | new_G5130_;
  assign new_G5126_ = G5069 & new_G5083_;
  assign new_G5127_ = ~G5069 & ~new_G5083_;
  assign new_G5128_ = G5069 & ~new_G5083_;
  assign new_G5129_ = G5069 & ~new_G5083_;
  assign new_G5130_ = ~G5069 & new_G5083_;
  assign new_G5137_ = new_G5144_ & new_G5143_;
  assign new_G5138_ = new_G5146_ | new_G5145_;
  assign new_G5139_ = new_G5148_ | new_G5147_;
  assign new_G5140_ = new_G5150_ & new_G5149_;
  assign new_G5141_ = new_G5150_ & new_G5151_;
  assign new_G5142_ = new_G5143_ | new_G5152_;
  assign new_G5143_ = G5132 | new_G5155_;
  assign new_G5144_ = new_G5154_ | new_G5153_;
  assign new_G5145_ = new_G5159_ & new_G5158_;
  assign new_G5146_ = new_G5157_ & new_G5156_;
  assign new_G5147_ = new_G5162_ | new_G5161_;
  assign new_G5148_ = new_G5157_ & new_G5160_;
  assign new_G5149_ = G5132 | new_G5165_;
  assign new_G5150_ = new_G5164_ | new_G5163_;
  assign new_G5151_ = new_G5167_ | new_G5166_;
  assign new_G5152_ = ~new_G5143_ & new_G5169_;
  assign new_G5153_ = ~new_G5145_ & new_G5157_;
  assign new_G5154_ = new_G5145_ & ~new_G5157_;
  assign new_G5155_ = G5131 & ~G5132;
  assign new_G5156_ = ~new_G5178_ | ~new_G5179_;
  assign new_G5157_ = new_G5171_ | new_G5173_;
  assign new_G5158_ = new_G5181_ | new_G5180_;
  assign new_G5159_ = new_G5175_ | new_G5174_;
  assign new_G5160_ = ~new_G5183_ | ~new_G5182_;
  assign new_G5161_ = ~new_G5184_ & new_G5185_;
  assign new_G5162_ = new_G5184_ & ~new_G5185_;
  assign new_G5163_ = ~G5131 & G5132;
  assign new_G5164_ = G5131 & ~G5132;
  assign new_G5165_ = ~new_G5147_ | new_G5157_;
  assign new_G5166_ = new_G5147_ & new_G5157_;
  assign new_G5167_ = ~new_G5147_ & ~new_G5157_;
  assign new_G5168_ = new_G5189_ | new_G5188_;
  assign new_G5169_ = G5135 | new_G5168_;
  assign new_G5170_ = new_G5193_ | new_G5192_;
  assign new_G5171_ = ~G5135 & new_G5170_;
  assign new_G5172_ = new_G5191_ | new_G5190_;
  assign new_G5173_ = G5135 & new_G5172_;
  assign new_G5174_ = G5133 & ~new_G5143_;
  assign new_G5175_ = ~G5133 & new_G5143_;
  assign new_G5176_ = ~G5132 | ~new_G5157_;
  assign new_G5177_ = new_G5143_ & new_G5176_;
  assign new_G5178_ = ~new_G5143_ & ~new_G5177_;
  assign new_G5179_ = new_G5143_ | new_G5176_;
  assign new_G5180_ = ~G5133 & G5134;
  assign new_G5181_ = G5133 & ~G5134;
  assign new_G5182_ = new_G5150_ | new_G5187_;
  assign new_G5183_ = ~new_G5150_ & ~new_G5186_;
  assign new_G5184_ = G5133 | new_G5150_;
  assign new_G5185_ = G5133 | G5134;
  assign new_G5186_ = new_G5150_ & new_G5187_;
  assign new_G5187_ = ~G5132 | ~new_G5157_;
  assign new_G5188_ = new_G5165_ & new_G5185_;
  assign new_G5189_ = ~new_G5165_ & ~new_G5185_;
  assign new_G5190_ = new_G5194_ | new_G5195_;
  assign new_G5191_ = ~G5136 & new_G5150_;
  assign new_G5192_ = new_G5196_ | new_G5197_;
  assign new_G5193_ = G5136 & new_G5150_;
  assign new_G5194_ = ~G5136 & ~new_G5150_;
  assign new_G5195_ = G5136 & ~new_G5150_;
  assign new_G5196_ = G5136 & ~new_G5150_;
  assign new_G5197_ = ~G5136 & new_G5150_;
  assign new_G5204_ = new_G5211_ & new_G5210_;
  assign new_G5205_ = new_G5213_ | new_G5212_;
  assign new_G5206_ = new_G5215_ | new_G5214_;
  assign new_G5207_ = new_G5217_ & new_G5216_;
  assign new_G5208_ = new_G5217_ & new_G5218_;
  assign new_G5209_ = new_G5210_ | new_G5219_;
  assign new_G5210_ = G5199 | new_G5222_;
  assign new_G5211_ = new_G5221_ | new_G5220_;
  assign new_G5212_ = new_G5226_ & new_G5225_;
  assign new_G5213_ = new_G5224_ & new_G5223_;
  assign new_G5214_ = new_G5229_ | new_G5228_;
  assign new_G5215_ = new_G5224_ & new_G5227_;
  assign new_G5216_ = G5199 | new_G5232_;
  assign new_G5217_ = new_G5231_ | new_G5230_;
  assign new_G5218_ = new_G5234_ | new_G5233_;
  assign new_G5219_ = ~new_G5210_ & new_G5236_;
  assign new_G5220_ = ~new_G5212_ & new_G5224_;
  assign new_G5221_ = new_G5212_ & ~new_G5224_;
  assign new_G5222_ = G5198 & ~G5199;
  assign new_G5223_ = ~new_G5245_ | ~new_G5246_;
  assign new_G5224_ = new_G5238_ | new_G5240_;
  assign new_G5225_ = new_G5248_ | new_G5247_;
  assign new_G5226_ = new_G5242_ | new_G5241_;
  assign new_G5227_ = ~new_G5250_ | ~new_G5249_;
  assign new_G5228_ = ~new_G5251_ & new_G5252_;
  assign new_G5229_ = new_G5251_ & ~new_G5252_;
  assign new_G5230_ = ~G5198 & G5199;
  assign new_G5231_ = G5198 & ~G5199;
  assign new_G5232_ = ~new_G5214_ | new_G5224_;
  assign new_G5233_ = new_G5214_ & new_G5224_;
  assign new_G5234_ = ~new_G5214_ & ~new_G5224_;
  assign new_G5235_ = new_G5256_ | new_G5255_;
  assign new_G5236_ = G5202 | new_G5235_;
  assign new_G5237_ = new_G5260_ | new_G5259_;
  assign new_G5238_ = ~G5202 & new_G5237_;
  assign new_G5239_ = new_G5258_ | new_G5257_;
  assign new_G5240_ = G5202 & new_G5239_;
  assign new_G5241_ = G5200 & ~new_G5210_;
  assign new_G5242_ = ~G5200 & new_G5210_;
  assign new_G5243_ = ~G5199 | ~new_G5224_;
  assign new_G5244_ = new_G5210_ & new_G5243_;
  assign new_G5245_ = ~new_G5210_ & ~new_G5244_;
  assign new_G5246_ = new_G5210_ | new_G5243_;
  assign new_G5247_ = ~G5200 & G5201;
  assign new_G5248_ = G5200 & ~G5201;
  assign new_G5249_ = new_G5217_ | new_G5254_;
  assign new_G5250_ = ~new_G5217_ & ~new_G5253_;
  assign new_G5251_ = G5200 | new_G5217_;
  assign new_G5252_ = G5200 | G5201;
  assign new_G5253_ = new_G5217_ & new_G5254_;
  assign new_G5254_ = ~G5199 | ~new_G5224_;
  assign new_G5255_ = new_G5232_ & new_G5252_;
  assign new_G5256_ = ~new_G5232_ & ~new_G5252_;
  assign new_G5257_ = new_G5261_ | new_G5262_;
  assign new_G5258_ = ~G5203 & new_G5217_;
  assign new_G5259_ = new_G5263_ | new_G5264_;
  assign new_G5260_ = G5203 & new_G5217_;
  assign new_G5261_ = ~G5203 & ~new_G5217_;
  assign new_G5262_ = G5203 & ~new_G5217_;
  assign new_G5263_ = G5203 & ~new_G5217_;
  assign new_G5264_ = ~G5203 & new_G5217_;
  assign new_G5271_ = new_G5278_ & new_G5277_;
  assign new_G5272_ = new_G5280_ | new_G5279_;
  assign new_G5273_ = new_G5282_ | new_G5281_;
  assign new_G5274_ = new_G5284_ & new_G5283_;
  assign new_G5275_ = new_G5284_ & new_G5285_;
  assign new_G5276_ = new_G5277_ | new_G5286_;
  assign new_G5277_ = G5266 | new_G5289_;
  assign new_G5278_ = new_G5288_ | new_G5287_;
  assign new_G5279_ = new_G5293_ & new_G5292_;
  assign new_G5280_ = new_G5291_ & new_G5290_;
  assign new_G5281_ = new_G5296_ | new_G5295_;
  assign new_G5282_ = new_G5291_ & new_G5294_;
  assign new_G5283_ = G5266 | new_G5299_;
  assign new_G5284_ = new_G5298_ | new_G5297_;
  assign new_G5285_ = new_G5301_ | new_G5300_;
  assign new_G5286_ = ~new_G5277_ & new_G5303_;
  assign new_G5287_ = ~new_G5279_ & new_G5291_;
  assign new_G5288_ = new_G5279_ & ~new_G5291_;
  assign new_G5289_ = G5265 & ~G5266;
  assign new_G5290_ = ~new_G5312_ | ~new_G5313_;
  assign new_G5291_ = new_G5305_ | new_G5307_;
  assign new_G5292_ = new_G5315_ | new_G5314_;
  assign new_G5293_ = new_G5309_ | new_G5308_;
  assign new_G5294_ = ~new_G5317_ | ~new_G5316_;
  assign new_G5295_ = ~new_G5318_ & new_G5319_;
  assign new_G5296_ = new_G5318_ & ~new_G5319_;
  assign new_G5297_ = ~G5265 & G5266;
  assign new_G5298_ = G5265 & ~G5266;
  assign new_G5299_ = ~new_G5281_ | new_G5291_;
  assign new_G5300_ = new_G5281_ & new_G5291_;
  assign new_G5301_ = ~new_G5281_ & ~new_G5291_;
  assign new_G5302_ = new_G5323_ | new_G5322_;
  assign new_G5303_ = G5269 | new_G5302_;
  assign new_G5304_ = new_G5327_ | new_G5326_;
  assign new_G5305_ = ~G5269 & new_G5304_;
  assign new_G5306_ = new_G5325_ | new_G5324_;
  assign new_G5307_ = G5269 & new_G5306_;
  assign new_G5308_ = G5267 & ~new_G5277_;
  assign new_G5309_ = ~G5267 & new_G5277_;
  assign new_G5310_ = ~G5266 | ~new_G5291_;
  assign new_G5311_ = new_G5277_ & new_G5310_;
  assign new_G5312_ = ~new_G5277_ & ~new_G5311_;
  assign new_G5313_ = new_G5277_ | new_G5310_;
  assign new_G5314_ = ~G5267 & G5268;
  assign new_G5315_ = G5267 & ~G5268;
  assign new_G5316_ = new_G5284_ | new_G5321_;
  assign new_G5317_ = ~new_G5284_ & ~new_G5320_;
  assign new_G5318_ = G5267 | new_G5284_;
  assign new_G5319_ = G5267 | G5268;
  assign new_G5320_ = new_G5284_ & new_G5321_;
  assign new_G5321_ = ~G5266 | ~new_G5291_;
  assign new_G5322_ = new_G5299_ & new_G5319_;
  assign new_G5323_ = ~new_G5299_ & ~new_G5319_;
  assign new_G5324_ = new_G5328_ | new_G5329_;
  assign new_G5325_ = ~G5270 & new_G5284_;
  assign new_G5326_ = new_G5330_ | new_G5331_;
  assign new_G5327_ = G5270 & new_G5284_;
  assign new_G5328_ = ~G5270 & ~new_G5284_;
  assign new_G5329_ = G5270 & ~new_G5284_;
  assign new_G5330_ = G5270 & ~new_G5284_;
  assign new_G5331_ = ~G5270 & new_G5284_;
  assign new_G5338_ = new_G5345_ & new_G5344_;
  assign new_G5339_ = new_G5347_ | new_G5346_;
  assign new_G5340_ = new_G5349_ | new_G5348_;
  assign new_G5341_ = new_G5351_ & new_G5350_;
  assign new_G5342_ = new_G5351_ & new_G5352_;
  assign new_G5343_ = new_G5344_ | new_G5353_;
  assign new_G5344_ = G5333 | new_G5356_;
  assign new_G5345_ = new_G5355_ | new_G5354_;
  assign new_G5346_ = new_G5360_ & new_G5359_;
  assign new_G5347_ = new_G5358_ & new_G5357_;
  assign new_G5348_ = new_G5363_ | new_G5362_;
  assign new_G5349_ = new_G5358_ & new_G5361_;
  assign new_G5350_ = G5333 | new_G5366_;
  assign new_G5351_ = new_G5365_ | new_G5364_;
  assign new_G5352_ = new_G5368_ | new_G5367_;
  assign new_G5353_ = ~new_G5344_ & new_G5370_;
  assign new_G5354_ = ~new_G5346_ & new_G5358_;
  assign new_G5355_ = new_G5346_ & ~new_G5358_;
  assign new_G5356_ = G5332 & ~G5333;
  assign new_G5357_ = ~new_G5379_ | ~new_G5380_;
  assign new_G5358_ = new_G5372_ | new_G5374_;
  assign new_G5359_ = new_G5382_ | new_G5381_;
  assign new_G5360_ = new_G5376_ | new_G5375_;
  assign new_G5361_ = ~new_G5384_ | ~new_G5383_;
  assign new_G5362_ = ~new_G5385_ & new_G5386_;
  assign new_G5363_ = new_G5385_ & ~new_G5386_;
  assign new_G5364_ = ~G5332 & G5333;
  assign new_G5365_ = G5332 & ~G5333;
  assign new_G5366_ = ~new_G5348_ | new_G5358_;
  assign new_G5367_ = new_G5348_ & new_G5358_;
  assign new_G5368_ = ~new_G5348_ & ~new_G5358_;
  assign new_G5369_ = new_G5390_ | new_G5389_;
  assign new_G5370_ = G5336 | new_G5369_;
  assign new_G5371_ = new_G5394_ | new_G5393_;
  assign new_G5372_ = ~G5336 & new_G5371_;
  assign new_G5373_ = new_G5392_ | new_G5391_;
  assign new_G5374_ = G5336 & new_G5373_;
  assign new_G5375_ = G5334 & ~new_G5344_;
  assign new_G5376_ = ~G5334 & new_G5344_;
  assign new_G5377_ = ~G5333 | ~new_G5358_;
  assign new_G5378_ = new_G5344_ & new_G5377_;
  assign new_G5379_ = ~new_G5344_ & ~new_G5378_;
  assign new_G5380_ = new_G5344_ | new_G5377_;
  assign new_G5381_ = ~G5334 & G5335;
  assign new_G5382_ = G5334 & ~G5335;
  assign new_G5383_ = new_G5351_ | new_G5388_;
  assign new_G5384_ = ~new_G5351_ & ~new_G5387_;
  assign new_G5385_ = G5334 | new_G5351_;
  assign new_G5386_ = G5334 | G5335;
  assign new_G5387_ = new_G5351_ & new_G5388_;
  assign new_G5388_ = ~G5333 | ~new_G5358_;
  assign new_G5389_ = new_G5366_ & new_G5386_;
  assign new_G5390_ = ~new_G5366_ & ~new_G5386_;
  assign new_G5391_ = new_G5395_ | new_G5396_;
  assign new_G5392_ = ~G5337 & new_G5351_;
  assign new_G5393_ = new_G5397_ | new_G5398_;
  assign new_G5394_ = G5337 & new_G5351_;
  assign new_G5395_ = ~G5337 & ~new_G5351_;
  assign new_G5396_ = G5337 & ~new_G5351_;
  assign new_G5397_ = G5337 & ~new_G5351_;
  assign new_G5398_ = ~G5337 & new_G5351_;
  assign new_G5405_ = new_G5412_ & new_G5411_;
  assign new_G5406_ = new_G5414_ | new_G5413_;
  assign new_G5407_ = new_G5416_ | new_G5415_;
  assign new_G5408_ = new_G5418_ & new_G5417_;
  assign new_G5409_ = new_G5418_ & new_G5419_;
  assign new_G5410_ = new_G5411_ | new_G5420_;
  assign new_G5411_ = G5400 | new_G5423_;
  assign new_G5412_ = new_G5422_ | new_G5421_;
  assign new_G5413_ = new_G5427_ & new_G5426_;
  assign new_G5414_ = new_G5425_ & new_G5424_;
  assign new_G5415_ = new_G5430_ | new_G5429_;
  assign new_G5416_ = new_G5425_ & new_G5428_;
  assign new_G5417_ = G5400 | new_G5433_;
  assign new_G5418_ = new_G5432_ | new_G5431_;
  assign new_G5419_ = new_G5435_ | new_G5434_;
  assign new_G5420_ = ~new_G5411_ & new_G5437_;
  assign new_G5421_ = ~new_G5413_ & new_G5425_;
  assign new_G5422_ = new_G5413_ & ~new_G5425_;
  assign new_G5423_ = G5399 & ~G5400;
  assign new_G5424_ = ~new_G5446_ | ~new_G5447_;
  assign new_G5425_ = new_G5439_ | new_G5441_;
  assign new_G5426_ = new_G5449_ | new_G5448_;
  assign new_G5427_ = new_G5443_ | new_G5442_;
  assign new_G5428_ = ~new_G5451_ | ~new_G5450_;
  assign new_G5429_ = ~new_G5452_ & new_G5453_;
  assign new_G5430_ = new_G5452_ & ~new_G5453_;
  assign new_G5431_ = ~G5399 & G5400;
  assign new_G5432_ = G5399 & ~G5400;
  assign new_G5433_ = ~new_G5415_ | new_G5425_;
  assign new_G5434_ = new_G5415_ & new_G5425_;
  assign new_G5435_ = ~new_G5415_ & ~new_G5425_;
  assign new_G5436_ = new_G5457_ | new_G5456_;
  assign new_G5437_ = G5403 | new_G5436_;
  assign new_G5438_ = new_G5461_ | new_G5460_;
  assign new_G5439_ = ~G5403 & new_G5438_;
  assign new_G5440_ = new_G5459_ | new_G5458_;
  assign new_G5441_ = G5403 & new_G5440_;
  assign new_G5442_ = G5401 & ~new_G5411_;
  assign new_G5443_ = ~G5401 & new_G5411_;
  assign new_G5444_ = ~G5400 | ~new_G5425_;
  assign new_G5445_ = new_G5411_ & new_G5444_;
  assign new_G5446_ = ~new_G5411_ & ~new_G5445_;
  assign new_G5447_ = new_G5411_ | new_G5444_;
  assign new_G5448_ = ~G5401 & G5402;
  assign new_G5449_ = G5401 & ~G5402;
  assign new_G5450_ = new_G5418_ | new_G5455_;
  assign new_G5451_ = ~new_G5418_ & ~new_G5454_;
  assign new_G5452_ = G5401 | new_G5418_;
  assign new_G5453_ = G5401 | G5402;
  assign new_G5454_ = new_G5418_ & new_G5455_;
  assign new_G5455_ = ~G5400 | ~new_G5425_;
  assign new_G5456_ = new_G5433_ & new_G5453_;
  assign new_G5457_ = ~new_G5433_ & ~new_G5453_;
  assign new_G5458_ = new_G5462_ | new_G5463_;
  assign new_G5459_ = ~G5404 & new_G5418_;
  assign new_G5460_ = new_G5464_ | new_G5465_;
  assign new_G5461_ = G5404 & new_G5418_;
  assign new_G5462_ = ~G5404 & ~new_G5418_;
  assign new_G5463_ = G5404 & ~new_G5418_;
  assign new_G5464_ = G5404 & ~new_G5418_;
  assign new_G5465_ = ~G5404 & new_G5418_;
  assign new_G5472_ = new_G5479_ & new_G5478_;
  assign new_G5473_ = new_G5481_ | new_G5480_;
  assign new_G5474_ = new_G5483_ | new_G5482_;
  assign new_G5475_ = new_G5485_ & new_G5484_;
  assign new_G5476_ = new_G5485_ & new_G5486_;
  assign new_G5477_ = new_G5478_ | new_G5487_;
  assign new_G5478_ = G5467 | new_G5490_;
  assign new_G5479_ = new_G5489_ | new_G5488_;
  assign new_G5480_ = new_G5494_ & new_G5493_;
  assign new_G5481_ = new_G5492_ & new_G5491_;
  assign new_G5482_ = new_G5497_ | new_G5496_;
  assign new_G5483_ = new_G5492_ & new_G5495_;
  assign new_G5484_ = G5467 | new_G5500_;
  assign new_G5485_ = new_G5499_ | new_G5498_;
  assign new_G5486_ = new_G5502_ | new_G5501_;
  assign new_G5487_ = ~new_G5478_ & new_G5504_;
  assign new_G5488_ = ~new_G5480_ & new_G5492_;
  assign new_G5489_ = new_G5480_ & ~new_G5492_;
  assign new_G5490_ = G5466 & ~G5467;
  assign new_G5491_ = ~new_G5513_ | ~new_G5514_;
  assign new_G5492_ = new_G5506_ | new_G5508_;
  assign new_G5493_ = new_G5516_ | new_G5515_;
  assign new_G5494_ = new_G5510_ | new_G5509_;
  assign new_G5495_ = ~new_G5518_ | ~new_G5517_;
  assign new_G5496_ = ~new_G5519_ & new_G5520_;
  assign new_G5497_ = new_G5519_ & ~new_G5520_;
  assign new_G5498_ = ~G5466 & G5467;
  assign new_G5499_ = G5466 & ~G5467;
  assign new_G5500_ = ~new_G5482_ | new_G5492_;
  assign new_G5501_ = new_G5482_ & new_G5492_;
  assign new_G5502_ = ~new_G5482_ & ~new_G5492_;
  assign new_G5503_ = new_G5524_ | new_G5523_;
  assign new_G5504_ = G5470 | new_G5503_;
  assign new_G5505_ = new_G5528_ | new_G5527_;
  assign new_G5506_ = ~G5470 & new_G5505_;
  assign new_G5507_ = new_G5526_ | new_G5525_;
  assign new_G5508_ = G5470 & new_G5507_;
  assign new_G5509_ = G5468 & ~new_G5478_;
  assign new_G5510_ = ~G5468 & new_G5478_;
  assign new_G5511_ = ~G5467 | ~new_G5492_;
  assign new_G5512_ = new_G5478_ & new_G5511_;
  assign new_G5513_ = ~new_G5478_ & ~new_G5512_;
  assign new_G5514_ = new_G5478_ | new_G5511_;
  assign new_G5515_ = ~G5468 & G5469;
  assign new_G5516_ = G5468 & ~G5469;
  assign new_G5517_ = new_G5485_ | new_G5522_;
  assign new_G5518_ = ~new_G5485_ & ~new_G5521_;
  assign new_G5519_ = G5468 | new_G5485_;
  assign new_G5520_ = G5468 | G5469;
  assign new_G5521_ = new_G5485_ & new_G5522_;
  assign new_G5522_ = ~G5467 | ~new_G5492_;
  assign new_G5523_ = new_G5500_ & new_G5520_;
  assign new_G5524_ = ~new_G5500_ & ~new_G5520_;
  assign new_G5525_ = new_G5529_ | new_G5530_;
  assign new_G5526_ = ~G5471 & new_G5485_;
  assign new_G5527_ = new_G5531_ | new_G5532_;
  assign new_G5528_ = G5471 & new_G5485_;
  assign new_G5529_ = ~G5471 & ~new_G5485_;
  assign new_G5530_ = G5471 & ~new_G5485_;
  assign new_G5531_ = G5471 & ~new_G5485_;
  assign new_G5532_ = ~G5471 & new_G5485_;
  assign new_G5539_ = new_G5546_ & new_G5545_;
  assign new_G5540_ = new_G5548_ | new_G5547_;
  assign new_G5541_ = new_G5550_ | new_G5549_;
  assign new_G5542_ = new_G5552_ & new_G5551_;
  assign new_G5543_ = new_G5552_ & new_G5553_;
  assign new_G5544_ = new_G5545_ | new_G5554_;
  assign new_G5545_ = G5534 | new_G5557_;
  assign new_G5546_ = new_G5556_ | new_G5555_;
  assign new_G5547_ = new_G5561_ & new_G5560_;
  assign new_G5548_ = new_G5559_ & new_G5558_;
  assign new_G5549_ = new_G5564_ | new_G5563_;
  assign new_G5550_ = new_G5559_ & new_G5562_;
  assign new_G5551_ = G5534 | new_G5567_;
  assign new_G5552_ = new_G5566_ | new_G5565_;
  assign new_G5553_ = new_G5569_ | new_G5568_;
  assign new_G5554_ = ~new_G5545_ & new_G5571_;
  assign new_G5555_ = ~new_G5547_ & new_G5559_;
  assign new_G5556_ = new_G5547_ & ~new_G5559_;
  assign new_G5557_ = G5533 & ~G5534;
  assign new_G5558_ = ~new_G5580_ | ~new_G5581_;
  assign new_G5559_ = new_G5573_ | new_G5575_;
  assign new_G5560_ = new_G5583_ | new_G5582_;
  assign new_G5561_ = new_G5577_ | new_G5576_;
  assign new_G5562_ = ~new_G5585_ | ~new_G5584_;
  assign new_G5563_ = ~new_G5586_ & new_G5587_;
  assign new_G5564_ = new_G5586_ & ~new_G5587_;
  assign new_G5565_ = ~G5533 & G5534;
  assign new_G5566_ = G5533 & ~G5534;
  assign new_G5567_ = ~new_G5549_ | new_G5559_;
  assign new_G5568_ = new_G5549_ & new_G5559_;
  assign new_G5569_ = ~new_G5549_ & ~new_G5559_;
  assign new_G5570_ = new_G5591_ | new_G5590_;
  assign new_G5571_ = G5537 | new_G5570_;
  assign new_G5572_ = new_G5595_ | new_G5594_;
  assign new_G5573_ = ~G5537 & new_G5572_;
  assign new_G5574_ = new_G5593_ | new_G5592_;
  assign new_G5575_ = G5537 & new_G5574_;
  assign new_G5576_ = G5535 & ~new_G5545_;
  assign new_G5577_ = ~G5535 & new_G5545_;
  assign new_G5578_ = ~G5534 | ~new_G5559_;
  assign new_G5579_ = new_G5545_ & new_G5578_;
  assign new_G5580_ = ~new_G5545_ & ~new_G5579_;
  assign new_G5581_ = new_G5545_ | new_G5578_;
  assign new_G5582_ = ~G5535 & G5536;
  assign new_G5583_ = G5535 & ~G5536;
  assign new_G5584_ = new_G5552_ | new_G5589_;
  assign new_G5585_ = ~new_G5552_ & ~new_G5588_;
  assign new_G5586_ = G5535 | new_G5552_;
  assign new_G5587_ = G5535 | G5536;
  assign new_G5588_ = new_G5552_ & new_G5589_;
  assign new_G5589_ = ~G5534 | ~new_G5559_;
  assign new_G5590_ = new_G5567_ & new_G5587_;
  assign new_G5591_ = ~new_G5567_ & ~new_G5587_;
  assign new_G5592_ = new_G5596_ | new_G5597_;
  assign new_G5593_ = ~G5538 & new_G5552_;
  assign new_G5594_ = new_G5598_ | new_G5599_;
  assign new_G5595_ = G5538 & new_G5552_;
  assign new_G5596_ = ~G5538 & ~new_G5552_;
  assign new_G5597_ = G5538 & ~new_G5552_;
  assign new_G5598_ = G5538 & ~new_G5552_;
  assign new_G5599_ = ~G5538 & new_G5552_;
  assign new_G5606_ = new_G5613_ & new_G5612_;
  assign new_G5607_ = new_G5615_ | new_G5614_;
  assign new_G5608_ = new_G5617_ | new_G5616_;
  assign new_G5609_ = new_G5619_ & new_G5618_;
  assign new_G5610_ = new_G5619_ & new_G5620_;
  assign new_G5611_ = new_G5612_ | new_G5621_;
  assign new_G5612_ = G5601 | new_G5624_;
  assign new_G5613_ = new_G5623_ | new_G5622_;
  assign new_G5614_ = new_G5628_ & new_G5627_;
  assign new_G5615_ = new_G5626_ & new_G5625_;
  assign new_G5616_ = new_G5631_ | new_G5630_;
  assign new_G5617_ = new_G5626_ & new_G5629_;
  assign new_G5618_ = G5601 | new_G5634_;
  assign new_G5619_ = new_G5633_ | new_G5632_;
  assign new_G5620_ = new_G5636_ | new_G5635_;
  assign new_G5621_ = ~new_G5612_ & new_G5638_;
  assign new_G5622_ = ~new_G5614_ & new_G5626_;
  assign new_G5623_ = new_G5614_ & ~new_G5626_;
  assign new_G5624_ = G5600 & ~G5601;
  assign new_G5625_ = ~new_G5647_ | ~new_G5648_;
  assign new_G5626_ = new_G5640_ | new_G5642_;
  assign new_G5627_ = new_G5650_ | new_G5649_;
  assign new_G5628_ = new_G5644_ | new_G5643_;
  assign new_G5629_ = ~new_G5652_ | ~new_G5651_;
  assign new_G5630_ = ~new_G5653_ & new_G5654_;
  assign new_G5631_ = new_G5653_ & ~new_G5654_;
  assign new_G5632_ = ~G5600 & G5601;
  assign new_G5633_ = G5600 & ~G5601;
  assign new_G5634_ = ~new_G5616_ | new_G5626_;
  assign new_G5635_ = new_G5616_ & new_G5626_;
  assign new_G5636_ = ~new_G5616_ & ~new_G5626_;
  assign new_G5637_ = new_G5658_ | new_G5657_;
  assign new_G5638_ = G5604 | new_G5637_;
  assign new_G5639_ = new_G5662_ | new_G5661_;
  assign new_G5640_ = ~G5604 & new_G5639_;
  assign new_G5641_ = new_G5660_ | new_G5659_;
  assign new_G5642_ = G5604 & new_G5641_;
  assign new_G5643_ = G5602 & ~new_G5612_;
  assign new_G5644_ = ~G5602 & new_G5612_;
  assign new_G5645_ = ~G5601 | ~new_G5626_;
  assign new_G5646_ = new_G5612_ & new_G5645_;
  assign new_G5647_ = ~new_G5612_ & ~new_G5646_;
  assign new_G5648_ = new_G5612_ | new_G5645_;
  assign new_G5649_ = ~G5602 & G5603;
  assign new_G5650_ = G5602 & ~G5603;
  assign new_G5651_ = new_G5619_ | new_G5656_;
  assign new_G5652_ = ~new_G5619_ & ~new_G5655_;
  assign new_G5653_ = G5602 | new_G5619_;
  assign new_G5654_ = G5602 | G5603;
  assign new_G5655_ = new_G5619_ & new_G5656_;
  assign new_G5656_ = ~G5601 | ~new_G5626_;
  assign new_G5657_ = new_G5634_ & new_G5654_;
  assign new_G5658_ = ~new_G5634_ & ~new_G5654_;
  assign new_G5659_ = new_G5663_ | new_G5664_;
  assign new_G5660_ = ~G5605 & new_G5619_;
  assign new_G5661_ = new_G5665_ | new_G5666_;
  assign new_G5662_ = G5605 & new_G5619_;
  assign new_G5663_ = ~G5605 & ~new_G5619_;
  assign new_G5664_ = G5605 & ~new_G5619_;
  assign new_G5665_ = G5605 & ~new_G5619_;
  assign new_G5666_ = ~G5605 & new_G5619_;
  assign new_G5673_ = new_G5680_ & new_G5679_;
  assign new_G5674_ = new_G5682_ | new_G5681_;
  assign new_G5675_ = new_G5684_ | new_G5683_;
  assign new_G5676_ = new_G5686_ & new_G5685_;
  assign new_G5677_ = new_G5686_ & new_G5687_;
  assign new_G5678_ = new_G5679_ | new_G5688_;
  assign new_G5679_ = G5668 | new_G5691_;
  assign new_G5680_ = new_G5690_ | new_G5689_;
  assign new_G5681_ = new_G5695_ & new_G5694_;
  assign new_G5682_ = new_G5693_ & new_G5692_;
  assign new_G5683_ = new_G5698_ | new_G5697_;
  assign new_G5684_ = new_G5693_ & new_G5696_;
  assign new_G5685_ = G5668 | new_G5701_;
  assign new_G5686_ = new_G5700_ | new_G5699_;
  assign new_G5687_ = new_G5703_ | new_G5702_;
  assign new_G5688_ = ~new_G5679_ & new_G5705_;
  assign new_G5689_ = ~new_G5681_ & new_G5693_;
  assign new_G5690_ = new_G5681_ & ~new_G5693_;
  assign new_G5691_ = G5667 & ~G5668;
  assign new_G5692_ = ~new_G5714_ | ~new_G5715_;
  assign new_G5693_ = new_G5707_ | new_G5709_;
  assign new_G5694_ = new_G5717_ | new_G5716_;
  assign new_G5695_ = new_G5711_ | new_G5710_;
  assign new_G5696_ = ~new_G5719_ | ~new_G5718_;
  assign new_G5697_ = ~new_G5720_ & new_G5721_;
  assign new_G5698_ = new_G5720_ & ~new_G5721_;
  assign new_G5699_ = ~G5667 & G5668;
  assign new_G5700_ = G5667 & ~G5668;
  assign new_G5701_ = ~new_G5683_ | new_G5693_;
  assign new_G5702_ = new_G5683_ & new_G5693_;
  assign new_G5703_ = ~new_G5683_ & ~new_G5693_;
  assign new_G5704_ = new_G5725_ | new_G5724_;
  assign new_G5705_ = G5671 | new_G5704_;
  assign new_G5706_ = new_G5729_ | new_G5728_;
  assign new_G5707_ = ~G5671 & new_G5706_;
  assign new_G5708_ = new_G5727_ | new_G5726_;
  assign new_G5709_ = G5671 & new_G5708_;
  assign new_G5710_ = G5669 & ~new_G5679_;
  assign new_G5711_ = ~G5669 & new_G5679_;
  assign new_G5712_ = ~G5668 | ~new_G5693_;
  assign new_G5713_ = new_G5679_ & new_G5712_;
  assign new_G5714_ = ~new_G5679_ & ~new_G5713_;
  assign new_G5715_ = new_G5679_ | new_G5712_;
  assign new_G5716_ = ~G5669 & G5670;
  assign new_G5717_ = G5669 & ~G5670;
  assign new_G5718_ = new_G5686_ | new_G5723_;
  assign new_G5719_ = ~new_G5686_ & ~new_G5722_;
  assign new_G5720_ = G5669 | new_G5686_;
  assign new_G5721_ = G5669 | G5670;
  assign new_G5722_ = new_G5686_ & new_G5723_;
  assign new_G5723_ = ~G5668 | ~new_G5693_;
  assign new_G5724_ = new_G5701_ & new_G5721_;
  assign new_G5725_ = ~new_G5701_ & ~new_G5721_;
  assign new_G5726_ = new_G5730_ | new_G5731_;
  assign new_G5727_ = ~G5672 & new_G5686_;
  assign new_G5728_ = new_G5732_ | new_G5733_;
  assign new_G5729_ = G5672 & new_G5686_;
  assign new_G5730_ = ~G5672 & ~new_G5686_;
  assign new_G5731_ = G5672 & ~new_G5686_;
  assign new_G5732_ = G5672 & ~new_G5686_;
  assign new_G5733_ = ~G5672 & new_G5686_;
  assign new_G5740_ = new_G5747_ & new_G5746_;
  assign new_G5741_ = new_G5749_ | new_G5748_;
  assign new_G5742_ = new_G5751_ | new_G5750_;
  assign new_G5743_ = new_G5753_ & new_G5752_;
  assign new_G5744_ = new_G5753_ & new_G5754_;
  assign new_G5745_ = new_G5746_ | new_G5755_;
  assign new_G5746_ = G5735 | new_G5758_;
  assign new_G5747_ = new_G5757_ | new_G5756_;
  assign new_G5748_ = new_G5762_ & new_G5761_;
  assign new_G5749_ = new_G5760_ & new_G5759_;
  assign new_G5750_ = new_G5765_ | new_G5764_;
  assign new_G5751_ = new_G5760_ & new_G5763_;
  assign new_G5752_ = G5735 | new_G5768_;
  assign new_G5753_ = new_G5767_ | new_G5766_;
  assign new_G5754_ = new_G5770_ | new_G5769_;
  assign new_G5755_ = ~new_G5746_ & new_G5772_;
  assign new_G5756_ = ~new_G5748_ & new_G5760_;
  assign new_G5757_ = new_G5748_ & ~new_G5760_;
  assign new_G5758_ = G5734 & ~G5735;
  assign new_G5759_ = ~new_G5781_ | ~new_G5782_;
  assign new_G5760_ = new_G5774_ | new_G5776_;
  assign new_G5761_ = new_G5784_ | new_G5783_;
  assign new_G5762_ = new_G5778_ | new_G5777_;
  assign new_G5763_ = ~new_G5786_ | ~new_G5785_;
  assign new_G5764_ = ~new_G5787_ & new_G5788_;
  assign new_G5765_ = new_G5787_ & ~new_G5788_;
  assign new_G5766_ = ~G5734 & G5735;
  assign new_G5767_ = G5734 & ~G5735;
  assign new_G5768_ = ~new_G5750_ | new_G5760_;
  assign new_G5769_ = new_G5750_ & new_G5760_;
  assign new_G5770_ = ~new_G5750_ & ~new_G5760_;
  assign new_G5771_ = new_G5792_ | new_G5791_;
  assign new_G5772_ = G5738 | new_G5771_;
  assign new_G5773_ = new_G5796_ | new_G5795_;
  assign new_G5774_ = ~G5738 & new_G5773_;
  assign new_G5775_ = new_G5794_ | new_G5793_;
  assign new_G5776_ = G5738 & new_G5775_;
  assign new_G5777_ = G5736 & ~new_G5746_;
  assign new_G5778_ = ~G5736 & new_G5746_;
  assign new_G5779_ = ~G5735 | ~new_G5760_;
  assign new_G5780_ = new_G5746_ & new_G5779_;
  assign new_G5781_ = ~new_G5746_ & ~new_G5780_;
  assign new_G5782_ = new_G5746_ | new_G5779_;
  assign new_G5783_ = ~G5736 & G5737;
  assign new_G5784_ = G5736 & ~G5737;
  assign new_G5785_ = new_G5753_ | new_G5790_;
  assign new_G5786_ = ~new_G5753_ & ~new_G5789_;
  assign new_G5787_ = G5736 | new_G5753_;
  assign new_G5788_ = G5736 | G5737;
  assign new_G5789_ = new_G5753_ & new_G5790_;
  assign new_G5790_ = ~G5735 | ~new_G5760_;
  assign new_G5791_ = new_G5768_ & new_G5788_;
  assign new_G5792_ = ~new_G5768_ & ~new_G5788_;
  assign new_G5793_ = new_G5797_ | new_G5798_;
  assign new_G5794_ = ~G5739 & new_G5753_;
  assign new_G5795_ = new_G5799_ | new_G5800_;
  assign new_G5796_ = G5739 & new_G5753_;
  assign new_G5797_ = ~G5739 & ~new_G5753_;
  assign new_G5798_ = G5739 & ~new_G5753_;
  assign new_G5799_ = G5739 & ~new_G5753_;
  assign new_G5800_ = ~G5739 & new_G5753_;
  assign new_G5807_ = new_G5814_ & new_G5813_;
  assign new_G5808_ = new_G5816_ | new_G5815_;
  assign new_G5809_ = new_G5818_ | new_G5817_;
  assign new_G5810_ = new_G5820_ & new_G5819_;
  assign new_G5811_ = new_G5820_ & new_G5821_;
  assign new_G5812_ = new_G5813_ | new_G5822_;
  assign new_G5813_ = G5802 | new_G5825_;
  assign new_G5814_ = new_G5824_ | new_G5823_;
  assign new_G5815_ = new_G5829_ & new_G5828_;
  assign new_G5816_ = new_G5827_ & new_G5826_;
  assign new_G5817_ = new_G5832_ | new_G5831_;
  assign new_G5818_ = new_G5827_ & new_G5830_;
  assign new_G5819_ = G5802 | new_G5835_;
  assign new_G5820_ = new_G5834_ | new_G5833_;
  assign new_G5821_ = new_G5837_ | new_G5836_;
  assign new_G5822_ = ~new_G5813_ & new_G5839_;
  assign new_G5823_ = ~new_G5815_ & new_G5827_;
  assign new_G5824_ = new_G5815_ & ~new_G5827_;
  assign new_G5825_ = G5801 & ~G5802;
  assign new_G5826_ = ~new_G5848_ | ~new_G5849_;
  assign new_G5827_ = new_G5841_ | new_G5843_;
  assign new_G5828_ = new_G5851_ | new_G5850_;
  assign new_G5829_ = new_G5845_ | new_G5844_;
  assign new_G5830_ = ~new_G5853_ | ~new_G5852_;
  assign new_G5831_ = ~new_G5854_ & new_G5855_;
  assign new_G5832_ = new_G5854_ & ~new_G5855_;
  assign new_G5833_ = ~G5801 & G5802;
  assign new_G5834_ = G5801 & ~G5802;
  assign new_G5835_ = ~new_G5817_ | new_G5827_;
  assign new_G5836_ = new_G5817_ & new_G5827_;
  assign new_G5837_ = ~new_G5817_ & ~new_G5827_;
  assign new_G5838_ = new_G5859_ | new_G5858_;
  assign new_G5839_ = G5805 | new_G5838_;
  assign new_G5840_ = new_G5863_ | new_G5862_;
  assign new_G5841_ = ~G5805 & new_G5840_;
  assign new_G5842_ = new_G5861_ | new_G5860_;
  assign new_G5843_ = G5805 & new_G5842_;
  assign new_G5844_ = G5803 & ~new_G5813_;
  assign new_G5845_ = ~G5803 & new_G5813_;
  assign new_G5846_ = ~G5802 | ~new_G5827_;
  assign new_G5847_ = new_G5813_ & new_G5846_;
  assign new_G5848_ = ~new_G5813_ & ~new_G5847_;
  assign new_G5849_ = new_G5813_ | new_G5846_;
  assign new_G5850_ = ~G5803 & G5804;
  assign new_G5851_ = G5803 & ~G5804;
  assign new_G5852_ = new_G5820_ | new_G5857_;
  assign new_G5853_ = ~new_G5820_ & ~new_G5856_;
  assign new_G5854_ = G5803 | new_G5820_;
  assign new_G5855_ = G5803 | G5804;
  assign new_G5856_ = new_G5820_ & new_G5857_;
  assign new_G5857_ = ~G5802 | ~new_G5827_;
  assign new_G5858_ = new_G5835_ & new_G5855_;
  assign new_G5859_ = ~new_G5835_ & ~new_G5855_;
  assign new_G5860_ = new_G5864_ | new_G5865_;
  assign new_G5861_ = ~G5806 & new_G5820_;
  assign new_G5862_ = new_G5866_ | new_G5867_;
  assign new_G5863_ = G5806 & new_G5820_;
  assign new_G5864_ = ~G5806 & ~new_G5820_;
  assign new_G5865_ = G5806 & ~new_G5820_;
  assign new_G5866_ = G5806 & ~new_G5820_;
  assign new_G5867_ = ~G5806 & new_G5820_;
  assign new_G5874_ = new_G5881_ & new_G5880_;
  assign new_G5875_ = new_G5883_ | new_G5882_;
  assign new_G5876_ = new_G5885_ | new_G5884_;
  assign new_G5877_ = new_G5887_ & new_G5886_;
  assign new_G5878_ = new_G5887_ & new_G5888_;
  assign new_G5879_ = new_G5880_ | new_G5889_;
  assign new_G5880_ = G5869 | new_G5892_;
  assign new_G5881_ = new_G5891_ | new_G5890_;
  assign new_G5882_ = new_G5896_ & new_G5895_;
  assign new_G5883_ = new_G5894_ & new_G5893_;
  assign new_G5884_ = new_G5899_ | new_G5898_;
  assign new_G5885_ = new_G5894_ & new_G5897_;
  assign new_G5886_ = G5869 | new_G5902_;
  assign new_G5887_ = new_G5901_ | new_G5900_;
  assign new_G5888_ = new_G5904_ | new_G5903_;
  assign new_G5889_ = ~new_G5880_ & new_G5906_;
  assign new_G5890_ = ~new_G5882_ & new_G5894_;
  assign new_G5891_ = new_G5882_ & ~new_G5894_;
  assign new_G5892_ = G5868 & ~G5869;
  assign new_G5893_ = ~new_G5915_ | ~new_G5916_;
  assign new_G5894_ = new_G5908_ | new_G5910_;
  assign new_G5895_ = new_G5918_ | new_G5917_;
  assign new_G5896_ = new_G5912_ | new_G5911_;
  assign new_G5897_ = ~new_G5920_ | ~new_G5919_;
  assign new_G5898_ = ~new_G5921_ & new_G5922_;
  assign new_G5899_ = new_G5921_ & ~new_G5922_;
  assign new_G5900_ = ~G5868 & G5869;
  assign new_G5901_ = G5868 & ~G5869;
  assign new_G5902_ = ~new_G5884_ | new_G5894_;
  assign new_G5903_ = new_G5884_ & new_G5894_;
  assign new_G5904_ = ~new_G5884_ & ~new_G5894_;
  assign new_G5905_ = new_G5926_ | new_G5925_;
  assign new_G5906_ = G5872 | new_G5905_;
  assign new_G5907_ = new_G5930_ | new_G5929_;
  assign new_G5908_ = ~G5872 & new_G5907_;
  assign new_G5909_ = new_G5928_ | new_G5927_;
  assign new_G5910_ = G5872 & new_G5909_;
  assign new_G5911_ = G5870 & ~new_G5880_;
  assign new_G5912_ = ~G5870 & new_G5880_;
  assign new_G5913_ = ~G5869 | ~new_G5894_;
  assign new_G5914_ = new_G5880_ & new_G5913_;
  assign new_G5915_ = ~new_G5880_ & ~new_G5914_;
  assign new_G5916_ = new_G5880_ | new_G5913_;
  assign new_G5917_ = ~G5870 & G5871;
  assign new_G5918_ = G5870 & ~G5871;
  assign new_G5919_ = new_G5887_ | new_G5924_;
  assign new_G5920_ = ~new_G5887_ & ~new_G5923_;
  assign new_G5921_ = G5870 | new_G5887_;
  assign new_G5922_ = G5870 | G5871;
  assign new_G5923_ = new_G5887_ & new_G5924_;
  assign new_G5924_ = ~G5869 | ~new_G5894_;
  assign new_G5925_ = new_G5902_ & new_G5922_;
  assign new_G5926_ = ~new_G5902_ & ~new_G5922_;
  assign new_G5927_ = new_G5931_ | new_G5932_;
  assign new_G5928_ = ~G5873 & new_G5887_;
  assign new_G5929_ = new_G5933_ | new_G5934_;
  assign new_G5930_ = G5873 & new_G5887_;
  assign new_G5931_ = ~G5873 & ~new_G5887_;
  assign new_G5932_ = G5873 & ~new_G5887_;
  assign new_G5933_ = G5873 & ~new_G5887_;
  assign new_G5934_ = ~G5873 & new_G5887_;
  assign new_D7054_ = ~new_D6993_ & new_D7007_;
  assign new_D7053_ = new_D6993_ & ~new_D7007_;
  assign new_D7052_ = new_D6993_ & ~new_D7007_;
  assign new_D7051_ = ~new_D6993_ & ~new_D7007_;
  assign new_D7050_ = new_D6993_ & new_D7007_;
  assign new_D7049_ = new_D7053_ | new_D7054_;
  assign new_D7048_ = ~new_D6993_ & new_D7007_;
  assign new_D7047_ = new_D7051_ | new_D7052_;
  assign new_D7046_ = ~new_D7022_ & ~new_D7042_;
  assign new_D7045_ = new_D7022_ & new_D7042_;
  assign new_D7044_ = ~new_D6989_ | ~new_D7014_;
  assign new_D7043_ = new_D7007_ & new_D7044_;
  assign new_D7042_ = new_D6990_ | new_D6991_;
  assign new_D7041_ = new_D6990_ | new_D7007_;
  assign new_D7040_ = ~new_D7007_ & ~new_D7043_;
  assign new_D7039_ = new_D7007_ | new_D7044_;
  assign new_D7038_ = new_D6990_ & ~new_D6991_;
  assign new_D7037_ = ~new_D6990_ & new_D6991_;
  assign new_D7036_ = new_D7000_ | new_D7033_;
  assign new_D7035_ = ~new_D7000_ & ~new_D7034_;
  assign new_D7034_ = new_D7000_ & new_D7033_;
  assign new_D7033_ = ~new_D6989_ | ~new_D7014_;
  assign new_D7032_ = ~new_D6990_ & new_D7000_;
  assign new_D7031_ = new_D6990_ & ~new_D7000_;
  assign new_D7030_ = new_D6992_ & new_D7029_;
  assign new_D7029_ = new_D7048_ | new_D7047_;
  assign new_D7028_ = ~new_D6992_ & new_D7027_;
  assign new_D7027_ = new_D7050_ | new_D7049_;
  assign new_D7026_ = new_D6992_ | new_D7025_;
  assign new_D7025_ = new_D7046_ | new_D7045_;
  assign new_D7024_ = ~new_D7004_ & ~new_D7014_;
  assign new_D7023_ = new_D7004_ & new_D7014_;
  assign new_D7022_ = ~new_D7004_ | new_D7014_;
  assign new_D7021_ = new_D6988_ & ~new_D6989_;
  assign new_D7020_ = ~new_D6988_ & new_D6989_;
  assign new_D7019_ = new_D7041_ & ~new_D7042_;
  assign new_D7018_ = ~new_D7041_ & new_D7042_;
  assign new_D7017_ = ~new_D7040_ | ~new_D7039_;
  assign new_D7016_ = new_D7032_ | new_D7031_;
  assign new_D7015_ = new_D7038_ | new_D7037_;
  assign new_D7014_ = new_D7028_ | new_D7030_;
  assign new_D7013_ = ~new_D7035_ | ~new_D7036_;
  assign new_D7012_ = new_D6988_ & ~new_D6989_;
  assign new_D7011_ = new_D7002_ & ~new_D7014_;
  assign new_D7010_ = ~new_D7002_ & new_D7014_;
  assign new_D7009_ = ~new_D7000_ & new_D7026_;
  assign new_D7008_ = new_D7024_ | new_D7023_;
  assign new_D7007_ = new_D7021_ | new_D7020_;
  assign new_D7006_ = new_D6989_ | new_D7022_;
  assign new_D7005_ = new_D7014_ & new_D7017_;
  assign new_D7004_ = new_D7019_ | new_D7018_;
  assign new_D7003_ = new_D7014_ & new_D7013_;
  assign new_D7002_ = new_D7016_ & new_D7015_;
  assign new_D7001_ = new_D7011_ | new_D7010_;
  assign new_D7000_ = new_D6989_ | new_D7012_;
  assign new_D6999_ = new_D7000_ | new_D7009_;
  assign new_D6998_ = new_D7007_ & new_D7008_;
  assign new_D6997_ = new_D7007_ & new_D7006_;
  assign new_D6996_ = new_D7005_ | new_D7004_;
  assign new_D6995_ = new_D7003_ | new_D7002_;
  assign new_D6994_ = new_D7001_ & new_D7000_;
  assign new_D6993_ = new_F1473_;
  assign new_D6992_ = new_F1535_;
  assign new_D6991_ = new_F1602_;
  assign new_D6990_ = new_F1669_;
  assign new_D6989_ = new_F1736_;
  assign new_D6988_ = new_F1803_;
  assign new_D7055_ = new_F1870_;
  assign new_D7056_ = new_F1937_;
  assign new_D7057_ = new_F2004_;
  assign new_D7058_ = new_F2071_;
  assign new_D7059_ = new_F2138_;
  assign new_D7060_ = new_F2205_;
  assign new_D7061_ = new_D7068_ & new_D7067_;
  assign new_D7062_ = new_D7070_ | new_D7069_;
  assign new_D7063_ = new_D7072_ | new_D7071_;
  assign new_D7064_ = new_D7074_ & new_D7073_;
  assign new_D7065_ = new_D7074_ & new_D7075_;
  assign new_D7066_ = new_D7067_ | new_D7076_;
  assign new_D7067_ = new_D7056_ | new_D7079_;
  assign new_D7068_ = new_D7078_ | new_D7077_;
  assign new_D7069_ = new_D7083_ & new_D7082_;
  assign new_D7070_ = new_D7081_ & new_D7080_;
  assign new_D7071_ = new_D7086_ | new_D7085_;
  assign new_D7072_ = new_D7081_ & new_D7084_;
  assign new_D7073_ = new_D7056_ | new_D7089_;
  assign new_D7074_ = new_D7088_ | new_D7087_;
  assign new_D7075_ = new_D7091_ | new_D7090_;
  assign new_D7076_ = ~new_D7067_ & new_D7093_;
  assign new_D7077_ = ~new_D7069_ & new_D7081_;
  assign new_D7078_ = new_D7069_ & ~new_D7081_;
  assign new_D7079_ = new_D7055_ & ~new_D7056_;
  assign new_D7080_ = ~new_D7102_ | ~new_D7103_;
  assign new_D7081_ = new_D7095_ | new_D7097_;
  assign new_D7082_ = new_D7105_ | new_D7104_;
  assign new_D7083_ = new_D7099_ | new_D7098_;
  assign new_D7084_ = ~new_D7107_ | ~new_D7106_;
  assign new_D7085_ = ~new_D7108_ & new_D7109_;
  assign new_D7086_ = new_D7108_ & ~new_D7109_;
  assign new_D7087_ = ~new_D7055_ & new_D7056_;
  assign new_D7088_ = new_D7055_ & ~new_D7056_;
  assign new_D7089_ = ~new_D7071_ | new_D7081_;
  assign new_D7090_ = new_D7071_ & new_D7081_;
  assign new_D7091_ = ~new_D7071_ & ~new_D7081_;
  assign new_D7092_ = new_D7113_ | new_D7112_;
  assign new_D7093_ = new_D7059_ | new_D7092_;
  assign new_D7094_ = new_D7117_ | new_D7116_;
  assign new_D7095_ = ~new_D7059_ & new_D7094_;
  assign new_D7096_ = new_D7115_ | new_D7114_;
  assign new_D7097_ = new_D7059_ & new_D7096_;
  assign new_D7098_ = new_D7057_ & ~new_D7067_;
  assign new_D7099_ = ~new_D7057_ & new_D7067_;
  assign new_D7100_ = ~new_D7056_ | ~new_D7081_;
  assign new_D7101_ = new_D7067_ & new_D7100_;
  assign new_D7102_ = ~new_D7067_ & ~new_D7101_;
  assign new_D7103_ = new_D7067_ | new_D7100_;
  assign new_D7104_ = ~new_D7057_ & new_D7058_;
  assign new_D7105_ = new_D7057_ & ~new_D7058_;
  assign new_D7106_ = new_D7074_ | new_D7111_;
  assign new_D7107_ = ~new_D7074_ & ~new_D7110_;
  assign new_D7108_ = new_D7057_ | new_D7074_;
  assign new_D7109_ = new_D7057_ | new_D7058_;
  assign new_D7110_ = new_D7074_ & new_D7111_;
  assign new_D7111_ = ~new_D7056_ | ~new_D7081_;
  assign new_D7112_ = new_D7089_ & new_D7109_;
  assign new_D7113_ = ~new_D7089_ & ~new_D7109_;
  assign new_D7114_ = new_D7118_ | new_D7119_;
  assign new_D7115_ = ~new_D7060_ & new_D7074_;
  assign new_D7116_ = new_D7120_ | new_D7121_;
  assign new_D7117_ = new_D7060_ & new_D7074_;
  assign new_D7118_ = ~new_D7060_ & ~new_D7074_;
  assign new_D7119_ = new_D7060_ & ~new_D7074_;
  assign new_D7120_ = new_D7060_ & ~new_D7074_;
  assign new_D7121_ = ~new_D7060_ & new_D7074_;
  assign new_D7122_ = new_F2272_;
  assign new_D7123_ = new_F2339_;
  assign new_D7124_ = new_F2406_;
  assign new_D7125_ = new_F2473_;
  assign new_D7126_ = new_F2540_;
  assign new_D7127_ = new_F2607_;
  assign new_D7128_ = new_D7135_ & new_D7134_;
  assign new_D7129_ = new_D7137_ | new_D7136_;
  assign new_D7130_ = new_D7139_ | new_D7138_;
  assign new_D7131_ = new_D7141_ & new_D7140_;
  assign new_D7132_ = new_D7141_ & new_D7142_;
  assign new_D7133_ = new_D7134_ | new_D7143_;
  assign new_D7134_ = new_D7123_ | new_D7146_;
  assign new_D7135_ = new_D7145_ | new_D7144_;
  assign new_D7136_ = new_D7150_ & new_D7149_;
  assign new_D7137_ = new_D7148_ & new_D7147_;
  assign new_D7138_ = new_D7153_ | new_D7152_;
  assign new_D7139_ = new_D7148_ & new_D7151_;
  assign new_D7140_ = new_D7123_ | new_D7156_;
  assign new_D7141_ = new_D7155_ | new_D7154_;
  assign new_D7142_ = new_D7158_ | new_D7157_;
  assign new_D7143_ = ~new_D7134_ & new_D7160_;
  assign new_D7144_ = ~new_D7136_ & new_D7148_;
  assign new_D7145_ = new_D7136_ & ~new_D7148_;
  assign new_D7146_ = new_D7122_ & ~new_D7123_;
  assign new_D7147_ = ~new_D7169_ | ~new_D7170_;
  assign new_D7148_ = new_D7162_ | new_D7164_;
  assign new_D7149_ = new_D7172_ | new_D7171_;
  assign new_D7150_ = new_D7166_ | new_D7165_;
  assign new_D7151_ = ~new_D7174_ | ~new_D7173_;
  assign new_D7152_ = ~new_D7175_ & new_D7176_;
  assign new_D7153_ = new_D7175_ & ~new_D7176_;
  assign new_D7154_ = ~new_D7122_ & new_D7123_;
  assign new_D7155_ = new_D7122_ & ~new_D7123_;
  assign new_D7156_ = ~new_D7138_ | new_D7148_;
  assign new_D7157_ = new_D7138_ & new_D7148_;
  assign new_D7158_ = ~new_D7138_ & ~new_D7148_;
  assign new_D7159_ = new_D7180_ | new_D7179_;
  assign new_D7160_ = new_D7126_ | new_D7159_;
  assign new_D7161_ = new_D7184_ | new_D7183_;
  assign new_D7162_ = ~new_D7126_ & new_D7161_;
  assign new_D7163_ = new_D7182_ | new_D7181_;
  assign new_D7164_ = new_D7126_ & new_D7163_;
  assign new_D7165_ = new_D7124_ & ~new_D7134_;
  assign new_D7166_ = ~new_D7124_ & new_D7134_;
  assign new_D7167_ = ~new_D7123_ | ~new_D7148_;
  assign new_D7168_ = new_D7134_ & new_D7167_;
  assign new_D7169_ = ~new_D7134_ & ~new_D7168_;
  assign new_D7170_ = new_D7134_ | new_D7167_;
  assign new_D7171_ = ~new_D7124_ & new_D7125_;
  assign new_D7172_ = new_D7124_ & ~new_D7125_;
  assign new_D7173_ = new_D7141_ | new_D7178_;
  assign new_D7174_ = ~new_D7141_ & ~new_D7177_;
  assign new_D7175_ = new_D7124_ | new_D7141_;
  assign new_D7176_ = new_D7124_ | new_D7125_;
  assign new_D7177_ = new_D7141_ & new_D7178_;
  assign new_D7178_ = ~new_D7123_ | ~new_D7148_;
  assign new_D7179_ = new_D7156_ & new_D7176_;
  assign new_D7180_ = ~new_D7156_ & ~new_D7176_;
  assign new_D7181_ = new_D7185_ | new_D7186_;
  assign new_D7182_ = ~new_D7127_ & new_D7141_;
  assign new_D7183_ = new_D7187_ | new_D7188_;
  assign new_D7184_ = new_D7127_ & new_D7141_;
  assign new_D7185_ = ~new_D7127_ & ~new_D7141_;
  assign new_D7186_ = new_D7127_ & ~new_D7141_;
  assign new_D7187_ = new_D7127_ & ~new_D7141_;
  assign new_D7188_ = ~new_D7127_ & new_D7141_;
  assign new_D7189_ = new_F2674_;
  assign new_D7190_ = new_F2741_;
  assign new_D7191_ = new_F2808_;
  assign new_D7192_ = new_F2875_;
  assign new_D7193_ = new_F2942_;
  assign new_D7194_ = new_F3009_;
  assign new_D7195_ = new_D7202_ & new_D7201_;
  assign new_D7196_ = new_D7204_ | new_D7203_;
  assign new_D7197_ = new_D7206_ | new_D7205_;
  assign new_D7198_ = new_D7208_ & new_D7207_;
  assign new_D7199_ = new_D7208_ & new_D7209_;
  assign new_D7200_ = new_D7201_ | new_D7210_;
  assign new_D7201_ = new_D7190_ | new_D7213_;
  assign new_D7202_ = new_D7212_ | new_D7211_;
  assign new_D7203_ = new_D7217_ & new_D7216_;
  assign new_D7204_ = new_D7215_ & new_D7214_;
  assign new_D7205_ = new_D7220_ | new_D7219_;
  assign new_D7206_ = new_D7215_ & new_D7218_;
  assign new_D7207_ = new_D7190_ | new_D7223_;
  assign new_D7208_ = new_D7222_ | new_D7221_;
  assign new_D7209_ = new_D7225_ | new_D7224_;
  assign new_D7210_ = ~new_D7201_ & new_D7227_;
  assign new_D7211_ = ~new_D7203_ & new_D7215_;
  assign new_D7212_ = new_D7203_ & ~new_D7215_;
  assign new_D7213_ = new_D7189_ & ~new_D7190_;
  assign new_D7214_ = ~new_D7236_ | ~new_D7237_;
  assign new_D7215_ = new_D7229_ | new_D7231_;
  assign new_D7216_ = new_D7239_ | new_D7238_;
  assign new_D7217_ = new_D7233_ | new_D7232_;
  assign new_D7218_ = ~new_D7241_ | ~new_D7240_;
  assign new_D7219_ = ~new_D7242_ & new_D7243_;
  assign new_D7220_ = new_D7242_ & ~new_D7243_;
  assign new_D7221_ = ~new_D7189_ & new_D7190_;
  assign new_D7222_ = new_D7189_ & ~new_D7190_;
  assign new_D7223_ = ~new_D7205_ | new_D7215_;
  assign new_D7224_ = new_D7205_ & new_D7215_;
  assign new_D7225_ = ~new_D7205_ & ~new_D7215_;
  assign new_D7226_ = new_D7247_ | new_D7246_;
  assign new_D7227_ = new_D7193_ | new_D7226_;
  assign new_D7228_ = new_D7251_ | new_D7250_;
  assign new_D7229_ = ~new_D7193_ & new_D7228_;
  assign new_D7230_ = new_D7249_ | new_D7248_;
  assign new_D7231_ = new_D7193_ & new_D7230_;
  assign new_D7232_ = new_D7191_ & ~new_D7201_;
  assign new_D7233_ = ~new_D7191_ & new_D7201_;
  assign new_D7234_ = ~new_D7190_ | ~new_D7215_;
  assign new_D7235_ = new_D7201_ & new_D7234_;
  assign new_D7236_ = ~new_D7201_ & ~new_D7235_;
  assign new_D7237_ = new_D7201_ | new_D7234_;
  assign new_D7238_ = ~new_D7191_ & new_D7192_;
  assign new_D7239_ = new_D7191_ & ~new_D7192_;
  assign new_D7240_ = new_D7208_ | new_D7245_;
  assign new_D7241_ = ~new_D7208_ & ~new_D7244_;
  assign new_D7242_ = new_D7191_ | new_D7208_;
  assign new_D7243_ = new_D7191_ | new_D7192_;
  assign new_D7244_ = new_D7208_ & new_D7245_;
  assign new_D7245_ = ~new_D7190_ | ~new_D7215_;
  assign new_D7246_ = new_D7223_ & new_D7243_;
  assign new_D7247_ = ~new_D7223_ & ~new_D7243_;
  assign new_D7248_ = new_D7252_ | new_D7253_;
  assign new_D7249_ = ~new_D7194_ & new_D7208_;
  assign new_D7250_ = new_D7254_ | new_D7255_;
  assign new_D7251_ = new_D7194_ & new_D7208_;
  assign new_D7252_ = ~new_D7194_ & ~new_D7208_;
  assign new_D7253_ = new_D7194_ & ~new_D7208_;
  assign new_D7254_ = new_D7194_ & ~new_D7208_;
  assign new_D7255_ = ~new_D7194_ & new_D7208_;
  assign new_D7256_ = new_F3076_;
  assign new_D7257_ = new_F3143_;
  assign new_D7258_ = new_F3210_;
  assign new_D7259_ = new_F3277_;
  assign new_D7260_ = new_F3344_;
  assign new_D7261_ = new_F3411_;
  assign new_D7262_ = new_D7269_ & new_D7268_;
  assign new_D7263_ = new_D7271_ | new_D7270_;
  assign new_D7264_ = new_D7273_ | new_D7272_;
  assign new_D7265_ = new_D7275_ & new_D7274_;
  assign new_D7266_ = new_D7275_ & new_D7276_;
  assign new_D7267_ = new_D7268_ | new_D7277_;
  assign new_D7268_ = new_D7257_ | new_D7280_;
  assign new_D7269_ = new_D7279_ | new_D7278_;
  assign new_D7270_ = new_D7284_ & new_D7283_;
  assign new_D7271_ = new_D7282_ & new_D7281_;
  assign new_D7272_ = new_D7287_ | new_D7286_;
  assign new_D7273_ = new_D7282_ & new_D7285_;
  assign new_D7274_ = new_D7257_ | new_D7290_;
  assign new_D7275_ = new_D7289_ | new_D7288_;
  assign new_D7276_ = new_D7292_ | new_D7291_;
  assign new_D7277_ = ~new_D7268_ & new_D7294_;
  assign new_D7278_ = ~new_D7270_ & new_D7282_;
  assign new_D7279_ = new_D7270_ & ~new_D7282_;
  assign new_D7280_ = new_D7256_ & ~new_D7257_;
  assign new_D7281_ = ~new_D7303_ | ~new_D7304_;
  assign new_D7282_ = new_D7296_ | new_D7298_;
  assign new_D7283_ = new_D7306_ | new_D7305_;
  assign new_D7284_ = new_D7300_ | new_D7299_;
  assign new_D7285_ = ~new_D7308_ | ~new_D7307_;
  assign new_D7286_ = ~new_D7309_ & new_D7310_;
  assign new_D7287_ = new_D7309_ & ~new_D7310_;
  assign new_D7288_ = ~new_D7256_ & new_D7257_;
  assign new_D7289_ = new_D7256_ & ~new_D7257_;
  assign new_D7290_ = ~new_D7272_ | new_D7282_;
  assign new_D7291_ = new_D7272_ & new_D7282_;
  assign new_D7292_ = ~new_D7272_ & ~new_D7282_;
  assign new_D7293_ = new_D7314_ | new_D7313_;
  assign new_D7294_ = new_D7260_ | new_D7293_;
  assign new_D7295_ = new_D7318_ | new_D7317_;
  assign new_D7296_ = ~new_D7260_ & new_D7295_;
  assign new_D7297_ = new_D7316_ | new_D7315_;
  assign new_D7298_ = new_D7260_ & new_D7297_;
  assign new_D7299_ = new_D7258_ & ~new_D7268_;
  assign new_D7300_ = ~new_D7258_ & new_D7268_;
  assign new_D7301_ = ~new_D7257_ | ~new_D7282_;
  assign new_D7302_ = new_D7268_ & new_D7301_;
  assign new_D7303_ = ~new_D7268_ & ~new_D7302_;
  assign new_D7304_ = new_D7268_ | new_D7301_;
  assign new_D7305_ = ~new_D7258_ & new_D7259_;
  assign new_D7306_ = new_D7258_ & ~new_D7259_;
  assign new_D7307_ = new_D7275_ | new_D7312_;
  assign new_D7308_ = ~new_D7275_ & ~new_D7311_;
  assign new_D7309_ = new_D7258_ | new_D7275_;
  assign new_D7310_ = new_D7258_ | new_D7259_;
  assign new_D7311_ = new_D7275_ & new_D7312_;
  assign new_D7312_ = ~new_D7257_ | ~new_D7282_;
  assign new_D7313_ = new_D7290_ & new_D7310_;
  assign new_D7314_ = ~new_D7290_ & ~new_D7310_;
  assign new_D7315_ = new_D7319_ | new_D7320_;
  assign new_D7316_ = ~new_D7261_ & new_D7275_;
  assign new_D7317_ = new_D7321_ | new_D7322_;
  assign new_D7318_ = new_D7261_ & new_D7275_;
  assign new_D7319_ = ~new_D7261_ & ~new_D7275_;
  assign new_D7320_ = new_D7261_ & ~new_D7275_;
  assign new_D7321_ = new_D7261_ & ~new_D7275_;
  assign new_D7322_ = ~new_D7261_ & new_D7275_;
  assign new_D7323_ = new_F3478_;
  assign new_D7324_ = new_F3545_;
  assign new_D7325_ = new_F3612_;
  assign new_D7326_ = new_F3679_;
  assign new_D7327_ = new_F3746_;
  assign new_D7328_ = new_F3813_;
  assign new_D7329_ = new_D7336_ & new_D7335_;
  assign new_D7330_ = new_D7338_ | new_D7337_;
  assign new_D7331_ = new_D7340_ | new_D7339_;
  assign new_D7332_ = new_D7342_ & new_D7341_;
  assign new_D7333_ = new_D7342_ & new_D7343_;
  assign new_D7334_ = new_D7335_ | new_D7344_;
  assign new_D7335_ = new_D7324_ | new_D7347_;
  assign new_D7336_ = new_D7346_ | new_D7345_;
  assign new_D7337_ = new_D7351_ & new_D7350_;
  assign new_D7338_ = new_D7349_ & new_D7348_;
  assign new_D7339_ = new_D7354_ | new_D7353_;
  assign new_D7340_ = new_D7349_ & new_D7352_;
  assign new_D7341_ = new_D7324_ | new_D7357_;
  assign new_D7342_ = new_D7356_ | new_D7355_;
  assign new_D7343_ = new_D7359_ | new_D7358_;
  assign new_D7344_ = ~new_D7335_ & new_D7361_;
  assign new_D7345_ = ~new_D7337_ & new_D7349_;
  assign new_D7346_ = new_D7337_ & ~new_D7349_;
  assign new_D7347_ = new_D7323_ & ~new_D7324_;
  assign new_D7348_ = ~new_D7370_ | ~new_D7371_;
  assign new_D7349_ = new_D7363_ | new_D7365_;
  assign new_D7350_ = new_D7373_ | new_D7372_;
  assign new_D7351_ = new_D7367_ | new_D7366_;
  assign new_D7352_ = ~new_D7375_ | ~new_D7374_;
  assign new_D7353_ = ~new_D7376_ & new_D7377_;
  assign new_D7354_ = new_D7376_ & ~new_D7377_;
  assign new_D7355_ = ~new_D7323_ & new_D7324_;
  assign new_D7356_ = new_D7323_ & ~new_D7324_;
  assign new_D7357_ = ~new_D7339_ | new_D7349_;
  assign new_D7358_ = new_D7339_ & new_D7349_;
  assign new_D7359_ = ~new_D7339_ & ~new_D7349_;
  assign new_D7360_ = new_D7381_ | new_D7380_;
  assign new_D7361_ = new_D7327_ | new_D7360_;
  assign new_D7362_ = new_D7385_ | new_D7384_;
  assign new_D7363_ = ~new_D7327_ & new_D7362_;
  assign new_D7364_ = new_D7383_ | new_D7382_;
  assign new_D7365_ = new_D7327_ & new_D7364_;
  assign new_D7366_ = new_D7325_ & ~new_D7335_;
  assign new_D7367_ = ~new_D7325_ & new_D7335_;
  assign new_D7368_ = ~new_D7324_ | ~new_D7349_;
  assign new_D7369_ = new_D7335_ & new_D7368_;
  assign new_D7370_ = ~new_D7335_ & ~new_D7369_;
  assign new_D7371_ = new_D7335_ | new_D7368_;
  assign new_D7372_ = ~new_D7325_ & new_D7326_;
  assign new_D7373_ = new_D7325_ & ~new_D7326_;
  assign new_D7374_ = new_D7342_ | new_D7379_;
  assign new_D7375_ = ~new_D7342_ & ~new_D7378_;
  assign new_D7376_ = new_D7325_ | new_D7342_;
  assign new_D7377_ = new_D7325_ | new_D7326_;
  assign new_D7378_ = new_D7342_ & new_D7379_;
  assign new_D7379_ = ~new_D7324_ | ~new_D7349_;
  assign new_D7380_ = new_D7357_ & new_D7377_;
  assign new_D7381_ = ~new_D7357_ & ~new_D7377_;
  assign new_D7382_ = new_D7386_ | new_D7387_;
  assign new_D7383_ = ~new_D7328_ & new_D7342_;
  assign new_D7384_ = new_D7388_ | new_D7389_;
  assign new_D7385_ = new_D7328_ & new_D7342_;
  assign new_D7386_ = ~new_D7328_ & ~new_D7342_;
  assign new_D7387_ = new_D7328_ & ~new_D7342_;
  assign new_D7388_ = new_D7328_ & ~new_D7342_;
  assign new_D7389_ = ~new_D7328_ & new_D7342_;
  assign new_D7390_ = new_F3880_;
  assign new_D7391_ = new_F3947_;
  assign new_D7392_ = new_F4014_;
  assign new_D7393_ = new_F4081_;
  assign new_D7394_ = new_F4148_;
  assign new_D7395_ = new_F4215_;
  assign new_D7396_ = new_D7403_ & new_D7402_;
  assign new_D7397_ = new_D7405_ | new_D7404_;
  assign new_D7398_ = new_D7407_ | new_D7406_;
  assign new_D7399_ = new_D7409_ & new_D7408_;
  assign new_D7400_ = new_D7409_ & new_D7410_;
  assign new_D7401_ = new_D7402_ | new_D7411_;
  assign new_D7402_ = new_D7391_ | new_D7414_;
  assign new_D7403_ = new_D7413_ | new_D7412_;
  assign new_D7404_ = new_D7418_ & new_D7417_;
  assign new_D7405_ = new_D7416_ & new_D7415_;
  assign new_D7406_ = new_D7421_ | new_D7420_;
  assign new_D7407_ = new_D7416_ & new_D7419_;
  assign new_D7408_ = new_D7391_ | new_D7424_;
  assign new_D7409_ = new_D7423_ | new_D7422_;
  assign new_D7410_ = new_D7426_ | new_D7425_;
  assign new_D7411_ = ~new_D7402_ & new_D7428_;
  assign new_D7412_ = ~new_D7404_ & new_D7416_;
  assign new_D7413_ = new_D7404_ & ~new_D7416_;
  assign new_D7414_ = new_D7390_ & ~new_D7391_;
  assign new_D7415_ = ~new_D7437_ | ~new_D7438_;
  assign new_D7416_ = new_D7430_ | new_D7432_;
  assign new_D7417_ = new_D7440_ | new_D7439_;
  assign new_D7418_ = new_D7434_ | new_D7433_;
  assign new_D7419_ = ~new_D7442_ | ~new_D7441_;
  assign new_D7420_ = ~new_D7443_ & new_D7444_;
  assign new_D7421_ = new_D7443_ & ~new_D7444_;
  assign new_D7422_ = ~new_D7390_ & new_D7391_;
  assign new_D7423_ = new_D7390_ & ~new_D7391_;
  assign new_D7424_ = ~new_D7406_ | new_D7416_;
  assign new_D7425_ = new_D7406_ & new_D7416_;
  assign new_D7426_ = ~new_D7406_ & ~new_D7416_;
  assign new_D7427_ = new_D7448_ | new_D7447_;
  assign new_D7428_ = new_D7394_ | new_D7427_;
  assign new_D7429_ = new_D7452_ | new_D7451_;
  assign new_D7430_ = ~new_D7394_ & new_D7429_;
  assign new_D7431_ = new_D7450_ | new_D7449_;
  assign new_D7432_ = new_D7394_ & new_D7431_;
  assign new_D7433_ = new_D7392_ & ~new_D7402_;
  assign new_D7434_ = ~new_D7392_ & new_D7402_;
  assign new_D7435_ = ~new_D7391_ | ~new_D7416_;
  assign new_D7436_ = new_D7402_ & new_D7435_;
  assign new_D7437_ = ~new_D7402_ & ~new_D7436_;
  assign new_D7438_ = new_D7402_ | new_D7435_;
  assign new_D7439_ = ~new_D7392_ & new_D7393_;
  assign new_D7440_ = new_D7392_ & ~new_D7393_;
  assign new_D7441_ = new_D7409_ | new_D7446_;
  assign new_D7442_ = ~new_D7409_ & ~new_D7445_;
  assign new_D7443_ = new_D7392_ | new_D7409_;
  assign new_D7444_ = new_D7392_ | new_D7393_;
  assign new_D7445_ = new_D7409_ & new_D7446_;
  assign new_D7446_ = ~new_D7391_ | ~new_D7416_;
  assign new_D7447_ = new_D7424_ & new_D7444_;
  assign new_D7448_ = ~new_D7424_ & ~new_D7444_;
  assign new_D7449_ = new_D7453_ | new_D7454_;
  assign new_D7450_ = ~new_D7395_ & new_D7409_;
  assign new_D7451_ = new_D7455_ | new_D7456_;
  assign new_D7452_ = new_D7395_ & new_D7409_;
  assign new_D7453_ = ~new_D7395_ & ~new_D7409_;
  assign new_D7454_ = new_D7395_ & ~new_D7409_;
  assign new_D7455_ = new_D7395_ & ~new_D7409_;
  assign new_D7456_ = ~new_D7395_ & new_D7409_;
  assign new_D7457_ = new_F4282_;
  assign new_D7458_ = new_F4349_;
  assign new_D7459_ = new_F4416_;
  assign new_D7460_ = new_F4483_;
  assign new_D7461_ = new_F4550_;
  assign new_D7462_ = new_F4617_;
  assign new_D7463_ = new_D7470_ & new_D7469_;
  assign new_D7464_ = new_D7472_ | new_D7471_;
  assign new_D7465_ = new_D7474_ | new_D7473_;
  assign new_D7466_ = new_D7476_ & new_D7475_;
  assign new_D7467_ = new_D7476_ & new_D7477_;
  assign new_D7468_ = new_D7469_ | new_D7478_;
  assign new_D7469_ = new_D7458_ | new_D7481_;
  assign new_D7470_ = new_D7480_ | new_D7479_;
  assign new_D7471_ = new_D7485_ & new_D7484_;
  assign new_D7472_ = new_D7483_ & new_D7482_;
  assign new_D7473_ = new_D7488_ | new_D7487_;
  assign new_D7474_ = new_D7483_ & new_D7486_;
  assign new_D7475_ = new_D7458_ | new_D7491_;
  assign new_D7476_ = new_D7490_ | new_D7489_;
  assign new_D7477_ = new_D7493_ | new_D7492_;
  assign new_D7478_ = ~new_D7469_ & new_D7495_;
  assign new_D7479_ = ~new_D7471_ & new_D7483_;
  assign new_D7480_ = new_D7471_ & ~new_D7483_;
  assign new_D7481_ = new_D7457_ & ~new_D7458_;
  assign new_D7482_ = ~new_D7504_ | ~new_D7505_;
  assign new_D7483_ = new_D7497_ | new_D7499_;
  assign new_D7484_ = new_D7507_ | new_D7506_;
  assign new_D7485_ = new_D7501_ | new_D7500_;
  assign new_D7486_ = ~new_D7509_ | ~new_D7508_;
  assign new_D7487_ = ~new_D7510_ & new_D7511_;
  assign new_D7488_ = new_D7510_ & ~new_D7511_;
  assign new_D7489_ = ~new_D7457_ & new_D7458_;
  assign new_D7490_ = new_D7457_ & ~new_D7458_;
  assign new_D7491_ = ~new_D7473_ | new_D7483_;
  assign new_D7492_ = new_D7473_ & new_D7483_;
  assign new_D7493_ = ~new_D7473_ & ~new_D7483_;
  assign new_D7494_ = new_D7515_ | new_D7514_;
  assign new_D7495_ = new_D7461_ | new_D7494_;
  assign new_D7496_ = new_D7519_ | new_D7518_;
  assign new_D7497_ = ~new_D7461_ & new_D7496_;
  assign new_D7498_ = new_D7517_ | new_D7516_;
  assign new_D7499_ = new_D7461_ & new_D7498_;
  assign new_D7500_ = new_D7459_ & ~new_D7469_;
  assign new_D7501_ = ~new_D7459_ & new_D7469_;
  assign new_D7502_ = ~new_D7458_ | ~new_D7483_;
  assign new_D7503_ = new_D7469_ & new_D7502_;
  assign new_D7504_ = ~new_D7469_ & ~new_D7503_;
  assign new_D7505_ = new_D7469_ | new_D7502_;
  assign new_D7506_ = ~new_D7459_ & new_D7460_;
  assign new_D7507_ = new_D7459_ & ~new_D7460_;
  assign new_D7508_ = new_D7476_ | new_D7513_;
  assign new_D7509_ = ~new_D7476_ & ~new_D7512_;
  assign new_D7510_ = new_D7459_ | new_D7476_;
  assign new_D7511_ = new_D7459_ | new_D7460_;
  assign new_D7512_ = new_D7476_ & new_D7513_;
  assign new_D7513_ = ~new_D7458_ | ~new_D7483_;
  assign new_D7514_ = new_D7491_ & new_D7511_;
  assign new_D7515_ = ~new_D7491_ & ~new_D7511_;
  assign new_D7516_ = new_D7520_ | new_D7521_;
  assign new_D7517_ = ~new_D7462_ & new_D7476_;
  assign new_D7518_ = new_D7522_ | new_D7523_;
  assign new_D7519_ = new_D7462_ & new_D7476_;
  assign new_D7520_ = ~new_D7462_ & ~new_D7476_;
  assign new_D7521_ = new_D7462_ & ~new_D7476_;
  assign new_D7522_ = new_D7462_ & ~new_D7476_;
  assign new_D7523_ = ~new_D7462_ & new_D7476_;
  assign new_D7524_ = new_F4684_;
  assign new_D7525_ = new_F4751_;
  assign new_D7526_ = new_F4818_;
  assign new_D7527_ = new_F4885_;
  assign new_D7528_ = new_F4952_;
  assign new_D7529_ = new_F5019_;
  assign new_D7530_ = new_D7537_ & new_D7536_;
  assign new_D7531_ = new_D7539_ | new_D7538_;
  assign new_D7532_ = new_D7541_ | new_D7540_;
  assign new_D7533_ = new_D7543_ & new_D7542_;
  assign new_D7534_ = new_D7543_ & new_D7544_;
  assign new_D7535_ = new_D7536_ | new_D7545_;
  assign new_D7536_ = new_D7525_ | new_D7548_;
  assign new_D7537_ = new_D7547_ | new_D7546_;
  assign new_D7538_ = new_D7552_ & new_D7551_;
  assign new_D7539_ = new_D7550_ & new_D7549_;
  assign new_D7540_ = new_D7555_ | new_D7554_;
  assign new_D7541_ = new_D7550_ & new_D7553_;
  assign new_D7542_ = new_D7525_ | new_D7558_;
  assign new_D7543_ = new_D7557_ | new_D7556_;
  assign new_D7544_ = new_D7560_ | new_D7559_;
  assign new_D7545_ = ~new_D7536_ & new_D7562_;
  assign new_D7546_ = ~new_D7538_ & new_D7550_;
  assign new_D7547_ = new_D7538_ & ~new_D7550_;
  assign new_D7548_ = new_D7524_ & ~new_D7525_;
  assign new_D7549_ = ~new_D7571_ | ~new_D7572_;
  assign new_D7550_ = new_D7564_ | new_D7566_;
  assign new_D7551_ = new_D7574_ | new_D7573_;
  assign new_D7552_ = new_D7568_ | new_D7567_;
  assign new_D7553_ = ~new_D7576_ | ~new_D7575_;
  assign new_D7554_ = ~new_D7577_ & new_D7578_;
  assign new_D7555_ = new_D7577_ & ~new_D7578_;
  assign new_D7556_ = ~new_D7524_ & new_D7525_;
  assign new_D7557_ = new_D7524_ & ~new_D7525_;
  assign new_D7558_ = ~new_D7540_ | new_D7550_;
  assign new_D7559_ = new_D7540_ & new_D7550_;
  assign new_D7560_ = ~new_D7540_ & ~new_D7550_;
  assign new_D7561_ = new_D7582_ | new_D7581_;
  assign new_D7562_ = new_D7528_ | new_D7561_;
  assign new_D7563_ = new_D7586_ | new_D7585_;
  assign new_D7564_ = ~new_D7528_ & new_D7563_;
  assign new_D7565_ = new_D7584_ | new_D7583_;
  assign new_D7566_ = new_D7528_ & new_D7565_;
  assign new_D7567_ = new_D7526_ & ~new_D7536_;
  assign new_D7568_ = ~new_D7526_ & new_D7536_;
  assign new_D7569_ = ~new_D7525_ | ~new_D7550_;
  assign new_D7570_ = new_D7536_ & new_D7569_;
  assign new_D7571_ = ~new_D7536_ & ~new_D7570_;
  assign new_D7572_ = new_D7536_ | new_D7569_;
  assign new_D7573_ = ~new_D7526_ & new_D7527_;
  assign new_D7574_ = new_D7526_ & ~new_D7527_;
  assign new_D7575_ = new_D7543_ | new_D7580_;
  assign new_D7576_ = ~new_D7543_ & ~new_D7579_;
  assign new_D7577_ = new_D7526_ | new_D7543_;
  assign new_D7578_ = new_D7526_ | new_D7527_;
  assign new_D7579_ = new_D7543_ & new_D7580_;
  assign new_D7580_ = ~new_D7525_ | ~new_D7550_;
  assign new_D7581_ = new_D7558_ & new_D7578_;
  assign new_D7582_ = ~new_D7558_ & ~new_D7578_;
  assign new_D7583_ = new_D7587_ | new_D7588_;
  assign new_D7584_ = ~new_D7529_ & new_D7543_;
  assign new_D7585_ = new_D7589_ | new_D7590_;
  assign new_D7586_ = new_D7529_ & new_D7543_;
  assign new_D7587_ = ~new_D7529_ & ~new_D7543_;
  assign new_D7588_ = new_D7529_ & ~new_D7543_;
  assign new_D7589_ = new_D7529_ & ~new_D7543_;
  assign new_D7590_ = ~new_D7529_ & new_D7543_;
  assign new_D7591_ = new_F5086_;
  assign new_D7592_ = new_F5153_;
  assign new_D7593_ = new_F5220_;
  assign new_D7594_ = new_F5287_;
  assign new_D7595_ = new_F5354_;
  assign new_D7596_ = new_F5421_;
  assign new_D7597_ = new_D7604_ & new_D7603_;
  assign new_D7598_ = new_D7606_ | new_D7605_;
  assign new_D7599_ = new_D7608_ | new_D7607_;
  assign new_D7600_ = new_D7610_ & new_D7609_;
  assign new_D7601_ = new_D7610_ & new_D7611_;
  assign new_D7602_ = new_D7603_ | new_D7612_;
  assign new_D7603_ = new_D7592_ | new_D7615_;
  assign new_D7604_ = new_D7614_ | new_D7613_;
  assign new_D7605_ = new_D7619_ & new_D7618_;
  assign new_D7606_ = new_D7617_ & new_D7616_;
  assign new_D7607_ = new_D7622_ | new_D7621_;
  assign new_D7608_ = new_D7617_ & new_D7620_;
  assign new_D7609_ = new_D7592_ | new_D7625_;
  assign new_D7610_ = new_D7624_ | new_D7623_;
  assign new_D7611_ = new_D7627_ | new_D7626_;
  assign new_D7612_ = ~new_D7603_ & new_D7629_;
  assign new_D7613_ = ~new_D7605_ & new_D7617_;
  assign new_D7614_ = new_D7605_ & ~new_D7617_;
  assign new_D7615_ = new_D7591_ & ~new_D7592_;
  assign new_D7616_ = ~new_D7638_ | ~new_D7639_;
  assign new_D7617_ = new_D7631_ | new_D7633_;
  assign new_D7618_ = new_D7641_ | new_D7640_;
  assign new_D7619_ = new_D7635_ | new_D7634_;
  assign new_D7620_ = ~new_D7643_ | ~new_D7642_;
  assign new_D7621_ = ~new_D7644_ & new_D7645_;
  assign new_D7622_ = new_D7644_ & ~new_D7645_;
  assign new_D7623_ = ~new_D7591_ & new_D7592_;
  assign new_D7624_ = new_D7591_ & ~new_D7592_;
  assign new_D7625_ = ~new_D7607_ | new_D7617_;
  assign new_D7626_ = new_D7607_ & new_D7617_;
  assign new_D7627_ = ~new_D7607_ & ~new_D7617_;
  assign new_D7628_ = new_D7649_ | new_D7648_;
  assign new_D7629_ = new_D7595_ | new_D7628_;
  assign new_D7630_ = new_D7653_ | new_D7652_;
  assign new_D7631_ = ~new_D7595_ & new_D7630_;
  assign new_D7632_ = new_D7651_ | new_D7650_;
  assign new_D7633_ = new_D7595_ & new_D7632_;
  assign new_D7634_ = new_D7593_ & ~new_D7603_;
  assign new_D7635_ = ~new_D7593_ & new_D7603_;
  assign new_D7636_ = ~new_D7592_ | ~new_D7617_;
  assign new_D7637_ = new_D7603_ & new_D7636_;
  assign new_D7638_ = ~new_D7603_ & ~new_D7637_;
  assign new_D7639_ = new_D7603_ | new_D7636_;
  assign new_D7640_ = ~new_D7593_ & new_D7594_;
  assign new_D7641_ = new_D7593_ & ~new_D7594_;
  assign new_D7642_ = new_D7610_ | new_D7647_;
  assign new_D7643_ = ~new_D7610_ & ~new_D7646_;
  assign new_D7644_ = new_D7593_ | new_D7610_;
  assign new_D7645_ = new_D7593_ | new_D7594_;
  assign new_D7646_ = new_D7610_ & new_D7647_;
  assign new_D7647_ = ~new_D7592_ | ~new_D7617_;
  assign new_D7648_ = new_D7625_ & new_D7645_;
  assign new_D7649_ = ~new_D7625_ & ~new_D7645_;
  assign new_D7650_ = new_D7654_ | new_D7655_;
  assign new_D7651_ = ~new_D7596_ & new_D7610_;
  assign new_D7652_ = new_D7656_ | new_D7657_;
  assign new_D7653_ = new_D7596_ & new_D7610_;
  assign new_D7654_ = ~new_D7596_ & ~new_D7610_;
  assign new_D7655_ = new_D7596_ & ~new_D7610_;
  assign new_D7656_ = new_D7596_ & ~new_D7610_;
  assign new_D7657_ = ~new_D7596_ & new_D7610_;
  assign new_D7658_ = new_F5488_;
  assign new_D7659_ = new_F5555_;
  assign new_D7660_ = new_F5622_;
  assign new_D7661_ = new_F5689_;
  assign new_D7662_ = new_F5756_;
  assign new_D7663_ = new_F5823_;
  assign new_D7664_ = new_D7671_ & new_D7670_;
  assign new_D7665_ = new_D7673_ | new_D7672_;
  assign new_D7666_ = new_D7675_ | new_D7674_;
  assign new_D7667_ = new_D7677_ & new_D7676_;
  assign new_D7668_ = new_D7677_ & new_D7678_;
  assign new_D7669_ = new_D7670_ | new_D7679_;
  assign new_D7670_ = new_D7659_ | new_D7682_;
  assign new_D7671_ = new_D7681_ | new_D7680_;
  assign new_D7672_ = new_D7686_ & new_D7685_;
  assign new_D7673_ = new_D7684_ & new_D7683_;
  assign new_D7674_ = new_D7689_ | new_D7688_;
  assign new_D7675_ = new_D7684_ & new_D7687_;
  assign new_D7676_ = new_D7659_ | new_D7692_;
  assign new_D7677_ = new_D7691_ | new_D7690_;
  assign new_D7678_ = new_D7694_ | new_D7693_;
  assign new_D7679_ = ~new_D7670_ & new_D7696_;
  assign new_D7680_ = ~new_D7672_ & new_D7684_;
  assign new_D7681_ = new_D7672_ & ~new_D7684_;
  assign new_D7682_ = new_D7658_ & ~new_D7659_;
  assign new_D7683_ = ~new_D7705_ | ~new_D7706_;
  assign new_D7684_ = new_D7698_ | new_D7700_;
  assign new_D7685_ = new_D7708_ | new_D7707_;
  assign new_D7686_ = new_D7702_ | new_D7701_;
  assign new_D7687_ = ~new_D7710_ | ~new_D7709_;
  assign new_D7688_ = ~new_D7711_ & new_D7712_;
  assign new_D7689_ = new_D7711_ & ~new_D7712_;
  assign new_D7690_ = ~new_D7658_ & new_D7659_;
  assign new_D7691_ = new_D7658_ & ~new_D7659_;
  assign new_D7692_ = ~new_D7674_ | new_D7684_;
  assign new_D7693_ = new_D7674_ & new_D7684_;
  assign new_D7694_ = ~new_D7674_ & ~new_D7684_;
  assign new_D7695_ = new_D7716_ | new_D7715_;
  assign new_D7696_ = new_D7662_ | new_D7695_;
  assign new_D7697_ = new_D7720_ | new_D7719_;
  assign new_D7698_ = ~new_D7662_ & new_D7697_;
  assign new_D7699_ = new_D7718_ | new_D7717_;
  assign new_D7700_ = new_D7662_ & new_D7699_;
  assign new_D7701_ = new_D7660_ & ~new_D7670_;
  assign new_D7702_ = ~new_D7660_ & new_D7670_;
  assign new_D7703_ = ~new_D7659_ | ~new_D7684_;
  assign new_D7704_ = new_D7670_ & new_D7703_;
  assign new_D7705_ = ~new_D7670_ & ~new_D7704_;
  assign new_D7706_ = new_D7670_ | new_D7703_;
  assign new_D7707_ = ~new_D7660_ & new_D7661_;
  assign new_D7708_ = new_D7660_ & ~new_D7661_;
  assign new_D7709_ = new_D7677_ | new_D7714_;
  assign new_D7710_ = ~new_D7677_ & ~new_D7713_;
  assign new_D7711_ = new_D7660_ | new_D7677_;
  assign new_D7712_ = new_D7660_ | new_D7661_;
  assign new_D7713_ = new_D7677_ & new_D7714_;
  assign new_D7714_ = ~new_D7659_ | ~new_D7684_;
  assign new_D7715_ = new_D7692_ & new_D7712_;
  assign new_D7716_ = ~new_D7692_ & ~new_D7712_;
  assign new_D7717_ = new_D7721_ | new_D7722_;
  assign new_D7718_ = ~new_D7663_ & new_D7677_;
  assign new_D7719_ = new_D7723_ | new_D7724_;
  assign new_D7720_ = new_D7663_ & new_D7677_;
  assign new_D7721_ = ~new_D7663_ & ~new_D7677_;
  assign new_D7722_ = new_D7663_ & ~new_D7677_;
  assign new_D7723_ = new_D7663_ & ~new_D7677_;
  assign new_D7724_ = ~new_D7663_ & new_D7677_;
  assign new_D7725_ = new_F5890_;
  assign new_D7726_ = new_F5957_;
  assign new_D7727_ = new_F6024_;
  assign new_D7728_ = new_F6091_;
  assign new_D7729_ = new_F6158_;
  assign new_D7730_ = new_F6225_;
  assign new_D7731_ = new_D7738_ & new_D7737_;
  assign new_D7732_ = new_D7740_ | new_D7739_;
  assign new_D7733_ = new_D7742_ | new_D7741_;
  assign new_D7734_ = new_D7744_ & new_D7743_;
  assign new_D7735_ = new_D7744_ & new_D7745_;
  assign new_D7736_ = new_D7737_ | new_D7746_;
  assign new_D7737_ = new_D7726_ | new_D7749_;
  assign new_D7738_ = new_D7748_ | new_D7747_;
  assign new_D7739_ = new_D7753_ & new_D7752_;
  assign new_D7740_ = new_D7751_ & new_D7750_;
  assign new_D7741_ = new_D7756_ | new_D7755_;
  assign new_D7742_ = new_D7751_ & new_D7754_;
  assign new_D7743_ = new_D7726_ | new_D7759_;
  assign new_D7744_ = new_D7758_ | new_D7757_;
  assign new_D7745_ = new_D7761_ | new_D7760_;
  assign new_D7746_ = ~new_D7737_ & new_D7763_;
  assign new_D7747_ = ~new_D7739_ & new_D7751_;
  assign new_D7748_ = new_D7739_ & ~new_D7751_;
  assign new_D7749_ = new_D7725_ & ~new_D7726_;
  assign new_D7750_ = ~new_D7772_ | ~new_D7773_;
  assign new_D7751_ = new_D7765_ | new_D7767_;
  assign new_D7752_ = new_D7775_ | new_D7774_;
  assign new_D7753_ = new_D7769_ | new_D7768_;
  assign new_D7754_ = ~new_D7777_ | ~new_D7776_;
  assign new_D7755_ = ~new_D7778_ & new_D7779_;
  assign new_D7756_ = new_D7778_ & ~new_D7779_;
  assign new_D7757_ = ~new_D7725_ & new_D7726_;
  assign new_D7758_ = new_D7725_ & ~new_D7726_;
  assign new_D7759_ = ~new_D7741_ | new_D7751_;
  assign new_D7760_ = new_D7741_ & new_D7751_;
  assign new_D7761_ = ~new_D7741_ & ~new_D7751_;
  assign new_D7762_ = new_D7783_ | new_D7782_;
  assign new_D7763_ = new_D7729_ | new_D7762_;
  assign new_D7764_ = new_D7787_ | new_D7786_;
  assign new_D7765_ = ~new_D7729_ & new_D7764_;
  assign new_D7766_ = new_D7785_ | new_D7784_;
  assign new_D7767_ = new_D7729_ & new_D7766_;
  assign new_D7768_ = new_D7727_ & ~new_D7737_;
  assign new_D7769_ = ~new_D7727_ & new_D7737_;
  assign new_D7770_ = ~new_D7726_ | ~new_D7751_;
  assign new_D7771_ = new_D7737_ & new_D7770_;
  assign new_D7772_ = ~new_D7737_ & ~new_D7771_;
  assign new_D7773_ = new_D7737_ | new_D7770_;
  assign new_D7774_ = ~new_D7727_ & new_D7728_;
  assign new_D7775_ = new_D7727_ & ~new_D7728_;
  assign new_D7776_ = new_D7744_ | new_D7781_;
  assign new_D7777_ = ~new_D7744_ & ~new_D7780_;
  assign new_D7778_ = new_D7727_ | new_D7744_;
  assign new_D7779_ = new_D7727_ | new_D7728_;
  assign new_D7780_ = new_D7744_ & new_D7781_;
  assign new_D7781_ = ~new_D7726_ | ~new_D7751_;
  assign new_D7782_ = new_D7759_ & new_D7779_;
  assign new_D7783_ = ~new_D7759_ & ~new_D7779_;
  assign new_D7784_ = new_D7788_ | new_D7789_;
  assign new_D7785_ = ~new_D7730_ & new_D7744_;
  assign new_D7786_ = new_D7790_ | new_D7791_;
  assign new_D7787_ = new_D7730_ & new_D7744_;
  assign new_D7788_ = ~new_D7730_ & ~new_D7744_;
  assign new_D7789_ = new_D7730_ & ~new_D7744_;
  assign new_D7790_ = new_D7730_ & ~new_D7744_;
  assign new_D7791_ = ~new_D7730_ & new_D7744_;
  assign new_D7792_ = new_F6292_;
  assign new_D7793_ = new_F6359_;
  assign new_D7794_ = new_F6426_;
  assign new_D7795_ = new_F6493_;
  assign new_D7796_ = new_F6560_;
  assign new_D7797_ = new_F6627_;
  assign new_D7798_ = new_D7805_ & new_D7804_;
  assign new_D7799_ = new_D7807_ | new_D7806_;
  assign new_D7800_ = new_D7809_ | new_D7808_;
  assign new_D7801_ = new_D7811_ & new_D7810_;
  assign new_D7802_ = new_D7811_ & new_D7812_;
  assign new_D7803_ = new_D7804_ | new_D7813_;
  assign new_D7804_ = new_D7793_ | new_D7816_;
  assign new_D7805_ = new_D7815_ | new_D7814_;
  assign new_D7806_ = new_D7820_ & new_D7819_;
  assign new_D7807_ = new_D7818_ & new_D7817_;
  assign new_D7808_ = new_D7823_ | new_D7822_;
  assign new_D7809_ = new_D7818_ & new_D7821_;
  assign new_D7810_ = new_D7793_ | new_D7826_;
  assign new_D7811_ = new_D7825_ | new_D7824_;
  assign new_D7812_ = new_D7828_ | new_D7827_;
  assign new_D7813_ = ~new_D7804_ & new_D7830_;
  assign new_D7814_ = ~new_D7806_ & new_D7818_;
  assign new_D7815_ = new_D7806_ & ~new_D7818_;
  assign new_D7816_ = new_D7792_ & ~new_D7793_;
  assign new_D7817_ = ~new_D7839_ | ~new_D7840_;
  assign new_D7818_ = new_D7832_ | new_D7834_;
  assign new_D7819_ = new_D7842_ | new_D7841_;
  assign new_D7820_ = new_D7836_ | new_D7835_;
  assign new_D7821_ = ~new_D7844_ | ~new_D7843_;
  assign new_D7822_ = ~new_D7845_ & new_D7846_;
  assign new_D7823_ = new_D7845_ & ~new_D7846_;
  assign new_D7824_ = ~new_D7792_ & new_D7793_;
  assign new_D7825_ = new_D7792_ & ~new_D7793_;
  assign new_D7826_ = ~new_D7808_ | new_D7818_;
  assign new_D7827_ = new_D7808_ & new_D7818_;
  assign new_D7828_ = ~new_D7808_ & ~new_D7818_;
  assign new_D7829_ = new_D7850_ | new_D7849_;
  assign new_D7830_ = new_D7796_ | new_D7829_;
  assign new_D7831_ = new_D7854_ | new_D7853_;
  assign new_D7832_ = ~new_D7796_ & new_D7831_;
  assign new_D7833_ = new_D7852_ | new_D7851_;
  assign new_D7834_ = new_D7796_ & new_D7833_;
  assign new_D7835_ = new_D7794_ & ~new_D7804_;
  assign new_D7836_ = ~new_D7794_ & new_D7804_;
  assign new_D7837_ = ~new_D7793_ | ~new_D7818_;
  assign new_D7838_ = new_D7804_ & new_D7837_;
  assign new_D7839_ = ~new_D7804_ & ~new_D7838_;
  assign new_D7840_ = new_D7804_ | new_D7837_;
  assign new_D7841_ = ~new_D7794_ & new_D7795_;
  assign new_D7842_ = new_D7794_ & ~new_D7795_;
  assign new_D7843_ = new_D7811_ | new_D7848_;
  assign new_D7844_ = ~new_D7811_ & ~new_D7847_;
  assign new_D7845_ = new_D7794_ | new_D7811_;
  assign new_D7846_ = new_D7794_ | new_D7795_;
  assign new_D7847_ = new_D7811_ & new_D7848_;
  assign new_D7848_ = ~new_D7793_ | ~new_D7818_;
  assign new_D7849_ = new_D7826_ & new_D7846_;
  assign new_D7850_ = ~new_D7826_ & ~new_D7846_;
  assign new_D7851_ = new_D7855_ | new_D7856_;
  assign new_D7852_ = ~new_D7797_ & new_D7811_;
  assign new_D7853_ = new_D7857_ | new_D7858_;
  assign new_D7854_ = new_D7797_ & new_D7811_;
  assign new_D7855_ = ~new_D7797_ & ~new_D7811_;
  assign new_D7856_ = new_D7797_ & ~new_D7811_;
  assign new_D7857_ = new_D7797_ & ~new_D7811_;
  assign new_D7858_ = ~new_D7797_ & new_D7811_;
  assign new_D7859_ = new_F6694_;
  assign new_D7860_ = new_F6761_;
  assign new_D7861_ = new_F6828_;
  assign new_D7862_ = new_F6895_;
  assign new_D7863_ = new_F6962_;
  assign new_D7864_ = new_F7029_;
  assign new_D7865_ = new_D7872_ & new_D7871_;
  assign new_D7866_ = new_D7874_ | new_D7873_;
  assign new_D7867_ = new_D7876_ | new_D7875_;
  assign new_D7868_ = new_D7878_ & new_D7877_;
  assign new_D7869_ = new_D7878_ & new_D7879_;
  assign new_D7870_ = new_D7871_ | new_D7880_;
  assign new_D7871_ = new_D7860_ | new_D7883_;
  assign new_D7872_ = new_D7882_ | new_D7881_;
  assign new_D7873_ = new_D7887_ & new_D7886_;
  assign new_D7874_ = new_D7885_ & new_D7884_;
  assign new_D7875_ = new_D7890_ | new_D7889_;
  assign new_D7876_ = new_D7885_ & new_D7888_;
  assign new_D7877_ = new_D7860_ | new_D7893_;
  assign new_D7878_ = new_D7892_ | new_D7891_;
  assign new_D7879_ = new_D7895_ | new_D7894_;
  assign new_D7880_ = ~new_D7871_ & new_D7897_;
  assign new_D7881_ = ~new_D7873_ & new_D7885_;
  assign new_D7882_ = new_D7873_ & ~new_D7885_;
  assign new_D7883_ = new_D7859_ & ~new_D7860_;
  assign new_D7884_ = ~new_D7906_ | ~new_D7907_;
  assign new_D7885_ = new_D7899_ | new_D7901_;
  assign new_D7886_ = new_D7909_ | new_D7908_;
  assign new_D7887_ = new_D7903_ | new_D7902_;
  assign new_D7888_ = ~new_D7911_ | ~new_D7910_;
  assign new_D7889_ = ~new_D7912_ & new_D7913_;
  assign new_D7890_ = new_D7912_ & ~new_D7913_;
  assign new_D7891_ = ~new_D7859_ & new_D7860_;
  assign new_D7892_ = new_D7859_ & ~new_D7860_;
  assign new_D7893_ = ~new_D7875_ | new_D7885_;
  assign new_D7894_ = new_D7875_ & new_D7885_;
  assign new_D7895_ = ~new_D7875_ & ~new_D7885_;
  assign new_D7896_ = new_D7917_ | new_D7916_;
  assign new_D7897_ = new_D7863_ | new_D7896_;
  assign new_D7898_ = new_D7921_ | new_D7920_;
  assign new_D7899_ = ~new_D7863_ & new_D7898_;
  assign new_D7900_ = new_D7919_ | new_D7918_;
  assign new_D7901_ = new_D7863_ & new_D7900_;
  assign new_D7902_ = new_D7861_ & ~new_D7871_;
  assign new_D7903_ = ~new_D7861_ & new_D7871_;
  assign new_D7904_ = ~new_D7860_ | ~new_D7885_;
  assign new_D7905_ = new_D7871_ & new_D7904_;
  assign new_D7906_ = ~new_D7871_ & ~new_D7905_;
  assign new_D7907_ = new_D7871_ | new_D7904_;
  assign new_D7908_ = ~new_D7861_ & new_D7862_;
  assign new_D7909_ = new_D7861_ & ~new_D7862_;
  assign new_D7910_ = new_D7878_ | new_D7915_;
  assign new_D7911_ = ~new_D7878_ & ~new_D7914_;
  assign new_D7912_ = new_D7861_ | new_D7878_;
  assign new_D7913_ = new_D7861_ | new_D7862_;
  assign new_D7914_ = new_D7878_ & new_D7915_;
  assign new_D7915_ = ~new_D7860_ | ~new_D7885_;
  assign new_D7916_ = new_D7893_ & new_D7913_;
  assign new_D7917_ = ~new_D7893_ & ~new_D7913_;
  assign new_D7918_ = new_D7922_ | new_D7923_;
  assign new_D7919_ = ~new_D7864_ & new_D7878_;
  assign new_D7920_ = new_D7924_ | new_D7925_;
  assign new_D7921_ = new_D7864_ & new_D7878_;
  assign new_D7922_ = ~new_D7864_ & ~new_D7878_;
  assign new_D7923_ = new_D7864_ & ~new_D7878_;
  assign new_D7924_ = new_D7864_ & ~new_D7878_;
  assign new_D7925_ = ~new_D7864_ & new_D7878_;
  assign new_D7926_ = new_F7096_;
  assign new_D7927_ = new_F7163_;
  assign new_D7928_ = new_F7230_;
  assign new_D7929_ = new_F7297_;
  assign new_D7930_ = new_F7364_;
  assign new_D7931_ = new_F7431_;
  assign new_D7932_ = new_D7939_ & new_D7938_;
  assign new_D7933_ = new_D7941_ | new_D7940_;
  assign new_D7934_ = new_D7943_ | new_D7942_;
  assign new_D7935_ = new_D7945_ & new_D7944_;
  assign new_D7936_ = new_D7945_ & new_D7946_;
  assign new_D7937_ = new_D7938_ | new_D7947_;
  assign new_D7938_ = new_D7927_ | new_D7950_;
  assign new_D7939_ = new_D7949_ | new_D7948_;
  assign new_D7940_ = new_D7954_ & new_D7953_;
  assign new_D7941_ = new_D7952_ & new_D7951_;
  assign new_D7942_ = new_D7957_ | new_D7956_;
  assign new_D7943_ = new_D7952_ & new_D7955_;
  assign new_D7944_ = new_D7927_ | new_D7960_;
  assign new_D7945_ = new_D7959_ | new_D7958_;
  assign new_D7946_ = new_D7962_ | new_D7961_;
  assign new_D7947_ = ~new_D7938_ & new_D7964_;
  assign new_D7948_ = ~new_D7940_ & new_D7952_;
  assign new_D7949_ = new_D7940_ & ~new_D7952_;
  assign new_D7950_ = new_D7926_ & ~new_D7927_;
  assign new_D7951_ = ~new_D7973_ | ~new_D7974_;
  assign new_D7952_ = new_D7966_ | new_D7968_;
  assign new_D7953_ = new_D7976_ | new_D7975_;
  assign new_D7954_ = new_D7970_ | new_D7969_;
  assign new_D7955_ = ~new_D7978_ | ~new_D7977_;
  assign new_D7956_ = ~new_D7979_ & new_D7980_;
  assign new_D7957_ = new_D7979_ & ~new_D7980_;
  assign new_D7958_ = ~new_D7926_ & new_D7927_;
  assign new_D7959_ = new_D7926_ & ~new_D7927_;
  assign new_D7960_ = ~new_D7942_ | new_D7952_;
  assign new_D7961_ = new_D7942_ & new_D7952_;
  assign new_D7962_ = ~new_D7942_ & ~new_D7952_;
  assign new_D7963_ = new_D7984_ | new_D7983_;
  assign new_D7964_ = new_D7930_ | new_D7963_;
  assign new_D7965_ = new_D7988_ | new_D7987_;
  assign new_D7966_ = ~new_D7930_ & new_D7965_;
  assign new_D7967_ = new_D7986_ | new_D7985_;
  assign new_D7968_ = new_D7930_ & new_D7967_;
  assign new_D7969_ = new_D7928_ & ~new_D7938_;
  assign new_D7970_ = ~new_D7928_ & new_D7938_;
  assign new_D7971_ = ~new_D7927_ | ~new_D7952_;
  assign new_D7972_ = new_D7938_ & new_D7971_;
  assign new_D7973_ = ~new_D7938_ & ~new_D7972_;
  assign new_D7974_ = new_D7938_ | new_D7971_;
  assign new_D7975_ = ~new_D7928_ & new_D7929_;
  assign new_D7976_ = new_D7928_ & ~new_D7929_;
  assign new_D7977_ = new_D7945_ | new_D7982_;
  assign new_D7978_ = ~new_D7945_ & ~new_D7981_;
  assign new_D7979_ = new_D7928_ | new_D7945_;
  assign new_D7980_ = new_D7928_ | new_D7929_;
  assign new_D7981_ = new_D7945_ & new_D7982_;
  assign new_D7982_ = ~new_D7927_ | ~new_D7952_;
  assign new_D7983_ = new_D7960_ & new_D7980_;
  assign new_D7984_ = ~new_D7960_ & ~new_D7980_;
  assign new_D7985_ = new_D7989_ | new_D7990_;
  assign new_D7986_ = ~new_D7931_ & new_D7945_;
  assign new_D7987_ = new_D7991_ | new_D7992_;
  assign new_D7988_ = new_D7931_ & new_D7945_;
  assign new_D7989_ = ~new_D7931_ & ~new_D7945_;
  assign new_D7990_ = new_D7931_ & ~new_D7945_;
  assign new_D7991_ = new_D7931_ & ~new_D7945_;
  assign new_D7992_ = ~new_D7931_ & new_D7945_;
  assign new_D7993_ = new_F7498_;
  assign new_D7994_ = new_F7565_;
  assign new_D7995_ = new_F7632_;
  assign new_D7996_ = new_F7699_;
  assign new_D7997_ = new_F7766_;
  assign new_D7998_ = new_F7833_;
  assign new_D7999_ = new_D8006_ & new_D8005_;
  assign new_D8000_ = new_D8008_ | new_D8007_;
  assign new_D8001_ = new_D8010_ | new_D8009_;
  assign new_D8002_ = new_D8012_ & new_D8011_;
  assign new_D8003_ = new_D8012_ & new_D8013_;
  assign new_D8004_ = new_D8005_ | new_D8014_;
  assign new_D8005_ = new_D7994_ | new_D8017_;
  assign new_D8006_ = new_D8016_ | new_D8015_;
  assign new_D8007_ = new_D8021_ & new_D8020_;
  assign new_D8008_ = new_D8019_ & new_D8018_;
  assign new_D8009_ = new_D8024_ | new_D8023_;
  assign new_D8010_ = new_D8019_ & new_D8022_;
  assign new_D8011_ = new_D7994_ | new_D8027_;
  assign new_D8012_ = new_D8026_ | new_D8025_;
  assign new_D8013_ = new_D8029_ | new_D8028_;
  assign new_D8014_ = ~new_D8005_ & new_D8031_;
  assign new_D8015_ = ~new_D8007_ & new_D8019_;
  assign new_D8016_ = new_D8007_ & ~new_D8019_;
  assign new_D8017_ = new_D7993_ & ~new_D7994_;
  assign new_D8018_ = ~new_D8040_ | ~new_D8041_;
  assign new_D8019_ = new_D8033_ | new_D8035_;
  assign new_D8020_ = new_D8043_ | new_D8042_;
  assign new_D8021_ = new_D8037_ | new_D8036_;
  assign new_D8022_ = ~new_D8045_ | ~new_D8044_;
  assign new_D8023_ = ~new_D8046_ & new_D8047_;
  assign new_D8024_ = new_D8046_ & ~new_D8047_;
  assign new_D8025_ = ~new_D7993_ & new_D7994_;
  assign new_D8026_ = new_D7993_ & ~new_D7994_;
  assign new_D8027_ = ~new_D8009_ | new_D8019_;
  assign new_D8028_ = new_D8009_ & new_D8019_;
  assign new_D8029_ = ~new_D8009_ & ~new_D8019_;
  assign new_D8030_ = new_D8051_ | new_D8050_;
  assign new_D8031_ = new_D7997_ | new_D8030_;
  assign new_D8032_ = new_D8055_ | new_D8054_;
  assign new_D8033_ = ~new_D7997_ & new_D8032_;
  assign new_D8034_ = new_D8053_ | new_D8052_;
  assign new_D8035_ = new_D7997_ & new_D8034_;
  assign new_D8036_ = new_D7995_ & ~new_D8005_;
  assign new_D8037_ = ~new_D7995_ & new_D8005_;
  assign new_D8038_ = ~new_D7994_ | ~new_D8019_;
  assign new_D8039_ = new_D8005_ & new_D8038_;
  assign new_D8040_ = ~new_D8005_ & ~new_D8039_;
  assign new_D8041_ = new_D8005_ | new_D8038_;
  assign new_D8042_ = ~new_D7995_ & new_D7996_;
  assign new_D8043_ = new_D7995_ & ~new_D7996_;
  assign new_D8044_ = new_D8012_ | new_D8049_;
  assign new_D8045_ = ~new_D8012_ & ~new_D8048_;
  assign new_D8046_ = new_D7995_ | new_D8012_;
  assign new_D8047_ = new_D7995_ | new_D7996_;
  assign new_D8048_ = new_D8012_ & new_D8049_;
  assign new_D8049_ = ~new_D7994_ | ~new_D8019_;
  assign new_D8050_ = new_D8027_ & new_D8047_;
  assign new_D8051_ = ~new_D8027_ & ~new_D8047_;
  assign new_D8052_ = new_D8056_ | new_D8057_;
  assign new_D8053_ = ~new_D7998_ & new_D8012_;
  assign new_D8054_ = new_D8058_ | new_D8059_;
  assign new_D8055_ = new_D7998_ & new_D8012_;
  assign new_D8056_ = ~new_D7998_ & ~new_D8012_;
  assign new_D8057_ = new_D7998_ & ~new_D8012_;
  assign new_D8058_ = new_D7998_ & ~new_D8012_;
  assign new_D8059_ = ~new_D7998_ & new_D8012_;
  assign new_D8060_ = new_F7900_;
  assign new_D8061_ = new_F7967_;
  assign new_D8062_ = new_F8034_;
  assign new_D8063_ = new_F8101_;
  assign new_D8064_ = new_F8168_;
  assign new_D8065_ = new_F8235_;
  assign new_D8066_ = new_D8073_ & new_D8072_;
  assign new_D8067_ = new_D8075_ | new_D8074_;
  assign new_D8068_ = new_D8077_ | new_D8076_;
  assign new_D8069_ = new_D8079_ & new_D8078_;
  assign new_D8070_ = new_D8079_ & new_D8080_;
  assign new_D8071_ = new_D8072_ | new_D8081_;
  assign new_D8072_ = new_D8061_ | new_D8084_;
  assign new_D8073_ = new_D8083_ | new_D8082_;
  assign new_D8074_ = new_D8088_ & new_D8087_;
  assign new_D8075_ = new_D8086_ & new_D8085_;
  assign new_D8076_ = new_D8091_ | new_D8090_;
  assign new_D8077_ = new_D8086_ & new_D8089_;
  assign new_D8078_ = new_D8061_ | new_D8094_;
  assign new_D8079_ = new_D8093_ | new_D8092_;
  assign new_D8080_ = new_D8096_ | new_D8095_;
  assign new_D8081_ = ~new_D8072_ & new_D8098_;
  assign new_D8082_ = ~new_D8074_ & new_D8086_;
  assign new_D8083_ = new_D8074_ & ~new_D8086_;
  assign new_D8084_ = new_D8060_ & ~new_D8061_;
  assign new_D8085_ = ~new_D8107_ | ~new_D8108_;
  assign new_D8086_ = new_D8100_ | new_D8102_;
  assign new_D8087_ = new_D8110_ | new_D8109_;
  assign new_D8088_ = new_D8104_ | new_D8103_;
  assign new_D8089_ = ~new_D8112_ | ~new_D8111_;
  assign new_D8090_ = ~new_D8113_ & new_D8114_;
  assign new_D8091_ = new_D8113_ & ~new_D8114_;
  assign new_D8092_ = ~new_D8060_ & new_D8061_;
  assign new_D8093_ = new_D8060_ & ~new_D8061_;
  assign new_D8094_ = ~new_D8076_ | new_D8086_;
  assign new_D8095_ = new_D8076_ & new_D8086_;
  assign new_D8096_ = ~new_D8076_ & ~new_D8086_;
  assign new_D8097_ = new_D8118_ | new_D8117_;
  assign new_D8098_ = new_D8064_ | new_D8097_;
  assign new_D8099_ = new_D8122_ | new_D8121_;
  assign new_D8100_ = ~new_D8064_ & new_D8099_;
  assign new_D8101_ = new_D8120_ | new_D8119_;
  assign new_D8102_ = new_D8064_ & new_D8101_;
  assign new_D8103_ = new_D8062_ & ~new_D8072_;
  assign new_D8104_ = ~new_D8062_ & new_D8072_;
  assign new_D8105_ = ~new_D8061_ | ~new_D8086_;
  assign new_D8106_ = new_D8072_ & new_D8105_;
  assign new_D8107_ = ~new_D8072_ & ~new_D8106_;
  assign new_D8108_ = new_D8072_ | new_D8105_;
  assign new_D8109_ = ~new_D8062_ & new_D8063_;
  assign new_D8110_ = new_D8062_ & ~new_D8063_;
  assign new_D8111_ = new_D8079_ | new_D8116_;
  assign new_D8112_ = ~new_D8079_ & ~new_D8115_;
  assign new_D8113_ = new_D8062_ | new_D8079_;
  assign new_D8114_ = new_D8062_ | new_D8063_;
  assign new_D8115_ = new_D8079_ & new_D8116_;
  assign new_D8116_ = ~new_D8061_ | ~new_D8086_;
  assign new_D8117_ = new_D8094_ & new_D8114_;
  assign new_D8118_ = ~new_D8094_ & ~new_D8114_;
  assign new_D8119_ = new_D8123_ | new_D8124_;
  assign new_D8120_ = ~new_D8065_ & new_D8079_;
  assign new_D8121_ = new_D8125_ | new_D8126_;
  assign new_D8122_ = new_D8065_ & new_D8079_;
  assign new_D8123_ = ~new_D8065_ & ~new_D8079_;
  assign new_D8124_ = new_D8065_ & ~new_D8079_;
  assign new_D8125_ = new_D8065_ & ~new_D8079_;
  assign new_D8126_ = ~new_D8065_ & new_D8079_;
  assign new_D8127_ = new_F8302_;
  assign new_D8128_ = new_F8369_;
  assign new_D8129_ = new_F8436_;
  assign new_D8130_ = new_F8503_;
  assign new_D8131_ = new_F8570_;
  assign new_D8132_ = new_F8637_;
  assign new_D8133_ = new_D8140_ & new_D8139_;
  assign new_D8134_ = new_D8142_ | new_D8141_;
  assign new_D8135_ = new_D8144_ | new_D8143_;
  assign new_D8136_ = new_D8146_ & new_D8145_;
  assign new_D8137_ = new_D8146_ & new_D8147_;
  assign new_D8138_ = new_D8139_ | new_D8148_;
  assign new_D8139_ = new_D8128_ | new_D8151_;
  assign new_D8140_ = new_D8150_ | new_D8149_;
  assign new_D8141_ = new_D8155_ & new_D8154_;
  assign new_D8142_ = new_D8153_ & new_D8152_;
  assign new_D8143_ = new_D8158_ | new_D8157_;
  assign new_D8144_ = new_D8153_ & new_D8156_;
  assign new_D8145_ = new_D8128_ | new_D8161_;
  assign new_D8146_ = new_D8160_ | new_D8159_;
  assign new_D8147_ = new_D8163_ | new_D8162_;
  assign new_D8148_ = ~new_D8139_ & new_D8165_;
  assign new_D8149_ = ~new_D8141_ & new_D8153_;
  assign new_D8150_ = new_D8141_ & ~new_D8153_;
  assign new_D8151_ = new_D8127_ & ~new_D8128_;
  assign new_D8152_ = ~new_D8174_ | ~new_D8175_;
  assign new_D8153_ = new_D8167_ | new_D8169_;
  assign new_D8154_ = new_D8177_ | new_D8176_;
  assign new_D8155_ = new_D8171_ | new_D8170_;
  assign new_D8156_ = ~new_D8179_ | ~new_D8178_;
  assign new_D8157_ = ~new_D8180_ & new_D8181_;
  assign new_D8158_ = new_D8180_ & ~new_D8181_;
  assign new_D8159_ = ~new_D8127_ & new_D8128_;
  assign new_D8160_ = new_D8127_ & ~new_D8128_;
  assign new_D8161_ = ~new_D8143_ | new_D8153_;
  assign new_D8162_ = new_D8143_ & new_D8153_;
  assign new_D8163_ = ~new_D8143_ & ~new_D8153_;
  assign new_D8164_ = new_D8185_ | new_D8184_;
  assign new_D8165_ = new_D8131_ | new_D8164_;
  assign new_D8166_ = new_D8189_ | new_D8188_;
  assign new_D8167_ = ~new_D8131_ & new_D8166_;
  assign new_D8168_ = new_D8187_ | new_D8186_;
  assign new_D8169_ = new_D8131_ & new_D8168_;
  assign new_D8170_ = new_D8129_ & ~new_D8139_;
  assign new_D8171_ = ~new_D8129_ & new_D8139_;
  assign new_D8172_ = ~new_D8128_ | ~new_D8153_;
  assign new_D8173_ = new_D8139_ & new_D8172_;
  assign new_D8174_ = ~new_D8139_ & ~new_D8173_;
  assign new_D8175_ = new_D8139_ | new_D8172_;
  assign new_D8176_ = ~new_D8129_ & new_D8130_;
  assign new_D8177_ = new_D8129_ & ~new_D8130_;
  assign new_D8178_ = new_D8146_ | new_D8183_;
  assign new_D8179_ = ~new_D8146_ & ~new_D8182_;
  assign new_D8180_ = new_D8129_ | new_D8146_;
  assign new_D8181_ = new_D8129_ | new_D8130_;
  assign new_D8182_ = new_D8146_ & new_D8183_;
  assign new_D8183_ = ~new_D8128_ | ~new_D8153_;
  assign new_D8184_ = new_D8161_ & new_D8181_;
  assign new_D8185_ = ~new_D8161_ & ~new_D8181_;
  assign new_D8186_ = new_D8190_ | new_D8191_;
  assign new_D8187_ = ~new_D8132_ & new_D8146_;
  assign new_D8188_ = new_D8192_ | new_D8193_;
  assign new_D8189_ = new_D8132_ & new_D8146_;
  assign new_D8190_ = ~new_D8132_ & ~new_D8146_;
  assign new_D8191_ = new_D8132_ & ~new_D8146_;
  assign new_D8192_ = new_D8132_ & ~new_D8146_;
  assign new_D8193_ = ~new_D8132_ & new_D8146_;
  assign new_D8194_ = new_F8704_;
  assign new_D8195_ = new_F8771_;
  assign new_D8196_ = new_F8838_;
  assign new_D8197_ = new_F8905_;
  assign new_D8198_ = new_F8972_;
  assign new_D8199_ = new_F9039_;
  assign new_D8200_ = new_D8207_ & new_D8206_;
  assign new_D8201_ = new_D8209_ | new_D8208_;
  assign new_D8202_ = new_D8211_ | new_D8210_;
  assign new_D8203_ = new_D8213_ & new_D8212_;
  assign new_D8204_ = new_D8213_ & new_D8214_;
  assign new_D8205_ = new_D8206_ | new_D8215_;
  assign new_D8206_ = new_D8195_ | new_D8218_;
  assign new_D8207_ = new_D8217_ | new_D8216_;
  assign new_D8208_ = new_D8222_ & new_D8221_;
  assign new_D8209_ = new_D8220_ & new_D8219_;
  assign new_D8210_ = new_D8225_ | new_D8224_;
  assign new_D8211_ = new_D8220_ & new_D8223_;
  assign new_D8212_ = new_D8195_ | new_D8228_;
  assign new_D8213_ = new_D8227_ | new_D8226_;
  assign new_D8214_ = new_D8230_ | new_D8229_;
  assign new_D8215_ = ~new_D8206_ & new_D8232_;
  assign new_D8216_ = ~new_D8208_ & new_D8220_;
  assign new_D8217_ = new_D8208_ & ~new_D8220_;
  assign new_D8218_ = new_D8194_ & ~new_D8195_;
  assign new_D8219_ = ~new_D8241_ | ~new_D8242_;
  assign new_D8220_ = new_D8234_ | new_D8236_;
  assign new_D8221_ = new_D8244_ | new_D8243_;
  assign new_D8222_ = new_D8238_ | new_D8237_;
  assign new_D8223_ = ~new_D8246_ | ~new_D8245_;
  assign new_D8224_ = ~new_D8247_ & new_D8248_;
  assign new_D8225_ = new_D8247_ & ~new_D8248_;
  assign new_D8226_ = ~new_D8194_ & new_D8195_;
  assign new_D8227_ = new_D8194_ & ~new_D8195_;
  assign new_D8228_ = ~new_D8210_ | new_D8220_;
  assign new_D8229_ = new_D8210_ & new_D8220_;
  assign new_D8230_ = ~new_D8210_ & ~new_D8220_;
  assign new_D8231_ = new_D8252_ | new_D8251_;
  assign new_D8232_ = new_D8198_ | new_D8231_;
  assign new_D8233_ = new_D8256_ | new_D8255_;
  assign new_D8234_ = ~new_D8198_ & new_D8233_;
  assign new_D8235_ = new_D8254_ | new_D8253_;
  assign new_D8236_ = new_D8198_ & new_D8235_;
  assign new_D8237_ = new_D8196_ & ~new_D8206_;
  assign new_D8238_ = ~new_D8196_ & new_D8206_;
  assign new_D8239_ = ~new_D8195_ | ~new_D8220_;
  assign new_D8240_ = new_D8206_ & new_D8239_;
  assign new_D8241_ = ~new_D8206_ & ~new_D8240_;
  assign new_D8242_ = new_D8206_ | new_D8239_;
  assign new_D8243_ = ~new_D8196_ & new_D8197_;
  assign new_D8244_ = new_D8196_ & ~new_D8197_;
  assign new_D8245_ = new_D8213_ | new_D8250_;
  assign new_D8246_ = ~new_D8213_ & ~new_D8249_;
  assign new_D8247_ = new_D8196_ | new_D8213_;
  assign new_D8248_ = new_D8196_ | new_D8197_;
  assign new_D8249_ = new_D8213_ & new_D8250_;
  assign new_D8250_ = ~new_D8195_ | ~new_D8220_;
  assign new_D8251_ = new_D8228_ & new_D8248_;
  assign new_D8252_ = ~new_D8228_ & ~new_D8248_;
  assign new_D8253_ = new_D8257_ | new_D8258_;
  assign new_D8254_ = ~new_D8199_ & new_D8213_;
  assign new_D8255_ = new_D8259_ | new_D8260_;
  assign new_D8256_ = new_D8199_ & new_D8213_;
  assign new_D8257_ = ~new_D8199_ & ~new_D8213_;
  assign new_D8258_ = new_D8199_ & ~new_D8213_;
  assign new_D8259_ = new_D8199_ & ~new_D8213_;
  assign new_D8260_ = ~new_D8199_ & new_D8213_;
  assign new_D8261_ = new_F9106_;
  assign new_D8262_ = new_F9173_;
  assign new_D8263_ = new_F9240_;
  assign new_D8264_ = new_F9307_;
  assign new_D8265_ = new_F9374_;
  assign new_D8266_ = new_F9441_;
  assign new_D8267_ = new_D8274_ & new_D8273_;
  assign new_D8268_ = new_D8276_ | new_D8275_;
  assign new_D8269_ = new_D8278_ | new_D8277_;
  assign new_D8270_ = new_D8280_ & new_D8279_;
  assign new_D8271_ = new_D8280_ & new_D8281_;
  assign new_D8272_ = new_D8273_ | new_D8282_;
  assign new_D8273_ = new_D8262_ | new_D8285_;
  assign new_D8274_ = new_D8284_ | new_D8283_;
  assign new_D8275_ = new_D8289_ & new_D8288_;
  assign new_D8276_ = new_D8287_ & new_D8286_;
  assign new_D8277_ = new_D8292_ | new_D8291_;
  assign new_D8278_ = new_D8287_ & new_D8290_;
  assign new_D8279_ = new_D8262_ | new_D8295_;
  assign new_D8280_ = new_D8294_ | new_D8293_;
  assign new_D8281_ = new_D8297_ | new_D8296_;
  assign new_D8282_ = ~new_D8273_ & new_D8299_;
  assign new_D8283_ = ~new_D8275_ & new_D8287_;
  assign new_D8284_ = new_D8275_ & ~new_D8287_;
  assign new_D8285_ = new_D8261_ & ~new_D8262_;
  assign new_D8286_ = ~new_D8308_ | ~new_D8309_;
  assign new_D8287_ = new_D8301_ | new_D8303_;
  assign new_D8288_ = new_D8311_ | new_D8310_;
  assign new_D8289_ = new_D8305_ | new_D8304_;
  assign new_D8290_ = ~new_D8313_ | ~new_D8312_;
  assign new_D8291_ = ~new_D8314_ & new_D8315_;
  assign new_D8292_ = new_D8314_ & ~new_D8315_;
  assign new_D8293_ = ~new_D8261_ & new_D8262_;
  assign new_D8294_ = new_D8261_ & ~new_D8262_;
  assign new_D8295_ = ~new_D8277_ | new_D8287_;
  assign new_D8296_ = new_D8277_ & new_D8287_;
  assign new_D8297_ = ~new_D8277_ & ~new_D8287_;
  assign new_D8298_ = new_D8319_ | new_D8318_;
  assign new_D8299_ = new_D8265_ | new_D8298_;
  assign new_D8300_ = new_D8323_ | new_D8322_;
  assign new_D8301_ = ~new_D8265_ & new_D8300_;
  assign new_D8302_ = new_D8321_ | new_D8320_;
  assign new_D8303_ = new_D8265_ & new_D8302_;
  assign new_D8304_ = new_D8263_ & ~new_D8273_;
  assign new_D8305_ = ~new_D8263_ & new_D8273_;
  assign new_D8306_ = ~new_D8262_ | ~new_D8287_;
  assign new_D8307_ = new_D8273_ & new_D8306_;
  assign new_D8308_ = ~new_D8273_ & ~new_D8307_;
  assign new_D8309_ = new_D8273_ | new_D8306_;
  assign new_D8310_ = ~new_D8263_ & new_D8264_;
  assign new_D8311_ = new_D8263_ & ~new_D8264_;
  assign new_D8312_ = new_D8280_ | new_D8317_;
  assign new_D8313_ = ~new_D8280_ & ~new_D8316_;
  assign new_D8314_ = new_D8263_ | new_D8280_;
  assign new_D8315_ = new_D8263_ | new_D8264_;
  assign new_D8316_ = new_D8280_ & new_D8317_;
  assign new_D8317_ = ~new_D8262_ | ~new_D8287_;
  assign new_D8318_ = new_D8295_ & new_D8315_;
  assign new_D8319_ = ~new_D8295_ & ~new_D8315_;
  assign new_D8320_ = new_D8324_ | new_D8325_;
  assign new_D8321_ = ~new_D8266_ & new_D8280_;
  assign new_D8322_ = new_D8326_ | new_D8327_;
  assign new_D8323_ = new_D8266_ & new_D8280_;
  assign new_D8324_ = ~new_D8266_ & ~new_D8280_;
  assign new_D8325_ = new_D8266_ & ~new_D8280_;
  assign new_D8326_ = new_D8266_ & ~new_D8280_;
  assign new_D8327_ = ~new_D8266_ & new_D8280_;
  assign new_D8328_ = new_F9508_;
  assign new_D8329_ = new_F9575_;
  assign new_D8330_ = new_F9642_;
  assign new_D8331_ = new_F9709_;
  assign new_D8332_ = new_F9776_;
  assign new_D8333_ = new_F9843_;
  assign new_D8334_ = new_D8341_ & new_D8340_;
  assign new_D8335_ = new_D8343_ | new_D8342_;
  assign new_D8336_ = new_D8345_ | new_D8344_;
  assign new_D8337_ = new_D8347_ & new_D8346_;
  assign new_D8338_ = new_D8347_ & new_D8348_;
  assign new_D8339_ = new_D8340_ | new_D8349_;
  assign new_D8340_ = new_D8329_ | new_D8352_;
  assign new_D8341_ = new_D8351_ | new_D8350_;
  assign new_D8342_ = new_D8356_ & new_D8355_;
  assign new_D8343_ = new_D8354_ & new_D8353_;
  assign new_D8344_ = new_D8359_ | new_D8358_;
  assign new_D8345_ = new_D8354_ & new_D8357_;
  assign new_D8346_ = new_D8329_ | new_D8362_;
  assign new_D8347_ = new_D8361_ | new_D8360_;
  assign new_D8348_ = new_D8364_ | new_D8363_;
  assign new_D8349_ = ~new_D8340_ & new_D8366_;
  assign new_D8350_ = ~new_D8342_ & new_D8354_;
  assign new_D8351_ = new_D8342_ & ~new_D8354_;
  assign new_D8352_ = new_D8328_ & ~new_D8329_;
  assign new_D8353_ = ~new_D8375_ | ~new_D8376_;
  assign new_D8354_ = new_D8368_ | new_D8370_;
  assign new_D8355_ = new_D8378_ | new_D8377_;
  assign new_D8356_ = new_D8372_ | new_D8371_;
  assign new_D8357_ = ~new_D8380_ | ~new_D8379_;
  assign new_D8358_ = ~new_D8381_ & new_D8382_;
  assign new_D8359_ = new_D8381_ & ~new_D8382_;
  assign new_D8360_ = ~new_D8328_ & new_D8329_;
  assign new_D8361_ = new_D8328_ & ~new_D8329_;
  assign new_D8362_ = ~new_D8344_ | new_D8354_;
  assign new_D8363_ = new_D8344_ & new_D8354_;
  assign new_D8364_ = ~new_D8344_ & ~new_D8354_;
  assign new_D8365_ = new_D8386_ | new_D8385_;
  assign new_D8366_ = new_D8332_ | new_D8365_;
  assign new_D8367_ = new_D8390_ | new_D8389_;
  assign new_D8368_ = ~new_D8332_ & new_D8367_;
  assign new_D8369_ = new_D8388_ | new_D8387_;
  assign new_D8370_ = new_D8332_ & new_D8369_;
  assign new_D8371_ = new_D8330_ & ~new_D8340_;
  assign new_D8372_ = ~new_D8330_ & new_D8340_;
  assign new_D8373_ = ~new_D8329_ | ~new_D8354_;
  assign new_D8374_ = new_D8340_ & new_D8373_;
  assign new_D8375_ = ~new_D8340_ & ~new_D8374_;
  assign new_D8376_ = new_D8340_ | new_D8373_;
  assign new_D8377_ = ~new_D8330_ & new_D8331_;
  assign new_D8378_ = new_D8330_ & ~new_D8331_;
  assign new_D8379_ = new_D8347_ | new_D8384_;
  assign new_D8380_ = ~new_D8347_ & ~new_D8383_;
  assign new_D8381_ = new_D8330_ | new_D8347_;
  assign new_D8382_ = new_D8330_ | new_D8331_;
  assign new_D8383_ = new_D8347_ & new_D8384_;
  assign new_D8384_ = ~new_D8329_ | ~new_D8354_;
  assign new_D8385_ = new_D8362_ & new_D8382_;
  assign new_D8386_ = ~new_D8362_ & ~new_D8382_;
  assign new_D8387_ = new_D8391_ | new_D8392_;
  assign new_D8388_ = ~new_D8333_ & new_D8347_;
  assign new_D8389_ = new_D8393_ | new_D8394_;
  assign new_D8390_ = new_D8333_ & new_D8347_;
  assign new_D8391_ = ~new_D8333_ & ~new_D8347_;
  assign new_D8392_ = new_D8333_ & ~new_D8347_;
  assign new_D8393_ = new_D8333_ & ~new_D8347_;
  assign new_D8394_ = ~new_D8333_ & new_D8347_;
  assign new_D8395_ = new_F9910_;
  assign new_D8396_ = new_F9977_;
  assign new_D8397_ = new_G45_;
  assign new_D8398_ = new_G112_;
  assign new_D8399_ = new_G179_;
  assign new_D8400_ = new_G246_;
  assign new_D8401_ = new_D8408_ & new_D8407_;
  assign new_D8402_ = new_D8410_ | new_D8409_;
  assign new_D8403_ = new_D8412_ | new_D8411_;
  assign new_D8404_ = new_D8414_ & new_D8413_;
  assign new_D8405_ = new_D8414_ & new_D8415_;
  assign new_D8406_ = new_D8407_ | new_D8416_;
  assign new_D8407_ = new_D8396_ | new_D8419_;
  assign new_D8408_ = new_D8418_ | new_D8417_;
  assign new_D8409_ = new_D8423_ & new_D8422_;
  assign new_D8410_ = new_D8421_ & new_D8420_;
  assign new_D8411_ = new_D8426_ | new_D8425_;
  assign new_D8412_ = new_D8421_ & new_D8424_;
  assign new_D8413_ = new_D8396_ | new_D8429_;
  assign new_D8414_ = new_D8428_ | new_D8427_;
  assign new_D8415_ = new_D8431_ | new_D8430_;
  assign new_D8416_ = ~new_D8407_ & new_D8433_;
  assign new_D8417_ = ~new_D8409_ & new_D8421_;
  assign new_D8418_ = new_D8409_ & ~new_D8421_;
  assign new_D8419_ = new_D8395_ & ~new_D8396_;
  assign new_D8420_ = ~new_D8442_ | ~new_D8443_;
  assign new_D8421_ = new_D8435_ | new_D8437_;
  assign new_D8422_ = new_D8445_ | new_D8444_;
  assign new_D8423_ = new_D8439_ | new_D8438_;
  assign new_D8424_ = ~new_D8447_ | ~new_D8446_;
  assign new_D8425_ = ~new_D8448_ & new_D8449_;
  assign new_D8426_ = new_D8448_ & ~new_D8449_;
  assign new_D8427_ = ~new_D8395_ & new_D8396_;
  assign new_D8428_ = new_D8395_ & ~new_D8396_;
  assign new_D8429_ = ~new_D8411_ | new_D8421_;
  assign new_D8430_ = new_D8411_ & new_D8421_;
  assign new_D8431_ = ~new_D8411_ & ~new_D8421_;
  assign new_D8432_ = new_D8453_ | new_D8452_;
  assign new_D8433_ = new_D8399_ | new_D8432_;
  assign new_D8434_ = new_D8457_ | new_D8456_;
  assign new_D8435_ = ~new_D8399_ & new_D8434_;
  assign new_D8436_ = new_D8455_ | new_D8454_;
  assign new_D8437_ = new_D8399_ & new_D8436_;
  assign new_D8438_ = new_D8397_ & ~new_D8407_;
  assign new_D8439_ = ~new_D8397_ & new_D8407_;
  assign new_D8440_ = ~new_D8396_ | ~new_D8421_;
  assign new_D8441_ = new_D8407_ & new_D8440_;
  assign new_D8442_ = ~new_D8407_ & ~new_D8441_;
  assign new_D8443_ = new_D8407_ | new_D8440_;
  assign new_D8444_ = ~new_D8397_ & new_D8398_;
  assign new_D8445_ = new_D8397_ & ~new_D8398_;
  assign new_D8446_ = new_D8414_ | new_D8451_;
  assign new_D8447_ = ~new_D8414_ & ~new_D8450_;
  assign new_D8448_ = new_D8397_ | new_D8414_;
  assign new_D8449_ = new_D8397_ | new_D8398_;
  assign new_D8450_ = new_D8414_ & new_D8451_;
  assign new_D8451_ = ~new_D8396_ | ~new_D8421_;
  assign new_D8452_ = new_D8429_ & new_D8449_;
  assign new_D8453_ = ~new_D8429_ & ~new_D8449_;
  assign new_D8454_ = new_D8458_ | new_D8459_;
  assign new_D8455_ = ~new_D8400_ & new_D8414_;
  assign new_D8456_ = new_D8460_ | new_D8461_;
  assign new_D8457_ = new_D8400_ & new_D8414_;
  assign new_D8458_ = ~new_D8400_ & ~new_D8414_;
  assign new_D8459_ = new_D8400_ & ~new_D8414_;
  assign new_D8460_ = new_D8400_ & ~new_D8414_;
  assign new_D8461_ = ~new_D8400_ & new_D8414_;
  assign new_D8462_ = new_G313_;
  assign new_D8463_ = new_G380_;
  assign new_D8464_ = new_G447_;
  assign new_D8465_ = new_G514_;
  assign new_D8466_ = new_G581_;
  assign new_D8467_ = new_G648_;
  assign new_D8468_ = new_D8475_ & new_D8474_;
  assign new_D8469_ = new_D8477_ | new_D8476_;
  assign new_D8470_ = new_D8479_ | new_D8478_;
  assign new_D8471_ = new_D8481_ & new_D8480_;
  assign new_D8472_ = new_D8481_ & new_D8482_;
  assign new_D8473_ = new_D8474_ | new_D8483_;
  assign new_D8474_ = new_D8463_ | new_D8486_;
  assign new_D8475_ = new_D8485_ | new_D8484_;
  assign new_D8476_ = new_D8490_ & new_D8489_;
  assign new_D8477_ = new_D8488_ & new_D8487_;
  assign new_D8478_ = new_D8493_ | new_D8492_;
  assign new_D8479_ = new_D8488_ & new_D8491_;
  assign new_D8480_ = new_D8463_ | new_D8496_;
  assign new_D8481_ = new_D8495_ | new_D8494_;
  assign new_D8482_ = new_D8498_ | new_D8497_;
  assign new_D8483_ = ~new_D8474_ & new_D8500_;
  assign new_D8484_ = ~new_D8476_ & new_D8488_;
  assign new_D8485_ = new_D8476_ & ~new_D8488_;
  assign new_D8486_ = new_D8462_ & ~new_D8463_;
  assign new_D8487_ = ~new_D8509_ | ~new_D8510_;
  assign new_D8488_ = new_D8502_ | new_D8504_;
  assign new_D8489_ = new_D8512_ | new_D8511_;
  assign new_D8490_ = new_D8506_ | new_D8505_;
  assign new_D8491_ = ~new_D8514_ | ~new_D8513_;
  assign new_D8492_ = ~new_D8515_ & new_D8516_;
  assign new_D8493_ = new_D8515_ & ~new_D8516_;
  assign new_D8494_ = ~new_D8462_ & new_D8463_;
  assign new_D8495_ = new_D8462_ & ~new_D8463_;
  assign new_D8496_ = ~new_D8478_ | new_D8488_;
  assign new_D8497_ = new_D8478_ & new_D8488_;
  assign new_D8498_ = ~new_D8478_ & ~new_D8488_;
  assign new_D8499_ = new_D8520_ | new_D8519_;
  assign new_D8500_ = new_D8466_ | new_D8499_;
  assign new_D8501_ = new_D8524_ | new_D8523_;
  assign new_D8502_ = ~new_D8466_ & new_D8501_;
  assign new_D8503_ = new_D8522_ | new_D8521_;
  assign new_D8504_ = new_D8466_ & new_D8503_;
  assign new_D8505_ = new_D8464_ & ~new_D8474_;
  assign new_D8506_ = ~new_D8464_ & new_D8474_;
  assign new_D8507_ = ~new_D8463_ | ~new_D8488_;
  assign new_D8508_ = new_D8474_ & new_D8507_;
  assign new_D8509_ = ~new_D8474_ & ~new_D8508_;
  assign new_D8510_ = new_D8474_ | new_D8507_;
  assign new_D8511_ = ~new_D8464_ & new_D8465_;
  assign new_D8512_ = new_D8464_ & ~new_D8465_;
  assign new_D8513_ = new_D8481_ | new_D8518_;
  assign new_D8514_ = ~new_D8481_ & ~new_D8517_;
  assign new_D8515_ = new_D8464_ | new_D8481_;
  assign new_D8516_ = new_D8464_ | new_D8465_;
  assign new_D8517_ = new_D8481_ & new_D8518_;
  assign new_D8518_ = ~new_D8463_ | ~new_D8488_;
  assign new_D8519_ = new_D8496_ & new_D8516_;
  assign new_D8520_ = ~new_D8496_ & ~new_D8516_;
  assign new_D8521_ = new_D8525_ | new_D8526_;
  assign new_D8522_ = ~new_D8467_ & new_D8481_;
  assign new_D8523_ = new_D8527_ | new_D8528_;
  assign new_D8524_ = new_D8467_ & new_D8481_;
  assign new_D8525_ = ~new_D8467_ & ~new_D8481_;
  assign new_D8526_ = new_D8467_ & ~new_D8481_;
  assign new_D8527_ = new_D8467_ & ~new_D8481_;
  assign new_D8528_ = ~new_D8467_ & new_D8481_;
  assign new_D8529_ = new_G715_;
  assign new_D8530_ = new_G782_;
  assign new_D8531_ = new_G849_;
  assign new_D8532_ = new_G916_;
  assign new_D8533_ = new_G983_;
  assign new_D8534_ = new_G1050_;
  assign new_D8535_ = new_D8542_ & new_D8541_;
  assign new_D8536_ = new_D8544_ | new_D8543_;
  assign new_D8537_ = new_D8546_ | new_D8545_;
  assign new_D8538_ = new_D8548_ & new_D8547_;
  assign new_D8539_ = new_D8548_ & new_D8549_;
  assign new_D8540_ = new_D8541_ | new_D8550_;
  assign new_D8541_ = new_D8530_ | new_D8553_;
  assign new_D8542_ = new_D8552_ | new_D8551_;
  assign new_D8543_ = new_D8557_ & new_D8556_;
  assign new_D8544_ = new_D8555_ & new_D8554_;
  assign new_D8545_ = new_D8560_ | new_D8559_;
  assign new_D8546_ = new_D8555_ & new_D8558_;
  assign new_D8547_ = new_D8530_ | new_D8563_;
  assign new_D8548_ = new_D8562_ | new_D8561_;
  assign new_D8549_ = new_D8565_ | new_D8564_;
  assign new_D8550_ = ~new_D8541_ & new_D8567_;
  assign new_D8551_ = ~new_D8543_ & new_D8555_;
  assign new_D8552_ = new_D8543_ & ~new_D8555_;
  assign new_D8553_ = new_D8529_ & ~new_D8530_;
  assign new_D8554_ = ~new_D8576_ | ~new_D8577_;
  assign new_D8555_ = new_D8569_ | new_D8571_;
  assign new_D8556_ = new_D8579_ | new_D8578_;
  assign new_D8557_ = new_D8573_ | new_D8572_;
  assign new_D8558_ = ~new_D8581_ | ~new_D8580_;
  assign new_D8559_ = ~new_D8582_ & new_D8583_;
  assign new_D8560_ = new_D8582_ & ~new_D8583_;
  assign new_D8561_ = ~new_D8529_ & new_D8530_;
  assign new_D8562_ = new_D8529_ & ~new_D8530_;
  assign new_D8563_ = ~new_D8545_ | new_D8555_;
  assign new_D8564_ = new_D8545_ & new_D8555_;
  assign new_D8565_ = ~new_D8545_ & ~new_D8555_;
  assign new_D8566_ = new_D8587_ | new_D8586_;
  assign new_D8567_ = new_D8533_ | new_D8566_;
  assign new_D8568_ = new_D8591_ | new_D8590_;
  assign new_D8569_ = ~new_D8533_ & new_D8568_;
  assign new_D8570_ = new_D8589_ | new_D8588_;
  assign new_D8571_ = new_D8533_ & new_D8570_;
  assign new_D8572_ = new_D8531_ & ~new_D8541_;
  assign new_D8573_ = ~new_D8531_ & new_D8541_;
  assign new_D8574_ = ~new_D8530_ | ~new_D8555_;
  assign new_D8575_ = new_D8541_ & new_D8574_;
  assign new_D8576_ = ~new_D8541_ & ~new_D8575_;
  assign new_D8577_ = new_D8541_ | new_D8574_;
  assign new_D8578_ = ~new_D8531_ & new_D8532_;
  assign new_D8579_ = new_D8531_ & ~new_D8532_;
  assign new_D8580_ = new_D8548_ | new_D8585_;
  assign new_D8581_ = ~new_D8548_ & ~new_D8584_;
  assign new_D8582_ = new_D8531_ | new_D8548_;
  assign new_D8583_ = new_D8531_ | new_D8532_;
  assign new_D8584_ = new_D8548_ & new_D8585_;
  assign new_D8585_ = ~new_D8530_ | ~new_D8555_;
  assign new_D8586_ = new_D8563_ & new_D8583_;
  assign new_D8587_ = ~new_D8563_ & ~new_D8583_;
  assign new_D8588_ = new_D8592_ | new_D8593_;
  assign new_D8589_ = ~new_D8534_ & new_D8548_;
  assign new_D8590_ = new_D8594_ | new_D8595_;
  assign new_D8591_ = new_D8534_ & new_D8548_;
  assign new_D8592_ = ~new_D8534_ & ~new_D8548_;
  assign new_D8593_ = new_D8534_ & ~new_D8548_;
  assign new_D8594_ = new_D8534_ & ~new_D8548_;
  assign new_D8595_ = ~new_D8534_ & new_D8548_;
  assign new_D8596_ = new_G1117_;
  assign new_D8597_ = new_G1184_;
  assign new_D8598_ = new_G1251_;
  assign new_D8599_ = new_G1318_;
  assign new_D8600_ = new_G1385_;
  assign new_D8601_ = new_G1452_;
  assign new_D8602_ = new_D8609_ & new_D8608_;
  assign new_D8603_ = new_D8611_ | new_D8610_;
  assign new_D8604_ = new_D8613_ | new_D8612_;
  assign new_D8605_ = new_D8615_ & new_D8614_;
  assign new_D8606_ = new_D8615_ & new_D8616_;
  assign new_D8607_ = new_D8608_ | new_D8617_;
  assign new_D8608_ = new_D8597_ | new_D8620_;
  assign new_D8609_ = new_D8619_ | new_D8618_;
  assign new_D8610_ = new_D8624_ & new_D8623_;
  assign new_D8611_ = new_D8622_ & new_D8621_;
  assign new_D8612_ = new_D8627_ | new_D8626_;
  assign new_D8613_ = new_D8622_ & new_D8625_;
  assign new_D8614_ = new_D8597_ | new_D8630_;
  assign new_D8615_ = new_D8629_ | new_D8628_;
  assign new_D8616_ = new_D8632_ | new_D8631_;
  assign new_D8617_ = ~new_D8608_ & new_D8634_;
  assign new_D8618_ = ~new_D8610_ & new_D8622_;
  assign new_D8619_ = new_D8610_ & ~new_D8622_;
  assign new_D8620_ = new_D8596_ & ~new_D8597_;
  assign new_D8621_ = ~new_D8643_ | ~new_D8644_;
  assign new_D8622_ = new_D8636_ | new_D8638_;
  assign new_D8623_ = new_D8646_ | new_D8645_;
  assign new_D8624_ = new_D8640_ | new_D8639_;
  assign new_D8625_ = ~new_D8648_ | ~new_D8647_;
  assign new_D8626_ = ~new_D8649_ & new_D8650_;
  assign new_D8627_ = new_D8649_ & ~new_D8650_;
  assign new_D8628_ = ~new_D8596_ & new_D8597_;
  assign new_D8629_ = new_D8596_ & ~new_D8597_;
  assign new_D8630_ = ~new_D8612_ | new_D8622_;
  assign new_D8631_ = new_D8612_ & new_D8622_;
  assign new_D8632_ = ~new_D8612_ & ~new_D8622_;
  assign new_D8633_ = new_D8654_ | new_D8653_;
  assign new_D8634_ = new_D8600_ | new_D8633_;
  assign new_D8635_ = new_D8658_ | new_D8657_;
  assign new_D8636_ = ~new_D8600_ & new_D8635_;
  assign new_D8637_ = new_D8656_ | new_D8655_;
  assign new_D8638_ = new_D8600_ & new_D8637_;
  assign new_D8639_ = new_D8598_ & ~new_D8608_;
  assign new_D8640_ = ~new_D8598_ & new_D8608_;
  assign new_D8641_ = ~new_D8597_ | ~new_D8622_;
  assign new_D8642_ = new_D8608_ & new_D8641_;
  assign new_D8643_ = ~new_D8608_ & ~new_D8642_;
  assign new_D8644_ = new_D8608_ | new_D8641_;
  assign new_D8645_ = ~new_D8598_ & new_D8599_;
  assign new_D8646_ = new_D8598_ & ~new_D8599_;
  assign new_D8647_ = new_D8615_ | new_D8652_;
  assign new_D8648_ = ~new_D8615_ & ~new_D8651_;
  assign new_D8649_ = new_D8598_ | new_D8615_;
  assign new_D8650_ = new_D8598_ | new_D8599_;
  assign new_D8651_ = new_D8615_ & new_D8652_;
  assign new_D8652_ = ~new_D8597_ | ~new_D8622_;
  assign new_D8653_ = new_D8630_ & new_D8650_;
  assign new_D8654_ = ~new_D8630_ & ~new_D8650_;
  assign new_D8655_ = new_D8659_ | new_D8660_;
  assign new_D8656_ = ~new_D8601_ & new_D8615_;
  assign new_D8657_ = new_D8661_ | new_D8662_;
  assign new_D8658_ = new_D8601_ & new_D8615_;
  assign new_D8659_ = ~new_D8601_ & ~new_D8615_;
  assign new_D8660_ = new_D8601_ & ~new_D8615_;
  assign new_D8661_ = new_D8601_ & ~new_D8615_;
  assign new_D8662_ = ~new_D8601_ & new_D8615_;
  assign new_D8663_ = new_G1519_;
  assign new_D8664_ = new_G1586_;
  assign new_D8665_ = new_G1653_;
  assign new_D8666_ = new_G1720_;
  assign new_D8667_ = new_G1787_;
  assign new_D8668_ = new_G1854_;
  assign new_D8669_ = new_D8676_ & new_D8675_;
  assign new_D8670_ = new_D8678_ | new_D8677_;
  assign new_D8671_ = new_D8680_ | new_D8679_;
  assign new_D8672_ = new_D8682_ & new_D8681_;
  assign new_D8673_ = new_D8682_ & new_D8683_;
  assign new_D8674_ = new_D8675_ | new_D8684_;
  assign new_D8675_ = new_D8664_ | new_D8687_;
  assign new_D8676_ = new_D8686_ | new_D8685_;
  assign new_D8677_ = new_D8691_ & new_D8690_;
  assign new_D8678_ = new_D8689_ & new_D8688_;
  assign new_D8679_ = new_D8694_ | new_D8693_;
  assign new_D8680_ = new_D8689_ & new_D8692_;
  assign new_D8681_ = new_D8664_ | new_D8697_;
  assign new_D8682_ = new_D8696_ | new_D8695_;
  assign new_D8683_ = new_D8699_ | new_D8698_;
  assign new_D8684_ = ~new_D8675_ & new_D8701_;
  assign new_D8685_ = ~new_D8677_ & new_D8689_;
  assign new_D8686_ = new_D8677_ & ~new_D8689_;
  assign new_D8687_ = new_D8663_ & ~new_D8664_;
  assign new_D8688_ = ~new_D8710_ | ~new_D8711_;
  assign new_D8689_ = new_D8703_ | new_D8705_;
  assign new_D8690_ = new_D8713_ | new_D8712_;
  assign new_D8691_ = new_D8707_ | new_D8706_;
  assign new_D8692_ = ~new_D8715_ | ~new_D8714_;
  assign new_D8693_ = ~new_D8716_ & new_D8717_;
  assign new_D8694_ = new_D8716_ & ~new_D8717_;
  assign new_D8695_ = ~new_D8663_ & new_D8664_;
  assign new_D8696_ = new_D8663_ & ~new_D8664_;
  assign new_D8697_ = ~new_D8679_ | new_D8689_;
  assign new_D8698_ = new_D8679_ & new_D8689_;
  assign new_D8699_ = ~new_D8679_ & ~new_D8689_;
  assign new_D8700_ = new_D8721_ | new_D8720_;
  assign new_D8701_ = new_D8667_ | new_D8700_;
  assign new_D8702_ = new_D8725_ | new_D8724_;
  assign new_D8703_ = ~new_D8667_ & new_D8702_;
  assign new_D8704_ = new_D8723_ | new_D8722_;
  assign new_D8705_ = new_D8667_ & new_D8704_;
  assign new_D8706_ = new_D8665_ & ~new_D8675_;
  assign new_D8707_ = ~new_D8665_ & new_D8675_;
  assign new_D8708_ = ~new_D8664_ | ~new_D8689_;
  assign new_D8709_ = new_D8675_ & new_D8708_;
  assign new_D8710_ = ~new_D8675_ & ~new_D8709_;
  assign new_D8711_ = new_D8675_ | new_D8708_;
  assign new_D8712_ = ~new_D8665_ & new_D8666_;
  assign new_D8713_ = new_D8665_ & ~new_D8666_;
  assign new_D8714_ = new_D8682_ | new_D8719_;
  assign new_D8715_ = ~new_D8682_ & ~new_D8718_;
  assign new_D8716_ = new_D8665_ | new_D8682_;
  assign new_D8717_ = new_D8665_ | new_D8666_;
  assign new_D8718_ = new_D8682_ & new_D8719_;
  assign new_D8719_ = ~new_D8664_ | ~new_D8689_;
  assign new_D8720_ = new_D8697_ & new_D8717_;
  assign new_D8721_ = ~new_D8697_ & ~new_D8717_;
  assign new_D8722_ = new_D8726_ | new_D8727_;
  assign new_D8723_ = ~new_D8668_ & new_D8682_;
  assign new_D8724_ = new_D8728_ | new_D8729_;
  assign new_D8725_ = new_D8668_ & new_D8682_;
  assign new_D8726_ = ~new_D8668_ & ~new_D8682_;
  assign new_D8727_ = new_D8668_ & ~new_D8682_;
  assign new_D8728_ = new_D8668_ & ~new_D8682_;
  assign new_D8729_ = ~new_D8668_ & new_D8682_;
  assign new_D8730_ = new_G1921_;
  assign new_D8731_ = new_G1988_;
  assign new_D8732_ = new_G2055_;
  assign new_D8733_ = new_G2122_;
  assign new_D8734_ = new_G2189_;
  assign new_D8735_ = new_G2256_;
  assign new_D8736_ = new_D8743_ & new_D8742_;
  assign new_D8737_ = new_D8745_ | new_D8744_;
  assign new_D8738_ = new_D8747_ | new_D8746_;
  assign new_D8739_ = new_D8749_ & new_D8748_;
  assign new_D8740_ = new_D8749_ & new_D8750_;
  assign new_D8741_ = new_D8742_ | new_D8751_;
  assign new_D8742_ = new_D8731_ | new_D8754_;
  assign new_D8743_ = new_D8753_ | new_D8752_;
  assign new_D8744_ = new_D8758_ & new_D8757_;
  assign new_D8745_ = new_D8756_ & new_D8755_;
  assign new_D8746_ = new_D8761_ | new_D8760_;
  assign new_D8747_ = new_D8756_ & new_D8759_;
  assign new_D8748_ = new_D8731_ | new_D8764_;
  assign new_D8749_ = new_D8763_ | new_D8762_;
  assign new_D8750_ = new_D8766_ | new_D8765_;
  assign new_D8751_ = ~new_D8742_ & new_D8768_;
  assign new_D8752_ = ~new_D8744_ & new_D8756_;
  assign new_D8753_ = new_D8744_ & ~new_D8756_;
  assign new_D8754_ = new_D8730_ & ~new_D8731_;
  assign new_D8755_ = ~new_D8777_ | ~new_D8778_;
  assign new_D8756_ = new_D8770_ | new_D8772_;
  assign new_D8757_ = new_D8780_ | new_D8779_;
  assign new_D8758_ = new_D8774_ | new_D8773_;
  assign new_D8759_ = ~new_D8782_ | ~new_D8781_;
  assign new_D8760_ = ~new_D8783_ & new_D8784_;
  assign new_D8761_ = new_D8783_ & ~new_D8784_;
  assign new_D8762_ = ~new_D8730_ & new_D8731_;
  assign new_D8763_ = new_D8730_ & ~new_D8731_;
  assign new_D8764_ = ~new_D8746_ | new_D8756_;
  assign new_D8765_ = new_D8746_ & new_D8756_;
  assign new_D8766_ = ~new_D8746_ & ~new_D8756_;
  assign new_D8767_ = new_D8788_ | new_D8787_;
  assign new_D8768_ = new_D8734_ | new_D8767_;
  assign new_D8769_ = new_D8792_ | new_D8791_;
  assign new_D8770_ = ~new_D8734_ & new_D8769_;
  assign new_D8771_ = new_D8790_ | new_D8789_;
  assign new_D8772_ = new_D8734_ & new_D8771_;
  assign new_D8773_ = new_D8732_ & ~new_D8742_;
  assign new_D8774_ = ~new_D8732_ & new_D8742_;
  assign new_D8775_ = ~new_D8731_ | ~new_D8756_;
  assign new_D8776_ = new_D8742_ & new_D8775_;
  assign new_D8777_ = ~new_D8742_ & ~new_D8776_;
  assign new_D8778_ = new_D8742_ | new_D8775_;
  assign new_D8779_ = ~new_D8732_ & new_D8733_;
  assign new_D8780_ = new_D8732_ & ~new_D8733_;
  assign new_D8781_ = new_D8749_ | new_D8786_;
  assign new_D8782_ = ~new_D8749_ & ~new_D8785_;
  assign new_D8783_ = new_D8732_ | new_D8749_;
  assign new_D8784_ = new_D8732_ | new_D8733_;
  assign new_D8785_ = new_D8749_ & new_D8786_;
  assign new_D8786_ = ~new_D8731_ | ~new_D8756_;
  assign new_D8787_ = new_D8764_ & new_D8784_;
  assign new_D8788_ = ~new_D8764_ & ~new_D8784_;
  assign new_D8789_ = new_D8793_ | new_D8794_;
  assign new_D8790_ = ~new_D8735_ & new_D8749_;
  assign new_D8791_ = new_D8795_ | new_D8796_;
  assign new_D8792_ = new_D8735_ & new_D8749_;
  assign new_D8793_ = ~new_D8735_ & ~new_D8749_;
  assign new_D8794_ = new_D8735_ & ~new_D8749_;
  assign new_D8795_ = new_D8735_ & ~new_D8749_;
  assign new_D8796_ = ~new_D8735_ & new_D8749_;
  assign new_D8797_ = new_G2323_;
  assign new_D8798_ = new_G2390_;
  assign new_D8799_ = new_G2457_;
  assign new_D8800_ = new_G2524_;
  assign new_D8801_ = new_G2591_;
  assign new_D8802_ = new_G2658_;
  assign new_D8803_ = new_D8810_ & new_D8809_;
  assign new_D8804_ = new_D8812_ | new_D8811_;
  assign new_D8805_ = new_D8814_ | new_D8813_;
  assign new_D8806_ = new_D8816_ & new_D8815_;
  assign new_D8807_ = new_D8816_ & new_D8817_;
  assign new_D8808_ = new_D8809_ | new_D8818_;
  assign new_D8809_ = new_D8798_ | new_D8821_;
  assign new_D8810_ = new_D8820_ | new_D8819_;
  assign new_D8811_ = new_D8825_ & new_D8824_;
  assign new_D8812_ = new_D8823_ & new_D8822_;
  assign new_D8813_ = new_D8828_ | new_D8827_;
  assign new_D8814_ = new_D8823_ & new_D8826_;
  assign new_D8815_ = new_D8798_ | new_D8831_;
  assign new_D8816_ = new_D8830_ | new_D8829_;
  assign new_D8817_ = new_D8833_ | new_D8832_;
  assign new_D8818_ = ~new_D8809_ & new_D8835_;
  assign new_D8819_ = ~new_D8811_ & new_D8823_;
  assign new_D8820_ = new_D8811_ & ~new_D8823_;
  assign new_D8821_ = new_D8797_ & ~new_D8798_;
  assign new_D8822_ = ~new_D8844_ | ~new_D8845_;
  assign new_D8823_ = new_D8837_ | new_D8839_;
  assign new_D8824_ = new_D8847_ | new_D8846_;
  assign new_D8825_ = new_D8841_ | new_D8840_;
  assign new_D8826_ = ~new_D8849_ | ~new_D8848_;
  assign new_D8827_ = ~new_D8850_ & new_D8851_;
  assign new_D8828_ = new_D8850_ & ~new_D8851_;
  assign new_D8829_ = ~new_D8797_ & new_D8798_;
  assign new_D8830_ = new_D8797_ & ~new_D8798_;
  assign new_D8831_ = ~new_D8813_ | new_D8823_;
  assign new_D8832_ = new_D8813_ & new_D8823_;
  assign new_D8833_ = ~new_D8813_ & ~new_D8823_;
  assign new_D8834_ = new_D8855_ | new_D8854_;
  assign new_D8835_ = new_D8801_ | new_D8834_;
  assign new_D8836_ = new_D8859_ | new_D8858_;
  assign new_D8837_ = ~new_D8801_ & new_D8836_;
  assign new_D8838_ = new_D8857_ | new_D8856_;
  assign new_D8839_ = new_D8801_ & new_D8838_;
  assign new_D8840_ = new_D8799_ & ~new_D8809_;
  assign new_D8841_ = ~new_D8799_ & new_D8809_;
  assign new_D8842_ = ~new_D8798_ | ~new_D8823_;
  assign new_D8843_ = new_D8809_ & new_D8842_;
  assign new_D8844_ = ~new_D8809_ & ~new_D8843_;
  assign new_D8845_ = new_D8809_ | new_D8842_;
  assign new_D8846_ = ~new_D8799_ & new_D8800_;
  assign new_D8847_ = new_D8799_ & ~new_D8800_;
  assign new_D8848_ = new_D8816_ | new_D8853_;
  assign new_D8849_ = ~new_D8816_ & ~new_D8852_;
  assign new_D8850_ = new_D8799_ | new_D8816_;
  assign new_D8851_ = new_D8799_ | new_D8800_;
  assign new_D8852_ = new_D8816_ & new_D8853_;
  assign new_D8853_ = ~new_D8798_ | ~new_D8823_;
  assign new_D8854_ = new_D8831_ & new_D8851_;
  assign new_D8855_ = ~new_D8831_ & ~new_D8851_;
  assign new_D8856_ = new_D8860_ | new_D8861_;
  assign new_D8857_ = ~new_D8802_ & new_D8816_;
  assign new_D8858_ = new_D8862_ | new_D8863_;
  assign new_D8859_ = new_D8802_ & new_D8816_;
  assign new_D8860_ = ~new_D8802_ & ~new_D8816_;
  assign new_D8861_ = new_D8802_ & ~new_D8816_;
  assign new_D8862_ = new_D8802_ & ~new_D8816_;
  assign new_D8863_ = ~new_D8802_ & new_D8816_;
  assign new_D8864_ = new_G2725_;
  assign new_D8865_ = new_G2792_;
  assign new_D8866_ = new_G2859_;
  assign new_D8867_ = new_G2926_;
  assign new_D8868_ = new_G2993_;
  assign new_D8869_ = new_G3060_;
  assign new_D8870_ = new_D8877_ & new_D8876_;
  assign new_D8871_ = new_D8879_ | new_D8878_;
  assign new_D8872_ = new_D8881_ | new_D8880_;
  assign new_D8873_ = new_D8883_ & new_D8882_;
  assign new_D8874_ = new_D8883_ & new_D8884_;
  assign new_D8875_ = new_D8876_ | new_D8885_;
  assign new_D8876_ = new_D8865_ | new_D8888_;
  assign new_D8877_ = new_D8887_ | new_D8886_;
  assign new_D8878_ = new_D8892_ & new_D8891_;
  assign new_D8879_ = new_D8890_ & new_D8889_;
  assign new_D8880_ = new_D8895_ | new_D8894_;
  assign new_D8881_ = new_D8890_ & new_D8893_;
  assign new_D8882_ = new_D8865_ | new_D8898_;
  assign new_D8883_ = new_D8897_ | new_D8896_;
  assign new_D8884_ = new_D8900_ | new_D8899_;
  assign new_D8885_ = ~new_D8876_ & new_D8902_;
  assign new_D8886_ = ~new_D8878_ & new_D8890_;
  assign new_D8887_ = new_D8878_ & ~new_D8890_;
  assign new_D8888_ = new_D8864_ & ~new_D8865_;
  assign new_D8889_ = ~new_D8911_ | ~new_D8912_;
  assign new_D8890_ = new_D8904_ | new_D8906_;
  assign new_D8891_ = new_D8914_ | new_D8913_;
  assign new_D8892_ = new_D8908_ | new_D8907_;
  assign new_D8893_ = ~new_D8916_ | ~new_D8915_;
  assign new_D8894_ = ~new_D8917_ & new_D8918_;
  assign new_D8895_ = new_D8917_ & ~new_D8918_;
  assign new_D8896_ = ~new_D8864_ & new_D8865_;
  assign new_D8897_ = new_D8864_ & ~new_D8865_;
  assign new_D8898_ = ~new_D8880_ | new_D8890_;
  assign new_D8899_ = new_D8880_ & new_D8890_;
  assign new_D8900_ = ~new_D8880_ & ~new_D8890_;
  assign new_D8901_ = new_D8922_ | new_D8921_;
  assign new_D8902_ = new_D8868_ | new_D8901_;
  assign new_D8903_ = new_D8926_ | new_D8925_;
  assign new_D8904_ = ~new_D8868_ & new_D8903_;
  assign new_D8905_ = new_D8924_ | new_D8923_;
  assign new_D8906_ = new_D8868_ & new_D8905_;
  assign new_D8907_ = new_D8866_ & ~new_D8876_;
  assign new_D8908_ = ~new_D8866_ & new_D8876_;
  assign new_D8909_ = ~new_D8865_ | ~new_D8890_;
  assign new_D8910_ = new_D8876_ & new_D8909_;
  assign new_D8911_ = ~new_D8876_ & ~new_D8910_;
  assign new_D8912_ = new_D8876_ | new_D8909_;
  assign new_D8913_ = ~new_D8866_ & new_D8867_;
  assign new_D8914_ = new_D8866_ & ~new_D8867_;
  assign new_D8915_ = new_D8883_ | new_D8920_;
  assign new_D8916_ = ~new_D8883_ & ~new_D8919_;
  assign new_D8917_ = new_D8866_ | new_D8883_;
  assign new_D8918_ = new_D8866_ | new_D8867_;
  assign new_D8919_ = new_D8883_ & new_D8920_;
  assign new_D8920_ = ~new_D8865_ | ~new_D8890_;
  assign new_D8921_ = new_D8898_ & new_D8918_;
  assign new_D8922_ = ~new_D8898_ & ~new_D8918_;
  assign new_D8923_ = new_D8927_ | new_D8928_;
  assign new_D8924_ = ~new_D8869_ & new_D8883_;
  assign new_D8925_ = new_D8929_ | new_D8930_;
  assign new_D8926_ = new_D8869_ & new_D8883_;
  assign new_D8927_ = ~new_D8869_ & ~new_D8883_;
  assign new_D8928_ = new_D8869_ & ~new_D8883_;
  assign new_D8929_ = new_D8869_ & ~new_D8883_;
  assign new_D8930_ = ~new_D8869_ & new_D8883_;
  assign new_D8931_ = new_G3127_;
  assign new_D8932_ = new_G3194_;
  assign new_D8933_ = new_G3261_;
  assign new_D8934_ = new_G3328_;
  assign new_D8935_ = new_G3395_;
  assign new_D8936_ = new_G3462_;
  assign new_D8937_ = new_D8944_ & new_D8943_;
  assign new_D8938_ = new_D8946_ | new_D8945_;
  assign new_D8939_ = new_D8948_ | new_D8947_;
  assign new_D8940_ = new_D8950_ & new_D8949_;
  assign new_D8941_ = new_D8950_ & new_D8951_;
  assign new_D8942_ = new_D8943_ | new_D8952_;
  assign new_D8943_ = new_D8932_ | new_D8955_;
  assign new_D8944_ = new_D8954_ | new_D8953_;
  assign new_D8945_ = new_D8959_ & new_D8958_;
  assign new_D8946_ = new_D8957_ & new_D8956_;
  assign new_D8947_ = new_D8962_ | new_D8961_;
  assign new_D8948_ = new_D8957_ & new_D8960_;
  assign new_D8949_ = new_D8932_ | new_D8965_;
  assign new_D8950_ = new_D8964_ | new_D8963_;
  assign new_D8951_ = new_D8967_ | new_D8966_;
  assign new_D8952_ = ~new_D8943_ & new_D8969_;
  assign new_D8953_ = ~new_D8945_ & new_D8957_;
  assign new_D8954_ = new_D8945_ & ~new_D8957_;
  assign new_D8955_ = new_D8931_ & ~new_D8932_;
  assign new_D8956_ = ~new_D8978_ | ~new_D8979_;
  assign new_D8957_ = new_D8971_ | new_D8973_;
  assign new_D8958_ = new_D8981_ | new_D8980_;
  assign new_D8959_ = new_D8975_ | new_D8974_;
  assign new_D8960_ = ~new_D8983_ | ~new_D8982_;
  assign new_D8961_ = ~new_D8984_ & new_D8985_;
  assign new_D8962_ = new_D8984_ & ~new_D8985_;
  assign new_D8963_ = ~new_D8931_ & new_D8932_;
  assign new_D8964_ = new_D8931_ & ~new_D8932_;
  assign new_D8965_ = ~new_D8947_ | new_D8957_;
  assign new_D8966_ = new_D8947_ & new_D8957_;
  assign new_D8967_ = ~new_D8947_ & ~new_D8957_;
  assign new_D8968_ = new_D8989_ | new_D8988_;
  assign new_D8969_ = new_D8935_ | new_D8968_;
  assign new_D8970_ = new_D8993_ | new_D8992_;
  assign new_D8971_ = ~new_D8935_ & new_D8970_;
  assign new_D8972_ = new_D8991_ | new_D8990_;
  assign new_D8973_ = new_D8935_ & new_D8972_;
  assign new_D8974_ = new_D8933_ & ~new_D8943_;
  assign new_D8975_ = ~new_D8933_ & new_D8943_;
  assign new_D8976_ = ~new_D8932_ | ~new_D8957_;
  assign new_D8977_ = new_D8943_ & new_D8976_;
  assign new_D8978_ = ~new_D8943_ & ~new_D8977_;
  assign new_D8979_ = new_D8943_ | new_D8976_;
  assign new_D8980_ = ~new_D8933_ & new_D8934_;
  assign new_D8981_ = new_D8933_ & ~new_D8934_;
  assign new_D8982_ = new_D8950_ | new_D8987_;
  assign new_D8983_ = ~new_D8950_ & ~new_D8986_;
  assign new_D8984_ = new_D8933_ | new_D8950_;
  assign new_D8985_ = new_D8933_ | new_D8934_;
  assign new_D8986_ = new_D8950_ & new_D8987_;
  assign new_D8987_ = ~new_D8932_ | ~new_D8957_;
  assign new_D8988_ = new_D8965_ & new_D8985_;
  assign new_D8989_ = ~new_D8965_ & ~new_D8985_;
  assign new_D8990_ = new_D8994_ | new_D8995_;
  assign new_D8991_ = ~new_D8936_ & new_D8950_;
  assign new_D8992_ = new_D8996_ | new_D8997_;
  assign new_D8993_ = new_D8936_ & new_D8950_;
  assign new_D8994_ = ~new_D8936_ & ~new_D8950_;
  assign new_D8995_ = new_D8936_ & ~new_D8950_;
  assign new_D8996_ = new_D8936_ & ~new_D8950_;
  assign new_D8997_ = ~new_D8936_ & new_D8950_;
  assign new_D8998_ = new_G3529_;
  assign new_D8999_ = new_G3596_;
  assign new_D9000_ = new_G3663_;
  assign new_D9001_ = new_G3730_;
  assign new_D9002_ = new_G3797_;
  assign new_D9003_ = new_G3864_;
  assign new_D9004_ = new_D9011_ & new_D9010_;
  assign new_D9005_ = new_D9013_ | new_D9012_;
  assign new_D9006_ = new_D9015_ | new_D9014_;
  assign new_D9007_ = new_D9017_ & new_D9016_;
  assign new_D9008_ = new_D9017_ & new_D9018_;
  assign new_D9009_ = new_D9010_ | new_D9019_;
  assign new_D9010_ = new_D8999_ | new_D9022_;
  assign new_D9011_ = new_D9021_ | new_D9020_;
  assign new_D9012_ = new_D9026_ & new_D9025_;
  assign new_D9013_ = new_D9024_ & new_D9023_;
  assign new_D9014_ = new_D9029_ | new_D9028_;
  assign new_D9015_ = new_D9024_ & new_D9027_;
  assign new_D9016_ = new_D8999_ | new_D9032_;
  assign new_D9017_ = new_D9031_ | new_D9030_;
  assign new_D9018_ = new_D9034_ | new_D9033_;
  assign new_D9019_ = ~new_D9010_ & new_D9036_;
  assign new_D9020_ = ~new_D9012_ & new_D9024_;
  assign new_D9021_ = new_D9012_ & ~new_D9024_;
  assign new_D9022_ = new_D8998_ & ~new_D8999_;
  assign new_D9023_ = ~new_D9045_ | ~new_D9046_;
  assign new_D9024_ = new_D9038_ | new_D9040_;
  assign new_D9025_ = new_D9048_ | new_D9047_;
  assign new_D9026_ = new_D9042_ | new_D9041_;
  assign new_D9027_ = ~new_D9050_ | ~new_D9049_;
  assign new_D9028_ = ~new_D9051_ & new_D9052_;
  assign new_D9029_ = new_D9051_ & ~new_D9052_;
  assign new_D9030_ = ~new_D8998_ & new_D8999_;
  assign new_D9031_ = new_D8998_ & ~new_D8999_;
  assign new_D9032_ = ~new_D9014_ | new_D9024_;
  assign new_D9033_ = new_D9014_ & new_D9024_;
  assign new_D9034_ = ~new_D9014_ & ~new_D9024_;
  assign new_D9035_ = new_D9056_ | new_D9055_;
  assign new_D9036_ = new_D9002_ | new_D9035_;
  assign new_D9037_ = new_D9060_ | new_D9059_;
  assign new_D9038_ = ~new_D9002_ & new_D9037_;
  assign new_D9039_ = new_D9058_ | new_D9057_;
  assign new_D9040_ = new_D9002_ & new_D9039_;
  assign new_D9041_ = new_D9000_ & ~new_D9010_;
  assign new_D9042_ = ~new_D9000_ & new_D9010_;
  assign new_D9043_ = ~new_D8999_ | ~new_D9024_;
  assign new_D9044_ = new_D9010_ & new_D9043_;
  assign new_D9045_ = ~new_D9010_ & ~new_D9044_;
  assign new_D9046_ = new_D9010_ | new_D9043_;
  assign new_D9047_ = ~new_D9000_ & new_D9001_;
  assign new_D9048_ = new_D9000_ & ~new_D9001_;
  assign new_D9049_ = new_D9017_ | new_D9054_;
  assign new_D9050_ = ~new_D9017_ & ~new_D9053_;
  assign new_D9051_ = new_D9000_ | new_D9017_;
  assign new_D9052_ = new_D9000_ | new_D9001_;
  assign new_D9053_ = new_D9017_ & new_D9054_;
  assign new_D9054_ = ~new_D8999_ | ~new_D9024_;
  assign new_D9055_ = new_D9032_ & new_D9052_;
  assign new_D9056_ = ~new_D9032_ & ~new_D9052_;
  assign new_D9057_ = new_D9061_ | new_D9062_;
  assign new_D9058_ = ~new_D9003_ & new_D9017_;
  assign new_D9059_ = new_D9063_ | new_D9064_;
  assign new_D9060_ = new_D9003_ & new_D9017_;
  assign new_D9061_ = ~new_D9003_ & ~new_D9017_;
  assign new_D9062_ = new_D9003_ & ~new_D9017_;
  assign new_D9063_ = new_D9003_ & ~new_D9017_;
  assign new_D9064_ = ~new_D9003_ & new_D9017_;
  assign new_D9065_ = new_G3931_;
  assign new_D9066_ = new_G3998_;
  assign new_D9067_ = new_G4065_;
  assign new_D9068_ = new_G4132_;
  assign new_D9069_ = new_G4199_;
  assign new_D9070_ = new_G4266_;
  assign new_D9071_ = new_D9078_ & new_D9077_;
  assign new_D9072_ = new_D9080_ | new_D9079_;
  assign new_D9073_ = new_D9082_ | new_D9081_;
  assign new_D9074_ = new_D9084_ & new_D9083_;
  assign new_D9075_ = new_D9084_ & new_D9085_;
  assign new_D9076_ = new_D9077_ | new_D9086_;
  assign new_D9077_ = new_D9066_ | new_D9089_;
  assign new_D9078_ = new_D9088_ | new_D9087_;
  assign new_D9079_ = new_D9093_ & new_D9092_;
  assign new_D9080_ = new_D9091_ & new_D9090_;
  assign new_D9081_ = new_D9096_ | new_D9095_;
  assign new_D9082_ = new_D9091_ & new_D9094_;
  assign new_D9083_ = new_D9066_ | new_D9099_;
  assign new_D9084_ = new_D9098_ | new_D9097_;
  assign new_D9085_ = new_D9101_ | new_D9100_;
  assign new_D9086_ = ~new_D9077_ & new_D9103_;
  assign new_D9087_ = ~new_D9079_ & new_D9091_;
  assign new_D9088_ = new_D9079_ & ~new_D9091_;
  assign new_D9089_ = new_D9065_ & ~new_D9066_;
  assign new_D9090_ = ~new_D9112_ | ~new_D9113_;
  assign new_D9091_ = new_D9105_ | new_D9107_;
  assign new_D9092_ = new_D9115_ | new_D9114_;
  assign new_D9093_ = new_D9109_ | new_D9108_;
  assign new_D9094_ = ~new_D9117_ | ~new_D9116_;
  assign new_D9095_ = ~new_D9118_ & new_D9119_;
  assign new_D9096_ = new_D9118_ & ~new_D9119_;
  assign new_D9097_ = ~new_D9065_ & new_D9066_;
  assign new_D9098_ = new_D9065_ & ~new_D9066_;
  assign new_D9099_ = ~new_D9081_ | new_D9091_;
  assign new_D9100_ = new_D9081_ & new_D9091_;
  assign new_D9101_ = ~new_D9081_ & ~new_D9091_;
  assign new_D9102_ = new_D9123_ | new_D9122_;
  assign new_D9103_ = new_D9069_ | new_D9102_;
  assign new_D9104_ = new_D9127_ | new_D9126_;
  assign new_D9105_ = ~new_D9069_ & new_D9104_;
  assign new_D9106_ = new_D9125_ | new_D9124_;
  assign new_D9107_ = new_D9069_ & new_D9106_;
  assign new_D9108_ = new_D9067_ & ~new_D9077_;
  assign new_D9109_ = ~new_D9067_ & new_D9077_;
  assign new_D9110_ = ~new_D9066_ | ~new_D9091_;
  assign new_D9111_ = new_D9077_ & new_D9110_;
  assign new_D9112_ = ~new_D9077_ & ~new_D9111_;
  assign new_D9113_ = new_D9077_ | new_D9110_;
  assign new_D9114_ = ~new_D9067_ & new_D9068_;
  assign new_D9115_ = new_D9067_ & ~new_D9068_;
  assign new_D9116_ = new_D9084_ | new_D9121_;
  assign new_D9117_ = ~new_D9084_ & ~new_D9120_;
  assign new_D9118_ = new_D9067_ | new_D9084_;
  assign new_D9119_ = new_D9067_ | new_D9068_;
  assign new_D9120_ = new_D9084_ & new_D9121_;
  assign new_D9121_ = ~new_D9066_ | ~new_D9091_;
  assign new_D9122_ = new_D9099_ & new_D9119_;
  assign new_D9123_ = ~new_D9099_ & ~new_D9119_;
  assign new_D9124_ = new_D9128_ | new_D9129_;
  assign new_D9125_ = ~new_D9070_ & new_D9084_;
  assign new_D9126_ = new_D9130_ | new_D9131_;
  assign new_D9127_ = new_D9070_ & new_D9084_;
  assign new_D9128_ = ~new_D9070_ & ~new_D9084_;
  assign new_D9129_ = new_D9070_ & ~new_D9084_;
  assign new_D9130_ = new_D9070_ & ~new_D9084_;
  assign new_D9131_ = ~new_D9070_ & new_D9084_;
  assign new_D9132_ = new_G4333_;
  assign new_D9133_ = new_G4400_;
  assign new_D9134_ = new_G4467_;
  assign new_D9135_ = new_G4534_;
  assign new_D9136_ = new_G4601_;
  assign new_D9137_ = new_G4668_;
  assign new_D9138_ = new_D9145_ & new_D9144_;
  assign new_D9139_ = new_D9147_ | new_D9146_;
  assign new_D9140_ = new_D9149_ | new_D9148_;
  assign new_D9141_ = new_D9151_ & new_D9150_;
  assign new_D9142_ = new_D9151_ & new_D9152_;
  assign new_D9143_ = new_D9144_ | new_D9153_;
  assign new_D9144_ = new_D9133_ | new_D9156_;
  assign new_D9145_ = new_D9155_ | new_D9154_;
  assign new_D9146_ = new_D9160_ & new_D9159_;
  assign new_D9147_ = new_D9158_ & new_D9157_;
  assign new_D9148_ = new_D9163_ | new_D9162_;
  assign new_D9149_ = new_D9158_ & new_D9161_;
  assign new_D9150_ = new_D9133_ | new_D9166_;
  assign new_D9151_ = new_D9165_ | new_D9164_;
  assign new_D9152_ = new_D9168_ | new_D9167_;
  assign new_D9153_ = ~new_D9144_ & new_D9170_;
  assign new_D9154_ = ~new_D9146_ & new_D9158_;
  assign new_D9155_ = new_D9146_ & ~new_D9158_;
  assign new_D9156_ = new_D9132_ & ~new_D9133_;
  assign new_D9157_ = ~new_D9179_ | ~new_D9180_;
  assign new_D9158_ = new_D9172_ | new_D9174_;
  assign new_D9159_ = new_D9182_ | new_D9181_;
  assign new_D9160_ = new_D9176_ | new_D9175_;
  assign new_D9161_ = ~new_D9184_ | ~new_D9183_;
  assign new_D9162_ = ~new_D9185_ & new_D9186_;
  assign new_D9163_ = new_D9185_ & ~new_D9186_;
  assign new_D9164_ = ~new_D9132_ & new_D9133_;
  assign new_D9165_ = new_D9132_ & ~new_D9133_;
  assign new_D9166_ = ~new_D9148_ | new_D9158_;
  assign new_D9167_ = new_D9148_ & new_D9158_;
  assign new_D9168_ = ~new_D9148_ & ~new_D9158_;
  assign new_D9169_ = new_D9190_ | new_D9189_;
  assign new_D9170_ = new_D9136_ | new_D9169_;
  assign new_D9171_ = new_D9194_ | new_D9193_;
  assign new_D9172_ = ~new_D9136_ & new_D9171_;
  assign new_D9173_ = new_D9192_ | new_D9191_;
  assign new_D9174_ = new_D9136_ & new_D9173_;
  assign new_D9175_ = new_D9134_ & ~new_D9144_;
  assign new_D9176_ = ~new_D9134_ & new_D9144_;
  assign new_D9177_ = ~new_D9133_ | ~new_D9158_;
  assign new_D9178_ = new_D9144_ & new_D9177_;
  assign new_D9179_ = ~new_D9144_ & ~new_D9178_;
  assign new_D9180_ = new_D9144_ | new_D9177_;
  assign new_D9181_ = ~new_D9134_ & new_D9135_;
  assign new_D9182_ = new_D9134_ & ~new_D9135_;
  assign new_D9183_ = new_D9151_ | new_D9188_;
  assign new_D9184_ = ~new_D9151_ & ~new_D9187_;
  assign new_D9185_ = new_D9134_ | new_D9151_;
  assign new_D9186_ = new_D9134_ | new_D9135_;
  assign new_D9187_ = new_D9151_ & new_D9188_;
  assign new_D9188_ = ~new_D9133_ | ~new_D9158_;
  assign new_D9189_ = new_D9166_ & new_D9186_;
  assign new_D9190_ = ~new_D9166_ & ~new_D9186_;
  assign new_D9191_ = new_D9195_ | new_D9196_;
  assign new_D9192_ = ~new_D9137_ & new_D9151_;
  assign new_D9193_ = new_D9197_ | new_D9198_;
  assign new_D9194_ = new_D9137_ & new_D9151_;
  assign new_D9195_ = ~new_D9137_ & ~new_D9151_;
  assign new_D9196_ = new_D9137_ & ~new_D9151_;
  assign new_D9197_ = new_D9137_ & ~new_D9151_;
  assign new_D9198_ = ~new_D9137_ & new_D9151_;
  assign new_D9199_ = new_G4735_;
  assign new_D9200_ = new_G4802_;
  assign new_D9201_ = new_G4869_;
  assign new_D9202_ = new_G4936_;
  assign new_D9203_ = new_G5003_;
  assign new_D9204_ = new_G5070_;
  assign new_D9205_ = new_D9212_ & new_D9211_;
  assign new_D9206_ = new_D9214_ | new_D9213_;
  assign new_D9207_ = new_D9216_ | new_D9215_;
  assign new_D9208_ = new_D9218_ & new_D9217_;
  assign new_D9209_ = new_D9218_ & new_D9219_;
  assign new_D9210_ = new_D9211_ | new_D9220_;
  assign new_D9211_ = new_D9200_ | new_D9223_;
  assign new_D9212_ = new_D9222_ | new_D9221_;
  assign new_D9213_ = new_D9227_ & new_D9226_;
  assign new_D9214_ = new_D9225_ & new_D9224_;
  assign new_D9215_ = new_D9230_ | new_D9229_;
  assign new_D9216_ = new_D9225_ & new_D9228_;
  assign new_D9217_ = new_D9200_ | new_D9233_;
  assign new_D9218_ = new_D9232_ | new_D9231_;
  assign new_D9219_ = new_D9235_ | new_D9234_;
  assign new_D9220_ = ~new_D9211_ & new_D9237_;
  assign new_D9221_ = ~new_D9213_ & new_D9225_;
  assign new_D9222_ = new_D9213_ & ~new_D9225_;
  assign new_D9223_ = new_D9199_ & ~new_D9200_;
  assign new_D9224_ = ~new_D9246_ | ~new_D9247_;
  assign new_D9225_ = new_D9239_ | new_D9241_;
  assign new_D9226_ = new_D9249_ | new_D9248_;
  assign new_D9227_ = new_D9243_ | new_D9242_;
  assign new_D9228_ = ~new_D9251_ | ~new_D9250_;
  assign new_D9229_ = ~new_D9252_ & new_D9253_;
  assign new_D9230_ = new_D9252_ & ~new_D9253_;
  assign new_D9231_ = ~new_D9199_ & new_D9200_;
  assign new_D9232_ = new_D9199_ & ~new_D9200_;
  assign new_D9233_ = ~new_D9215_ | new_D9225_;
  assign new_D9234_ = new_D9215_ & new_D9225_;
  assign new_D9235_ = ~new_D9215_ & ~new_D9225_;
  assign new_D9236_ = new_D9257_ | new_D9256_;
  assign new_D9237_ = new_D9203_ | new_D9236_;
  assign new_D9238_ = new_D9261_ | new_D9260_;
  assign new_D9239_ = ~new_D9203_ & new_D9238_;
  assign new_D9240_ = new_D9259_ | new_D9258_;
  assign new_D9241_ = new_D9203_ & new_D9240_;
  assign new_D9242_ = new_D9201_ & ~new_D9211_;
  assign new_D9243_ = ~new_D9201_ & new_D9211_;
  assign new_D9244_ = ~new_D9200_ | ~new_D9225_;
  assign new_D9245_ = new_D9211_ & new_D9244_;
  assign new_D9246_ = ~new_D9211_ & ~new_D9245_;
  assign new_D9247_ = new_D9211_ | new_D9244_;
  assign new_D9248_ = ~new_D9201_ & new_D9202_;
  assign new_D9249_ = new_D9201_ & ~new_D9202_;
  assign new_D9250_ = new_D9218_ | new_D9255_;
  assign new_D9251_ = ~new_D9218_ & ~new_D9254_;
  assign new_D9252_ = new_D9201_ | new_D9218_;
  assign new_D9253_ = new_D9201_ | new_D9202_;
  assign new_D9254_ = new_D9218_ & new_D9255_;
  assign new_D9255_ = ~new_D9200_ | ~new_D9225_;
  assign new_D9256_ = new_D9233_ & new_D9253_;
  assign new_D9257_ = ~new_D9233_ & ~new_D9253_;
  assign new_D9258_ = new_D9262_ | new_D9263_;
  assign new_D9259_ = ~new_D9204_ & new_D9218_;
  assign new_D9260_ = new_D9264_ | new_D9265_;
  assign new_D9261_ = new_D9204_ & new_D9218_;
  assign new_D9262_ = ~new_D9204_ & ~new_D9218_;
  assign new_D9263_ = new_D9204_ & ~new_D9218_;
  assign new_D9264_ = new_D9204_ & ~new_D9218_;
  assign new_D9265_ = ~new_D9204_ & new_D9218_;
  assign new_D9266_ = new_G5137_;
  assign new_D9267_ = new_G5204_;
  assign new_D9268_ = new_G5271_;
  assign new_D9269_ = new_G5338_;
  assign new_D9270_ = new_G5405_;
  assign new_D9271_ = new_G5472_;
  assign new_D9272_ = new_D9279_ & new_D9278_;
  assign new_D9273_ = new_D9281_ | new_D9280_;
  assign new_D9274_ = new_D9283_ | new_D9282_;
  assign new_D9275_ = new_D9285_ & new_D9284_;
  assign new_D9276_ = new_D9285_ & new_D9286_;
  assign new_D9277_ = new_D9278_ | new_D9287_;
  assign new_D9278_ = new_D9267_ | new_D9290_;
  assign new_D9279_ = new_D9289_ | new_D9288_;
  assign new_D9280_ = new_D9294_ & new_D9293_;
  assign new_D9281_ = new_D9292_ & new_D9291_;
  assign new_D9282_ = new_D9297_ | new_D9296_;
  assign new_D9283_ = new_D9292_ & new_D9295_;
  assign new_D9284_ = new_D9267_ | new_D9300_;
  assign new_D9285_ = new_D9299_ | new_D9298_;
  assign new_D9286_ = new_D9302_ | new_D9301_;
  assign new_D9287_ = ~new_D9278_ & new_D9304_;
  assign new_D9288_ = ~new_D9280_ & new_D9292_;
  assign new_D9289_ = new_D9280_ & ~new_D9292_;
  assign new_D9290_ = new_D9266_ & ~new_D9267_;
  assign new_D9291_ = ~new_D9313_ | ~new_D9314_;
  assign new_D9292_ = new_D9306_ | new_D9308_;
  assign new_D9293_ = new_D9316_ | new_D9315_;
  assign new_D9294_ = new_D9310_ | new_D9309_;
  assign new_D9295_ = ~new_D9318_ | ~new_D9317_;
  assign new_D9296_ = ~new_D9319_ & new_D9320_;
  assign new_D9297_ = new_D9319_ & ~new_D9320_;
  assign new_D9298_ = ~new_D9266_ & new_D9267_;
  assign new_D9299_ = new_D9266_ & ~new_D9267_;
  assign new_D9300_ = ~new_D9282_ | new_D9292_;
  assign new_D9301_ = new_D9282_ & new_D9292_;
  assign new_D9302_ = ~new_D9282_ & ~new_D9292_;
  assign new_D9303_ = new_D9324_ | new_D9323_;
  assign new_D9304_ = new_D9270_ | new_D9303_;
  assign new_D9305_ = new_D9328_ | new_D9327_;
  assign new_D9306_ = ~new_D9270_ & new_D9305_;
  assign new_D9307_ = new_D9326_ | new_D9325_;
  assign new_D9308_ = new_D9270_ & new_D9307_;
  assign new_D9309_ = new_D9268_ & ~new_D9278_;
  assign new_D9310_ = ~new_D9268_ & new_D9278_;
  assign new_D9311_ = ~new_D9267_ | ~new_D9292_;
  assign new_D9312_ = new_D9278_ & new_D9311_;
  assign new_D9313_ = ~new_D9278_ & ~new_D9312_;
  assign new_D9314_ = new_D9278_ | new_D9311_;
  assign new_D9315_ = ~new_D9268_ & new_D9269_;
  assign new_D9316_ = new_D9268_ & ~new_D9269_;
  assign new_D9317_ = new_D9285_ | new_D9322_;
  assign new_D9318_ = ~new_D9285_ & ~new_D9321_;
  assign new_D9319_ = new_D9268_ | new_D9285_;
  assign new_D9320_ = new_D9268_ | new_D9269_;
  assign new_D9321_ = new_D9285_ & new_D9322_;
  assign new_D9322_ = ~new_D9267_ | ~new_D9292_;
  assign new_D9323_ = new_D9300_ & new_D9320_;
  assign new_D9324_ = ~new_D9300_ & ~new_D9320_;
  assign new_D9325_ = new_D9329_ | new_D9330_;
  assign new_D9326_ = ~new_D9271_ & new_D9285_;
  assign new_D9327_ = new_D9331_ | new_D9332_;
  assign new_D9328_ = new_D9271_ & new_D9285_;
  assign new_D9329_ = ~new_D9271_ & ~new_D9285_;
  assign new_D9330_ = new_D9271_ & ~new_D9285_;
  assign new_D9331_ = new_D9271_ & ~new_D9285_;
  assign new_D9332_ = ~new_D9271_ & new_D9285_;
  assign new_D9333_ = new_G5539_;
  assign new_D9334_ = new_G5606_;
  assign new_D9335_ = new_G5673_;
  assign new_D9336_ = new_G5740_;
  assign new_D9337_ = new_G5807_;
  assign new_D9338_ = new_G5874_;
  assign new_D9339_ = new_D9346_ & new_D9345_;
  assign new_D9340_ = new_D9348_ | new_D9347_;
  assign new_D9341_ = new_D9350_ | new_D9349_;
  assign new_D9342_ = new_D9352_ & new_D9351_;
  assign new_D9343_ = new_D9352_ & new_D9353_;
  assign new_D9344_ = new_D9345_ | new_D9354_;
  assign new_D9345_ = new_D9334_ | new_D9357_;
  assign new_D9346_ = new_D9356_ | new_D9355_;
  assign new_D9347_ = new_D9361_ & new_D9360_;
  assign new_D9348_ = new_D9359_ & new_D9358_;
  assign new_D9349_ = new_D9364_ | new_D9363_;
  assign new_D9350_ = new_D9359_ & new_D9362_;
  assign new_D9351_ = new_D9334_ | new_D9367_;
  assign new_D9352_ = new_D9366_ | new_D9365_;
  assign new_D9353_ = new_D9369_ | new_D9368_;
  assign new_D9354_ = ~new_D9345_ & new_D9371_;
  assign new_D9355_ = ~new_D9347_ & new_D9359_;
  assign new_D9356_ = new_D9347_ & ~new_D9359_;
  assign new_D9357_ = new_D9333_ & ~new_D9334_;
  assign new_D9358_ = ~new_D9380_ | ~new_D9381_;
  assign new_D9359_ = new_D9373_ | new_D9375_;
  assign new_D9360_ = new_D9383_ | new_D9382_;
  assign new_D9361_ = new_D9377_ | new_D9376_;
  assign new_D9362_ = ~new_D9385_ | ~new_D9384_;
  assign new_D9363_ = ~new_D9386_ & new_D9387_;
  assign new_D9364_ = new_D9386_ & ~new_D9387_;
  assign new_D9365_ = ~new_D9333_ & new_D9334_;
  assign new_D9366_ = new_D9333_ & ~new_D9334_;
  assign new_D9367_ = ~new_D9349_ | new_D9359_;
  assign new_D9368_ = new_D9349_ & new_D9359_;
  assign new_D9369_ = ~new_D9349_ & ~new_D9359_;
  assign new_D9370_ = new_D9391_ | new_D9390_;
  assign new_D9371_ = new_D9337_ | new_D9370_;
  assign new_D9372_ = new_D9395_ | new_D9394_;
  assign new_D9373_ = ~new_D9337_ & new_D9372_;
  assign new_D9374_ = new_D9393_ | new_D9392_;
  assign new_D9375_ = new_D9337_ & new_D9374_;
  assign new_D9376_ = new_D9335_ & ~new_D9345_;
  assign new_D9377_ = ~new_D9335_ & new_D9345_;
  assign new_D9378_ = ~new_D9334_ | ~new_D9359_;
  assign new_D9379_ = new_D9345_ & new_D9378_;
  assign new_D9380_ = ~new_D9345_ & ~new_D9379_;
  assign new_D9381_ = new_D9345_ | new_D9378_;
  assign new_D9382_ = ~new_D9335_ & new_D9336_;
  assign new_D9383_ = new_D9335_ & ~new_D9336_;
  assign new_D9384_ = new_D9352_ | new_D9389_;
  assign new_D9385_ = ~new_D9352_ & ~new_D9388_;
  assign new_D9386_ = new_D9335_ | new_D9352_;
  assign new_D9387_ = new_D9335_ | new_D9336_;
  assign new_D9388_ = new_D9352_ & new_D9389_;
  assign new_D9389_ = ~new_D9334_ | ~new_D9359_;
  assign new_D9390_ = new_D9367_ & new_D9387_;
  assign new_D9391_ = ~new_D9367_ & ~new_D9387_;
  assign new_D9392_ = new_D9396_ | new_D9397_;
  assign new_D9393_ = ~new_D9338_ & new_D9352_;
  assign new_D9394_ = new_D9398_ | new_D9399_;
  assign new_D9395_ = new_D9338_ & new_D9352_;
  assign new_D9396_ = ~new_D9338_ & ~new_D9352_;
  assign new_D9397_ = new_D9338_ & ~new_D9352_;
  assign new_D9398_ = new_D9338_ & ~new_D9352_;
  assign new_D9399_ = ~new_D9338_ & new_D9352_;
  assign new_D9400_ = new_F1472_;
  assign new_D9401_ = new_F1536_;
  assign new_D9402_ = new_F1603_;
  assign new_D9403_ = new_F1670_;
  assign new_D9404_ = new_F1737_;
  assign new_D9405_ = new_F1804_;
  assign new_D9406_ = new_D9413_ & new_D9412_;
  assign new_D9407_ = new_D9415_ | new_D9414_;
  assign new_D9408_ = new_D9417_ | new_D9416_;
  assign new_D9409_ = new_D9419_ & new_D9418_;
  assign new_D9410_ = new_D9419_ & new_D9420_;
  assign new_D9411_ = new_D9412_ | new_D9421_;
  assign new_D9412_ = new_D9401_ | new_D9424_;
  assign new_D9413_ = new_D9423_ | new_D9422_;
  assign new_D9414_ = new_D9428_ & new_D9427_;
  assign new_D9415_ = new_D9426_ & new_D9425_;
  assign new_D9416_ = new_D9431_ | new_D9430_;
  assign new_D9417_ = new_D9426_ & new_D9429_;
  assign new_D9418_ = new_D9401_ | new_D9434_;
  assign new_D9419_ = new_D9433_ | new_D9432_;
  assign new_D9420_ = new_D9436_ | new_D9435_;
  assign new_D9421_ = ~new_D9412_ & new_D9438_;
  assign new_D9422_ = ~new_D9414_ & new_D9426_;
  assign new_D9423_ = new_D9414_ & ~new_D9426_;
  assign new_D9424_ = new_D9400_ & ~new_D9401_;
  assign new_D9425_ = ~new_D9447_ | ~new_D9448_;
  assign new_D9426_ = new_D9440_ | new_D9442_;
  assign new_D9427_ = new_D9450_ | new_D9449_;
  assign new_D9428_ = new_D9444_ | new_D9443_;
  assign new_D9429_ = ~new_D9452_ | ~new_D9451_;
  assign new_D9430_ = ~new_D9453_ & new_D9454_;
  assign new_D9431_ = new_D9453_ & ~new_D9454_;
  assign new_D9432_ = ~new_D9400_ & new_D9401_;
  assign new_D9433_ = new_D9400_ & ~new_D9401_;
  assign new_D9434_ = ~new_D9416_ | new_D9426_;
  assign new_D9435_ = new_D9416_ & new_D9426_;
  assign new_D9436_ = ~new_D9416_ & ~new_D9426_;
  assign new_D9437_ = new_D9458_ | new_D9457_;
  assign new_D9438_ = new_D9404_ | new_D9437_;
  assign new_D9439_ = new_D9462_ | new_D9461_;
  assign new_D9440_ = ~new_D9404_ & new_D9439_;
  assign new_D9441_ = new_D9460_ | new_D9459_;
  assign new_D9442_ = new_D9404_ & new_D9441_;
  assign new_D9443_ = new_D9402_ & ~new_D9412_;
  assign new_D9444_ = ~new_D9402_ & new_D9412_;
  assign new_D9445_ = ~new_D9401_ | ~new_D9426_;
  assign new_D9446_ = new_D9412_ & new_D9445_;
  assign new_D9447_ = ~new_D9412_ & ~new_D9446_;
  assign new_D9448_ = new_D9412_ | new_D9445_;
  assign new_D9449_ = ~new_D9402_ & new_D9403_;
  assign new_D9450_ = new_D9402_ & ~new_D9403_;
  assign new_D9451_ = new_D9419_ | new_D9456_;
  assign new_D9452_ = ~new_D9419_ & ~new_D9455_;
  assign new_D9453_ = new_D9402_ | new_D9419_;
  assign new_D9454_ = new_D9402_ | new_D9403_;
  assign new_D9455_ = new_D9419_ & new_D9456_;
  assign new_D9456_ = ~new_D9401_ | ~new_D9426_;
  assign new_D9457_ = new_D9434_ & new_D9454_;
  assign new_D9458_ = ~new_D9434_ & ~new_D9454_;
  assign new_D9459_ = new_D9463_ | new_D9464_;
  assign new_D9460_ = ~new_D9405_ & new_D9419_;
  assign new_D9461_ = new_D9465_ | new_D9466_;
  assign new_D9462_ = new_D9405_ & new_D9419_;
  assign new_D9463_ = ~new_D9405_ & ~new_D9419_;
  assign new_D9464_ = new_D9405_ & ~new_D9419_;
  assign new_D9465_ = new_D9405_ & ~new_D9419_;
  assign new_D9466_ = ~new_D9405_ & new_D9419_;
  assign new_D9467_ = new_F1871_;
  assign new_D9468_ = new_F1938_;
  assign new_D9469_ = new_F2005_;
  assign new_D9470_ = new_F2072_;
  assign new_D9471_ = new_F2139_;
  assign new_D9472_ = new_F2206_;
  assign new_D9473_ = new_D9480_ & new_D9479_;
  assign new_D9474_ = new_D9482_ | new_D9481_;
  assign new_D9475_ = new_D9484_ | new_D9483_;
  assign new_D9476_ = new_D9486_ & new_D9485_;
  assign new_D9477_ = new_D9486_ & new_D9487_;
  assign new_D9478_ = new_D9479_ | new_D9488_;
  assign new_D9479_ = new_D9468_ | new_D9491_;
  assign new_D9480_ = new_D9490_ | new_D9489_;
  assign new_D9481_ = new_D9495_ & new_D9494_;
  assign new_D9482_ = new_D9493_ & new_D9492_;
  assign new_D9483_ = new_D9498_ | new_D9497_;
  assign new_D9484_ = new_D9493_ & new_D9496_;
  assign new_D9485_ = new_D9468_ | new_D9501_;
  assign new_D9486_ = new_D9500_ | new_D9499_;
  assign new_D9487_ = new_D9503_ | new_D9502_;
  assign new_D9488_ = ~new_D9479_ & new_D9505_;
  assign new_D9489_ = ~new_D9481_ & new_D9493_;
  assign new_D9490_ = new_D9481_ & ~new_D9493_;
  assign new_D9491_ = new_D9467_ & ~new_D9468_;
  assign new_D9492_ = ~new_D9514_ | ~new_D9515_;
  assign new_D9493_ = new_D9507_ | new_D9509_;
  assign new_D9494_ = new_D9517_ | new_D9516_;
  assign new_D9495_ = new_D9511_ | new_D9510_;
  assign new_D9496_ = ~new_D9519_ | ~new_D9518_;
  assign new_D9497_ = ~new_D9520_ & new_D9521_;
  assign new_D9498_ = new_D9520_ & ~new_D9521_;
  assign new_D9499_ = ~new_D9467_ & new_D9468_;
  assign new_D9500_ = new_D9467_ & ~new_D9468_;
  assign new_D9501_ = ~new_D9483_ | new_D9493_;
  assign new_D9502_ = new_D9483_ & new_D9493_;
  assign new_D9503_ = ~new_D9483_ & ~new_D9493_;
  assign new_D9504_ = new_D9525_ | new_D9524_;
  assign new_D9505_ = new_D9471_ | new_D9504_;
  assign new_D9506_ = new_D9529_ | new_D9528_;
  assign new_D9507_ = ~new_D9471_ & new_D9506_;
  assign new_D9508_ = new_D9527_ | new_D9526_;
  assign new_D9509_ = new_D9471_ & new_D9508_;
  assign new_D9510_ = new_D9469_ & ~new_D9479_;
  assign new_D9511_ = ~new_D9469_ & new_D9479_;
  assign new_D9512_ = ~new_D9468_ | ~new_D9493_;
  assign new_D9513_ = new_D9479_ & new_D9512_;
  assign new_D9514_ = ~new_D9479_ & ~new_D9513_;
  assign new_D9515_ = new_D9479_ | new_D9512_;
  assign new_D9516_ = ~new_D9469_ & new_D9470_;
  assign new_D9517_ = new_D9469_ & ~new_D9470_;
  assign new_D9518_ = new_D9486_ | new_D9523_;
  assign new_D9519_ = ~new_D9486_ & ~new_D9522_;
  assign new_D9520_ = new_D9469_ | new_D9486_;
  assign new_D9521_ = new_D9469_ | new_D9470_;
  assign new_D9522_ = new_D9486_ & new_D9523_;
  assign new_D9523_ = ~new_D9468_ | ~new_D9493_;
  assign new_D9524_ = new_D9501_ & new_D9521_;
  assign new_D9525_ = ~new_D9501_ & ~new_D9521_;
  assign new_D9526_ = new_D9530_ | new_D9531_;
  assign new_D9527_ = ~new_D9472_ & new_D9486_;
  assign new_D9528_ = new_D9532_ | new_D9533_;
  assign new_D9529_ = new_D9472_ & new_D9486_;
  assign new_D9530_ = ~new_D9472_ & ~new_D9486_;
  assign new_D9531_ = new_D9472_ & ~new_D9486_;
  assign new_D9532_ = new_D9472_ & ~new_D9486_;
  assign new_D9533_ = ~new_D9472_ & new_D9486_;
  assign new_D9534_ = new_F2273_;
  assign new_D9535_ = new_F2340_;
  assign new_D9536_ = new_F2407_;
  assign new_D9537_ = new_F2474_;
  assign new_D9538_ = new_F2541_;
  assign new_D9539_ = new_F2608_;
  assign new_D9540_ = new_D9547_ & new_D9546_;
  assign new_D9541_ = new_D9549_ | new_D9548_;
  assign new_D9542_ = new_D9551_ | new_D9550_;
  assign new_D9543_ = new_D9553_ & new_D9552_;
  assign new_D9544_ = new_D9553_ & new_D9554_;
  assign new_D9545_ = new_D9546_ | new_D9555_;
  assign new_D9546_ = new_D9535_ | new_D9558_;
  assign new_D9547_ = new_D9557_ | new_D9556_;
  assign new_D9548_ = new_D9562_ & new_D9561_;
  assign new_D9549_ = new_D9560_ & new_D9559_;
  assign new_D9550_ = new_D9565_ | new_D9564_;
  assign new_D9551_ = new_D9560_ & new_D9563_;
  assign new_D9552_ = new_D9535_ | new_D9568_;
  assign new_D9553_ = new_D9567_ | new_D9566_;
  assign new_D9554_ = new_D9570_ | new_D9569_;
  assign new_D9555_ = ~new_D9546_ & new_D9572_;
  assign new_D9556_ = ~new_D9548_ & new_D9560_;
  assign new_D9557_ = new_D9548_ & ~new_D9560_;
  assign new_D9558_ = new_D9534_ & ~new_D9535_;
  assign new_D9559_ = ~new_D9581_ | ~new_D9582_;
  assign new_D9560_ = new_D9574_ | new_D9576_;
  assign new_D9561_ = new_D9584_ | new_D9583_;
  assign new_D9562_ = new_D9578_ | new_D9577_;
  assign new_D9563_ = ~new_D9586_ | ~new_D9585_;
  assign new_D9564_ = ~new_D9587_ & new_D9588_;
  assign new_D9565_ = new_D9587_ & ~new_D9588_;
  assign new_D9566_ = ~new_D9534_ & new_D9535_;
  assign new_D9567_ = new_D9534_ & ~new_D9535_;
  assign new_D9568_ = ~new_D9550_ | new_D9560_;
  assign new_D9569_ = new_D9550_ & new_D9560_;
  assign new_D9570_ = ~new_D9550_ & ~new_D9560_;
  assign new_D9571_ = new_D9592_ | new_D9591_;
  assign new_D9572_ = new_D9538_ | new_D9571_;
  assign new_D9573_ = new_D9596_ | new_D9595_;
  assign new_D9574_ = ~new_D9538_ & new_D9573_;
  assign new_D9575_ = new_D9594_ | new_D9593_;
  assign new_D9576_ = new_D9538_ & new_D9575_;
  assign new_D9577_ = new_D9536_ & ~new_D9546_;
  assign new_D9578_ = ~new_D9536_ & new_D9546_;
  assign new_D9579_ = ~new_D9535_ | ~new_D9560_;
  assign new_D9580_ = new_D9546_ & new_D9579_;
  assign new_D9581_ = ~new_D9546_ & ~new_D9580_;
  assign new_D9582_ = new_D9546_ | new_D9579_;
  assign new_D9583_ = ~new_D9536_ & new_D9537_;
  assign new_D9584_ = new_D9536_ & ~new_D9537_;
  assign new_D9585_ = new_D9553_ | new_D9590_;
  assign new_D9586_ = ~new_D9553_ & ~new_D9589_;
  assign new_D9587_ = new_D9536_ | new_D9553_;
  assign new_D9588_ = new_D9536_ | new_D9537_;
  assign new_D9589_ = new_D9553_ & new_D9590_;
  assign new_D9590_ = ~new_D9535_ | ~new_D9560_;
  assign new_D9591_ = new_D9568_ & new_D9588_;
  assign new_D9592_ = ~new_D9568_ & ~new_D9588_;
  assign new_D9593_ = new_D9597_ | new_D9598_;
  assign new_D9594_ = ~new_D9539_ & new_D9553_;
  assign new_D9595_ = new_D9599_ | new_D9600_;
  assign new_D9596_ = new_D9539_ & new_D9553_;
  assign new_D9597_ = ~new_D9539_ & ~new_D9553_;
  assign new_D9598_ = new_D9539_ & ~new_D9553_;
  assign new_D9599_ = new_D9539_ & ~new_D9553_;
  assign new_D9600_ = ~new_D9539_ & new_D9553_;
  assign new_D9601_ = new_F2675_;
  assign new_D9602_ = new_F2742_;
  assign new_D9603_ = new_F2809_;
  assign new_D9604_ = new_F2876_;
  assign new_D9605_ = new_F2943_;
  assign new_D9606_ = new_F3010_;
  assign new_D9607_ = new_D9614_ & new_D9613_;
  assign new_D9608_ = new_D9616_ | new_D9615_;
  assign new_D9609_ = new_D9618_ | new_D9617_;
  assign new_D9610_ = new_D9620_ & new_D9619_;
  assign new_D9611_ = new_D9620_ & new_D9621_;
  assign new_D9612_ = new_D9613_ | new_D9622_;
  assign new_D9613_ = new_D9602_ | new_D9625_;
  assign new_D9614_ = new_D9624_ | new_D9623_;
  assign new_D9615_ = new_D9629_ & new_D9628_;
  assign new_D9616_ = new_D9627_ & new_D9626_;
  assign new_D9617_ = new_D9632_ | new_D9631_;
  assign new_D9618_ = new_D9627_ & new_D9630_;
  assign new_D9619_ = new_D9602_ | new_D9635_;
  assign new_D9620_ = new_D9634_ | new_D9633_;
  assign new_D9621_ = new_D9637_ | new_D9636_;
  assign new_D9622_ = ~new_D9613_ & new_D9639_;
  assign new_D9623_ = ~new_D9615_ & new_D9627_;
  assign new_D9624_ = new_D9615_ & ~new_D9627_;
  assign new_D9625_ = new_D9601_ & ~new_D9602_;
  assign new_D9626_ = ~new_D9648_ | ~new_D9649_;
  assign new_D9627_ = new_D9641_ | new_D9643_;
  assign new_D9628_ = new_D9651_ | new_D9650_;
  assign new_D9629_ = new_D9645_ | new_D9644_;
  assign new_D9630_ = ~new_D9653_ | ~new_D9652_;
  assign new_D9631_ = ~new_D9654_ & new_D9655_;
  assign new_D9632_ = new_D9654_ & ~new_D9655_;
  assign new_D9633_ = ~new_D9601_ & new_D9602_;
  assign new_D9634_ = new_D9601_ & ~new_D9602_;
  assign new_D9635_ = ~new_D9617_ | new_D9627_;
  assign new_D9636_ = new_D9617_ & new_D9627_;
  assign new_D9637_ = ~new_D9617_ & ~new_D9627_;
  assign new_D9638_ = new_D9659_ | new_D9658_;
  assign new_D9639_ = new_D9605_ | new_D9638_;
  assign new_D9640_ = new_D9663_ | new_D9662_;
  assign new_D9641_ = ~new_D9605_ & new_D9640_;
  assign new_D9642_ = new_D9661_ | new_D9660_;
  assign new_D9643_ = new_D9605_ & new_D9642_;
  assign new_D9644_ = new_D9603_ & ~new_D9613_;
  assign new_D9645_ = ~new_D9603_ & new_D9613_;
  assign new_D9646_ = ~new_D9602_ | ~new_D9627_;
  assign new_D9647_ = new_D9613_ & new_D9646_;
  assign new_D9648_ = ~new_D9613_ & ~new_D9647_;
  assign new_D9649_ = new_D9613_ | new_D9646_;
  assign new_D9650_ = ~new_D9603_ & new_D9604_;
  assign new_D9651_ = new_D9603_ & ~new_D9604_;
  assign new_D9652_ = new_D9620_ | new_D9657_;
  assign new_D9653_ = ~new_D9620_ & ~new_D9656_;
  assign new_D9654_ = new_D9603_ | new_D9620_;
  assign new_D9655_ = new_D9603_ | new_D9604_;
  assign new_D9656_ = new_D9620_ & new_D9657_;
  assign new_D9657_ = ~new_D9602_ | ~new_D9627_;
  assign new_D9658_ = new_D9635_ & new_D9655_;
  assign new_D9659_ = ~new_D9635_ & ~new_D9655_;
  assign new_D9660_ = new_D9664_ | new_D9665_;
  assign new_D9661_ = ~new_D9606_ & new_D9620_;
  assign new_D9662_ = new_D9666_ | new_D9667_;
  assign new_D9663_ = new_D9606_ & new_D9620_;
  assign new_D9664_ = ~new_D9606_ & ~new_D9620_;
  assign new_D9665_ = new_D9606_ & ~new_D9620_;
  assign new_D9666_ = new_D9606_ & ~new_D9620_;
  assign new_D9667_ = ~new_D9606_ & new_D9620_;
  assign new_D9668_ = new_F3077_;
  assign new_D9669_ = new_F3144_;
  assign new_D9670_ = new_F3211_;
  assign new_D9671_ = new_F3278_;
  assign new_D9672_ = new_F3345_;
  assign new_D9673_ = new_F3412_;
  assign new_D9674_ = new_D9681_ & new_D9680_;
  assign new_D9675_ = new_D9683_ | new_D9682_;
  assign new_D9676_ = new_D9685_ | new_D9684_;
  assign new_D9677_ = new_D9687_ & new_D9686_;
  assign new_D9678_ = new_D9687_ & new_D9688_;
  assign new_D9679_ = new_D9680_ | new_D9689_;
  assign new_D9680_ = new_D9669_ | new_D9692_;
  assign new_D9681_ = new_D9691_ | new_D9690_;
  assign new_D9682_ = new_D9696_ & new_D9695_;
  assign new_D9683_ = new_D9694_ & new_D9693_;
  assign new_D9684_ = new_D9699_ | new_D9698_;
  assign new_D9685_ = new_D9694_ & new_D9697_;
  assign new_D9686_ = new_D9669_ | new_D9702_;
  assign new_D9687_ = new_D9701_ | new_D9700_;
  assign new_D9688_ = new_D9704_ | new_D9703_;
  assign new_D9689_ = ~new_D9680_ & new_D9706_;
  assign new_D9690_ = ~new_D9682_ & new_D9694_;
  assign new_D9691_ = new_D9682_ & ~new_D9694_;
  assign new_D9692_ = new_D9668_ & ~new_D9669_;
  assign new_D9693_ = ~new_D9715_ | ~new_D9716_;
  assign new_D9694_ = new_D9708_ | new_D9710_;
  assign new_D9695_ = new_D9718_ | new_D9717_;
  assign new_D9696_ = new_D9712_ | new_D9711_;
  assign new_D9697_ = ~new_D9720_ | ~new_D9719_;
  assign new_D9698_ = ~new_D9721_ & new_D9722_;
  assign new_D9699_ = new_D9721_ & ~new_D9722_;
  assign new_D9700_ = ~new_D9668_ & new_D9669_;
  assign new_D9701_ = new_D9668_ & ~new_D9669_;
  assign new_D9702_ = ~new_D9684_ | new_D9694_;
  assign new_D9703_ = new_D9684_ & new_D9694_;
  assign new_D9704_ = ~new_D9684_ & ~new_D9694_;
  assign new_D9705_ = new_D9726_ | new_D9725_;
  assign new_D9706_ = new_D9672_ | new_D9705_;
  assign new_D9707_ = new_D9730_ | new_D9729_;
  assign new_D9708_ = ~new_D9672_ & new_D9707_;
  assign new_D9709_ = new_D9728_ | new_D9727_;
  assign new_D9710_ = new_D9672_ & new_D9709_;
  assign new_D9711_ = new_D9670_ & ~new_D9680_;
  assign new_D9712_ = ~new_D9670_ & new_D9680_;
  assign new_D9713_ = ~new_D9669_ | ~new_D9694_;
  assign new_D9714_ = new_D9680_ & new_D9713_;
  assign new_D9715_ = ~new_D9680_ & ~new_D9714_;
  assign new_D9716_ = new_D9680_ | new_D9713_;
  assign new_D9717_ = ~new_D9670_ & new_D9671_;
  assign new_D9718_ = new_D9670_ & ~new_D9671_;
  assign new_D9719_ = new_D9687_ | new_D9724_;
  assign new_D9720_ = ~new_D9687_ & ~new_D9723_;
  assign new_D9721_ = new_D9670_ | new_D9687_;
  assign new_D9722_ = new_D9670_ | new_D9671_;
  assign new_D9723_ = new_D9687_ & new_D9724_;
  assign new_D9724_ = ~new_D9669_ | ~new_D9694_;
  assign new_D9725_ = new_D9702_ & new_D9722_;
  assign new_D9726_ = ~new_D9702_ & ~new_D9722_;
  assign new_D9727_ = new_D9731_ | new_D9732_;
  assign new_D9728_ = ~new_D9673_ & new_D9687_;
  assign new_D9729_ = new_D9733_ | new_D9734_;
  assign new_D9730_ = new_D9673_ & new_D9687_;
  assign new_D9731_ = ~new_D9673_ & ~new_D9687_;
  assign new_D9732_ = new_D9673_ & ~new_D9687_;
  assign new_D9733_ = new_D9673_ & ~new_D9687_;
  assign new_D9734_ = ~new_D9673_ & new_D9687_;
  assign new_D9735_ = new_F3479_;
  assign new_D9736_ = new_F3546_;
  assign new_D9737_ = new_F3613_;
  assign new_D9738_ = new_F3680_;
  assign new_D9739_ = new_F3747_;
  assign new_D9740_ = new_F3814_;
  assign new_D9741_ = new_D9748_ & new_D9747_;
  assign new_D9742_ = new_D9750_ | new_D9749_;
  assign new_D9743_ = new_D9752_ | new_D9751_;
  assign new_D9744_ = new_D9754_ & new_D9753_;
  assign new_D9745_ = new_D9754_ & new_D9755_;
  assign new_D9746_ = new_D9747_ | new_D9756_;
  assign new_D9747_ = new_D9736_ | new_D9759_;
  assign new_D9748_ = new_D9758_ | new_D9757_;
  assign new_D9749_ = new_D9763_ & new_D9762_;
  assign new_D9750_ = new_D9761_ & new_D9760_;
  assign new_D9751_ = new_D9766_ | new_D9765_;
  assign new_D9752_ = new_D9761_ & new_D9764_;
  assign new_D9753_ = new_D9736_ | new_D9769_;
  assign new_D9754_ = new_D9768_ | new_D9767_;
  assign new_D9755_ = new_D9771_ | new_D9770_;
  assign new_D9756_ = ~new_D9747_ & new_D9773_;
  assign new_D9757_ = ~new_D9749_ & new_D9761_;
  assign new_D9758_ = new_D9749_ & ~new_D9761_;
  assign new_D9759_ = new_D9735_ & ~new_D9736_;
  assign new_D9760_ = ~new_D9782_ | ~new_D9783_;
  assign new_D9761_ = new_D9775_ | new_D9777_;
  assign new_D9762_ = new_D9785_ | new_D9784_;
  assign new_D9763_ = new_D9779_ | new_D9778_;
  assign new_D9764_ = ~new_D9787_ | ~new_D9786_;
  assign new_D9765_ = ~new_D9788_ & new_D9789_;
  assign new_D9766_ = new_D9788_ & ~new_D9789_;
  assign new_D9767_ = ~new_D9735_ & new_D9736_;
  assign new_D9768_ = new_D9735_ & ~new_D9736_;
  assign new_D9769_ = ~new_D9751_ | new_D9761_;
  assign new_D9770_ = new_D9751_ & new_D9761_;
  assign new_D9771_ = ~new_D9751_ & ~new_D9761_;
  assign new_D9772_ = new_D9793_ | new_D9792_;
  assign new_D9773_ = new_D9739_ | new_D9772_;
  assign new_D9774_ = new_D9797_ | new_D9796_;
  assign new_D9775_ = ~new_D9739_ & new_D9774_;
  assign new_D9776_ = new_D9795_ | new_D9794_;
  assign new_D9777_ = new_D9739_ & new_D9776_;
  assign new_D9778_ = new_D9737_ & ~new_D9747_;
  assign new_D9779_ = ~new_D9737_ & new_D9747_;
  assign new_D9780_ = ~new_D9736_ | ~new_D9761_;
  assign new_D9781_ = new_D9747_ & new_D9780_;
  assign new_D9782_ = ~new_D9747_ & ~new_D9781_;
  assign new_D9783_ = new_D9747_ | new_D9780_;
  assign new_D9784_ = ~new_D9737_ & new_D9738_;
  assign new_D9785_ = new_D9737_ & ~new_D9738_;
  assign new_D9786_ = new_D9754_ | new_D9791_;
  assign new_D9787_ = ~new_D9754_ & ~new_D9790_;
  assign new_D9788_ = new_D9737_ | new_D9754_;
  assign new_D9789_ = new_D9737_ | new_D9738_;
  assign new_D9790_ = new_D9754_ & new_D9791_;
  assign new_D9791_ = ~new_D9736_ | ~new_D9761_;
  assign new_D9792_ = new_D9769_ & new_D9789_;
  assign new_D9793_ = ~new_D9769_ & ~new_D9789_;
  assign new_D9794_ = new_D9798_ | new_D9799_;
  assign new_D9795_ = ~new_D9740_ & new_D9754_;
  assign new_D9796_ = new_D9800_ | new_D9801_;
  assign new_D9797_ = new_D9740_ & new_D9754_;
  assign new_D9798_ = ~new_D9740_ & ~new_D9754_;
  assign new_D9799_ = new_D9740_ & ~new_D9754_;
  assign new_D9800_ = new_D9740_ & ~new_D9754_;
  assign new_D9801_ = ~new_D9740_ & new_D9754_;
  assign new_D9802_ = new_F3881_;
  assign new_D9803_ = new_F3948_;
  assign new_D9804_ = new_F4015_;
  assign new_D9805_ = new_F4082_;
  assign new_D9806_ = new_F4149_;
  assign new_D9807_ = new_F4216_;
  assign new_D9808_ = new_D9815_ & new_D9814_;
  assign new_D9809_ = new_D9817_ | new_D9816_;
  assign new_D9810_ = new_D9819_ | new_D9818_;
  assign new_D9811_ = new_D9821_ & new_D9820_;
  assign new_D9812_ = new_D9821_ & new_D9822_;
  assign new_D9813_ = new_D9814_ | new_D9823_;
  assign new_D9814_ = new_D9803_ | new_D9826_;
  assign new_D9815_ = new_D9825_ | new_D9824_;
  assign new_D9816_ = new_D9830_ & new_D9829_;
  assign new_D9817_ = new_D9828_ & new_D9827_;
  assign new_D9818_ = new_D9833_ | new_D9832_;
  assign new_D9819_ = new_D9828_ & new_D9831_;
  assign new_D9820_ = new_D9803_ | new_D9836_;
  assign new_D9821_ = new_D9835_ | new_D9834_;
  assign new_D9822_ = new_D9838_ | new_D9837_;
  assign new_D9823_ = ~new_D9814_ & new_D9840_;
  assign new_D9824_ = ~new_D9816_ & new_D9828_;
  assign new_D9825_ = new_D9816_ & ~new_D9828_;
  assign new_D9826_ = new_D9802_ & ~new_D9803_;
  assign new_D9827_ = ~new_D9849_ | ~new_D9850_;
  assign new_D9828_ = new_D9842_ | new_D9844_;
  assign new_D9829_ = new_D9852_ | new_D9851_;
  assign new_D9830_ = new_D9846_ | new_D9845_;
  assign new_D9831_ = ~new_D9854_ | ~new_D9853_;
  assign new_D9832_ = ~new_D9855_ & new_D9856_;
  assign new_D9833_ = new_D9855_ & ~new_D9856_;
  assign new_D9834_ = ~new_D9802_ & new_D9803_;
  assign new_D9835_ = new_D9802_ & ~new_D9803_;
  assign new_D9836_ = ~new_D9818_ | new_D9828_;
  assign new_D9837_ = new_D9818_ & new_D9828_;
  assign new_D9838_ = ~new_D9818_ & ~new_D9828_;
  assign new_D9839_ = new_D9860_ | new_D9859_;
  assign new_D9840_ = new_D9806_ | new_D9839_;
  assign new_D9841_ = new_D9864_ | new_D9863_;
  assign new_D9842_ = ~new_D9806_ & new_D9841_;
  assign new_D9843_ = new_D9862_ | new_D9861_;
  assign new_D9844_ = new_D9806_ & new_D9843_;
  assign new_D9845_ = new_D9804_ & ~new_D9814_;
  assign new_D9846_ = ~new_D9804_ & new_D9814_;
  assign new_D9847_ = ~new_D9803_ | ~new_D9828_;
  assign new_D9848_ = new_D9814_ & new_D9847_;
  assign new_D9849_ = ~new_D9814_ & ~new_D9848_;
  assign new_D9850_ = new_D9814_ | new_D9847_;
  assign new_D9851_ = ~new_D9804_ & new_D9805_;
  assign new_D9852_ = new_D9804_ & ~new_D9805_;
  assign new_D9853_ = new_D9821_ | new_D9858_;
  assign new_D9854_ = ~new_D9821_ & ~new_D9857_;
  assign new_D9855_ = new_D9804_ | new_D9821_;
  assign new_D9856_ = new_D9804_ | new_D9805_;
  assign new_D9857_ = new_D9821_ & new_D9858_;
  assign new_D9858_ = ~new_D9803_ | ~new_D9828_;
  assign new_D9859_ = new_D9836_ & new_D9856_;
  assign new_D9860_ = ~new_D9836_ & ~new_D9856_;
  assign new_D9861_ = new_D9865_ | new_D9866_;
  assign new_D9862_ = ~new_D9807_ & new_D9821_;
  assign new_D9863_ = new_D9867_ | new_D9868_;
  assign new_D9864_ = new_D9807_ & new_D9821_;
  assign new_D9865_ = ~new_D9807_ & ~new_D9821_;
  assign new_D9866_ = new_D9807_ & ~new_D9821_;
  assign new_D9867_ = new_D9807_ & ~new_D9821_;
  assign new_D9868_ = ~new_D9807_ & new_D9821_;
  assign new_D9869_ = new_F4283_;
  assign new_D9870_ = new_F4350_;
  assign new_D9871_ = new_F4417_;
  assign new_D9872_ = new_F4484_;
  assign new_D9873_ = new_F4551_;
  assign new_D9874_ = new_F4618_;
  assign new_D9875_ = new_D9882_ & new_D9881_;
  assign new_D9876_ = new_D9884_ | new_D9883_;
  assign new_D9877_ = new_D9886_ | new_D9885_;
  assign new_D9878_ = new_D9888_ & new_D9887_;
  assign new_D9879_ = new_D9888_ & new_D9889_;
  assign new_D9880_ = new_D9881_ | new_D9890_;
  assign new_D9881_ = new_D9870_ | new_D9893_;
  assign new_D9882_ = new_D9892_ | new_D9891_;
  assign new_D9883_ = new_D9897_ & new_D9896_;
  assign new_D9884_ = new_D9895_ & new_D9894_;
  assign new_D9885_ = new_D9900_ | new_D9899_;
  assign new_D9886_ = new_D9895_ & new_D9898_;
  assign new_D9887_ = new_D9870_ | new_D9903_;
  assign new_D9888_ = new_D9902_ | new_D9901_;
  assign new_D9889_ = new_D9905_ | new_D9904_;
  assign new_D9890_ = ~new_D9881_ & new_D9907_;
  assign new_D9891_ = ~new_D9883_ & new_D9895_;
  assign new_D9892_ = new_D9883_ & ~new_D9895_;
  assign new_D9893_ = new_D9869_ & ~new_D9870_;
  assign new_D9894_ = ~new_D9916_ | ~new_D9917_;
  assign new_D9895_ = new_D9909_ | new_D9911_;
  assign new_D9896_ = new_D9919_ | new_D9918_;
  assign new_D9897_ = new_D9913_ | new_D9912_;
  assign new_D9898_ = ~new_D9921_ | ~new_D9920_;
  assign new_D9899_ = ~new_D9922_ & new_D9923_;
  assign new_D9900_ = new_D9922_ & ~new_D9923_;
  assign new_D9901_ = ~new_D9869_ & new_D9870_;
  assign new_D9902_ = new_D9869_ & ~new_D9870_;
  assign new_D9903_ = ~new_D9885_ | new_D9895_;
  assign new_D9904_ = new_D9885_ & new_D9895_;
  assign new_D9905_ = ~new_D9885_ & ~new_D9895_;
  assign new_D9906_ = new_D9927_ | new_D9926_;
  assign new_D9907_ = new_D9873_ | new_D9906_;
  assign new_D9908_ = new_D9931_ | new_D9930_;
  assign new_D9909_ = ~new_D9873_ & new_D9908_;
  assign new_D9910_ = new_D9929_ | new_D9928_;
  assign new_D9911_ = new_D9873_ & new_D9910_;
  assign new_D9912_ = new_D9871_ & ~new_D9881_;
  assign new_D9913_ = ~new_D9871_ & new_D9881_;
  assign new_D9914_ = ~new_D9870_ | ~new_D9895_;
  assign new_D9915_ = new_D9881_ & new_D9914_;
  assign new_D9916_ = ~new_D9881_ & ~new_D9915_;
  assign new_D9917_ = new_D9881_ | new_D9914_;
  assign new_D9918_ = ~new_D9871_ & new_D9872_;
  assign new_D9919_ = new_D9871_ & ~new_D9872_;
  assign new_D9920_ = new_D9888_ | new_D9925_;
  assign new_D9921_ = ~new_D9888_ & ~new_D9924_;
  assign new_D9922_ = new_D9871_ | new_D9888_;
  assign new_D9923_ = new_D9871_ | new_D9872_;
  assign new_D9924_ = new_D9888_ & new_D9925_;
  assign new_D9925_ = ~new_D9870_ | ~new_D9895_;
  assign new_D9926_ = new_D9903_ & new_D9923_;
  assign new_D9927_ = ~new_D9903_ & ~new_D9923_;
  assign new_D9928_ = new_D9932_ | new_D9933_;
  assign new_D9929_ = ~new_D9874_ & new_D9888_;
  assign new_D9930_ = new_D9934_ | new_D9935_;
  assign new_D9931_ = new_D9874_ & new_D9888_;
  assign new_D9932_ = ~new_D9874_ & ~new_D9888_;
  assign new_D9933_ = new_D9874_ & ~new_D9888_;
  assign new_D9934_ = new_D9874_ & ~new_D9888_;
  assign new_D9935_ = ~new_D9874_ & new_D9888_;
  assign new_D9936_ = new_F4685_;
  assign new_D9937_ = new_F4752_;
  assign new_D9938_ = new_F4819_;
  assign new_D9939_ = new_F4886_;
  assign new_D9940_ = new_F4953_;
  assign new_D9941_ = new_F5020_;
  assign new_D9942_ = new_D9949_ & new_D9948_;
  assign new_D9943_ = new_D9951_ | new_D9950_;
  assign new_D9944_ = new_D9953_ | new_D9952_;
  assign new_D9945_ = new_D9955_ & new_D9954_;
  assign new_D9946_ = new_D9955_ & new_D9956_;
  assign new_D9947_ = new_D9948_ | new_D9957_;
  assign new_D9948_ = new_D9937_ | new_D9960_;
  assign new_D9949_ = new_D9959_ | new_D9958_;
  assign new_D9950_ = new_D9964_ & new_D9963_;
  assign new_D9951_ = new_D9962_ & new_D9961_;
  assign new_D9952_ = new_D9967_ | new_D9966_;
  assign new_D9953_ = new_D9962_ & new_D9965_;
  assign new_D9954_ = new_D9937_ | new_D9970_;
  assign new_D9955_ = new_D9969_ | new_D9968_;
  assign new_D9956_ = new_D9972_ | new_D9971_;
  assign new_D9957_ = ~new_D9948_ & new_D9974_;
  assign new_D9958_ = ~new_D9950_ & new_D9962_;
  assign new_D9959_ = new_D9950_ & ~new_D9962_;
  assign new_D9960_ = new_D9936_ & ~new_D9937_;
  assign new_D9961_ = ~new_D9983_ | ~new_D9984_;
  assign new_D9962_ = new_D9976_ | new_D9978_;
  assign new_D9963_ = new_D9986_ | new_D9985_;
  assign new_D9964_ = new_D9980_ | new_D9979_;
  assign new_D9965_ = ~new_D9988_ | ~new_D9987_;
  assign new_D9966_ = ~new_D9989_ & new_D9990_;
  assign new_D9967_ = new_D9989_ & ~new_D9990_;
  assign new_D9968_ = ~new_D9936_ & new_D9937_;
  assign new_D9969_ = new_D9936_ & ~new_D9937_;
  assign new_D9970_ = ~new_D9952_ | new_D9962_;
  assign new_D9971_ = new_D9952_ & new_D9962_;
  assign new_D9972_ = ~new_D9952_ & ~new_D9962_;
  assign new_D9973_ = new_D9994_ | new_D9993_;
  assign new_D9974_ = new_D9940_ | new_D9973_;
  assign new_D9975_ = new_D9998_ | new_D9997_;
  assign new_D9976_ = ~new_D9940_ & new_D9975_;
  assign new_D9977_ = new_D9996_ | new_D9995_;
  assign new_D9978_ = new_D9940_ & new_D9977_;
  assign new_D9979_ = new_D9938_ & ~new_D9948_;
  assign new_D9980_ = ~new_D9938_ & new_D9948_;
  assign new_D9981_ = ~new_D9937_ | ~new_D9962_;
  assign new_D9982_ = new_D9948_ & new_D9981_;
  assign new_D9983_ = ~new_D9948_ & ~new_D9982_;
  assign new_D9984_ = new_D9948_ | new_D9981_;
  assign new_D9985_ = ~new_D9938_ & new_D9939_;
  assign new_D9986_ = new_D9938_ & ~new_D9939_;
  assign new_D9987_ = new_D9955_ | new_D9992_;
  assign new_D9988_ = ~new_D9955_ & ~new_D9991_;
  assign new_D9989_ = new_D9938_ | new_D9955_;
  assign new_D9990_ = new_D9938_ | new_D9939_;
  assign new_D9991_ = new_D9955_ & new_D9992_;
  assign new_D9992_ = ~new_D9937_ | ~new_D9962_;
  assign new_D9993_ = new_D9970_ & new_D9990_;
  assign new_D9994_ = ~new_D9970_ & ~new_D9990_;
  assign new_D9995_ = new_D9999_ | new_E1_;
  assign new_D9996_ = ~new_D9941_ & new_D9955_;
  assign new_D9997_ = new_E2_ | new_E3_;
  assign new_D9998_ = new_D9941_ & new_D9955_;
  assign new_D9999_ = ~new_D9941_ & ~new_D9955_;
  assign new_E1_ = new_D9941_ & ~new_D9955_;
  assign new_E2_ = new_D9941_ & ~new_D9955_;
  assign new_E3_ = ~new_D9941_ & new_D9955_;
  assign new_E4_ = new_F5087_;
  assign new_E5_ = new_F5154_;
  assign new_E6_ = new_F5221_;
  assign new_E7_ = new_F5288_;
  assign new_E8_ = new_F5355_;
  assign new_E9_ = new_F5422_;
  assign new_E10_ = new_E17_ & new_E16_;
  assign new_E11_ = new_E19_ | new_E18_;
  assign new_E12_ = new_E21_ | new_E20_;
  assign new_E13_ = new_E23_ & new_E22_;
  assign new_E14_ = new_E23_ & new_E24_;
  assign new_E15_ = new_E16_ | new_E25_;
  assign new_E16_ = new_E5_ | new_E28_;
  assign new_E17_ = new_E27_ | new_E26_;
  assign new_E18_ = new_E32_ & new_E31_;
  assign new_E19_ = new_E30_ & new_E29_;
  assign new_E20_ = new_E35_ | new_E34_;
  assign new_E21_ = new_E30_ & new_E33_;
  assign new_E22_ = new_E5_ | new_E38_;
  assign new_E23_ = new_E37_ | new_E36_;
  assign new_E24_ = new_E40_ | new_E39_;
  assign new_E25_ = ~new_E16_ & new_E42_;
  assign new_E26_ = ~new_E18_ & new_E30_;
  assign new_E27_ = new_E18_ & ~new_E30_;
  assign new_E28_ = new_E4_ & ~new_E5_;
  assign new_E29_ = ~new_E51_ | ~new_E52_;
  assign new_E30_ = new_E44_ | new_E46_;
  assign new_E31_ = new_E54_ | new_E53_;
  assign new_E32_ = new_E48_ | new_E47_;
  assign new_E33_ = ~new_E56_ | ~new_E55_;
  assign new_E34_ = ~new_E57_ & new_E58_;
  assign new_E35_ = new_E57_ & ~new_E58_;
  assign new_E36_ = ~new_E4_ & new_E5_;
  assign new_E37_ = new_E4_ & ~new_E5_;
  assign new_E38_ = ~new_E20_ | new_E30_;
  assign new_E39_ = new_E20_ & new_E30_;
  assign new_E40_ = ~new_E20_ & ~new_E30_;
  assign new_E41_ = new_E62_ | new_E61_;
  assign new_E42_ = new_E8_ | new_E41_;
  assign new_E43_ = new_E66_ | new_E65_;
  assign new_E44_ = ~new_E8_ & new_E43_;
  assign new_E45_ = new_E64_ | new_E63_;
  assign new_E46_ = new_E8_ & new_E45_;
  assign new_E47_ = new_E6_ & ~new_E16_;
  assign new_E48_ = ~new_E6_ & new_E16_;
  assign new_E49_ = ~new_E5_ | ~new_E30_;
  assign new_E50_ = new_E16_ & new_E49_;
  assign new_E51_ = ~new_E16_ & ~new_E50_;
  assign new_E52_ = new_E16_ | new_E49_;
  assign new_E53_ = ~new_E6_ & new_E7_;
  assign new_E54_ = new_E6_ & ~new_E7_;
  assign new_E55_ = new_E23_ | new_E60_;
  assign new_E56_ = ~new_E23_ & ~new_E59_;
  assign new_E57_ = new_E6_ | new_E23_;
  assign new_E58_ = new_E6_ | new_E7_;
  assign new_E59_ = new_E23_ & new_E60_;
  assign new_E60_ = ~new_E5_ | ~new_E30_;
  assign new_E61_ = new_E38_ & new_E58_;
  assign new_E62_ = ~new_E38_ & ~new_E58_;
  assign new_E63_ = new_E67_ | new_E68_;
  assign new_E64_ = ~new_E9_ & new_E23_;
  assign new_E65_ = new_E69_ | new_E70_;
  assign new_E66_ = new_E9_ & new_E23_;
  assign new_E67_ = ~new_E9_ & ~new_E23_;
  assign new_E68_ = new_E9_ & ~new_E23_;
  assign new_E69_ = new_E9_ & ~new_E23_;
  assign new_E70_ = ~new_E9_ & new_E23_;
  assign new_E71_ = new_F5489_;
  assign new_E72_ = new_F5556_;
  assign new_E73_ = new_F5623_;
  assign new_E74_ = new_F5690_;
  assign new_E75_ = new_F5757_;
  assign new_E76_ = new_F5824_;
  assign new_E77_ = new_E84_ & new_E83_;
  assign new_E78_ = new_E86_ | new_E85_;
  assign new_E79_ = new_E88_ | new_E87_;
  assign new_E80_ = new_E90_ & new_E89_;
  assign new_E81_ = new_E90_ & new_E91_;
  assign new_E82_ = new_E83_ | new_E92_;
  assign new_E83_ = new_E72_ | new_E95_;
  assign new_E84_ = new_E94_ | new_E93_;
  assign new_E85_ = new_E99_ & new_E98_;
  assign new_E86_ = new_E97_ & new_E96_;
  assign new_E87_ = new_E102_ | new_E101_;
  assign new_E88_ = new_E97_ & new_E100_;
  assign new_E89_ = new_E72_ | new_E105_;
  assign new_E90_ = new_E104_ | new_E103_;
  assign new_E91_ = new_E107_ | new_E106_;
  assign new_E92_ = ~new_E83_ & new_E109_;
  assign new_E93_ = ~new_E85_ & new_E97_;
  assign new_E94_ = new_E85_ & ~new_E97_;
  assign new_E95_ = new_E71_ & ~new_E72_;
  assign new_E96_ = ~new_E118_ | ~new_E119_;
  assign new_E97_ = new_E111_ | new_E113_;
  assign new_E98_ = new_E121_ | new_E120_;
  assign new_E99_ = new_E115_ | new_E114_;
  assign new_E100_ = ~new_E123_ | ~new_E122_;
  assign new_E101_ = ~new_E124_ & new_E125_;
  assign new_E102_ = new_E124_ & ~new_E125_;
  assign new_E103_ = ~new_E71_ & new_E72_;
  assign new_E104_ = new_E71_ & ~new_E72_;
  assign new_E105_ = ~new_E87_ | new_E97_;
  assign new_E106_ = new_E87_ & new_E97_;
  assign new_E107_ = ~new_E87_ & ~new_E97_;
  assign new_E108_ = new_E129_ | new_E128_;
  assign new_E109_ = new_E75_ | new_E108_;
  assign new_E110_ = new_E133_ | new_E132_;
  assign new_E111_ = ~new_E75_ & new_E110_;
  assign new_E112_ = new_E131_ | new_E130_;
  assign new_E113_ = new_E75_ & new_E112_;
  assign new_E114_ = new_E73_ & ~new_E83_;
  assign new_E115_ = ~new_E73_ & new_E83_;
  assign new_E116_ = ~new_E72_ | ~new_E97_;
  assign new_E117_ = new_E83_ & new_E116_;
  assign new_E118_ = ~new_E83_ & ~new_E117_;
  assign new_E119_ = new_E83_ | new_E116_;
  assign new_E120_ = ~new_E73_ & new_E74_;
  assign new_E121_ = new_E73_ & ~new_E74_;
  assign new_E122_ = new_E90_ | new_E127_;
  assign new_E123_ = ~new_E90_ & ~new_E126_;
  assign new_E124_ = new_E73_ | new_E90_;
  assign new_E125_ = new_E73_ | new_E74_;
  assign new_E126_ = new_E90_ & new_E127_;
  assign new_E127_ = ~new_E72_ | ~new_E97_;
  assign new_E128_ = new_E105_ & new_E125_;
  assign new_E129_ = ~new_E105_ & ~new_E125_;
  assign new_E130_ = new_E134_ | new_E135_;
  assign new_E131_ = ~new_E76_ & new_E90_;
  assign new_E132_ = new_E136_ | new_E137_;
  assign new_E133_ = new_E76_ & new_E90_;
  assign new_E134_ = ~new_E76_ & ~new_E90_;
  assign new_E135_ = new_E76_ & ~new_E90_;
  assign new_E136_ = new_E76_ & ~new_E90_;
  assign new_E137_ = ~new_E76_ & new_E90_;
  assign new_E138_ = new_F5891_;
  assign new_E139_ = new_F5958_;
  assign new_E140_ = new_F6025_;
  assign new_E141_ = new_F6092_;
  assign new_E142_ = new_F6159_;
  assign new_E143_ = new_F6226_;
  assign new_E144_ = new_E151_ & new_E150_;
  assign new_E145_ = new_E153_ | new_E152_;
  assign new_E146_ = new_E155_ | new_E154_;
  assign new_E147_ = new_E157_ & new_E156_;
  assign new_E148_ = new_E157_ & new_E158_;
  assign new_E149_ = new_E150_ | new_E159_;
  assign new_E150_ = new_E139_ | new_E162_;
  assign new_E151_ = new_E161_ | new_E160_;
  assign new_E152_ = new_E166_ & new_E165_;
  assign new_E153_ = new_E164_ & new_E163_;
  assign new_E154_ = new_E169_ | new_E168_;
  assign new_E155_ = new_E164_ & new_E167_;
  assign new_E156_ = new_E139_ | new_E172_;
  assign new_E157_ = new_E171_ | new_E170_;
  assign new_E158_ = new_E174_ | new_E173_;
  assign new_E159_ = ~new_E150_ & new_E176_;
  assign new_E160_ = ~new_E152_ & new_E164_;
  assign new_E161_ = new_E152_ & ~new_E164_;
  assign new_E162_ = new_E138_ & ~new_E139_;
  assign new_E163_ = ~new_E185_ | ~new_E186_;
  assign new_E164_ = new_E178_ | new_E180_;
  assign new_E165_ = new_E188_ | new_E187_;
  assign new_E166_ = new_E182_ | new_E181_;
  assign new_E167_ = ~new_E190_ | ~new_E189_;
  assign new_E168_ = ~new_E191_ & new_E192_;
  assign new_E169_ = new_E191_ & ~new_E192_;
  assign new_E170_ = ~new_E138_ & new_E139_;
  assign new_E171_ = new_E138_ & ~new_E139_;
  assign new_E172_ = ~new_E154_ | new_E164_;
  assign new_E173_ = new_E154_ & new_E164_;
  assign new_E174_ = ~new_E154_ & ~new_E164_;
  assign new_E175_ = new_E196_ | new_E195_;
  assign new_E176_ = new_E142_ | new_E175_;
  assign new_E177_ = new_E200_ | new_E199_;
  assign new_E178_ = ~new_E142_ & new_E177_;
  assign new_E179_ = new_E198_ | new_E197_;
  assign new_E180_ = new_E142_ & new_E179_;
  assign new_E181_ = new_E140_ & ~new_E150_;
  assign new_E182_ = ~new_E140_ & new_E150_;
  assign new_E183_ = ~new_E139_ | ~new_E164_;
  assign new_E184_ = new_E150_ & new_E183_;
  assign new_E185_ = ~new_E150_ & ~new_E184_;
  assign new_E186_ = new_E150_ | new_E183_;
  assign new_E187_ = ~new_E140_ & new_E141_;
  assign new_E188_ = new_E140_ & ~new_E141_;
  assign new_E189_ = new_E157_ | new_E194_;
  assign new_E190_ = ~new_E157_ & ~new_E193_;
  assign new_E191_ = new_E140_ | new_E157_;
  assign new_E192_ = new_E140_ | new_E141_;
  assign new_E193_ = new_E157_ & new_E194_;
  assign new_E194_ = ~new_E139_ | ~new_E164_;
  assign new_E195_ = new_E172_ & new_E192_;
  assign new_E196_ = ~new_E172_ & ~new_E192_;
  assign new_E197_ = new_E201_ | new_E202_;
  assign new_E198_ = ~new_E143_ & new_E157_;
  assign new_E199_ = new_E203_ | new_E204_;
  assign new_E200_ = new_E143_ & new_E157_;
  assign new_E201_ = ~new_E143_ & ~new_E157_;
  assign new_E202_ = new_E143_ & ~new_E157_;
  assign new_E203_ = new_E143_ & ~new_E157_;
  assign new_E204_ = ~new_E143_ & new_E157_;
  assign new_E205_ = new_F6293_;
  assign new_E206_ = new_F6360_;
  assign new_E207_ = new_F6427_;
  assign new_E208_ = new_F6494_;
  assign new_E209_ = new_F6561_;
  assign new_E210_ = new_F6628_;
  assign new_E211_ = new_E218_ & new_E217_;
  assign new_E212_ = new_E220_ | new_E219_;
  assign new_E213_ = new_E222_ | new_E221_;
  assign new_E214_ = new_E224_ & new_E223_;
  assign new_E215_ = new_E224_ & new_E225_;
  assign new_E216_ = new_E217_ | new_E226_;
  assign new_E217_ = new_E206_ | new_E229_;
  assign new_E218_ = new_E228_ | new_E227_;
  assign new_E219_ = new_E233_ & new_E232_;
  assign new_E220_ = new_E231_ & new_E230_;
  assign new_E221_ = new_E236_ | new_E235_;
  assign new_E222_ = new_E231_ & new_E234_;
  assign new_E223_ = new_E206_ | new_E239_;
  assign new_E224_ = new_E238_ | new_E237_;
  assign new_E225_ = new_E241_ | new_E240_;
  assign new_E226_ = ~new_E217_ & new_E243_;
  assign new_E227_ = ~new_E219_ & new_E231_;
  assign new_E228_ = new_E219_ & ~new_E231_;
  assign new_E229_ = new_E205_ & ~new_E206_;
  assign new_E230_ = ~new_E252_ | ~new_E253_;
  assign new_E231_ = new_E245_ | new_E247_;
  assign new_E232_ = new_E255_ | new_E254_;
  assign new_E233_ = new_E249_ | new_E248_;
  assign new_E234_ = ~new_E257_ | ~new_E256_;
  assign new_E235_ = ~new_E258_ & new_E259_;
  assign new_E236_ = new_E258_ & ~new_E259_;
  assign new_E237_ = ~new_E205_ & new_E206_;
  assign new_E238_ = new_E205_ & ~new_E206_;
  assign new_E239_ = ~new_E221_ | new_E231_;
  assign new_E240_ = new_E221_ & new_E231_;
  assign new_E241_ = ~new_E221_ & ~new_E231_;
  assign new_E242_ = new_E263_ | new_E262_;
  assign new_E243_ = new_E209_ | new_E242_;
  assign new_E244_ = new_E267_ | new_E266_;
  assign new_E245_ = ~new_E209_ & new_E244_;
  assign new_E246_ = new_E265_ | new_E264_;
  assign new_E247_ = new_E209_ & new_E246_;
  assign new_E248_ = new_E207_ & ~new_E217_;
  assign new_E249_ = ~new_E207_ & new_E217_;
  assign new_E250_ = ~new_E206_ | ~new_E231_;
  assign new_E251_ = new_E217_ & new_E250_;
  assign new_E252_ = ~new_E217_ & ~new_E251_;
  assign new_E253_ = new_E217_ | new_E250_;
  assign new_E254_ = ~new_E207_ & new_E208_;
  assign new_E255_ = new_E207_ & ~new_E208_;
  assign new_E256_ = new_E224_ | new_E261_;
  assign new_E257_ = ~new_E224_ & ~new_E260_;
  assign new_E258_ = new_E207_ | new_E224_;
  assign new_E259_ = new_E207_ | new_E208_;
  assign new_E260_ = new_E224_ & new_E261_;
  assign new_E261_ = ~new_E206_ | ~new_E231_;
  assign new_E262_ = new_E239_ & new_E259_;
  assign new_E263_ = ~new_E239_ & ~new_E259_;
  assign new_E264_ = new_E268_ | new_E269_;
  assign new_E265_ = ~new_E210_ & new_E224_;
  assign new_E266_ = new_E270_ | new_E271_;
  assign new_E267_ = new_E210_ & new_E224_;
  assign new_E268_ = ~new_E210_ & ~new_E224_;
  assign new_E269_ = new_E210_ & ~new_E224_;
  assign new_E270_ = new_E210_ & ~new_E224_;
  assign new_E271_ = ~new_E210_ & new_E224_;
  assign new_E272_ = new_F6695_;
  assign new_E273_ = new_F6762_;
  assign new_E274_ = new_F6829_;
  assign new_E275_ = new_F6896_;
  assign new_E276_ = new_F6963_;
  assign new_E277_ = new_F7030_;
  assign new_E278_ = new_E285_ & new_E284_;
  assign new_E279_ = new_E287_ | new_E286_;
  assign new_E280_ = new_E289_ | new_E288_;
  assign new_E281_ = new_E291_ & new_E290_;
  assign new_E282_ = new_E291_ & new_E292_;
  assign new_E283_ = new_E284_ | new_E293_;
  assign new_E284_ = new_E273_ | new_E296_;
  assign new_E285_ = new_E295_ | new_E294_;
  assign new_E286_ = new_E300_ & new_E299_;
  assign new_E287_ = new_E298_ & new_E297_;
  assign new_E288_ = new_E303_ | new_E302_;
  assign new_E289_ = new_E298_ & new_E301_;
  assign new_E290_ = new_E273_ | new_E306_;
  assign new_E291_ = new_E305_ | new_E304_;
  assign new_E292_ = new_E308_ | new_E307_;
  assign new_E293_ = ~new_E284_ & new_E310_;
  assign new_E294_ = ~new_E286_ & new_E298_;
  assign new_E295_ = new_E286_ & ~new_E298_;
  assign new_E296_ = new_E272_ & ~new_E273_;
  assign new_E297_ = ~new_E319_ | ~new_E320_;
  assign new_E298_ = new_E312_ | new_E314_;
  assign new_E299_ = new_E322_ | new_E321_;
  assign new_E300_ = new_E316_ | new_E315_;
  assign new_E301_ = ~new_E324_ | ~new_E323_;
  assign new_E302_ = ~new_E325_ & new_E326_;
  assign new_E303_ = new_E325_ & ~new_E326_;
  assign new_E304_ = ~new_E272_ & new_E273_;
  assign new_E305_ = new_E272_ & ~new_E273_;
  assign new_E306_ = ~new_E288_ | new_E298_;
  assign new_E307_ = new_E288_ & new_E298_;
  assign new_E308_ = ~new_E288_ & ~new_E298_;
  assign new_E309_ = new_E330_ | new_E329_;
  assign new_E310_ = new_E276_ | new_E309_;
  assign new_E311_ = new_E334_ | new_E333_;
  assign new_E312_ = ~new_E276_ & new_E311_;
  assign new_E313_ = new_E332_ | new_E331_;
  assign new_E314_ = new_E276_ & new_E313_;
  assign new_E315_ = new_E274_ & ~new_E284_;
  assign new_E316_ = ~new_E274_ & new_E284_;
  assign new_E317_ = ~new_E273_ | ~new_E298_;
  assign new_E318_ = new_E284_ & new_E317_;
  assign new_E319_ = ~new_E284_ & ~new_E318_;
  assign new_E320_ = new_E284_ | new_E317_;
  assign new_E321_ = ~new_E274_ & new_E275_;
  assign new_E322_ = new_E274_ & ~new_E275_;
  assign new_E323_ = new_E291_ | new_E328_;
  assign new_E324_ = ~new_E291_ & ~new_E327_;
  assign new_E325_ = new_E274_ | new_E291_;
  assign new_E326_ = new_E274_ | new_E275_;
  assign new_E327_ = new_E291_ & new_E328_;
  assign new_E328_ = ~new_E273_ | ~new_E298_;
  assign new_E329_ = new_E306_ & new_E326_;
  assign new_E330_ = ~new_E306_ & ~new_E326_;
  assign new_E331_ = new_E335_ | new_E336_;
  assign new_E332_ = ~new_E277_ & new_E291_;
  assign new_E333_ = new_E337_ | new_E338_;
  assign new_E334_ = new_E277_ & new_E291_;
  assign new_E335_ = ~new_E277_ & ~new_E291_;
  assign new_E336_ = new_E277_ & ~new_E291_;
  assign new_E337_ = new_E277_ & ~new_E291_;
  assign new_E338_ = ~new_E277_ & new_E291_;
  assign new_E339_ = new_F7097_;
  assign new_E340_ = new_F7164_;
  assign new_E341_ = new_F7231_;
  assign new_E342_ = new_F7298_;
  assign new_E343_ = new_F7365_;
  assign new_E344_ = new_F7432_;
  assign new_E345_ = new_E352_ & new_E351_;
  assign new_E346_ = new_E354_ | new_E353_;
  assign new_E347_ = new_E356_ | new_E355_;
  assign new_E348_ = new_E358_ & new_E357_;
  assign new_E349_ = new_E358_ & new_E359_;
  assign new_E350_ = new_E351_ | new_E360_;
  assign new_E351_ = new_E340_ | new_E363_;
  assign new_E352_ = new_E362_ | new_E361_;
  assign new_E353_ = new_E367_ & new_E366_;
  assign new_E354_ = new_E365_ & new_E364_;
  assign new_E355_ = new_E370_ | new_E369_;
  assign new_E356_ = new_E365_ & new_E368_;
  assign new_E357_ = new_E340_ | new_E373_;
  assign new_E358_ = new_E372_ | new_E371_;
  assign new_E359_ = new_E375_ | new_E374_;
  assign new_E360_ = ~new_E351_ & new_E377_;
  assign new_E361_ = ~new_E353_ & new_E365_;
  assign new_E362_ = new_E353_ & ~new_E365_;
  assign new_E363_ = new_E339_ & ~new_E340_;
  assign new_E364_ = ~new_E386_ | ~new_E387_;
  assign new_E365_ = new_E379_ | new_E381_;
  assign new_E366_ = new_E389_ | new_E388_;
  assign new_E367_ = new_E383_ | new_E382_;
  assign new_E368_ = ~new_E391_ | ~new_E390_;
  assign new_E369_ = ~new_E392_ & new_E393_;
  assign new_E370_ = new_E392_ & ~new_E393_;
  assign new_E371_ = ~new_E339_ & new_E340_;
  assign new_E372_ = new_E339_ & ~new_E340_;
  assign new_E373_ = ~new_E355_ | new_E365_;
  assign new_E374_ = new_E355_ & new_E365_;
  assign new_E375_ = ~new_E355_ & ~new_E365_;
  assign new_E376_ = new_E397_ | new_E396_;
  assign new_E377_ = new_E343_ | new_E376_;
  assign new_E378_ = new_E401_ | new_E400_;
  assign new_E379_ = ~new_E343_ & new_E378_;
  assign new_E380_ = new_E399_ | new_E398_;
  assign new_E381_ = new_E343_ & new_E380_;
  assign new_E382_ = new_E341_ & ~new_E351_;
  assign new_E383_ = ~new_E341_ & new_E351_;
  assign new_E384_ = ~new_E340_ | ~new_E365_;
  assign new_E385_ = new_E351_ & new_E384_;
  assign new_E386_ = ~new_E351_ & ~new_E385_;
  assign new_E387_ = new_E351_ | new_E384_;
  assign new_E388_ = ~new_E341_ & new_E342_;
  assign new_E389_ = new_E341_ & ~new_E342_;
  assign new_E390_ = new_E358_ | new_E395_;
  assign new_E391_ = ~new_E358_ & ~new_E394_;
  assign new_E392_ = new_E341_ | new_E358_;
  assign new_E393_ = new_E341_ | new_E342_;
  assign new_E394_ = new_E358_ & new_E395_;
  assign new_E395_ = ~new_E340_ | ~new_E365_;
  assign new_E396_ = new_E373_ & new_E393_;
  assign new_E397_ = ~new_E373_ & ~new_E393_;
  assign new_E398_ = new_E402_ | new_E403_;
  assign new_E399_ = ~new_E344_ & new_E358_;
  assign new_E400_ = new_E404_ | new_E405_;
  assign new_E401_ = new_E344_ & new_E358_;
  assign new_E402_ = ~new_E344_ & ~new_E358_;
  assign new_E403_ = new_E344_ & ~new_E358_;
  assign new_E404_ = new_E344_ & ~new_E358_;
  assign new_E405_ = ~new_E344_ & new_E358_;
  assign new_E406_ = new_F7499_;
  assign new_E407_ = new_F7566_;
  assign new_E408_ = new_F7633_;
  assign new_E409_ = new_F7700_;
  assign new_E410_ = new_F7767_;
  assign new_E411_ = new_F7834_;
  assign new_E412_ = new_E419_ & new_E418_;
  assign new_E413_ = new_E421_ | new_E420_;
  assign new_E414_ = new_E423_ | new_E422_;
  assign new_E415_ = new_E425_ & new_E424_;
  assign new_E416_ = new_E425_ & new_E426_;
  assign new_E417_ = new_E418_ | new_E427_;
  assign new_E418_ = new_E407_ | new_E430_;
  assign new_E419_ = new_E429_ | new_E428_;
  assign new_E420_ = new_E434_ & new_E433_;
  assign new_E421_ = new_E432_ & new_E431_;
  assign new_E422_ = new_E437_ | new_E436_;
  assign new_E423_ = new_E432_ & new_E435_;
  assign new_E424_ = new_E407_ | new_E440_;
  assign new_E425_ = new_E439_ | new_E438_;
  assign new_E426_ = new_E442_ | new_E441_;
  assign new_E427_ = ~new_E418_ & new_E444_;
  assign new_E428_ = ~new_E420_ & new_E432_;
  assign new_E429_ = new_E420_ & ~new_E432_;
  assign new_E430_ = new_E406_ & ~new_E407_;
  assign new_E431_ = ~new_E453_ | ~new_E454_;
  assign new_E432_ = new_E446_ | new_E448_;
  assign new_E433_ = new_E456_ | new_E455_;
  assign new_E434_ = new_E450_ | new_E449_;
  assign new_E435_ = ~new_E458_ | ~new_E457_;
  assign new_E436_ = ~new_E459_ & new_E460_;
  assign new_E437_ = new_E459_ & ~new_E460_;
  assign new_E438_ = ~new_E406_ & new_E407_;
  assign new_E439_ = new_E406_ & ~new_E407_;
  assign new_E440_ = ~new_E422_ | new_E432_;
  assign new_E441_ = new_E422_ & new_E432_;
  assign new_E442_ = ~new_E422_ & ~new_E432_;
  assign new_E443_ = new_E464_ | new_E463_;
  assign new_E444_ = new_E410_ | new_E443_;
  assign new_E445_ = new_E468_ | new_E467_;
  assign new_E446_ = ~new_E410_ & new_E445_;
  assign new_E447_ = new_E466_ | new_E465_;
  assign new_E448_ = new_E410_ & new_E447_;
  assign new_E449_ = new_E408_ & ~new_E418_;
  assign new_E450_ = ~new_E408_ & new_E418_;
  assign new_E451_ = ~new_E407_ | ~new_E432_;
  assign new_E452_ = new_E418_ & new_E451_;
  assign new_E453_ = ~new_E418_ & ~new_E452_;
  assign new_E454_ = new_E418_ | new_E451_;
  assign new_E455_ = ~new_E408_ & new_E409_;
  assign new_E456_ = new_E408_ & ~new_E409_;
  assign new_E457_ = new_E425_ | new_E462_;
  assign new_E458_ = ~new_E425_ & ~new_E461_;
  assign new_E459_ = new_E408_ | new_E425_;
  assign new_E460_ = new_E408_ | new_E409_;
  assign new_E461_ = new_E425_ & new_E462_;
  assign new_E462_ = ~new_E407_ | ~new_E432_;
  assign new_E463_ = new_E440_ & new_E460_;
  assign new_E464_ = ~new_E440_ & ~new_E460_;
  assign new_E465_ = new_E469_ | new_E470_;
  assign new_E466_ = ~new_E411_ & new_E425_;
  assign new_E467_ = new_E471_ | new_E472_;
  assign new_E468_ = new_E411_ & new_E425_;
  assign new_E469_ = ~new_E411_ & ~new_E425_;
  assign new_E470_ = new_E411_ & ~new_E425_;
  assign new_E471_ = new_E411_ & ~new_E425_;
  assign new_E472_ = ~new_E411_ & new_E425_;
  assign new_E473_ = new_F7901_;
  assign new_E474_ = new_F7968_;
  assign new_E475_ = new_F8035_;
  assign new_E476_ = new_F8102_;
  assign new_E477_ = new_F8169_;
  assign new_E478_ = new_F8236_;
  assign new_E479_ = new_E486_ & new_E485_;
  assign new_E480_ = new_E488_ | new_E487_;
  assign new_E481_ = new_E490_ | new_E489_;
  assign new_E482_ = new_E492_ & new_E491_;
  assign new_E483_ = new_E492_ & new_E493_;
  assign new_E484_ = new_E485_ | new_E494_;
  assign new_E485_ = new_E474_ | new_E497_;
  assign new_E486_ = new_E496_ | new_E495_;
  assign new_E487_ = new_E501_ & new_E500_;
  assign new_E488_ = new_E499_ & new_E498_;
  assign new_E489_ = new_E504_ | new_E503_;
  assign new_E490_ = new_E499_ & new_E502_;
  assign new_E491_ = new_E474_ | new_E507_;
  assign new_E492_ = new_E506_ | new_E505_;
  assign new_E493_ = new_E509_ | new_E508_;
  assign new_E494_ = ~new_E485_ & new_E511_;
  assign new_E495_ = ~new_E487_ & new_E499_;
  assign new_E496_ = new_E487_ & ~new_E499_;
  assign new_E497_ = new_E473_ & ~new_E474_;
  assign new_E498_ = ~new_E520_ | ~new_E521_;
  assign new_E499_ = new_E513_ | new_E515_;
  assign new_E500_ = new_E523_ | new_E522_;
  assign new_E501_ = new_E517_ | new_E516_;
  assign new_E502_ = ~new_E525_ | ~new_E524_;
  assign new_E503_ = ~new_E526_ & new_E527_;
  assign new_E504_ = new_E526_ & ~new_E527_;
  assign new_E505_ = ~new_E473_ & new_E474_;
  assign new_E506_ = new_E473_ & ~new_E474_;
  assign new_E507_ = ~new_E489_ | new_E499_;
  assign new_E508_ = new_E489_ & new_E499_;
  assign new_E509_ = ~new_E489_ & ~new_E499_;
  assign new_E510_ = new_E531_ | new_E530_;
  assign new_E511_ = new_E477_ | new_E510_;
  assign new_E512_ = new_E535_ | new_E534_;
  assign new_E513_ = ~new_E477_ & new_E512_;
  assign new_E514_ = new_E533_ | new_E532_;
  assign new_E515_ = new_E477_ & new_E514_;
  assign new_E516_ = new_E475_ & ~new_E485_;
  assign new_E517_ = ~new_E475_ & new_E485_;
  assign new_E518_ = ~new_E474_ | ~new_E499_;
  assign new_E519_ = new_E485_ & new_E518_;
  assign new_E520_ = ~new_E485_ & ~new_E519_;
  assign new_E521_ = new_E485_ | new_E518_;
  assign new_E522_ = ~new_E475_ & new_E476_;
  assign new_E523_ = new_E475_ & ~new_E476_;
  assign new_E524_ = new_E492_ | new_E529_;
  assign new_E525_ = ~new_E492_ & ~new_E528_;
  assign new_E526_ = new_E475_ | new_E492_;
  assign new_E527_ = new_E475_ | new_E476_;
  assign new_E528_ = new_E492_ & new_E529_;
  assign new_E529_ = ~new_E474_ | ~new_E499_;
  assign new_E530_ = new_E507_ & new_E527_;
  assign new_E531_ = ~new_E507_ & ~new_E527_;
  assign new_E532_ = new_E536_ | new_E537_;
  assign new_E533_ = ~new_E478_ & new_E492_;
  assign new_E534_ = new_E538_ | new_E539_;
  assign new_E535_ = new_E478_ & new_E492_;
  assign new_E536_ = ~new_E478_ & ~new_E492_;
  assign new_E537_ = new_E478_ & ~new_E492_;
  assign new_E538_ = new_E478_ & ~new_E492_;
  assign new_E539_ = ~new_E478_ & new_E492_;
  assign new_E540_ = new_F8303_;
  assign new_E541_ = new_F8370_;
  assign new_E542_ = new_F8437_;
  assign new_E543_ = new_F8504_;
  assign new_E544_ = new_F8571_;
  assign new_E545_ = new_F8638_;
  assign new_E546_ = new_E553_ & new_E552_;
  assign new_E547_ = new_E555_ | new_E554_;
  assign new_E548_ = new_E557_ | new_E556_;
  assign new_E549_ = new_E559_ & new_E558_;
  assign new_E550_ = new_E559_ & new_E560_;
  assign new_E551_ = new_E552_ | new_E561_;
  assign new_E552_ = new_E541_ | new_E564_;
  assign new_E553_ = new_E563_ | new_E562_;
  assign new_E554_ = new_E568_ & new_E567_;
  assign new_E555_ = new_E566_ & new_E565_;
  assign new_E556_ = new_E571_ | new_E570_;
  assign new_E557_ = new_E566_ & new_E569_;
  assign new_E558_ = new_E541_ | new_E574_;
  assign new_E559_ = new_E573_ | new_E572_;
  assign new_E560_ = new_E576_ | new_E575_;
  assign new_E561_ = ~new_E552_ & new_E578_;
  assign new_E562_ = ~new_E554_ & new_E566_;
  assign new_E563_ = new_E554_ & ~new_E566_;
  assign new_E564_ = new_E540_ & ~new_E541_;
  assign new_E565_ = ~new_E587_ | ~new_E588_;
  assign new_E566_ = new_E580_ | new_E582_;
  assign new_E567_ = new_E590_ | new_E589_;
  assign new_E568_ = new_E584_ | new_E583_;
  assign new_E569_ = ~new_E592_ | ~new_E591_;
  assign new_E570_ = ~new_E593_ & new_E594_;
  assign new_E571_ = new_E593_ & ~new_E594_;
  assign new_E572_ = ~new_E540_ & new_E541_;
  assign new_E573_ = new_E540_ & ~new_E541_;
  assign new_E574_ = ~new_E556_ | new_E566_;
  assign new_E575_ = new_E556_ & new_E566_;
  assign new_E576_ = ~new_E556_ & ~new_E566_;
  assign new_E577_ = new_E598_ | new_E597_;
  assign new_E578_ = new_E544_ | new_E577_;
  assign new_E579_ = new_E602_ | new_E601_;
  assign new_E580_ = ~new_E544_ & new_E579_;
  assign new_E581_ = new_E600_ | new_E599_;
  assign new_E582_ = new_E544_ & new_E581_;
  assign new_E583_ = new_E542_ & ~new_E552_;
  assign new_E584_ = ~new_E542_ & new_E552_;
  assign new_E585_ = ~new_E541_ | ~new_E566_;
  assign new_E586_ = new_E552_ & new_E585_;
  assign new_E587_ = ~new_E552_ & ~new_E586_;
  assign new_E588_ = new_E552_ | new_E585_;
  assign new_E589_ = ~new_E542_ & new_E543_;
  assign new_E590_ = new_E542_ & ~new_E543_;
  assign new_E591_ = new_E559_ | new_E596_;
  assign new_E592_ = ~new_E559_ & ~new_E595_;
  assign new_E593_ = new_E542_ | new_E559_;
  assign new_E594_ = new_E542_ | new_E543_;
  assign new_E595_ = new_E559_ & new_E596_;
  assign new_E596_ = ~new_E541_ | ~new_E566_;
  assign new_E597_ = new_E574_ & new_E594_;
  assign new_E598_ = ~new_E574_ & ~new_E594_;
  assign new_E599_ = new_E603_ | new_E604_;
  assign new_E600_ = ~new_E545_ & new_E559_;
  assign new_E601_ = new_E605_ | new_E606_;
  assign new_E602_ = new_E545_ & new_E559_;
  assign new_E603_ = ~new_E545_ & ~new_E559_;
  assign new_E604_ = new_E545_ & ~new_E559_;
  assign new_E605_ = new_E545_ & ~new_E559_;
  assign new_E606_ = ~new_E545_ & new_E559_;
  assign new_E607_ = new_F8705_;
  assign new_E608_ = new_F8772_;
  assign new_E609_ = new_F8839_;
  assign new_E610_ = new_F8906_;
  assign new_E611_ = new_F8973_;
  assign new_E612_ = new_F9040_;
  assign new_E613_ = new_E620_ & new_E619_;
  assign new_E614_ = new_E622_ | new_E621_;
  assign new_E615_ = new_E624_ | new_E623_;
  assign new_E616_ = new_E626_ & new_E625_;
  assign new_E617_ = new_E626_ & new_E627_;
  assign new_E618_ = new_E619_ | new_E628_;
  assign new_E619_ = new_E608_ | new_E631_;
  assign new_E620_ = new_E630_ | new_E629_;
  assign new_E621_ = new_E635_ & new_E634_;
  assign new_E622_ = new_E633_ & new_E632_;
  assign new_E623_ = new_E638_ | new_E637_;
  assign new_E624_ = new_E633_ & new_E636_;
  assign new_E625_ = new_E608_ | new_E641_;
  assign new_E626_ = new_E640_ | new_E639_;
  assign new_E627_ = new_E643_ | new_E642_;
  assign new_E628_ = ~new_E619_ & new_E645_;
  assign new_E629_ = ~new_E621_ & new_E633_;
  assign new_E630_ = new_E621_ & ~new_E633_;
  assign new_E631_ = new_E607_ & ~new_E608_;
  assign new_E632_ = ~new_E654_ | ~new_E655_;
  assign new_E633_ = new_E647_ | new_E649_;
  assign new_E634_ = new_E657_ | new_E656_;
  assign new_E635_ = new_E651_ | new_E650_;
  assign new_E636_ = ~new_E659_ | ~new_E658_;
  assign new_E637_ = ~new_E660_ & new_E661_;
  assign new_E638_ = new_E660_ & ~new_E661_;
  assign new_E639_ = ~new_E607_ & new_E608_;
  assign new_E640_ = new_E607_ & ~new_E608_;
  assign new_E641_ = ~new_E623_ | new_E633_;
  assign new_E642_ = new_E623_ & new_E633_;
  assign new_E643_ = ~new_E623_ & ~new_E633_;
  assign new_E644_ = new_E665_ | new_E664_;
  assign new_E645_ = new_E611_ | new_E644_;
  assign new_E646_ = new_E669_ | new_E668_;
  assign new_E647_ = ~new_E611_ & new_E646_;
  assign new_E648_ = new_E667_ | new_E666_;
  assign new_E649_ = new_E611_ & new_E648_;
  assign new_E650_ = new_E609_ & ~new_E619_;
  assign new_E651_ = ~new_E609_ & new_E619_;
  assign new_E652_ = ~new_E608_ | ~new_E633_;
  assign new_E653_ = new_E619_ & new_E652_;
  assign new_E654_ = ~new_E619_ & ~new_E653_;
  assign new_E655_ = new_E619_ | new_E652_;
  assign new_E656_ = ~new_E609_ & new_E610_;
  assign new_E657_ = new_E609_ & ~new_E610_;
  assign new_E658_ = new_E626_ | new_E663_;
  assign new_E659_ = ~new_E626_ & ~new_E662_;
  assign new_E660_ = new_E609_ | new_E626_;
  assign new_E661_ = new_E609_ | new_E610_;
  assign new_E662_ = new_E626_ & new_E663_;
  assign new_E663_ = ~new_E608_ | ~new_E633_;
  assign new_E664_ = new_E641_ & new_E661_;
  assign new_E665_ = ~new_E641_ & ~new_E661_;
  assign new_E666_ = new_E670_ | new_E671_;
  assign new_E667_ = ~new_E612_ & new_E626_;
  assign new_E668_ = new_E672_ | new_E673_;
  assign new_E669_ = new_E612_ & new_E626_;
  assign new_E670_ = ~new_E612_ & ~new_E626_;
  assign new_E671_ = new_E612_ & ~new_E626_;
  assign new_E672_ = new_E612_ & ~new_E626_;
  assign new_E673_ = ~new_E612_ & new_E626_;
  assign new_E674_ = new_F9107_;
  assign new_E675_ = new_F9174_;
  assign new_E676_ = new_F9241_;
  assign new_E677_ = new_F9308_;
  assign new_E678_ = new_F9375_;
  assign new_E679_ = new_F9442_;
  assign new_E680_ = new_E687_ & new_E686_;
  assign new_E681_ = new_E689_ | new_E688_;
  assign new_E682_ = new_E691_ | new_E690_;
  assign new_E683_ = new_E693_ & new_E692_;
  assign new_E684_ = new_E693_ & new_E694_;
  assign new_E685_ = new_E686_ | new_E695_;
  assign new_E686_ = new_E675_ | new_E698_;
  assign new_E687_ = new_E697_ | new_E696_;
  assign new_E688_ = new_E702_ & new_E701_;
  assign new_E689_ = new_E700_ & new_E699_;
  assign new_E690_ = new_E705_ | new_E704_;
  assign new_E691_ = new_E700_ & new_E703_;
  assign new_E692_ = new_E675_ | new_E708_;
  assign new_E693_ = new_E707_ | new_E706_;
  assign new_E694_ = new_E710_ | new_E709_;
  assign new_E695_ = ~new_E686_ & new_E712_;
  assign new_E696_ = ~new_E688_ & new_E700_;
  assign new_E697_ = new_E688_ & ~new_E700_;
  assign new_E698_ = new_E674_ & ~new_E675_;
  assign new_E699_ = ~new_E721_ | ~new_E722_;
  assign new_E700_ = new_E714_ | new_E716_;
  assign new_E701_ = new_E724_ | new_E723_;
  assign new_E702_ = new_E718_ | new_E717_;
  assign new_E703_ = ~new_E726_ | ~new_E725_;
  assign new_E704_ = ~new_E727_ & new_E728_;
  assign new_E705_ = new_E727_ & ~new_E728_;
  assign new_E706_ = ~new_E674_ & new_E675_;
  assign new_E707_ = new_E674_ & ~new_E675_;
  assign new_E708_ = ~new_E690_ | new_E700_;
  assign new_E709_ = new_E690_ & new_E700_;
  assign new_E710_ = ~new_E690_ & ~new_E700_;
  assign new_E711_ = new_E732_ | new_E731_;
  assign new_E712_ = new_E678_ | new_E711_;
  assign new_E713_ = new_E736_ | new_E735_;
  assign new_E714_ = ~new_E678_ & new_E713_;
  assign new_E715_ = new_E734_ | new_E733_;
  assign new_E716_ = new_E678_ & new_E715_;
  assign new_E717_ = new_E676_ & ~new_E686_;
  assign new_E718_ = ~new_E676_ & new_E686_;
  assign new_E719_ = ~new_E675_ | ~new_E700_;
  assign new_E720_ = new_E686_ & new_E719_;
  assign new_E721_ = ~new_E686_ & ~new_E720_;
  assign new_E722_ = new_E686_ | new_E719_;
  assign new_E723_ = ~new_E676_ & new_E677_;
  assign new_E724_ = new_E676_ & ~new_E677_;
  assign new_E725_ = new_E693_ | new_E730_;
  assign new_E726_ = ~new_E693_ & ~new_E729_;
  assign new_E727_ = new_E676_ | new_E693_;
  assign new_E728_ = new_E676_ | new_E677_;
  assign new_E729_ = new_E693_ & new_E730_;
  assign new_E730_ = ~new_E675_ | ~new_E700_;
  assign new_E731_ = new_E708_ & new_E728_;
  assign new_E732_ = ~new_E708_ & ~new_E728_;
  assign new_E733_ = new_E737_ | new_E738_;
  assign new_E734_ = ~new_E679_ & new_E693_;
  assign new_E735_ = new_E739_ | new_E740_;
  assign new_E736_ = new_E679_ & new_E693_;
  assign new_E737_ = ~new_E679_ & ~new_E693_;
  assign new_E738_ = new_E679_ & ~new_E693_;
  assign new_E739_ = new_E679_ & ~new_E693_;
  assign new_E740_ = ~new_E679_ & new_E693_;
  assign new_E741_ = new_F9509_;
  assign new_E742_ = new_F9576_;
  assign new_E743_ = new_F9643_;
  assign new_E744_ = new_F9710_;
  assign new_E745_ = new_F9777_;
  assign new_E746_ = new_F9844_;
  assign new_E747_ = new_E754_ & new_E753_;
  assign new_E748_ = new_E756_ | new_E755_;
  assign new_E749_ = new_E758_ | new_E757_;
  assign new_E750_ = new_E760_ & new_E759_;
  assign new_E751_ = new_E760_ & new_E761_;
  assign new_E752_ = new_E753_ | new_E762_;
  assign new_E753_ = new_E742_ | new_E765_;
  assign new_E754_ = new_E764_ | new_E763_;
  assign new_E755_ = new_E769_ & new_E768_;
  assign new_E756_ = new_E767_ & new_E766_;
  assign new_E757_ = new_E772_ | new_E771_;
  assign new_E758_ = new_E767_ & new_E770_;
  assign new_E759_ = new_E742_ | new_E775_;
  assign new_E760_ = new_E774_ | new_E773_;
  assign new_E761_ = new_E777_ | new_E776_;
  assign new_E762_ = ~new_E753_ & new_E779_;
  assign new_E763_ = ~new_E755_ & new_E767_;
  assign new_E764_ = new_E755_ & ~new_E767_;
  assign new_E765_ = new_E741_ & ~new_E742_;
  assign new_E766_ = ~new_E788_ | ~new_E789_;
  assign new_E767_ = new_E781_ | new_E783_;
  assign new_E768_ = new_E791_ | new_E790_;
  assign new_E769_ = new_E785_ | new_E784_;
  assign new_E770_ = ~new_E793_ | ~new_E792_;
  assign new_E771_ = ~new_E794_ & new_E795_;
  assign new_E772_ = new_E794_ & ~new_E795_;
  assign new_E773_ = ~new_E741_ & new_E742_;
  assign new_E774_ = new_E741_ & ~new_E742_;
  assign new_E775_ = ~new_E757_ | new_E767_;
  assign new_E776_ = new_E757_ & new_E767_;
  assign new_E777_ = ~new_E757_ & ~new_E767_;
  assign new_E778_ = new_E799_ | new_E798_;
  assign new_E779_ = new_E745_ | new_E778_;
  assign new_E780_ = new_E803_ | new_E802_;
  assign new_E781_ = ~new_E745_ & new_E780_;
  assign new_E782_ = new_E801_ | new_E800_;
  assign new_E783_ = new_E745_ & new_E782_;
  assign new_E784_ = new_E743_ & ~new_E753_;
  assign new_E785_ = ~new_E743_ & new_E753_;
  assign new_E786_ = ~new_E742_ | ~new_E767_;
  assign new_E787_ = new_E753_ & new_E786_;
  assign new_E788_ = ~new_E753_ & ~new_E787_;
  assign new_E789_ = new_E753_ | new_E786_;
  assign new_E790_ = ~new_E743_ & new_E744_;
  assign new_E791_ = new_E743_ & ~new_E744_;
  assign new_E792_ = new_E760_ | new_E797_;
  assign new_E793_ = ~new_E760_ & ~new_E796_;
  assign new_E794_ = new_E743_ | new_E760_;
  assign new_E795_ = new_E743_ | new_E744_;
  assign new_E796_ = new_E760_ & new_E797_;
  assign new_E797_ = ~new_E742_ | ~new_E767_;
  assign new_E798_ = new_E775_ & new_E795_;
  assign new_E799_ = ~new_E775_ & ~new_E795_;
  assign new_E800_ = new_E804_ | new_E805_;
  assign new_E801_ = ~new_E746_ & new_E760_;
  assign new_E802_ = new_E806_ | new_E807_;
  assign new_E803_ = new_E746_ & new_E760_;
  assign new_E804_ = ~new_E746_ & ~new_E760_;
  assign new_E805_ = new_E746_ & ~new_E760_;
  assign new_E806_ = new_E746_ & ~new_E760_;
  assign new_E807_ = ~new_E746_ & new_E760_;
  assign new_E808_ = new_F9911_;
  assign new_E809_ = new_F9978_;
  assign new_E810_ = new_G46_;
  assign new_E811_ = new_G113_;
  assign new_E812_ = new_G180_;
  assign new_E813_ = new_G247_;
  assign new_E814_ = new_E821_ & new_E820_;
  assign new_E815_ = new_E823_ | new_E822_;
  assign new_E816_ = new_E825_ | new_E824_;
  assign new_E817_ = new_E827_ & new_E826_;
  assign new_E818_ = new_E827_ & new_E828_;
  assign new_E819_ = new_E820_ | new_E829_;
  assign new_E820_ = new_E809_ | new_E832_;
  assign new_E821_ = new_E831_ | new_E830_;
  assign new_E822_ = new_E836_ & new_E835_;
  assign new_E823_ = new_E834_ & new_E833_;
  assign new_E824_ = new_E839_ | new_E838_;
  assign new_E825_ = new_E834_ & new_E837_;
  assign new_E826_ = new_E809_ | new_E842_;
  assign new_E827_ = new_E841_ | new_E840_;
  assign new_E828_ = new_E844_ | new_E843_;
  assign new_E829_ = ~new_E820_ & new_E846_;
  assign new_E830_ = ~new_E822_ & new_E834_;
  assign new_E831_ = new_E822_ & ~new_E834_;
  assign new_E832_ = new_E808_ & ~new_E809_;
  assign new_E833_ = ~new_E855_ | ~new_E856_;
  assign new_E834_ = new_E848_ | new_E850_;
  assign new_E835_ = new_E858_ | new_E857_;
  assign new_E836_ = new_E852_ | new_E851_;
  assign new_E837_ = ~new_E860_ | ~new_E859_;
  assign new_E838_ = ~new_E861_ & new_E862_;
  assign new_E839_ = new_E861_ & ~new_E862_;
  assign new_E840_ = ~new_E808_ & new_E809_;
  assign new_E841_ = new_E808_ & ~new_E809_;
  assign new_E842_ = ~new_E824_ | new_E834_;
  assign new_E843_ = new_E824_ & new_E834_;
  assign new_E844_ = ~new_E824_ & ~new_E834_;
  assign new_E845_ = new_E866_ | new_E865_;
  assign new_E846_ = new_E812_ | new_E845_;
  assign new_E847_ = new_E870_ | new_E869_;
  assign new_E848_ = ~new_E812_ & new_E847_;
  assign new_E849_ = new_E868_ | new_E867_;
  assign new_E850_ = new_E812_ & new_E849_;
  assign new_E851_ = new_E810_ & ~new_E820_;
  assign new_E852_ = ~new_E810_ & new_E820_;
  assign new_E853_ = ~new_E809_ | ~new_E834_;
  assign new_E854_ = new_E820_ & new_E853_;
  assign new_E855_ = ~new_E820_ & ~new_E854_;
  assign new_E856_ = new_E820_ | new_E853_;
  assign new_E857_ = ~new_E810_ & new_E811_;
  assign new_E858_ = new_E810_ & ~new_E811_;
  assign new_E859_ = new_E827_ | new_E864_;
  assign new_E860_ = ~new_E827_ & ~new_E863_;
  assign new_E861_ = new_E810_ | new_E827_;
  assign new_E862_ = new_E810_ | new_E811_;
  assign new_E863_ = new_E827_ & new_E864_;
  assign new_E864_ = ~new_E809_ | ~new_E834_;
  assign new_E865_ = new_E842_ & new_E862_;
  assign new_E866_ = ~new_E842_ & ~new_E862_;
  assign new_E867_ = new_E871_ | new_E872_;
  assign new_E868_ = ~new_E813_ & new_E827_;
  assign new_E869_ = new_E873_ | new_E874_;
  assign new_E870_ = new_E813_ & new_E827_;
  assign new_E871_ = ~new_E813_ & ~new_E827_;
  assign new_E872_ = new_E813_ & ~new_E827_;
  assign new_E873_ = new_E813_ & ~new_E827_;
  assign new_E874_ = ~new_E813_ & new_E827_;
  assign new_E875_ = new_G314_;
  assign new_E876_ = new_G381_;
  assign new_E877_ = new_G448_;
  assign new_E878_ = new_G515_;
  assign new_E879_ = new_G582_;
  assign new_E880_ = new_G649_;
  assign new_E881_ = new_E888_ & new_E887_;
  assign new_E882_ = new_E890_ | new_E889_;
  assign new_E883_ = new_E892_ | new_E891_;
  assign new_E884_ = new_E894_ & new_E893_;
  assign new_E885_ = new_E894_ & new_E895_;
  assign new_E886_ = new_E887_ | new_E896_;
  assign new_E887_ = new_E876_ | new_E899_;
  assign new_E888_ = new_E898_ | new_E897_;
  assign new_E889_ = new_E903_ & new_E902_;
  assign new_E890_ = new_E901_ & new_E900_;
  assign new_E891_ = new_E906_ | new_E905_;
  assign new_E892_ = new_E901_ & new_E904_;
  assign new_E893_ = new_E876_ | new_E909_;
  assign new_E894_ = new_E908_ | new_E907_;
  assign new_E895_ = new_E911_ | new_E910_;
  assign new_E896_ = ~new_E887_ & new_E913_;
  assign new_E897_ = ~new_E889_ & new_E901_;
  assign new_E898_ = new_E889_ & ~new_E901_;
  assign new_E899_ = new_E875_ & ~new_E876_;
  assign new_E900_ = ~new_E922_ | ~new_E923_;
  assign new_E901_ = new_E915_ | new_E917_;
  assign new_E902_ = new_E925_ | new_E924_;
  assign new_E903_ = new_E919_ | new_E918_;
  assign new_E904_ = ~new_E927_ | ~new_E926_;
  assign new_E905_ = ~new_E928_ & new_E929_;
  assign new_E906_ = new_E928_ & ~new_E929_;
  assign new_E907_ = ~new_E875_ & new_E876_;
  assign new_E908_ = new_E875_ & ~new_E876_;
  assign new_E909_ = ~new_E891_ | new_E901_;
  assign new_E910_ = new_E891_ & new_E901_;
  assign new_E911_ = ~new_E891_ & ~new_E901_;
  assign new_E912_ = new_E933_ | new_E932_;
  assign new_E913_ = new_E879_ | new_E912_;
  assign new_E914_ = new_E937_ | new_E936_;
  assign new_E915_ = ~new_E879_ & new_E914_;
  assign new_E916_ = new_E935_ | new_E934_;
  assign new_E917_ = new_E879_ & new_E916_;
  assign new_E918_ = new_E877_ & ~new_E887_;
  assign new_E919_ = ~new_E877_ & new_E887_;
  assign new_E920_ = ~new_E876_ | ~new_E901_;
  assign new_E921_ = new_E887_ & new_E920_;
  assign new_E922_ = ~new_E887_ & ~new_E921_;
  assign new_E923_ = new_E887_ | new_E920_;
  assign new_E924_ = ~new_E877_ & new_E878_;
  assign new_E925_ = new_E877_ & ~new_E878_;
  assign new_E926_ = new_E894_ | new_E931_;
  assign new_E927_ = ~new_E894_ & ~new_E930_;
  assign new_E928_ = new_E877_ | new_E894_;
  assign new_E929_ = new_E877_ | new_E878_;
  assign new_E930_ = new_E894_ & new_E931_;
  assign new_E931_ = ~new_E876_ | ~new_E901_;
  assign new_E932_ = new_E909_ & new_E929_;
  assign new_E933_ = ~new_E909_ & ~new_E929_;
  assign new_E934_ = new_E938_ | new_E939_;
  assign new_E935_ = ~new_E880_ & new_E894_;
  assign new_E936_ = new_E940_ | new_E941_;
  assign new_E937_ = new_E880_ & new_E894_;
  assign new_E938_ = ~new_E880_ & ~new_E894_;
  assign new_E939_ = new_E880_ & ~new_E894_;
  assign new_E940_ = new_E880_ & ~new_E894_;
  assign new_E941_ = ~new_E880_ & new_E894_;
  assign new_E942_ = new_G716_;
  assign new_E943_ = new_G783_;
  assign new_E944_ = new_G850_;
  assign new_E945_ = new_G917_;
  assign new_E946_ = new_G984_;
  assign new_E947_ = new_G1051_;
  assign new_E948_ = new_E955_ & new_E954_;
  assign new_E949_ = new_E957_ | new_E956_;
  assign new_E950_ = new_E959_ | new_E958_;
  assign new_E951_ = new_E961_ & new_E960_;
  assign new_E952_ = new_E961_ & new_E962_;
  assign new_E953_ = new_E954_ | new_E963_;
  assign new_E954_ = new_E943_ | new_E966_;
  assign new_E955_ = new_E965_ | new_E964_;
  assign new_E956_ = new_E970_ & new_E969_;
  assign new_E957_ = new_E968_ & new_E967_;
  assign new_E958_ = new_E973_ | new_E972_;
  assign new_E959_ = new_E968_ & new_E971_;
  assign new_E960_ = new_E943_ | new_E976_;
  assign new_E961_ = new_E975_ | new_E974_;
  assign new_E962_ = new_E978_ | new_E977_;
  assign new_E963_ = ~new_E954_ & new_E980_;
  assign new_E964_ = ~new_E956_ & new_E968_;
  assign new_E965_ = new_E956_ & ~new_E968_;
  assign new_E966_ = new_E942_ & ~new_E943_;
  assign new_E967_ = ~new_E989_ | ~new_E990_;
  assign new_E968_ = new_E982_ | new_E984_;
  assign new_E969_ = new_E992_ | new_E991_;
  assign new_E970_ = new_E986_ | new_E985_;
  assign new_E971_ = ~new_E994_ | ~new_E993_;
  assign new_E972_ = ~new_E995_ & new_E996_;
  assign new_E973_ = new_E995_ & ~new_E996_;
  assign new_E974_ = ~new_E942_ & new_E943_;
  assign new_E975_ = new_E942_ & ~new_E943_;
  assign new_E976_ = ~new_E958_ | new_E968_;
  assign new_E977_ = new_E958_ & new_E968_;
  assign new_E978_ = ~new_E958_ & ~new_E968_;
  assign new_E979_ = new_E1000_ | new_E999_;
  assign new_E980_ = new_E946_ | new_E979_;
  assign new_E981_ = new_E1004_ | new_E1003_;
  assign new_E982_ = ~new_E946_ & new_E981_;
  assign new_E983_ = new_E1002_ | new_E1001_;
  assign new_E984_ = new_E946_ & new_E983_;
  assign new_E985_ = new_E944_ & ~new_E954_;
  assign new_E986_ = ~new_E944_ & new_E954_;
  assign new_E987_ = ~new_E943_ | ~new_E968_;
  assign new_E988_ = new_E954_ & new_E987_;
  assign new_E989_ = ~new_E954_ & ~new_E988_;
  assign new_E990_ = new_E954_ | new_E987_;
  assign new_E991_ = ~new_E944_ & new_E945_;
  assign new_E992_ = new_E944_ & ~new_E945_;
  assign new_E993_ = new_E961_ | new_E998_;
  assign new_E994_ = ~new_E961_ & ~new_E997_;
  assign new_E995_ = new_E944_ | new_E961_;
  assign new_E996_ = new_E944_ | new_E945_;
  assign new_E997_ = new_E961_ & new_E998_;
  assign new_E998_ = ~new_E943_ | ~new_E968_;
  assign new_E999_ = new_E976_ & new_E996_;
  assign new_E1000_ = ~new_E976_ & ~new_E996_;
  assign new_E1001_ = new_E1005_ | new_E1006_;
  assign new_E1002_ = ~new_E947_ & new_E961_;
  assign new_E1003_ = new_E1007_ | new_E1008_;
  assign new_E1004_ = new_E947_ & new_E961_;
  assign new_E1005_ = ~new_E947_ & ~new_E961_;
  assign new_E1006_ = new_E947_ & ~new_E961_;
  assign new_E1007_ = new_E947_ & ~new_E961_;
  assign new_E1008_ = ~new_E947_ & new_E961_;
  assign new_E1009_ = new_G1118_;
  assign new_E1010_ = new_G1185_;
  assign new_E1011_ = new_G1252_;
  assign new_E1012_ = new_G1319_;
  assign new_E1013_ = new_G1386_;
  assign new_E1014_ = new_G1453_;
  assign new_E1015_ = new_E1022_ & new_E1021_;
  assign new_E1016_ = new_E1024_ | new_E1023_;
  assign new_E1017_ = new_E1026_ | new_E1025_;
  assign new_E1018_ = new_E1028_ & new_E1027_;
  assign new_E1019_ = new_E1028_ & new_E1029_;
  assign new_E1020_ = new_E1021_ | new_E1030_;
  assign new_E1021_ = new_E1010_ | new_E1033_;
  assign new_E1022_ = new_E1032_ | new_E1031_;
  assign new_E1023_ = new_E1037_ & new_E1036_;
  assign new_E1024_ = new_E1035_ & new_E1034_;
  assign new_E1025_ = new_E1040_ | new_E1039_;
  assign new_E1026_ = new_E1035_ & new_E1038_;
  assign new_E1027_ = new_E1010_ | new_E1043_;
  assign new_E1028_ = new_E1042_ | new_E1041_;
  assign new_E1029_ = new_E1045_ | new_E1044_;
  assign new_E1030_ = ~new_E1021_ & new_E1047_;
  assign new_E1031_ = ~new_E1023_ & new_E1035_;
  assign new_E1032_ = new_E1023_ & ~new_E1035_;
  assign new_E1033_ = new_E1009_ & ~new_E1010_;
  assign new_E1034_ = ~new_E1056_ | ~new_E1057_;
  assign new_E1035_ = new_E1049_ | new_E1051_;
  assign new_E1036_ = new_E1059_ | new_E1058_;
  assign new_E1037_ = new_E1053_ | new_E1052_;
  assign new_E1038_ = ~new_E1061_ | ~new_E1060_;
  assign new_E1039_ = ~new_E1062_ & new_E1063_;
  assign new_E1040_ = new_E1062_ & ~new_E1063_;
  assign new_E1041_ = ~new_E1009_ & new_E1010_;
  assign new_E1042_ = new_E1009_ & ~new_E1010_;
  assign new_E1043_ = ~new_E1025_ | new_E1035_;
  assign new_E1044_ = new_E1025_ & new_E1035_;
  assign new_E1045_ = ~new_E1025_ & ~new_E1035_;
  assign new_E1046_ = new_E1067_ | new_E1066_;
  assign new_E1047_ = new_E1013_ | new_E1046_;
  assign new_E1048_ = new_E1071_ | new_E1070_;
  assign new_E1049_ = ~new_E1013_ & new_E1048_;
  assign new_E1050_ = new_E1069_ | new_E1068_;
  assign new_E1051_ = new_E1013_ & new_E1050_;
  assign new_E1052_ = new_E1011_ & ~new_E1021_;
  assign new_E1053_ = ~new_E1011_ & new_E1021_;
  assign new_E1054_ = ~new_E1010_ | ~new_E1035_;
  assign new_E1055_ = new_E1021_ & new_E1054_;
  assign new_E1056_ = ~new_E1021_ & ~new_E1055_;
  assign new_E1057_ = new_E1021_ | new_E1054_;
  assign new_E1058_ = ~new_E1011_ & new_E1012_;
  assign new_E1059_ = new_E1011_ & ~new_E1012_;
  assign new_E1060_ = new_E1028_ | new_E1065_;
  assign new_E1061_ = ~new_E1028_ & ~new_E1064_;
  assign new_E1062_ = new_E1011_ | new_E1028_;
  assign new_E1063_ = new_E1011_ | new_E1012_;
  assign new_E1064_ = new_E1028_ & new_E1065_;
  assign new_E1065_ = ~new_E1010_ | ~new_E1035_;
  assign new_E1066_ = new_E1043_ & new_E1063_;
  assign new_E1067_ = ~new_E1043_ & ~new_E1063_;
  assign new_E1068_ = new_E1072_ | new_E1073_;
  assign new_E1069_ = ~new_E1014_ & new_E1028_;
  assign new_E1070_ = new_E1074_ | new_E1075_;
  assign new_E1071_ = new_E1014_ & new_E1028_;
  assign new_E1072_ = ~new_E1014_ & ~new_E1028_;
  assign new_E1073_ = new_E1014_ & ~new_E1028_;
  assign new_E1074_ = new_E1014_ & ~new_E1028_;
  assign new_E1075_ = ~new_E1014_ & new_E1028_;
  assign new_E1076_ = new_G1520_;
  assign new_E1077_ = new_G1587_;
  assign new_E1078_ = new_G1654_;
  assign new_E1079_ = new_G1721_;
  assign new_E1080_ = new_G1788_;
  assign new_E1081_ = new_G1855_;
  assign new_E1082_ = new_E1089_ & new_E1088_;
  assign new_E1083_ = new_E1091_ | new_E1090_;
  assign new_E1084_ = new_E1093_ | new_E1092_;
  assign new_E1085_ = new_E1095_ & new_E1094_;
  assign new_E1086_ = new_E1095_ & new_E1096_;
  assign new_E1087_ = new_E1088_ | new_E1097_;
  assign new_E1088_ = new_E1077_ | new_E1100_;
  assign new_E1089_ = new_E1099_ | new_E1098_;
  assign new_E1090_ = new_E1104_ & new_E1103_;
  assign new_E1091_ = new_E1102_ & new_E1101_;
  assign new_E1092_ = new_E1107_ | new_E1106_;
  assign new_E1093_ = new_E1102_ & new_E1105_;
  assign new_E1094_ = new_E1077_ | new_E1110_;
  assign new_E1095_ = new_E1109_ | new_E1108_;
  assign new_E1096_ = new_E1112_ | new_E1111_;
  assign new_E1097_ = ~new_E1088_ & new_E1114_;
  assign new_E1098_ = ~new_E1090_ & new_E1102_;
  assign new_E1099_ = new_E1090_ & ~new_E1102_;
  assign new_E1100_ = new_E1076_ & ~new_E1077_;
  assign new_E1101_ = ~new_E1123_ | ~new_E1124_;
  assign new_E1102_ = new_E1116_ | new_E1118_;
  assign new_E1103_ = new_E1126_ | new_E1125_;
  assign new_E1104_ = new_E1120_ | new_E1119_;
  assign new_E1105_ = ~new_E1128_ | ~new_E1127_;
  assign new_E1106_ = ~new_E1129_ & new_E1130_;
  assign new_E1107_ = new_E1129_ & ~new_E1130_;
  assign new_E1108_ = ~new_E1076_ & new_E1077_;
  assign new_E1109_ = new_E1076_ & ~new_E1077_;
  assign new_E1110_ = ~new_E1092_ | new_E1102_;
  assign new_E1111_ = new_E1092_ & new_E1102_;
  assign new_E1112_ = ~new_E1092_ & ~new_E1102_;
  assign new_E1113_ = new_E1134_ | new_E1133_;
  assign new_E1114_ = new_E1080_ | new_E1113_;
  assign new_E1115_ = new_E1138_ | new_E1137_;
  assign new_E1116_ = ~new_E1080_ & new_E1115_;
  assign new_E1117_ = new_E1136_ | new_E1135_;
  assign new_E1118_ = new_E1080_ & new_E1117_;
  assign new_E1119_ = new_E1078_ & ~new_E1088_;
  assign new_E1120_ = ~new_E1078_ & new_E1088_;
  assign new_E1121_ = ~new_E1077_ | ~new_E1102_;
  assign new_E1122_ = new_E1088_ & new_E1121_;
  assign new_E1123_ = ~new_E1088_ & ~new_E1122_;
  assign new_E1124_ = new_E1088_ | new_E1121_;
  assign new_E1125_ = ~new_E1078_ & new_E1079_;
  assign new_E1126_ = new_E1078_ & ~new_E1079_;
  assign new_E1127_ = new_E1095_ | new_E1132_;
  assign new_E1128_ = ~new_E1095_ & ~new_E1131_;
  assign new_E1129_ = new_E1078_ | new_E1095_;
  assign new_E1130_ = new_E1078_ | new_E1079_;
  assign new_E1131_ = new_E1095_ & new_E1132_;
  assign new_E1132_ = ~new_E1077_ | ~new_E1102_;
  assign new_E1133_ = new_E1110_ & new_E1130_;
  assign new_E1134_ = ~new_E1110_ & ~new_E1130_;
  assign new_E1135_ = new_E1139_ | new_E1140_;
  assign new_E1136_ = ~new_E1081_ & new_E1095_;
  assign new_E1137_ = new_E1141_ | new_E1142_;
  assign new_E1138_ = new_E1081_ & new_E1095_;
  assign new_E1139_ = ~new_E1081_ & ~new_E1095_;
  assign new_E1140_ = new_E1081_ & ~new_E1095_;
  assign new_E1141_ = new_E1081_ & ~new_E1095_;
  assign new_E1142_ = ~new_E1081_ & new_E1095_;
  assign new_E1143_ = new_G1922_;
  assign new_E1144_ = new_G1989_;
  assign new_E1145_ = new_G2056_;
  assign new_E1146_ = new_G2123_;
  assign new_E1147_ = new_G2190_;
  assign new_E1148_ = new_G2257_;
  assign new_E1149_ = new_E1156_ & new_E1155_;
  assign new_E1150_ = new_E1158_ | new_E1157_;
  assign new_E1151_ = new_E1160_ | new_E1159_;
  assign new_E1152_ = new_E1162_ & new_E1161_;
  assign new_E1153_ = new_E1162_ & new_E1163_;
  assign new_E1154_ = new_E1155_ | new_E1164_;
  assign new_E1155_ = new_E1144_ | new_E1167_;
  assign new_E1156_ = new_E1166_ | new_E1165_;
  assign new_E1157_ = new_E1171_ & new_E1170_;
  assign new_E1158_ = new_E1169_ & new_E1168_;
  assign new_E1159_ = new_E1174_ | new_E1173_;
  assign new_E1160_ = new_E1169_ & new_E1172_;
  assign new_E1161_ = new_E1144_ | new_E1177_;
  assign new_E1162_ = new_E1176_ | new_E1175_;
  assign new_E1163_ = new_E1179_ | new_E1178_;
  assign new_E1164_ = ~new_E1155_ & new_E1181_;
  assign new_E1165_ = ~new_E1157_ & new_E1169_;
  assign new_E1166_ = new_E1157_ & ~new_E1169_;
  assign new_E1167_ = new_E1143_ & ~new_E1144_;
  assign new_E1168_ = ~new_E1190_ | ~new_E1191_;
  assign new_E1169_ = new_E1183_ | new_E1185_;
  assign new_E1170_ = new_E1193_ | new_E1192_;
  assign new_E1171_ = new_E1187_ | new_E1186_;
  assign new_E1172_ = ~new_E1195_ | ~new_E1194_;
  assign new_E1173_ = ~new_E1196_ & new_E1197_;
  assign new_E1174_ = new_E1196_ & ~new_E1197_;
  assign new_E1175_ = ~new_E1143_ & new_E1144_;
  assign new_E1176_ = new_E1143_ & ~new_E1144_;
  assign new_E1177_ = ~new_E1159_ | new_E1169_;
  assign new_E1178_ = new_E1159_ & new_E1169_;
  assign new_E1179_ = ~new_E1159_ & ~new_E1169_;
  assign new_E1180_ = new_E1201_ | new_E1200_;
  assign new_E1181_ = new_E1147_ | new_E1180_;
  assign new_E1182_ = new_E1205_ | new_E1204_;
  assign new_E1183_ = ~new_E1147_ & new_E1182_;
  assign new_E1184_ = new_E1203_ | new_E1202_;
  assign new_E1185_ = new_E1147_ & new_E1184_;
  assign new_E1186_ = new_E1145_ & ~new_E1155_;
  assign new_E1187_ = ~new_E1145_ & new_E1155_;
  assign new_E1188_ = ~new_E1144_ | ~new_E1169_;
  assign new_E1189_ = new_E1155_ & new_E1188_;
  assign new_E1190_ = ~new_E1155_ & ~new_E1189_;
  assign new_E1191_ = new_E1155_ | new_E1188_;
  assign new_E1192_ = ~new_E1145_ & new_E1146_;
  assign new_E1193_ = new_E1145_ & ~new_E1146_;
  assign new_E1194_ = new_E1162_ | new_E1199_;
  assign new_E1195_ = ~new_E1162_ & ~new_E1198_;
  assign new_E1196_ = new_E1145_ | new_E1162_;
  assign new_E1197_ = new_E1145_ | new_E1146_;
  assign new_E1198_ = new_E1162_ & new_E1199_;
  assign new_E1199_ = ~new_E1144_ | ~new_E1169_;
  assign new_E1200_ = new_E1177_ & new_E1197_;
  assign new_E1201_ = ~new_E1177_ & ~new_E1197_;
  assign new_E1202_ = new_E1206_ | new_E1207_;
  assign new_E1203_ = ~new_E1148_ & new_E1162_;
  assign new_E1204_ = new_E1208_ | new_E1209_;
  assign new_E1205_ = new_E1148_ & new_E1162_;
  assign new_E1206_ = ~new_E1148_ & ~new_E1162_;
  assign new_E1207_ = new_E1148_ & ~new_E1162_;
  assign new_E1208_ = new_E1148_ & ~new_E1162_;
  assign new_E1209_ = ~new_E1148_ & new_E1162_;
  assign new_E1210_ = new_G2324_;
  assign new_E1211_ = new_G2391_;
  assign new_E1212_ = new_G2458_;
  assign new_E1213_ = new_G2525_;
  assign new_E1214_ = new_G2592_;
  assign new_E1215_ = new_G2659_;
  assign new_E1216_ = new_E1223_ & new_E1222_;
  assign new_E1217_ = new_E1225_ | new_E1224_;
  assign new_E1218_ = new_E1227_ | new_E1226_;
  assign new_E1219_ = new_E1229_ & new_E1228_;
  assign new_E1220_ = new_E1229_ & new_E1230_;
  assign new_E1221_ = new_E1222_ | new_E1231_;
  assign new_E1222_ = new_E1211_ | new_E1234_;
  assign new_E1223_ = new_E1233_ | new_E1232_;
  assign new_E1224_ = new_E1238_ & new_E1237_;
  assign new_E1225_ = new_E1236_ & new_E1235_;
  assign new_E1226_ = new_E1241_ | new_E1240_;
  assign new_E1227_ = new_E1236_ & new_E1239_;
  assign new_E1228_ = new_E1211_ | new_E1244_;
  assign new_E1229_ = new_E1243_ | new_E1242_;
  assign new_E1230_ = new_E1246_ | new_E1245_;
  assign new_E1231_ = ~new_E1222_ & new_E1248_;
  assign new_E1232_ = ~new_E1224_ & new_E1236_;
  assign new_E1233_ = new_E1224_ & ~new_E1236_;
  assign new_E1234_ = new_E1210_ & ~new_E1211_;
  assign new_E1235_ = ~new_E1257_ | ~new_E1258_;
  assign new_E1236_ = new_E1250_ | new_E1252_;
  assign new_E1237_ = new_E1260_ | new_E1259_;
  assign new_E1238_ = new_E1254_ | new_E1253_;
  assign new_E1239_ = ~new_E1262_ | ~new_E1261_;
  assign new_E1240_ = ~new_E1263_ & new_E1264_;
  assign new_E1241_ = new_E1263_ & ~new_E1264_;
  assign new_E1242_ = ~new_E1210_ & new_E1211_;
  assign new_E1243_ = new_E1210_ & ~new_E1211_;
  assign new_E1244_ = ~new_E1226_ | new_E1236_;
  assign new_E1245_ = new_E1226_ & new_E1236_;
  assign new_E1246_ = ~new_E1226_ & ~new_E1236_;
  assign new_E1247_ = new_E1268_ | new_E1267_;
  assign new_E1248_ = new_E1214_ | new_E1247_;
  assign new_E1249_ = new_E1272_ | new_E1271_;
  assign new_E1250_ = ~new_E1214_ & new_E1249_;
  assign new_E1251_ = new_E1270_ | new_E1269_;
  assign new_E1252_ = new_E1214_ & new_E1251_;
  assign new_E1253_ = new_E1212_ & ~new_E1222_;
  assign new_E1254_ = ~new_E1212_ & new_E1222_;
  assign new_E1255_ = ~new_E1211_ | ~new_E1236_;
  assign new_E1256_ = new_E1222_ & new_E1255_;
  assign new_E1257_ = ~new_E1222_ & ~new_E1256_;
  assign new_E1258_ = new_E1222_ | new_E1255_;
  assign new_E1259_ = ~new_E1212_ & new_E1213_;
  assign new_E1260_ = new_E1212_ & ~new_E1213_;
  assign new_E1261_ = new_E1229_ | new_E1266_;
  assign new_E1262_ = ~new_E1229_ & ~new_E1265_;
  assign new_E1263_ = new_E1212_ | new_E1229_;
  assign new_E1264_ = new_E1212_ | new_E1213_;
  assign new_E1265_ = new_E1229_ & new_E1266_;
  assign new_E1266_ = ~new_E1211_ | ~new_E1236_;
  assign new_E1267_ = new_E1244_ & new_E1264_;
  assign new_E1268_ = ~new_E1244_ & ~new_E1264_;
  assign new_E1269_ = new_E1273_ | new_E1274_;
  assign new_E1270_ = ~new_E1215_ & new_E1229_;
  assign new_E1271_ = new_E1275_ | new_E1276_;
  assign new_E1272_ = new_E1215_ & new_E1229_;
  assign new_E1273_ = ~new_E1215_ & ~new_E1229_;
  assign new_E1274_ = new_E1215_ & ~new_E1229_;
  assign new_E1275_ = new_E1215_ & ~new_E1229_;
  assign new_E1276_ = ~new_E1215_ & new_E1229_;
  assign new_E1277_ = new_G2726_;
  assign new_E1278_ = new_G2793_;
  assign new_E1279_ = new_G2860_;
  assign new_E1280_ = new_G2927_;
  assign new_E1281_ = new_G2994_;
  assign new_E1282_ = new_G3061_;
  assign new_E1283_ = new_E1290_ & new_E1289_;
  assign new_E1284_ = new_E1292_ | new_E1291_;
  assign new_E1285_ = new_E1294_ | new_E1293_;
  assign new_E1286_ = new_E1296_ & new_E1295_;
  assign new_E1287_ = new_E1296_ & new_E1297_;
  assign new_E1288_ = new_E1289_ | new_E1298_;
  assign new_E1289_ = new_E1278_ | new_E1301_;
  assign new_E1290_ = new_E1300_ | new_E1299_;
  assign new_E1291_ = new_E1305_ & new_E1304_;
  assign new_E1292_ = new_E1303_ & new_E1302_;
  assign new_E1293_ = new_E1308_ | new_E1307_;
  assign new_E1294_ = new_E1303_ & new_E1306_;
  assign new_E1295_ = new_E1278_ | new_E1311_;
  assign new_E1296_ = new_E1310_ | new_E1309_;
  assign new_E1297_ = new_E1313_ | new_E1312_;
  assign new_E1298_ = ~new_E1289_ & new_E1315_;
  assign new_E1299_ = ~new_E1291_ & new_E1303_;
  assign new_E1300_ = new_E1291_ & ~new_E1303_;
  assign new_E1301_ = new_E1277_ & ~new_E1278_;
  assign new_E1302_ = ~new_E1324_ | ~new_E1325_;
  assign new_E1303_ = new_E1317_ | new_E1319_;
  assign new_E1304_ = new_E1327_ | new_E1326_;
  assign new_E1305_ = new_E1321_ | new_E1320_;
  assign new_E1306_ = ~new_E1329_ | ~new_E1328_;
  assign new_E1307_ = ~new_E1330_ & new_E1331_;
  assign new_E1308_ = new_E1330_ & ~new_E1331_;
  assign new_E1309_ = ~new_E1277_ & new_E1278_;
  assign new_E1310_ = new_E1277_ & ~new_E1278_;
  assign new_E1311_ = ~new_E1293_ | new_E1303_;
  assign new_E1312_ = new_E1293_ & new_E1303_;
  assign new_E1313_ = ~new_E1293_ & ~new_E1303_;
  assign new_E1314_ = new_E1335_ | new_E1334_;
  assign new_E1315_ = new_E1281_ | new_E1314_;
  assign new_E1316_ = new_E1339_ | new_E1338_;
  assign new_E1317_ = ~new_E1281_ & new_E1316_;
  assign new_E1318_ = new_E1337_ | new_E1336_;
  assign new_E1319_ = new_E1281_ & new_E1318_;
  assign new_E1320_ = new_E1279_ & ~new_E1289_;
  assign new_E1321_ = ~new_E1279_ & new_E1289_;
  assign new_E1322_ = ~new_E1278_ | ~new_E1303_;
  assign new_E1323_ = new_E1289_ & new_E1322_;
  assign new_E1324_ = ~new_E1289_ & ~new_E1323_;
  assign new_E1325_ = new_E1289_ | new_E1322_;
  assign new_E1326_ = ~new_E1279_ & new_E1280_;
  assign new_E1327_ = new_E1279_ & ~new_E1280_;
  assign new_E1328_ = new_E1296_ | new_E1333_;
  assign new_E1329_ = ~new_E1296_ & ~new_E1332_;
  assign new_E1330_ = new_E1279_ | new_E1296_;
  assign new_E1331_ = new_E1279_ | new_E1280_;
  assign new_E1332_ = new_E1296_ & new_E1333_;
  assign new_E1333_ = ~new_E1278_ | ~new_E1303_;
  assign new_E1334_ = new_E1311_ & new_E1331_;
  assign new_E1335_ = ~new_E1311_ & ~new_E1331_;
  assign new_E1336_ = new_E1340_ | new_E1341_;
  assign new_E1337_ = ~new_E1282_ & new_E1296_;
  assign new_E1338_ = new_E1342_ | new_E1343_;
  assign new_E1339_ = new_E1282_ & new_E1296_;
  assign new_E1340_ = ~new_E1282_ & ~new_E1296_;
  assign new_E1341_ = new_E1282_ & ~new_E1296_;
  assign new_E1342_ = new_E1282_ & ~new_E1296_;
  assign new_E1343_ = ~new_E1282_ & new_E1296_;
  assign new_E1344_ = new_G3128_;
  assign new_E1345_ = new_G3195_;
  assign new_E1346_ = new_G3262_;
  assign new_E1347_ = new_G3329_;
  assign new_E1348_ = new_G3396_;
  assign new_E1349_ = new_G3463_;
  assign new_E1350_ = new_E1357_ & new_E1356_;
  assign new_E1351_ = new_E1359_ | new_E1358_;
  assign new_E1352_ = new_E1361_ | new_E1360_;
  assign new_E1353_ = new_E1363_ & new_E1362_;
  assign new_E1354_ = new_E1363_ & new_E1364_;
  assign new_E1355_ = new_E1356_ | new_E1365_;
  assign new_E1356_ = new_E1345_ | new_E1368_;
  assign new_E1357_ = new_E1367_ | new_E1366_;
  assign new_E1358_ = new_E1372_ & new_E1371_;
  assign new_E1359_ = new_E1370_ & new_E1369_;
  assign new_E1360_ = new_E1375_ | new_E1374_;
  assign new_E1361_ = new_E1370_ & new_E1373_;
  assign new_E1362_ = new_E1345_ | new_E1378_;
  assign new_E1363_ = new_E1377_ | new_E1376_;
  assign new_E1364_ = new_E1380_ | new_E1379_;
  assign new_E1365_ = ~new_E1356_ & new_E1382_;
  assign new_E1366_ = ~new_E1358_ & new_E1370_;
  assign new_E1367_ = new_E1358_ & ~new_E1370_;
  assign new_E1368_ = new_E1344_ & ~new_E1345_;
  assign new_E1369_ = ~new_E1391_ | ~new_E1392_;
  assign new_E1370_ = new_E1384_ | new_E1386_;
  assign new_E1371_ = new_E1394_ | new_E1393_;
  assign new_E1372_ = new_E1388_ | new_E1387_;
  assign new_E1373_ = ~new_E1396_ | ~new_E1395_;
  assign new_E1374_ = ~new_E1397_ & new_E1398_;
  assign new_E1375_ = new_E1397_ & ~new_E1398_;
  assign new_E1376_ = ~new_E1344_ & new_E1345_;
  assign new_E1377_ = new_E1344_ & ~new_E1345_;
  assign new_E1378_ = ~new_E1360_ | new_E1370_;
  assign new_E1379_ = new_E1360_ & new_E1370_;
  assign new_E1380_ = ~new_E1360_ & ~new_E1370_;
  assign new_E1381_ = new_E1402_ | new_E1401_;
  assign new_E1382_ = new_E1348_ | new_E1381_;
  assign new_E1383_ = new_E1406_ | new_E1405_;
  assign new_E1384_ = ~new_E1348_ & new_E1383_;
  assign new_E1385_ = new_E1404_ | new_E1403_;
  assign new_E1386_ = new_E1348_ & new_E1385_;
  assign new_E1387_ = new_E1346_ & ~new_E1356_;
  assign new_E1388_ = ~new_E1346_ & new_E1356_;
  assign new_E1389_ = ~new_E1345_ | ~new_E1370_;
  assign new_E1390_ = new_E1356_ & new_E1389_;
  assign new_E1391_ = ~new_E1356_ & ~new_E1390_;
  assign new_E1392_ = new_E1356_ | new_E1389_;
  assign new_E1393_ = ~new_E1346_ & new_E1347_;
  assign new_E1394_ = new_E1346_ & ~new_E1347_;
  assign new_E1395_ = new_E1363_ | new_E1400_;
  assign new_E1396_ = ~new_E1363_ & ~new_E1399_;
  assign new_E1397_ = new_E1346_ | new_E1363_;
  assign new_E1398_ = new_E1346_ | new_E1347_;
  assign new_E1399_ = new_E1363_ & new_E1400_;
  assign new_E1400_ = ~new_E1345_ | ~new_E1370_;
  assign new_E1401_ = new_E1378_ & new_E1398_;
  assign new_E1402_ = ~new_E1378_ & ~new_E1398_;
  assign new_E1403_ = new_E1407_ | new_E1408_;
  assign new_E1404_ = ~new_E1349_ & new_E1363_;
  assign new_E1405_ = new_E1409_ | new_E1410_;
  assign new_E1406_ = new_E1349_ & new_E1363_;
  assign new_E1407_ = ~new_E1349_ & ~new_E1363_;
  assign new_E1408_ = new_E1349_ & ~new_E1363_;
  assign new_E1409_ = new_E1349_ & ~new_E1363_;
  assign new_E1410_ = ~new_E1349_ & new_E1363_;
  assign new_E1411_ = new_G3530_;
  assign new_E1412_ = new_G3597_;
  assign new_E1413_ = new_G3664_;
  assign new_E1414_ = new_G3731_;
  assign new_E1415_ = new_G3798_;
  assign new_E1416_ = new_G3865_;
  assign new_E1417_ = new_E1424_ & new_E1423_;
  assign new_E1418_ = new_E1426_ | new_E1425_;
  assign new_E1419_ = new_E1428_ | new_E1427_;
  assign new_E1420_ = new_E1430_ & new_E1429_;
  assign new_E1421_ = new_E1430_ & new_E1431_;
  assign new_E1422_ = new_E1423_ | new_E1432_;
  assign new_E1423_ = new_E1412_ | new_E1435_;
  assign new_E1424_ = new_E1434_ | new_E1433_;
  assign new_E1425_ = new_E1439_ & new_E1438_;
  assign new_E1426_ = new_E1437_ & new_E1436_;
  assign new_E1427_ = new_E1442_ | new_E1441_;
  assign new_E1428_ = new_E1437_ & new_E1440_;
  assign new_E1429_ = new_E1412_ | new_E1445_;
  assign new_E1430_ = new_E1444_ | new_E1443_;
  assign new_E1431_ = new_E1447_ | new_E1446_;
  assign new_E1432_ = ~new_E1423_ & new_E1449_;
  assign new_E1433_ = ~new_E1425_ & new_E1437_;
  assign new_E1434_ = new_E1425_ & ~new_E1437_;
  assign new_E1435_ = new_E1411_ & ~new_E1412_;
  assign new_E1436_ = ~new_E1458_ | ~new_E1459_;
  assign new_E1437_ = new_E1451_ | new_E1453_;
  assign new_E1438_ = new_E1461_ | new_E1460_;
  assign new_E1439_ = new_E1455_ | new_E1454_;
  assign new_E1440_ = ~new_E1463_ | ~new_E1462_;
  assign new_E1441_ = ~new_E1464_ & new_E1465_;
  assign new_E1442_ = new_E1464_ & ~new_E1465_;
  assign new_E1443_ = ~new_E1411_ & new_E1412_;
  assign new_E1444_ = new_E1411_ & ~new_E1412_;
  assign new_E1445_ = ~new_E1427_ | new_E1437_;
  assign new_E1446_ = new_E1427_ & new_E1437_;
  assign new_E1447_ = ~new_E1427_ & ~new_E1437_;
  assign new_E1448_ = new_E1469_ | new_E1468_;
  assign new_E1449_ = new_E1415_ | new_E1448_;
  assign new_E1450_ = new_E1473_ | new_E1472_;
  assign new_E1451_ = ~new_E1415_ & new_E1450_;
  assign new_E1452_ = new_E1471_ | new_E1470_;
  assign new_E1453_ = new_E1415_ & new_E1452_;
  assign new_E1454_ = new_E1413_ & ~new_E1423_;
  assign new_E1455_ = ~new_E1413_ & new_E1423_;
  assign new_E1456_ = ~new_E1412_ | ~new_E1437_;
  assign new_E1457_ = new_E1423_ & new_E1456_;
  assign new_E1458_ = ~new_E1423_ & ~new_E1457_;
  assign new_E1459_ = new_E1423_ | new_E1456_;
  assign new_E1460_ = ~new_E1413_ & new_E1414_;
  assign new_E1461_ = new_E1413_ & ~new_E1414_;
  assign new_E1462_ = new_E1430_ | new_E1467_;
  assign new_E1463_ = ~new_E1430_ & ~new_E1466_;
  assign new_E1464_ = new_E1413_ | new_E1430_;
  assign new_E1465_ = new_E1413_ | new_E1414_;
  assign new_E1466_ = new_E1430_ & new_E1467_;
  assign new_E1467_ = ~new_E1412_ | ~new_E1437_;
  assign new_E1468_ = new_E1445_ & new_E1465_;
  assign new_E1469_ = ~new_E1445_ & ~new_E1465_;
  assign new_E1470_ = new_E1474_ | new_E1475_;
  assign new_E1471_ = ~new_E1416_ & new_E1430_;
  assign new_E1472_ = new_E1476_ | new_E1477_;
  assign new_E1473_ = new_E1416_ & new_E1430_;
  assign new_E1474_ = ~new_E1416_ & ~new_E1430_;
  assign new_E1475_ = new_E1416_ & ~new_E1430_;
  assign new_E1476_ = new_E1416_ & ~new_E1430_;
  assign new_E1477_ = ~new_E1416_ & new_E1430_;
  assign new_E1478_ = new_G3932_;
  assign new_E1479_ = new_G3999_;
  assign new_E1480_ = new_G4066_;
  assign new_E1481_ = new_G4133_;
  assign new_E1482_ = new_G4200_;
  assign new_E1483_ = new_G4267_;
  assign new_E1484_ = new_E1491_ & new_E1490_;
  assign new_E1485_ = new_E1493_ | new_E1492_;
  assign new_E1486_ = new_E1495_ | new_E1494_;
  assign new_E1487_ = new_E1497_ & new_E1496_;
  assign new_E1488_ = new_E1497_ & new_E1498_;
  assign new_E1489_ = new_E1490_ | new_E1499_;
  assign new_E1490_ = new_E1479_ | new_E1502_;
  assign new_E1491_ = new_E1501_ | new_E1500_;
  assign new_E1492_ = new_E1506_ & new_E1505_;
  assign new_E1493_ = new_E1504_ & new_E1503_;
  assign new_E1494_ = new_E1509_ | new_E1508_;
  assign new_E1495_ = new_E1504_ & new_E1507_;
  assign new_E1496_ = new_E1479_ | new_E1512_;
  assign new_E1497_ = new_E1511_ | new_E1510_;
  assign new_E1498_ = new_E1514_ | new_E1513_;
  assign new_E1499_ = ~new_E1490_ & new_E1516_;
  assign new_E1500_ = ~new_E1492_ & new_E1504_;
  assign new_E1501_ = new_E1492_ & ~new_E1504_;
  assign new_E1502_ = new_E1478_ & ~new_E1479_;
  assign new_E1503_ = ~new_E1525_ | ~new_E1526_;
  assign new_E1504_ = new_E1518_ | new_E1520_;
  assign new_E1505_ = new_E1528_ | new_E1527_;
  assign new_E1506_ = new_E1522_ | new_E1521_;
  assign new_E1507_ = ~new_E1530_ | ~new_E1529_;
  assign new_E1508_ = ~new_E1531_ & new_E1532_;
  assign new_E1509_ = new_E1531_ & ~new_E1532_;
  assign new_E1510_ = ~new_E1478_ & new_E1479_;
  assign new_E1511_ = new_E1478_ & ~new_E1479_;
  assign new_E1512_ = ~new_E1494_ | new_E1504_;
  assign new_E1513_ = new_E1494_ & new_E1504_;
  assign new_E1514_ = ~new_E1494_ & ~new_E1504_;
  assign new_E1515_ = new_E1536_ | new_E1535_;
  assign new_E1516_ = new_E1482_ | new_E1515_;
  assign new_E1517_ = new_E1540_ | new_E1539_;
  assign new_E1518_ = ~new_E1482_ & new_E1517_;
  assign new_E1519_ = new_E1538_ | new_E1537_;
  assign new_E1520_ = new_E1482_ & new_E1519_;
  assign new_E1521_ = new_E1480_ & ~new_E1490_;
  assign new_E1522_ = ~new_E1480_ & new_E1490_;
  assign new_E1523_ = ~new_E1479_ | ~new_E1504_;
  assign new_E1524_ = new_E1490_ & new_E1523_;
  assign new_E1525_ = ~new_E1490_ & ~new_E1524_;
  assign new_E1526_ = new_E1490_ | new_E1523_;
  assign new_E1527_ = ~new_E1480_ & new_E1481_;
  assign new_E1528_ = new_E1480_ & ~new_E1481_;
  assign new_E1529_ = new_E1497_ | new_E1534_;
  assign new_E1530_ = ~new_E1497_ & ~new_E1533_;
  assign new_E1531_ = new_E1480_ | new_E1497_;
  assign new_E1532_ = new_E1480_ | new_E1481_;
  assign new_E1533_ = new_E1497_ & new_E1534_;
  assign new_E1534_ = ~new_E1479_ | ~new_E1504_;
  assign new_E1535_ = new_E1512_ & new_E1532_;
  assign new_E1536_ = ~new_E1512_ & ~new_E1532_;
  assign new_E1537_ = new_E1541_ | new_E1542_;
  assign new_E1538_ = ~new_E1483_ & new_E1497_;
  assign new_E1539_ = new_E1543_ | new_E1544_;
  assign new_E1540_ = new_E1483_ & new_E1497_;
  assign new_E1541_ = ~new_E1483_ & ~new_E1497_;
  assign new_E1542_ = new_E1483_ & ~new_E1497_;
  assign new_E1543_ = new_E1483_ & ~new_E1497_;
  assign new_E1544_ = ~new_E1483_ & new_E1497_;
  assign new_E1545_ = new_G4334_;
  assign new_E1546_ = new_G4401_;
  assign new_E1547_ = new_G4468_;
  assign new_E1548_ = new_G4535_;
  assign new_E1549_ = new_G4602_;
  assign new_E1550_ = new_G4669_;
  assign new_E1551_ = new_E1558_ & new_E1557_;
  assign new_E1552_ = new_E1560_ | new_E1559_;
  assign new_E1553_ = new_E1562_ | new_E1561_;
  assign new_E1554_ = new_E1564_ & new_E1563_;
  assign new_E1555_ = new_E1564_ & new_E1565_;
  assign new_E1556_ = new_E1557_ | new_E1566_;
  assign new_E1557_ = new_E1546_ | new_E1569_;
  assign new_E1558_ = new_E1568_ | new_E1567_;
  assign new_E1559_ = new_E1573_ & new_E1572_;
  assign new_E1560_ = new_E1571_ & new_E1570_;
  assign new_E1561_ = new_E1576_ | new_E1575_;
  assign new_E1562_ = new_E1571_ & new_E1574_;
  assign new_E1563_ = new_E1546_ | new_E1579_;
  assign new_E1564_ = new_E1578_ | new_E1577_;
  assign new_E1565_ = new_E1581_ | new_E1580_;
  assign new_E1566_ = ~new_E1557_ & new_E1583_;
  assign new_E1567_ = ~new_E1559_ & new_E1571_;
  assign new_E1568_ = new_E1559_ & ~new_E1571_;
  assign new_E1569_ = new_E1545_ & ~new_E1546_;
  assign new_E1570_ = ~new_E1592_ | ~new_E1593_;
  assign new_E1571_ = new_E1585_ | new_E1587_;
  assign new_E1572_ = new_E1595_ | new_E1594_;
  assign new_E1573_ = new_E1589_ | new_E1588_;
  assign new_E1574_ = ~new_E1597_ | ~new_E1596_;
  assign new_E1575_ = ~new_E1598_ & new_E1599_;
  assign new_E1576_ = new_E1598_ & ~new_E1599_;
  assign new_E1577_ = ~new_E1545_ & new_E1546_;
  assign new_E1578_ = new_E1545_ & ~new_E1546_;
  assign new_E1579_ = ~new_E1561_ | new_E1571_;
  assign new_E1580_ = new_E1561_ & new_E1571_;
  assign new_E1581_ = ~new_E1561_ & ~new_E1571_;
  assign new_E1582_ = new_E1603_ | new_E1602_;
  assign new_E1583_ = new_E1549_ | new_E1582_;
  assign new_E1584_ = new_E1607_ | new_E1606_;
  assign new_E1585_ = ~new_E1549_ & new_E1584_;
  assign new_E1586_ = new_E1605_ | new_E1604_;
  assign new_E1587_ = new_E1549_ & new_E1586_;
  assign new_E1588_ = new_E1547_ & ~new_E1557_;
  assign new_E1589_ = ~new_E1547_ & new_E1557_;
  assign new_E1590_ = ~new_E1546_ | ~new_E1571_;
  assign new_E1591_ = new_E1557_ & new_E1590_;
  assign new_E1592_ = ~new_E1557_ & ~new_E1591_;
  assign new_E1593_ = new_E1557_ | new_E1590_;
  assign new_E1594_ = ~new_E1547_ & new_E1548_;
  assign new_E1595_ = new_E1547_ & ~new_E1548_;
  assign new_E1596_ = new_E1564_ | new_E1601_;
  assign new_E1597_ = ~new_E1564_ & ~new_E1600_;
  assign new_E1598_ = new_E1547_ | new_E1564_;
  assign new_E1599_ = new_E1547_ | new_E1548_;
  assign new_E1600_ = new_E1564_ & new_E1601_;
  assign new_E1601_ = ~new_E1546_ | ~new_E1571_;
  assign new_E1602_ = new_E1579_ & new_E1599_;
  assign new_E1603_ = ~new_E1579_ & ~new_E1599_;
  assign new_E1604_ = new_E1608_ | new_E1609_;
  assign new_E1605_ = ~new_E1550_ & new_E1564_;
  assign new_E1606_ = new_E1610_ | new_E1611_;
  assign new_E1607_ = new_E1550_ & new_E1564_;
  assign new_E1608_ = ~new_E1550_ & ~new_E1564_;
  assign new_E1609_ = new_E1550_ & ~new_E1564_;
  assign new_E1610_ = new_E1550_ & ~new_E1564_;
  assign new_E1611_ = ~new_E1550_ & new_E1564_;
  assign new_E1612_ = new_G4736_;
  assign new_E1613_ = new_G4803_;
  assign new_E1614_ = new_G4870_;
  assign new_E1615_ = new_G4937_;
  assign new_E1616_ = new_G5004_;
  assign new_E1617_ = new_G5071_;
  assign new_E1618_ = new_E1625_ & new_E1624_;
  assign new_E1619_ = new_E1627_ | new_E1626_;
  assign new_E1620_ = new_E1629_ | new_E1628_;
  assign new_E1621_ = new_E1631_ & new_E1630_;
  assign new_E1622_ = new_E1631_ & new_E1632_;
  assign new_E1623_ = new_E1624_ | new_E1633_;
  assign new_E1624_ = new_E1613_ | new_E1636_;
  assign new_E1625_ = new_E1635_ | new_E1634_;
  assign new_E1626_ = new_E1640_ & new_E1639_;
  assign new_E1627_ = new_E1638_ & new_E1637_;
  assign new_E1628_ = new_E1643_ | new_E1642_;
  assign new_E1629_ = new_E1638_ & new_E1641_;
  assign new_E1630_ = new_E1613_ | new_E1646_;
  assign new_E1631_ = new_E1645_ | new_E1644_;
  assign new_E1632_ = new_E1648_ | new_E1647_;
  assign new_E1633_ = ~new_E1624_ & new_E1650_;
  assign new_E1634_ = ~new_E1626_ & new_E1638_;
  assign new_E1635_ = new_E1626_ & ~new_E1638_;
  assign new_E1636_ = new_E1612_ & ~new_E1613_;
  assign new_E1637_ = ~new_E1659_ | ~new_E1660_;
  assign new_E1638_ = new_E1652_ | new_E1654_;
  assign new_E1639_ = new_E1662_ | new_E1661_;
  assign new_E1640_ = new_E1656_ | new_E1655_;
  assign new_E1641_ = ~new_E1664_ | ~new_E1663_;
  assign new_E1642_ = ~new_E1665_ & new_E1666_;
  assign new_E1643_ = new_E1665_ & ~new_E1666_;
  assign new_E1644_ = ~new_E1612_ & new_E1613_;
  assign new_E1645_ = new_E1612_ & ~new_E1613_;
  assign new_E1646_ = ~new_E1628_ | new_E1638_;
  assign new_E1647_ = new_E1628_ & new_E1638_;
  assign new_E1648_ = ~new_E1628_ & ~new_E1638_;
  assign new_E1649_ = new_E1670_ | new_E1669_;
  assign new_E1650_ = new_E1616_ | new_E1649_;
  assign new_E1651_ = new_E1674_ | new_E1673_;
  assign new_E1652_ = ~new_E1616_ & new_E1651_;
  assign new_E1653_ = new_E1672_ | new_E1671_;
  assign new_E1654_ = new_E1616_ & new_E1653_;
  assign new_E1655_ = new_E1614_ & ~new_E1624_;
  assign new_E1656_ = ~new_E1614_ & new_E1624_;
  assign new_E1657_ = ~new_E1613_ | ~new_E1638_;
  assign new_E1658_ = new_E1624_ & new_E1657_;
  assign new_E1659_ = ~new_E1624_ & ~new_E1658_;
  assign new_E1660_ = new_E1624_ | new_E1657_;
  assign new_E1661_ = ~new_E1614_ & new_E1615_;
  assign new_E1662_ = new_E1614_ & ~new_E1615_;
  assign new_E1663_ = new_E1631_ | new_E1668_;
  assign new_E1664_ = ~new_E1631_ & ~new_E1667_;
  assign new_E1665_ = new_E1614_ | new_E1631_;
  assign new_E1666_ = new_E1614_ | new_E1615_;
  assign new_E1667_ = new_E1631_ & new_E1668_;
  assign new_E1668_ = ~new_E1613_ | ~new_E1638_;
  assign new_E1669_ = new_E1646_ & new_E1666_;
  assign new_E1670_ = ~new_E1646_ & ~new_E1666_;
  assign new_E1671_ = new_E1675_ | new_E1676_;
  assign new_E1672_ = ~new_E1617_ & new_E1631_;
  assign new_E1673_ = new_E1677_ | new_E1678_;
  assign new_E1674_ = new_E1617_ & new_E1631_;
  assign new_E1675_ = ~new_E1617_ & ~new_E1631_;
  assign new_E1676_ = new_E1617_ & ~new_E1631_;
  assign new_E1677_ = new_E1617_ & ~new_E1631_;
  assign new_E1678_ = ~new_E1617_ & new_E1631_;
  assign new_E1679_ = new_G5138_;
  assign new_E1680_ = new_G5205_;
  assign new_E1681_ = new_G5272_;
  assign new_E1682_ = new_G5339_;
  assign new_E1683_ = new_G5406_;
  assign new_E1684_ = new_G5473_;
  assign new_E1685_ = new_E1692_ & new_E1691_;
  assign new_E1686_ = new_E1694_ | new_E1693_;
  assign new_E1687_ = new_E1696_ | new_E1695_;
  assign new_E1688_ = new_E1698_ & new_E1697_;
  assign new_E1689_ = new_E1698_ & new_E1699_;
  assign new_E1690_ = new_E1691_ | new_E1700_;
  assign new_E1691_ = new_E1680_ | new_E1703_;
  assign new_E1692_ = new_E1702_ | new_E1701_;
  assign new_E1693_ = new_E1707_ & new_E1706_;
  assign new_E1694_ = new_E1705_ & new_E1704_;
  assign new_E1695_ = new_E1710_ | new_E1709_;
  assign new_E1696_ = new_E1705_ & new_E1708_;
  assign new_E1697_ = new_E1680_ | new_E1713_;
  assign new_E1698_ = new_E1712_ | new_E1711_;
  assign new_E1699_ = new_E1715_ | new_E1714_;
  assign new_E1700_ = ~new_E1691_ & new_E1717_;
  assign new_E1701_ = ~new_E1693_ & new_E1705_;
  assign new_E1702_ = new_E1693_ & ~new_E1705_;
  assign new_E1703_ = new_E1679_ & ~new_E1680_;
  assign new_E1704_ = ~new_E1726_ | ~new_E1727_;
  assign new_E1705_ = new_E1719_ | new_E1721_;
  assign new_E1706_ = new_E1729_ | new_E1728_;
  assign new_E1707_ = new_E1723_ | new_E1722_;
  assign new_E1708_ = ~new_E1731_ | ~new_E1730_;
  assign new_E1709_ = ~new_E1732_ & new_E1733_;
  assign new_E1710_ = new_E1732_ & ~new_E1733_;
  assign new_E1711_ = ~new_E1679_ & new_E1680_;
  assign new_E1712_ = new_E1679_ & ~new_E1680_;
  assign new_E1713_ = ~new_E1695_ | new_E1705_;
  assign new_E1714_ = new_E1695_ & new_E1705_;
  assign new_E1715_ = ~new_E1695_ & ~new_E1705_;
  assign new_E1716_ = new_E1737_ | new_E1736_;
  assign new_E1717_ = new_E1683_ | new_E1716_;
  assign new_E1718_ = new_E1741_ | new_E1740_;
  assign new_E1719_ = ~new_E1683_ & new_E1718_;
  assign new_E1720_ = new_E1739_ | new_E1738_;
  assign new_E1721_ = new_E1683_ & new_E1720_;
  assign new_E1722_ = new_E1681_ & ~new_E1691_;
  assign new_E1723_ = ~new_E1681_ & new_E1691_;
  assign new_E1724_ = ~new_E1680_ | ~new_E1705_;
  assign new_E1725_ = new_E1691_ & new_E1724_;
  assign new_E1726_ = ~new_E1691_ & ~new_E1725_;
  assign new_E1727_ = new_E1691_ | new_E1724_;
  assign new_E1728_ = ~new_E1681_ & new_E1682_;
  assign new_E1729_ = new_E1681_ & ~new_E1682_;
  assign new_E1730_ = new_E1698_ | new_E1735_;
  assign new_E1731_ = ~new_E1698_ & ~new_E1734_;
  assign new_E1732_ = new_E1681_ | new_E1698_;
  assign new_E1733_ = new_E1681_ | new_E1682_;
  assign new_E1734_ = new_E1698_ & new_E1735_;
  assign new_E1735_ = ~new_E1680_ | ~new_E1705_;
  assign new_E1736_ = new_E1713_ & new_E1733_;
  assign new_E1737_ = ~new_E1713_ & ~new_E1733_;
  assign new_E1738_ = new_E1742_ | new_E1743_;
  assign new_E1739_ = ~new_E1684_ & new_E1698_;
  assign new_E1740_ = new_E1744_ | new_E1745_;
  assign new_E1741_ = new_E1684_ & new_E1698_;
  assign new_E1742_ = ~new_E1684_ & ~new_E1698_;
  assign new_E1743_ = new_E1684_ & ~new_E1698_;
  assign new_E1744_ = new_E1684_ & ~new_E1698_;
  assign new_E1745_ = ~new_E1684_ & new_E1698_;
  assign new_E1746_ = new_G5540_;
  assign new_E1747_ = new_G5607_;
  assign new_E1748_ = new_G5674_;
  assign new_E1749_ = new_G5741_;
  assign new_E1750_ = new_G5808_;
  assign new_E1751_ = new_G5875_;
  assign new_E1752_ = new_E1759_ & new_E1758_;
  assign new_E1753_ = new_E1761_ | new_E1760_;
  assign new_E1754_ = new_E1763_ | new_E1762_;
  assign new_E1755_ = new_E1765_ & new_E1764_;
  assign new_E1756_ = new_E1765_ & new_E1766_;
  assign new_E1757_ = new_E1758_ | new_E1767_;
  assign new_E1758_ = new_E1747_ | new_E1770_;
  assign new_E1759_ = new_E1769_ | new_E1768_;
  assign new_E1760_ = new_E1774_ & new_E1773_;
  assign new_E1761_ = new_E1772_ & new_E1771_;
  assign new_E1762_ = new_E1777_ | new_E1776_;
  assign new_E1763_ = new_E1772_ & new_E1775_;
  assign new_E1764_ = new_E1747_ | new_E1780_;
  assign new_E1765_ = new_E1779_ | new_E1778_;
  assign new_E1766_ = new_E1782_ | new_E1781_;
  assign new_E1767_ = ~new_E1758_ & new_E1784_;
  assign new_E1768_ = ~new_E1760_ & new_E1772_;
  assign new_E1769_ = new_E1760_ & ~new_E1772_;
  assign new_E1770_ = new_E1746_ & ~new_E1747_;
  assign new_E1771_ = ~new_E1793_ | ~new_E1794_;
  assign new_E1772_ = new_E1786_ | new_E1788_;
  assign new_E1773_ = new_E1796_ | new_E1795_;
  assign new_E1774_ = new_E1790_ | new_E1789_;
  assign new_E1775_ = ~new_E1798_ | ~new_E1797_;
  assign new_E1776_ = ~new_E1799_ & new_E1800_;
  assign new_E1777_ = new_E1799_ & ~new_E1800_;
  assign new_E1778_ = ~new_E1746_ & new_E1747_;
  assign new_E1779_ = new_E1746_ & ~new_E1747_;
  assign new_E1780_ = ~new_E1762_ | new_E1772_;
  assign new_E1781_ = new_E1762_ & new_E1772_;
  assign new_E1782_ = ~new_E1762_ & ~new_E1772_;
  assign new_E1783_ = new_E1804_ | new_E1803_;
  assign new_E1784_ = new_E1750_ | new_E1783_;
  assign new_E1785_ = new_E1808_ | new_E1807_;
  assign new_E1786_ = ~new_E1750_ & new_E1785_;
  assign new_E1787_ = new_E1806_ | new_E1805_;
  assign new_E1788_ = new_E1750_ & new_E1787_;
  assign new_E1789_ = new_E1748_ & ~new_E1758_;
  assign new_E1790_ = ~new_E1748_ & new_E1758_;
  assign new_E1791_ = ~new_E1747_ | ~new_E1772_;
  assign new_E1792_ = new_E1758_ & new_E1791_;
  assign new_E1793_ = ~new_E1758_ & ~new_E1792_;
  assign new_E1794_ = new_E1758_ | new_E1791_;
  assign new_E1795_ = ~new_E1748_ & new_E1749_;
  assign new_E1796_ = new_E1748_ & ~new_E1749_;
  assign new_E1797_ = new_E1765_ | new_E1802_;
  assign new_E1798_ = ~new_E1765_ & ~new_E1801_;
  assign new_E1799_ = new_E1748_ | new_E1765_;
  assign new_E1800_ = new_E1748_ | new_E1749_;
  assign new_E1801_ = new_E1765_ & new_E1802_;
  assign new_E1802_ = ~new_E1747_ | ~new_E1772_;
  assign new_E1803_ = new_E1780_ & new_E1800_;
  assign new_E1804_ = ~new_E1780_ & ~new_E1800_;
  assign new_E1805_ = new_E1809_ | new_E1810_;
  assign new_E1806_ = ~new_E1751_ & new_E1765_;
  assign new_E1807_ = new_E1811_ | new_E1812_;
  assign new_E1808_ = new_E1751_ & new_E1765_;
  assign new_E1809_ = ~new_E1751_ & ~new_E1765_;
  assign new_E1810_ = new_E1751_ & ~new_E1765_;
  assign new_E1811_ = new_E1751_ & ~new_E1765_;
  assign new_E1812_ = ~new_E1751_ & new_E1765_;
  assign new_E1813_ = new_F1471_;
  assign new_E1814_ = new_F1537_;
  assign new_E1815_ = new_F1604_;
  assign new_E1816_ = new_F1671_;
  assign new_E1817_ = new_F1738_;
  assign new_E1818_ = new_F1805_;
  assign new_E1819_ = new_E1826_ & new_E1825_;
  assign new_E1820_ = new_E1828_ | new_E1827_;
  assign new_E1821_ = new_E1830_ | new_E1829_;
  assign new_E1822_ = new_E1832_ & new_E1831_;
  assign new_E1823_ = new_E1832_ & new_E1833_;
  assign new_E1824_ = new_E1825_ | new_E1834_;
  assign new_E1825_ = new_E1814_ | new_E1837_;
  assign new_E1826_ = new_E1836_ | new_E1835_;
  assign new_E1827_ = new_E1841_ & new_E1840_;
  assign new_E1828_ = new_E1839_ & new_E1838_;
  assign new_E1829_ = new_E1844_ | new_E1843_;
  assign new_E1830_ = new_E1839_ & new_E1842_;
  assign new_E1831_ = new_E1814_ | new_E1847_;
  assign new_E1832_ = new_E1846_ | new_E1845_;
  assign new_E1833_ = new_E1849_ | new_E1848_;
  assign new_E1834_ = ~new_E1825_ & new_E1851_;
  assign new_E1835_ = ~new_E1827_ & new_E1839_;
  assign new_E1836_ = new_E1827_ & ~new_E1839_;
  assign new_E1837_ = new_E1813_ & ~new_E1814_;
  assign new_E1838_ = ~new_E1860_ | ~new_E1861_;
  assign new_E1839_ = new_E1853_ | new_E1855_;
  assign new_E1840_ = new_E1863_ | new_E1862_;
  assign new_E1841_ = new_E1857_ | new_E1856_;
  assign new_E1842_ = ~new_E1865_ | ~new_E1864_;
  assign new_E1843_ = ~new_E1866_ & new_E1867_;
  assign new_E1844_ = new_E1866_ & ~new_E1867_;
  assign new_E1845_ = ~new_E1813_ & new_E1814_;
  assign new_E1846_ = new_E1813_ & ~new_E1814_;
  assign new_E1847_ = ~new_E1829_ | new_E1839_;
  assign new_E1848_ = new_E1829_ & new_E1839_;
  assign new_E1849_ = ~new_E1829_ & ~new_E1839_;
  assign new_E1850_ = new_E1871_ | new_E1870_;
  assign new_E1851_ = new_E1817_ | new_E1850_;
  assign new_E1852_ = new_E1875_ | new_E1874_;
  assign new_E1853_ = ~new_E1817_ & new_E1852_;
  assign new_E1854_ = new_E1873_ | new_E1872_;
  assign new_E1855_ = new_E1817_ & new_E1854_;
  assign new_E1856_ = new_E1815_ & ~new_E1825_;
  assign new_E1857_ = ~new_E1815_ & new_E1825_;
  assign new_E1858_ = ~new_E1814_ | ~new_E1839_;
  assign new_E1859_ = new_E1825_ & new_E1858_;
  assign new_E1860_ = ~new_E1825_ & ~new_E1859_;
  assign new_E1861_ = new_E1825_ | new_E1858_;
  assign new_E1862_ = ~new_E1815_ & new_E1816_;
  assign new_E1863_ = new_E1815_ & ~new_E1816_;
  assign new_E1864_ = new_E1832_ | new_E1869_;
  assign new_E1865_ = ~new_E1832_ & ~new_E1868_;
  assign new_E1866_ = new_E1815_ | new_E1832_;
  assign new_E1867_ = new_E1815_ | new_E1816_;
  assign new_E1868_ = new_E1832_ & new_E1869_;
  assign new_E1869_ = ~new_E1814_ | ~new_E1839_;
  assign new_E1870_ = new_E1847_ & new_E1867_;
  assign new_E1871_ = ~new_E1847_ & ~new_E1867_;
  assign new_E1872_ = new_E1876_ | new_E1877_;
  assign new_E1873_ = ~new_E1818_ & new_E1832_;
  assign new_E1874_ = new_E1878_ | new_E1879_;
  assign new_E1875_ = new_E1818_ & new_E1832_;
  assign new_E1876_ = ~new_E1818_ & ~new_E1832_;
  assign new_E1877_ = new_E1818_ & ~new_E1832_;
  assign new_E1878_ = new_E1818_ & ~new_E1832_;
  assign new_E1879_ = ~new_E1818_ & new_E1832_;
  assign new_E1880_ = new_F1872_;
  assign new_E1881_ = new_F1939_;
  assign new_E1882_ = new_F2006_;
  assign new_E1883_ = new_F2073_;
  assign new_E1884_ = new_F2140_;
  assign new_E1885_ = new_F2207_;
  assign new_E1886_ = new_E1893_ & new_E1892_;
  assign new_E1887_ = new_E1895_ | new_E1894_;
  assign new_E1888_ = new_E1897_ | new_E1896_;
  assign new_E1889_ = new_E1899_ & new_E1898_;
  assign new_E1890_ = new_E1899_ & new_E1900_;
  assign new_E1891_ = new_E1892_ | new_E1901_;
  assign new_E1892_ = new_E1881_ | new_E1904_;
  assign new_E1893_ = new_E1903_ | new_E1902_;
  assign new_E1894_ = new_E1908_ & new_E1907_;
  assign new_E1895_ = new_E1906_ & new_E1905_;
  assign new_E1896_ = new_E1911_ | new_E1910_;
  assign new_E1897_ = new_E1906_ & new_E1909_;
  assign new_E1898_ = new_E1881_ | new_E1914_;
  assign new_E1899_ = new_E1913_ | new_E1912_;
  assign new_E1900_ = new_E1916_ | new_E1915_;
  assign new_E1901_ = ~new_E1892_ & new_E1918_;
  assign new_E1902_ = ~new_E1894_ & new_E1906_;
  assign new_E1903_ = new_E1894_ & ~new_E1906_;
  assign new_E1904_ = new_E1880_ & ~new_E1881_;
  assign new_E1905_ = ~new_E1927_ | ~new_E1928_;
  assign new_E1906_ = new_E1920_ | new_E1922_;
  assign new_E1907_ = new_E1930_ | new_E1929_;
  assign new_E1908_ = new_E1924_ | new_E1923_;
  assign new_E1909_ = ~new_E1932_ | ~new_E1931_;
  assign new_E1910_ = ~new_E1933_ & new_E1934_;
  assign new_E1911_ = new_E1933_ & ~new_E1934_;
  assign new_E1912_ = ~new_E1880_ & new_E1881_;
  assign new_E1913_ = new_E1880_ & ~new_E1881_;
  assign new_E1914_ = ~new_E1896_ | new_E1906_;
  assign new_E1915_ = new_E1896_ & new_E1906_;
  assign new_E1916_ = ~new_E1896_ & ~new_E1906_;
  assign new_E1917_ = new_E1938_ | new_E1937_;
  assign new_E1918_ = new_E1884_ | new_E1917_;
  assign new_E1919_ = new_E1942_ | new_E1941_;
  assign new_E1920_ = ~new_E1884_ & new_E1919_;
  assign new_E1921_ = new_E1940_ | new_E1939_;
  assign new_E1922_ = new_E1884_ & new_E1921_;
  assign new_E1923_ = new_E1882_ & ~new_E1892_;
  assign new_E1924_ = ~new_E1882_ & new_E1892_;
  assign new_E1925_ = ~new_E1881_ | ~new_E1906_;
  assign new_E1926_ = new_E1892_ & new_E1925_;
  assign new_E1927_ = ~new_E1892_ & ~new_E1926_;
  assign new_E1928_ = new_E1892_ | new_E1925_;
  assign new_E1929_ = ~new_E1882_ & new_E1883_;
  assign new_E1930_ = new_E1882_ & ~new_E1883_;
  assign new_E1931_ = new_E1899_ | new_E1936_;
  assign new_E1932_ = ~new_E1899_ & ~new_E1935_;
  assign new_E1933_ = new_E1882_ | new_E1899_;
  assign new_E1934_ = new_E1882_ | new_E1883_;
  assign new_E1935_ = new_E1899_ & new_E1936_;
  assign new_E1936_ = ~new_E1881_ | ~new_E1906_;
  assign new_E1937_ = new_E1914_ & new_E1934_;
  assign new_E1938_ = ~new_E1914_ & ~new_E1934_;
  assign new_E1939_ = new_E1943_ | new_E1944_;
  assign new_E1940_ = ~new_E1885_ & new_E1899_;
  assign new_E1941_ = new_E1945_ | new_E1946_;
  assign new_E1942_ = new_E1885_ & new_E1899_;
  assign new_E1943_ = ~new_E1885_ & ~new_E1899_;
  assign new_E1944_ = new_E1885_ & ~new_E1899_;
  assign new_E1945_ = new_E1885_ & ~new_E1899_;
  assign new_E1946_ = ~new_E1885_ & new_E1899_;
  assign new_E1947_ = new_F2274_;
  assign new_E1948_ = new_F2341_;
  assign new_E1949_ = new_F2408_;
  assign new_E1950_ = new_F2475_;
  assign new_E1951_ = new_F2542_;
  assign new_E1952_ = new_F2609_;
  assign new_E1953_ = new_E1960_ & new_E1959_;
  assign new_E1954_ = new_E1962_ | new_E1961_;
  assign new_E1955_ = new_E1964_ | new_E1963_;
  assign new_E1956_ = new_E1966_ & new_E1965_;
  assign new_E1957_ = new_E1966_ & new_E1967_;
  assign new_E1958_ = new_E1959_ | new_E1968_;
  assign new_E1959_ = new_E1948_ | new_E1971_;
  assign new_E1960_ = new_E1970_ | new_E1969_;
  assign new_E1961_ = new_E1975_ & new_E1974_;
  assign new_E1962_ = new_E1973_ & new_E1972_;
  assign new_E1963_ = new_E1978_ | new_E1977_;
  assign new_E1964_ = new_E1973_ & new_E1976_;
  assign new_E1965_ = new_E1948_ | new_E1981_;
  assign new_E1966_ = new_E1980_ | new_E1979_;
  assign new_E1967_ = new_E1983_ | new_E1982_;
  assign new_E1968_ = ~new_E1959_ & new_E1985_;
  assign new_E1969_ = ~new_E1961_ & new_E1973_;
  assign new_E1970_ = new_E1961_ & ~new_E1973_;
  assign new_E1971_ = new_E1947_ & ~new_E1948_;
  assign new_E1972_ = ~new_E1994_ | ~new_E1995_;
  assign new_E1973_ = new_E1987_ | new_E1989_;
  assign new_E1974_ = new_E1997_ | new_E1996_;
  assign new_E1975_ = new_E1991_ | new_E1990_;
  assign new_E1976_ = ~new_E1999_ | ~new_E1998_;
  assign new_E1977_ = ~new_E2000_ & new_E2001_;
  assign new_E1978_ = new_E2000_ & ~new_E2001_;
  assign new_E1979_ = ~new_E1947_ & new_E1948_;
  assign new_E1980_ = new_E1947_ & ~new_E1948_;
  assign new_E1981_ = ~new_E1963_ | new_E1973_;
  assign new_E1982_ = new_E1963_ & new_E1973_;
  assign new_E1983_ = ~new_E1963_ & ~new_E1973_;
  assign new_E1984_ = new_E2005_ | new_E2004_;
  assign new_E1985_ = new_E1951_ | new_E1984_;
  assign new_E1986_ = new_E2009_ | new_E2008_;
  assign new_E1987_ = ~new_E1951_ & new_E1986_;
  assign new_E1988_ = new_E2007_ | new_E2006_;
  assign new_E1989_ = new_E1951_ & new_E1988_;
  assign new_E1990_ = new_E1949_ & ~new_E1959_;
  assign new_E1991_ = ~new_E1949_ & new_E1959_;
  assign new_E1992_ = ~new_E1948_ | ~new_E1973_;
  assign new_E1993_ = new_E1959_ & new_E1992_;
  assign new_E1994_ = ~new_E1959_ & ~new_E1993_;
  assign new_E1995_ = new_E1959_ | new_E1992_;
  assign new_E1996_ = ~new_E1949_ & new_E1950_;
  assign new_E1997_ = new_E1949_ & ~new_E1950_;
  assign new_E1998_ = new_E1966_ | new_E2003_;
  assign new_E1999_ = ~new_E1966_ & ~new_E2002_;
  assign new_E2000_ = new_E1949_ | new_E1966_;
  assign new_E2001_ = new_E1949_ | new_E1950_;
  assign new_E2002_ = new_E1966_ & new_E2003_;
  assign new_E2003_ = ~new_E1948_ | ~new_E1973_;
  assign new_E2004_ = new_E1981_ & new_E2001_;
  assign new_E2005_ = ~new_E1981_ & ~new_E2001_;
  assign new_E2006_ = new_E2010_ | new_E2011_;
  assign new_E2007_ = ~new_E1952_ & new_E1966_;
  assign new_E2008_ = new_E2012_ | new_E2013_;
  assign new_E2009_ = new_E1952_ & new_E1966_;
  assign new_E2010_ = ~new_E1952_ & ~new_E1966_;
  assign new_E2011_ = new_E1952_ & ~new_E1966_;
  assign new_E2012_ = new_E1952_ & ~new_E1966_;
  assign new_E2013_ = ~new_E1952_ & new_E1966_;
  assign new_E2014_ = new_F2676_;
  assign new_E2015_ = new_F2743_;
  assign new_E2016_ = new_F2810_;
  assign new_E2017_ = new_F2877_;
  assign new_E2018_ = new_F2944_;
  assign new_E2019_ = new_F3011_;
  assign new_E2020_ = new_E2027_ & new_E2026_;
  assign new_E2021_ = new_E2029_ | new_E2028_;
  assign new_E2022_ = new_E2031_ | new_E2030_;
  assign new_E2023_ = new_E2033_ & new_E2032_;
  assign new_E2024_ = new_E2033_ & new_E2034_;
  assign new_E2025_ = new_E2026_ | new_E2035_;
  assign new_E2026_ = new_E2015_ | new_E2038_;
  assign new_E2027_ = new_E2037_ | new_E2036_;
  assign new_E2028_ = new_E2042_ & new_E2041_;
  assign new_E2029_ = new_E2040_ & new_E2039_;
  assign new_E2030_ = new_E2045_ | new_E2044_;
  assign new_E2031_ = new_E2040_ & new_E2043_;
  assign new_E2032_ = new_E2015_ | new_E2048_;
  assign new_E2033_ = new_E2047_ | new_E2046_;
  assign new_E2034_ = new_E2050_ | new_E2049_;
  assign new_E2035_ = ~new_E2026_ & new_E2052_;
  assign new_E2036_ = ~new_E2028_ & new_E2040_;
  assign new_E2037_ = new_E2028_ & ~new_E2040_;
  assign new_E2038_ = new_E2014_ & ~new_E2015_;
  assign new_E2039_ = ~new_E2061_ | ~new_E2062_;
  assign new_E2040_ = new_E2054_ | new_E2056_;
  assign new_E2041_ = new_E2064_ | new_E2063_;
  assign new_E2042_ = new_E2058_ | new_E2057_;
  assign new_E2043_ = ~new_E2066_ | ~new_E2065_;
  assign new_E2044_ = ~new_E2067_ & new_E2068_;
  assign new_E2045_ = new_E2067_ & ~new_E2068_;
  assign new_E2046_ = ~new_E2014_ & new_E2015_;
  assign new_E2047_ = new_E2014_ & ~new_E2015_;
  assign new_E2048_ = ~new_E2030_ | new_E2040_;
  assign new_E2049_ = new_E2030_ & new_E2040_;
  assign new_E2050_ = ~new_E2030_ & ~new_E2040_;
  assign new_E2051_ = new_E2072_ | new_E2071_;
  assign new_E2052_ = new_E2018_ | new_E2051_;
  assign new_E2053_ = new_E2076_ | new_E2075_;
  assign new_E2054_ = ~new_E2018_ & new_E2053_;
  assign new_E2055_ = new_E2074_ | new_E2073_;
  assign new_E2056_ = new_E2018_ & new_E2055_;
  assign new_E2057_ = new_E2016_ & ~new_E2026_;
  assign new_E2058_ = ~new_E2016_ & new_E2026_;
  assign new_E2059_ = ~new_E2015_ | ~new_E2040_;
  assign new_E2060_ = new_E2026_ & new_E2059_;
  assign new_E2061_ = ~new_E2026_ & ~new_E2060_;
  assign new_E2062_ = new_E2026_ | new_E2059_;
  assign new_E2063_ = ~new_E2016_ & new_E2017_;
  assign new_E2064_ = new_E2016_ & ~new_E2017_;
  assign new_E2065_ = new_E2033_ | new_E2070_;
  assign new_E2066_ = ~new_E2033_ & ~new_E2069_;
  assign new_E2067_ = new_E2016_ | new_E2033_;
  assign new_E2068_ = new_E2016_ | new_E2017_;
  assign new_E2069_ = new_E2033_ & new_E2070_;
  assign new_E2070_ = ~new_E2015_ | ~new_E2040_;
  assign new_E2071_ = new_E2048_ & new_E2068_;
  assign new_E2072_ = ~new_E2048_ & ~new_E2068_;
  assign new_E2073_ = new_E2077_ | new_E2078_;
  assign new_E2074_ = ~new_E2019_ & new_E2033_;
  assign new_E2075_ = new_E2079_ | new_E2080_;
  assign new_E2076_ = new_E2019_ & new_E2033_;
  assign new_E2077_ = ~new_E2019_ & ~new_E2033_;
  assign new_E2078_ = new_E2019_ & ~new_E2033_;
  assign new_E2079_ = new_E2019_ & ~new_E2033_;
  assign new_E2080_ = ~new_E2019_ & new_E2033_;
  assign new_E2081_ = new_F3078_;
  assign new_E2082_ = new_F3145_;
  assign new_E2083_ = new_F3212_;
  assign new_E2084_ = new_F3279_;
  assign new_E2085_ = new_F3346_;
  assign new_E2086_ = new_F3413_;
  assign new_E2087_ = new_E2094_ & new_E2093_;
  assign new_E2088_ = new_E2096_ | new_E2095_;
  assign new_E2089_ = new_E2098_ | new_E2097_;
  assign new_E2090_ = new_E2100_ & new_E2099_;
  assign new_E2091_ = new_E2100_ & new_E2101_;
  assign new_E2092_ = new_E2093_ | new_E2102_;
  assign new_E2093_ = new_E2082_ | new_E2105_;
  assign new_E2094_ = new_E2104_ | new_E2103_;
  assign new_E2095_ = new_E2109_ & new_E2108_;
  assign new_E2096_ = new_E2107_ & new_E2106_;
  assign new_E2097_ = new_E2112_ | new_E2111_;
  assign new_E2098_ = new_E2107_ & new_E2110_;
  assign new_E2099_ = new_E2082_ | new_E2115_;
  assign new_E2100_ = new_E2114_ | new_E2113_;
  assign new_E2101_ = new_E2117_ | new_E2116_;
  assign new_E2102_ = ~new_E2093_ & new_E2119_;
  assign new_E2103_ = ~new_E2095_ & new_E2107_;
  assign new_E2104_ = new_E2095_ & ~new_E2107_;
  assign new_E2105_ = new_E2081_ & ~new_E2082_;
  assign new_E2106_ = ~new_E2128_ | ~new_E2129_;
  assign new_E2107_ = new_E2121_ | new_E2123_;
  assign new_E2108_ = new_E2131_ | new_E2130_;
  assign new_E2109_ = new_E2125_ | new_E2124_;
  assign new_E2110_ = ~new_E2133_ | ~new_E2132_;
  assign new_E2111_ = ~new_E2134_ & new_E2135_;
  assign new_E2112_ = new_E2134_ & ~new_E2135_;
  assign new_E2113_ = ~new_E2081_ & new_E2082_;
  assign new_E2114_ = new_E2081_ & ~new_E2082_;
  assign new_E2115_ = ~new_E2097_ | new_E2107_;
  assign new_E2116_ = new_E2097_ & new_E2107_;
  assign new_E2117_ = ~new_E2097_ & ~new_E2107_;
  assign new_E2118_ = new_E2139_ | new_E2138_;
  assign new_E2119_ = new_E2085_ | new_E2118_;
  assign new_E2120_ = new_E2143_ | new_E2142_;
  assign new_E2121_ = ~new_E2085_ & new_E2120_;
  assign new_E2122_ = new_E2141_ | new_E2140_;
  assign new_E2123_ = new_E2085_ & new_E2122_;
  assign new_E2124_ = new_E2083_ & ~new_E2093_;
  assign new_E2125_ = ~new_E2083_ & new_E2093_;
  assign new_E2126_ = ~new_E2082_ | ~new_E2107_;
  assign new_E2127_ = new_E2093_ & new_E2126_;
  assign new_E2128_ = ~new_E2093_ & ~new_E2127_;
  assign new_E2129_ = new_E2093_ | new_E2126_;
  assign new_E2130_ = ~new_E2083_ & new_E2084_;
  assign new_E2131_ = new_E2083_ & ~new_E2084_;
  assign new_E2132_ = new_E2100_ | new_E2137_;
  assign new_E2133_ = ~new_E2100_ & ~new_E2136_;
  assign new_E2134_ = new_E2083_ | new_E2100_;
  assign new_E2135_ = new_E2083_ | new_E2084_;
  assign new_E2136_ = new_E2100_ & new_E2137_;
  assign new_E2137_ = ~new_E2082_ | ~new_E2107_;
  assign new_E2138_ = new_E2115_ & new_E2135_;
  assign new_E2139_ = ~new_E2115_ & ~new_E2135_;
  assign new_E2140_ = new_E2144_ | new_E2145_;
  assign new_E2141_ = ~new_E2086_ & new_E2100_;
  assign new_E2142_ = new_E2146_ | new_E2147_;
  assign new_E2143_ = new_E2086_ & new_E2100_;
  assign new_E2144_ = ~new_E2086_ & ~new_E2100_;
  assign new_E2145_ = new_E2086_ & ~new_E2100_;
  assign new_E2146_ = new_E2086_ & ~new_E2100_;
  assign new_E2147_ = ~new_E2086_ & new_E2100_;
  assign new_E2148_ = new_F3480_;
  assign new_E2149_ = new_F3547_;
  assign new_E2150_ = new_F3614_;
  assign new_E2151_ = new_F3681_;
  assign new_E2152_ = new_F3748_;
  assign new_E2153_ = new_F3815_;
  assign new_E2154_ = new_E2161_ & new_E2160_;
  assign new_E2155_ = new_E2163_ | new_E2162_;
  assign new_E2156_ = new_E2165_ | new_E2164_;
  assign new_E2157_ = new_E2167_ & new_E2166_;
  assign new_E2158_ = new_E2167_ & new_E2168_;
  assign new_E2159_ = new_E2160_ | new_E2169_;
  assign new_E2160_ = new_E2149_ | new_E2172_;
  assign new_E2161_ = new_E2171_ | new_E2170_;
  assign new_E2162_ = new_E2176_ & new_E2175_;
  assign new_E2163_ = new_E2174_ & new_E2173_;
  assign new_E2164_ = new_E2179_ | new_E2178_;
  assign new_E2165_ = new_E2174_ & new_E2177_;
  assign new_E2166_ = new_E2149_ | new_E2182_;
  assign new_E2167_ = new_E2181_ | new_E2180_;
  assign new_E2168_ = new_E2184_ | new_E2183_;
  assign new_E2169_ = ~new_E2160_ & new_E2186_;
  assign new_E2170_ = ~new_E2162_ & new_E2174_;
  assign new_E2171_ = new_E2162_ & ~new_E2174_;
  assign new_E2172_ = new_E2148_ & ~new_E2149_;
  assign new_E2173_ = ~new_E2195_ | ~new_E2196_;
  assign new_E2174_ = new_E2188_ | new_E2190_;
  assign new_E2175_ = new_E2198_ | new_E2197_;
  assign new_E2176_ = new_E2192_ | new_E2191_;
  assign new_E2177_ = ~new_E2200_ | ~new_E2199_;
  assign new_E2178_ = ~new_E2201_ & new_E2202_;
  assign new_E2179_ = new_E2201_ & ~new_E2202_;
  assign new_E2180_ = ~new_E2148_ & new_E2149_;
  assign new_E2181_ = new_E2148_ & ~new_E2149_;
  assign new_E2182_ = ~new_E2164_ | new_E2174_;
  assign new_E2183_ = new_E2164_ & new_E2174_;
  assign new_E2184_ = ~new_E2164_ & ~new_E2174_;
  assign new_E2185_ = new_E2206_ | new_E2205_;
  assign new_E2186_ = new_E2152_ | new_E2185_;
  assign new_E2187_ = new_E2210_ | new_E2209_;
  assign new_E2188_ = ~new_E2152_ & new_E2187_;
  assign new_E2189_ = new_E2208_ | new_E2207_;
  assign new_E2190_ = new_E2152_ & new_E2189_;
  assign new_E2191_ = new_E2150_ & ~new_E2160_;
  assign new_E2192_ = ~new_E2150_ & new_E2160_;
  assign new_E2193_ = ~new_E2149_ | ~new_E2174_;
  assign new_E2194_ = new_E2160_ & new_E2193_;
  assign new_E2195_ = ~new_E2160_ & ~new_E2194_;
  assign new_E2196_ = new_E2160_ | new_E2193_;
  assign new_E2197_ = ~new_E2150_ & new_E2151_;
  assign new_E2198_ = new_E2150_ & ~new_E2151_;
  assign new_E2199_ = new_E2167_ | new_E2204_;
  assign new_E2200_ = ~new_E2167_ & ~new_E2203_;
  assign new_E2201_ = new_E2150_ | new_E2167_;
  assign new_E2202_ = new_E2150_ | new_E2151_;
  assign new_E2203_ = new_E2167_ & new_E2204_;
  assign new_E2204_ = ~new_E2149_ | ~new_E2174_;
  assign new_E2205_ = new_E2182_ & new_E2202_;
  assign new_E2206_ = ~new_E2182_ & ~new_E2202_;
  assign new_E2207_ = new_E2211_ | new_E2212_;
  assign new_E2208_ = ~new_E2153_ & new_E2167_;
  assign new_E2209_ = new_E2213_ | new_E2214_;
  assign new_E2210_ = new_E2153_ & new_E2167_;
  assign new_E2211_ = ~new_E2153_ & ~new_E2167_;
  assign new_E2212_ = new_E2153_ & ~new_E2167_;
  assign new_E2213_ = new_E2153_ & ~new_E2167_;
  assign new_E2214_ = ~new_E2153_ & new_E2167_;
  assign new_E2215_ = new_F3882_;
  assign new_E2216_ = new_F3949_;
  assign new_E2217_ = new_F4016_;
  assign new_E2218_ = new_F4083_;
  assign new_E2219_ = new_F4150_;
  assign new_E2220_ = new_F4217_;
  assign new_E2221_ = new_E2228_ & new_E2227_;
  assign new_E2222_ = new_E2230_ | new_E2229_;
  assign new_E2223_ = new_E2232_ | new_E2231_;
  assign new_E2224_ = new_E2234_ & new_E2233_;
  assign new_E2225_ = new_E2234_ & new_E2235_;
  assign new_E2226_ = new_E2227_ | new_E2236_;
  assign new_E2227_ = new_E2216_ | new_E2239_;
  assign new_E2228_ = new_E2238_ | new_E2237_;
  assign new_E2229_ = new_E2243_ & new_E2242_;
  assign new_E2230_ = new_E2241_ & new_E2240_;
  assign new_E2231_ = new_E2246_ | new_E2245_;
  assign new_E2232_ = new_E2241_ & new_E2244_;
  assign new_E2233_ = new_E2216_ | new_E2249_;
  assign new_E2234_ = new_E2248_ | new_E2247_;
  assign new_E2235_ = new_E2251_ | new_E2250_;
  assign new_E2236_ = ~new_E2227_ & new_E2253_;
  assign new_E2237_ = ~new_E2229_ & new_E2241_;
  assign new_E2238_ = new_E2229_ & ~new_E2241_;
  assign new_E2239_ = new_E2215_ & ~new_E2216_;
  assign new_E2240_ = ~new_E2262_ | ~new_E2263_;
  assign new_E2241_ = new_E2255_ | new_E2257_;
  assign new_E2242_ = new_E2265_ | new_E2264_;
  assign new_E2243_ = new_E2259_ | new_E2258_;
  assign new_E2244_ = ~new_E2267_ | ~new_E2266_;
  assign new_E2245_ = ~new_E2268_ & new_E2269_;
  assign new_E2246_ = new_E2268_ & ~new_E2269_;
  assign new_E2247_ = ~new_E2215_ & new_E2216_;
  assign new_E2248_ = new_E2215_ & ~new_E2216_;
  assign new_E2249_ = ~new_E2231_ | new_E2241_;
  assign new_E2250_ = new_E2231_ & new_E2241_;
  assign new_E2251_ = ~new_E2231_ & ~new_E2241_;
  assign new_E2252_ = new_E2273_ | new_E2272_;
  assign new_E2253_ = new_E2219_ | new_E2252_;
  assign new_E2254_ = new_E2277_ | new_E2276_;
  assign new_E2255_ = ~new_E2219_ & new_E2254_;
  assign new_E2256_ = new_E2275_ | new_E2274_;
  assign new_E2257_ = new_E2219_ & new_E2256_;
  assign new_E2258_ = new_E2217_ & ~new_E2227_;
  assign new_E2259_ = ~new_E2217_ & new_E2227_;
  assign new_E2260_ = ~new_E2216_ | ~new_E2241_;
  assign new_E2261_ = new_E2227_ & new_E2260_;
  assign new_E2262_ = ~new_E2227_ & ~new_E2261_;
  assign new_E2263_ = new_E2227_ | new_E2260_;
  assign new_E2264_ = ~new_E2217_ & new_E2218_;
  assign new_E2265_ = new_E2217_ & ~new_E2218_;
  assign new_E2266_ = new_E2234_ | new_E2271_;
  assign new_E2267_ = ~new_E2234_ & ~new_E2270_;
  assign new_E2268_ = new_E2217_ | new_E2234_;
  assign new_E2269_ = new_E2217_ | new_E2218_;
  assign new_E2270_ = new_E2234_ & new_E2271_;
  assign new_E2271_ = ~new_E2216_ | ~new_E2241_;
  assign new_E2272_ = new_E2249_ & new_E2269_;
  assign new_E2273_ = ~new_E2249_ & ~new_E2269_;
  assign new_E2274_ = new_E2278_ | new_E2279_;
  assign new_E2275_ = ~new_E2220_ & new_E2234_;
  assign new_E2276_ = new_E2280_ | new_E2281_;
  assign new_E2277_ = new_E2220_ & new_E2234_;
  assign new_E2278_ = ~new_E2220_ & ~new_E2234_;
  assign new_E2279_ = new_E2220_ & ~new_E2234_;
  assign new_E2280_ = new_E2220_ & ~new_E2234_;
  assign new_E2281_ = ~new_E2220_ & new_E2234_;
  assign new_E2282_ = new_F4284_;
  assign new_E2283_ = new_F4351_;
  assign new_E2284_ = new_F4418_;
  assign new_E2285_ = new_F4485_;
  assign new_E2286_ = new_F4552_;
  assign new_E2287_ = new_F4619_;
  assign new_E2288_ = new_E2295_ & new_E2294_;
  assign new_E2289_ = new_E2297_ | new_E2296_;
  assign new_E2290_ = new_E2299_ | new_E2298_;
  assign new_E2291_ = new_E2301_ & new_E2300_;
  assign new_E2292_ = new_E2301_ & new_E2302_;
  assign new_E2293_ = new_E2294_ | new_E2303_;
  assign new_E2294_ = new_E2283_ | new_E2306_;
  assign new_E2295_ = new_E2305_ | new_E2304_;
  assign new_E2296_ = new_E2310_ & new_E2309_;
  assign new_E2297_ = new_E2308_ & new_E2307_;
  assign new_E2298_ = new_E2313_ | new_E2312_;
  assign new_E2299_ = new_E2308_ & new_E2311_;
  assign new_E2300_ = new_E2283_ | new_E2316_;
  assign new_E2301_ = new_E2315_ | new_E2314_;
  assign new_E2302_ = new_E2318_ | new_E2317_;
  assign new_E2303_ = ~new_E2294_ & new_E2320_;
  assign new_E2304_ = ~new_E2296_ & new_E2308_;
  assign new_E2305_ = new_E2296_ & ~new_E2308_;
  assign new_E2306_ = new_E2282_ & ~new_E2283_;
  assign new_E2307_ = ~new_E2329_ | ~new_E2330_;
  assign new_E2308_ = new_E2322_ | new_E2324_;
  assign new_E2309_ = new_E2332_ | new_E2331_;
  assign new_E2310_ = new_E2326_ | new_E2325_;
  assign new_E2311_ = ~new_E2334_ | ~new_E2333_;
  assign new_E2312_ = ~new_E2335_ & new_E2336_;
  assign new_E2313_ = new_E2335_ & ~new_E2336_;
  assign new_E2314_ = ~new_E2282_ & new_E2283_;
  assign new_E2315_ = new_E2282_ & ~new_E2283_;
  assign new_E2316_ = ~new_E2298_ | new_E2308_;
  assign new_E2317_ = new_E2298_ & new_E2308_;
  assign new_E2318_ = ~new_E2298_ & ~new_E2308_;
  assign new_E2319_ = new_E2340_ | new_E2339_;
  assign new_E2320_ = new_E2286_ | new_E2319_;
  assign new_E2321_ = new_E2344_ | new_E2343_;
  assign new_E2322_ = ~new_E2286_ & new_E2321_;
  assign new_E2323_ = new_E2342_ | new_E2341_;
  assign new_E2324_ = new_E2286_ & new_E2323_;
  assign new_E2325_ = new_E2284_ & ~new_E2294_;
  assign new_E2326_ = ~new_E2284_ & new_E2294_;
  assign new_E2327_ = ~new_E2283_ | ~new_E2308_;
  assign new_E2328_ = new_E2294_ & new_E2327_;
  assign new_E2329_ = ~new_E2294_ & ~new_E2328_;
  assign new_E2330_ = new_E2294_ | new_E2327_;
  assign new_E2331_ = ~new_E2284_ & new_E2285_;
  assign new_E2332_ = new_E2284_ & ~new_E2285_;
  assign new_E2333_ = new_E2301_ | new_E2338_;
  assign new_E2334_ = ~new_E2301_ & ~new_E2337_;
  assign new_E2335_ = new_E2284_ | new_E2301_;
  assign new_E2336_ = new_E2284_ | new_E2285_;
  assign new_E2337_ = new_E2301_ & new_E2338_;
  assign new_E2338_ = ~new_E2283_ | ~new_E2308_;
  assign new_E2339_ = new_E2316_ & new_E2336_;
  assign new_E2340_ = ~new_E2316_ & ~new_E2336_;
  assign new_E2341_ = new_E2345_ | new_E2346_;
  assign new_E2342_ = ~new_E2287_ & new_E2301_;
  assign new_E2343_ = new_E2347_ | new_E2348_;
  assign new_E2344_ = new_E2287_ & new_E2301_;
  assign new_E2345_ = ~new_E2287_ & ~new_E2301_;
  assign new_E2346_ = new_E2287_ & ~new_E2301_;
  assign new_E2347_ = new_E2287_ & ~new_E2301_;
  assign new_E2348_ = ~new_E2287_ & new_E2301_;
  assign new_E2349_ = new_F4686_;
  assign new_E2350_ = new_F4753_;
  assign new_E2351_ = new_F4820_;
  assign new_E2352_ = new_F4887_;
  assign new_E2353_ = new_F4954_;
  assign new_E2354_ = new_F5021_;
  assign new_E2355_ = new_E2362_ & new_E2361_;
  assign new_E2356_ = new_E2364_ | new_E2363_;
  assign new_E2357_ = new_E2366_ | new_E2365_;
  assign new_E2358_ = new_E2368_ & new_E2367_;
  assign new_E2359_ = new_E2368_ & new_E2369_;
  assign new_E2360_ = new_E2361_ | new_E2370_;
  assign new_E2361_ = new_E2350_ | new_E2373_;
  assign new_E2362_ = new_E2372_ | new_E2371_;
  assign new_E2363_ = new_E2377_ & new_E2376_;
  assign new_E2364_ = new_E2375_ & new_E2374_;
  assign new_E2365_ = new_E2380_ | new_E2379_;
  assign new_E2366_ = new_E2375_ & new_E2378_;
  assign new_E2367_ = new_E2350_ | new_E2383_;
  assign new_E2368_ = new_E2382_ | new_E2381_;
  assign new_E2369_ = new_E2385_ | new_E2384_;
  assign new_E2370_ = ~new_E2361_ & new_E2387_;
  assign new_E2371_ = ~new_E2363_ & new_E2375_;
  assign new_E2372_ = new_E2363_ & ~new_E2375_;
  assign new_E2373_ = new_E2349_ & ~new_E2350_;
  assign new_E2374_ = ~new_E2396_ | ~new_E2397_;
  assign new_E2375_ = new_E2389_ | new_E2391_;
  assign new_E2376_ = new_E2399_ | new_E2398_;
  assign new_E2377_ = new_E2393_ | new_E2392_;
  assign new_E2378_ = ~new_E2401_ | ~new_E2400_;
  assign new_E2379_ = ~new_E2402_ & new_E2403_;
  assign new_E2380_ = new_E2402_ & ~new_E2403_;
  assign new_E2381_ = ~new_E2349_ & new_E2350_;
  assign new_E2382_ = new_E2349_ & ~new_E2350_;
  assign new_E2383_ = ~new_E2365_ | new_E2375_;
  assign new_E2384_ = new_E2365_ & new_E2375_;
  assign new_E2385_ = ~new_E2365_ & ~new_E2375_;
  assign new_E2386_ = new_E2407_ | new_E2406_;
  assign new_E2387_ = new_E2353_ | new_E2386_;
  assign new_E2388_ = new_E2411_ | new_E2410_;
  assign new_E2389_ = ~new_E2353_ & new_E2388_;
  assign new_E2390_ = new_E2409_ | new_E2408_;
  assign new_E2391_ = new_E2353_ & new_E2390_;
  assign new_E2392_ = new_E2351_ & ~new_E2361_;
  assign new_E2393_ = ~new_E2351_ & new_E2361_;
  assign new_E2394_ = ~new_E2350_ | ~new_E2375_;
  assign new_E2395_ = new_E2361_ & new_E2394_;
  assign new_E2396_ = ~new_E2361_ & ~new_E2395_;
  assign new_E2397_ = new_E2361_ | new_E2394_;
  assign new_E2398_ = ~new_E2351_ & new_E2352_;
  assign new_E2399_ = new_E2351_ & ~new_E2352_;
  assign new_E2400_ = new_E2368_ | new_E2405_;
  assign new_E2401_ = ~new_E2368_ & ~new_E2404_;
  assign new_E2402_ = new_E2351_ | new_E2368_;
  assign new_E2403_ = new_E2351_ | new_E2352_;
  assign new_E2404_ = new_E2368_ & new_E2405_;
  assign new_E2405_ = ~new_E2350_ | ~new_E2375_;
  assign new_E2406_ = new_E2383_ & new_E2403_;
  assign new_E2407_ = ~new_E2383_ & ~new_E2403_;
  assign new_E2408_ = new_E2412_ | new_E2413_;
  assign new_E2409_ = ~new_E2354_ & new_E2368_;
  assign new_E2410_ = new_E2414_ | new_E2415_;
  assign new_E2411_ = new_E2354_ & new_E2368_;
  assign new_E2412_ = ~new_E2354_ & ~new_E2368_;
  assign new_E2413_ = new_E2354_ & ~new_E2368_;
  assign new_E2414_ = new_E2354_ & ~new_E2368_;
  assign new_E2415_ = ~new_E2354_ & new_E2368_;
  assign new_E2416_ = new_F5088_;
  assign new_E2417_ = new_F5155_;
  assign new_E2418_ = new_F5222_;
  assign new_E2419_ = new_F5289_;
  assign new_E2420_ = new_F5356_;
  assign new_E2421_ = new_F5423_;
  assign new_E2422_ = new_E2429_ & new_E2428_;
  assign new_E2423_ = new_E2431_ | new_E2430_;
  assign new_E2424_ = new_E2433_ | new_E2432_;
  assign new_E2425_ = new_E2435_ & new_E2434_;
  assign new_E2426_ = new_E2435_ & new_E2436_;
  assign new_E2427_ = new_E2428_ | new_E2437_;
  assign new_E2428_ = new_E2417_ | new_E2440_;
  assign new_E2429_ = new_E2439_ | new_E2438_;
  assign new_E2430_ = new_E2444_ & new_E2443_;
  assign new_E2431_ = new_E2442_ & new_E2441_;
  assign new_E2432_ = new_E2447_ | new_E2446_;
  assign new_E2433_ = new_E2442_ & new_E2445_;
  assign new_E2434_ = new_E2417_ | new_E2450_;
  assign new_E2435_ = new_E2449_ | new_E2448_;
  assign new_E2436_ = new_E2452_ | new_E2451_;
  assign new_E2437_ = ~new_E2428_ & new_E2454_;
  assign new_E2438_ = ~new_E2430_ & new_E2442_;
  assign new_E2439_ = new_E2430_ & ~new_E2442_;
  assign new_E2440_ = new_E2416_ & ~new_E2417_;
  assign new_E2441_ = ~new_E2463_ | ~new_E2464_;
  assign new_E2442_ = new_E2456_ | new_E2458_;
  assign new_E2443_ = new_E2466_ | new_E2465_;
  assign new_E2444_ = new_E2460_ | new_E2459_;
  assign new_E2445_ = ~new_E2468_ | ~new_E2467_;
  assign new_E2446_ = ~new_E2469_ & new_E2470_;
  assign new_E2447_ = new_E2469_ & ~new_E2470_;
  assign new_E2448_ = ~new_E2416_ & new_E2417_;
  assign new_E2449_ = new_E2416_ & ~new_E2417_;
  assign new_E2450_ = ~new_E2432_ | new_E2442_;
  assign new_E2451_ = new_E2432_ & new_E2442_;
  assign new_E2452_ = ~new_E2432_ & ~new_E2442_;
  assign new_E2453_ = new_E2474_ | new_E2473_;
  assign new_E2454_ = new_E2420_ | new_E2453_;
  assign new_E2455_ = new_E2478_ | new_E2477_;
  assign new_E2456_ = ~new_E2420_ & new_E2455_;
  assign new_E2457_ = new_E2476_ | new_E2475_;
  assign new_E2458_ = new_E2420_ & new_E2457_;
  assign new_E2459_ = new_E2418_ & ~new_E2428_;
  assign new_E2460_ = ~new_E2418_ & new_E2428_;
  assign new_E2461_ = ~new_E2417_ | ~new_E2442_;
  assign new_E2462_ = new_E2428_ & new_E2461_;
  assign new_E2463_ = ~new_E2428_ & ~new_E2462_;
  assign new_E2464_ = new_E2428_ | new_E2461_;
  assign new_E2465_ = ~new_E2418_ & new_E2419_;
  assign new_E2466_ = new_E2418_ & ~new_E2419_;
  assign new_E2467_ = new_E2435_ | new_E2472_;
  assign new_E2468_ = ~new_E2435_ & ~new_E2471_;
  assign new_E2469_ = new_E2418_ | new_E2435_;
  assign new_E2470_ = new_E2418_ | new_E2419_;
  assign new_E2471_ = new_E2435_ & new_E2472_;
  assign new_E2472_ = ~new_E2417_ | ~new_E2442_;
  assign new_E2473_ = new_E2450_ & new_E2470_;
  assign new_E2474_ = ~new_E2450_ & ~new_E2470_;
  assign new_E2475_ = new_E2479_ | new_E2480_;
  assign new_E2476_ = ~new_E2421_ & new_E2435_;
  assign new_E2477_ = new_E2481_ | new_E2482_;
  assign new_E2478_ = new_E2421_ & new_E2435_;
  assign new_E2479_ = ~new_E2421_ & ~new_E2435_;
  assign new_E2480_ = new_E2421_ & ~new_E2435_;
  assign new_E2481_ = new_E2421_ & ~new_E2435_;
  assign new_E2482_ = ~new_E2421_ & new_E2435_;
  assign new_E2483_ = new_F5490_;
  assign new_E2484_ = new_F5557_;
  assign new_E2485_ = new_F5624_;
  assign new_E2486_ = new_F5691_;
  assign new_E2487_ = new_F5758_;
  assign new_E2488_ = new_F5825_;
  assign new_E2489_ = new_E2496_ & new_E2495_;
  assign new_E2490_ = new_E2498_ | new_E2497_;
  assign new_E2491_ = new_E2500_ | new_E2499_;
  assign new_E2492_ = new_E2502_ & new_E2501_;
  assign new_E2493_ = new_E2502_ & new_E2503_;
  assign new_E2494_ = new_E2495_ | new_E2504_;
  assign new_E2495_ = new_E2484_ | new_E2507_;
  assign new_E2496_ = new_E2506_ | new_E2505_;
  assign new_E2497_ = new_E2511_ & new_E2510_;
  assign new_E2498_ = new_E2509_ & new_E2508_;
  assign new_E2499_ = new_E2514_ | new_E2513_;
  assign new_E2500_ = new_E2509_ & new_E2512_;
  assign new_E2501_ = new_E2484_ | new_E2517_;
  assign new_E2502_ = new_E2516_ | new_E2515_;
  assign new_E2503_ = new_E2519_ | new_E2518_;
  assign new_E2504_ = ~new_E2495_ & new_E2521_;
  assign new_E2505_ = ~new_E2497_ & new_E2509_;
  assign new_E2506_ = new_E2497_ & ~new_E2509_;
  assign new_E2507_ = new_E2483_ & ~new_E2484_;
  assign new_E2508_ = ~new_E2530_ | ~new_E2531_;
  assign new_E2509_ = new_E2523_ | new_E2525_;
  assign new_E2510_ = new_E2533_ | new_E2532_;
  assign new_E2511_ = new_E2527_ | new_E2526_;
  assign new_E2512_ = ~new_E2535_ | ~new_E2534_;
  assign new_E2513_ = ~new_E2536_ & new_E2537_;
  assign new_E2514_ = new_E2536_ & ~new_E2537_;
  assign new_E2515_ = ~new_E2483_ & new_E2484_;
  assign new_E2516_ = new_E2483_ & ~new_E2484_;
  assign new_E2517_ = ~new_E2499_ | new_E2509_;
  assign new_E2518_ = new_E2499_ & new_E2509_;
  assign new_E2519_ = ~new_E2499_ & ~new_E2509_;
  assign new_E2520_ = new_E2541_ | new_E2540_;
  assign new_E2521_ = new_E2487_ | new_E2520_;
  assign new_E2522_ = new_E2545_ | new_E2544_;
  assign new_E2523_ = ~new_E2487_ & new_E2522_;
  assign new_E2524_ = new_E2543_ | new_E2542_;
  assign new_E2525_ = new_E2487_ & new_E2524_;
  assign new_E2526_ = new_E2485_ & ~new_E2495_;
  assign new_E2527_ = ~new_E2485_ & new_E2495_;
  assign new_E2528_ = ~new_E2484_ | ~new_E2509_;
  assign new_E2529_ = new_E2495_ & new_E2528_;
  assign new_E2530_ = ~new_E2495_ & ~new_E2529_;
  assign new_E2531_ = new_E2495_ | new_E2528_;
  assign new_E2532_ = ~new_E2485_ & new_E2486_;
  assign new_E2533_ = new_E2485_ & ~new_E2486_;
  assign new_E2534_ = new_E2502_ | new_E2539_;
  assign new_E2535_ = ~new_E2502_ & ~new_E2538_;
  assign new_E2536_ = new_E2485_ | new_E2502_;
  assign new_E2537_ = new_E2485_ | new_E2486_;
  assign new_E2538_ = new_E2502_ & new_E2539_;
  assign new_E2539_ = ~new_E2484_ | ~new_E2509_;
  assign new_E2540_ = new_E2517_ & new_E2537_;
  assign new_E2541_ = ~new_E2517_ & ~new_E2537_;
  assign new_E2542_ = new_E2546_ | new_E2547_;
  assign new_E2543_ = ~new_E2488_ & new_E2502_;
  assign new_E2544_ = new_E2548_ | new_E2549_;
  assign new_E2545_ = new_E2488_ & new_E2502_;
  assign new_E2546_ = ~new_E2488_ & ~new_E2502_;
  assign new_E2547_ = new_E2488_ & ~new_E2502_;
  assign new_E2548_ = new_E2488_ & ~new_E2502_;
  assign new_E2549_ = ~new_E2488_ & new_E2502_;
  assign new_E2550_ = new_F5892_;
  assign new_E2551_ = new_F5959_;
  assign new_E2552_ = new_F6026_;
  assign new_E2553_ = new_F6093_;
  assign new_E2554_ = new_F6160_;
  assign new_E2555_ = new_F6227_;
  assign new_E2556_ = new_E2563_ & new_E2562_;
  assign new_E2557_ = new_E2565_ | new_E2564_;
  assign new_E2558_ = new_E2567_ | new_E2566_;
  assign new_E2559_ = new_E2569_ & new_E2568_;
  assign new_E2560_ = new_E2569_ & new_E2570_;
  assign new_E2561_ = new_E2562_ | new_E2571_;
  assign new_E2562_ = new_E2551_ | new_E2574_;
  assign new_E2563_ = new_E2573_ | new_E2572_;
  assign new_E2564_ = new_E2578_ & new_E2577_;
  assign new_E2565_ = new_E2576_ & new_E2575_;
  assign new_E2566_ = new_E2581_ | new_E2580_;
  assign new_E2567_ = new_E2576_ & new_E2579_;
  assign new_E2568_ = new_E2551_ | new_E2584_;
  assign new_E2569_ = new_E2583_ | new_E2582_;
  assign new_E2570_ = new_E2586_ | new_E2585_;
  assign new_E2571_ = ~new_E2562_ & new_E2588_;
  assign new_E2572_ = ~new_E2564_ & new_E2576_;
  assign new_E2573_ = new_E2564_ & ~new_E2576_;
  assign new_E2574_ = new_E2550_ & ~new_E2551_;
  assign new_E2575_ = ~new_E2597_ | ~new_E2598_;
  assign new_E2576_ = new_E2590_ | new_E2592_;
  assign new_E2577_ = new_E2600_ | new_E2599_;
  assign new_E2578_ = new_E2594_ | new_E2593_;
  assign new_E2579_ = ~new_E2602_ | ~new_E2601_;
  assign new_E2580_ = ~new_E2603_ & new_E2604_;
  assign new_E2581_ = new_E2603_ & ~new_E2604_;
  assign new_E2582_ = ~new_E2550_ & new_E2551_;
  assign new_E2583_ = new_E2550_ & ~new_E2551_;
  assign new_E2584_ = ~new_E2566_ | new_E2576_;
  assign new_E2585_ = new_E2566_ & new_E2576_;
  assign new_E2586_ = ~new_E2566_ & ~new_E2576_;
  assign new_E2587_ = new_E2608_ | new_E2607_;
  assign new_E2588_ = new_E2554_ | new_E2587_;
  assign new_E2589_ = new_E2612_ | new_E2611_;
  assign new_E2590_ = ~new_E2554_ & new_E2589_;
  assign new_E2591_ = new_E2610_ | new_E2609_;
  assign new_E2592_ = new_E2554_ & new_E2591_;
  assign new_E2593_ = new_E2552_ & ~new_E2562_;
  assign new_E2594_ = ~new_E2552_ & new_E2562_;
  assign new_E2595_ = ~new_E2551_ | ~new_E2576_;
  assign new_E2596_ = new_E2562_ & new_E2595_;
  assign new_E2597_ = ~new_E2562_ & ~new_E2596_;
  assign new_E2598_ = new_E2562_ | new_E2595_;
  assign new_E2599_ = ~new_E2552_ & new_E2553_;
  assign new_E2600_ = new_E2552_ & ~new_E2553_;
  assign new_E2601_ = new_E2569_ | new_E2606_;
  assign new_E2602_ = ~new_E2569_ & ~new_E2605_;
  assign new_E2603_ = new_E2552_ | new_E2569_;
  assign new_E2604_ = new_E2552_ | new_E2553_;
  assign new_E2605_ = new_E2569_ & new_E2606_;
  assign new_E2606_ = ~new_E2551_ | ~new_E2576_;
  assign new_E2607_ = new_E2584_ & new_E2604_;
  assign new_E2608_ = ~new_E2584_ & ~new_E2604_;
  assign new_E2609_ = new_E2613_ | new_E2614_;
  assign new_E2610_ = ~new_E2555_ & new_E2569_;
  assign new_E2611_ = new_E2615_ | new_E2616_;
  assign new_E2612_ = new_E2555_ & new_E2569_;
  assign new_E2613_ = ~new_E2555_ & ~new_E2569_;
  assign new_E2614_ = new_E2555_ & ~new_E2569_;
  assign new_E2615_ = new_E2555_ & ~new_E2569_;
  assign new_E2616_ = ~new_E2555_ & new_E2569_;
  assign new_E2617_ = new_F6294_;
  assign new_E2618_ = new_F6361_;
  assign new_E2619_ = new_F6428_;
  assign new_E2620_ = new_F6495_;
  assign new_E2621_ = new_F6562_;
  assign new_E2622_ = new_F6629_;
  assign new_E2623_ = new_E2630_ & new_E2629_;
  assign new_E2624_ = new_E2632_ | new_E2631_;
  assign new_E2625_ = new_E2634_ | new_E2633_;
  assign new_E2626_ = new_E2636_ & new_E2635_;
  assign new_E2627_ = new_E2636_ & new_E2637_;
  assign new_E2628_ = new_E2629_ | new_E2638_;
  assign new_E2629_ = new_E2618_ | new_E2641_;
  assign new_E2630_ = new_E2640_ | new_E2639_;
  assign new_E2631_ = new_E2645_ & new_E2644_;
  assign new_E2632_ = new_E2643_ & new_E2642_;
  assign new_E2633_ = new_E2648_ | new_E2647_;
  assign new_E2634_ = new_E2643_ & new_E2646_;
  assign new_E2635_ = new_E2618_ | new_E2651_;
  assign new_E2636_ = new_E2650_ | new_E2649_;
  assign new_E2637_ = new_E2653_ | new_E2652_;
  assign new_E2638_ = ~new_E2629_ & new_E2655_;
  assign new_E2639_ = ~new_E2631_ & new_E2643_;
  assign new_E2640_ = new_E2631_ & ~new_E2643_;
  assign new_E2641_ = new_E2617_ & ~new_E2618_;
  assign new_E2642_ = ~new_E2664_ | ~new_E2665_;
  assign new_E2643_ = new_E2657_ | new_E2659_;
  assign new_E2644_ = new_E2667_ | new_E2666_;
  assign new_E2645_ = new_E2661_ | new_E2660_;
  assign new_E2646_ = ~new_E2669_ | ~new_E2668_;
  assign new_E2647_ = ~new_E2670_ & new_E2671_;
  assign new_E2648_ = new_E2670_ & ~new_E2671_;
  assign new_E2649_ = ~new_E2617_ & new_E2618_;
  assign new_E2650_ = new_E2617_ & ~new_E2618_;
  assign new_E2651_ = ~new_E2633_ | new_E2643_;
  assign new_E2652_ = new_E2633_ & new_E2643_;
  assign new_E2653_ = ~new_E2633_ & ~new_E2643_;
  assign new_E2654_ = new_E2675_ | new_E2674_;
  assign new_E2655_ = new_E2621_ | new_E2654_;
  assign new_E2656_ = new_E2679_ | new_E2678_;
  assign new_E2657_ = ~new_E2621_ & new_E2656_;
  assign new_E2658_ = new_E2677_ | new_E2676_;
  assign new_E2659_ = new_E2621_ & new_E2658_;
  assign new_E2660_ = new_E2619_ & ~new_E2629_;
  assign new_E2661_ = ~new_E2619_ & new_E2629_;
  assign new_E2662_ = ~new_E2618_ | ~new_E2643_;
  assign new_E2663_ = new_E2629_ & new_E2662_;
  assign new_E2664_ = ~new_E2629_ & ~new_E2663_;
  assign new_E2665_ = new_E2629_ | new_E2662_;
  assign new_E2666_ = ~new_E2619_ & new_E2620_;
  assign new_E2667_ = new_E2619_ & ~new_E2620_;
  assign new_E2668_ = new_E2636_ | new_E2673_;
  assign new_E2669_ = ~new_E2636_ & ~new_E2672_;
  assign new_E2670_ = new_E2619_ | new_E2636_;
  assign new_E2671_ = new_E2619_ | new_E2620_;
  assign new_E2672_ = new_E2636_ & new_E2673_;
  assign new_E2673_ = ~new_E2618_ | ~new_E2643_;
  assign new_E2674_ = new_E2651_ & new_E2671_;
  assign new_E2675_ = ~new_E2651_ & ~new_E2671_;
  assign new_E2676_ = new_E2680_ | new_E2681_;
  assign new_E2677_ = ~new_E2622_ & new_E2636_;
  assign new_E2678_ = new_E2682_ | new_E2683_;
  assign new_E2679_ = new_E2622_ & new_E2636_;
  assign new_E2680_ = ~new_E2622_ & ~new_E2636_;
  assign new_E2681_ = new_E2622_ & ~new_E2636_;
  assign new_E2682_ = new_E2622_ & ~new_E2636_;
  assign new_E2683_ = ~new_E2622_ & new_E2636_;
  assign new_E2684_ = new_F6696_;
  assign new_E2685_ = new_F6763_;
  assign new_E2686_ = new_F6830_;
  assign new_E2687_ = new_F6897_;
  assign new_E2688_ = new_F6964_;
  assign new_E2689_ = new_F7031_;
  assign new_E2690_ = new_E2697_ & new_E2696_;
  assign new_E2691_ = new_E2699_ | new_E2698_;
  assign new_E2692_ = new_E2701_ | new_E2700_;
  assign new_E2693_ = new_E2703_ & new_E2702_;
  assign new_E2694_ = new_E2703_ & new_E2704_;
  assign new_E2695_ = new_E2696_ | new_E2705_;
  assign new_E2696_ = new_E2685_ | new_E2708_;
  assign new_E2697_ = new_E2707_ | new_E2706_;
  assign new_E2698_ = new_E2712_ & new_E2711_;
  assign new_E2699_ = new_E2710_ & new_E2709_;
  assign new_E2700_ = new_E2715_ | new_E2714_;
  assign new_E2701_ = new_E2710_ & new_E2713_;
  assign new_E2702_ = new_E2685_ | new_E2718_;
  assign new_E2703_ = new_E2717_ | new_E2716_;
  assign new_E2704_ = new_E2720_ | new_E2719_;
  assign new_E2705_ = ~new_E2696_ & new_E2722_;
  assign new_E2706_ = ~new_E2698_ & new_E2710_;
  assign new_E2707_ = new_E2698_ & ~new_E2710_;
  assign new_E2708_ = new_E2684_ & ~new_E2685_;
  assign new_E2709_ = ~new_E2731_ | ~new_E2732_;
  assign new_E2710_ = new_E2724_ | new_E2726_;
  assign new_E2711_ = new_E2734_ | new_E2733_;
  assign new_E2712_ = new_E2728_ | new_E2727_;
  assign new_E2713_ = ~new_E2736_ | ~new_E2735_;
  assign new_E2714_ = ~new_E2737_ & new_E2738_;
  assign new_E2715_ = new_E2737_ & ~new_E2738_;
  assign new_E2716_ = ~new_E2684_ & new_E2685_;
  assign new_E2717_ = new_E2684_ & ~new_E2685_;
  assign new_E2718_ = ~new_E2700_ | new_E2710_;
  assign new_E2719_ = new_E2700_ & new_E2710_;
  assign new_E2720_ = ~new_E2700_ & ~new_E2710_;
  assign new_E2721_ = new_E2742_ | new_E2741_;
  assign new_E2722_ = new_E2688_ | new_E2721_;
  assign new_E2723_ = new_E2746_ | new_E2745_;
  assign new_E2724_ = ~new_E2688_ & new_E2723_;
  assign new_E2725_ = new_E2744_ | new_E2743_;
  assign new_E2726_ = new_E2688_ & new_E2725_;
  assign new_E2727_ = new_E2686_ & ~new_E2696_;
  assign new_E2728_ = ~new_E2686_ & new_E2696_;
  assign new_E2729_ = ~new_E2685_ | ~new_E2710_;
  assign new_E2730_ = new_E2696_ & new_E2729_;
  assign new_E2731_ = ~new_E2696_ & ~new_E2730_;
  assign new_E2732_ = new_E2696_ | new_E2729_;
  assign new_E2733_ = ~new_E2686_ & new_E2687_;
  assign new_E2734_ = new_E2686_ & ~new_E2687_;
  assign new_E2735_ = new_E2703_ | new_E2740_;
  assign new_E2736_ = ~new_E2703_ & ~new_E2739_;
  assign new_E2737_ = new_E2686_ | new_E2703_;
  assign new_E2738_ = new_E2686_ | new_E2687_;
  assign new_E2739_ = new_E2703_ & new_E2740_;
  assign new_E2740_ = ~new_E2685_ | ~new_E2710_;
  assign new_E2741_ = new_E2718_ & new_E2738_;
  assign new_E2742_ = ~new_E2718_ & ~new_E2738_;
  assign new_E2743_ = new_E2747_ | new_E2748_;
  assign new_E2744_ = ~new_E2689_ & new_E2703_;
  assign new_E2745_ = new_E2749_ | new_E2750_;
  assign new_E2746_ = new_E2689_ & new_E2703_;
  assign new_E2747_ = ~new_E2689_ & ~new_E2703_;
  assign new_E2748_ = new_E2689_ & ~new_E2703_;
  assign new_E2749_ = new_E2689_ & ~new_E2703_;
  assign new_E2750_ = ~new_E2689_ & new_E2703_;
  assign new_E2751_ = new_F7098_;
  assign new_E2752_ = new_F7165_;
  assign new_E2753_ = new_F7232_;
  assign new_E2754_ = new_F7299_;
  assign new_E2755_ = new_F7366_;
  assign new_E2756_ = new_F7433_;
  assign new_E2757_ = new_E2764_ & new_E2763_;
  assign new_E2758_ = new_E2766_ | new_E2765_;
  assign new_E2759_ = new_E2768_ | new_E2767_;
  assign new_E2760_ = new_E2770_ & new_E2769_;
  assign new_E2761_ = new_E2770_ & new_E2771_;
  assign new_E2762_ = new_E2763_ | new_E2772_;
  assign new_E2763_ = new_E2752_ | new_E2775_;
  assign new_E2764_ = new_E2774_ | new_E2773_;
  assign new_E2765_ = new_E2779_ & new_E2778_;
  assign new_E2766_ = new_E2777_ & new_E2776_;
  assign new_E2767_ = new_E2782_ | new_E2781_;
  assign new_E2768_ = new_E2777_ & new_E2780_;
  assign new_E2769_ = new_E2752_ | new_E2785_;
  assign new_E2770_ = new_E2784_ | new_E2783_;
  assign new_E2771_ = new_E2787_ | new_E2786_;
  assign new_E2772_ = ~new_E2763_ & new_E2789_;
  assign new_E2773_ = ~new_E2765_ & new_E2777_;
  assign new_E2774_ = new_E2765_ & ~new_E2777_;
  assign new_E2775_ = new_E2751_ & ~new_E2752_;
  assign new_E2776_ = ~new_E2798_ | ~new_E2799_;
  assign new_E2777_ = new_E2791_ | new_E2793_;
  assign new_E2778_ = new_E2801_ | new_E2800_;
  assign new_E2779_ = new_E2795_ | new_E2794_;
  assign new_E2780_ = ~new_E2803_ | ~new_E2802_;
  assign new_E2781_ = ~new_E2804_ & new_E2805_;
  assign new_E2782_ = new_E2804_ & ~new_E2805_;
  assign new_E2783_ = ~new_E2751_ & new_E2752_;
  assign new_E2784_ = new_E2751_ & ~new_E2752_;
  assign new_E2785_ = ~new_E2767_ | new_E2777_;
  assign new_E2786_ = new_E2767_ & new_E2777_;
  assign new_E2787_ = ~new_E2767_ & ~new_E2777_;
  assign new_E2788_ = new_E2809_ | new_E2808_;
  assign new_E2789_ = new_E2755_ | new_E2788_;
  assign new_E2790_ = new_E2813_ | new_E2812_;
  assign new_E2791_ = ~new_E2755_ & new_E2790_;
  assign new_E2792_ = new_E2811_ | new_E2810_;
  assign new_E2793_ = new_E2755_ & new_E2792_;
  assign new_E2794_ = new_E2753_ & ~new_E2763_;
  assign new_E2795_ = ~new_E2753_ & new_E2763_;
  assign new_E2796_ = ~new_E2752_ | ~new_E2777_;
  assign new_E2797_ = new_E2763_ & new_E2796_;
  assign new_E2798_ = ~new_E2763_ & ~new_E2797_;
  assign new_E2799_ = new_E2763_ | new_E2796_;
  assign new_E2800_ = ~new_E2753_ & new_E2754_;
  assign new_E2801_ = new_E2753_ & ~new_E2754_;
  assign new_E2802_ = new_E2770_ | new_E2807_;
  assign new_E2803_ = ~new_E2770_ & ~new_E2806_;
  assign new_E2804_ = new_E2753_ | new_E2770_;
  assign new_E2805_ = new_E2753_ | new_E2754_;
  assign new_E2806_ = new_E2770_ & new_E2807_;
  assign new_E2807_ = ~new_E2752_ | ~new_E2777_;
  assign new_E2808_ = new_E2785_ & new_E2805_;
  assign new_E2809_ = ~new_E2785_ & ~new_E2805_;
  assign new_E2810_ = new_E2814_ | new_E2815_;
  assign new_E2811_ = ~new_E2756_ & new_E2770_;
  assign new_E2812_ = new_E2816_ | new_E2817_;
  assign new_E2813_ = new_E2756_ & new_E2770_;
  assign new_E2814_ = ~new_E2756_ & ~new_E2770_;
  assign new_E2815_ = new_E2756_ & ~new_E2770_;
  assign new_E2816_ = new_E2756_ & ~new_E2770_;
  assign new_E2817_ = ~new_E2756_ & new_E2770_;
  assign new_E2818_ = new_F7500_;
  assign new_E2819_ = new_F7567_;
  assign new_E2820_ = new_F7634_;
  assign new_E2821_ = new_F7701_;
  assign new_E2822_ = new_F7768_;
  assign new_E2823_ = new_F7835_;
  assign new_E2824_ = new_E2831_ & new_E2830_;
  assign new_E2825_ = new_E2833_ | new_E2832_;
  assign new_E2826_ = new_E2835_ | new_E2834_;
  assign new_E2827_ = new_E2837_ & new_E2836_;
  assign new_E2828_ = new_E2837_ & new_E2838_;
  assign new_E2829_ = new_E2830_ | new_E2839_;
  assign new_E2830_ = new_E2819_ | new_E2842_;
  assign new_E2831_ = new_E2841_ | new_E2840_;
  assign new_E2832_ = new_E2846_ & new_E2845_;
  assign new_E2833_ = new_E2844_ & new_E2843_;
  assign new_E2834_ = new_E2849_ | new_E2848_;
  assign new_E2835_ = new_E2844_ & new_E2847_;
  assign new_E2836_ = new_E2819_ | new_E2852_;
  assign new_E2837_ = new_E2851_ | new_E2850_;
  assign new_E2838_ = new_E2854_ | new_E2853_;
  assign new_E2839_ = ~new_E2830_ & new_E2856_;
  assign new_E2840_ = ~new_E2832_ & new_E2844_;
  assign new_E2841_ = new_E2832_ & ~new_E2844_;
  assign new_E2842_ = new_E2818_ & ~new_E2819_;
  assign new_E2843_ = ~new_E2865_ | ~new_E2866_;
  assign new_E2844_ = new_E2858_ | new_E2860_;
  assign new_E2845_ = new_E2868_ | new_E2867_;
  assign new_E2846_ = new_E2862_ | new_E2861_;
  assign new_E2847_ = ~new_E2870_ | ~new_E2869_;
  assign new_E2848_ = ~new_E2871_ & new_E2872_;
  assign new_E2849_ = new_E2871_ & ~new_E2872_;
  assign new_E2850_ = ~new_E2818_ & new_E2819_;
  assign new_E2851_ = new_E2818_ & ~new_E2819_;
  assign new_E2852_ = ~new_E2834_ | new_E2844_;
  assign new_E2853_ = new_E2834_ & new_E2844_;
  assign new_E2854_ = ~new_E2834_ & ~new_E2844_;
  assign new_E2855_ = new_E2876_ | new_E2875_;
  assign new_E2856_ = new_E2822_ | new_E2855_;
  assign new_E2857_ = new_E2880_ | new_E2879_;
  assign new_E2858_ = ~new_E2822_ & new_E2857_;
  assign new_E2859_ = new_E2878_ | new_E2877_;
  assign new_E2860_ = new_E2822_ & new_E2859_;
  assign new_E2861_ = new_E2820_ & ~new_E2830_;
  assign new_E2862_ = ~new_E2820_ & new_E2830_;
  assign new_E2863_ = ~new_E2819_ | ~new_E2844_;
  assign new_E2864_ = new_E2830_ & new_E2863_;
  assign new_E2865_ = ~new_E2830_ & ~new_E2864_;
  assign new_E2866_ = new_E2830_ | new_E2863_;
  assign new_E2867_ = ~new_E2820_ & new_E2821_;
  assign new_E2868_ = new_E2820_ & ~new_E2821_;
  assign new_E2869_ = new_E2837_ | new_E2874_;
  assign new_E2870_ = ~new_E2837_ & ~new_E2873_;
  assign new_E2871_ = new_E2820_ | new_E2837_;
  assign new_E2872_ = new_E2820_ | new_E2821_;
  assign new_E2873_ = new_E2837_ & new_E2874_;
  assign new_E2874_ = ~new_E2819_ | ~new_E2844_;
  assign new_E2875_ = new_E2852_ & new_E2872_;
  assign new_E2876_ = ~new_E2852_ & ~new_E2872_;
  assign new_E2877_ = new_E2881_ | new_E2882_;
  assign new_E2878_ = ~new_E2823_ & new_E2837_;
  assign new_E2879_ = new_E2883_ | new_E2884_;
  assign new_E2880_ = new_E2823_ & new_E2837_;
  assign new_E2881_ = ~new_E2823_ & ~new_E2837_;
  assign new_E2882_ = new_E2823_ & ~new_E2837_;
  assign new_E2883_ = new_E2823_ & ~new_E2837_;
  assign new_E2884_ = ~new_E2823_ & new_E2837_;
  assign new_E2885_ = new_F7902_;
  assign new_E2886_ = new_F7969_;
  assign new_E2887_ = new_F8036_;
  assign new_E2888_ = new_F8103_;
  assign new_E2889_ = new_F8170_;
  assign new_E2890_ = new_F8237_;
  assign new_E2891_ = new_E2898_ & new_E2897_;
  assign new_E2892_ = new_E2900_ | new_E2899_;
  assign new_E2893_ = new_E2902_ | new_E2901_;
  assign new_E2894_ = new_E2904_ & new_E2903_;
  assign new_E2895_ = new_E2904_ & new_E2905_;
  assign new_E2896_ = new_E2897_ | new_E2906_;
  assign new_E2897_ = new_E2886_ | new_E2909_;
  assign new_E2898_ = new_E2908_ | new_E2907_;
  assign new_E2899_ = new_E2913_ & new_E2912_;
  assign new_E2900_ = new_E2911_ & new_E2910_;
  assign new_E2901_ = new_E2916_ | new_E2915_;
  assign new_E2902_ = new_E2911_ & new_E2914_;
  assign new_E2903_ = new_E2886_ | new_E2919_;
  assign new_E2904_ = new_E2918_ | new_E2917_;
  assign new_E2905_ = new_E2921_ | new_E2920_;
  assign new_E2906_ = ~new_E2897_ & new_E2923_;
  assign new_E2907_ = ~new_E2899_ & new_E2911_;
  assign new_E2908_ = new_E2899_ & ~new_E2911_;
  assign new_E2909_ = new_E2885_ & ~new_E2886_;
  assign new_E2910_ = ~new_E2932_ | ~new_E2933_;
  assign new_E2911_ = new_E2925_ | new_E2927_;
  assign new_E2912_ = new_E2935_ | new_E2934_;
  assign new_E2913_ = new_E2929_ | new_E2928_;
  assign new_E2914_ = ~new_E2937_ | ~new_E2936_;
  assign new_E2915_ = ~new_E2938_ & new_E2939_;
  assign new_E2916_ = new_E2938_ & ~new_E2939_;
  assign new_E2917_ = ~new_E2885_ & new_E2886_;
  assign new_E2918_ = new_E2885_ & ~new_E2886_;
  assign new_E2919_ = ~new_E2901_ | new_E2911_;
  assign new_E2920_ = new_E2901_ & new_E2911_;
  assign new_E2921_ = ~new_E2901_ & ~new_E2911_;
  assign new_E2922_ = new_E2943_ | new_E2942_;
  assign new_E2923_ = new_E2889_ | new_E2922_;
  assign new_E2924_ = new_E2947_ | new_E2946_;
  assign new_E2925_ = ~new_E2889_ & new_E2924_;
  assign new_E2926_ = new_E2945_ | new_E2944_;
  assign new_E2927_ = new_E2889_ & new_E2926_;
  assign new_E2928_ = new_E2887_ & ~new_E2897_;
  assign new_E2929_ = ~new_E2887_ & new_E2897_;
  assign new_E2930_ = ~new_E2886_ | ~new_E2911_;
  assign new_E2931_ = new_E2897_ & new_E2930_;
  assign new_E2932_ = ~new_E2897_ & ~new_E2931_;
  assign new_E2933_ = new_E2897_ | new_E2930_;
  assign new_E2934_ = ~new_E2887_ & new_E2888_;
  assign new_E2935_ = new_E2887_ & ~new_E2888_;
  assign new_E2936_ = new_E2904_ | new_E2941_;
  assign new_E2937_ = ~new_E2904_ & ~new_E2940_;
  assign new_E2938_ = new_E2887_ | new_E2904_;
  assign new_E2939_ = new_E2887_ | new_E2888_;
  assign new_E2940_ = new_E2904_ & new_E2941_;
  assign new_E2941_ = ~new_E2886_ | ~new_E2911_;
  assign new_E2942_ = new_E2919_ & new_E2939_;
  assign new_E2943_ = ~new_E2919_ & ~new_E2939_;
  assign new_E2944_ = new_E2948_ | new_E2949_;
  assign new_E2945_ = ~new_E2890_ & new_E2904_;
  assign new_E2946_ = new_E2950_ | new_E2951_;
  assign new_E2947_ = new_E2890_ & new_E2904_;
  assign new_E2948_ = ~new_E2890_ & ~new_E2904_;
  assign new_E2949_ = new_E2890_ & ~new_E2904_;
  assign new_E2950_ = new_E2890_ & ~new_E2904_;
  assign new_E2951_ = ~new_E2890_ & new_E2904_;
  assign new_E2952_ = new_F8304_;
  assign new_E2953_ = new_F8371_;
  assign new_E2954_ = new_F8438_;
  assign new_E2955_ = new_F8505_;
  assign new_E2956_ = new_F8572_;
  assign new_E2957_ = new_F8639_;
  assign new_E2958_ = new_E2965_ & new_E2964_;
  assign new_E2959_ = new_E2967_ | new_E2966_;
  assign new_E2960_ = new_E2969_ | new_E2968_;
  assign new_E2961_ = new_E2971_ & new_E2970_;
  assign new_E2962_ = new_E2971_ & new_E2972_;
  assign new_E2963_ = new_E2964_ | new_E2973_;
  assign new_E2964_ = new_E2953_ | new_E2976_;
  assign new_E2965_ = new_E2975_ | new_E2974_;
  assign new_E2966_ = new_E2980_ & new_E2979_;
  assign new_E2967_ = new_E2978_ & new_E2977_;
  assign new_E2968_ = new_E2983_ | new_E2982_;
  assign new_E2969_ = new_E2978_ & new_E2981_;
  assign new_E2970_ = new_E2953_ | new_E2986_;
  assign new_E2971_ = new_E2985_ | new_E2984_;
  assign new_E2972_ = new_E2988_ | new_E2987_;
  assign new_E2973_ = ~new_E2964_ & new_E2990_;
  assign new_E2974_ = ~new_E2966_ & new_E2978_;
  assign new_E2975_ = new_E2966_ & ~new_E2978_;
  assign new_E2976_ = new_E2952_ & ~new_E2953_;
  assign new_E2977_ = ~new_E2999_ | ~new_E3000_;
  assign new_E2978_ = new_E2992_ | new_E2994_;
  assign new_E2979_ = new_E3002_ | new_E3001_;
  assign new_E2980_ = new_E2996_ | new_E2995_;
  assign new_E2981_ = ~new_E3004_ | ~new_E3003_;
  assign new_E2982_ = ~new_E3005_ & new_E3006_;
  assign new_E2983_ = new_E3005_ & ~new_E3006_;
  assign new_E2984_ = ~new_E2952_ & new_E2953_;
  assign new_E2985_ = new_E2952_ & ~new_E2953_;
  assign new_E2986_ = ~new_E2968_ | new_E2978_;
  assign new_E2987_ = new_E2968_ & new_E2978_;
  assign new_E2988_ = ~new_E2968_ & ~new_E2978_;
  assign new_E2989_ = new_E3010_ | new_E3009_;
  assign new_E2990_ = new_E2956_ | new_E2989_;
  assign new_E2991_ = new_E3014_ | new_E3013_;
  assign new_E2992_ = ~new_E2956_ & new_E2991_;
  assign new_E2993_ = new_E3012_ | new_E3011_;
  assign new_E2994_ = new_E2956_ & new_E2993_;
  assign new_E2995_ = new_E2954_ & ~new_E2964_;
  assign new_E2996_ = ~new_E2954_ & new_E2964_;
  assign new_E2997_ = ~new_E2953_ | ~new_E2978_;
  assign new_E2998_ = new_E2964_ & new_E2997_;
  assign new_E2999_ = ~new_E2964_ & ~new_E2998_;
  assign new_E3000_ = new_E2964_ | new_E2997_;
  assign new_E3001_ = ~new_E2954_ & new_E2955_;
  assign new_E3002_ = new_E2954_ & ~new_E2955_;
  assign new_E3003_ = new_E2971_ | new_E3008_;
  assign new_E3004_ = ~new_E2971_ & ~new_E3007_;
  assign new_E3005_ = new_E2954_ | new_E2971_;
  assign new_E3006_ = new_E2954_ | new_E2955_;
  assign new_E3007_ = new_E2971_ & new_E3008_;
  assign new_E3008_ = ~new_E2953_ | ~new_E2978_;
  assign new_E3009_ = new_E2986_ & new_E3006_;
  assign new_E3010_ = ~new_E2986_ & ~new_E3006_;
  assign new_E3011_ = new_E3015_ | new_E3016_;
  assign new_E3012_ = ~new_E2957_ & new_E2971_;
  assign new_E3013_ = new_E3017_ | new_E3018_;
  assign new_E3014_ = new_E2957_ & new_E2971_;
  assign new_E3015_ = ~new_E2957_ & ~new_E2971_;
  assign new_E3016_ = new_E2957_ & ~new_E2971_;
  assign new_E3017_ = new_E2957_ & ~new_E2971_;
  assign new_E3018_ = ~new_E2957_ & new_E2971_;
  assign new_E3019_ = new_F8706_;
  assign new_E3020_ = new_F8773_;
  assign new_E3021_ = new_F8840_;
  assign new_E3022_ = new_F8907_;
  assign new_E3023_ = new_F8974_;
  assign new_E3024_ = new_F9041_;
  assign new_E3025_ = new_E3032_ & new_E3031_;
  assign new_E3026_ = new_E3034_ | new_E3033_;
  assign new_E3027_ = new_E3036_ | new_E3035_;
  assign new_E3028_ = new_E3038_ & new_E3037_;
  assign new_E3029_ = new_E3038_ & new_E3039_;
  assign new_E3030_ = new_E3031_ | new_E3040_;
  assign new_E3031_ = new_E3020_ | new_E3043_;
  assign new_E3032_ = new_E3042_ | new_E3041_;
  assign new_E3033_ = new_E3047_ & new_E3046_;
  assign new_E3034_ = new_E3045_ & new_E3044_;
  assign new_E3035_ = new_E3050_ | new_E3049_;
  assign new_E3036_ = new_E3045_ & new_E3048_;
  assign new_E3037_ = new_E3020_ | new_E3053_;
  assign new_E3038_ = new_E3052_ | new_E3051_;
  assign new_E3039_ = new_E3055_ | new_E3054_;
  assign new_E3040_ = ~new_E3031_ & new_E3057_;
  assign new_E3041_ = ~new_E3033_ & new_E3045_;
  assign new_E3042_ = new_E3033_ & ~new_E3045_;
  assign new_E3043_ = new_E3019_ & ~new_E3020_;
  assign new_E3044_ = ~new_E3066_ | ~new_E3067_;
  assign new_E3045_ = new_E3059_ | new_E3061_;
  assign new_E3046_ = new_E3069_ | new_E3068_;
  assign new_E3047_ = new_E3063_ | new_E3062_;
  assign new_E3048_ = ~new_E3071_ | ~new_E3070_;
  assign new_E3049_ = ~new_E3072_ & new_E3073_;
  assign new_E3050_ = new_E3072_ & ~new_E3073_;
  assign new_E3051_ = ~new_E3019_ & new_E3020_;
  assign new_E3052_ = new_E3019_ & ~new_E3020_;
  assign new_E3053_ = ~new_E3035_ | new_E3045_;
  assign new_E3054_ = new_E3035_ & new_E3045_;
  assign new_E3055_ = ~new_E3035_ & ~new_E3045_;
  assign new_E3056_ = new_E3077_ | new_E3076_;
  assign new_E3057_ = new_E3023_ | new_E3056_;
  assign new_E3058_ = new_E3081_ | new_E3080_;
  assign new_E3059_ = ~new_E3023_ & new_E3058_;
  assign new_E3060_ = new_E3079_ | new_E3078_;
  assign new_E3061_ = new_E3023_ & new_E3060_;
  assign new_E3062_ = new_E3021_ & ~new_E3031_;
  assign new_E3063_ = ~new_E3021_ & new_E3031_;
  assign new_E3064_ = ~new_E3020_ | ~new_E3045_;
  assign new_E3065_ = new_E3031_ & new_E3064_;
  assign new_E3066_ = ~new_E3031_ & ~new_E3065_;
  assign new_E3067_ = new_E3031_ | new_E3064_;
  assign new_E3068_ = ~new_E3021_ & new_E3022_;
  assign new_E3069_ = new_E3021_ & ~new_E3022_;
  assign new_E3070_ = new_E3038_ | new_E3075_;
  assign new_E3071_ = ~new_E3038_ & ~new_E3074_;
  assign new_E3072_ = new_E3021_ | new_E3038_;
  assign new_E3073_ = new_E3021_ | new_E3022_;
  assign new_E3074_ = new_E3038_ & new_E3075_;
  assign new_E3075_ = ~new_E3020_ | ~new_E3045_;
  assign new_E3076_ = new_E3053_ & new_E3073_;
  assign new_E3077_ = ~new_E3053_ & ~new_E3073_;
  assign new_E3078_ = new_E3082_ | new_E3083_;
  assign new_E3079_ = ~new_E3024_ & new_E3038_;
  assign new_E3080_ = new_E3084_ | new_E3085_;
  assign new_E3081_ = new_E3024_ & new_E3038_;
  assign new_E3082_ = ~new_E3024_ & ~new_E3038_;
  assign new_E3083_ = new_E3024_ & ~new_E3038_;
  assign new_E3084_ = new_E3024_ & ~new_E3038_;
  assign new_E3085_ = ~new_E3024_ & new_E3038_;
  assign new_E3086_ = new_F9108_;
  assign new_E3087_ = new_F9175_;
  assign new_E3088_ = new_F9242_;
  assign new_E3089_ = new_F9309_;
  assign new_E3090_ = new_F9376_;
  assign new_E3091_ = new_F9443_;
  assign new_E3092_ = new_E3099_ & new_E3098_;
  assign new_E3093_ = new_E3101_ | new_E3100_;
  assign new_E3094_ = new_E3103_ | new_E3102_;
  assign new_E3095_ = new_E3105_ & new_E3104_;
  assign new_E3096_ = new_E3105_ & new_E3106_;
  assign new_E3097_ = new_E3098_ | new_E3107_;
  assign new_E3098_ = new_E3087_ | new_E3110_;
  assign new_E3099_ = new_E3109_ | new_E3108_;
  assign new_E3100_ = new_E3114_ & new_E3113_;
  assign new_E3101_ = new_E3112_ & new_E3111_;
  assign new_E3102_ = new_E3117_ | new_E3116_;
  assign new_E3103_ = new_E3112_ & new_E3115_;
  assign new_E3104_ = new_E3087_ | new_E3120_;
  assign new_E3105_ = new_E3119_ | new_E3118_;
  assign new_E3106_ = new_E3122_ | new_E3121_;
  assign new_E3107_ = ~new_E3098_ & new_E3124_;
  assign new_E3108_ = ~new_E3100_ & new_E3112_;
  assign new_E3109_ = new_E3100_ & ~new_E3112_;
  assign new_E3110_ = new_E3086_ & ~new_E3087_;
  assign new_E3111_ = ~new_E3133_ | ~new_E3134_;
  assign new_E3112_ = new_E3126_ | new_E3128_;
  assign new_E3113_ = new_E3136_ | new_E3135_;
  assign new_E3114_ = new_E3130_ | new_E3129_;
  assign new_E3115_ = ~new_E3138_ | ~new_E3137_;
  assign new_E3116_ = ~new_E3139_ & new_E3140_;
  assign new_E3117_ = new_E3139_ & ~new_E3140_;
  assign new_E3118_ = ~new_E3086_ & new_E3087_;
  assign new_E3119_ = new_E3086_ & ~new_E3087_;
  assign new_E3120_ = ~new_E3102_ | new_E3112_;
  assign new_E3121_ = new_E3102_ & new_E3112_;
  assign new_E3122_ = ~new_E3102_ & ~new_E3112_;
  assign new_E3123_ = new_E3144_ | new_E3143_;
  assign new_E3124_ = new_E3090_ | new_E3123_;
  assign new_E3125_ = new_E3148_ | new_E3147_;
  assign new_E3126_ = ~new_E3090_ & new_E3125_;
  assign new_E3127_ = new_E3146_ | new_E3145_;
  assign new_E3128_ = new_E3090_ & new_E3127_;
  assign new_E3129_ = new_E3088_ & ~new_E3098_;
  assign new_E3130_ = ~new_E3088_ & new_E3098_;
  assign new_E3131_ = ~new_E3087_ | ~new_E3112_;
  assign new_E3132_ = new_E3098_ & new_E3131_;
  assign new_E3133_ = ~new_E3098_ & ~new_E3132_;
  assign new_E3134_ = new_E3098_ | new_E3131_;
  assign new_E3135_ = ~new_E3088_ & new_E3089_;
  assign new_E3136_ = new_E3088_ & ~new_E3089_;
  assign new_E3137_ = new_E3105_ | new_E3142_;
  assign new_E3138_ = ~new_E3105_ & ~new_E3141_;
  assign new_E3139_ = new_E3088_ | new_E3105_;
  assign new_E3140_ = new_E3088_ | new_E3089_;
  assign new_E3141_ = new_E3105_ & new_E3142_;
  assign new_E3142_ = ~new_E3087_ | ~new_E3112_;
  assign new_E3143_ = new_E3120_ & new_E3140_;
  assign new_E3144_ = ~new_E3120_ & ~new_E3140_;
  assign new_E3145_ = new_E3149_ | new_E3150_;
  assign new_E3146_ = ~new_E3091_ & new_E3105_;
  assign new_E3147_ = new_E3151_ | new_E3152_;
  assign new_E3148_ = new_E3091_ & new_E3105_;
  assign new_E3149_ = ~new_E3091_ & ~new_E3105_;
  assign new_E3150_ = new_E3091_ & ~new_E3105_;
  assign new_E3151_ = new_E3091_ & ~new_E3105_;
  assign new_E3152_ = ~new_E3091_ & new_E3105_;
  assign new_E3153_ = new_F9510_;
  assign new_E3154_ = new_F9577_;
  assign new_E3155_ = new_F9644_;
  assign new_E3156_ = new_F9711_;
  assign new_E3157_ = new_F9778_;
  assign new_E3158_ = new_F9845_;
  assign new_E3159_ = new_E3166_ & new_E3165_;
  assign new_E3160_ = new_E3168_ | new_E3167_;
  assign new_E3161_ = new_E3170_ | new_E3169_;
  assign new_E3162_ = new_E3172_ & new_E3171_;
  assign new_E3163_ = new_E3172_ & new_E3173_;
  assign new_E3164_ = new_E3165_ | new_E3174_;
  assign new_E3165_ = new_E3154_ | new_E3177_;
  assign new_E3166_ = new_E3176_ | new_E3175_;
  assign new_E3167_ = new_E3181_ & new_E3180_;
  assign new_E3168_ = new_E3179_ & new_E3178_;
  assign new_E3169_ = new_E3184_ | new_E3183_;
  assign new_E3170_ = new_E3179_ & new_E3182_;
  assign new_E3171_ = new_E3154_ | new_E3187_;
  assign new_E3172_ = new_E3186_ | new_E3185_;
  assign new_E3173_ = new_E3189_ | new_E3188_;
  assign new_E3174_ = ~new_E3165_ & new_E3191_;
  assign new_E3175_ = ~new_E3167_ & new_E3179_;
  assign new_E3176_ = new_E3167_ & ~new_E3179_;
  assign new_E3177_ = new_E3153_ & ~new_E3154_;
  assign new_E3178_ = ~new_E3200_ | ~new_E3201_;
  assign new_E3179_ = new_E3193_ | new_E3195_;
  assign new_E3180_ = new_E3203_ | new_E3202_;
  assign new_E3181_ = new_E3197_ | new_E3196_;
  assign new_E3182_ = ~new_E3205_ | ~new_E3204_;
  assign new_E3183_ = ~new_E3206_ & new_E3207_;
  assign new_E3184_ = new_E3206_ & ~new_E3207_;
  assign new_E3185_ = ~new_E3153_ & new_E3154_;
  assign new_E3186_ = new_E3153_ & ~new_E3154_;
  assign new_E3187_ = ~new_E3169_ | new_E3179_;
  assign new_E3188_ = new_E3169_ & new_E3179_;
  assign new_E3189_ = ~new_E3169_ & ~new_E3179_;
  assign new_E3190_ = new_E3211_ | new_E3210_;
  assign new_E3191_ = new_E3157_ | new_E3190_;
  assign new_E3192_ = new_E3215_ | new_E3214_;
  assign new_E3193_ = ~new_E3157_ & new_E3192_;
  assign new_E3194_ = new_E3213_ | new_E3212_;
  assign new_E3195_ = new_E3157_ & new_E3194_;
  assign new_E3196_ = new_E3155_ & ~new_E3165_;
  assign new_E3197_ = ~new_E3155_ & new_E3165_;
  assign new_E3198_ = ~new_E3154_ | ~new_E3179_;
  assign new_E3199_ = new_E3165_ & new_E3198_;
  assign new_E3200_ = ~new_E3165_ & ~new_E3199_;
  assign new_E3201_ = new_E3165_ | new_E3198_;
  assign new_E3202_ = ~new_E3155_ & new_E3156_;
  assign new_E3203_ = new_E3155_ & ~new_E3156_;
  assign new_E3204_ = new_E3172_ | new_E3209_;
  assign new_E3205_ = ~new_E3172_ & ~new_E3208_;
  assign new_E3206_ = new_E3155_ | new_E3172_;
  assign new_E3207_ = new_E3155_ | new_E3156_;
  assign new_E3208_ = new_E3172_ & new_E3209_;
  assign new_E3209_ = ~new_E3154_ | ~new_E3179_;
  assign new_E3210_ = new_E3187_ & new_E3207_;
  assign new_E3211_ = ~new_E3187_ & ~new_E3207_;
  assign new_E3212_ = new_E3216_ | new_E3217_;
  assign new_E3213_ = ~new_E3158_ & new_E3172_;
  assign new_E3214_ = new_E3218_ | new_E3219_;
  assign new_E3215_ = new_E3158_ & new_E3172_;
  assign new_E3216_ = ~new_E3158_ & ~new_E3172_;
  assign new_E3217_ = new_E3158_ & ~new_E3172_;
  assign new_E3218_ = new_E3158_ & ~new_E3172_;
  assign new_E3219_ = ~new_E3158_ & new_E3172_;
  assign new_E3220_ = new_F9912_;
  assign new_E3221_ = new_F9979_;
  assign new_E3222_ = new_G47_;
  assign new_E3223_ = new_G114_;
  assign new_E3224_ = new_G181_;
  assign new_E3225_ = new_G248_;
  assign new_E3226_ = new_E3233_ & new_E3232_;
  assign new_E3227_ = new_E3235_ | new_E3234_;
  assign new_E3228_ = new_E3237_ | new_E3236_;
  assign new_E3229_ = new_E3239_ & new_E3238_;
  assign new_E3230_ = new_E3239_ & new_E3240_;
  assign new_E3231_ = new_E3232_ | new_E3241_;
  assign new_E3232_ = new_E3221_ | new_E3244_;
  assign new_E3233_ = new_E3243_ | new_E3242_;
  assign new_E3234_ = new_E3248_ & new_E3247_;
  assign new_E3235_ = new_E3246_ & new_E3245_;
  assign new_E3236_ = new_E3251_ | new_E3250_;
  assign new_E3237_ = new_E3246_ & new_E3249_;
  assign new_E3238_ = new_E3221_ | new_E3254_;
  assign new_E3239_ = new_E3253_ | new_E3252_;
  assign new_E3240_ = new_E3256_ | new_E3255_;
  assign new_E3241_ = ~new_E3232_ & new_E3258_;
  assign new_E3242_ = ~new_E3234_ & new_E3246_;
  assign new_E3243_ = new_E3234_ & ~new_E3246_;
  assign new_E3244_ = new_E3220_ & ~new_E3221_;
  assign new_E3245_ = ~new_E3267_ | ~new_E3268_;
  assign new_E3246_ = new_E3260_ | new_E3262_;
  assign new_E3247_ = new_E3270_ | new_E3269_;
  assign new_E3248_ = new_E3264_ | new_E3263_;
  assign new_E3249_ = ~new_E3272_ | ~new_E3271_;
  assign new_E3250_ = ~new_E3273_ & new_E3274_;
  assign new_E3251_ = new_E3273_ & ~new_E3274_;
  assign new_E3252_ = ~new_E3220_ & new_E3221_;
  assign new_E3253_ = new_E3220_ & ~new_E3221_;
  assign new_E3254_ = ~new_E3236_ | new_E3246_;
  assign new_E3255_ = new_E3236_ & new_E3246_;
  assign new_E3256_ = ~new_E3236_ & ~new_E3246_;
  assign new_E3257_ = new_E3278_ | new_E3277_;
  assign new_E3258_ = new_E3224_ | new_E3257_;
  assign new_E3259_ = new_E3282_ | new_E3281_;
  assign new_E3260_ = ~new_E3224_ & new_E3259_;
  assign new_E3261_ = new_E3280_ | new_E3279_;
  assign new_E3262_ = new_E3224_ & new_E3261_;
  assign new_E3263_ = new_E3222_ & ~new_E3232_;
  assign new_E3264_ = ~new_E3222_ & new_E3232_;
  assign new_E3265_ = ~new_E3221_ | ~new_E3246_;
  assign new_E3266_ = new_E3232_ & new_E3265_;
  assign new_E3267_ = ~new_E3232_ & ~new_E3266_;
  assign new_E3268_ = new_E3232_ | new_E3265_;
  assign new_E3269_ = ~new_E3222_ & new_E3223_;
  assign new_E3270_ = new_E3222_ & ~new_E3223_;
  assign new_E3271_ = new_E3239_ | new_E3276_;
  assign new_E3272_ = ~new_E3239_ & ~new_E3275_;
  assign new_E3273_ = new_E3222_ | new_E3239_;
  assign new_E3274_ = new_E3222_ | new_E3223_;
  assign new_E3275_ = new_E3239_ & new_E3276_;
  assign new_E3276_ = ~new_E3221_ | ~new_E3246_;
  assign new_E3277_ = new_E3254_ & new_E3274_;
  assign new_E3278_ = ~new_E3254_ & ~new_E3274_;
  assign new_E3279_ = new_E3283_ | new_E3284_;
  assign new_E3280_ = ~new_E3225_ & new_E3239_;
  assign new_E3281_ = new_E3285_ | new_E3286_;
  assign new_E3282_ = new_E3225_ & new_E3239_;
  assign new_E3283_ = ~new_E3225_ & ~new_E3239_;
  assign new_E3284_ = new_E3225_ & ~new_E3239_;
  assign new_E3285_ = new_E3225_ & ~new_E3239_;
  assign new_E3286_ = ~new_E3225_ & new_E3239_;
  assign new_E3287_ = new_G315_;
  assign new_E3288_ = new_G382_;
  assign new_E3289_ = new_G449_;
  assign new_E3290_ = new_G516_;
  assign new_E3291_ = new_G583_;
  assign new_E3292_ = new_G650_;
  assign new_E3293_ = new_E3300_ & new_E3299_;
  assign new_E3294_ = new_E3302_ | new_E3301_;
  assign new_E3295_ = new_E3304_ | new_E3303_;
  assign new_E3296_ = new_E3306_ & new_E3305_;
  assign new_E3297_ = new_E3306_ & new_E3307_;
  assign new_E3298_ = new_E3299_ | new_E3308_;
  assign new_E3299_ = new_E3288_ | new_E3311_;
  assign new_E3300_ = new_E3310_ | new_E3309_;
  assign new_E3301_ = new_E3315_ & new_E3314_;
  assign new_E3302_ = new_E3313_ & new_E3312_;
  assign new_E3303_ = new_E3318_ | new_E3317_;
  assign new_E3304_ = new_E3313_ & new_E3316_;
  assign new_E3305_ = new_E3288_ | new_E3321_;
  assign new_E3306_ = new_E3320_ | new_E3319_;
  assign new_E3307_ = new_E3323_ | new_E3322_;
  assign new_E3308_ = ~new_E3299_ & new_E3325_;
  assign new_E3309_ = ~new_E3301_ & new_E3313_;
  assign new_E3310_ = new_E3301_ & ~new_E3313_;
  assign new_E3311_ = new_E3287_ & ~new_E3288_;
  assign new_E3312_ = ~new_E3334_ | ~new_E3335_;
  assign new_E3313_ = new_E3327_ | new_E3329_;
  assign new_E3314_ = new_E3337_ | new_E3336_;
  assign new_E3315_ = new_E3331_ | new_E3330_;
  assign new_E3316_ = ~new_E3339_ | ~new_E3338_;
  assign new_E3317_ = ~new_E3340_ & new_E3341_;
  assign new_E3318_ = new_E3340_ & ~new_E3341_;
  assign new_E3319_ = ~new_E3287_ & new_E3288_;
  assign new_E3320_ = new_E3287_ & ~new_E3288_;
  assign new_E3321_ = ~new_E3303_ | new_E3313_;
  assign new_E3322_ = new_E3303_ & new_E3313_;
  assign new_E3323_ = ~new_E3303_ & ~new_E3313_;
  assign new_E3324_ = new_E3345_ | new_E3344_;
  assign new_E3325_ = new_E3291_ | new_E3324_;
  assign new_E3326_ = new_E3349_ | new_E3348_;
  assign new_E3327_ = ~new_E3291_ & new_E3326_;
  assign new_E3328_ = new_E3347_ | new_E3346_;
  assign new_E3329_ = new_E3291_ & new_E3328_;
  assign new_E3330_ = new_E3289_ & ~new_E3299_;
  assign new_E3331_ = ~new_E3289_ & new_E3299_;
  assign new_E3332_ = ~new_E3288_ | ~new_E3313_;
  assign new_E3333_ = new_E3299_ & new_E3332_;
  assign new_E3334_ = ~new_E3299_ & ~new_E3333_;
  assign new_E3335_ = new_E3299_ | new_E3332_;
  assign new_E3336_ = ~new_E3289_ & new_E3290_;
  assign new_E3337_ = new_E3289_ & ~new_E3290_;
  assign new_E3338_ = new_E3306_ | new_E3343_;
  assign new_E3339_ = ~new_E3306_ & ~new_E3342_;
  assign new_E3340_ = new_E3289_ | new_E3306_;
  assign new_E3341_ = new_E3289_ | new_E3290_;
  assign new_E3342_ = new_E3306_ & new_E3343_;
  assign new_E3343_ = ~new_E3288_ | ~new_E3313_;
  assign new_E3344_ = new_E3321_ & new_E3341_;
  assign new_E3345_ = ~new_E3321_ & ~new_E3341_;
  assign new_E3346_ = new_E3350_ | new_E3351_;
  assign new_E3347_ = ~new_E3292_ & new_E3306_;
  assign new_E3348_ = new_E3352_ | new_E3353_;
  assign new_E3349_ = new_E3292_ & new_E3306_;
  assign new_E3350_ = ~new_E3292_ & ~new_E3306_;
  assign new_E3351_ = new_E3292_ & ~new_E3306_;
  assign new_E3352_ = new_E3292_ & ~new_E3306_;
  assign new_E3353_ = ~new_E3292_ & new_E3306_;
  assign new_E3354_ = new_G717_;
  assign new_E3355_ = new_G784_;
  assign new_E3356_ = new_G851_;
  assign new_E3357_ = new_G918_;
  assign new_E3358_ = new_G985_;
  assign new_E3359_ = new_G1052_;
  assign new_E3360_ = new_E3367_ & new_E3366_;
  assign new_E3361_ = new_E3369_ | new_E3368_;
  assign new_E3362_ = new_E3371_ | new_E3370_;
  assign new_E3363_ = new_E3373_ & new_E3372_;
  assign new_E3364_ = new_E3373_ & new_E3374_;
  assign new_E3365_ = new_E3366_ | new_E3375_;
  assign new_E3366_ = new_E3355_ | new_E3378_;
  assign new_E3367_ = new_E3377_ | new_E3376_;
  assign new_E3368_ = new_E3382_ & new_E3381_;
  assign new_E3369_ = new_E3380_ & new_E3379_;
  assign new_E3370_ = new_E3385_ | new_E3384_;
  assign new_E3371_ = new_E3380_ & new_E3383_;
  assign new_E3372_ = new_E3355_ | new_E3388_;
  assign new_E3373_ = new_E3387_ | new_E3386_;
  assign new_E3374_ = new_E3390_ | new_E3389_;
  assign new_E3375_ = ~new_E3366_ & new_E3392_;
  assign new_E3376_ = ~new_E3368_ & new_E3380_;
  assign new_E3377_ = new_E3368_ & ~new_E3380_;
  assign new_E3378_ = new_E3354_ & ~new_E3355_;
  assign new_E3379_ = ~new_E3401_ | ~new_E3402_;
  assign new_E3380_ = new_E3394_ | new_E3396_;
  assign new_E3381_ = new_E3404_ | new_E3403_;
  assign new_E3382_ = new_E3398_ | new_E3397_;
  assign new_E3383_ = ~new_E3406_ | ~new_E3405_;
  assign new_E3384_ = ~new_E3407_ & new_E3408_;
  assign new_E3385_ = new_E3407_ & ~new_E3408_;
  assign new_E3386_ = ~new_E3354_ & new_E3355_;
  assign new_E3387_ = new_E3354_ & ~new_E3355_;
  assign new_E3388_ = ~new_E3370_ | new_E3380_;
  assign new_E3389_ = new_E3370_ & new_E3380_;
  assign new_E3390_ = ~new_E3370_ & ~new_E3380_;
  assign new_E3391_ = new_E3412_ | new_E3411_;
  assign new_E3392_ = new_E3358_ | new_E3391_;
  assign new_E3393_ = new_E3416_ | new_E3415_;
  assign new_E3394_ = ~new_E3358_ & new_E3393_;
  assign new_E3395_ = new_E3414_ | new_E3413_;
  assign new_E3396_ = new_E3358_ & new_E3395_;
  assign new_E3397_ = new_E3356_ & ~new_E3366_;
  assign new_E3398_ = ~new_E3356_ & new_E3366_;
  assign new_E3399_ = ~new_E3355_ | ~new_E3380_;
  assign new_E3400_ = new_E3366_ & new_E3399_;
  assign new_E3401_ = ~new_E3366_ & ~new_E3400_;
  assign new_E3402_ = new_E3366_ | new_E3399_;
  assign new_E3403_ = ~new_E3356_ & new_E3357_;
  assign new_E3404_ = new_E3356_ & ~new_E3357_;
  assign new_E3405_ = new_E3373_ | new_E3410_;
  assign new_E3406_ = ~new_E3373_ & ~new_E3409_;
  assign new_E3407_ = new_E3356_ | new_E3373_;
  assign new_E3408_ = new_E3356_ | new_E3357_;
  assign new_E3409_ = new_E3373_ & new_E3410_;
  assign new_E3410_ = ~new_E3355_ | ~new_E3380_;
  assign new_E3411_ = new_E3388_ & new_E3408_;
  assign new_E3412_ = ~new_E3388_ & ~new_E3408_;
  assign new_E3413_ = new_E3417_ | new_E3418_;
  assign new_E3414_ = ~new_E3359_ & new_E3373_;
  assign new_E3415_ = new_E3419_ | new_E3420_;
  assign new_E3416_ = new_E3359_ & new_E3373_;
  assign new_E3417_ = ~new_E3359_ & ~new_E3373_;
  assign new_E3418_ = new_E3359_ & ~new_E3373_;
  assign new_E3419_ = new_E3359_ & ~new_E3373_;
  assign new_E3420_ = ~new_E3359_ & new_E3373_;
  assign new_E3421_ = new_G1119_;
  assign new_E3422_ = new_G1186_;
  assign new_E3423_ = new_G1253_;
  assign new_E3424_ = new_G1320_;
  assign new_E3425_ = new_G1387_;
  assign new_E3426_ = new_G1454_;
  assign new_E3427_ = new_E3434_ & new_E3433_;
  assign new_E3428_ = new_E3436_ | new_E3435_;
  assign new_E3429_ = new_E3438_ | new_E3437_;
  assign new_E3430_ = new_E3440_ & new_E3439_;
  assign new_E3431_ = new_E3440_ & new_E3441_;
  assign new_E3432_ = new_E3433_ | new_E3442_;
  assign new_E3433_ = new_E3422_ | new_E3445_;
  assign new_E3434_ = new_E3444_ | new_E3443_;
  assign new_E3435_ = new_E3449_ & new_E3448_;
  assign new_E3436_ = new_E3447_ & new_E3446_;
  assign new_E3437_ = new_E3452_ | new_E3451_;
  assign new_E3438_ = new_E3447_ & new_E3450_;
  assign new_E3439_ = new_E3422_ | new_E3455_;
  assign new_E3440_ = new_E3454_ | new_E3453_;
  assign new_E3441_ = new_E3457_ | new_E3456_;
  assign new_E3442_ = ~new_E3433_ & new_E3459_;
  assign new_E3443_ = ~new_E3435_ & new_E3447_;
  assign new_E3444_ = new_E3435_ & ~new_E3447_;
  assign new_E3445_ = new_E3421_ & ~new_E3422_;
  assign new_E3446_ = ~new_E3468_ | ~new_E3469_;
  assign new_E3447_ = new_E3461_ | new_E3463_;
  assign new_E3448_ = new_E3471_ | new_E3470_;
  assign new_E3449_ = new_E3465_ | new_E3464_;
  assign new_E3450_ = ~new_E3473_ | ~new_E3472_;
  assign new_E3451_ = ~new_E3474_ & new_E3475_;
  assign new_E3452_ = new_E3474_ & ~new_E3475_;
  assign new_E3453_ = ~new_E3421_ & new_E3422_;
  assign new_E3454_ = new_E3421_ & ~new_E3422_;
  assign new_E3455_ = ~new_E3437_ | new_E3447_;
  assign new_E3456_ = new_E3437_ & new_E3447_;
  assign new_E3457_ = ~new_E3437_ & ~new_E3447_;
  assign new_E3458_ = new_E3479_ | new_E3478_;
  assign new_E3459_ = new_E3425_ | new_E3458_;
  assign new_E3460_ = new_E3483_ | new_E3482_;
  assign new_E3461_ = ~new_E3425_ & new_E3460_;
  assign new_E3462_ = new_E3481_ | new_E3480_;
  assign new_E3463_ = new_E3425_ & new_E3462_;
  assign new_E3464_ = new_E3423_ & ~new_E3433_;
  assign new_E3465_ = ~new_E3423_ & new_E3433_;
  assign new_E3466_ = ~new_E3422_ | ~new_E3447_;
  assign new_E3467_ = new_E3433_ & new_E3466_;
  assign new_E3468_ = ~new_E3433_ & ~new_E3467_;
  assign new_E3469_ = new_E3433_ | new_E3466_;
  assign new_E3470_ = ~new_E3423_ & new_E3424_;
  assign new_E3471_ = new_E3423_ & ~new_E3424_;
  assign new_E3472_ = new_E3440_ | new_E3477_;
  assign new_E3473_ = ~new_E3440_ & ~new_E3476_;
  assign new_E3474_ = new_E3423_ | new_E3440_;
  assign new_E3475_ = new_E3423_ | new_E3424_;
  assign new_E3476_ = new_E3440_ & new_E3477_;
  assign new_E3477_ = ~new_E3422_ | ~new_E3447_;
  assign new_E3478_ = new_E3455_ & new_E3475_;
  assign new_E3479_ = ~new_E3455_ & ~new_E3475_;
  assign new_E3480_ = new_E3484_ | new_E3485_;
  assign new_E3481_ = ~new_E3426_ & new_E3440_;
  assign new_E3482_ = new_E3486_ | new_E3487_;
  assign new_E3483_ = new_E3426_ & new_E3440_;
  assign new_E3484_ = ~new_E3426_ & ~new_E3440_;
  assign new_E3485_ = new_E3426_ & ~new_E3440_;
  assign new_E3486_ = new_E3426_ & ~new_E3440_;
  assign new_E3487_ = ~new_E3426_ & new_E3440_;
  assign new_E3488_ = new_G1521_;
  assign new_E3489_ = new_G1588_;
  assign new_E3490_ = new_G1655_;
  assign new_E3491_ = new_G1722_;
  assign new_E3492_ = new_G1789_;
  assign new_E3493_ = new_G1856_;
  assign new_E3494_ = new_E3501_ & new_E3500_;
  assign new_E3495_ = new_E3503_ | new_E3502_;
  assign new_E3496_ = new_E3505_ | new_E3504_;
  assign new_E3497_ = new_E3507_ & new_E3506_;
  assign new_E3498_ = new_E3507_ & new_E3508_;
  assign new_E3499_ = new_E3500_ | new_E3509_;
  assign new_E3500_ = new_E3489_ | new_E3512_;
  assign new_E3501_ = new_E3511_ | new_E3510_;
  assign new_E3502_ = new_E3516_ & new_E3515_;
  assign new_E3503_ = new_E3514_ & new_E3513_;
  assign new_E3504_ = new_E3519_ | new_E3518_;
  assign new_E3505_ = new_E3514_ & new_E3517_;
  assign new_E3506_ = new_E3489_ | new_E3522_;
  assign new_E3507_ = new_E3521_ | new_E3520_;
  assign new_E3508_ = new_E3524_ | new_E3523_;
  assign new_E3509_ = ~new_E3500_ & new_E3526_;
  assign new_E3510_ = ~new_E3502_ & new_E3514_;
  assign new_E3511_ = new_E3502_ & ~new_E3514_;
  assign new_E3512_ = new_E3488_ & ~new_E3489_;
  assign new_E3513_ = ~new_E3535_ | ~new_E3536_;
  assign new_E3514_ = new_E3528_ | new_E3530_;
  assign new_E3515_ = new_E3538_ | new_E3537_;
  assign new_E3516_ = new_E3532_ | new_E3531_;
  assign new_E3517_ = ~new_E3540_ | ~new_E3539_;
  assign new_E3518_ = ~new_E3541_ & new_E3542_;
  assign new_E3519_ = new_E3541_ & ~new_E3542_;
  assign new_E3520_ = ~new_E3488_ & new_E3489_;
  assign new_E3521_ = new_E3488_ & ~new_E3489_;
  assign new_E3522_ = ~new_E3504_ | new_E3514_;
  assign new_E3523_ = new_E3504_ & new_E3514_;
  assign new_E3524_ = ~new_E3504_ & ~new_E3514_;
  assign new_E3525_ = new_E3546_ | new_E3545_;
  assign new_E3526_ = new_E3492_ | new_E3525_;
  assign new_E3527_ = new_E3550_ | new_E3549_;
  assign new_E3528_ = ~new_E3492_ & new_E3527_;
  assign new_E3529_ = new_E3548_ | new_E3547_;
  assign new_E3530_ = new_E3492_ & new_E3529_;
  assign new_E3531_ = new_E3490_ & ~new_E3500_;
  assign new_E3532_ = ~new_E3490_ & new_E3500_;
  assign new_E3533_ = ~new_E3489_ | ~new_E3514_;
  assign new_E3534_ = new_E3500_ & new_E3533_;
  assign new_E3535_ = ~new_E3500_ & ~new_E3534_;
  assign new_E3536_ = new_E3500_ | new_E3533_;
  assign new_E3537_ = ~new_E3490_ & new_E3491_;
  assign new_E3538_ = new_E3490_ & ~new_E3491_;
  assign new_E3539_ = new_E3507_ | new_E3544_;
  assign new_E3540_ = ~new_E3507_ & ~new_E3543_;
  assign new_E3541_ = new_E3490_ | new_E3507_;
  assign new_E3542_ = new_E3490_ | new_E3491_;
  assign new_E3543_ = new_E3507_ & new_E3544_;
  assign new_E3544_ = ~new_E3489_ | ~new_E3514_;
  assign new_E3545_ = new_E3522_ & new_E3542_;
  assign new_E3546_ = ~new_E3522_ & ~new_E3542_;
  assign new_E3547_ = new_E3551_ | new_E3552_;
  assign new_E3548_ = ~new_E3493_ & new_E3507_;
  assign new_E3549_ = new_E3553_ | new_E3554_;
  assign new_E3550_ = new_E3493_ & new_E3507_;
  assign new_E3551_ = ~new_E3493_ & ~new_E3507_;
  assign new_E3552_ = new_E3493_ & ~new_E3507_;
  assign new_E3553_ = new_E3493_ & ~new_E3507_;
  assign new_E3554_ = ~new_E3493_ & new_E3507_;
  assign new_E3555_ = new_G1923_;
  assign new_E3556_ = new_G1990_;
  assign new_E3557_ = new_G2057_;
  assign new_E3558_ = new_G2124_;
  assign new_E3559_ = new_G2191_;
  assign new_E3560_ = new_G2258_;
  assign new_E3561_ = new_E3568_ & new_E3567_;
  assign new_E3562_ = new_E3570_ | new_E3569_;
  assign new_E3563_ = new_E3572_ | new_E3571_;
  assign new_E3564_ = new_E3574_ & new_E3573_;
  assign new_E3565_ = new_E3574_ & new_E3575_;
  assign new_E3566_ = new_E3567_ | new_E3576_;
  assign new_E3567_ = new_E3556_ | new_E3579_;
  assign new_E3568_ = new_E3578_ | new_E3577_;
  assign new_E3569_ = new_E3583_ & new_E3582_;
  assign new_E3570_ = new_E3581_ & new_E3580_;
  assign new_E3571_ = new_E3586_ | new_E3585_;
  assign new_E3572_ = new_E3581_ & new_E3584_;
  assign new_E3573_ = new_E3556_ | new_E3589_;
  assign new_E3574_ = new_E3588_ | new_E3587_;
  assign new_E3575_ = new_E3591_ | new_E3590_;
  assign new_E3576_ = ~new_E3567_ & new_E3593_;
  assign new_E3577_ = ~new_E3569_ & new_E3581_;
  assign new_E3578_ = new_E3569_ & ~new_E3581_;
  assign new_E3579_ = new_E3555_ & ~new_E3556_;
  assign new_E3580_ = ~new_E3602_ | ~new_E3603_;
  assign new_E3581_ = new_E3595_ | new_E3597_;
  assign new_E3582_ = new_E3605_ | new_E3604_;
  assign new_E3583_ = new_E3599_ | new_E3598_;
  assign new_E3584_ = ~new_E3607_ | ~new_E3606_;
  assign new_E3585_ = ~new_E3608_ & new_E3609_;
  assign new_E3586_ = new_E3608_ & ~new_E3609_;
  assign new_E3587_ = ~new_E3555_ & new_E3556_;
  assign new_E3588_ = new_E3555_ & ~new_E3556_;
  assign new_E3589_ = ~new_E3571_ | new_E3581_;
  assign new_E3590_ = new_E3571_ & new_E3581_;
  assign new_E3591_ = ~new_E3571_ & ~new_E3581_;
  assign new_E3592_ = new_E3613_ | new_E3612_;
  assign new_E3593_ = new_E3559_ | new_E3592_;
  assign new_E3594_ = new_E3617_ | new_E3616_;
  assign new_E3595_ = ~new_E3559_ & new_E3594_;
  assign new_E3596_ = new_E3615_ | new_E3614_;
  assign new_E3597_ = new_E3559_ & new_E3596_;
  assign new_E3598_ = new_E3557_ & ~new_E3567_;
  assign new_E3599_ = ~new_E3557_ & new_E3567_;
  assign new_E3600_ = ~new_E3556_ | ~new_E3581_;
  assign new_E3601_ = new_E3567_ & new_E3600_;
  assign new_E3602_ = ~new_E3567_ & ~new_E3601_;
  assign new_E3603_ = new_E3567_ | new_E3600_;
  assign new_E3604_ = ~new_E3557_ & new_E3558_;
  assign new_E3605_ = new_E3557_ & ~new_E3558_;
  assign new_E3606_ = new_E3574_ | new_E3611_;
  assign new_E3607_ = ~new_E3574_ & ~new_E3610_;
  assign new_E3608_ = new_E3557_ | new_E3574_;
  assign new_E3609_ = new_E3557_ | new_E3558_;
  assign new_E3610_ = new_E3574_ & new_E3611_;
  assign new_E3611_ = ~new_E3556_ | ~new_E3581_;
  assign new_E3612_ = new_E3589_ & new_E3609_;
  assign new_E3613_ = ~new_E3589_ & ~new_E3609_;
  assign new_E3614_ = new_E3618_ | new_E3619_;
  assign new_E3615_ = ~new_E3560_ & new_E3574_;
  assign new_E3616_ = new_E3620_ | new_E3621_;
  assign new_E3617_ = new_E3560_ & new_E3574_;
  assign new_E3618_ = ~new_E3560_ & ~new_E3574_;
  assign new_E3619_ = new_E3560_ & ~new_E3574_;
  assign new_E3620_ = new_E3560_ & ~new_E3574_;
  assign new_E3621_ = ~new_E3560_ & new_E3574_;
  assign new_E3622_ = new_G2325_;
  assign new_E3623_ = new_G2392_;
  assign new_E3624_ = new_G2459_;
  assign new_E3625_ = new_G2526_;
  assign new_E3626_ = new_G2593_;
  assign new_E3627_ = new_G2660_;
  assign new_E3628_ = new_E3635_ & new_E3634_;
  assign new_E3629_ = new_E3637_ | new_E3636_;
  assign new_E3630_ = new_E3639_ | new_E3638_;
  assign new_E3631_ = new_E3641_ & new_E3640_;
  assign new_E3632_ = new_E3641_ & new_E3642_;
  assign new_E3633_ = new_E3634_ | new_E3643_;
  assign new_E3634_ = new_E3623_ | new_E3646_;
  assign new_E3635_ = new_E3645_ | new_E3644_;
  assign new_E3636_ = new_E3650_ & new_E3649_;
  assign new_E3637_ = new_E3648_ & new_E3647_;
  assign new_E3638_ = new_E3653_ | new_E3652_;
  assign new_E3639_ = new_E3648_ & new_E3651_;
  assign new_E3640_ = new_E3623_ | new_E3656_;
  assign new_E3641_ = new_E3655_ | new_E3654_;
  assign new_E3642_ = new_E3658_ | new_E3657_;
  assign new_E3643_ = ~new_E3634_ & new_E3660_;
  assign new_E3644_ = ~new_E3636_ & new_E3648_;
  assign new_E3645_ = new_E3636_ & ~new_E3648_;
  assign new_E3646_ = new_E3622_ & ~new_E3623_;
  assign new_E3647_ = ~new_E3669_ | ~new_E3670_;
  assign new_E3648_ = new_E3662_ | new_E3664_;
  assign new_E3649_ = new_E3672_ | new_E3671_;
  assign new_E3650_ = new_E3666_ | new_E3665_;
  assign new_E3651_ = ~new_E3674_ | ~new_E3673_;
  assign new_E3652_ = ~new_E3675_ & new_E3676_;
  assign new_E3653_ = new_E3675_ & ~new_E3676_;
  assign new_E3654_ = ~new_E3622_ & new_E3623_;
  assign new_E3655_ = new_E3622_ & ~new_E3623_;
  assign new_E3656_ = ~new_E3638_ | new_E3648_;
  assign new_E3657_ = new_E3638_ & new_E3648_;
  assign new_E3658_ = ~new_E3638_ & ~new_E3648_;
  assign new_E3659_ = new_E3680_ | new_E3679_;
  assign new_E3660_ = new_E3626_ | new_E3659_;
  assign new_E3661_ = new_E3684_ | new_E3683_;
  assign new_E3662_ = ~new_E3626_ & new_E3661_;
  assign new_E3663_ = new_E3682_ | new_E3681_;
  assign new_E3664_ = new_E3626_ & new_E3663_;
  assign new_E3665_ = new_E3624_ & ~new_E3634_;
  assign new_E3666_ = ~new_E3624_ & new_E3634_;
  assign new_E3667_ = ~new_E3623_ | ~new_E3648_;
  assign new_E3668_ = new_E3634_ & new_E3667_;
  assign new_E3669_ = ~new_E3634_ & ~new_E3668_;
  assign new_E3670_ = new_E3634_ | new_E3667_;
  assign new_E3671_ = ~new_E3624_ & new_E3625_;
  assign new_E3672_ = new_E3624_ & ~new_E3625_;
  assign new_E3673_ = new_E3641_ | new_E3678_;
  assign new_E3674_ = ~new_E3641_ & ~new_E3677_;
  assign new_E3675_ = new_E3624_ | new_E3641_;
  assign new_E3676_ = new_E3624_ | new_E3625_;
  assign new_E3677_ = new_E3641_ & new_E3678_;
  assign new_E3678_ = ~new_E3623_ | ~new_E3648_;
  assign new_E3679_ = new_E3656_ & new_E3676_;
  assign new_E3680_ = ~new_E3656_ & ~new_E3676_;
  assign new_E3681_ = new_E3685_ | new_E3686_;
  assign new_E3682_ = ~new_E3627_ & new_E3641_;
  assign new_E3683_ = new_E3687_ | new_E3688_;
  assign new_E3684_ = new_E3627_ & new_E3641_;
  assign new_E3685_ = ~new_E3627_ & ~new_E3641_;
  assign new_E3686_ = new_E3627_ & ~new_E3641_;
  assign new_E3687_ = new_E3627_ & ~new_E3641_;
  assign new_E3688_ = ~new_E3627_ & new_E3641_;
  assign new_E3689_ = new_G2727_;
  assign new_E3690_ = new_G2794_;
  assign new_E3691_ = new_G2861_;
  assign new_E3692_ = new_G2928_;
  assign new_E3693_ = new_G2995_;
  assign new_E3694_ = new_G3062_;
  assign new_E3695_ = new_E3702_ & new_E3701_;
  assign new_E3696_ = new_E3704_ | new_E3703_;
  assign new_E3697_ = new_E3706_ | new_E3705_;
  assign new_E3698_ = new_E3708_ & new_E3707_;
  assign new_E3699_ = new_E3708_ & new_E3709_;
  assign new_E3700_ = new_E3701_ | new_E3710_;
  assign new_E3701_ = new_E3690_ | new_E3713_;
  assign new_E3702_ = new_E3712_ | new_E3711_;
  assign new_E3703_ = new_E3717_ & new_E3716_;
  assign new_E3704_ = new_E3715_ & new_E3714_;
  assign new_E3705_ = new_E3720_ | new_E3719_;
  assign new_E3706_ = new_E3715_ & new_E3718_;
  assign new_E3707_ = new_E3690_ | new_E3723_;
  assign new_E3708_ = new_E3722_ | new_E3721_;
  assign new_E3709_ = new_E3725_ | new_E3724_;
  assign new_E3710_ = ~new_E3701_ & new_E3727_;
  assign new_E3711_ = ~new_E3703_ & new_E3715_;
  assign new_E3712_ = new_E3703_ & ~new_E3715_;
  assign new_E3713_ = new_E3689_ & ~new_E3690_;
  assign new_E3714_ = ~new_E3736_ | ~new_E3737_;
  assign new_E3715_ = new_E3729_ | new_E3731_;
  assign new_E3716_ = new_E3739_ | new_E3738_;
  assign new_E3717_ = new_E3733_ | new_E3732_;
  assign new_E3718_ = ~new_E3741_ | ~new_E3740_;
  assign new_E3719_ = ~new_E3742_ & new_E3743_;
  assign new_E3720_ = new_E3742_ & ~new_E3743_;
  assign new_E3721_ = ~new_E3689_ & new_E3690_;
  assign new_E3722_ = new_E3689_ & ~new_E3690_;
  assign new_E3723_ = ~new_E3705_ | new_E3715_;
  assign new_E3724_ = new_E3705_ & new_E3715_;
  assign new_E3725_ = ~new_E3705_ & ~new_E3715_;
  assign new_E3726_ = new_E3747_ | new_E3746_;
  assign new_E3727_ = new_E3693_ | new_E3726_;
  assign new_E3728_ = new_E3751_ | new_E3750_;
  assign new_E3729_ = ~new_E3693_ & new_E3728_;
  assign new_E3730_ = new_E3749_ | new_E3748_;
  assign new_E3731_ = new_E3693_ & new_E3730_;
  assign new_E3732_ = new_E3691_ & ~new_E3701_;
  assign new_E3733_ = ~new_E3691_ & new_E3701_;
  assign new_E3734_ = ~new_E3690_ | ~new_E3715_;
  assign new_E3735_ = new_E3701_ & new_E3734_;
  assign new_E3736_ = ~new_E3701_ & ~new_E3735_;
  assign new_E3737_ = new_E3701_ | new_E3734_;
  assign new_E3738_ = ~new_E3691_ & new_E3692_;
  assign new_E3739_ = new_E3691_ & ~new_E3692_;
  assign new_E3740_ = new_E3708_ | new_E3745_;
  assign new_E3741_ = ~new_E3708_ & ~new_E3744_;
  assign new_E3742_ = new_E3691_ | new_E3708_;
  assign new_E3743_ = new_E3691_ | new_E3692_;
  assign new_E3744_ = new_E3708_ & new_E3745_;
  assign new_E3745_ = ~new_E3690_ | ~new_E3715_;
  assign new_E3746_ = new_E3723_ & new_E3743_;
  assign new_E3747_ = ~new_E3723_ & ~new_E3743_;
  assign new_E3748_ = new_E3752_ | new_E3753_;
  assign new_E3749_ = ~new_E3694_ & new_E3708_;
  assign new_E3750_ = new_E3754_ | new_E3755_;
  assign new_E3751_ = new_E3694_ & new_E3708_;
  assign new_E3752_ = ~new_E3694_ & ~new_E3708_;
  assign new_E3753_ = new_E3694_ & ~new_E3708_;
  assign new_E3754_ = new_E3694_ & ~new_E3708_;
  assign new_E3755_ = ~new_E3694_ & new_E3708_;
  assign new_E3756_ = new_G3129_;
  assign new_E3757_ = new_G3196_;
  assign new_E3758_ = new_G3263_;
  assign new_E3759_ = new_G3330_;
  assign new_E3760_ = new_G3397_;
  assign new_E3761_ = new_G3464_;
  assign new_E3762_ = new_E3769_ & new_E3768_;
  assign new_E3763_ = new_E3771_ | new_E3770_;
  assign new_E3764_ = new_E3773_ | new_E3772_;
  assign new_E3765_ = new_E3775_ & new_E3774_;
  assign new_E3766_ = new_E3775_ & new_E3776_;
  assign new_E3767_ = new_E3768_ | new_E3777_;
  assign new_E3768_ = new_E3757_ | new_E3780_;
  assign new_E3769_ = new_E3779_ | new_E3778_;
  assign new_E3770_ = new_E3784_ & new_E3783_;
  assign new_E3771_ = new_E3782_ & new_E3781_;
  assign new_E3772_ = new_E3787_ | new_E3786_;
  assign new_E3773_ = new_E3782_ & new_E3785_;
  assign new_E3774_ = new_E3757_ | new_E3790_;
  assign new_E3775_ = new_E3789_ | new_E3788_;
  assign new_E3776_ = new_E3792_ | new_E3791_;
  assign new_E3777_ = ~new_E3768_ & new_E3794_;
  assign new_E3778_ = ~new_E3770_ & new_E3782_;
  assign new_E3779_ = new_E3770_ & ~new_E3782_;
  assign new_E3780_ = new_E3756_ & ~new_E3757_;
  assign new_E3781_ = ~new_E3803_ | ~new_E3804_;
  assign new_E3782_ = new_E3796_ | new_E3798_;
  assign new_E3783_ = new_E3806_ | new_E3805_;
  assign new_E3784_ = new_E3800_ | new_E3799_;
  assign new_E3785_ = ~new_E3808_ | ~new_E3807_;
  assign new_E3786_ = ~new_E3809_ & new_E3810_;
  assign new_E3787_ = new_E3809_ & ~new_E3810_;
  assign new_E3788_ = ~new_E3756_ & new_E3757_;
  assign new_E3789_ = new_E3756_ & ~new_E3757_;
  assign new_E3790_ = ~new_E3772_ | new_E3782_;
  assign new_E3791_ = new_E3772_ & new_E3782_;
  assign new_E3792_ = ~new_E3772_ & ~new_E3782_;
  assign new_E3793_ = new_E3814_ | new_E3813_;
  assign new_E3794_ = new_E3760_ | new_E3793_;
  assign new_E3795_ = new_E3818_ | new_E3817_;
  assign new_E3796_ = ~new_E3760_ & new_E3795_;
  assign new_E3797_ = new_E3816_ | new_E3815_;
  assign new_E3798_ = new_E3760_ & new_E3797_;
  assign new_E3799_ = new_E3758_ & ~new_E3768_;
  assign new_E3800_ = ~new_E3758_ & new_E3768_;
  assign new_E3801_ = ~new_E3757_ | ~new_E3782_;
  assign new_E3802_ = new_E3768_ & new_E3801_;
  assign new_E3803_ = ~new_E3768_ & ~new_E3802_;
  assign new_E3804_ = new_E3768_ | new_E3801_;
  assign new_E3805_ = ~new_E3758_ & new_E3759_;
  assign new_E3806_ = new_E3758_ & ~new_E3759_;
  assign new_E3807_ = new_E3775_ | new_E3812_;
  assign new_E3808_ = ~new_E3775_ & ~new_E3811_;
  assign new_E3809_ = new_E3758_ | new_E3775_;
  assign new_E3810_ = new_E3758_ | new_E3759_;
  assign new_E3811_ = new_E3775_ & new_E3812_;
  assign new_E3812_ = ~new_E3757_ | ~new_E3782_;
  assign new_E3813_ = new_E3790_ & new_E3810_;
  assign new_E3814_ = ~new_E3790_ & ~new_E3810_;
  assign new_E3815_ = new_E3819_ | new_E3820_;
  assign new_E3816_ = ~new_E3761_ & new_E3775_;
  assign new_E3817_ = new_E3821_ | new_E3822_;
  assign new_E3818_ = new_E3761_ & new_E3775_;
  assign new_E3819_ = ~new_E3761_ & ~new_E3775_;
  assign new_E3820_ = new_E3761_ & ~new_E3775_;
  assign new_E3821_ = new_E3761_ & ~new_E3775_;
  assign new_E3822_ = ~new_E3761_ & new_E3775_;
  assign new_E3823_ = new_G3531_;
  assign new_E3824_ = new_G3598_;
  assign new_E3825_ = new_G3665_;
  assign new_E3826_ = new_G3732_;
  assign new_E3827_ = new_G3799_;
  assign new_E3828_ = new_G3866_;
  assign new_E3829_ = new_E3836_ & new_E3835_;
  assign new_E3830_ = new_E3838_ | new_E3837_;
  assign new_E3831_ = new_E3840_ | new_E3839_;
  assign new_E3832_ = new_E3842_ & new_E3841_;
  assign new_E3833_ = new_E3842_ & new_E3843_;
  assign new_E3834_ = new_E3835_ | new_E3844_;
  assign new_E3835_ = new_E3824_ | new_E3847_;
  assign new_E3836_ = new_E3846_ | new_E3845_;
  assign new_E3837_ = new_E3851_ & new_E3850_;
  assign new_E3838_ = new_E3849_ & new_E3848_;
  assign new_E3839_ = new_E3854_ | new_E3853_;
  assign new_E3840_ = new_E3849_ & new_E3852_;
  assign new_E3841_ = new_E3824_ | new_E3857_;
  assign new_E3842_ = new_E3856_ | new_E3855_;
  assign new_E3843_ = new_E3859_ | new_E3858_;
  assign new_E3844_ = ~new_E3835_ & new_E3861_;
  assign new_E3845_ = ~new_E3837_ & new_E3849_;
  assign new_E3846_ = new_E3837_ & ~new_E3849_;
  assign new_E3847_ = new_E3823_ & ~new_E3824_;
  assign new_E3848_ = ~new_E3870_ | ~new_E3871_;
  assign new_E3849_ = new_E3863_ | new_E3865_;
  assign new_E3850_ = new_E3873_ | new_E3872_;
  assign new_E3851_ = new_E3867_ | new_E3866_;
  assign new_E3852_ = ~new_E3875_ | ~new_E3874_;
  assign new_E3853_ = ~new_E3876_ & new_E3877_;
  assign new_E3854_ = new_E3876_ & ~new_E3877_;
  assign new_E3855_ = ~new_E3823_ & new_E3824_;
  assign new_E3856_ = new_E3823_ & ~new_E3824_;
  assign new_E3857_ = ~new_E3839_ | new_E3849_;
  assign new_E3858_ = new_E3839_ & new_E3849_;
  assign new_E3859_ = ~new_E3839_ & ~new_E3849_;
  assign new_E3860_ = new_E3881_ | new_E3880_;
  assign new_E3861_ = new_E3827_ | new_E3860_;
  assign new_E3862_ = new_E3885_ | new_E3884_;
  assign new_E3863_ = ~new_E3827_ & new_E3862_;
  assign new_E3864_ = new_E3883_ | new_E3882_;
  assign new_E3865_ = new_E3827_ & new_E3864_;
  assign new_E3866_ = new_E3825_ & ~new_E3835_;
  assign new_E3867_ = ~new_E3825_ & new_E3835_;
  assign new_E3868_ = ~new_E3824_ | ~new_E3849_;
  assign new_E3869_ = new_E3835_ & new_E3868_;
  assign new_E3870_ = ~new_E3835_ & ~new_E3869_;
  assign new_E3871_ = new_E3835_ | new_E3868_;
  assign new_E3872_ = ~new_E3825_ & new_E3826_;
  assign new_E3873_ = new_E3825_ & ~new_E3826_;
  assign new_E3874_ = new_E3842_ | new_E3879_;
  assign new_E3875_ = ~new_E3842_ & ~new_E3878_;
  assign new_E3876_ = new_E3825_ | new_E3842_;
  assign new_E3877_ = new_E3825_ | new_E3826_;
  assign new_E3878_ = new_E3842_ & new_E3879_;
  assign new_E3879_ = ~new_E3824_ | ~new_E3849_;
  assign new_E3880_ = new_E3857_ & new_E3877_;
  assign new_E3881_ = ~new_E3857_ & ~new_E3877_;
  assign new_E3882_ = new_E3886_ | new_E3887_;
  assign new_E3883_ = ~new_E3828_ & new_E3842_;
  assign new_E3884_ = new_E3888_ | new_E3889_;
  assign new_E3885_ = new_E3828_ & new_E3842_;
  assign new_E3886_ = ~new_E3828_ & ~new_E3842_;
  assign new_E3887_ = new_E3828_ & ~new_E3842_;
  assign new_E3888_ = new_E3828_ & ~new_E3842_;
  assign new_E3889_ = ~new_E3828_ & new_E3842_;
  assign new_E3890_ = new_G3933_;
  assign new_E3891_ = new_G4000_;
  assign new_E3892_ = new_G4067_;
  assign new_E3893_ = new_G4134_;
  assign new_E3894_ = new_G4201_;
  assign new_E3895_ = new_G4268_;
  assign new_E3896_ = new_E3903_ & new_E3902_;
  assign new_E3897_ = new_E3905_ | new_E3904_;
  assign new_E3898_ = new_E3907_ | new_E3906_;
  assign new_E3899_ = new_E3909_ & new_E3908_;
  assign new_E3900_ = new_E3909_ & new_E3910_;
  assign new_E3901_ = new_E3902_ | new_E3911_;
  assign new_E3902_ = new_E3891_ | new_E3914_;
  assign new_E3903_ = new_E3913_ | new_E3912_;
  assign new_E3904_ = new_E3918_ & new_E3917_;
  assign new_E3905_ = new_E3916_ & new_E3915_;
  assign new_E3906_ = new_E3921_ | new_E3920_;
  assign new_E3907_ = new_E3916_ & new_E3919_;
  assign new_E3908_ = new_E3891_ | new_E3924_;
  assign new_E3909_ = new_E3923_ | new_E3922_;
  assign new_E3910_ = new_E3926_ | new_E3925_;
  assign new_E3911_ = ~new_E3902_ & new_E3928_;
  assign new_E3912_ = ~new_E3904_ & new_E3916_;
  assign new_E3913_ = new_E3904_ & ~new_E3916_;
  assign new_E3914_ = new_E3890_ & ~new_E3891_;
  assign new_E3915_ = ~new_E3937_ | ~new_E3938_;
  assign new_E3916_ = new_E3930_ | new_E3932_;
  assign new_E3917_ = new_E3940_ | new_E3939_;
  assign new_E3918_ = new_E3934_ | new_E3933_;
  assign new_E3919_ = ~new_E3942_ | ~new_E3941_;
  assign new_E3920_ = ~new_E3943_ & new_E3944_;
  assign new_E3921_ = new_E3943_ & ~new_E3944_;
  assign new_E3922_ = ~new_E3890_ & new_E3891_;
  assign new_E3923_ = new_E3890_ & ~new_E3891_;
  assign new_E3924_ = ~new_E3906_ | new_E3916_;
  assign new_E3925_ = new_E3906_ & new_E3916_;
  assign new_E3926_ = ~new_E3906_ & ~new_E3916_;
  assign new_E3927_ = new_E3948_ | new_E3947_;
  assign new_E3928_ = new_E3894_ | new_E3927_;
  assign new_E3929_ = new_E3952_ | new_E3951_;
  assign new_E3930_ = ~new_E3894_ & new_E3929_;
  assign new_E3931_ = new_E3950_ | new_E3949_;
  assign new_E3932_ = new_E3894_ & new_E3931_;
  assign new_E3933_ = new_E3892_ & ~new_E3902_;
  assign new_E3934_ = ~new_E3892_ & new_E3902_;
  assign new_E3935_ = ~new_E3891_ | ~new_E3916_;
  assign new_E3936_ = new_E3902_ & new_E3935_;
  assign new_E3937_ = ~new_E3902_ & ~new_E3936_;
  assign new_E3938_ = new_E3902_ | new_E3935_;
  assign new_E3939_ = ~new_E3892_ & new_E3893_;
  assign new_E3940_ = new_E3892_ & ~new_E3893_;
  assign new_E3941_ = new_E3909_ | new_E3946_;
  assign new_E3942_ = ~new_E3909_ & ~new_E3945_;
  assign new_E3943_ = new_E3892_ | new_E3909_;
  assign new_E3944_ = new_E3892_ | new_E3893_;
  assign new_E3945_ = new_E3909_ & new_E3946_;
  assign new_E3946_ = ~new_E3891_ | ~new_E3916_;
  assign new_E3947_ = new_E3924_ & new_E3944_;
  assign new_E3948_ = ~new_E3924_ & ~new_E3944_;
  assign new_E3949_ = new_E3953_ | new_E3954_;
  assign new_E3950_ = ~new_E3895_ & new_E3909_;
  assign new_E3951_ = new_E3955_ | new_E3956_;
  assign new_E3952_ = new_E3895_ & new_E3909_;
  assign new_E3953_ = ~new_E3895_ & ~new_E3909_;
  assign new_E3954_ = new_E3895_ & ~new_E3909_;
  assign new_E3955_ = new_E3895_ & ~new_E3909_;
  assign new_E3956_ = ~new_E3895_ & new_E3909_;
  assign new_E3957_ = new_G4335_;
  assign new_E3958_ = new_G4402_;
  assign new_E3959_ = new_G4469_;
  assign new_E3960_ = new_G4536_;
  assign new_E3961_ = new_G4603_;
  assign new_E3962_ = new_G4670_;
  assign new_E3963_ = new_E3970_ & new_E3969_;
  assign new_E3964_ = new_E3972_ | new_E3971_;
  assign new_E3965_ = new_E3974_ | new_E3973_;
  assign new_E3966_ = new_E3976_ & new_E3975_;
  assign new_E3967_ = new_E3976_ & new_E3977_;
  assign new_E3968_ = new_E3969_ | new_E3978_;
  assign new_E3969_ = new_E3958_ | new_E3981_;
  assign new_E3970_ = new_E3980_ | new_E3979_;
  assign new_E3971_ = new_E3985_ & new_E3984_;
  assign new_E3972_ = new_E3983_ & new_E3982_;
  assign new_E3973_ = new_E3988_ | new_E3987_;
  assign new_E3974_ = new_E3983_ & new_E3986_;
  assign new_E3975_ = new_E3958_ | new_E3991_;
  assign new_E3976_ = new_E3990_ | new_E3989_;
  assign new_E3977_ = new_E3993_ | new_E3992_;
  assign new_E3978_ = ~new_E3969_ & new_E3995_;
  assign new_E3979_ = ~new_E3971_ & new_E3983_;
  assign new_E3980_ = new_E3971_ & ~new_E3983_;
  assign new_E3981_ = new_E3957_ & ~new_E3958_;
  assign new_E3982_ = ~new_E4004_ | ~new_E4005_;
  assign new_E3983_ = new_E3997_ | new_E3999_;
  assign new_E3984_ = new_E4007_ | new_E4006_;
  assign new_E3985_ = new_E4001_ | new_E4000_;
  assign new_E3986_ = ~new_E4009_ | ~new_E4008_;
  assign new_E3987_ = ~new_E4010_ & new_E4011_;
  assign new_E3988_ = new_E4010_ & ~new_E4011_;
  assign new_E3989_ = ~new_E3957_ & new_E3958_;
  assign new_E3990_ = new_E3957_ & ~new_E3958_;
  assign new_E3991_ = ~new_E3973_ | new_E3983_;
  assign new_E3992_ = new_E3973_ & new_E3983_;
  assign new_E3993_ = ~new_E3973_ & ~new_E3983_;
  assign new_E3994_ = new_E4015_ | new_E4014_;
  assign new_E3995_ = new_E3961_ | new_E3994_;
  assign new_E3996_ = new_E4019_ | new_E4018_;
  assign new_E3997_ = ~new_E3961_ & new_E3996_;
  assign new_E3998_ = new_E4017_ | new_E4016_;
  assign new_E3999_ = new_E3961_ & new_E3998_;
  assign new_E4000_ = new_E3959_ & ~new_E3969_;
  assign new_E4001_ = ~new_E3959_ & new_E3969_;
  assign new_E4002_ = ~new_E3958_ | ~new_E3983_;
  assign new_E4003_ = new_E3969_ & new_E4002_;
  assign new_E4004_ = ~new_E3969_ & ~new_E4003_;
  assign new_E4005_ = new_E3969_ | new_E4002_;
  assign new_E4006_ = ~new_E3959_ & new_E3960_;
  assign new_E4007_ = new_E3959_ & ~new_E3960_;
  assign new_E4008_ = new_E3976_ | new_E4013_;
  assign new_E4009_ = ~new_E3976_ & ~new_E4012_;
  assign new_E4010_ = new_E3959_ | new_E3976_;
  assign new_E4011_ = new_E3959_ | new_E3960_;
  assign new_E4012_ = new_E3976_ & new_E4013_;
  assign new_E4013_ = ~new_E3958_ | ~new_E3983_;
  assign new_E4014_ = new_E3991_ & new_E4011_;
  assign new_E4015_ = ~new_E3991_ & ~new_E4011_;
  assign new_E4016_ = new_E4020_ | new_E4021_;
  assign new_E4017_ = ~new_E3962_ & new_E3976_;
  assign new_E4018_ = new_E4022_ | new_E4023_;
  assign new_E4019_ = new_E3962_ & new_E3976_;
  assign new_E4020_ = ~new_E3962_ & ~new_E3976_;
  assign new_E4021_ = new_E3962_ & ~new_E3976_;
  assign new_E4022_ = new_E3962_ & ~new_E3976_;
  assign new_E4023_ = ~new_E3962_ & new_E3976_;
  assign new_E4024_ = new_G4737_;
  assign new_E4025_ = new_G4804_;
  assign new_E4026_ = new_G4871_;
  assign new_E4027_ = new_G4938_;
  assign new_E4028_ = new_G5005_;
  assign new_E4029_ = new_G5072_;
  assign new_E4030_ = new_E4037_ & new_E4036_;
  assign new_E4031_ = new_E4039_ | new_E4038_;
  assign new_E4032_ = new_E4041_ | new_E4040_;
  assign new_E4033_ = new_E4043_ & new_E4042_;
  assign new_E4034_ = new_E4043_ & new_E4044_;
  assign new_E4035_ = new_E4036_ | new_E4045_;
  assign new_E4036_ = new_E4025_ | new_E4048_;
  assign new_E4037_ = new_E4047_ | new_E4046_;
  assign new_E4038_ = new_E4052_ & new_E4051_;
  assign new_E4039_ = new_E4050_ & new_E4049_;
  assign new_E4040_ = new_E4055_ | new_E4054_;
  assign new_E4041_ = new_E4050_ & new_E4053_;
  assign new_E4042_ = new_E4025_ | new_E4058_;
  assign new_E4043_ = new_E4057_ | new_E4056_;
  assign new_E4044_ = new_E4060_ | new_E4059_;
  assign new_E4045_ = ~new_E4036_ & new_E4062_;
  assign new_E4046_ = ~new_E4038_ & new_E4050_;
  assign new_E4047_ = new_E4038_ & ~new_E4050_;
  assign new_E4048_ = new_E4024_ & ~new_E4025_;
  assign new_E4049_ = ~new_E4071_ | ~new_E4072_;
  assign new_E4050_ = new_E4064_ | new_E4066_;
  assign new_E4051_ = new_E4074_ | new_E4073_;
  assign new_E4052_ = new_E4068_ | new_E4067_;
  assign new_E4053_ = ~new_E4076_ | ~new_E4075_;
  assign new_E4054_ = ~new_E4077_ & new_E4078_;
  assign new_E4055_ = new_E4077_ & ~new_E4078_;
  assign new_E4056_ = ~new_E4024_ & new_E4025_;
  assign new_E4057_ = new_E4024_ & ~new_E4025_;
  assign new_E4058_ = ~new_E4040_ | new_E4050_;
  assign new_E4059_ = new_E4040_ & new_E4050_;
  assign new_E4060_ = ~new_E4040_ & ~new_E4050_;
  assign new_E4061_ = new_E4082_ | new_E4081_;
  assign new_E4062_ = new_E4028_ | new_E4061_;
  assign new_E4063_ = new_E4086_ | new_E4085_;
  assign new_E4064_ = ~new_E4028_ & new_E4063_;
  assign new_E4065_ = new_E4084_ | new_E4083_;
  assign new_E4066_ = new_E4028_ & new_E4065_;
  assign new_E4067_ = new_E4026_ & ~new_E4036_;
  assign new_E4068_ = ~new_E4026_ & new_E4036_;
  assign new_E4069_ = ~new_E4025_ | ~new_E4050_;
  assign new_E4070_ = new_E4036_ & new_E4069_;
  assign new_E4071_ = ~new_E4036_ & ~new_E4070_;
  assign new_E4072_ = new_E4036_ | new_E4069_;
  assign new_E4073_ = ~new_E4026_ & new_E4027_;
  assign new_E4074_ = new_E4026_ & ~new_E4027_;
  assign new_E4075_ = new_E4043_ | new_E4080_;
  assign new_E4076_ = ~new_E4043_ & ~new_E4079_;
  assign new_E4077_ = new_E4026_ | new_E4043_;
  assign new_E4078_ = new_E4026_ | new_E4027_;
  assign new_E4079_ = new_E4043_ & new_E4080_;
  assign new_E4080_ = ~new_E4025_ | ~new_E4050_;
  assign new_E4081_ = new_E4058_ & new_E4078_;
  assign new_E4082_ = ~new_E4058_ & ~new_E4078_;
  assign new_E4083_ = new_E4087_ | new_E4088_;
  assign new_E4084_ = ~new_E4029_ & new_E4043_;
  assign new_E4085_ = new_E4089_ | new_E4090_;
  assign new_E4086_ = new_E4029_ & new_E4043_;
  assign new_E4087_ = ~new_E4029_ & ~new_E4043_;
  assign new_E4088_ = new_E4029_ & ~new_E4043_;
  assign new_E4089_ = new_E4029_ & ~new_E4043_;
  assign new_E4090_ = ~new_E4029_ & new_E4043_;
  assign new_E4091_ = new_G5139_;
  assign new_E4092_ = new_G5206_;
  assign new_E4093_ = new_G5273_;
  assign new_E4094_ = new_G5340_;
  assign new_E4095_ = new_G5407_;
  assign new_E4096_ = new_G5474_;
  assign new_E4097_ = new_E4104_ & new_E4103_;
  assign new_E4098_ = new_E4106_ | new_E4105_;
  assign new_E4099_ = new_E4108_ | new_E4107_;
  assign new_E4100_ = new_E4110_ & new_E4109_;
  assign new_E4101_ = new_E4110_ & new_E4111_;
  assign new_E4102_ = new_E4103_ | new_E4112_;
  assign new_E4103_ = new_E4092_ | new_E4115_;
  assign new_E4104_ = new_E4114_ | new_E4113_;
  assign new_E4105_ = new_E4119_ & new_E4118_;
  assign new_E4106_ = new_E4117_ & new_E4116_;
  assign new_E4107_ = new_E4122_ | new_E4121_;
  assign new_E4108_ = new_E4117_ & new_E4120_;
  assign new_E4109_ = new_E4092_ | new_E4125_;
  assign new_E4110_ = new_E4124_ | new_E4123_;
  assign new_E4111_ = new_E4127_ | new_E4126_;
  assign new_E4112_ = ~new_E4103_ & new_E4129_;
  assign new_E4113_ = ~new_E4105_ & new_E4117_;
  assign new_E4114_ = new_E4105_ & ~new_E4117_;
  assign new_E4115_ = new_E4091_ & ~new_E4092_;
  assign new_E4116_ = ~new_E4138_ | ~new_E4139_;
  assign new_E4117_ = new_E4131_ | new_E4133_;
  assign new_E4118_ = new_E4141_ | new_E4140_;
  assign new_E4119_ = new_E4135_ | new_E4134_;
  assign new_E4120_ = ~new_E4143_ | ~new_E4142_;
  assign new_E4121_ = ~new_E4144_ & new_E4145_;
  assign new_E4122_ = new_E4144_ & ~new_E4145_;
  assign new_E4123_ = ~new_E4091_ & new_E4092_;
  assign new_E4124_ = new_E4091_ & ~new_E4092_;
  assign new_E4125_ = ~new_E4107_ | new_E4117_;
  assign new_E4126_ = new_E4107_ & new_E4117_;
  assign new_E4127_ = ~new_E4107_ & ~new_E4117_;
  assign new_E4128_ = new_E4149_ | new_E4148_;
  assign new_E4129_ = new_E4095_ | new_E4128_;
  assign new_E4130_ = new_E4153_ | new_E4152_;
  assign new_E4131_ = ~new_E4095_ & new_E4130_;
  assign new_E4132_ = new_E4151_ | new_E4150_;
  assign new_E4133_ = new_E4095_ & new_E4132_;
  assign new_E4134_ = new_E4093_ & ~new_E4103_;
  assign new_E4135_ = ~new_E4093_ & new_E4103_;
  assign new_E4136_ = ~new_E4092_ | ~new_E4117_;
  assign new_E4137_ = new_E4103_ & new_E4136_;
  assign new_E4138_ = ~new_E4103_ & ~new_E4137_;
  assign new_E4139_ = new_E4103_ | new_E4136_;
  assign new_E4140_ = ~new_E4093_ & new_E4094_;
  assign new_E4141_ = new_E4093_ & ~new_E4094_;
  assign new_E4142_ = new_E4110_ | new_E4147_;
  assign new_E4143_ = ~new_E4110_ & ~new_E4146_;
  assign new_E4144_ = new_E4093_ | new_E4110_;
  assign new_E4145_ = new_E4093_ | new_E4094_;
  assign new_E4146_ = new_E4110_ & new_E4147_;
  assign new_E4147_ = ~new_E4092_ | ~new_E4117_;
  assign new_E4148_ = new_E4125_ & new_E4145_;
  assign new_E4149_ = ~new_E4125_ & ~new_E4145_;
  assign new_E4150_ = new_E4154_ | new_E4155_;
  assign new_E4151_ = ~new_E4096_ & new_E4110_;
  assign new_E4152_ = new_E4156_ | new_E4157_;
  assign new_E4153_ = new_E4096_ & new_E4110_;
  assign new_E4154_ = ~new_E4096_ & ~new_E4110_;
  assign new_E4155_ = new_E4096_ & ~new_E4110_;
  assign new_E4156_ = new_E4096_ & ~new_E4110_;
  assign new_E4157_ = ~new_E4096_ & new_E4110_;
  assign new_E4158_ = new_G5541_;
  assign new_E4159_ = new_G5608_;
  assign new_E4160_ = new_G5675_;
  assign new_E4161_ = new_G5742_;
  assign new_E4162_ = new_G5809_;
  assign new_E4163_ = new_G5876_;
  assign new_E4164_ = new_E4171_ & new_E4170_;
  assign new_E4165_ = new_E4173_ | new_E4172_;
  assign new_E4166_ = new_E4175_ | new_E4174_;
  assign new_E4167_ = new_E4177_ & new_E4176_;
  assign new_E4168_ = new_E4177_ & new_E4178_;
  assign new_E4169_ = new_E4170_ | new_E4179_;
  assign new_E4170_ = new_E4159_ | new_E4182_;
  assign new_E4171_ = new_E4181_ | new_E4180_;
  assign new_E4172_ = new_E4186_ & new_E4185_;
  assign new_E4173_ = new_E4184_ & new_E4183_;
  assign new_E4174_ = new_E4189_ | new_E4188_;
  assign new_E4175_ = new_E4184_ & new_E4187_;
  assign new_E4176_ = new_E4159_ | new_E4192_;
  assign new_E4177_ = new_E4191_ | new_E4190_;
  assign new_E4178_ = new_E4194_ | new_E4193_;
  assign new_E4179_ = ~new_E4170_ & new_E4196_;
  assign new_E4180_ = ~new_E4172_ & new_E4184_;
  assign new_E4181_ = new_E4172_ & ~new_E4184_;
  assign new_E4182_ = new_E4158_ & ~new_E4159_;
  assign new_E4183_ = ~new_E4205_ | ~new_E4206_;
  assign new_E4184_ = new_E4198_ | new_E4200_;
  assign new_E4185_ = new_E4208_ | new_E4207_;
  assign new_E4186_ = new_E4202_ | new_E4201_;
  assign new_E4187_ = ~new_E4210_ | ~new_E4209_;
  assign new_E4188_ = ~new_E4211_ & new_E4212_;
  assign new_E4189_ = new_E4211_ & ~new_E4212_;
  assign new_E4190_ = ~new_E4158_ & new_E4159_;
  assign new_E4191_ = new_E4158_ & ~new_E4159_;
  assign new_E4192_ = ~new_E4174_ | new_E4184_;
  assign new_E4193_ = new_E4174_ & new_E4184_;
  assign new_E4194_ = ~new_E4174_ & ~new_E4184_;
  assign new_E4195_ = new_E4216_ | new_E4215_;
  assign new_E4196_ = new_E4162_ | new_E4195_;
  assign new_E4197_ = new_E4220_ | new_E4219_;
  assign new_E4198_ = ~new_E4162_ & new_E4197_;
  assign new_E4199_ = new_E4218_ | new_E4217_;
  assign new_E4200_ = new_E4162_ & new_E4199_;
  assign new_E4201_ = new_E4160_ & ~new_E4170_;
  assign new_E4202_ = ~new_E4160_ & new_E4170_;
  assign new_E4203_ = ~new_E4159_ | ~new_E4184_;
  assign new_E4204_ = new_E4170_ & new_E4203_;
  assign new_E4205_ = ~new_E4170_ & ~new_E4204_;
  assign new_E4206_ = new_E4170_ | new_E4203_;
  assign new_E4207_ = ~new_E4160_ & new_E4161_;
  assign new_E4208_ = new_E4160_ & ~new_E4161_;
  assign new_E4209_ = new_E4177_ | new_E4214_;
  assign new_E4210_ = ~new_E4177_ & ~new_E4213_;
  assign new_E4211_ = new_E4160_ | new_E4177_;
  assign new_E4212_ = new_E4160_ | new_E4161_;
  assign new_E4213_ = new_E4177_ & new_E4214_;
  assign new_E4214_ = ~new_E4159_ | ~new_E4184_;
  assign new_E4215_ = new_E4192_ & new_E4212_;
  assign new_E4216_ = ~new_E4192_ & ~new_E4212_;
  assign new_E4217_ = new_E4221_ | new_E4222_;
  assign new_E4218_ = ~new_E4163_ & new_E4177_;
  assign new_E4219_ = new_E4223_ | new_E4224_;
  assign new_E4220_ = new_E4163_ & new_E4177_;
  assign new_E4221_ = ~new_E4163_ & ~new_E4177_;
  assign new_E4222_ = new_E4163_ & ~new_E4177_;
  assign new_E4223_ = new_E4163_ & ~new_E4177_;
  assign new_E4224_ = ~new_E4163_ & new_E4177_;
  assign new_E4225_ = new_F1470_;
  assign new_E4226_ = new_F1538_;
  assign new_E4227_ = new_F1605_;
  assign new_E4228_ = new_F1672_;
  assign new_E4229_ = new_F1739_;
  assign new_E4230_ = new_F1806_;
  assign new_E4231_ = new_E4238_ & new_E4237_;
  assign new_E4232_ = new_E4240_ | new_E4239_;
  assign new_E4233_ = new_E4242_ | new_E4241_;
  assign new_E4234_ = new_E4244_ & new_E4243_;
  assign new_E4235_ = new_E4244_ & new_E4245_;
  assign new_E4236_ = new_E4237_ | new_E4246_;
  assign new_E4237_ = new_E4226_ | new_E4249_;
  assign new_E4238_ = new_E4248_ | new_E4247_;
  assign new_E4239_ = new_E4253_ & new_E4252_;
  assign new_E4240_ = new_E4251_ & new_E4250_;
  assign new_E4241_ = new_E4256_ | new_E4255_;
  assign new_E4242_ = new_E4251_ & new_E4254_;
  assign new_E4243_ = new_E4226_ | new_E4259_;
  assign new_E4244_ = new_E4258_ | new_E4257_;
  assign new_E4245_ = new_E4261_ | new_E4260_;
  assign new_E4246_ = ~new_E4237_ & new_E4263_;
  assign new_E4247_ = ~new_E4239_ & new_E4251_;
  assign new_E4248_ = new_E4239_ & ~new_E4251_;
  assign new_E4249_ = new_E4225_ & ~new_E4226_;
  assign new_E4250_ = ~new_E4272_ | ~new_E4273_;
  assign new_E4251_ = new_E4265_ | new_E4267_;
  assign new_E4252_ = new_E4275_ | new_E4274_;
  assign new_E4253_ = new_E4269_ | new_E4268_;
  assign new_E4254_ = ~new_E4277_ | ~new_E4276_;
  assign new_E4255_ = ~new_E4278_ & new_E4279_;
  assign new_E4256_ = new_E4278_ & ~new_E4279_;
  assign new_E4257_ = ~new_E4225_ & new_E4226_;
  assign new_E4258_ = new_E4225_ & ~new_E4226_;
  assign new_E4259_ = ~new_E4241_ | new_E4251_;
  assign new_E4260_ = new_E4241_ & new_E4251_;
  assign new_E4261_ = ~new_E4241_ & ~new_E4251_;
  assign new_E4262_ = new_E4283_ | new_E4282_;
  assign new_E4263_ = new_E4229_ | new_E4262_;
  assign new_E4264_ = new_E4287_ | new_E4286_;
  assign new_E4265_ = ~new_E4229_ & new_E4264_;
  assign new_E4266_ = new_E4285_ | new_E4284_;
  assign new_E4267_ = new_E4229_ & new_E4266_;
  assign new_E4268_ = new_E4227_ & ~new_E4237_;
  assign new_E4269_ = ~new_E4227_ & new_E4237_;
  assign new_E4270_ = ~new_E4226_ | ~new_E4251_;
  assign new_E4271_ = new_E4237_ & new_E4270_;
  assign new_E4272_ = ~new_E4237_ & ~new_E4271_;
  assign new_E4273_ = new_E4237_ | new_E4270_;
  assign new_E4274_ = ~new_E4227_ & new_E4228_;
  assign new_E4275_ = new_E4227_ & ~new_E4228_;
  assign new_E4276_ = new_E4244_ | new_E4281_;
  assign new_E4277_ = ~new_E4244_ & ~new_E4280_;
  assign new_E4278_ = new_E4227_ | new_E4244_;
  assign new_E4279_ = new_E4227_ | new_E4228_;
  assign new_E4280_ = new_E4244_ & new_E4281_;
  assign new_E4281_ = ~new_E4226_ | ~new_E4251_;
  assign new_E4282_ = new_E4259_ & new_E4279_;
  assign new_E4283_ = ~new_E4259_ & ~new_E4279_;
  assign new_E4284_ = new_E4288_ | new_E4289_;
  assign new_E4285_ = ~new_E4230_ & new_E4244_;
  assign new_E4286_ = new_E4290_ | new_E4291_;
  assign new_E4287_ = new_E4230_ & new_E4244_;
  assign new_E4288_ = ~new_E4230_ & ~new_E4244_;
  assign new_E4289_ = new_E4230_ & ~new_E4244_;
  assign new_E4290_ = new_E4230_ & ~new_E4244_;
  assign new_E4291_ = ~new_E4230_ & new_E4244_;
  assign new_E4292_ = new_F1873_;
  assign new_E4293_ = new_F1940_;
  assign new_E4294_ = new_F2007_;
  assign new_E4295_ = new_F2074_;
  assign new_E4296_ = new_F2141_;
  assign new_E4297_ = new_F2208_;
  assign new_E4298_ = new_E4305_ & new_E4304_;
  assign new_E4299_ = new_E4307_ | new_E4306_;
  assign new_E4300_ = new_E4309_ | new_E4308_;
  assign new_E4301_ = new_E4311_ & new_E4310_;
  assign new_E4302_ = new_E4311_ & new_E4312_;
  assign new_E4303_ = new_E4304_ | new_E4313_;
  assign new_E4304_ = new_E4293_ | new_E4316_;
  assign new_E4305_ = new_E4315_ | new_E4314_;
  assign new_E4306_ = new_E4320_ & new_E4319_;
  assign new_E4307_ = new_E4318_ & new_E4317_;
  assign new_E4308_ = new_E4323_ | new_E4322_;
  assign new_E4309_ = new_E4318_ & new_E4321_;
  assign new_E4310_ = new_E4293_ | new_E4326_;
  assign new_E4311_ = new_E4325_ | new_E4324_;
  assign new_E4312_ = new_E4328_ | new_E4327_;
  assign new_E4313_ = ~new_E4304_ & new_E4330_;
  assign new_E4314_ = ~new_E4306_ & new_E4318_;
  assign new_E4315_ = new_E4306_ & ~new_E4318_;
  assign new_E4316_ = new_E4292_ & ~new_E4293_;
  assign new_E4317_ = ~new_E4339_ | ~new_E4340_;
  assign new_E4318_ = new_E4332_ | new_E4334_;
  assign new_E4319_ = new_E4342_ | new_E4341_;
  assign new_E4320_ = new_E4336_ | new_E4335_;
  assign new_E4321_ = ~new_E4344_ | ~new_E4343_;
  assign new_E4322_ = ~new_E4345_ & new_E4346_;
  assign new_E4323_ = new_E4345_ & ~new_E4346_;
  assign new_E4324_ = ~new_E4292_ & new_E4293_;
  assign new_E4325_ = new_E4292_ & ~new_E4293_;
  assign new_E4326_ = ~new_E4308_ | new_E4318_;
  assign new_E4327_ = new_E4308_ & new_E4318_;
  assign new_E4328_ = ~new_E4308_ & ~new_E4318_;
  assign new_E4329_ = new_E4350_ | new_E4349_;
  assign new_E4330_ = new_E4296_ | new_E4329_;
  assign new_E4331_ = new_E4354_ | new_E4353_;
  assign new_E4332_ = ~new_E4296_ & new_E4331_;
  assign new_E4333_ = new_E4352_ | new_E4351_;
  assign new_E4334_ = new_E4296_ & new_E4333_;
  assign new_E4335_ = new_E4294_ & ~new_E4304_;
  assign new_E4336_ = ~new_E4294_ & new_E4304_;
  assign new_E4337_ = ~new_E4293_ | ~new_E4318_;
  assign new_E4338_ = new_E4304_ & new_E4337_;
  assign new_E4339_ = ~new_E4304_ & ~new_E4338_;
  assign new_E4340_ = new_E4304_ | new_E4337_;
  assign new_E4341_ = ~new_E4294_ & new_E4295_;
  assign new_E4342_ = new_E4294_ & ~new_E4295_;
  assign new_E4343_ = new_E4311_ | new_E4348_;
  assign new_E4344_ = ~new_E4311_ & ~new_E4347_;
  assign new_E4345_ = new_E4294_ | new_E4311_;
  assign new_E4346_ = new_E4294_ | new_E4295_;
  assign new_E4347_ = new_E4311_ & new_E4348_;
  assign new_E4348_ = ~new_E4293_ | ~new_E4318_;
  assign new_E4349_ = new_E4326_ & new_E4346_;
  assign new_E4350_ = ~new_E4326_ & ~new_E4346_;
  assign new_E4351_ = new_E4355_ | new_E4356_;
  assign new_E4352_ = ~new_E4297_ & new_E4311_;
  assign new_E4353_ = new_E4357_ | new_E4358_;
  assign new_E4354_ = new_E4297_ & new_E4311_;
  assign new_E4355_ = ~new_E4297_ & ~new_E4311_;
  assign new_E4356_ = new_E4297_ & ~new_E4311_;
  assign new_E4357_ = new_E4297_ & ~new_E4311_;
  assign new_E4358_ = ~new_E4297_ & new_E4311_;
  assign new_E4359_ = new_F2275_;
  assign new_E4360_ = new_F2342_;
  assign new_E4361_ = new_F2409_;
  assign new_E4362_ = new_F2476_;
  assign new_E4363_ = new_F2543_;
  assign new_E4364_ = new_F2610_;
  assign new_E4365_ = new_E4372_ & new_E4371_;
  assign new_E4366_ = new_E4374_ | new_E4373_;
  assign new_E4367_ = new_E4376_ | new_E4375_;
  assign new_E4368_ = new_E4378_ & new_E4377_;
  assign new_E4369_ = new_E4378_ & new_E4379_;
  assign new_E4370_ = new_E4371_ | new_E4380_;
  assign new_E4371_ = new_E4360_ | new_E4383_;
  assign new_E4372_ = new_E4382_ | new_E4381_;
  assign new_E4373_ = new_E4387_ & new_E4386_;
  assign new_E4374_ = new_E4385_ & new_E4384_;
  assign new_E4375_ = new_E4390_ | new_E4389_;
  assign new_E4376_ = new_E4385_ & new_E4388_;
  assign new_E4377_ = new_E4360_ | new_E4393_;
  assign new_E4378_ = new_E4392_ | new_E4391_;
  assign new_E4379_ = new_E4395_ | new_E4394_;
  assign new_E4380_ = ~new_E4371_ & new_E4397_;
  assign new_E4381_ = ~new_E4373_ & new_E4385_;
  assign new_E4382_ = new_E4373_ & ~new_E4385_;
  assign new_E4383_ = new_E4359_ & ~new_E4360_;
  assign new_E4384_ = ~new_E4406_ | ~new_E4407_;
  assign new_E4385_ = new_E4399_ | new_E4401_;
  assign new_E4386_ = new_E4409_ | new_E4408_;
  assign new_E4387_ = new_E4403_ | new_E4402_;
  assign new_E4388_ = ~new_E4411_ | ~new_E4410_;
  assign new_E4389_ = ~new_E4412_ & new_E4413_;
  assign new_E4390_ = new_E4412_ & ~new_E4413_;
  assign new_E4391_ = ~new_E4359_ & new_E4360_;
  assign new_E4392_ = new_E4359_ & ~new_E4360_;
  assign new_E4393_ = ~new_E4375_ | new_E4385_;
  assign new_E4394_ = new_E4375_ & new_E4385_;
  assign new_E4395_ = ~new_E4375_ & ~new_E4385_;
  assign new_E4396_ = new_E4417_ | new_E4416_;
  assign new_E4397_ = new_E4363_ | new_E4396_;
  assign new_E4398_ = new_E4421_ | new_E4420_;
  assign new_E4399_ = ~new_E4363_ & new_E4398_;
  assign new_E4400_ = new_E4419_ | new_E4418_;
  assign new_E4401_ = new_E4363_ & new_E4400_;
  assign new_E4402_ = new_E4361_ & ~new_E4371_;
  assign new_E4403_ = ~new_E4361_ & new_E4371_;
  assign new_E4404_ = ~new_E4360_ | ~new_E4385_;
  assign new_E4405_ = new_E4371_ & new_E4404_;
  assign new_E4406_ = ~new_E4371_ & ~new_E4405_;
  assign new_E4407_ = new_E4371_ | new_E4404_;
  assign new_E4408_ = ~new_E4361_ & new_E4362_;
  assign new_E4409_ = new_E4361_ & ~new_E4362_;
  assign new_E4410_ = new_E4378_ | new_E4415_;
  assign new_E4411_ = ~new_E4378_ & ~new_E4414_;
  assign new_E4412_ = new_E4361_ | new_E4378_;
  assign new_E4413_ = new_E4361_ | new_E4362_;
  assign new_E4414_ = new_E4378_ & new_E4415_;
  assign new_E4415_ = ~new_E4360_ | ~new_E4385_;
  assign new_E4416_ = new_E4393_ & new_E4413_;
  assign new_E4417_ = ~new_E4393_ & ~new_E4413_;
  assign new_E4418_ = new_E4422_ | new_E4423_;
  assign new_E4419_ = ~new_E4364_ & new_E4378_;
  assign new_E4420_ = new_E4424_ | new_E4425_;
  assign new_E4421_ = new_E4364_ & new_E4378_;
  assign new_E4422_ = ~new_E4364_ & ~new_E4378_;
  assign new_E4423_ = new_E4364_ & ~new_E4378_;
  assign new_E4424_ = new_E4364_ & ~new_E4378_;
  assign new_E4425_ = ~new_E4364_ & new_E4378_;
  assign new_E4426_ = new_F2677_;
  assign new_E4427_ = new_F2744_;
  assign new_E4428_ = new_F2811_;
  assign new_E4429_ = new_F2878_;
  assign new_E4430_ = new_F2945_;
  assign new_E4431_ = new_F3012_;
  assign new_E4432_ = new_E4439_ & new_E4438_;
  assign new_E4433_ = new_E4441_ | new_E4440_;
  assign new_E4434_ = new_E4443_ | new_E4442_;
  assign new_E4435_ = new_E4445_ & new_E4444_;
  assign new_E4436_ = new_E4445_ & new_E4446_;
  assign new_E4437_ = new_E4438_ | new_E4447_;
  assign new_E4438_ = new_E4427_ | new_E4450_;
  assign new_E4439_ = new_E4449_ | new_E4448_;
  assign new_E4440_ = new_E4454_ & new_E4453_;
  assign new_E4441_ = new_E4452_ & new_E4451_;
  assign new_E4442_ = new_E4457_ | new_E4456_;
  assign new_E4443_ = new_E4452_ & new_E4455_;
  assign new_E4444_ = new_E4427_ | new_E4460_;
  assign new_E4445_ = new_E4459_ | new_E4458_;
  assign new_E4446_ = new_E4462_ | new_E4461_;
  assign new_E4447_ = ~new_E4438_ & new_E4464_;
  assign new_E4448_ = ~new_E4440_ & new_E4452_;
  assign new_E4449_ = new_E4440_ & ~new_E4452_;
  assign new_E4450_ = new_E4426_ & ~new_E4427_;
  assign new_E4451_ = ~new_E4473_ | ~new_E4474_;
  assign new_E4452_ = new_E4466_ | new_E4468_;
  assign new_E4453_ = new_E4476_ | new_E4475_;
  assign new_E4454_ = new_E4470_ | new_E4469_;
  assign new_E4455_ = ~new_E4478_ | ~new_E4477_;
  assign new_E4456_ = ~new_E4479_ & new_E4480_;
  assign new_E4457_ = new_E4479_ & ~new_E4480_;
  assign new_E4458_ = ~new_E4426_ & new_E4427_;
  assign new_E4459_ = new_E4426_ & ~new_E4427_;
  assign new_E4460_ = ~new_E4442_ | new_E4452_;
  assign new_E4461_ = new_E4442_ & new_E4452_;
  assign new_E4462_ = ~new_E4442_ & ~new_E4452_;
  assign new_E4463_ = new_E4484_ | new_E4483_;
  assign new_E4464_ = new_E4430_ | new_E4463_;
  assign new_E4465_ = new_E4488_ | new_E4487_;
  assign new_E4466_ = ~new_E4430_ & new_E4465_;
  assign new_E4467_ = new_E4486_ | new_E4485_;
  assign new_E4468_ = new_E4430_ & new_E4467_;
  assign new_E4469_ = new_E4428_ & ~new_E4438_;
  assign new_E4470_ = ~new_E4428_ & new_E4438_;
  assign new_E4471_ = ~new_E4427_ | ~new_E4452_;
  assign new_E4472_ = new_E4438_ & new_E4471_;
  assign new_E4473_ = ~new_E4438_ & ~new_E4472_;
  assign new_E4474_ = new_E4438_ | new_E4471_;
  assign new_E4475_ = ~new_E4428_ & new_E4429_;
  assign new_E4476_ = new_E4428_ & ~new_E4429_;
  assign new_E4477_ = new_E4445_ | new_E4482_;
  assign new_E4478_ = ~new_E4445_ & ~new_E4481_;
  assign new_E4479_ = new_E4428_ | new_E4445_;
  assign new_E4480_ = new_E4428_ | new_E4429_;
  assign new_E4481_ = new_E4445_ & new_E4482_;
  assign new_E4482_ = ~new_E4427_ | ~new_E4452_;
  assign new_E4483_ = new_E4460_ & new_E4480_;
  assign new_E4484_ = ~new_E4460_ & ~new_E4480_;
  assign new_E4485_ = new_E4489_ | new_E4490_;
  assign new_E4486_ = ~new_E4431_ & new_E4445_;
  assign new_E4487_ = new_E4491_ | new_E4492_;
  assign new_E4488_ = new_E4431_ & new_E4445_;
  assign new_E4489_ = ~new_E4431_ & ~new_E4445_;
  assign new_E4490_ = new_E4431_ & ~new_E4445_;
  assign new_E4491_ = new_E4431_ & ~new_E4445_;
  assign new_E4492_ = ~new_E4431_ & new_E4445_;
  assign new_E4493_ = new_F3079_;
  assign new_E4494_ = new_F3146_;
  assign new_E4495_ = new_F3213_;
  assign new_E4496_ = new_F3280_;
  assign new_E4497_ = new_F3347_;
  assign new_E4498_ = new_F3414_;
  assign new_E4499_ = new_E4506_ & new_E4505_;
  assign new_E4500_ = new_E4508_ | new_E4507_;
  assign new_E4501_ = new_E4510_ | new_E4509_;
  assign new_E4502_ = new_E4512_ & new_E4511_;
  assign new_E4503_ = new_E4512_ & new_E4513_;
  assign new_E4504_ = new_E4505_ | new_E4514_;
  assign new_E4505_ = new_E4494_ | new_E4517_;
  assign new_E4506_ = new_E4516_ | new_E4515_;
  assign new_E4507_ = new_E4521_ & new_E4520_;
  assign new_E4508_ = new_E4519_ & new_E4518_;
  assign new_E4509_ = new_E4524_ | new_E4523_;
  assign new_E4510_ = new_E4519_ & new_E4522_;
  assign new_E4511_ = new_E4494_ | new_E4527_;
  assign new_E4512_ = new_E4526_ | new_E4525_;
  assign new_E4513_ = new_E4529_ | new_E4528_;
  assign new_E4514_ = ~new_E4505_ & new_E4531_;
  assign new_E4515_ = ~new_E4507_ & new_E4519_;
  assign new_E4516_ = new_E4507_ & ~new_E4519_;
  assign new_E4517_ = new_E4493_ & ~new_E4494_;
  assign new_E4518_ = ~new_E4540_ | ~new_E4541_;
  assign new_E4519_ = new_E4533_ | new_E4535_;
  assign new_E4520_ = new_E4543_ | new_E4542_;
  assign new_E4521_ = new_E4537_ | new_E4536_;
  assign new_E4522_ = ~new_E4545_ | ~new_E4544_;
  assign new_E4523_ = ~new_E4546_ & new_E4547_;
  assign new_E4524_ = new_E4546_ & ~new_E4547_;
  assign new_E4525_ = ~new_E4493_ & new_E4494_;
  assign new_E4526_ = new_E4493_ & ~new_E4494_;
  assign new_E4527_ = ~new_E4509_ | new_E4519_;
  assign new_E4528_ = new_E4509_ & new_E4519_;
  assign new_E4529_ = ~new_E4509_ & ~new_E4519_;
  assign new_E4530_ = new_E4551_ | new_E4550_;
  assign new_E4531_ = new_E4497_ | new_E4530_;
  assign new_E4532_ = new_E4555_ | new_E4554_;
  assign new_E4533_ = ~new_E4497_ & new_E4532_;
  assign new_E4534_ = new_E4553_ | new_E4552_;
  assign new_E4535_ = new_E4497_ & new_E4534_;
  assign new_E4536_ = new_E4495_ & ~new_E4505_;
  assign new_E4537_ = ~new_E4495_ & new_E4505_;
  assign new_E4538_ = ~new_E4494_ | ~new_E4519_;
  assign new_E4539_ = new_E4505_ & new_E4538_;
  assign new_E4540_ = ~new_E4505_ & ~new_E4539_;
  assign new_E4541_ = new_E4505_ | new_E4538_;
  assign new_E4542_ = ~new_E4495_ & new_E4496_;
  assign new_E4543_ = new_E4495_ & ~new_E4496_;
  assign new_E4544_ = new_E4512_ | new_E4549_;
  assign new_E4545_ = ~new_E4512_ & ~new_E4548_;
  assign new_E4546_ = new_E4495_ | new_E4512_;
  assign new_E4547_ = new_E4495_ | new_E4496_;
  assign new_E4548_ = new_E4512_ & new_E4549_;
  assign new_E4549_ = ~new_E4494_ | ~new_E4519_;
  assign new_E4550_ = new_E4527_ & new_E4547_;
  assign new_E4551_ = ~new_E4527_ & ~new_E4547_;
  assign new_E4552_ = new_E4556_ | new_E4557_;
  assign new_E4553_ = ~new_E4498_ & new_E4512_;
  assign new_E4554_ = new_E4558_ | new_E4559_;
  assign new_E4555_ = new_E4498_ & new_E4512_;
  assign new_E4556_ = ~new_E4498_ & ~new_E4512_;
  assign new_E4557_ = new_E4498_ & ~new_E4512_;
  assign new_E4558_ = new_E4498_ & ~new_E4512_;
  assign new_E4559_ = ~new_E4498_ & new_E4512_;
  assign new_E4560_ = new_F3481_;
  assign new_E4561_ = new_F3548_;
  assign new_E4562_ = new_F3615_;
  assign new_E4563_ = new_F3682_;
  assign new_E4564_ = new_F3749_;
  assign new_E4565_ = new_F3816_;
  assign new_E4566_ = new_E4573_ & new_E4572_;
  assign new_E4567_ = new_E4575_ | new_E4574_;
  assign new_E4568_ = new_E4577_ | new_E4576_;
  assign new_E4569_ = new_E4579_ & new_E4578_;
  assign new_E4570_ = new_E4579_ & new_E4580_;
  assign new_E4571_ = new_E4572_ | new_E4581_;
  assign new_E4572_ = new_E4561_ | new_E4584_;
  assign new_E4573_ = new_E4583_ | new_E4582_;
  assign new_E4574_ = new_E4588_ & new_E4587_;
  assign new_E4575_ = new_E4586_ & new_E4585_;
  assign new_E4576_ = new_E4591_ | new_E4590_;
  assign new_E4577_ = new_E4586_ & new_E4589_;
  assign new_E4578_ = new_E4561_ | new_E4594_;
  assign new_E4579_ = new_E4593_ | new_E4592_;
  assign new_E4580_ = new_E4596_ | new_E4595_;
  assign new_E4581_ = ~new_E4572_ & new_E4598_;
  assign new_E4582_ = ~new_E4574_ & new_E4586_;
  assign new_E4583_ = new_E4574_ & ~new_E4586_;
  assign new_E4584_ = new_E4560_ & ~new_E4561_;
  assign new_E4585_ = ~new_E4607_ | ~new_E4608_;
  assign new_E4586_ = new_E4600_ | new_E4602_;
  assign new_E4587_ = new_E4610_ | new_E4609_;
  assign new_E4588_ = new_E4604_ | new_E4603_;
  assign new_E4589_ = ~new_E4612_ | ~new_E4611_;
  assign new_E4590_ = ~new_E4613_ & new_E4614_;
  assign new_E4591_ = new_E4613_ & ~new_E4614_;
  assign new_E4592_ = ~new_E4560_ & new_E4561_;
  assign new_E4593_ = new_E4560_ & ~new_E4561_;
  assign new_E4594_ = ~new_E4576_ | new_E4586_;
  assign new_E4595_ = new_E4576_ & new_E4586_;
  assign new_E4596_ = ~new_E4576_ & ~new_E4586_;
  assign new_E4597_ = new_E4618_ | new_E4617_;
  assign new_E4598_ = new_E4564_ | new_E4597_;
  assign new_E4599_ = new_E4622_ | new_E4621_;
  assign new_E4600_ = ~new_E4564_ & new_E4599_;
  assign new_E4601_ = new_E4620_ | new_E4619_;
  assign new_E4602_ = new_E4564_ & new_E4601_;
  assign new_E4603_ = new_E4562_ & ~new_E4572_;
  assign new_E4604_ = ~new_E4562_ & new_E4572_;
  assign new_E4605_ = ~new_E4561_ | ~new_E4586_;
  assign new_E4606_ = new_E4572_ & new_E4605_;
  assign new_E4607_ = ~new_E4572_ & ~new_E4606_;
  assign new_E4608_ = new_E4572_ | new_E4605_;
  assign new_E4609_ = ~new_E4562_ & new_E4563_;
  assign new_E4610_ = new_E4562_ & ~new_E4563_;
  assign new_E4611_ = new_E4579_ | new_E4616_;
  assign new_E4612_ = ~new_E4579_ & ~new_E4615_;
  assign new_E4613_ = new_E4562_ | new_E4579_;
  assign new_E4614_ = new_E4562_ | new_E4563_;
  assign new_E4615_ = new_E4579_ & new_E4616_;
  assign new_E4616_ = ~new_E4561_ | ~new_E4586_;
  assign new_E4617_ = new_E4594_ & new_E4614_;
  assign new_E4618_ = ~new_E4594_ & ~new_E4614_;
  assign new_E4619_ = new_E4623_ | new_E4624_;
  assign new_E4620_ = ~new_E4565_ & new_E4579_;
  assign new_E4621_ = new_E4625_ | new_E4626_;
  assign new_E4622_ = new_E4565_ & new_E4579_;
  assign new_E4623_ = ~new_E4565_ & ~new_E4579_;
  assign new_E4624_ = new_E4565_ & ~new_E4579_;
  assign new_E4625_ = new_E4565_ & ~new_E4579_;
  assign new_E4626_ = ~new_E4565_ & new_E4579_;
  assign new_E4627_ = new_F3883_;
  assign new_E4628_ = new_F3950_;
  assign new_E4629_ = new_F4017_;
  assign new_E4630_ = new_F4084_;
  assign new_E4631_ = new_F4151_;
  assign new_E4632_ = new_F4218_;
  assign new_E4633_ = new_E4640_ & new_E4639_;
  assign new_E4634_ = new_E4642_ | new_E4641_;
  assign new_E4635_ = new_E4644_ | new_E4643_;
  assign new_E4636_ = new_E4646_ & new_E4645_;
  assign new_E4637_ = new_E4646_ & new_E4647_;
  assign new_E4638_ = new_E4639_ | new_E4648_;
  assign new_E4639_ = new_E4628_ | new_E4651_;
  assign new_E4640_ = new_E4650_ | new_E4649_;
  assign new_E4641_ = new_E4655_ & new_E4654_;
  assign new_E4642_ = new_E4653_ & new_E4652_;
  assign new_E4643_ = new_E4658_ | new_E4657_;
  assign new_E4644_ = new_E4653_ & new_E4656_;
  assign new_E4645_ = new_E4628_ | new_E4661_;
  assign new_E4646_ = new_E4660_ | new_E4659_;
  assign new_E4647_ = new_E4663_ | new_E4662_;
  assign new_E4648_ = ~new_E4639_ & new_E4665_;
  assign new_E4649_ = ~new_E4641_ & new_E4653_;
  assign new_E4650_ = new_E4641_ & ~new_E4653_;
  assign new_E4651_ = new_E4627_ & ~new_E4628_;
  assign new_E4652_ = ~new_E4674_ | ~new_E4675_;
  assign new_E4653_ = new_E4667_ | new_E4669_;
  assign new_E4654_ = new_E4677_ | new_E4676_;
  assign new_E4655_ = new_E4671_ | new_E4670_;
  assign new_E4656_ = ~new_E4679_ | ~new_E4678_;
  assign new_E4657_ = ~new_E4680_ & new_E4681_;
  assign new_E4658_ = new_E4680_ & ~new_E4681_;
  assign new_E4659_ = ~new_E4627_ & new_E4628_;
  assign new_E4660_ = new_E4627_ & ~new_E4628_;
  assign new_E4661_ = ~new_E4643_ | new_E4653_;
  assign new_E4662_ = new_E4643_ & new_E4653_;
  assign new_E4663_ = ~new_E4643_ & ~new_E4653_;
  assign new_E4664_ = new_E4685_ | new_E4684_;
  assign new_E4665_ = new_E4631_ | new_E4664_;
  assign new_E4666_ = new_E4689_ | new_E4688_;
  assign new_E4667_ = ~new_E4631_ & new_E4666_;
  assign new_E4668_ = new_E4687_ | new_E4686_;
  assign new_E4669_ = new_E4631_ & new_E4668_;
  assign new_E4670_ = new_E4629_ & ~new_E4639_;
  assign new_E4671_ = ~new_E4629_ & new_E4639_;
  assign new_E4672_ = ~new_E4628_ | ~new_E4653_;
  assign new_E4673_ = new_E4639_ & new_E4672_;
  assign new_E4674_ = ~new_E4639_ & ~new_E4673_;
  assign new_E4675_ = new_E4639_ | new_E4672_;
  assign new_E4676_ = ~new_E4629_ & new_E4630_;
  assign new_E4677_ = new_E4629_ & ~new_E4630_;
  assign new_E4678_ = new_E4646_ | new_E4683_;
  assign new_E4679_ = ~new_E4646_ & ~new_E4682_;
  assign new_E4680_ = new_E4629_ | new_E4646_;
  assign new_E4681_ = new_E4629_ | new_E4630_;
  assign new_E4682_ = new_E4646_ & new_E4683_;
  assign new_E4683_ = ~new_E4628_ | ~new_E4653_;
  assign new_E4684_ = new_E4661_ & new_E4681_;
  assign new_E4685_ = ~new_E4661_ & ~new_E4681_;
  assign new_E4686_ = new_E4690_ | new_E4691_;
  assign new_E4687_ = ~new_E4632_ & new_E4646_;
  assign new_E4688_ = new_E4692_ | new_E4693_;
  assign new_E4689_ = new_E4632_ & new_E4646_;
  assign new_E4690_ = ~new_E4632_ & ~new_E4646_;
  assign new_E4691_ = new_E4632_ & ~new_E4646_;
  assign new_E4692_ = new_E4632_ & ~new_E4646_;
  assign new_E4693_ = ~new_E4632_ & new_E4646_;
  assign new_E4694_ = new_F4285_;
  assign new_E4695_ = new_F4352_;
  assign new_E4696_ = new_F4419_;
  assign new_E4697_ = new_F4486_;
  assign new_E4698_ = new_F4553_;
  assign new_E4699_ = new_F4620_;
  assign new_E4700_ = new_E4707_ & new_E4706_;
  assign new_E4701_ = new_E4709_ | new_E4708_;
  assign new_E4702_ = new_E4711_ | new_E4710_;
  assign new_E4703_ = new_E4713_ & new_E4712_;
  assign new_E4704_ = new_E4713_ & new_E4714_;
  assign new_E4705_ = new_E4706_ | new_E4715_;
  assign new_E4706_ = new_E4695_ | new_E4718_;
  assign new_E4707_ = new_E4717_ | new_E4716_;
  assign new_E4708_ = new_E4722_ & new_E4721_;
  assign new_E4709_ = new_E4720_ & new_E4719_;
  assign new_E4710_ = new_E4725_ | new_E4724_;
  assign new_E4711_ = new_E4720_ & new_E4723_;
  assign new_E4712_ = new_E4695_ | new_E4728_;
  assign new_E4713_ = new_E4727_ | new_E4726_;
  assign new_E4714_ = new_E4730_ | new_E4729_;
  assign new_E4715_ = ~new_E4706_ & new_E4732_;
  assign new_E4716_ = ~new_E4708_ & new_E4720_;
  assign new_E4717_ = new_E4708_ & ~new_E4720_;
  assign new_E4718_ = new_E4694_ & ~new_E4695_;
  assign new_E4719_ = ~new_E4741_ | ~new_E4742_;
  assign new_E4720_ = new_E4734_ | new_E4736_;
  assign new_E4721_ = new_E4744_ | new_E4743_;
  assign new_E4722_ = new_E4738_ | new_E4737_;
  assign new_E4723_ = ~new_E4746_ | ~new_E4745_;
  assign new_E4724_ = ~new_E4747_ & new_E4748_;
  assign new_E4725_ = new_E4747_ & ~new_E4748_;
  assign new_E4726_ = ~new_E4694_ & new_E4695_;
  assign new_E4727_ = new_E4694_ & ~new_E4695_;
  assign new_E4728_ = ~new_E4710_ | new_E4720_;
  assign new_E4729_ = new_E4710_ & new_E4720_;
  assign new_E4730_ = ~new_E4710_ & ~new_E4720_;
  assign new_E4731_ = new_E4752_ | new_E4751_;
  assign new_E4732_ = new_E4698_ | new_E4731_;
  assign new_E4733_ = new_E4756_ | new_E4755_;
  assign new_E4734_ = ~new_E4698_ & new_E4733_;
  assign new_E4735_ = new_E4754_ | new_E4753_;
  assign new_E4736_ = new_E4698_ & new_E4735_;
  assign new_E4737_ = new_E4696_ & ~new_E4706_;
  assign new_E4738_ = ~new_E4696_ & new_E4706_;
  assign new_E4739_ = ~new_E4695_ | ~new_E4720_;
  assign new_E4740_ = new_E4706_ & new_E4739_;
  assign new_E4741_ = ~new_E4706_ & ~new_E4740_;
  assign new_E4742_ = new_E4706_ | new_E4739_;
  assign new_E4743_ = ~new_E4696_ & new_E4697_;
  assign new_E4744_ = new_E4696_ & ~new_E4697_;
  assign new_E4745_ = new_E4713_ | new_E4750_;
  assign new_E4746_ = ~new_E4713_ & ~new_E4749_;
  assign new_E4747_ = new_E4696_ | new_E4713_;
  assign new_E4748_ = new_E4696_ | new_E4697_;
  assign new_E4749_ = new_E4713_ & new_E4750_;
  assign new_E4750_ = ~new_E4695_ | ~new_E4720_;
  assign new_E4751_ = new_E4728_ & new_E4748_;
  assign new_E4752_ = ~new_E4728_ & ~new_E4748_;
  assign new_E4753_ = new_E4757_ | new_E4758_;
  assign new_E4754_ = ~new_E4699_ & new_E4713_;
  assign new_E4755_ = new_E4759_ | new_E4760_;
  assign new_E4756_ = new_E4699_ & new_E4713_;
  assign new_E4757_ = ~new_E4699_ & ~new_E4713_;
  assign new_E4758_ = new_E4699_ & ~new_E4713_;
  assign new_E4759_ = new_E4699_ & ~new_E4713_;
  assign new_E4760_ = ~new_E4699_ & new_E4713_;
  assign new_E4761_ = new_F4687_;
  assign new_E4762_ = new_F4754_;
  assign new_E4763_ = new_F4821_;
  assign new_E4764_ = new_F4888_;
  assign new_E4765_ = new_F4955_;
  assign new_E4766_ = new_F5022_;
  assign new_E4767_ = new_E4774_ & new_E4773_;
  assign new_E4768_ = new_E4776_ | new_E4775_;
  assign new_E4769_ = new_E4778_ | new_E4777_;
  assign new_E4770_ = new_E4780_ & new_E4779_;
  assign new_E4771_ = new_E4780_ & new_E4781_;
  assign new_E4772_ = new_E4773_ | new_E4782_;
  assign new_E4773_ = new_E4762_ | new_E4785_;
  assign new_E4774_ = new_E4784_ | new_E4783_;
  assign new_E4775_ = new_E4789_ & new_E4788_;
  assign new_E4776_ = new_E4787_ & new_E4786_;
  assign new_E4777_ = new_E4792_ | new_E4791_;
  assign new_E4778_ = new_E4787_ & new_E4790_;
  assign new_E4779_ = new_E4762_ | new_E4795_;
  assign new_E4780_ = new_E4794_ | new_E4793_;
  assign new_E4781_ = new_E4797_ | new_E4796_;
  assign new_E4782_ = ~new_E4773_ & new_E4799_;
  assign new_E4783_ = ~new_E4775_ & new_E4787_;
  assign new_E4784_ = new_E4775_ & ~new_E4787_;
  assign new_E4785_ = new_E4761_ & ~new_E4762_;
  assign new_E4786_ = ~new_E4808_ | ~new_E4809_;
  assign new_E4787_ = new_E4801_ | new_E4803_;
  assign new_E4788_ = new_E4811_ | new_E4810_;
  assign new_E4789_ = new_E4805_ | new_E4804_;
  assign new_E4790_ = ~new_E4813_ | ~new_E4812_;
  assign new_E4791_ = ~new_E4814_ & new_E4815_;
  assign new_E4792_ = new_E4814_ & ~new_E4815_;
  assign new_E4793_ = ~new_E4761_ & new_E4762_;
  assign new_E4794_ = new_E4761_ & ~new_E4762_;
  assign new_E4795_ = ~new_E4777_ | new_E4787_;
  assign new_E4796_ = new_E4777_ & new_E4787_;
  assign new_E4797_ = ~new_E4777_ & ~new_E4787_;
  assign new_E4798_ = new_E4819_ | new_E4818_;
  assign new_E4799_ = new_E4765_ | new_E4798_;
  assign new_E4800_ = new_E4823_ | new_E4822_;
  assign new_E4801_ = ~new_E4765_ & new_E4800_;
  assign new_E4802_ = new_E4821_ | new_E4820_;
  assign new_E4803_ = new_E4765_ & new_E4802_;
  assign new_E4804_ = new_E4763_ & ~new_E4773_;
  assign new_E4805_ = ~new_E4763_ & new_E4773_;
  assign new_E4806_ = ~new_E4762_ | ~new_E4787_;
  assign new_E4807_ = new_E4773_ & new_E4806_;
  assign new_E4808_ = ~new_E4773_ & ~new_E4807_;
  assign new_E4809_ = new_E4773_ | new_E4806_;
  assign new_E4810_ = ~new_E4763_ & new_E4764_;
  assign new_E4811_ = new_E4763_ & ~new_E4764_;
  assign new_E4812_ = new_E4780_ | new_E4817_;
  assign new_E4813_ = ~new_E4780_ & ~new_E4816_;
  assign new_E4814_ = new_E4763_ | new_E4780_;
  assign new_E4815_ = new_E4763_ | new_E4764_;
  assign new_E4816_ = new_E4780_ & new_E4817_;
  assign new_E4817_ = ~new_E4762_ | ~new_E4787_;
  assign new_E4818_ = new_E4795_ & new_E4815_;
  assign new_E4819_ = ~new_E4795_ & ~new_E4815_;
  assign new_E4820_ = new_E4824_ | new_E4825_;
  assign new_E4821_ = ~new_E4766_ & new_E4780_;
  assign new_E4822_ = new_E4826_ | new_E4827_;
  assign new_E4823_ = new_E4766_ & new_E4780_;
  assign new_E4824_ = ~new_E4766_ & ~new_E4780_;
  assign new_E4825_ = new_E4766_ & ~new_E4780_;
  assign new_E4826_ = new_E4766_ & ~new_E4780_;
  assign new_E4827_ = ~new_E4766_ & new_E4780_;
  assign new_E4828_ = new_F5089_;
  assign new_E4829_ = new_F5156_;
  assign new_E4830_ = new_F5223_;
  assign new_E4831_ = new_F5290_;
  assign new_E4832_ = new_F5357_;
  assign new_E4833_ = new_F5424_;
  assign new_E4834_ = new_E4841_ & new_E4840_;
  assign new_E4835_ = new_E4843_ | new_E4842_;
  assign new_E4836_ = new_E4845_ | new_E4844_;
  assign new_E4837_ = new_E4847_ & new_E4846_;
  assign new_E4838_ = new_E4847_ & new_E4848_;
  assign new_E4839_ = new_E4840_ | new_E4849_;
  assign new_E4840_ = new_E4829_ | new_E4852_;
  assign new_E4841_ = new_E4851_ | new_E4850_;
  assign new_E4842_ = new_E4856_ & new_E4855_;
  assign new_E4843_ = new_E4854_ & new_E4853_;
  assign new_E4844_ = new_E4859_ | new_E4858_;
  assign new_E4845_ = new_E4854_ & new_E4857_;
  assign new_E4846_ = new_E4829_ | new_E4862_;
  assign new_E4847_ = new_E4861_ | new_E4860_;
  assign new_E4848_ = new_E4864_ | new_E4863_;
  assign new_E4849_ = ~new_E4840_ & new_E4866_;
  assign new_E4850_ = ~new_E4842_ & new_E4854_;
  assign new_E4851_ = new_E4842_ & ~new_E4854_;
  assign new_E4852_ = new_E4828_ & ~new_E4829_;
  assign new_E4853_ = ~new_E4875_ | ~new_E4876_;
  assign new_E4854_ = new_E4868_ | new_E4870_;
  assign new_E4855_ = new_E4878_ | new_E4877_;
  assign new_E4856_ = new_E4872_ | new_E4871_;
  assign new_E4857_ = ~new_E4880_ | ~new_E4879_;
  assign new_E4858_ = ~new_E4881_ & new_E4882_;
  assign new_E4859_ = new_E4881_ & ~new_E4882_;
  assign new_E4860_ = ~new_E4828_ & new_E4829_;
  assign new_E4861_ = new_E4828_ & ~new_E4829_;
  assign new_E4862_ = ~new_E4844_ | new_E4854_;
  assign new_E4863_ = new_E4844_ & new_E4854_;
  assign new_E4864_ = ~new_E4844_ & ~new_E4854_;
  assign new_E4865_ = new_E4886_ | new_E4885_;
  assign new_E4866_ = new_E4832_ | new_E4865_;
  assign new_E4867_ = new_E4890_ | new_E4889_;
  assign new_E4868_ = ~new_E4832_ & new_E4867_;
  assign new_E4869_ = new_E4888_ | new_E4887_;
  assign new_E4870_ = new_E4832_ & new_E4869_;
  assign new_E4871_ = new_E4830_ & ~new_E4840_;
  assign new_E4872_ = ~new_E4830_ & new_E4840_;
  assign new_E4873_ = ~new_E4829_ | ~new_E4854_;
  assign new_E4874_ = new_E4840_ & new_E4873_;
  assign new_E4875_ = ~new_E4840_ & ~new_E4874_;
  assign new_E4876_ = new_E4840_ | new_E4873_;
  assign new_E4877_ = ~new_E4830_ & new_E4831_;
  assign new_E4878_ = new_E4830_ & ~new_E4831_;
  assign new_E4879_ = new_E4847_ | new_E4884_;
  assign new_E4880_ = ~new_E4847_ & ~new_E4883_;
  assign new_E4881_ = new_E4830_ | new_E4847_;
  assign new_E4882_ = new_E4830_ | new_E4831_;
  assign new_E4883_ = new_E4847_ & new_E4884_;
  assign new_E4884_ = ~new_E4829_ | ~new_E4854_;
  assign new_E4885_ = new_E4862_ & new_E4882_;
  assign new_E4886_ = ~new_E4862_ & ~new_E4882_;
  assign new_E4887_ = new_E4891_ | new_E4892_;
  assign new_E4888_ = ~new_E4833_ & new_E4847_;
  assign new_E4889_ = new_E4893_ | new_E4894_;
  assign new_E4890_ = new_E4833_ & new_E4847_;
  assign new_E4891_ = ~new_E4833_ & ~new_E4847_;
  assign new_E4892_ = new_E4833_ & ~new_E4847_;
  assign new_E4893_ = new_E4833_ & ~new_E4847_;
  assign new_E4894_ = ~new_E4833_ & new_E4847_;
  assign new_E4895_ = new_F5491_;
  assign new_E4896_ = new_F5558_;
  assign new_E4897_ = new_F5625_;
  assign new_E4898_ = new_F5692_;
  assign new_E4899_ = new_F5759_;
  assign new_E4900_ = new_F5826_;
  assign new_E4901_ = new_E4908_ & new_E4907_;
  assign new_E4902_ = new_E4910_ | new_E4909_;
  assign new_E4903_ = new_E4912_ | new_E4911_;
  assign new_E4904_ = new_E4914_ & new_E4913_;
  assign new_E4905_ = new_E4914_ & new_E4915_;
  assign new_E4906_ = new_E4907_ | new_E4916_;
  assign new_E4907_ = new_E4896_ | new_E4919_;
  assign new_E4908_ = new_E4918_ | new_E4917_;
  assign new_E4909_ = new_E4923_ & new_E4922_;
  assign new_E4910_ = new_E4921_ & new_E4920_;
  assign new_E4911_ = new_E4926_ | new_E4925_;
  assign new_E4912_ = new_E4921_ & new_E4924_;
  assign new_E4913_ = new_E4896_ | new_E4929_;
  assign new_E4914_ = new_E4928_ | new_E4927_;
  assign new_E4915_ = new_E4931_ | new_E4930_;
  assign new_E4916_ = ~new_E4907_ & new_E4933_;
  assign new_E4917_ = ~new_E4909_ & new_E4921_;
  assign new_E4918_ = new_E4909_ & ~new_E4921_;
  assign new_E4919_ = new_E4895_ & ~new_E4896_;
  assign new_E4920_ = ~new_E4942_ | ~new_E4943_;
  assign new_E4921_ = new_E4935_ | new_E4937_;
  assign new_E4922_ = new_E4945_ | new_E4944_;
  assign new_E4923_ = new_E4939_ | new_E4938_;
  assign new_E4924_ = ~new_E4947_ | ~new_E4946_;
  assign new_E4925_ = ~new_E4948_ & new_E4949_;
  assign new_E4926_ = new_E4948_ & ~new_E4949_;
  assign new_E4927_ = ~new_E4895_ & new_E4896_;
  assign new_E4928_ = new_E4895_ & ~new_E4896_;
  assign new_E4929_ = ~new_E4911_ | new_E4921_;
  assign new_E4930_ = new_E4911_ & new_E4921_;
  assign new_E4931_ = ~new_E4911_ & ~new_E4921_;
  assign new_E4932_ = new_E4953_ | new_E4952_;
  assign new_E4933_ = new_E4899_ | new_E4932_;
  assign new_E4934_ = new_E4957_ | new_E4956_;
  assign new_E4935_ = ~new_E4899_ & new_E4934_;
  assign new_E4936_ = new_E4955_ | new_E4954_;
  assign new_E4937_ = new_E4899_ & new_E4936_;
  assign new_E4938_ = new_E4897_ & ~new_E4907_;
  assign new_E4939_ = ~new_E4897_ & new_E4907_;
  assign new_E4940_ = ~new_E4896_ | ~new_E4921_;
  assign new_E4941_ = new_E4907_ & new_E4940_;
  assign new_E4942_ = ~new_E4907_ & ~new_E4941_;
  assign new_E4943_ = new_E4907_ | new_E4940_;
  assign new_E4944_ = ~new_E4897_ & new_E4898_;
  assign new_E4945_ = new_E4897_ & ~new_E4898_;
  assign new_E4946_ = new_E4914_ | new_E4951_;
  assign new_E4947_ = ~new_E4914_ & ~new_E4950_;
  assign new_E4948_ = new_E4897_ | new_E4914_;
  assign new_E4949_ = new_E4897_ | new_E4898_;
  assign new_E4950_ = new_E4914_ & new_E4951_;
  assign new_E4951_ = ~new_E4896_ | ~new_E4921_;
  assign new_E4952_ = new_E4929_ & new_E4949_;
  assign new_E4953_ = ~new_E4929_ & ~new_E4949_;
  assign new_E4954_ = new_E4958_ | new_E4959_;
  assign new_E4955_ = ~new_E4900_ & new_E4914_;
  assign new_E4956_ = new_E4960_ | new_E4961_;
  assign new_E4957_ = new_E4900_ & new_E4914_;
  assign new_E4958_ = ~new_E4900_ & ~new_E4914_;
  assign new_E4959_ = new_E4900_ & ~new_E4914_;
  assign new_E4960_ = new_E4900_ & ~new_E4914_;
  assign new_E4961_ = ~new_E4900_ & new_E4914_;
  assign new_E4962_ = new_F5893_;
  assign new_E4963_ = new_F5960_;
  assign new_E4964_ = new_F6027_;
  assign new_E4965_ = new_F6094_;
  assign new_E4966_ = new_F6161_;
  assign new_E4967_ = new_F6228_;
  assign new_E4968_ = new_E4975_ & new_E4974_;
  assign new_E4969_ = new_E4977_ | new_E4976_;
  assign new_E4970_ = new_E4979_ | new_E4978_;
  assign new_E4971_ = new_E4981_ & new_E4980_;
  assign new_E4972_ = new_E4981_ & new_E4982_;
  assign new_E4973_ = new_E4974_ | new_E4983_;
  assign new_E4974_ = new_E4963_ | new_E4986_;
  assign new_E4975_ = new_E4985_ | new_E4984_;
  assign new_E4976_ = new_E4990_ & new_E4989_;
  assign new_E4977_ = new_E4988_ & new_E4987_;
  assign new_E4978_ = new_E4993_ | new_E4992_;
  assign new_E4979_ = new_E4988_ & new_E4991_;
  assign new_E4980_ = new_E4963_ | new_E4996_;
  assign new_E4981_ = new_E4995_ | new_E4994_;
  assign new_E4982_ = new_E4998_ | new_E4997_;
  assign new_E4983_ = ~new_E4974_ & new_E5000_;
  assign new_E4984_ = ~new_E4976_ & new_E4988_;
  assign new_E4985_ = new_E4976_ & ~new_E4988_;
  assign new_E4986_ = new_E4962_ & ~new_E4963_;
  assign new_E4987_ = ~new_E5009_ | ~new_E5010_;
  assign new_E4988_ = new_E5002_ | new_E5004_;
  assign new_E4989_ = new_E5012_ | new_E5011_;
  assign new_E4990_ = new_E5006_ | new_E5005_;
  assign new_E4991_ = ~new_E5014_ | ~new_E5013_;
  assign new_E4992_ = ~new_E5015_ & new_E5016_;
  assign new_E4993_ = new_E5015_ & ~new_E5016_;
  assign new_E4994_ = ~new_E4962_ & new_E4963_;
  assign new_E4995_ = new_E4962_ & ~new_E4963_;
  assign new_E4996_ = ~new_E4978_ | new_E4988_;
  assign new_E4997_ = new_E4978_ & new_E4988_;
  assign new_E4998_ = ~new_E4978_ & ~new_E4988_;
  assign new_E4999_ = new_E5020_ | new_E5019_;
  assign new_E5000_ = new_E4966_ | new_E4999_;
  assign new_E5001_ = new_E5024_ | new_E5023_;
  assign new_E5002_ = ~new_E4966_ & new_E5001_;
  assign new_E5003_ = new_E5022_ | new_E5021_;
  assign new_E5004_ = new_E4966_ & new_E5003_;
  assign new_E5005_ = new_E4964_ & ~new_E4974_;
  assign new_E5006_ = ~new_E4964_ & new_E4974_;
  assign new_E5007_ = ~new_E4963_ | ~new_E4988_;
  assign new_E5008_ = new_E4974_ & new_E5007_;
  assign new_E5009_ = ~new_E4974_ & ~new_E5008_;
  assign new_E5010_ = new_E4974_ | new_E5007_;
  assign new_E5011_ = ~new_E4964_ & new_E4965_;
  assign new_E5012_ = new_E4964_ & ~new_E4965_;
  assign new_E5013_ = new_E4981_ | new_E5018_;
  assign new_E5014_ = ~new_E4981_ & ~new_E5017_;
  assign new_E5015_ = new_E4964_ | new_E4981_;
  assign new_E5016_ = new_E4964_ | new_E4965_;
  assign new_E5017_ = new_E4981_ & new_E5018_;
  assign new_E5018_ = ~new_E4963_ | ~new_E4988_;
  assign new_E5019_ = new_E4996_ & new_E5016_;
  assign new_E5020_ = ~new_E4996_ & ~new_E5016_;
  assign new_E5021_ = new_E5025_ | new_E5026_;
  assign new_E5022_ = ~new_E4967_ & new_E4981_;
  assign new_E5023_ = new_E5027_ | new_E5028_;
  assign new_E5024_ = new_E4967_ & new_E4981_;
  assign new_E5025_ = ~new_E4967_ & ~new_E4981_;
  assign new_E5026_ = new_E4967_ & ~new_E4981_;
  assign new_E5027_ = new_E4967_ & ~new_E4981_;
  assign new_E5028_ = ~new_E4967_ & new_E4981_;
  assign new_E5029_ = new_F6295_;
  assign new_E5030_ = new_F6362_;
  assign new_E5031_ = new_F6429_;
  assign new_E5032_ = new_F6496_;
  assign new_E5033_ = new_F6563_;
  assign new_E5034_ = new_F6630_;
  assign new_E5035_ = new_E5042_ & new_E5041_;
  assign new_E5036_ = new_E5044_ | new_E5043_;
  assign new_E5037_ = new_E5046_ | new_E5045_;
  assign new_E5038_ = new_E5048_ & new_E5047_;
  assign new_E5039_ = new_E5048_ & new_E5049_;
  assign new_E5040_ = new_E5041_ | new_E5050_;
  assign new_E5041_ = new_E5030_ | new_E5053_;
  assign new_E5042_ = new_E5052_ | new_E5051_;
  assign new_E5043_ = new_E5057_ & new_E5056_;
  assign new_E5044_ = new_E5055_ & new_E5054_;
  assign new_E5045_ = new_E5060_ | new_E5059_;
  assign new_E5046_ = new_E5055_ & new_E5058_;
  assign new_E5047_ = new_E5030_ | new_E5063_;
  assign new_E5048_ = new_E5062_ | new_E5061_;
  assign new_E5049_ = new_E5065_ | new_E5064_;
  assign new_E5050_ = ~new_E5041_ & new_E5067_;
  assign new_E5051_ = ~new_E5043_ & new_E5055_;
  assign new_E5052_ = new_E5043_ & ~new_E5055_;
  assign new_E5053_ = new_E5029_ & ~new_E5030_;
  assign new_E5054_ = ~new_E5076_ | ~new_E5077_;
  assign new_E5055_ = new_E5069_ | new_E5071_;
  assign new_E5056_ = new_E5079_ | new_E5078_;
  assign new_E5057_ = new_E5073_ | new_E5072_;
  assign new_E5058_ = ~new_E5081_ | ~new_E5080_;
  assign new_E5059_ = ~new_E5082_ & new_E5083_;
  assign new_E5060_ = new_E5082_ & ~new_E5083_;
  assign new_E5061_ = ~new_E5029_ & new_E5030_;
  assign new_E5062_ = new_E5029_ & ~new_E5030_;
  assign new_E5063_ = ~new_E5045_ | new_E5055_;
  assign new_E5064_ = new_E5045_ & new_E5055_;
  assign new_E5065_ = ~new_E5045_ & ~new_E5055_;
  assign new_E5066_ = new_E5087_ | new_E5086_;
  assign new_E5067_ = new_E5033_ | new_E5066_;
  assign new_E5068_ = new_E5091_ | new_E5090_;
  assign new_E5069_ = ~new_E5033_ & new_E5068_;
  assign new_E5070_ = new_E5089_ | new_E5088_;
  assign new_E5071_ = new_E5033_ & new_E5070_;
  assign new_E5072_ = new_E5031_ & ~new_E5041_;
  assign new_E5073_ = ~new_E5031_ & new_E5041_;
  assign new_E5074_ = ~new_E5030_ | ~new_E5055_;
  assign new_E5075_ = new_E5041_ & new_E5074_;
  assign new_E5076_ = ~new_E5041_ & ~new_E5075_;
  assign new_E5077_ = new_E5041_ | new_E5074_;
  assign new_E5078_ = ~new_E5031_ & new_E5032_;
  assign new_E5079_ = new_E5031_ & ~new_E5032_;
  assign new_E5080_ = new_E5048_ | new_E5085_;
  assign new_E5081_ = ~new_E5048_ & ~new_E5084_;
  assign new_E5082_ = new_E5031_ | new_E5048_;
  assign new_E5083_ = new_E5031_ | new_E5032_;
  assign new_E5084_ = new_E5048_ & new_E5085_;
  assign new_E5085_ = ~new_E5030_ | ~new_E5055_;
  assign new_E5086_ = new_E5063_ & new_E5083_;
  assign new_E5087_ = ~new_E5063_ & ~new_E5083_;
  assign new_E5088_ = new_E5092_ | new_E5093_;
  assign new_E5089_ = ~new_E5034_ & new_E5048_;
  assign new_E5090_ = new_E5094_ | new_E5095_;
  assign new_E5091_ = new_E5034_ & new_E5048_;
  assign new_E5092_ = ~new_E5034_ & ~new_E5048_;
  assign new_E5093_ = new_E5034_ & ~new_E5048_;
  assign new_E5094_ = new_E5034_ & ~new_E5048_;
  assign new_E5095_ = ~new_E5034_ & new_E5048_;
  assign new_E5096_ = new_F6697_;
  assign new_E5097_ = new_F6764_;
  assign new_E5098_ = new_F6831_;
  assign new_E5099_ = new_F6898_;
  assign new_E5100_ = new_F6965_;
  assign new_E5101_ = new_F7032_;
  assign new_E5102_ = new_E5109_ & new_E5108_;
  assign new_E5103_ = new_E5111_ | new_E5110_;
  assign new_E5104_ = new_E5113_ | new_E5112_;
  assign new_E5105_ = new_E5115_ & new_E5114_;
  assign new_E5106_ = new_E5115_ & new_E5116_;
  assign new_E5107_ = new_E5108_ | new_E5117_;
  assign new_E5108_ = new_E5097_ | new_E5120_;
  assign new_E5109_ = new_E5119_ | new_E5118_;
  assign new_E5110_ = new_E5124_ & new_E5123_;
  assign new_E5111_ = new_E5122_ & new_E5121_;
  assign new_E5112_ = new_E5127_ | new_E5126_;
  assign new_E5113_ = new_E5122_ & new_E5125_;
  assign new_E5114_ = new_E5097_ | new_E5130_;
  assign new_E5115_ = new_E5129_ | new_E5128_;
  assign new_E5116_ = new_E5132_ | new_E5131_;
  assign new_E5117_ = ~new_E5108_ & new_E5134_;
  assign new_E5118_ = ~new_E5110_ & new_E5122_;
  assign new_E5119_ = new_E5110_ & ~new_E5122_;
  assign new_E5120_ = new_E5096_ & ~new_E5097_;
  assign new_E5121_ = ~new_E5143_ | ~new_E5144_;
  assign new_E5122_ = new_E5136_ | new_E5138_;
  assign new_E5123_ = new_E5146_ | new_E5145_;
  assign new_E5124_ = new_E5140_ | new_E5139_;
  assign new_E5125_ = ~new_E5148_ | ~new_E5147_;
  assign new_E5126_ = ~new_E5149_ & new_E5150_;
  assign new_E5127_ = new_E5149_ & ~new_E5150_;
  assign new_E5128_ = ~new_E5096_ & new_E5097_;
  assign new_E5129_ = new_E5096_ & ~new_E5097_;
  assign new_E5130_ = ~new_E5112_ | new_E5122_;
  assign new_E5131_ = new_E5112_ & new_E5122_;
  assign new_E5132_ = ~new_E5112_ & ~new_E5122_;
  assign new_E5133_ = new_E5154_ | new_E5153_;
  assign new_E5134_ = new_E5100_ | new_E5133_;
  assign new_E5135_ = new_E5158_ | new_E5157_;
  assign new_E5136_ = ~new_E5100_ & new_E5135_;
  assign new_E5137_ = new_E5156_ | new_E5155_;
  assign new_E5138_ = new_E5100_ & new_E5137_;
  assign new_E5139_ = new_E5098_ & ~new_E5108_;
  assign new_E5140_ = ~new_E5098_ & new_E5108_;
  assign new_E5141_ = ~new_E5097_ | ~new_E5122_;
  assign new_E5142_ = new_E5108_ & new_E5141_;
  assign new_E5143_ = ~new_E5108_ & ~new_E5142_;
  assign new_E5144_ = new_E5108_ | new_E5141_;
  assign new_E5145_ = ~new_E5098_ & new_E5099_;
  assign new_E5146_ = new_E5098_ & ~new_E5099_;
  assign new_E5147_ = new_E5115_ | new_E5152_;
  assign new_E5148_ = ~new_E5115_ & ~new_E5151_;
  assign new_E5149_ = new_E5098_ | new_E5115_;
  assign new_E5150_ = new_E5098_ | new_E5099_;
  assign new_E5151_ = new_E5115_ & new_E5152_;
  assign new_E5152_ = ~new_E5097_ | ~new_E5122_;
  assign new_E5153_ = new_E5130_ & new_E5150_;
  assign new_E5154_ = ~new_E5130_ & ~new_E5150_;
  assign new_E5155_ = new_E5159_ | new_E5160_;
  assign new_E5156_ = ~new_E5101_ & new_E5115_;
  assign new_E5157_ = new_E5161_ | new_E5162_;
  assign new_E5158_ = new_E5101_ & new_E5115_;
  assign new_E5159_ = ~new_E5101_ & ~new_E5115_;
  assign new_E5160_ = new_E5101_ & ~new_E5115_;
  assign new_E5161_ = new_E5101_ & ~new_E5115_;
  assign new_E5162_ = ~new_E5101_ & new_E5115_;
  assign new_E5163_ = new_F7099_;
  assign new_E5164_ = new_F7166_;
  assign new_E5165_ = new_F7233_;
  assign new_E5166_ = new_F7300_;
  assign new_E5167_ = new_F7367_;
  assign new_E5168_ = new_F7434_;
  assign new_E5169_ = new_E5176_ & new_E5175_;
  assign new_E5170_ = new_E5178_ | new_E5177_;
  assign new_E5171_ = new_E5180_ | new_E5179_;
  assign new_E5172_ = new_E5182_ & new_E5181_;
  assign new_E5173_ = new_E5182_ & new_E5183_;
  assign new_E5174_ = new_E5175_ | new_E5184_;
  assign new_E5175_ = new_E5164_ | new_E5187_;
  assign new_E5176_ = new_E5186_ | new_E5185_;
  assign new_E5177_ = new_E5191_ & new_E5190_;
  assign new_E5178_ = new_E5189_ & new_E5188_;
  assign new_E5179_ = new_E5194_ | new_E5193_;
  assign new_E5180_ = new_E5189_ & new_E5192_;
  assign new_E5181_ = new_E5164_ | new_E5197_;
  assign new_E5182_ = new_E5196_ | new_E5195_;
  assign new_E5183_ = new_E5199_ | new_E5198_;
  assign new_E5184_ = ~new_E5175_ & new_E5201_;
  assign new_E5185_ = ~new_E5177_ & new_E5189_;
  assign new_E5186_ = new_E5177_ & ~new_E5189_;
  assign new_E5187_ = new_E5163_ & ~new_E5164_;
  assign new_E5188_ = ~new_E5210_ | ~new_E5211_;
  assign new_E5189_ = new_E5203_ | new_E5205_;
  assign new_E5190_ = new_E5213_ | new_E5212_;
  assign new_E5191_ = new_E5207_ | new_E5206_;
  assign new_E5192_ = ~new_E5215_ | ~new_E5214_;
  assign new_E5193_ = ~new_E5216_ & new_E5217_;
  assign new_E5194_ = new_E5216_ & ~new_E5217_;
  assign new_E5195_ = ~new_E5163_ & new_E5164_;
  assign new_E5196_ = new_E5163_ & ~new_E5164_;
  assign new_E5197_ = ~new_E5179_ | new_E5189_;
  assign new_E5198_ = new_E5179_ & new_E5189_;
  assign new_E5199_ = ~new_E5179_ & ~new_E5189_;
  assign new_E5200_ = new_E5221_ | new_E5220_;
  assign new_E5201_ = new_E5167_ | new_E5200_;
  assign new_E5202_ = new_E5225_ | new_E5224_;
  assign new_E5203_ = ~new_E5167_ & new_E5202_;
  assign new_E5204_ = new_E5223_ | new_E5222_;
  assign new_E5205_ = new_E5167_ & new_E5204_;
  assign new_E5206_ = new_E5165_ & ~new_E5175_;
  assign new_E5207_ = ~new_E5165_ & new_E5175_;
  assign new_E5208_ = ~new_E5164_ | ~new_E5189_;
  assign new_E5209_ = new_E5175_ & new_E5208_;
  assign new_E5210_ = ~new_E5175_ & ~new_E5209_;
  assign new_E5211_ = new_E5175_ | new_E5208_;
  assign new_E5212_ = ~new_E5165_ & new_E5166_;
  assign new_E5213_ = new_E5165_ & ~new_E5166_;
  assign new_E5214_ = new_E5182_ | new_E5219_;
  assign new_E5215_ = ~new_E5182_ & ~new_E5218_;
  assign new_E5216_ = new_E5165_ | new_E5182_;
  assign new_E5217_ = new_E5165_ | new_E5166_;
  assign new_E5218_ = new_E5182_ & new_E5219_;
  assign new_E5219_ = ~new_E5164_ | ~new_E5189_;
  assign new_E5220_ = new_E5197_ & new_E5217_;
  assign new_E5221_ = ~new_E5197_ & ~new_E5217_;
  assign new_E5222_ = new_E5226_ | new_E5227_;
  assign new_E5223_ = ~new_E5168_ & new_E5182_;
  assign new_E5224_ = new_E5228_ | new_E5229_;
  assign new_E5225_ = new_E5168_ & new_E5182_;
  assign new_E5226_ = ~new_E5168_ & ~new_E5182_;
  assign new_E5227_ = new_E5168_ & ~new_E5182_;
  assign new_E5228_ = new_E5168_ & ~new_E5182_;
  assign new_E5229_ = ~new_E5168_ & new_E5182_;
  assign new_E5230_ = new_F7501_;
  assign new_E5231_ = new_F7568_;
  assign new_E5232_ = new_F7635_;
  assign new_E5233_ = new_F7702_;
  assign new_E5234_ = new_F7769_;
  assign new_E5235_ = new_F7836_;
  assign new_E5236_ = new_E5243_ & new_E5242_;
  assign new_E5237_ = new_E5245_ | new_E5244_;
  assign new_E5238_ = new_E5247_ | new_E5246_;
  assign new_E5239_ = new_E5249_ & new_E5248_;
  assign new_E5240_ = new_E5249_ & new_E5250_;
  assign new_E5241_ = new_E5242_ | new_E5251_;
  assign new_E5242_ = new_E5231_ | new_E5254_;
  assign new_E5243_ = new_E5253_ | new_E5252_;
  assign new_E5244_ = new_E5258_ & new_E5257_;
  assign new_E5245_ = new_E5256_ & new_E5255_;
  assign new_E5246_ = new_E5261_ | new_E5260_;
  assign new_E5247_ = new_E5256_ & new_E5259_;
  assign new_E5248_ = new_E5231_ | new_E5264_;
  assign new_E5249_ = new_E5263_ | new_E5262_;
  assign new_E5250_ = new_E5266_ | new_E5265_;
  assign new_E5251_ = ~new_E5242_ & new_E5268_;
  assign new_E5252_ = ~new_E5244_ & new_E5256_;
  assign new_E5253_ = new_E5244_ & ~new_E5256_;
  assign new_E5254_ = new_E5230_ & ~new_E5231_;
  assign new_E5255_ = ~new_E5277_ | ~new_E5278_;
  assign new_E5256_ = new_E5270_ | new_E5272_;
  assign new_E5257_ = new_E5280_ | new_E5279_;
  assign new_E5258_ = new_E5274_ | new_E5273_;
  assign new_E5259_ = ~new_E5282_ | ~new_E5281_;
  assign new_E5260_ = ~new_E5283_ & new_E5284_;
  assign new_E5261_ = new_E5283_ & ~new_E5284_;
  assign new_E5262_ = ~new_E5230_ & new_E5231_;
  assign new_E5263_ = new_E5230_ & ~new_E5231_;
  assign new_E5264_ = ~new_E5246_ | new_E5256_;
  assign new_E5265_ = new_E5246_ & new_E5256_;
  assign new_E5266_ = ~new_E5246_ & ~new_E5256_;
  assign new_E5267_ = new_E5288_ | new_E5287_;
  assign new_E5268_ = new_E5234_ | new_E5267_;
  assign new_E5269_ = new_E5292_ | new_E5291_;
  assign new_E5270_ = ~new_E5234_ & new_E5269_;
  assign new_E5271_ = new_E5290_ | new_E5289_;
  assign new_E5272_ = new_E5234_ & new_E5271_;
  assign new_E5273_ = new_E5232_ & ~new_E5242_;
  assign new_E5274_ = ~new_E5232_ & new_E5242_;
  assign new_E5275_ = ~new_E5231_ | ~new_E5256_;
  assign new_E5276_ = new_E5242_ & new_E5275_;
  assign new_E5277_ = ~new_E5242_ & ~new_E5276_;
  assign new_E5278_ = new_E5242_ | new_E5275_;
  assign new_E5279_ = ~new_E5232_ & new_E5233_;
  assign new_E5280_ = new_E5232_ & ~new_E5233_;
  assign new_E5281_ = new_E5249_ | new_E5286_;
  assign new_E5282_ = ~new_E5249_ & ~new_E5285_;
  assign new_E5283_ = new_E5232_ | new_E5249_;
  assign new_E5284_ = new_E5232_ | new_E5233_;
  assign new_E5285_ = new_E5249_ & new_E5286_;
  assign new_E5286_ = ~new_E5231_ | ~new_E5256_;
  assign new_E5287_ = new_E5264_ & new_E5284_;
  assign new_E5288_ = ~new_E5264_ & ~new_E5284_;
  assign new_E5289_ = new_E5293_ | new_E5294_;
  assign new_E5290_ = ~new_E5235_ & new_E5249_;
  assign new_E5291_ = new_E5295_ | new_E5296_;
  assign new_E5292_ = new_E5235_ & new_E5249_;
  assign new_E5293_ = ~new_E5235_ & ~new_E5249_;
  assign new_E5294_ = new_E5235_ & ~new_E5249_;
  assign new_E5295_ = new_E5235_ & ~new_E5249_;
  assign new_E5296_ = ~new_E5235_ & new_E5249_;
  assign new_E5297_ = new_F7903_;
  assign new_E5298_ = new_F7970_;
  assign new_E5299_ = new_F8037_;
  assign new_E5300_ = new_F8104_;
  assign new_E5301_ = new_F8171_;
  assign new_E5302_ = new_F8238_;
  assign new_E5303_ = new_E5310_ & new_E5309_;
  assign new_E5304_ = new_E5312_ | new_E5311_;
  assign new_E5305_ = new_E5314_ | new_E5313_;
  assign new_E5306_ = new_E5316_ & new_E5315_;
  assign new_E5307_ = new_E5316_ & new_E5317_;
  assign new_E5308_ = new_E5309_ | new_E5318_;
  assign new_E5309_ = new_E5298_ | new_E5321_;
  assign new_E5310_ = new_E5320_ | new_E5319_;
  assign new_E5311_ = new_E5325_ & new_E5324_;
  assign new_E5312_ = new_E5323_ & new_E5322_;
  assign new_E5313_ = new_E5328_ | new_E5327_;
  assign new_E5314_ = new_E5323_ & new_E5326_;
  assign new_E5315_ = new_E5298_ | new_E5331_;
  assign new_E5316_ = new_E5330_ | new_E5329_;
  assign new_E5317_ = new_E5333_ | new_E5332_;
  assign new_E5318_ = ~new_E5309_ & new_E5335_;
  assign new_E5319_ = ~new_E5311_ & new_E5323_;
  assign new_E5320_ = new_E5311_ & ~new_E5323_;
  assign new_E5321_ = new_E5297_ & ~new_E5298_;
  assign new_E5322_ = ~new_E5344_ | ~new_E5345_;
  assign new_E5323_ = new_E5337_ | new_E5339_;
  assign new_E5324_ = new_E5347_ | new_E5346_;
  assign new_E5325_ = new_E5341_ | new_E5340_;
  assign new_E5326_ = ~new_E5349_ | ~new_E5348_;
  assign new_E5327_ = ~new_E5350_ & new_E5351_;
  assign new_E5328_ = new_E5350_ & ~new_E5351_;
  assign new_E5329_ = ~new_E5297_ & new_E5298_;
  assign new_E5330_ = new_E5297_ & ~new_E5298_;
  assign new_E5331_ = ~new_E5313_ | new_E5323_;
  assign new_E5332_ = new_E5313_ & new_E5323_;
  assign new_E5333_ = ~new_E5313_ & ~new_E5323_;
  assign new_E5334_ = new_E5355_ | new_E5354_;
  assign new_E5335_ = new_E5301_ | new_E5334_;
  assign new_E5336_ = new_E5359_ | new_E5358_;
  assign new_E5337_ = ~new_E5301_ & new_E5336_;
  assign new_E5338_ = new_E5357_ | new_E5356_;
  assign new_E5339_ = new_E5301_ & new_E5338_;
  assign new_E5340_ = new_E5299_ & ~new_E5309_;
  assign new_E5341_ = ~new_E5299_ & new_E5309_;
  assign new_E5342_ = ~new_E5298_ | ~new_E5323_;
  assign new_E5343_ = new_E5309_ & new_E5342_;
  assign new_E5344_ = ~new_E5309_ & ~new_E5343_;
  assign new_E5345_ = new_E5309_ | new_E5342_;
  assign new_E5346_ = ~new_E5299_ & new_E5300_;
  assign new_E5347_ = new_E5299_ & ~new_E5300_;
  assign new_E5348_ = new_E5316_ | new_E5353_;
  assign new_E5349_ = ~new_E5316_ & ~new_E5352_;
  assign new_E5350_ = new_E5299_ | new_E5316_;
  assign new_E5351_ = new_E5299_ | new_E5300_;
  assign new_E5352_ = new_E5316_ & new_E5353_;
  assign new_E5353_ = ~new_E5298_ | ~new_E5323_;
  assign new_E5354_ = new_E5331_ & new_E5351_;
  assign new_E5355_ = ~new_E5331_ & ~new_E5351_;
  assign new_E5356_ = new_E5360_ | new_E5361_;
  assign new_E5357_ = ~new_E5302_ & new_E5316_;
  assign new_E5358_ = new_E5362_ | new_E5363_;
  assign new_E5359_ = new_E5302_ & new_E5316_;
  assign new_E5360_ = ~new_E5302_ & ~new_E5316_;
  assign new_E5361_ = new_E5302_ & ~new_E5316_;
  assign new_E5362_ = new_E5302_ & ~new_E5316_;
  assign new_E5363_ = ~new_E5302_ & new_E5316_;
  assign new_E5364_ = new_F8305_;
  assign new_E5365_ = new_F8372_;
  assign new_E5366_ = new_F8439_;
  assign new_E5367_ = new_F8506_;
  assign new_E5368_ = new_F8573_;
  assign new_E5369_ = new_F8640_;
  assign new_E5370_ = new_E5377_ & new_E5376_;
  assign new_E5371_ = new_E5379_ | new_E5378_;
  assign new_E5372_ = new_E5381_ | new_E5380_;
  assign new_E5373_ = new_E5383_ & new_E5382_;
  assign new_E5374_ = new_E5383_ & new_E5384_;
  assign new_E5375_ = new_E5376_ | new_E5385_;
  assign new_E5376_ = new_E5365_ | new_E5388_;
  assign new_E5377_ = new_E5387_ | new_E5386_;
  assign new_E5378_ = new_E5392_ & new_E5391_;
  assign new_E5379_ = new_E5390_ & new_E5389_;
  assign new_E5380_ = new_E5395_ | new_E5394_;
  assign new_E5381_ = new_E5390_ & new_E5393_;
  assign new_E5382_ = new_E5365_ | new_E5398_;
  assign new_E5383_ = new_E5397_ | new_E5396_;
  assign new_E5384_ = new_E5400_ | new_E5399_;
  assign new_E5385_ = ~new_E5376_ & new_E5402_;
  assign new_E5386_ = ~new_E5378_ & new_E5390_;
  assign new_E5387_ = new_E5378_ & ~new_E5390_;
  assign new_E5388_ = new_E5364_ & ~new_E5365_;
  assign new_E5389_ = ~new_E5411_ | ~new_E5412_;
  assign new_E5390_ = new_E5404_ | new_E5406_;
  assign new_E5391_ = new_E5414_ | new_E5413_;
  assign new_E5392_ = new_E5408_ | new_E5407_;
  assign new_E5393_ = ~new_E5416_ | ~new_E5415_;
  assign new_E5394_ = ~new_E5417_ & new_E5418_;
  assign new_E5395_ = new_E5417_ & ~new_E5418_;
  assign new_E5396_ = ~new_E5364_ & new_E5365_;
  assign new_E5397_ = new_E5364_ & ~new_E5365_;
  assign new_E5398_ = ~new_E5380_ | new_E5390_;
  assign new_E5399_ = new_E5380_ & new_E5390_;
  assign new_E5400_ = ~new_E5380_ & ~new_E5390_;
  assign new_E5401_ = new_E5422_ | new_E5421_;
  assign new_E5402_ = new_E5368_ | new_E5401_;
  assign new_E5403_ = new_E5426_ | new_E5425_;
  assign new_E5404_ = ~new_E5368_ & new_E5403_;
  assign new_E5405_ = new_E5424_ | new_E5423_;
  assign new_E5406_ = new_E5368_ & new_E5405_;
  assign new_E5407_ = new_E5366_ & ~new_E5376_;
  assign new_E5408_ = ~new_E5366_ & new_E5376_;
  assign new_E5409_ = ~new_E5365_ | ~new_E5390_;
  assign new_E5410_ = new_E5376_ & new_E5409_;
  assign new_E5411_ = ~new_E5376_ & ~new_E5410_;
  assign new_E5412_ = new_E5376_ | new_E5409_;
  assign new_E5413_ = ~new_E5366_ & new_E5367_;
  assign new_E5414_ = new_E5366_ & ~new_E5367_;
  assign new_E5415_ = new_E5383_ | new_E5420_;
  assign new_E5416_ = ~new_E5383_ & ~new_E5419_;
  assign new_E5417_ = new_E5366_ | new_E5383_;
  assign new_E5418_ = new_E5366_ | new_E5367_;
  assign new_E5419_ = new_E5383_ & new_E5420_;
  assign new_E5420_ = ~new_E5365_ | ~new_E5390_;
  assign new_E5421_ = new_E5398_ & new_E5418_;
  assign new_E5422_ = ~new_E5398_ & ~new_E5418_;
  assign new_E5423_ = new_E5427_ | new_E5428_;
  assign new_E5424_ = ~new_E5369_ & new_E5383_;
  assign new_E5425_ = new_E5429_ | new_E5430_;
  assign new_E5426_ = new_E5369_ & new_E5383_;
  assign new_E5427_ = ~new_E5369_ & ~new_E5383_;
  assign new_E5428_ = new_E5369_ & ~new_E5383_;
  assign new_E5429_ = new_E5369_ & ~new_E5383_;
  assign new_E5430_ = ~new_E5369_ & new_E5383_;
  assign new_E5431_ = new_F8707_;
  assign new_E5432_ = new_F8774_;
  assign new_E5433_ = new_F8841_;
  assign new_E5434_ = new_F8908_;
  assign new_E5435_ = new_F8975_;
  assign new_E5436_ = new_F9042_;
  assign new_E5437_ = new_E5444_ & new_E5443_;
  assign new_E5438_ = new_E5446_ | new_E5445_;
  assign new_E5439_ = new_E5448_ | new_E5447_;
  assign new_E5440_ = new_E5450_ & new_E5449_;
  assign new_E5441_ = new_E5450_ & new_E5451_;
  assign new_E5442_ = new_E5443_ | new_E5452_;
  assign new_E5443_ = new_E5432_ | new_E5455_;
  assign new_E5444_ = new_E5454_ | new_E5453_;
  assign new_E5445_ = new_E5459_ & new_E5458_;
  assign new_E5446_ = new_E5457_ & new_E5456_;
  assign new_E5447_ = new_E5462_ | new_E5461_;
  assign new_E5448_ = new_E5457_ & new_E5460_;
  assign new_E5449_ = new_E5432_ | new_E5465_;
  assign new_E5450_ = new_E5464_ | new_E5463_;
  assign new_E5451_ = new_E5467_ | new_E5466_;
  assign new_E5452_ = ~new_E5443_ & new_E5469_;
  assign new_E5453_ = ~new_E5445_ & new_E5457_;
  assign new_E5454_ = new_E5445_ & ~new_E5457_;
  assign new_E5455_ = new_E5431_ & ~new_E5432_;
  assign new_E5456_ = ~new_E5478_ | ~new_E5479_;
  assign new_E5457_ = new_E5471_ | new_E5473_;
  assign new_E5458_ = new_E5481_ | new_E5480_;
  assign new_E5459_ = new_E5475_ | new_E5474_;
  assign new_E5460_ = ~new_E5483_ | ~new_E5482_;
  assign new_E5461_ = ~new_E5484_ & new_E5485_;
  assign new_E5462_ = new_E5484_ & ~new_E5485_;
  assign new_E5463_ = ~new_E5431_ & new_E5432_;
  assign new_E5464_ = new_E5431_ & ~new_E5432_;
  assign new_E5465_ = ~new_E5447_ | new_E5457_;
  assign new_E5466_ = new_E5447_ & new_E5457_;
  assign new_E5467_ = ~new_E5447_ & ~new_E5457_;
  assign new_E5468_ = new_E5489_ | new_E5488_;
  assign new_E5469_ = new_E5435_ | new_E5468_;
  assign new_E5470_ = new_E5493_ | new_E5492_;
  assign new_E5471_ = ~new_E5435_ & new_E5470_;
  assign new_E5472_ = new_E5491_ | new_E5490_;
  assign new_E5473_ = new_E5435_ & new_E5472_;
  assign new_E5474_ = new_E5433_ & ~new_E5443_;
  assign new_E5475_ = ~new_E5433_ & new_E5443_;
  assign new_E5476_ = ~new_E5432_ | ~new_E5457_;
  assign new_E5477_ = new_E5443_ & new_E5476_;
  assign new_E5478_ = ~new_E5443_ & ~new_E5477_;
  assign new_E5479_ = new_E5443_ | new_E5476_;
  assign new_E5480_ = ~new_E5433_ & new_E5434_;
  assign new_E5481_ = new_E5433_ & ~new_E5434_;
  assign new_E5482_ = new_E5450_ | new_E5487_;
  assign new_E5483_ = ~new_E5450_ & ~new_E5486_;
  assign new_E5484_ = new_E5433_ | new_E5450_;
  assign new_E5485_ = new_E5433_ | new_E5434_;
  assign new_E5486_ = new_E5450_ & new_E5487_;
  assign new_E5487_ = ~new_E5432_ | ~new_E5457_;
  assign new_E5488_ = new_E5465_ & new_E5485_;
  assign new_E5489_ = ~new_E5465_ & ~new_E5485_;
  assign new_E5490_ = new_E5494_ | new_E5495_;
  assign new_E5491_ = ~new_E5436_ & new_E5450_;
  assign new_E5492_ = new_E5496_ | new_E5497_;
  assign new_E5493_ = new_E5436_ & new_E5450_;
  assign new_E5494_ = ~new_E5436_ & ~new_E5450_;
  assign new_E5495_ = new_E5436_ & ~new_E5450_;
  assign new_E5496_ = new_E5436_ & ~new_E5450_;
  assign new_E5497_ = ~new_E5436_ & new_E5450_;
  assign new_E5498_ = new_F9109_;
  assign new_E5499_ = new_F9176_;
  assign new_E5500_ = new_F9243_;
  assign new_E5501_ = new_F9310_;
  assign new_E5502_ = new_F9377_;
  assign new_E5503_ = new_F9444_;
  assign new_E5504_ = new_E5511_ & new_E5510_;
  assign new_E5505_ = new_E5513_ | new_E5512_;
  assign new_E5506_ = new_E5515_ | new_E5514_;
  assign new_E5507_ = new_E5517_ & new_E5516_;
  assign new_E5508_ = new_E5517_ & new_E5518_;
  assign new_E5509_ = new_E5510_ | new_E5519_;
  assign new_E5510_ = new_E5499_ | new_E5522_;
  assign new_E5511_ = new_E5521_ | new_E5520_;
  assign new_E5512_ = new_E5526_ & new_E5525_;
  assign new_E5513_ = new_E5524_ & new_E5523_;
  assign new_E5514_ = new_E5529_ | new_E5528_;
  assign new_E5515_ = new_E5524_ & new_E5527_;
  assign new_E5516_ = new_E5499_ | new_E5532_;
  assign new_E5517_ = new_E5531_ | new_E5530_;
  assign new_E5518_ = new_E5534_ | new_E5533_;
  assign new_E5519_ = ~new_E5510_ & new_E5536_;
  assign new_E5520_ = ~new_E5512_ & new_E5524_;
  assign new_E5521_ = new_E5512_ & ~new_E5524_;
  assign new_E5522_ = new_E5498_ & ~new_E5499_;
  assign new_E5523_ = ~new_E5545_ | ~new_E5546_;
  assign new_E5524_ = new_E5538_ | new_E5540_;
  assign new_E5525_ = new_E5548_ | new_E5547_;
  assign new_E5526_ = new_E5542_ | new_E5541_;
  assign new_E5527_ = ~new_E5550_ | ~new_E5549_;
  assign new_E5528_ = ~new_E5551_ & new_E5552_;
  assign new_E5529_ = new_E5551_ & ~new_E5552_;
  assign new_E5530_ = ~new_E5498_ & new_E5499_;
  assign new_E5531_ = new_E5498_ & ~new_E5499_;
  assign new_E5532_ = ~new_E5514_ | new_E5524_;
  assign new_E5533_ = new_E5514_ & new_E5524_;
  assign new_E5534_ = ~new_E5514_ & ~new_E5524_;
  assign new_E5535_ = new_E5556_ | new_E5555_;
  assign new_E5536_ = new_E5502_ | new_E5535_;
  assign new_E5537_ = new_E5560_ | new_E5559_;
  assign new_E5538_ = ~new_E5502_ & new_E5537_;
  assign new_E5539_ = new_E5558_ | new_E5557_;
  assign new_E5540_ = new_E5502_ & new_E5539_;
  assign new_E5541_ = new_E5500_ & ~new_E5510_;
  assign new_E5542_ = ~new_E5500_ & new_E5510_;
  assign new_E5543_ = ~new_E5499_ | ~new_E5524_;
  assign new_E5544_ = new_E5510_ & new_E5543_;
  assign new_E5545_ = ~new_E5510_ & ~new_E5544_;
  assign new_E5546_ = new_E5510_ | new_E5543_;
  assign new_E5547_ = ~new_E5500_ & new_E5501_;
  assign new_E5548_ = new_E5500_ & ~new_E5501_;
  assign new_E5549_ = new_E5517_ | new_E5554_;
  assign new_E5550_ = ~new_E5517_ & ~new_E5553_;
  assign new_E5551_ = new_E5500_ | new_E5517_;
  assign new_E5552_ = new_E5500_ | new_E5501_;
  assign new_E5553_ = new_E5517_ & new_E5554_;
  assign new_E5554_ = ~new_E5499_ | ~new_E5524_;
  assign new_E5555_ = new_E5532_ & new_E5552_;
  assign new_E5556_ = ~new_E5532_ & ~new_E5552_;
  assign new_E5557_ = new_E5561_ | new_E5562_;
  assign new_E5558_ = ~new_E5503_ & new_E5517_;
  assign new_E5559_ = new_E5563_ | new_E5564_;
  assign new_E5560_ = new_E5503_ & new_E5517_;
  assign new_E5561_ = ~new_E5503_ & ~new_E5517_;
  assign new_E5562_ = new_E5503_ & ~new_E5517_;
  assign new_E5563_ = new_E5503_ & ~new_E5517_;
  assign new_E5564_ = ~new_E5503_ & new_E5517_;
  assign new_E5565_ = new_F9511_;
  assign new_E5566_ = new_F9578_;
  assign new_E5567_ = new_F9645_;
  assign new_E5568_ = new_F9712_;
  assign new_E5569_ = new_F9779_;
  assign new_E5570_ = new_F9846_;
  assign new_E5571_ = new_E5578_ & new_E5577_;
  assign new_E5572_ = new_E5580_ | new_E5579_;
  assign new_E5573_ = new_E5582_ | new_E5581_;
  assign new_E5574_ = new_E5584_ & new_E5583_;
  assign new_E5575_ = new_E5584_ & new_E5585_;
  assign new_E5576_ = new_E5577_ | new_E5586_;
  assign new_E5577_ = new_E5566_ | new_E5589_;
  assign new_E5578_ = new_E5588_ | new_E5587_;
  assign new_E5579_ = new_E5593_ & new_E5592_;
  assign new_E5580_ = new_E5591_ & new_E5590_;
  assign new_E5581_ = new_E5596_ | new_E5595_;
  assign new_E5582_ = new_E5591_ & new_E5594_;
  assign new_E5583_ = new_E5566_ | new_E5599_;
  assign new_E5584_ = new_E5598_ | new_E5597_;
  assign new_E5585_ = new_E5601_ | new_E5600_;
  assign new_E5586_ = ~new_E5577_ & new_E5603_;
  assign new_E5587_ = ~new_E5579_ & new_E5591_;
  assign new_E5588_ = new_E5579_ & ~new_E5591_;
  assign new_E5589_ = new_E5565_ & ~new_E5566_;
  assign new_E5590_ = ~new_E5612_ | ~new_E5613_;
  assign new_E5591_ = new_E5605_ | new_E5607_;
  assign new_E5592_ = new_E5615_ | new_E5614_;
  assign new_E5593_ = new_E5609_ | new_E5608_;
  assign new_E5594_ = ~new_E5617_ | ~new_E5616_;
  assign new_E5595_ = ~new_E5618_ & new_E5619_;
  assign new_E5596_ = new_E5618_ & ~new_E5619_;
  assign new_E5597_ = ~new_E5565_ & new_E5566_;
  assign new_E5598_ = new_E5565_ & ~new_E5566_;
  assign new_E5599_ = ~new_E5581_ | new_E5591_;
  assign new_E5600_ = new_E5581_ & new_E5591_;
  assign new_E5601_ = ~new_E5581_ & ~new_E5591_;
  assign new_E5602_ = new_E5623_ | new_E5622_;
  assign new_E5603_ = new_E5569_ | new_E5602_;
  assign new_E5604_ = new_E5627_ | new_E5626_;
  assign new_E5605_ = ~new_E5569_ & new_E5604_;
  assign new_E5606_ = new_E5625_ | new_E5624_;
  assign new_E5607_ = new_E5569_ & new_E5606_;
  assign new_E5608_ = new_E5567_ & ~new_E5577_;
  assign new_E5609_ = ~new_E5567_ & new_E5577_;
  assign new_E5610_ = ~new_E5566_ | ~new_E5591_;
  assign new_E5611_ = new_E5577_ & new_E5610_;
  assign new_E5612_ = ~new_E5577_ & ~new_E5611_;
  assign new_E5613_ = new_E5577_ | new_E5610_;
  assign new_E5614_ = ~new_E5567_ & new_E5568_;
  assign new_E5615_ = new_E5567_ & ~new_E5568_;
  assign new_E5616_ = new_E5584_ | new_E5621_;
  assign new_E5617_ = ~new_E5584_ & ~new_E5620_;
  assign new_E5618_ = new_E5567_ | new_E5584_;
  assign new_E5619_ = new_E5567_ | new_E5568_;
  assign new_E5620_ = new_E5584_ & new_E5621_;
  assign new_E5621_ = ~new_E5566_ | ~new_E5591_;
  assign new_E5622_ = new_E5599_ & new_E5619_;
  assign new_E5623_ = ~new_E5599_ & ~new_E5619_;
  assign new_E5624_ = new_E5628_ | new_E5629_;
  assign new_E5625_ = ~new_E5570_ & new_E5584_;
  assign new_E5626_ = new_E5630_ | new_E5631_;
  assign new_E5627_ = new_E5570_ & new_E5584_;
  assign new_E5628_ = ~new_E5570_ & ~new_E5584_;
  assign new_E5629_ = new_E5570_ & ~new_E5584_;
  assign new_E5630_ = new_E5570_ & ~new_E5584_;
  assign new_E5631_ = ~new_E5570_ & new_E5584_;
  assign new_E5632_ = new_F9913_;
  assign new_E5633_ = new_F9980_;
  assign new_E5634_ = new_G48_;
  assign new_E5635_ = new_G115_;
  assign new_E5636_ = new_G182_;
  assign new_E5637_ = new_G249_;
  assign new_E5638_ = new_E5645_ & new_E5644_;
  assign new_E5639_ = new_E5647_ | new_E5646_;
  assign new_E5640_ = new_E5649_ | new_E5648_;
  assign new_E5641_ = new_E5651_ & new_E5650_;
  assign new_E5642_ = new_E5651_ & new_E5652_;
  assign new_E5643_ = new_E5644_ | new_E5653_;
  assign new_E5644_ = new_E5633_ | new_E5656_;
  assign new_E5645_ = new_E5655_ | new_E5654_;
  assign new_E5646_ = new_E5660_ & new_E5659_;
  assign new_E5647_ = new_E5658_ & new_E5657_;
  assign new_E5648_ = new_E5663_ | new_E5662_;
  assign new_E5649_ = new_E5658_ & new_E5661_;
  assign new_E5650_ = new_E5633_ | new_E5666_;
  assign new_E5651_ = new_E5665_ | new_E5664_;
  assign new_E5652_ = new_E5668_ | new_E5667_;
  assign new_E5653_ = ~new_E5644_ & new_E5670_;
  assign new_E5654_ = ~new_E5646_ & new_E5658_;
  assign new_E5655_ = new_E5646_ & ~new_E5658_;
  assign new_E5656_ = new_E5632_ & ~new_E5633_;
  assign new_E5657_ = ~new_E5679_ | ~new_E5680_;
  assign new_E5658_ = new_E5672_ | new_E5674_;
  assign new_E5659_ = new_E5682_ | new_E5681_;
  assign new_E5660_ = new_E5676_ | new_E5675_;
  assign new_E5661_ = ~new_E5684_ | ~new_E5683_;
  assign new_E5662_ = ~new_E5685_ & new_E5686_;
  assign new_E5663_ = new_E5685_ & ~new_E5686_;
  assign new_E5664_ = ~new_E5632_ & new_E5633_;
  assign new_E5665_ = new_E5632_ & ~new_E5633_;
  assign new_E5666_ = ~new_E5648_ | new_E5658_;
  assign new_E5667_ = new_E5648_ & new_E5658_;
  assign new_E5668_ = ~new_E5648_ & ~new_E5658_;
  assign new_E5669_ = new_E5690_ | new_E5689_;
  assign new_E5670_ = new_E5636_ | new_E5669_;
  assign new_E5671_ = new_E5694_ | new_E5693_;
  assign new_E5672_ = ~new_E5636_ & new_E5671_;
  assign new_E5673_ = new_E5692_ | new_E5691_;
  assign new_E5674_ = new_E5636_ & new_E5673_;
  assign new_E5675_ = new_E5634_ & ~new_E5644_;
  assign new_E5676_ = ~new_E5634_ & new_E5644_;
  assign new_E5677_ = ~new_E5633_ | ~new_E5658_;
  assign new_E5678_ = new_E5644_ & new_E5677_;
  assign new_E5679_ = ~new_E5644_ & ~new_E5678_;
  assign new_E5680_ = new_E5644_ | new_E5677_;
  assign new_E5681_ = ~new_E5634_ & new_E5635_;
  assign new_E5682_ = new_E5634_ & ~new_E5635_;
  assign new_E5683_ = new_E5651_ | new_E5688_;
  assign new_E5684_ = ~new_E5651_ & ~new_E5687_;
  assign new_E5685_ = new_E5634_ | new_E5651_;
  assign new_E5686_ = new_E5634_ | new_E5635_;
  assign new_E5687_ = new_E5651_ & new_E5688_;
  assign new_E5688_ = ~new_E5633_ | ~new_E5658_;
  assign new_E5689_ = new_E5666_ & new_E5686_;
  assign new_E5690_ = ~new_E5666_ & ~new_E5686_;
  assign new_E5691_ = new_E5695_ | new_E5696_;
  assign new_E5692_ = ~new_E5637_ & new_E5651_;
  assign new_E5693_ = new_E5697_ | new_E5698_;
  assign new_E5694_ = new_E5637_ & new_E5651_;
  assign new_E5695_ = ~new_E5637_ & ~new_E5651_;
  assign new_E5696_ = new_E5637_ & ~new_E5651_;
  assign new_E5697_ = new_E5637_ & ~new_E5651_;
  assign new_E5698_ = ~new_E5637_ & new_E5651_;
  assign new_E5699_ = new_G316_;
  assign new_E5700_ = new_G383_;
  assign new_E5701_ = new_G450_;
  assign new_E5702_ = new_G517_;
  assign new_E5703_ = new_G584_;
  assign new_E5704_ = new_G651_;
  assign new_E5705_ = new_E5712_ & new_E5711_;
  assign new_E5706_ = new_E5714_ | new_E5713_;
  assign new_E5707_ = new_E5716_ | new_E5715_;
  assign new_E5708_ = new_E5718_ & new_E5717_;
  assign new_E5709_ = new_E5718_ & new_E5719_;
  assign new_E5710_ = new_E5711_ | new_E5720_;
  assign new_E5711_ = new_E5700_ | new_E5723_;
  assign new_E5712_ = new_E5722_ | new_E5721_;
  assign new_E5713_ = new_E5727_ & new_E5726_;
  assign new_E5714_ = new_E5725_ & new_E5724_;
  assign new_E5715_ = new_E5730_ | new_E5729_;
  assign new_E5716_ = new_E5725_ & new_E5728_;
  assign new_E5717_ = new_E5700_ | new_E5733_;
  assign new_E5718_ = new_E5732_ | new_E5731_;
  assign new_E5719_ = new_E5735_ | new_E5734_;
  assign new_E5720_ = ~new_E5711_ & new_E5737_;
  assign new_E5721_ = ~new_E5713_ & new_E5725_;
  assign new_E5722_ = new_E5713_ & ~new_E5725_;
  assign new_E5723_ = new_E5699_ & ~new_E5700_;
  assign new_E5724_ = ~new_E5746_ | ~new_E5747_;
  assign new_E5725_ = new_E5739_ | new_E5741_;
  assign new_E5726_ = new_E5749_ | new_E5748_;
  assign new_E5727_ = new_E5743_ | new_E5742_;
  assign new_E5728_ = ~new_E5751_ | ~new_E5750_;
  assign new_E5729_ = ~new_E5752_ & new_E5753_;
  assign new_E5730_ = new_E5752_ & ~new_E5753_;
  assign new_E5731_ = ~new_E5699_ & new_E5700_;
  assign new_E5732_ = new_E5699_ & ~new_E5700_;
  assign new_E5733_ = ~new_E5715_ | new_E5725_;
  assign new_E5734_ = new_E5715_ & new_E5725_;
  assign new_E5735_ = ~new_E5715_ & ~new_E5725_;
  assign new_E5736_ = new_E5757_ | new_E5756_;
  assign new_E5737_ = new_E5703_ | new_E5736_;
  assign new_E5738_ = new_E5761_ | new_E5760_;
  assign new_E5739_ = ~new_E5703_ & new_E5738_;
  assign new_E5740_ = new_E5759_ | new_E5758_;
  assign new_E5741_ = new_E5703_ & new_E5740_;
  assign new_E5742_ = new_E5701_ & ~new_E5711_;
  assign new_E5743_ = ~new_E5701_ & new_E5711_;
  assign new_E5744_ = ~new_E5700_ | ~new_E5725_;
  assign new_E5745_ = new_E5711_ & new_E5744_;
  assign new_E5746_ = ~new_E5711_ & ~new_E5745_;
  assign new_E5747_ = new_E5711_ | new_E5744_;
  assign new_E5748_ = ~new_E5701_ & new_E5702_;
  assign new_E5749_ = new_E5701_ & ~new_E5702_;
  assign new_E5750_ = new_E5718_ | new_E5755_;
  assign new_E5751_ = ~new_E5718_ & ~new_E5754_;
  assign new_E5752_ = new_E5701_ | new_E5718_;
  assign new_E5753_ = new_E5701_ | new_E5702_;
  assign new_E5754_ = new_E5718_ & new_E5755_;
  assign new_E5755_ = ~new_E5700_ | ~new_E5725_;
  assign new_E5756_ = new_E5733_ & new_E5753_;
  assign new_E5757_ = ~new_E5733_ & ~new_E5753_;
  assign new_E5758_ = new_E5762_ | new_E5763_;
  assign new_E5759_ = ~new_E5704_ & new_E5718_;
  assign new_E5760_ = new_E5764_ | new_E5765_;
  assign new_E5761_ = new_E5704_ & new_E5718_;
  assign new_E5762_ = ~new_E5704_ & ~new_E5718_;
  assign new_E5763_ = new_E5704_ & ~new_E5718_;
  assign new_E5764_ = new_E5704_ & ~new_E5718_;
  assign new_E5765_ = ~new_E5704_ & new_E5718_;
  assign new_E5766_ = new_G718_;
  assign new_E5767_ = new_G785_;
  assign new_E5768_ = new_G852_;
  assign new_E5769_ = new_G919_;
  assign new_E5770_ = new_G986_;
  assign new_E5771_ = new_G1053_;
  assign new_E5772_ = new_E5779_ & new_E5778_;
  assign new_E5773_ = new_E5781_ | new_E5780_;
  assign new_E5774_ = new_E5783_ | new_E5782_;
  assign new_E5775_ = new_E5785_ & new_E5784_;
  assign new_E5776_ = new_E5785_ & new_E5786_;
  assign new_E5777_ = new_E5778_ | new_E5787_;
  assign new_E5778_ = new_E5767_ | new_E5790_;
  assign new_E5779_ = new_E5789_ | new_E5788_;
  assign new_E5780_ = new_E5794_ & new_E5793_;
  assign new_E5781_ = new_E5792_ & new_E5791_;
  assign new_E5782_ = new_E5797_ | new_E5796_;
  assign new_E5783_ = new_E5792_ & new_E5795_;
  assign new_E5784_ = new_E5767_ | new_E5800_;
  assign new_E5785_ = new_E5799_ | new_E5798_;
  assign new_E5786_ = new_E5802_ | new_E5801_;
  assign new_E5787_ = ~new_E5778_ & new_E5804_;
  assign new_E5788_ = ~new_E5780_ & new_E5792_;
  assign new_E5789_ = new_E5780_ & ~new_E5792_;
  assign new_E5790_ = new_E5766_ & ~new_E5767_;
  assign new_E5791_ = ~new_E5813_ | ~new_E5814_;
  assign new_E5792_ = new_E5806_ | new_E5808_;
  assign new_E5793_ = new_E5816_ | new_E5815_;
  assign new_E5794_ = new_E5810_ | new_E5809_;
  assign new_E5795_ = ~new_E5818_ | ~new_E5817_;
  assign new_E5796_ = ~new_E5819_ & new_E5820_;
  assign new_E5797_ = new_E5819_ & ~new_E5820_;
  assign new_E5798_ = ~new_E5766_ & new_E5767_;
  assign new_E5799_ = new_E5766_ & ~new_E5767_;
  assign new_E5800_ = ~new_E5782_ | new_E5792_;
  assign new_E5801_ = new_E5782_ & new_E5792_;
  assign new_E5802_ = ~new_E5782_ & ~new_E5792_;
  assign new_E5803_ = new_E5824_ | new_E5823_;
  assign new_E5804_ = new_E5770_ | new_E5803_;
  assign new_E5805_ = new_E5828_ | new_E5827_;
  assign new_E5806_ = ~new_E5770_ & new_E5805_;
  assign new_E5807_ = new_E5826_ | new_E5825_;
  assign new_E5808_ = new_E5770_ & new_E5807_;
  assign new_E5809_ = new_E5768_ & ~new_E5778_;
  assign new_E5810_ = ~new_E5768_ & new_E5778_;
  assign new_E5811_ = ~new_E5767_ | ~new_E5792_;
  assign new_E5812_ = new_E5778_ & new_E5811_;
  assign new_E5813_ = ~new_E5778_ & ~new_E5812_;
  assign new_E5814_ = new_E5778_ | new_E5811_;
  assign new_E5815_ = ~new_E5768_ & new_E5769_;
  assign new_E5816_ = new_E5768_ & ~new_E5769_;
  assign new_E5817_ = new_E5785_ | new_E5822_;
  assign new_E5818_ = ~new_E5785_ & ~new_E5821_;
  assign new_E5819_ = new_E5768_ | new_E5785_;
  assign new_E5820_ = new_E5768_ | new_E5769_;
  assign new_E5821_ = new_E5785_ & new_E5822_;
  assign new_E5822_ = ~new_E5767_ | ~new_E5792_;
  assign new_E5823_ = new_E5800_ & new_E5820_;
  assign new_E5824_ = ~new_E5800_ & ~new_E5820_;
  assign new_E5825_ = new_E5829_ | new_E5830_;
  assign new_E5826_ = ~new_E5771_ & new_E5785_;
  assign new_E5827_ = new_E5831_ | new_E5832_;
  assign new_E5828_ = new_E5771_ & new_E5785_;
  assign new_E5829_ = ~new_E5771_ & ~new_E5785_;
  assign new_E5830_ = new_E5771_ & ~new_E5785_;
  assign new_E5831_ = new_E5771_ & ~new_E5785_;
  assign new_E5832_ = ~new_E5771_ & new_E5785_;
  assign new_E5833_ = new_G1120_;
  assign new_E5834_ = new_G1187_;
  assign new_E5835_ = new_G1254_;
  assign new_E5836_ = new_G1321_;
  assign new_E5837_ = new_G1388_;
  assign new_E5838_ = new_G1455_;
  assign new_E5839_ = new_E5846_ & new_E5845_;
  assign new_E5840_ = new_E5848_ | new_E5847_;
  assign new_E5841_ = new_E5850_ | new_E5849_;
  assign new_E5842_ = new_E5852_ & new_E5851_;
  assign new_E5843_ = new_E5852_ & new_E5853_;
  assign new_E5844_ = new_E5845_ | new_E5854_;
  assign new_E5845_ = new_E5834_ | new_E5857_;
  assign new_E5846_ = new_E5856_ | new_E5855_;
  assign new_E5847_ = new_E5861_ & new_E5860_;
  assign new_E5848_ = new_E5859_ & new_E5858_;
  assign new_E5849_ = new_E5864_ | new_E5863_;
  assign new_E5850_ = new_E5859_ & new_E5862_;
  assign new_E5851_ = new_E5834_ | new_E5867_;
  assign new_E5852_ = new_E5866_ | new_E5865_;
  assign new_E5853_ = new_E5869_ | new_E5868_;
  assign new_E5854_ = ~new_E5845_ & new_E5871_;
  assign new_E5855_ = ~new_E5847_ & new_E5859_;
  assign new_E5856_ = new_E5847_ & ~new_E5859_;
  assign new_E5857_ = new_E5833_ & ~new_E5834_;
  assign new_E5858_ = ~new_E5880_ | ~new_E5881_;
  assign new_E5859_ = new_E5873_ | new_E5875_;
  assign new_E5860_ = new_E5883_ | new_E5882_;
  assign new_E5861_ = new_E5877_ | new_E5876_;
  assign new_E5862_ = ~new_E5885_ | ~new_E5884_;
  assign new_E5863_ = ~new_E5886_ & new_E5887_;
  assign new_E5864_ = new_E5886_ & ~new_E5887_;
  assign new_E5865_ = ~new_E5833_ & new_E5834_;
  assign new_E5866_ = new_E5833_ & ~new_E5834_;
  assign new_E5867_ = ~new_E5849_ | new_E5859_;
  assign new_E5868_ = new_E5849_ & new_E5859_;
  assign new_E5869_ = ~new_E5849_ & ~new_E5859_;
  assign new_E5870_ = new_E5891_ | new_E5890_;
  assign new_E5871_ = new_E5837_ | new_E5870_;
  assign new_E5872_ = new_E5895_ | new_E5894_;
  assign new_E5873_ = ~new_E5837_ & new_E5872_;
  assign new_E5874_ = new_E5893_ | new_E5892_;
  assign new_E5875_ = new_E5837_ & new_E5874_;
  assign new_E5876_ = new_E5835_ & ~new_E5845_;
  assign new_E5877_ = ~new_E5835_ & new_E5845_;
  assign new_E5878_ = ~new_E5834_ | ~new_E5859_;
  assign new_E5879_ = new_E5845_ & new_E5878_;
  assign new_E5880_ = ~new_E5845_ & ~new_E5879_;
  assign new_E5881_ = new_E5845_ | new_E5878_;
  assign new_E5882_ = ~new_E5835_ & new_E5836_;
  assign new_E5883_ = new_E5835_ & ~new_E5836_;
  assign new_E5884_ = new_E5852_ | new_E5889_;
  assign new_E5885_ = ~new_E5852_ & ~new_E5888_;
  assign new_E5886_ = new_E5835_ | new_E5852_;
  assign new_E5887_ = new_E5835_ | new_E5836_;
  assign new_E5888_ = new_E5852_ & new_E5889_;
  assign new_E5889_ = ~new_E5834_ | ~new_E5859_;
  assign new_E5890_ = new_E5867_ & new_E5887_;
  assign new_E5891_ = ~new_E5867_ & ~new_E5887_;
  assign new_E5892_ = new_E5896_ | new_E5897_;
  assign new_E5893_ = ~new_E5838_ & new_E5852_;
  assign new_E5894_ = new_E5898_ | new_E5899_;
  assign new_E5895_ = new_E5838_ & new_E5852_;
  assign new_E5896_ = ~new_E5838_ & ~new_E5852_;
  assign new_E5897_ = new_E5838_ & ~new_E5852_;
  assign new_E5898_ = new_E5838_ & ~new_E5852_;
  assign new_E5899_ = ~new_E5838_ & new_E5852_;
  assign new_E5900_ = new_G1522_;
  assign new_E5901_ = new_G1589_;
  assign new_E5902_ = new_G1656_;
  assign new_E5903_ = new_G1723_;
  assign new_E5904_ = new_G1790_;
  assign new_E5905_ = new_G1857_;
  assign new_E5906_ = new_E5913_ & new_E5912_;
  assign new_E5907_ = new_E5915_ | new_E5914_;
  assign new_E5908_ = new_E5917_ | new_E5916_;
  assign new_E5909_ = new_E5919_ & new_E5918_;
  assign new_E5910_ = new_E5919_ & new_E5920_;
  assign new_E5911_ = new_E5912_ | new_E5921_;
  assign new_E5912_ = new_E5901_ | new_E5924_;
  assign new_E5913_ = new_E5923_ | new_E5922_;
  assign new_E5914_ = new_E5928_ & new_E5927_;
  assign new_E5915_ = new_E5926_ & new_E5925_;
  assign new_E5916_ = new_E5931_ | new_E5930_;
  assign new_E5917_ = new_E5926_ & new_E5929_;
  assign new_E5918_ = new_E5901_ | new_E5934_;
  assign new_E5919_ = new_E5933_ | new_E5932_;
  assign new_E5920_ = new_E5936_ | new_E5935_;
  assign new_E5921_ = ~new_E5912_ & new_E5938_;
  assign new_E5922_ = ~new_E5914_ & new_E5926_;
  assign new_E5923_ = new_E5914_ & ~new_E5926_;
  assign new_E5924_ = new_E5900_ & ~new_E5901_;
  assign new_E5925_ = ~new_E5947_ | ~new_E5948_;
  assign new_E5926_ = new_E5940_ | new_E5942_;
  assign new_E5927_ = new_E5950_ | new_E5949_;
  assign new_E5928_ = new_E5944_ | new_E5943_;
  assign new_E5929_ = ~new_E5952_ | ~new_E5951_;
  assign new_E5930_ = ~new_E5953_ & new_E5954_;
  assign new_E5931_ = new_E5953_ & ~new_E5954_;
  assign new_E5932_ = ~new_E5900_ & new_E5901_;
  assign new_E5933_ = new_E5900_ & ~new_E5901_;
  assign new_E5934_ = ~new_E5916_ | new_E5926_;
  assign new_E5935_ = new_E5916_ & new_E5926_;
  assign new_E5936_ = ~new_E5916_ & ~new_E5926_;
  assign new_E5937_ = new_E5958_ | new_E5957_;
  assign new_E5938_ = new_E5904_ | new_E5937_;
  assign new_E5939_ = new_E5962_ | new_E5961_;
  assign new_E5940_ = ~new_E5904_ & new_E5939_;
  assign new_E5941_ = new_E5960_ | new_E5959_;
  assign new_E5942_ = new_E5904_ & new_E5941_;
  assign new_E5943_ = new_E5902_ & ~new_E5912_;
  assign new_E5944_ = ~new_E5902_ & new_E5912_;
  assign new_E5945_ = ~new_E5901_ | ~new_E5926_;
  assign new_E5946_ = new_E5912_ & new_E5945_;
  assign new_E5947_ = ~new_E5912_ & ~new_E5946_;
  assign new_E5948_ = new_E5912_ | new_E5945_;
  assign new_E5949_ = ~new_E5902_ & new_E5903_;
  assign new_E5950_ = new_E5902_ & ~new_E5903_;
  assign new_E5951_ = new_E5919_ | new_E5956_;
  assign new_E5952_ = ~new_E5919_ & ~new_E5955_;
  assign new_E5953_ = new_E5902_ | new_E5919_;
  assign new_E5954_ = new_E5902_ | new_E5903_;
  assign new_E5955_ = new_E5919_ & new_E5956_;
  assign new_E5956_ = ~new_E5901_ | ~new_E5926_;
  assign new_E5957_ = new_E5934_ & new_E5954_;
  assign new_E5958_ = ~new_E5934_ & ~new_E5954_;
  assign new_E5959_ = new_E5963_ | new_E5964_;
  assign new_E5960_ = ~new_E5905_ & new_E5919_;
  assign new_E5961_ = new_E5965_ | new_E5966_;
  assign new_E5962_ = new_E5905_ & new_E5919_;
  assign new_E5963_ = ~new_E5905_ & ~new_E5919_;
  assign new_E5964_ = new_E5905_ & ~new_E5919_;
  assign new_E5965_ = new_E5905_ & ~new_E5919_;
  assign new_E5966_ = ~new_E5905_ & new_E5919_;
  assign new_E5967_ = new_G1924_;
  assign new_E5968_ = new_G1991_;
  assign new_E5969_ = new_G2058_;
  assign new_E5970_ = new_G2125_;
  assign new_E5971_ = new_G2192_;
  assign new_E5972_ = new_G2259_;
  assign new_E5973_ = new_E5980_ & new_E5979_;
  assign new_E5974_ = new_E5982_ | new_E5981_;
  assign new_E5975_ = new_E5984_ | new_E5983_;
  assign new_E5976_ = new_E5986_ & new_E5985_;
  assign new_E5977_ = new_E5986_ & new_E5987_;
  assign new_E5978_ = new_E5979_ | new_E5988_;
  assign new_E5979_ = new_E5968_ | new_E5991_;
  assign new_E5980_ = new_E5990_ | new_E5989_;
  assign new_E5981_ = new_E5995_ & new_E5994_;
  assign new_E5982_ = new_E5993_ & new_E5992_;
  assign new_E5983_ = new_E5998_ | new_E5997_;
  assign new_E5984_ = new_E5993_ & new_E5996_;
  assign new_E5985_ = new_E5968_ | new_E6001_;
  assign new_E5986_ = new_E6000_ | new_E5999_;
  assign new_E5987_ = new_E6003_ | new_E6002_;
  assign new_E5988_ = ~new_E5979_ & new_E6005_;
  assign new_E5989_ = ~new_E5981_ & new_E5993_;
  assign new_E5990_ = new_E5981_ & ~new_E5993_;
  assign new_E5991_ = new_E5967_ & ~new_E5968_;
  assign new_E5992_ = ~new_E6014_ | ~new_E6015_;
  assign new_E5993_ = new_E6007_ | new_E6009_;
  assign new_E5994_ = new_E6017_ | new_E6016_;
  assign new_E5995_ = new_E6011_ | new_E6010_;
  assign new_E5996_ = ~new_E6019_ | ~new_E6018_;
  assign new_E5997_ = ~new_E6020_ & new_E6021_;
  assign new_E5998_ = new_E6020_ & ~new_E6021_;
  assign new_E5999_ = ~new_E5967_ & new_E5968_;
  assign new_E6000_ = new_E5967_ & ~new_E5968_;
  assign new_E6001_ = ~new_E5983_ | new_E5993_;
  assign new_E6002_ = new_E5983_ & new_E5993_;
  assign new_E6003_ = ~new_E5983_ & ~new_E5993_;
  assign new_E6004_ = new_E6025_ | new_E6024_;
  assign new_E6005_ = new_E5971_ | new_E6004_;
  assign new_E6006_ = new_E6029_ | new_E6028_;
  assign new_E6007_ = ~new_E5971_ & new_E6006_;
  assign new_E6008_ = new_E6027_ | new_E6026_;
  assign new_E6009_ = new_E5971_ & new_E6008_;
  assign new_E6010_ = new_E5969_ & ~new_E5979_;
  assign new_E6011_ = ~new_E5969_ & new_E5979_;
  assign new_E6012_ = ~new_E5968_ | ~new_E5993_;
  assign new_E6013_ = new_E5979_ & new_E6012_;
  assign new_E6014_ = ~new_E5979_ & ~new_E6013_;
  assign new_E6015_ = new_E5979_ | new_E6012_;
  assign new_E6016_ = ~new_E5969_ & new_E5970_;
  assign new_E6017_ = new_E5969_ & ~new_E5970_;
  assign new_E6018_ = new_E5986_ | new_E6023_;
  assign new_E6019_ = ~new_E5986_ & ~new_E6022_;
  assign new_E6020_ = new_E5969_ | new_E5986_;
  assign new_E6021_ = new_E5969_ | new_E5970_;
  assign new_E6022_ = new_E5986_ & new_E6023_;
  assign new_E6023_ = ~new_E5968_ | ~new_E5993_;
  assign new_E6024_ = new_E6001_ & new_E6021_;
  assign new_E6025_ = ~new_E6001_ & ~new_E6021_;
  assign new_E6026_ = new_E6030_ | new_E6031_;
  assign new_E6027_ = ~new_E5972_ & new_E5986_;
  assign new_E6028_ = new_E6032_ | new_E6033_;
  assign new_E6029_ = new_E5972_ & new_E5986_;
  assign new_E6030_ = ~new_E5972_ & ~new_E5986_;
  assign new_E6031_ = new_E5972_ & ~new_E5986_;
  assign new_E6032_ = new_E5972_ & ~new_E5986_;
  assign new_E6033_ = ~new_E5972_ & new_E5986_;
  assign new_E6034_ = new_G2326_;
  assign new_E6035_ = new_G2393_;
  assign new_E6036_ = new_G2460_;
  assign new_E6037_ = new_G2527_;
  assign new_E6038_ = new_G2594_;
  assign new_E6039_ = new_G2661_;
  assign new_E6040_ = new_E6047_ & new_E6046_;
  assign new_E6041_ = new_E6049_ | new_E6048_;
  assign new_E6042_ = new_E6051_ | new_E6050_;
  assign new_E6043_ = new_E6053_ & new_E6052_;
  assign new_E6044_ = new_E6053_ & new_E6054_;
  assign new_E6045_ = new_E6046_ | new_E6055_;
  assign new_E6046_ = new_E6035_ | new_E6058_;
  assign new_E6047_ = new_E6057_ | new_E6056_;
  assign new_E6048_ = new_E6062_ & new_E6061_;
  assign new_E6049_ = new_E6060_ & new_E6059_;
  assign new_E6050_ = new_E6065_ | new_E6064_;
  assign new_E6051_ = new_E6060_ & new_E6063_;
  assign new_E6052_ = new_E6035_ | new_E6068_;
  assign new_E6053_ = new_E6067_ | new_E6066_;
  assign new_E6054_ = new_E6070_ | new_E6069_;
  assign new_E6055_ = ~new_E6046_ & new_E6072_;
  assign new_E6056_ = ~new_E6048_ & new_E6060_;
  assign new_E6057_ = new_E6048_ & ~new_E6060_;
  assign new_E6058_ = new_E6034_ & ~new_E6035_;
  assign new_E6059_ = ~new_E6081_ | ~new_E6082_;
  assign new_E6060_ = new_E6074_ | new_E6076_;
  assign new_E6061_ = new_E6084_ | new_E6083_;
  assign new_E6062_ = new_E6078_ | new_E6077_;
  assign new_E6063_ = ~new_E6086_ | ~new_E6085_;
  assign new_E6064_ = ~new_E6087_ & new_E6088_;
  assign new_E6065_ = new_E6087_ & ~new_E6088_;
  assign new_E6066_ = ~new_E6034_ & new_E6035_;
  assign new_E6067_ = new_E6034_ & ~new_E6035_;
  assign new_E6068_ = ~new_E6050_ | new_E6060_;
  assign new_E6069_ = new_E6050_ & new_E6060_;
  assign new_E6070_ = ~new_E6050_ & ~new_E6060_;
  assign new_E6071_ = new_E6092_ | new_E6091_;
  assign new_E6072_ = new_E6038_ | new_E6071_;
  assign new_E6073_ = new_E6096_ | new_E6095_;
  assign new_E6074_ = ~new_E6038_ & new_E6073_;
  assign new_E6075_ = new_E6094_ | new_E6093_;
  assign new_E6076_ = new_E6038_ & new_E6075_;
  assign new_E6077_ = new_E6036_ & ~new_E6046_;
  assign new_E6078_ = ~new_E6036_ & new_E6046_;
  assign new_E6079_ = ~new_E6035_ | ~new_E6060_;
  assign new_E6080_ = new_E6046_ & new_E6079_;
  assign new_E6081_ = ~new_E6046_ & ~new_E6080_;
  assign new_E6082_ = new_E6046_ | new_E6079_;
  assign new_E6083_ = ~new_E6036_ & new_E6037_;
  assign new_E6084_ = new_E6036_ & ~new_E6037_;
  assign new_E6085_ = new_E6053_ | new_E6090_;
  assign new_E6086_ = ~new_E6053_ & ~new_E6089_;
  assign new_E6087_ = new_E6036_ | new_E6053_;
  assign new_E6088_ = new_E6036_ | new_E6037_;
  assign new_E6089_ = new_E6053_ & new_E6090_;
  assign new_E6090_ = ~new_E6035_ | ~new_E6060_;
  assign new_E6091_ = new_E6068_ & new_E6088_;
  assign new_E6092_ = ~new_E6068_ & ~new_E6088_;
  assign new_E6093_ = new_E6097_ | new_E6098_;
  assign new_E6094_ = ~new_E6039_ & new_E6053_;
  assign new_E6095_ = new_E6099_ | new_E6100_;
  assign new_E6096_ = new_E6039_ & new_E6053_;
  assign new_E6097_ = ~new_E6039_ & ~new_E6053_;
  assign new_E6098_ = new_E6039_ & ~new_E6053_;
  assign new_E6099_ = new_E6039_ & ~new_E6053_;
  assign new_E6100_ = ~new_E6039_ & new_E6053_;
  assign new_E6101_ = new_G2728_;
  assign new_E6102_ = new_G2795_;
  assign new_E6103_ = new_G2862_;
  assign new_E6104_ = new_G2929_;
  assign new_E6105_ = new_G2996_;
  assign new_E6106_ = new_G3063_;
  assign new_E6107_ = new_E6114_ & new_E6113_;
  assign new_E6108_ = new_E6116_ | new_E6115_;
  assign new_E6109_ = new_E6118_ | new_E6117_;
  assign new_E6110_ = new_E6120_ & new_E6119_;
  assign new_E6111_ = new_E6120_ & new_E6121_;
  assign new_E6112_ = new_E6113_ | new_E6122_;
  assign new_E6113_ = new_E6102_ | new_E6125_;
  assign new_E6114_ = new_E6124_ | new_E6123_;
  assign new_E6115_ = new_E6129_ & new_E6128_;
  assign new_E6116_ = new_E6127_ & new_E6126_;
  assign new_E6117_ = new_E6132_ | new_E6131_;
  assign new_E6118_ = new_E6127_ & new_E6130_;
  assign new_E6119_ = new_E6102_ | new_E6135_;
  assign new_E6120_ = new_E6134_ | new_E6133_;
  assign new_E6121_ = new_E6137_ | new_E6136_;
  assign new_E6122_ = ~new_E6113_ & new_E6139_;
  assign new_E6123_ = ~new_E6115_ & new_E6127_;
  assign new_E6124_ = new_E6115_ & ~new_E6127_;
  assign new_E6125_ = new_E6101_ & ~new_E6102_;
  assign new_E6126_ = ~new_E6148_ | ~new_E6149_;
  assign new_E6127_ = new_E6141_ | new_E6143_;
  assign new_E6128_ = new_E6151_ | new_E6150_;
  assign new_E6129_ = new_E6145_ | new_E6144_;
  assign new_E6130_ = ~new_E6153_ | ~new_E6152_;
  assign new_E6131_ = ~new_E6154_ & new_E6155_;
  assign new_E6132_ = new_E6154_ & ~new_E6155_;
  assign new_E6133_ = ~new_E6101_ & new_E6102_;
  assign new_E6134_ = new_E6101_ & ~new_E6102_;
  assign new_E6135_ = ~new_E6117_ | new_E6127_;
  assign new_E6136_ = new_E6117_ & new_E6127_;
  assign new_E6137_ = ~new_E6117_ & ~new_E6127_;
  assign new_E6138_ = new_E6159_ | new_E6158_;
  assign new_E6139_ = new_E6105_ | new_E6138_;
  assign new_E6140_ = new_E6163_ | new_E6162_;
  assign new_E6141_ = ~new_E6105_ & new_E6140_;
  assign new_E6142_ = new_E6161_ | new_E6160_;
  assign new_E6143_ = new_E6105_ & new_E6142_;
  assign new_E6144_ = new_E6103_ & ~new_E6113_;
  assign new_E6145_ = ~new_E6103_ & new_E6113_;
  assign new_E6146_ = ~new_E6102_ | ~new_E6127_;
  assign new_E6147_ = new_E6113_ & new_E6146_;
  assign new_E6148_ = ~new_E6113_ & ~new_E6147_;
  assign new_E6149_ = new_E6113_ | new_E6146_;
  assign new_E6150_ = ~new_E6103_ & new_E6104_;
  assign new_E6151_ = new_E6103_ & ~new_E6104_;
  assign new_E6152_ = new_E6120_ | new_E6157_;
  assign new_E6153_ = ~new_E6120_ & ~new_E6156_;
  assign new_E6154_ = new_E6103_ | new_E6120_;
  assign new_E6155_ = new_E6103_ | new_E6104_;
  assign new_E6156_ = new_E6120_ & new_E6157_;
  assign new_E6157_ = ~new_E6102_ | ~new_E6127_;
  assign new_E6158_ = new_E6135_ & new_E6155_;
  assign new_E6159_ = ~new_E6135_ & ~new_E6155_;
  assign new_E6160_ = new_E6164_ | new_E6165_;
  assign new_E6161_ = ~new_E6106_ & new_E6120_;
  assign new_E6162_ = new_E6166_ | new_E6167_;
  assign new_E6163_ = new_E6106_ & new_E6120_;
  assign new_E6164_ = ~new_E6106_ & ~new_E6120_;
  assign new_E6165_ = new_E6106_ & ~new_E6120_;
  assign new_E6166_ = new_E6106_ & ~new_E6120_;
  assign new_E6167_ = ~new_E6106_ & new_E6120_;
  assign new_E6168_ = new_G3130_;
  assign new_E6169_ = new_G3197_;
  assign new_E6170_ = new_G3264_;
  assign new_E6171_ = new_G3331_;
  assign new_E6172_ = new_G3398_;
  assign new_E6173_ = new_G3465_;
  assign new_E6174_ = new_E6181_ & new_E6180_;
  assign new_E6175_ = new_E6183_ | new_E6182_;
  assign new_E6176_ = new_E6185_ | new_E6184_;
  assign new_E6177_ = new_E6187_ & new_E6186_;
  assign new_E6178_ = new_E6187_ & new_E6188_;
  assign new_E6179_ = new_E6180_ | new_E6189_;
  assign new_E6180_ = new_E6169_ | new_E6192_;
  assign new_E6181_ = new_E6191_ | new_E6190_;
  assign new_E6182_ = new_E6196_ & new_E6195_;
  assign new_E6183_ = new_E6194_ & new_E6193_;
  assign new_E6184_ = new_E6199_ | new_E6198_;
  assign new_E6185_ = new_E6194_ & new_E6197_;
  assign new_E6186_ = new_E6169_ | new_E6202_;
  assign new_E6187_ = new_E6201_ | new_E6200_;
  assign new_E6188_ = new_E6204_ | new_E6203_;
  assign new_E6189_ = ~new_E6180_ & new_E6206_;
  assign new_E6190_ = ~new_E6182_ & new_E6194_;
  assign new_E6191_ = new_E6182_ & ~new_E6194_;
  assign new_E6192_ = new_E6168_ & ~new_E6169_;
  assign new_E6193_ = ~new_E6215_ | ~new_E6216_;
  assign new_E6194_ = new_E6208_ | new_E6210_;
  assign new_E6195_ = new_E6218_ | new_E6217_;
  assign new_E6196_ = new_E6212_ | new_E6211_;
  assign new_E6197_ = ~new_E6220_ | ~new_E6219_;
  assign new_E6198_ = ~new_E6221_ & new_E6222_;
  assign new_E6199_ = new_E6221_ & ~new_E6222_;
  assign new_E6200_ = ~new_E6168_ & new_E6169_;
  assign new_E6201_ = new_E6168_ & ~new_E6169_;
  assign new_E6202_ = ~new_E6184_ | new_E6194_;
  assign new_E6203_ = new_E6184_ & new_E6194_;
  assign new_E6204_ = ~new_E6184_ & ~new_E6194_;
  assign new_E6205_ = new_E6226_ | new_E6225_;
  assign new_E6206_ = new_E6172_ | new_E6205_;
  assign new_E6207_ = new_E6230_ | new_E6229_;
  assign new_E6208_ = ~new_E6172_ & new_E6207_;
  assign new_E6209_ = new_E6228_ | new_E6227_;
  assign new_E6210_ = new_E6172_ & new_E6209_;
  assign new_E6211_ = new_E6170_ & ~new_E6180_;
  assign new_E6212_ = ~new_E6170_ & new_E6180_;
  assign new_E6213_ = ~new_E6169_ | ~new_E6194_;
  assign new_E6214_ = new_E6180_ & new_E6213_;
  assign new_E6215_ = ~new_E6180_ & ~new_E6214_;
  assign new_E6216_ = new_E6180_ | new_E6213_;
  assign new_E6217_ = ~new_E6170_ & new_E6171_;
  assign new_E6218_ = new_E6170_ & ~new_E6171_;
  assign new_E6219_ = new_E6187_ | new_E6224_;
  assign new_E6220_ = ~new_E6187_ & ~new_E6223_;
  assign new_E6221_ = new_E6170_ | new_E6187_;
  assign new_E6222_ = new_E6170_ | new_E6171_;
  assign new_E6223_ = new_E6187_ & new_E6224_;
  assign new_E6224_ = ~new_E6169_ | ~new_E6194_;
  assign new_E6225_ = new_E6202_ & new_E6222_;
  assign new_E6226_ = ~new_E6202_ & ~new_E6222_;
  assign new_E6227_ = new_E6231_ | new_E6232_;
  assign new_E6228_ = ~new_E6173_ & new_E6187_;
  assign new_E6229_ = new_E6233_ | new_E6234_;
  assign new_E6230_ = new_E6173_ & new_E6187_;
  assign new_E6231_ = ~new_E6173_ & ~new_E6187_;
  assign new_E6232_ = new_E6173_ & ~new_E6187_;
  assign new_E6233_ = new_E6173_ & ~new_E6187_;
  assign new_E6234_ = ~new_E6173_ & new_E6187_;
  assign new_E6235_ = new_G3532_;
  assign new_E6236_ = new_G3599_;
  assign new_E6237_ = new_G3666_;
  assign new_E6238_ = new_G3733_;
  assign new_E6239_ = new_G3800_;
  assign new_E6240_ = new_G3867_;
  assign new_E6241_ = new_E6248_ & new_E6247_;
  assign new_E6242_ = new_E6250_ | new_E6249_;
  assign new_E6243_ = new_E6252_ | new_E6251_;
  assign new_E6244_ = new_E6254_ & new_E6253_;
  assign new_E6245_ = new_E6254_ & new_E6255_;
  assign new_E6246_ = new_E6247_ | new_E6256_;
  assign new_E6247_ = new_E6236_ | new_E6259_;
  assign new_E6248_ = new_E6258_ | new_E6257_;
  assign new_E6249_ = new_E6263_ & new_E6262_;
  assign new_E6250_ = new_E6261_ & new_E6260_;
  assign new_E6251_ = new_E6266_ | new_E6265_;
  assign new_E6252_ = new_E6261_ & new_E6264_;
  assign new_E6253_ = new_E6236_ | new_E6269_;
  assign new_E6254_ = new_E6268_ | new_E6267_;
  assign new_E6255_ = new_E6271_ | new_E6270_;
  assign new_E6256_ = ~new_E6247_ & new_E6273_;
  assign new_E6257_ = ~new_E6249_ & new_E6261_;
  assign new_E6258_ = new_E6249_ & ~new_E6261_;
  assign new_E6259_ = new_E6235_ & ~new_E6236_;
  assign new_E6260_ = ~new_E6282_ | ~new_E6283_;
  assign new_E6261_ = new_E6275_ | new_E6277_;
  assign new_E6262_ = new_E6285_ | new_E6284_;
  assign new_E6263_ = new_E6279_ | new_E6278_;
  assign new_E6264_ = ~new_E6287_ | ~new_E6286_;
  assign new_E6265_ = ~new_E6288_ & new_E6289_;
  assign new_E6266_ = new_E6288_ & ~new_E6289_;
  assign new_E6267_ = ~new_E6235_ & new_E6236_;
  assign new_E6268_ = new_E6235_ & ~new_E6236_;
  assign new_E6269_ = ~new_E6251_ | new_E6261_;
  assign new_E6270_ = new_E6251_ & new_E6261_;
  assign new_E6271_ = ~new_E6251_ & ~new_E6261_;
  assign new_E6272_ = new_E6293_ | new_E6292_;
  assign new_E6273_ = new_E6239_ | new_E6272_;
  assign new_E6274_ = new_E6297_ | new_E6296_;
  assign new_E6275_ = ~new_E6239_ & new_E6274_;
  assign new_E6276_ = new_E6295_ | new_E6294_;
  assign new_E6277_ = new_E6239_ & new_E6276_;
  assign new_E6278_ = new_E6237_ & ~new_E6247_;
  assign new_E6279_ = ~new_E6237_ & new_E6247_;
  assign new_E6280_ = ~new_E6236_ | ~new_E6261_;
  assign new_E6281_ = new_E6247_ & new_E6280_;
  assign new_E6282_ = ~new_E6247_ & ~new_E6281_;
  assign new_E6283_ = new_E6247_ | new_E6280_;
  assign new_E6284_ = ~new_E6237_ & new_E6238_;
  assign new_E6285_ = new_E6237_ & ~new_E6238_;
  assign new_E6286_ = new_E6254_ | new_E6291_;
  assign new_E6287_ = ~new_E6254_ & ~new_E6290_;
  assign new_E6288_ = new_E6237_ | new_E6254_;
  assign new_E6289_ = new_E6237_ | new_E6238_;
  assign new_E6290_ = new_E6254_ & new_E6291_;
  assign new_E6291_ = ~new_E6236_ | ~new_E6261_;
  assign new_E6292_ = new_E6269_ & new_E6289_;
  assign new_E6293_ = ~new_E6269_ & ~new_E6289_;
  assign new_E6294_ = new_E6298_ | new_E6299_;
  assign new_E6295_ = ~new_E6240_ & new_E6254_;
  assign new_E6296_ = new_E6300_ | new_E6301_;
  assign new_E6297_ = new_E6240_ & new_E6254_;
  assign new_E6298_ = ~new_E6240_ & ~new_E6254_;
  assign new_E6299_ = new_E6240_ & ~new_E6254_;
  assign new_E6300_ = new_E6240_ & ~new_E6254_;
  assign new_E6301_ = ~new_E6240_ & new_E6254_;
  assign new_E6302_ = new_G3934_;
  assign new_E6303_ = new_G4001_;
  assign new_E6304_ = new_G4068_;
  assign new_E6305_ = new_G4135_;
  assign new_E6306_ = new_G4202_;
  assign new_E6307_ = new_G4269_;
  assign new_E6308_ = new_E6315_ & new_E6314_;
  assign new_E6309_ = new_E6317_ | new_E6316_;
  assign new_E6310_ = new_E6319_ | new_E6318_;
  assign new_E6311_ = new_E6321_ & new_E6320_;
  assign new_E6312_ = new_E6321_ & new_E6322_;
  assign new_E6313_ = new_E6314_ | new_E6323_;
  assign new_E6314_ = new_E6303_ | new_E6326_;
  assign new_E6315_ = new_E6325_ | new_E6324_;
  assign new_E6316_ = new_E6330_ & new_E6329_;
  assign new_E6317_ = new_E6328_ & new_E6327_;
  assign new_E6318_ = new_E6333_ | new_E6332_;
  assign new_E6319_ = new_E6328_ & new_E6331_;
  assign new_E6320_ = new_E6303_ | new_E6336_;
  assign new_E6321_ = new_E6335_ | new_E6334_;
  assign new_E6322_ = new_E6338_ | new_E6337_;
  assign new_E6323_ = ~new_E6314_ & new_E6340_;
  assign new_E6324_ = ~new_E6316_ & new_E6328_;
  assign new_E6325_ = new_E6316_ & ~new_E6328_;
  assign new_E6326_ = new_E6302_ & ~new_E6303_;
  assign new_E6327_ = ~new_E6349_ | ~new_E6350_;
  assign new_E6328_ = new_E6342_ | new_E6344_;
  assign new_E6329_ = new_E6352_ | new_E6351_;
  assign new_E6330_ = new_E6346_ | new_E6345_;
  assign new_E6331_ = ~new_E6354_ | ~new_E6353_;
  assign new_E6332_ = ~new_E6355_ & new_E6356_;
  assign new_E6333_ = new_E6355_ & ~new_E6356_;
  assign new_E6334_ = ~new_E6302_ & new_E6303_;
  assign new_E6335_ = new_E6302_ & ~new_E6303_;
  assign new_E6336_ = ~new_E6318_ | new_E6328_;
  assign new_E6337_ = new_E6318_ & new_E6328_;
  assign new_E6338_ = ~new_E6318_ & ~new_E6328_;
  assign new_E6339_ = new_E6360_ | new_E6359_;
  assign new_E6340_ = new_E6306_ | new_E6339_;
  assign new_E6341_ = new_E6364_ | new_E6363_;
  assign new_E6342_ = ~new_E6306_ & new_E6341_;
  assign new_E6343_ = new_E6362_ | new_E6361_;
  assign new_E6344_ = new_E6306_ & new_E6343_;
  assign new_E6345_ = new_E6304_ & ~new_E6314_;
  assign new_E6346_ = ~new_E6304_ & new_E6314_;
  assign new_E6347_ = ~new_E6303_ | ~new_E6328_;
  assign new_E6348_ = new_E6314_ & new_E6347_;
  assign new_E6349_ = ~new_E6314_ & ~new_E6348_;
  assign new_E6350_ = new_E6314_ | new_E6347_;
  assign new_E6351_ = ~new_E6304_ & new_E6305_;
  assign new_E6352_ = new_E6304_ & ~new_E6305_;
  assign new_E6353_ = new_E6321_ | new_E6358_;
  assign new_E6354_ = ~new_E6321_ & ~new_E6357_;
  assign new_E6355_ = new_E6304_ | new_E6321_;
  assign new_E6356_ = new_E6304_ | new_E6305_;
  assign new_E6357_ = new_E6321_ & new_E6358_;
  assign new_E6358_ = ~new_E6303_ | ~new_E6328_;
  assign new_E6359_ = new_E6336_ & new_E6356_;
  assign new_E6360_ = ~new_E6336_ & ~new_E6356_;
  assign new_E6361_ = new_E6365_ | new_E6366_;
  assign new_E6362_ = ~new_E6307_ & new_E6321_;
  assign new_E6363_ = new_E6367_ | new_E6368_;
  assign new_E6364_ = new_E6307_ & new_E6321_;
  assign new_E6365_ = ~new_E6307_ & ~new_E6321_;
  assign new_E6366_ = new_E6307_ & ~new_E6321_;
  assign new_E6367_ = new_E6307_ & ~new_E6321_;
  assign new_E6368_ = ~new_E6307_ & new_E6321_;
  assign new_E6369_ = new_G4336_;
  assign new_E6370_ = new_G4403_;
  assign new_E6371_ = new_G4470_;
  assign new_E6372_ = new_G4537_;
  assign new_E6373_ = new_G4604_;
  assign new_E6374_ = new_G4671_;
  assign new_E6375_ = new_E6382_ & new_E6381_;
  assign new_E6376_ = new_E6384_ | new_E6383_;
  assign new_E6377_ = new_E6386_ | new_E6385_;
  assign new_E6378_ = new_E6388_ & new_E6387_;
  assign new_E6379_ = new_E6388_ & new_E6389_;
  assign new_E6380_ = new_E6381_ | new_E6390_;
  assign new_E6381_ = new_E6370_ | new_E6393_;
  assign new_E6382_ = new_E6392_ | new_E6391_;
  assign new_E6383_ = new_E6397_ & new_E6396_;
  assign new_E6384_ = new_E6395_ & new_E6394_;
  assign new_E6385_ = new_E6400_ | new_E6399_;
  assign new_E6386_ = new_E6395_ & new_E6398_;
  assign new_E6387_ = new_E6370_ | new_E6403_;
  assign new_E6388_ = new_E6402_ | new_E6401_;
  assign new_E6389_ = new_E6405_ | new_E6404_;
  assign new_E6390_ = ~new_E6381_ & new_E6407_;
  assign new_E6391_ = ~new_E6383_ & new_E6395_;
  assign new_E6392_ = new_E6383_ & ~new_E6395_;
  assign new_E6393_ = new_E6369_ & ~new_E6370_;
  assign new_E6394_ = ~new_E6416_ | ~new_E6417_;
  assign new_E6395_ = new_E6409_ | new_E6411_;
  assign new_E6396_ = new_E6419_ | new_E6418_;
  assign new_E6397_ = new_E6413_ | new_E6412_;
  assign new_E6398_ = ~new_E6421_ | ~new_E6420_;
  assign new_E6399_ = ~new_E6422_ & new_E6423_;
  assign new_E6400_ = new_E6422_ & ~new_E6423_;
  assign new_E6401_ = ~new_E6369_ & new_E6370_;
  assign new_E6402_ = new_E6369_ & ~new_E6370_;
  assign new_E6403_ = ~new_E6385_ | new_E6395_;
  assign new_E6404_ = new_E6385_ & new_E6395_;
  assign new_E6405_ = ~new_E6385_ & ~new_E6395_;
  assign new_E6406_ = new_E6427_ | new_E6426_;
  assign new_E6407_ = new_E6373_ | new_E6406_;
  assign new_E6408_ = new_E6431_ | new_E6430_;
  assign new_E6409_ = ~new_E6373_ & new_E6408_;
  assign new_E6410_ = new_E6429_ | new_E6428_;
  assign new_E6411_ = new_E6373_ & new_E6410_;
  assign new_E6412_ = new_E6371_ & ~new_E6381_;
  assign new_E6413_ = ~new_E6371_ & new_E6381_;
  assign new_E6414_ = ~new_E6370_ | ~new_E6395_;
  assign new_E6415_ = new_E6381_ & new_E6414_;
  assign new_E6416_ = ~new_E6381_ & ~new_E6415_;
  assign new_E6417_ = new_E6381_ | new_E6414_;
  assign new_E6418_ = ~new_E6371_ & new_E6372_;
  assign new_E6419_ = new_E6371_ & ~new_E6372_;
  assign new_E6420_ = new_E6388_ | new_E6425_;
  assign new_E6421_ = ~new_E6388_ & ~new_E6424_;
  assign new_E6422_ = new_E6371_ | new_E6388_;
  assign new_E6423_ = new_E6371_ | new_E6372_;
  assign new_E6424_ = new_E6388_ & new_E6425_;
  assign new_E6425_ = ~new_E6370_ | ~new_E6395_;
  assign new_E6426_ = new_E6403_ & new_E6423_;
  assign new_E6427_ = ~new_E6403_ & ~new_E6423_;
  assign new_E6428_ = new_E6432_ | new_E6433_;
  assign new_E6429_ = ~new_E6374_ & new_E6388_;
  assign new_E6430_ = new_E6434_ | new_E6435_;
  assign new_E6431_ = new_E6374_ & new_E6388_;
  assign new_E6432_ = ~new_E6374_ & ~new_E6388_;
  assign new_E6433_ = new_E6374_ & ~new_E6388_;
  assign new_E6434_ = new_E6374_ & ~new_E6388_;
  assign new_E6435_ = ~new_E6374_ & new_E6388_;
  assign new_E6436_ = new_G4738_;
  assign new_E6437_ = new_G4805_;
  assign new_E6438_ = new_G4872_;
  assign new_E6439_ = new_G4939_;
  assign new_E6440_ = new_G5006_;
  assign new_E6441_ = new_G5073_;
  assign new_E6442_ = new_E6449_ & new_E6448_;
  assign new_E6443_ = new_E6451_ | new_E6450_;
  assign new_E6444_ = new_E6453_ | new_E6452_;
  assign new_E6445_ = new_E6455_ & new_E6454_;
  assign new_E6446_ = new_E6455_ & new_E6456_;
  assign new_E6447_ = new_E6448_ | new_E6457_;
  assign new_E6448_ = new_E6437_ | new_E6460_;
  assign new_E6449_ = new_E6459_ | new_E6458_;
  assign new_E6450_ = new_E6464_ & new_E6463_;
  assign new_E6451_ = new_E6462_ & new_E6461_;
  assign new_E6452_ = new_E6467_ | new_E6466_;
  assign new_E6453_ = new_E6462_ & new_E6465_;
  assign new_E6454_ = new_E6437_ | new_E6470_;
  assign new_E6455_ = new_E6469_ | new_E6468_;
  assign new_E6456_ = new_E6472_ | new_E6471_;
  assign new_E6457_ = ~new_E6448_ & new_E6474_;
  assign new_E6458_ = ~new_E6450_ & new_E6462_;
  assign new_E6459_ = new_E6450_ & ~new_E6462_;
  assign new_E6460_ = new_E6436_ & ~new_E6437_;
  assign new_E6461_ = ~new_E6483_ | ~new_E6484_;
  assign new_E6462_ = new_E6476_ | new_E6478_;
  assign new_E6463_ = new_E6486_ | new_E6485_;
  assign new_E6464_ = new_E6480_ | new_E6479_;
  assign new_E6465_ = ~new_E6488_ | ~new_E6487_;
  assign new_E6466_ = ~new_E6489_ & new_E6490_;
  assign new_E6467_ = new_E6489_ & ~new_E6490_;
  assign new_E6468_ = ~new_E6436_ & new_E6437_;
  assign new_E6469_ = new_E6436_ & ~new_E6437_;
  assign new_E6470_ = ~new_E6452_ | new_E6462_;
  assign new_E6471_ = new_E6452_ & new_E6462_;
  assign new_E6472_ = ~new_E6452_ & ~new_E6462_;
  assign new_E6473_ = new_E6494_ | new_E6493_;
  assign new_E6474_ = new_E6440_ | new_E6473_;
  assign new_E6475_ = new_E6498_ | new_E6497_;
  assign new_E6476_ = ~new_E6440_ & new_E6475_;
  assign new_E6477_ = new_E6496_ | new_E6495_;
  assign new_E6478_ = new_E6440_ & new_E6477_;
  assign new_E6479_ = new_E6438_ & ~new_E6448_;
  assign new_E6480_ = ~new_E6438_ & new_E6448_;
  assign new_E6481_ = ~new_E6437_ | ~new_E6462_;
  assign new_E6482_ = new_E6448_ & new_E6481_;
  assign new_E6483_ = ~new_E6448_ & ~new_E6482_;
  assign new_E6484_ = new_E6448_ | new_E6481_;
  assign new_E6485_ = ~new_E6438_ & new_E6439_;
  assign new_E6486_ = new_E6438_ & ~new_E6439_;
  assign new_E6487_ = new_E6455_ | new_E6492_;
  assign new_E6488_ = ~new_E6455_ & ~new_E6491_;
  assign new_E6489_ = new_E6438_ | new_E6455_;
  assign new_E6490_ = new_E6438_ | new_E6439_;
  assign new_E6491_ = new_E6455_ & new_E6492_;
  assign new_E6492_ = ~new_E6437_ | ~new_E6462_;
  assign new_E6493_ = new_E6470_ & new_E6490_;
  assign new_E6494_ = ~new_E6470_ & ~new_E6490_;
  assign new_E6495_ = new_E6499_ | new_E6500_;
  assign new_E6496_ = ~new_E6441_ & new_E6455_;
  assign new_E6497_ = new_E6501_ | new_E6502_;
  assign new_E6498_ = new_E6441_ & new_E6455_;
  assign new_E6499_ = ~new_E6441_ & ~new_E6455_;
  assign new_E6500_ = new_E6441_ & ~new_E6455_;
  assign new_E6501_ = new_E6441_ & ~new_E6455_;
  assign new_E6502_ = ~new_E6441_ & new_E6455_;
  assign new_E6503_ = new_G5140_;
  assign new_E6504_ = new_G5207_;
  assign new_E6505_ = new_G5274_;
  assign new_E6506_ = new_G5341_;
  assign new_E6507_ = new_G5408_;
  assign new_E6508_ = new_G5475_;
  assign new_E6509_ = new_E6516_ & new_E6515_;
  assign new_E6510_ = new_E6518_ | new_E6517_;
  assign new_E6511_ = new_E6520_ | new_E6519_;
  assign new_E6512_ = new_E6522_ & new_E6521_;
  assign new_E6513_ = new_E6522_ & new_E6523_;
  assign new_E6514_ = new_E6515_ | new_E6524_;
  assign new_E6515_ = new_E6504_ | new_E6527_;
  assign new_E6516_ = new_E6526_ | new_E6525_;
  assign new_E6517_ = new_E6531_ & new_E6530_;
  assign new_E6518_ = new_E6529_ & new_E6528_;
  assign new_E6519_ = new_E6534_ | new_E6533_;
  assign new_E6520_ = new_E6529_ & new_E6532_;
  assign new_E6521_ = new_E6504_ | new_E6537_;
  assign new_E6522_ = new_E6536_ | new_E6535_;
  assign new_E6523_ = new_E6539_ | new_E6538_;
  assign new_E6524_ = ~new_E6515_ & new_E6541_;
  assign new_E6525_ = ~new_E6517_ & new_E6529_;
  assign new_E6526_ = new_E6517_ & ~new_E6529_;
  assign new_E6527_ = new_E6503_ & ~new_E6504_;
  assign new_E6528_ = ~new_E6550_ | ~new_E6551_;
  assign new_E6529_ = new_E6543_ | new_E6545_;
  assign new_E6530_ = new_E6553_ | new_E6552_;
  assign new_E6531_ = new_E6547_ | new_E6546_;
  assign new_E6532_ = ~new_E6555_ | ~new_E6554_;
  assign new_E6533_ = ~new_E6556_ & new_E6557_;
  assign new_E6534_ = new_E6556_ & ~new_E6557_;
  assign new_E6535_ = ~new_E6503_ & new_E6504_;
  assign new_E6536_ = new_E6503_ & ~new_E6504_;
  assign new_E6537_ = ~new_E6519_ | new_E6529_;
  assign new_E6538_ = new_E6519_ & new_E6529_;
  assign new_E6539_ = ~new_E6519_ & ~new_E6529_;
  assign new_E6540_ = new_E6561_ | new_E6560_;
  assign new_E6541_ = new_E6507_ | new_E6540_;
  assign new_E6542_ = new_E6565_ | new_E6564_;
  assign new_E6543_ = ~new_E6507_ & new_E6542_;
  assign new_E6544_ = new_E6563_ | new_E6562_;
  assign new_E6545_ = new_E6507_ & new_E6544_;
  assign new_E6546_ = new_E6505_ & ~new_E6515_;
  assign new_E6547_ = ~new_E6505_ & new_E6515_;
  assign new_E6548_ = ~new_E6504_ | ~new_E6529_;
  assign new_E6549_ = new_E6515_ & new_E6548_;
  assign new_E6550_ = ~new_E6515_ & ~new_E6549_;
  assign new_E6551_ = new_E6515_ | new_E6548_;
  assign new_E6552_ = ~new_E6505_ & new_E6506_;
  assign new_E6553_ = new_E6505_ & ~new_E6506_;
  assign new_E6554_ = new_E6522_ | new_E6559_;
  assign new_E6555_ = ~new_E6522_ & ~new_E6558_;
  assign new_E6556_ = new_E6505_ | new_E6522_;
  assign new_E6557_ = new_E6505_ | new_E6506_;
  assign new_E6558_ = new_E6522_ & new_E6559_;
  assign new_E6559_ = ~new_E6504_ | ~new_E6529_;
  assign new_E6560_ = new_E6537_ & new_E6557_;
  assign new_E6561_ = ~new_E6537_ & ~new_E6557_;
  assign new_E6562_ = new_E6566_ | new_E6567_;
  assign new_E6563_ = ~new_E6508_ & new_E6522_;
  assign new_E6564_ = new_E6568_ | new_E6569_;
  assign new_E6565_ = new_E6508_ & new_E6522_;
  assign new_E6566_ = ~new_E6508_ & ~new_E6522_;
  assign new_E6567_ = new_E6508_ & ~new_E6522_;
  assign new_E6568_ = new_E6508_ & ~new_E6522_;
  assign new_E6569_ = ~new_E6508_ & new_E6522_;
  assign new_E6570_ = new_G5542_;
  assign new_E6571_ = new_G5609_;
  assign new_E6572_ = new_G5676_;
  assign new_E6573_ = new_G5743_;
  assign new_E6574_ = new_G5810_;
  assign new_E6575_ = new_G5877_;
  assign new_E6576_ = new_E6583_ & new_E6582_;
  assign new_E6577_ = new_E6585_ | new_E6584_;
  assign new_E6578_ = new_E6587_ | new_E6586_;
  assign new_E6579_ = new_E6589_ & new_E6588_;
  assign new_E6580_ = new_E6589_ & new_E6590_;
  assign new_E6581_ = new_E6582_ | new_E6591_;
  assign new_E6582_ = new_E6571_ | new_E6594_;
  assign new_E6583_ = new_E6593_ | new_E6592_;
  assign new_E6584_ = new_E6598_ & new_E6597_;
  assign new_E6585_ = new_E6596_ & new_E6595_;
  assign new_E6586_ = new_E6601_ | new_E6600_;
  assign new_E6587_ = new_E6596_ & new_E6599_;
  assign new_E6588_ = new_E6571_ | new_E6604_;
  assign new_E6589_ = new_E6603_ | new_E6602_;
  assign new_E6590_ = new_E6606_ | new_E6605_;
  assign new_E6591_ = ~new_E6582_ & new_E6608_;
  assign new_E6592_ = ~new_E6584_ & new_E6596_;
  assign new_E6593_ = new_E6584_ & ~new_E6596_;
  assign new_E6594_ = new_E6570_ & ~new_E6571_;
  assign new_E6595_ = ~new_E6617_ | ~new_E6618_;
  assign new_E6596_ = new_E6610_ | new_E6612_;
  assign new_E6597_ = new_E6620_ | new_E6619_;
  assign new_E6598_ = new_E6614_ | new_E6613_;
  assign new_E6599_ = ~new_E6622_ | ~new_E6621_;
  assign new_E6600_ = ~new_E6623_ & new_E6624_;
  assign new_E6601_ = new_E6623_ & ~new_E6624_;
  assign new_E6602_ = ~new_E6570_ & new_E6571_;
  assign new_E6603_ = new_E6570_ & ~new_E6571_;
  assign new_E6604_ = ~new_E6586_ | new_E6596_;
  assign new_E6605_ = new_E6586_ & new_E6596_;
  assign new_E6606_ = ~new_E6586_ & ~new_E6596_;
  assign new_E6607_ = new_E6628_ | new_E6627_;
  assign new_E6608_ = new_E6574_ | new_E6607_;
  assign new_E6609_ = new_E6632_ | new_E6631_;
  assign new_E6610_ = ~new_E6574_ & new_E6609_;
  assign new_E6611_ = new_E6630_ | new_E6629_;
  assign new_E6612_ = new_E6574_ & new_E6611_;
  assign new_E6613_ = new_E6572_ & ~new_E6582_;
  assign new_E6614_ = ~new_E6572_ & new_E6582_;
  assign new_E6615_ = ~new_E6571_ | ~new_E6596_;
  assign new_E6616_ = new_E6582_ & new_E6615_;
  assign new_E6617_ = ~new_E6582_ & ~new_E6616_;
  assign new_E6618_ = new_E6582_ | new_E6615_;
  assign new_E6619_ = ~new_E6572_ & new_E6573_;
  assign new_E6620_ = new_E6572_ & ~new_E6573_;
  assign new_E6621_ = new_E6589_ | new_E6626_;
  assign new_E6622_ = ~new_E6589_ & ~new_E6625_;
  assign new_E6623_ = new_E6572_ | new_E6589_;
  assign new_E6624_ = new_E6572_ | new_E6573_;
  assign new_E6625_ = new_E6589_ & new_E6626_;
  assign new_E6626_ = ~new_E6571_ | ~new_E6596_;
  assign new_E6627_ = new_E6604_ & new_E6624_;
  assign new_E6628_ = ~new_E6604_ & ~new_E6624_;
  assign new_E6629_ = new_E6633_ | new_E6634_;
  assign new_E6630_ = ~new_E6575_ & new_E6589_;
  assign new_E6631_ = new_E6635_ | new_E6636_;
  assign new_E6632_ = new_E6575_ & new_E6589_;
  assign new_E6633_ = ~new_E6575_ & ~new_E6589_;
  assign new_E6634_ = new_E6575_ & ~new_E6589_;
  assign new_E6635_ = new_E6575_ & ~new_E6589_;
  assign new_E6636_ = ~new_E6575_ & new_E6589_;
  assign new_E6637_ = new_F1469_;
  assign new_E6638_ = new_F1539_;
  assign new_E6639_ = new_F1606_;
  assign new_E6640_ = new_F1673_;
  assign new_E6641_ = new_F1740_;
  assign new_E6642_ = new_F1807_;
  assign new_E6643_ = new_E6650_ & new_E6649_;
  assign new_E6644_ = new_E6652_ | new_E6651_;
  assign new_E6645_ = new_E6654_ | new_E6653_;
  assign new_E6646_ = new_E6656_ & new_E6655_;
  assign new_E6647_ = new_E6656_ & new_E6657_;
  assign new_E6648_ = new_E6649_ | new_E6658_;
  assign new_E6649_ = new_E6638_ | new_E6661_;
  assign new_E6650_ = new_E6660_ | new_E6659_;
  assign new_E6651_ = new_E6665_ & new_E6664_;
  assign new_E6652_ = new_E6663_ & new_E6662_;
  assign new_E6653_ = new_E6668_ | new_E6667_;
  assign new_E6654_ = new_E6663_ & new_E6666_;
  assign new_E6655_ = new_E6638_ | new_E6671_;
  assign new_E6656_ = new_E6670_ | new_E6669_;
  assign new_E6657_ = new_E6673_ | new_E6672_;
  assign new_E6658_ = ~new_E6649_ & new_E6675_;
  assign new_E6659_ = ~new_E6651_ & new_E6663_;
  assign new_E6660_ = new_E6651_ & ~new_E6663_;
  assign new_E6661_ = new_E6637_ & ~new_E6638_;
  assign new_E6662_ = ~new_E6684_ | ~new_E6685_;
  assign new_E6663_ = new_E6677_ | new_E6679_;
  assign new_E6664_ = new_E6687_ | new_E6686_;
  assign new_E6665_ = new_E6681_ | new_E6680_;
  assign new_E6666_ = ~new_E6689_ | ~new_E6688_;
  assign new_E6667_ = ~new_E6690_ & new_E6691_;
  assign new_E6668_ = new_E6690_ & ~new_E6691_;
  assign new_E6669_ = ~new_E6637_ & new_E6638_;
  assign new_E6670_ = new_E6637_ & ~new_E6638_;
  assign new_E6671_ = ~new_E6653_ | new_E6663_;
  assign new_E6672_ = new_E6653_ & new_E6663_;
  assign new_E6673_ = ~new_E6653_ & ~new_E6663_;
  assign new_E6674_ = new_E6695_ | new_E6694_;
  assign new_E6675_ = new_E6641_ | new_E6674_;
  assign new_E6676_ = new_E6699_ | new_E6698_;
  assign new_E6677_ = ~new_E6641_ & new_E6676_;
  assign new_E6678_ = new_E6697_ | new_E6696_;
  assign new_E6679_ = new_E6641_ & new_E6678_;
  assign new_E6680_ = new_E6639_ & ~new_E6649_;
  assign new_E6681_ = ~new_E6639_ & new_E6649_;
  assign new_E6682_ = ~new_E6638_ | ~new_E6663_;
  assign new_E6683_ = new_E6649_ & new_E6682_;
  assign new_E6684_ = ~new_E6649_ & ~new_E6683_;
  assign new_E6685_ = new_E6649_ | new_E6682_;
  assign new_E6686_ = ~new_E6639_ & new_E6640_;
  assign new_E6687_ = new_E6639_ & ~new_E6640_;
  assign new_E6688_ = new_E6656_ | new_E6693_;
  assign new_E6689_ = ~new_E6656_ & ~new_E6692_;
  assign new_E6690_ = new_E6639_ | new_E6656_;
  assign new_E6691_ = new_E6639_ | new_E6640_;
  assign new_E6692_ = new_E6656_ & new_E6693_;
  assign new_E6693_ = ~new_E6638_ | ~new_E6663_;
  assign new_E6694_ = new_E6671_ & new_E6691_;
  assign new_E6695_ = ~new_E6671_ & ~new_E6691_;
  assign new_E6696_ = new_E6700_ | new_E6701_;
  assign new_E6697_ = ~new_E6642_ & new_E6656_;
  assign new_E6698_ = new_E6702_ | new_E6703_;
  assign new_E6699_ = new_E6642_ & new_E6656_;
  assign new_E6700_ = ~new_E6642_ & ~new_E6656_;
  assign new_E6701_ = new_E6642_ & ~new_E6656_;
  assign new_E6702_ = new_E6642_ & ~new_E6656_;
  assign new_E6703_ = ~new_E6642_ & new_E6656_;
  assign new_E6704_ = new_F1874_;
  assign new_E6705_ = new_F1941_;
  assign new_E6706_ = new_F2008_;
  assign new_E6707_ = new_F2075_;
  assign new_E6708_ = new_F2142_;
  assign new_E6709_ = new_F2209_;
  assign new_E6710_ = new_E6717_ & new_E6716_;
  assign new_E6711_ = new_E6719_ | new_E6718_;
  assign new_E6712_ = new_E6721_ | new_E6720_;
  assign new_E6713_ = new_E6723_ & new_E6722_;
  assign new_E6714_ = new_E6723_ & new_E6724_;
  assign new_E6715_ = new_E6716_ | new_E6725_;
  assign new_E6716_ = new_E6705_ | new_E6728_;
  assign new_E6717_ = new_E6727_ | new_E6726_;
  assign new_E6718_ = new_E6732_ & new_E6731_;
  assign new_E6719_ = new_E6730_ & new_E6729_;
  assign new_E6720_ = new_E6735_ | new_E6734_;
  assign new_E6721_ = new_E6730_ & new_E6733_;
  assign new_E6722_ = new_E6705_ | new_E6738_;
  assign new_E6723_ = new_E6737_ | new_E6736_;
  assign new_E6724_ = new_E6740_ | new_E6739_;
  assign new_E6725_ = ~new_E6716_ & new_E6742_;
  assign new_E6726_ = ~new_E6718_ & new_E6730_;
  assign new_E6727_ = new_E6718_ & ~new_E6730_;
  assign new_E6728_ = new_E6704_ & ~new_E6705_;
  assign new_E6729_ = ~new_E6751_ | ~new_E6752_;
  assign new_E6730_ = new_E6744_ | new_E6746_;
  assign new_E6731_ = new_E6754_ | new_E6753_;
  assign new_E6732_ = new_E6748_ | new_E6747_;
  assign new_E6733_ = ~new_E6756_ | ~new_E6755_;
  assign new_E6734_ = ~new_E6757_ & new_E6758_;
  assign new_E6735_ = new_E6757_ & ~new_E6758_;
  assign new_E6736_ = ~new_E6704_ & new_E6705_;
  assign new_E6737_ = new_E6704_ & ~new_E6705_;
  assign new_E6738_ = ~new_E6720_ | new_E6730_;
  assign new_E6739_ = new_E6720_ & new_E6730_;
  assign new_E6740_ = ~new_E6720_ & ~new_E6730_;
  assign new_E6741_ = new_E6762_ | new_E6761_;
  assign new_E6742_ = new_E6708_ | new_E6741_;
  assign new_E6743_ = new_E6766_ | new_E6765_;
  assign new_E6744_ = ~new_E6708_ & new_E6743_;
  assign new_E6745_ = new_E6764_ | new_E6763_;
  assign new_E6746_ = new_E6708_ & new_E6745_;
  assign new_E6747_ = new_E6706_ & ~new_E6716_;
  assign new_E6748_ = ~new_E6706_ & new_E6716_;
  assign new_E6749_ = ~new_E6705_ | ~new_E6730_;
  assign new_E6750_ = new_E6716_ & new_E6749_;
  assign new_E6751_ = ~new_E6716_ & ~new_E6750_;
  assign new_E6752_ = new_E6716_ | new_E6749_;
  assign new_E6753_ = ~new_E6706_ & new_E6707_;
  assign new_E6754_ = new_E6706_ & ~new_E6707_;
  assign new_E6755_ = new_E6723_ | new_E6760_;
  assign new_E6756_ = ~new_E6723_ & ~new_E6759_;
  assign new_E6757_ = new_E6706_ | new_E6723_;
  assign new_E6758_ = new_E6706_ | new_E6707_;
  assign new_E6759_ = new_E6723_ & new_E6760_;
  assign new_E6760_ = ~new_E6705_ | ~new_E6730_;
  assign new_E6761_ = new_E6738_ & new_E6758_;
  assign new_E6762_ = ~new_E6738_ & ~new_E6758_;
  assign new_E6763_ = new_E6767_ | new_E6768_;
  assign new_E6764_ = ~new_E6709_ & new_E6723_;
  assign new_E6765_ = new_E6769_ | new_E6770_;
  assign new_E6766_ = new_E6709_ & new_E6723_;
  assign new_E6767_ = ~new_E6709_ & ~new_E6723_;
  assign new_E6768_ = new_E6709_ & ~new_E6723_;
  assign new_E6769_ = new_E6709_ & ~new_E6723_;
  assign new_E6770_ = ~new_E6709_ & new_E6723_;
  assign new_E6771_ = new_F2276_;
  assign new_E6772_ = new_F2343_;
  assign new_E6773_ = new_F2410_;
  assign new_E6774_ = new_F2477_;
  assign new_E6775_ = new_F2544_;
  assign new_E6776_ = new_F2611_;
  assign new_E6777_ = new_E6784_ & new_E6783_;
  assign new_E6778_ = new_E6786_ | new_E6785_;
  assign new_E6779_ = new_E6788_ | new_E6787_;
  assign new_E6780_ = new_E6790_ & new_E6789_;
  assign new_E6781_ = new_E6790_ & new_E6791_;
  assign new_E6782_ = new_E6783_ | new_E6792_;
  assign new_E6783_ = new_E6772_ | new_E6795_;
  assign new_E6784_ = new_E6794_ | new_E6793_;
  assign new_E6785_ = new_E6799_ & new_E6798_;
  assign new_E6786_ = new_E6797_ & new_E6796_;
  assign new_E6787_ = new_E6802_ | new_E6801_;
  assign new_E6788_ = new_E6797_ & new_E6800_;
  assign new_E6789_ = new_E6772_ | new_E6805_;
  assign new_E6790_ = new_E6804_ | new_E6803_;
  assign new_E6791_ = new_E6807_ | new_E6806_;
  assign new_E6792_ = ~new_E6783_ & new_E6809_;
  assign new_E6793_ = ~new_E6785_ & new_E6797_;
  assign new_E6794_ = new_E6785_ & ~new_E6797_;
  assign new_E6795_ = new_E6771_ & ~new_E6772_;
  assign new_E6796_ = ~new_E6818_ | ~new_E6819_;
  assign new_E6797_ = new_E6811_ | new_E6813_;
  assign new_E6798_ = new_E6821_ | new_E6820_;
  assign new_E6799_ = new_E6815_ | new_E6814_;
  assign new_E6800_ = ~new_E6823_ | ~new_E6822_;
  assign new_E6801_ = ~new_E6824_ & new_E6825_;
  assign new_E6802_ = new_E6824_ & ~new_E6825_;
  assign new_E6803_ = ~new_E6771_ & new_E6772_;
  assign new_E6804_ = new_E6771_ & ~new_E6772_;
  assign new_E6805_ = ~new_E6787_ | new_E6797_;
  assign new_E6806_ = new_E6787_ & new_E6797_;
  assign new_E6807_ = ~new_E6787_ & ~new_E6797_;
  assign new_E6808_ = new_E6829_ | new_E6828_;
  assign new_E6809_ = new_E6775_ | new_E6808_;
  assign new_E6810_ = new_E6833_ | new_E6832_;
  assign new_E6811_ = ~new_E6775_ & new_E6810_;
  assign new_E6812_ = new_E6831_ | new_E6830_;
  assign new_E6813_ = new_E6775_ & new_E6812_;
  assign new_E6814_ = new_E6773_ & ~new_E6783_;
  assign new_E6815_ = ~new_E6773_ & new_E6783_;
  assign new_E6816_ = ~new_E6772_ | ~new_E6797_;
  assign new_E6817_ = new_E6783_ & new_E6816_;
  assign new_E6818_ = ~new_E6783_ & ~new_E6817_;
  assign new_E6819_ = new_E6783_ | new_E6816_;
  assign new_E6820_ = ~new_E6773_ & new_E6774_;
  assign new_E6821_ = new_E6773_ & ~new_E6774_;
  assign new_E6822_ = new_E6790_ | new_E6827_;
  assign new_E6823_ = ~new_E6790_ & ~new_E6826_;
  assign new_E6824_ = new_E6773_ | new_E6790_;
  assign new_E6825_ = new_E6773_ | new_E6774_;
  assign new_E6826_ = new_E6790_ & new_E6827_;
  assign new_E6827_ = ~new_E6772_ | ~new_E6797_;
  assign new_E6828_ = new_E6805_ & new_E6825_;
  assign new_E6829_ = ~new_E6805_ & ~new_E6825_;
  assign new_E6830_ = new_E6834_ | new_E6835_;
  assign new_E6831_ = ~new_E6776_ & new_E6790_;
  assign new_E6832_ = new_E6836_ | new_E6837_;
  assign new_E6833_ = new_E6776_ & new_E6790_;
  assign new_E6834_ = ~new_E6776_ & ~new_E6790_;
  assign new_E6835_ = new_E6776_ & ~new_E6790_;
  assign new_E6836_ = new_E6776_ & ~new_E6790_;
  assign new_E6837_ = ~new_E6776_ & new_E6790_;
  assign new_E6838_ = new_F2678_;
  assign new_E6839_ = new_F2745_;
  assign new_E6840_ = new_F2812_;
  assign new_E6841_ = new_F2879_;
  assign new_E6842_ = new_F2946_;
  assign new_E6843_ = new_F3013_;
  assign new_E6844_ = new_E6851_ & new_E6850_;
  assign new_E6845_ = new_E6853_ | new_E6852_;
  assign new_E6846_ = new_E6855_ | new_E6854_;
  assign new_E6847_ = new_E6857_ & new_E6856_;
  assign new_E6848_ = new_E6857_ & new_E6858_;
  assign new_E6849_ = new_E6850_ | new_E6859_;
  assign new_E6850_ = new_E6839_ | new_E6862_;
  assign new_E6851_ = new_E6861_ | new_E6860_;
  assign new_E6852_ = new_E6866_ & new_E6865_;
  assign new_E6853_ = new_E6864_ & new_E6863_;
  assign new_E6854_ = new_E6869_ | new_E6868_;
  assign new_E6855_ = new_E6864_ & new_E6867_;
  assign new_E6856_ = new_E6839_ | new_E6872_;
  assign new_E6857_ = new_E6871_ | new_E6870_;
  assign new_E6858_ = new_E6874_ | new_E6873_;
  assign new_E6859_ = ~new_E6850_ & new_E6876_;
  assign new_E6860_ = ~new_E6852_ & new_E6864_;
  assign new_E6861_ = new_E6852_ & ~new_E6864_;
  assign new_E6862_ = new_E6838_ & ~new_E6839_;
  assign new_E6863_ = ~new_E6885_ | ~new_E6886_;
  assign new_E6864_ = new_E6878_ | new_E6880_;
  assign new_E6865_ = new_E6888_ | new_E6887_;
  assign new_E6866_ = new_E6882_ | new_E6881_;
  assign new_E6867_ = ~new_E6890_ | ~new_E6889_;
  assign new_E6868_ = ~new_E6891_ & new_E6892_;
  assign new_E6869_ = new_E6891_ & ~new_E6892_;
  assign new_E6870_ = ~new_E6838_ & new_E6839_;
  assign new_E6871_ = new_E6838_ & ~new_E6839_;
  assign new_E6872_ = ~new_E6854_ | new_E6864_;
  assign new_E6873_ = new_E6854_ & new_E6864_;
  assign new_E6874_ = ~new_E6854_ & ~new_E6864_;
  assign new_E6875_ = new_E6896_ | new_E6895_;
  assign new_E6876_ = new_E6842_ | new_E6875_;
  assign new_E6877_ = new_E6900_ | new_E6899_;
  assign new_E6878_ = ~new_E6842_ & new_E6877_;
  assign new_E6879_ = new_E6898_ | new_E6897_;
  assign new_E6880_ = new_E6842_ & new_E6879_;
  assign new_E6881_ = new_E6840_ & ~new_E6850_;
  assign new_E6882_ = ~new_E6840_ & new_E6850_;
  assign new_E6883_ = ~new_E6839_ | ~new_E6864_;
  assign new_E6884_ = new_E6850_ & new_E6883_;
  assign new_E6885_ = ~new_E6850_ & ~new_E6884_;
  assign new_E6886_ = new_E6850_ | new_E6883_;
  assign new_E6887_ = ~new_E6840_ & new_E6841_;
  assign new_E6888_ = new_E6840_ & ~new_E6841_;
  assign new_E6889_ = new_E6857_ | new_E6894_;
  assign new_E6890_ = ~new_E6857_ & ~new_E6893_;
  assign new_E6891_ = new_E6840_ | new_E6857_;
  assign new_E6892_ = new_E6840_ | new_E6841_;
  assign new_E6893_ = new_E6857_ & new_E6894_;
  assign new_E6894_ = ~new_E6839_ | ~new_E6864_;
  assign new_E6895_ = new_E6872_ & new_E6892_;
  assign new_E6896_ = ~new_E6872_ & ~new_E6892_;
  assign new_E6897_ = new_E6901_ | new_E6902_;
  assign new_E6898_ = ~new_E6843_ & new_E6857_;
  assign new_E6899_ = new_E6903_ | new_E6904_;
  assign new_E6900_ = new_E6843_ & new_E6857_;
  assign new_E6901_ = ~new_E6843_ & ~new_E6857_;
  assign new_E6902_ = new_E6843_ & ~new_E6857_;
  assign new_E6903_ = new_E6843_ & ~new_E6857_;
  assign new_E6904_ = ~new_E6843_ & new_E6857_;
  assign new_E6905_ = new_F3080_;
  assign new_E6906_ = new_F3147_;
  assign new_E6907_ = new_F3214_;
  assign new_E6908_ = new_F3281_;
  assign new_E6909_ = new_F3348_;
  assign new_E6910_ = new_F3415_;
  assign new_E6911_ = new_E6918_ & new_E6917_;
  assign new_E6912_ = new_E6920_ | new_E6919_;
  assign new_E6913_ = new_E6922_ | new_E6921_;
  assign new_E6914_ = new_E6924_ & new_E6923_;
  assign new_E6915_ = new_E6924_ & new_E6925_;
  assign new_E6916_ = new_E6917_ | new_E6926_;
  assign new_E6917_ = new_E6906_ | new_E6929_;
  assign new_E6918_ = new_E6928_ | new_E6927_;
  assign new_E6919_ = new_E6933_ & new_E6932_;
  assign new_E6920_ = new_E6931_ & new_E6930_;
  assign new_E6921_ = new_E6936_ | new_E6935_;
  assign new_E6922_ = new_E6931_ & new_E6934_;
  assign new_E6923_ = new_E6906_ | new_E6939_;
  assign new_E6924_ = new_E6938_ | new_E6937_;
  assign new_E6925_ = new_E6941_ | new_E6940_;
  assign new_E6926_ = ~new_E6917_ & new_E6943_;
  assign new_E6927_ = ~new_E6919_ & new_E6931_;
  assign new_E6928_ = new_E6919_ & ~new_E6931_;
  assign new_E6929_ = new_E6905_ & ~new_E6906_;
  assign new_E6930_ = ~new_E6952_ | ~new_E6953_;
  assign new_E6931_ = new_E6945_ | new_E6947_;
  assign new_E6932_ = new_E6955_ | new_E6954_;
  assign new_E6933_ = new_E6949_ | new_E6948_;
  assign new_E6934_ = ~new_E6957_ | ~new_E6956_;
  assign new_E6935_ = ~new_E6958_ & new_E6959_;
  assign new_E6936_ = new_E6958_ & ~new_E6959_;
  assign new_E6937_ = ~new_E6905_ & new_E6906_;
  assign new_E6938_ = new_E6905_ & ~new_E6906_;
  assign new_E6939_ = ~new_E6921_ | new_E6931_;
  assign new_E6940_ = new_E6921_ & new_E6931_;
  assign new_E6941_ = ~new_E6921_ & ~new_E6931_;
  assign new_E6942_ = new_E6963_ | new_E6962_;
  assign new_E6943_ = new_E6909_ | new_E6942_;
  assign new_E6944_ = new_E6967_ | new_E6966_;
  assign new_E6945_ = ~new_E6909_ & new_E6944_;
  assign new_E6946_ = new_E6965_ | new_E6964_;
  assign new_E6947_ = new_E6909_ & new_E6946_;
  assign new_E6948_ = new_E6907_ & ~new_E6917_;
  assign new_E6949_ = ~new_E6907_ & new_E6917_;
  assign new_E6950_ = ~new_E6906_ | ~new_E6931_;
  assign new_E6951_ = new_E6917_ & new_E6950_;
  assign new_E6952_ = ~new_E6917_ & ~new_E6951_;
  assign new_E6953_ = new_E6917_ | new_E6950_;
  assign new_E6954_ = ~new_E6907_ & new_E6908_;
  assign new_E6955_ = new_E6907_ & ~new_E6908_;
  assign new_E6956_ = new_E6924_ | new_E6961_;
  assign new_E6957_ = ~new_E6924_ & ~new_E6960_;
  assign new_E6958_ = new_E6907_ | new_E6924_;
  assign new_E6959_ = new_E6907_ | new_E6908_;
  assign new_E6960_ = new_E6924_ & new_E6961_;
  assign new_E6961_ = ~new_E6906_ | ~new_E6931_;
  assign new_E6962_ = new_E6939_ & new_E6959_;
  assign new_E6963_ = ~new_E6939_ & ~new_E6959_;
  assign new_E6964_ = new_E6968_ | new_E6969_;
  assign new_E6965_ = ~new_E6910_ & new_E6924_;
  assign new_E6966_ = new_E6970_ | new_E6971_;
  assign new_E6967_ = new_E6910_ & new_E6924_;
  assign new_E6968_ = ~new_E6910_ & ~new_E6924_;
  assign new_E6969_ = new_E6910_ & ~new_E6924_;
  assign new_E6970_ = new_E6910_ & ~new_E6924_;
  assign new_E6971_ = ~new_E6910_ & new_E6924_;
  assign new_E6972_ = new_F3482_;
  assign new_E6973_ = new_F3549_;
  assign new_E6974_ = new_F3616_;
  assign new_E6975_ = new_F3683_;
  assign new_E6976_ = new_F3750_;
  assign new_E6977_ = new_F3817_;
  assign new_E6978_ = new_E6985_ & new_E6984_;
  assign new_E6979_ = new_E6987_ | new_E6986_;
  assign new_E6980_ = new_E6989_ | new_E6988_;
  assign new_E6981_ = new_E6991_ & new_E6990_;
  assign new_E6982_ = new_E6991_ & new_E6992_;
  assign new_E6983_ = new_E6984_ | new_E6993_;
  assign new_E6984_ = new_E6973_ | new_E6996_;
  assign new_E6985_ = new_E6995_ | new_E6994_;
  assign new_E6986_ = new_E7000_ & new_E6999_;
  assign new_E6987_ = new_E6998_ & new_E6997_;
  assign new_E6988_ = new_E7003_ | new_E7002_;
  assign new_E6989_ = new_E6998_ & new_E7001_;
  assign new_E6990_ = new_E6973_ | new_E7006_;
  assign new_E6991_ = new_E7005_ | new_E7004_;
  assign new_E6992_ = new_E7008_ | new_E7007_;
  assign new_E6993_ = ~new_E6984_ & new_E7010_;
  assign new_E6994_ = ~new_E6986_ & new_E6998_;
  assign new_E6995_ = new_E6986_ & ~new_E6998_;
  assign new_E6996_ = new_E6972_ & ~new_E6973_;
  assign new_E6997_ = ~new_E7019_ | ~new_E7020_;
  assign new_E6998_ = new_E7012_ | new_E7014_;
  assign new_E6999_ = new_E7022_ | new_E7021_;
  assign new_E7000_ = new_E7016_ | new_E7015_;
  assign new_E7001_ = ~new_E7024_ | ~new_E7023_;
  assign new_E7002_ = ~new_E7025_ & new_E7026_;
  assign new_E7003_ = new_E7025_ & ~new_E7026_;
  assign new_E7004_ = ~new_E6972_ & new_E6973_;
  assign new_E7005_ = new_E6972_ & ~new_E6973_;
  assign new_E7006_ = ~new_E6988_ | new_E6998_;
  assign new_E7007_ = new_E6988_ & new_E6998_;
  assign new_E7008_ = ~new_E6988_ & ~new_E6998_;
  assign new_E7009_ = new_E7030_ | new_E7029_;
  assign new_E7010_ = new_E6976_ | new_E7009_;
  assign new_E7011_ = new_E7034_ | new_E7033_;
  assign new_E7012_ = ~new_E6976_ & new_E7011_;
  assign new_E7013_ = new_E7032_ | new_E7031_;
  assign new_E7014_ = new_E6976_ & new_E7013_;
  assign new_E7015_ = new_E6974_ & ~new_E6984_;
  assign new_E7016_ = ~new_E6974_ & new_E6984_;
  assign new_E7017_ = ~new_E6973_ | ~new_E6998_;
  assign new_E7018_ = new_E6984_ & new_E7017_;
  assign new_E7019_ = ~new_E6984_ & ~new_E7018_;
  assign new_E7020_ = new_E6984_ | new_E7017_;
  assign new_E7021_ = ~new_E6974_ & new_E6975_;
  assign new_E7022_ = new_E6974_ & ~new_E6975_;
  assign new_E7023_ = new_E6991_ | new_E7028_;
  assign new_E7024_ = ~new_E6991_ & ~new_E7027_;
  assign new_E7025_ = new_E6974_ | new_E6991_;
  assign new_E7026_ = new_E6974_ | new_E6975_;
  assign new_E7027_ = new_E6991_ & new_E7028_;
  assign new_E7028_ = ~new_E6973_ | ~new_E6998_;
  assign new_E7029_ = new_E7006_ & new_E7026_;
  assign new_E7030_ = ~new_E7006_ & ~new_E7026_;
  assign new_E7031_ = new_E7035_ | new_E7036_;
  assign new_E7032_ = ~new_E6977_ & new_E6991_;
  assign new_E7033_ = new_E7037_ | new_E7038_;
  assign new_E7034_ = new_E6977_ & new_E6991_;
  assign new_E7035_ = ~new_E6977_ & ~new_E6991_;
  assign new_E7036_ = new_E6977_ & ~new_E6991_;
  assign new_E7037_ = new_E6977_ & ~new_E6991_;
  assign new_E7038_ = ~new_E6977_ & new_E6991_;
  assign new_E7039_ = new_F3884_;
  assign new_E7040_ = new_F3951_;
  assign new_E7041_ = new_F4018_;
  assign new_E7042_ = new_F4085_;
  assign new_E7043_ = new_F4152_;
  assign new_E7044_ = new_F4219_;
  assign new_E7045_ = new_E7052_ & new_E7051_;
  assign new_E7046_ = new_E7054_ | new_E7053_;
  assign new_E7047_ = new_E7056_ | new_E7055_;
  assign new_E7048_ = new_E7058_ & new_E7057_;
  assign new_E7049_ = new_E7058_ & new_E7059_;
  assign new_E7050_ = new_E7051_ | new_E7060_;
  assign new_E7051_ = new_E7040_ | new_E7063_;
  assign new_E7052_ = new_E7062_ | new_E7061_;
  assign new_E7053_ = new_E7067_ & new_E7066_;
  assign new_E7054_ = new_E7065_ & new_E7064_;
  assign new_E7055_ = new_E7070_ | new_E7069_;
  assign new_E7056_ = new_E7065_ & new_E7068_;
  assign new_E7057_ = new_E7040_ | new_E7073_;
  assign new_E7058_ = new_E7072_ | new_E7071_;
  assign new_E7059_ = new_E7075_ | new_E7074_;
  assign new_E7060_ = ~new_E7051_ & new_E7077_;
  assign new_E7061_ = ~new_E7053_ & new_E7065_;
  assign new_E7062_ = new_E7053_ & ~new_E7065_;
  assign new_E7063_ = new_E7039_ & ~new_E7040_;
  assign new_E7064_ = ~new_E7086_ | ~new_E7087_;
  assign new_E7065_ = new_E7079_ | new_E7081_;
  assign new_E7066_ = new_E7089_ | new_E7088_;
  assign new_E7067_ = new_E7083_ | new_E7082_;
  assign new_E7068_ = ~new_E7091_ | ~new_E7090_;
  assign new_E7069_ = ~new_E7092_ & new_E7093_;
  assign new_E7070_ = new_E7092_ & ~new_E7093_;
  assign new_E7071_ = ~new_E7039_ & new_E7040_;
  assign new_E7072_ = new_E7039_ & ~new_E7040_;
  assign new_E7073_ = ~new_E7055_ | new_E7065_;
  assign new_E7074_ = new_E7055_ & new_E7065_;
  assign new_E7075_ = ~new_E7055_ & ~new_E7065_;
  assign new_E7076_ = new_E7097_ | new_E7096_;
  assign new_E7077_ = new_E7043_ | new_E7076_;
  assign new_E7078_ = new_E7101_ | new_E7100_;
  assign new_E7079_ = ~new_E7043_ & new_E7078_;
  assign new_E7080_ = new_E7099_ | new_E7098_;
  assign new_E7081_ = new_E7043_ & new_E7080_;
  assign new_E7082_ = new_E7041_ & ~new_E7051_;
  assign new_E7083_ = ~new_E7041_ & new_E7051_;
  assign new_E7084_ = ~new_E7040_ | ~new_E7065_;
  assign new_E7085_ = new_E7051_ & new_E7084_;
  assign new_E7086_ = ~new_E7051_ & ~new_E7085_;
  assign new_E7087_ = new_E7051_ | new_E7084_;
  assign new_E7088_ = ~new_E7041_ & new_E7042_;
  assign new_E7089_ = new_E7041_ & ~new_E7042_;
  assign new_E7090_ = new_E7058_ | new_E7095_;
  assign new_E7091_ = ~new_E7058_ & ~new_E7094_;
  assign new_E7092_ = new_E7041_ | new_E7058_;
  assign new_E7093_ = new_E7041_ | new_E7042_;
  assign new_E7094_ = new_E7058_ & new_E7095_;
  assign new_E7095_ = ~new_E7040_ | ~new_E7065_;
  assign new_E7096_ = new_E7073_ & new_E7093_;
  assign new_E7097_ = ~new_E7073_ & ~new_E7093_;
  assign new_E7098_ = new_E7102_ | new_E7103_;
  assign new_E7099_ = ~new_E7044_ & new_E7058_;
  assign new_E7100_ = new_E7104_ | new_E7105_;
  assign new_E7101_ = new_E7044_ & new_E7058_;
  assign new_E7102_ = ~new_E7044_ & ~new_E7058_;
  assign new_E7103_ = new_E7044_ & ~new_E7058_;
  assign new_E7104_ = new_E7044_ & ~new_E7058_;
  assign new_E7105_ = ~new_E7044_ & new_E7058_;
  assign new_E7106_ = new_F4286_;
  assign new_E7107_ = new_F4353_;
  assign new_E7108_ = new_F4420_;
  assign new_E7109_ = new_F4487_;
  assign new_E7110_ = new_F4554_;
  assign new_E7111_ = new_F4621_;
  assign new_E7112_ = new_E7119_ & new_E7118_;
  assign new_E7113_ = new_E7121_ | new_E7120_;
  assign new_E7114_ = new_E7123_ | new_E7122_;
  assign new_E7115_ = new_E7125_ & new_E7124_;
  assign new_E7116_ = new_E7125_ & new_E7126_;
  assign new_E7117_ = new_E7118_ | new_E7127_;
  assign new_E7118_ = new_E7107_ | new_E7130_;
  assign new_E7119_ = new_E7129_ | new_E7128_;
  assign new_E7120_ = new_E7134_ & new_E7133_;
  assign new_E7121_ = new_E7132_ & new_E7131_;
  assign new_E7122_ = new_E7137_ | new_E7136_;
  assign new_E7123_ = new_E7132_ & new_E7135_;
  assign new_E7124_ = new_E7107_ | new_E7140_;
  assign new_E7125_ = new_E7139_ | new_E7138_;
  assign new_E7126_ = new_E7142_ | new_E7141_;
  assign new_E7127_ = ~new_E7118_ & new_E7144_;
  assign new_E7128_ = ~new_E7120_ & new_E7132_;
  assign new_E7129_ = new_E7120_ & ~new_E7132_;
  assign new_E7130_ = new_E7106_ & ~new_E7107_;
  assign new_E7131_ = ~new_E7153_ | ~new_E7154_;
  assign new_E7132_ = new_E7146_ | new_E7148_;
  assign new_E7133_ = new_E7156_ | new_E7155_;
  assign new_E7134_ = new_E7150_ | new_E7149_;
  assign new_E7135_ = ~new_E7158_ | ~new_E7157_;
  assign new_E7136_ = ~new_E7159_ & new_E7160_;
  assign new_E7137_ = new_E7159_ & ~new_E7160_;
  assign new_E7138_ = ~new_E7106_ & new_E7107_;
  assign new_E7139_ = new_E7106_ & ~new_E7107_;
  assign new_E7140_ = ~new_E7122_ | new_E7132_;
  assign new_E7141_ = new_E7122_ & new_E7132_;
  assign new_E7142_ = ~new_E7122_ & ~new_E7132_;
  assign new_E7143_ = new_E7164_ | new_E7163_;
  assign new_E7144_ = new_E7110_ | new_E7143_;
  assign new_E7145_ = new_E7168_ | new_E7167_;
  assign new_E7146_ = ~new_E7110_ & new_E7145_;
  assign new_E7147_ = new_E7166_ | new_E7165_;
  assign new_E7148_ = new_E7110_ & new_E7147_;
  assign new_E7149_ = new_E7108_ & ~new_E7118_;
  assign new_E7150_ = ~new_E7108_ & new_E7118_;
  assign new_E7151_ = ~new_E7107_ | ~new_E7132_;
  assign new_E7152_ = new_E7118_ & new_E7151_;
  assign new_E7153_ = ~new_E7118_ & ~new_E7152_;
  assign new_E7154_ = new_E7118_ | new_E7151_;
  assign new_E7155_ = ~new_E7108_ & new_E7109_;
  assign new_E7156_ = new_E7108_ & ~new_E7109_;
  assign new_E7157_ = new_E7125_ | new_E7162_;
  assign new_E7158_ = ~new_E7125_ & ~new_E7161_;
  assign new_E7159_ = new_E7108_ | new_E7125_;
  assign new_E7160_ = new_E7108_ | new_E7109_;
  assign new_E7161_ = new_E7125_ & new_E7162_;
  assign new_E7162_ = ~new_E7107_ | ~new_E7132_;
  assign new_E7163_ = new_E7140_ & new_E7160_;
  assign new_E7164_ = ~new_E7140_ & ~new_E7160_;
  assign new_E7165_ = new_E7169_ | new_E7170_;
  assign new_E7166_ = ~new_E7111_ & new_E7125_;
  assign new_E7167_ = new_E7171_ | new_E7172_;
  assign new_E7168_ = new_E7111_ & new_E7125_;
  assign new_E7169_ = ~new_E7111_ & ~new_E7125_;
  assign new_E7170_ = new_E7111_ & ~new_E7125_;
  assign new_E7171_ = new_E7111_ & ~new_E7125_;
  assign new_E7172_ = ~new_E7111_ & new_E7125_;
  assign new_E7173_ = new_F4688_;
  assign new_E7174_ = new_F4755_;
  assign new_E7175_ = new_F4822_;
  assign new_E7176_ = new_F4889_;
  assign new_E7177_ = new_F4956_;
  assign new_E7178_ = new_F5023_;
  assign new_E7179_ = new_E7186_ & new_E7185_;
  assign new_E7180_ = new_E7188_ | new_E7187_;
  assign new_E7181_ = new_E7190_ | new_E7189_;
  assign new_E7182_ = new_E7192_ & new_E7191_;
  assign new_E7183_ = new_E7192_ & new_E7193_;
  assign new_E7184_ = new_E7185_ | new_E7194_;
  assign new_E7185_ = new_E7174_ | new_E7197_;
  assign new_E7186_ = new_E7196_ | new_E7195_;
  assign new_E7187_ = new_E7201_ & new_E7200_;
  assign new_E7188_ = new_E7199_ & new_E7198_;
  assign new_E7189_ = new_E7204_ | new_E7203_;
  assign new_E7190_ = new_E7199_ & new_E7202_;
  assign new_E7191_ = new_E7174_ | new_E7207_;
  assign new_E7192_ = new_E7206_ | new_E7205_;
  assign new_E7193_ = new_E7209_ | new_E7208_;
  assign new_E7194_ = ~new_E7185_ & new_E7211_;
  assign new_E7195_ = ~new_E7187_ & new_E7199_;
  assign new_E7196_ = new_E7187_ & ~new_E7199_;
  assign new_E7197_ = new_E7173_ & ~new_E7174_;
  assign new_E7198_ = ~new_E7220_ | ~new_E7221_;
  assign new_E7199_ = new_E7213_ | new_E7215_;
  assign new_E7200_ = new_E7223_ | new_E7222_;
  assign new_E7201_ = new_E7217_ | new_E7216_;
  assign new_E7202_ = ~new_E7225_ | ~new_E7224_;
  assign new_E7203_ = ~new_E7226_ & new_E7227_;
  assign new_E7204_ = new_E7226_ & ~new_E7227_;
  assign new_E7205_ = ~new_E7173_ & new_E7174_;
  assign new_E7206_ = new_E7173_ & ~new_E7174_;
  assign new_E7207_ = ~new_E7189_ | new_E7199_;
  assign new_E7208_ = new_E7189_ & new_E7199_;
  assign new_E7209_ = ~new_E7189_ & ~new_E7199_;
  assign new_E7210_ = new_E7231_ | new_E7230_;
  assign new_E7211_ = new_E7177_ | new_E7210_;
  assign new_E7212_ = new_E7235_ | new_E7234_;
  assign new_E7213_ = ~new_E7177_ & new_E7212_;
  assign new_E7214_ = new_E7233_ | new_E7232_;
  assign new_E7215_ = new_E7177_ & new_E7214_;
  assign new_E7216_ = new_E7175_ & ~new_E7185_;
  assign new_E7217_ = ~new_E7175_ & new_E7185_;
  assign new_E7218_ = ~new_E7174_ | ~new_E7199_;
  assign new_E7219_ = new_E7185_ & new_E7218_;
  assign new_E7220_ = ~new_E7185_ & ~new_E7219_;
  assign new_E7221_ = new_E7185_ | new_E7218_;
  assign new_E7222_ = ~new_E7175_ & new_E7176_;
  assign new_E7223_ = new_E7175_ & ~new_E7176_;
  assign new_E7224_ = new_E7192_ | new_E7229_;
  assign new_E7225_ = ~new_E7192_ & ~new_E7228_;
  assign new_E7226_ = new_E7175_ | new_E7192_;
  assign new_E7227_ = new_E7175_ | new_E7176_;
  assign new_E7228_ = new_E7192_ & new_E7229_;
  assign new_E7229_ = ~new_E7174_ | ~new_E7199_;
  assign new_E7230_ = new_E7207_ & new_E7227_;
  assign new_E7231_ = ~new_E7207_ & ~new_E7227_;
  assign new_E7232_ = new_E7236_ | new_E7237_;
  assign new_E7233_ = ~new_E7178_ & new_E7192_;
  assign new_E7234_ = new_E7238_ | new_E7239_;
  assign new_E7235_ = new_E7178_ & new_E7192_;
  assign new_E7236_ = ~new_E7178_ & ~new_E7192_;
  assign new_E7237_ = new_E7178_ & ~new_E7192_;
  assign new_E7238_ = new_E7178_ & ~new_E7192_;
  assign new_E7239_ = ~new_E7178_ & new_E7192_;
  assign new_E7240_ = new_F5090_;
  assign new_E7241_ = new_F5157_;
  assign new_E7242_ = new_F5224_;
  assign new_E7243_ = new_F5291_;
  assign new_E7244_ = new_F5358_;
  assign new_E7245_ = new_F5425_;
  assign new_E7246_ = new_E7253_ & new_E7252_;
  assign new_E7247_ = new_E7255_ | new_E7254_;
  assign new_E7248_ = new_E7257_ | new_E7256_;
  assign new_E7249_ = new_E7259_ & new_E7258_;
  assign new_E7250_ = new_E7259_ & new_E7260_;
  assign new_E7251_ = new_E7252_ | new_E7261_;
  assign new_E7252_ = new_E7241_ | new_E7264_;
  assign new_E7253_ = new_E7263_ | new_E7262_;
  assign new_E7254_ = new_E7268_ & new_E7267_;
  assign new_E7255_ = new_E7266_ & new_E7265_;
  assign new_E7256_ = new_E7271_ | new_E7270_;
  assign new_E7257_ = new_E7266_ & new_E7269_;
  assign new_E7258_ = new_E7241_ | new_E7274_;
  assign new_E7259_ = new_E7273_ | new_E7272_;
  assign new_E7260_ = new_E7276_ | new_E7275_;
  assign new_E7261_ = ~new_E7252_ & new_E7278_;
  assign new_E7262_ = ~new_E7254_ & new_E7266_;
  assign new_E7263_ = new_E7254_ & ~new_E7266_;
  assign new_E7264_ = new_E7240_ & ~new_E7241_;
  assign new_E7265_ = ~new_E7287_ | ~new_E7288_;
  assign new_E7266_ = new_E7280_ | new_E7282_;
  assign new_E7267_ = new_E7290_ | new_E7289_;
  assign new_E7268_ = new_E7284_ | new_E7283_;
  assign new_E7269_ = ~new_E7292_ | ~new_E7291_;
  assign new_E7270_ = ~new_E7293_ & new_E7294_;
  assign new_E7271_ = new_E7293_ & ~new_E7294_;
  assign new_E7272_ = ~new_E7240_ & new_E7241_;
  assign new_E7273_ = new_E7240_ & ~new_E7241_;
  assign new_E7274_ = ~new_E7256_ | new_E7266_;
  assign new_E7275_ = new_E7256_ & new_E7266_;
  assign new_E7276_ = ~new_E7256_ & ~new_E7266_;
  assign new_E7277_ = new_E7298_ | new_E7297_;
  assign new_E7278_ = new_E7244_ | new_E7277_;
  assign new_E7279_ = new_E7302_ | new_E7301_;
  assign new_E7280_ = ~new_E7244_ & new_E7279_;
  assign new_E7281_ = new_E7300_ | new_E7299_;
  assign new_E7282_ = new_E7244_ & new_E7281_;
  assign new_E7283_ = new_E7242_ & ~new_E7252_;
  assign new_E7284_ = ~new_E7242_ & new_E7252_;
  assign new_E7285_ = ~new_E7241_ | ~new_E7266_;
  assign new_E7286_ = new_E7252_ & new_E7285_;
  assign new_E7287_ = ~new_E7252_ & ~new_E7286_;
  assign new_E7288_ = new_E7252_ | new_E7285_;
  assign new_E7289_ = ~new_E7242_ & new_E7243_;
  assign new_E7290_ = new_E7242_ & ~new_E7243_;
  assign new_E7291_ = new_E7259_ | new_E7296_;
  assign new_E7292_ = ~new_E7259_ & ~new_E7295_;
  assign new_E7293_ = new_E7242_ | new_E7259_;
  assign new_E7294_ = new_E7242_ | new_E7243_;
  assign new_E7295_ = new_E7259_ & new_E7296_;
  assign new_E7296_ = ~new_E7241_ | ~new_E7266_;
  assign new_E7297_ = new_E7274_ & new_E7294_;
  assign new_E7298_ = ~new_E7274_ & ~new_E7294_;
  assign new_E7299_ = new_E7303_ | new_E7304_;
  assign new_E7300_ = ~new_E7245_ & new_E7259_;
  assign new_E7301_ = new_E7305_ | new_E7306_;
  assign new_E7302_ = new_E7245_ & new_E7259_;
  assign new_E7303_ = ~new_E7245_ & ~new_E7259_;
  assign new_E7304_ = new_E7245_ & ~new_E7259_;
  assign new_E7305_ = new_E7245_ & ~new_E7259_;
  assign new_E7306_ = ~new_E7245_ & new_E7259_;
  assign new_E7307_ = new_F5492_;
  assign new_E7308_ = new_F5559_;
  assign new_E7309_ = new_F5626_;
  assign new_E7310_ = new_F5693_;
  assign new_E7311_ = new_F5760_;
  assign new_E7312_ = new_F5827_;
  assign new_E7313_ = new_E7320_ & new_E7319_;
  assign new_E7314_ = new_E7322_ | new_E7321_;
  assign new_E7315_ = new_E7324_ | new_E7323_;
  assign new_E7316_ = new_E7326_ & new_E7325_;
  assign new_E7317_ = new_E7326_ & new_E7327_;
  assign new_E7318_ = new_E7319_ | new_E7328_;
  assign new_E7319_ = new_E7308_ | new_E7331_;
  assign new_E7320_ = new_E7330_ | new_E7329_;
  assign new_E7321_ = new_E7335_ & new_E7334_;
  assign new_E7322_ = new_E7333_ & new_E7332_;
  assign new_E7323_ = new_E7338_ | new_E7337_;
  assign new_E7324_ = new_E7333_ & new_E7336_;
  assign new_E7325_ = new_E7308_ | new_E7341_;
  assign new_E7326_ = new_E7340_ | new_E7339_;
  assign new_E7327_ = new_E7343_ | new_E7342_;
  assign new_E7328_ = ~new_E7319_ & new_E7345_;
  assign new_E7329_ = ~new_E7321_ & new_E7333_;
  assign new_E7330_ = new_E7321_ & ~new_E7333_;
  assign new_E7331_ = new_E7307_ & ~new_E7308_;
  assign new_E7332_ = ~new_E7354_ | ~new_E7355_;
  assign new_E7333_ = new_E7347_ | new_E7349_;
  assign new_E7334_ = new_E7357_ | new_E7356_;
  assign new_E7335_ = new_E7351_ | new_E7350_;
  assign new_E7336_ = ~new_E7359_ | ~new_E7358_;
  assign new_E7337_ = ~new_E7360_ & new_E7361_;
  assign new_E7338_ = new_E7360_ & ~new_E7361_;
  assign new_E7339_ = ~new_E7307_ & new_E7308_;
  assign new_E7340_ = new_E7307_ & ~new_E7308_;
  assign new_E7341_ = ~new_E7323_ | new_E7333_;
  assign new_E7342_ = new_E7323_ & new_E7333_;
  assign new_E7343_ = ~new_E7323_ & ~new_E7333_;
  assign new_E7344_ = new_E7365_ | new_E7364_;
  assign new_E7345_ = new_E7311_ | new_E7344_;
  assign new_E7346_ = new_E7369_ | new_E7368_;
  assign new_E7347_ = ~new_E7311_ & new_E7346_;
  assign new_E7348_ = new_E7367_ | new_E7366_;
  assign new_E7349_ = new_E7311_ & new_E7348_;
  assign new_E7350_ = new_E7309_ & ~new_E7319_;
  assign new_E7351_ = ~new_E7309_ & new_E7319_;
  assign new_E7352_ = ~new_E7308_ | ~new_E7333_;
  assign new_E7353_ = new_E7319_ & new_E7352_;
  assign new_E7354_ = ~new_E7319_ & ~new_E7353_;
  assign new_E7355_ = new_E7319_ | new_E7352_;
  assign new_E7356_ = ~new_E7309_ & new_E7310_;
  assign new_E7357_ = new_E7309_ & ~new_E7310_;
  assign new_E7358_ = new_E7326_ | new_E7363_;
  assign new_E7359_ = ~new_E7326_ & ~new_E7362_;
  assign new_E7360_ = new_E7309_ | new_E7326_;
  assign new_E7361_ = new_E7309_ | new_E7310_;
  assign new_E7362_ = new_E7326_ & new_E7363_;
  assign new_E7363_ = ~new_E7308_ | ~new_E7333_;
  assign new_E7364_ = new_E7341_ & new_E7361_;
  assign new_E7365_ = ~new_E7341_ & ~new_E7361_;
  assign new_E7366_ = new_E7370_ | new_E7371_;
  assign new_E7367_ = ~new_E7312_ & new_E7326_;
  assign new_E7368_ = new_E7372_ | new_E7373_;
  assign new_E7369_ = new_E7312_ & new_E7326_;
  assign new_E7370_ = ~new_E7312_ & ~new_E7326_;
  assign new_E7371_ = new_E7312_ & ~new_E7326_;
  assign new_E7372_ = new_E7312_ & ~new_E7326_;
  assign new_E7373_ = ~new_E7312_ & new_E7326_;
  assign new_E7374_ = new_F5894_;
  assign new_E7375_ = new_F5961_;
  assign new_E7376_ = new_F6028_;
  assign new_E7377_ = new_F6095_;
  assign new_E7378_ = new_F6162_;
  assign new_E7379_ = new_F6229_;
  assign new_E7380_ = new_E7387_ & new_E7386_;
  assign new_E7381_ = new_E7389_ | new_E7388_;
  assign new_E7382_ = new_E7391_ | new_E7390_;
  assign new_E7383_ = new_E7393_ & new_E7392_;
  assign new_E7384_ = new_E7393_ & new_E7394_;
  assign new_E7385_ = new_E7386_ | new_E7395_;
  assign new_E7386_ = new_E7375_ | new_E7398_;
  assign new_E7387_ = new_E7397_ | new_E7396_;
  assign new_E7388_ = new_E7402_ & new_E7401_;
  assign new_E7389_ = new_E7400_ & new_E7399_;
  assign new_E7390_ = new_E7405_ | new_E7404_;
  assign new_E7391_ = new_E7400_ & new_E7403_;
  assign new_E7392_ = new_E7375_ | new_E7408_;
  assign new_E7393_ = new_E7407_ | new_E7406_;
  assign new_E7394_ = new_E7410_ | new_E7409_;
  assign new_E7395_ = ~new_E7386_ & new_E7412_;
  assign new_E7396_ = ~new_E7388_ & new_E7400_;
  assign new_E7397_ = new_E7388_ & ~new_E7400_;
  assign new_E7398_ = new_E7374_ & ~new_E7375_;
  assign new_E7399_ = ~new_E7421_ | ~new_E7422_;
  assign new_E7400_ = new_E7414_ | new_E7416_;
  assign new_E7401_ = new_E7424_ | new_E7423_;
  assign new_E7402_ = new_E7418_ | new_E7417_;
  assign new_E7403_ = ~new_E7426_ | ~new_E7425_;
  assign new_E7404_ = ~new_E7427_ & new_E7428_;
  assign new_E7405_ = new_E7427_ & ~new_E7428_;
  assign new_E7406_ = ~new_E7374_ & new_E7375_;
  assign new_E7407_ = new_E7374_ & ~new_E7375_;
  assign new_E7408_ = ~new_E7390_ | new_E7400_;
  assign new_E7409_ = new_E7390_ & new_E7400_;
  assign new_E7410_ = ~new_E7390_ & ~new_E7400_;
  assign new_E7411_ = new_E7432_ | new_E7431_;
  assign new_E7412_ = new_E7378_ | new_E7411_;
  assign new_E7413_ = new_E7436_ | new_E7435_;
  assign new_E7414_ = ~new_E7378_ & new_E7413_;
  assign new_E7415_ = new_E7434_ | new_E7433_;
  assign new_E7416_ = new_E7378_ & new_E7415_;
  assign new_E7417_ = new_E7376_ & ~new_E7386_;
  assign new_E7418_ = ~new_E7376_ & new_E7386_;
  assign new_E7419_ = ~new_E7375_ | ~new_E7400_;
  assign new_E7420_ = new_E7386_ & new_E7419_;
  assign new_E7421_ = ~new_E7386_ & ~new_E7420_;
  assign new_E7422_ = new_E7386_ | new_E7419_;
  assign new_E7423_ = ~new_E7376_ & new_E7377_;
  assign new_E7424_ = new_E7376_ & ~new_E7377_;
  assign new_E7425_ = new_E7393_ | new_E7430_;
  assign new_E7426_ = ~new_E7393_ & ~new_E7429_;
  assign new_E7427_ = new_E7376_ | new_E7393_;
  assign new_E7428_ = new_E7376_ | new_E7377_;
  assign new_E7429_ = new_E7393_ & new_E7430_;
  assign new_E7430_ = ~new_E7375_ | ~new_E7400_;
  assign new_E7431_ = new_E7408_ & new_E7428_;
  assign new_E7432_ = ~new_E7408_ & ~new_E7428_;
  assign new_E7433_ = new_E7437_ | new_E7438_;
  assign new_E7434_ = ~new_E7379_ & new_E7393_;
  assign new_E7435_ = new_E7439_ | new_E7440_;
  assign new_E7436_ = new_E7379_ & new_E7393_;
  assign new_E7437_ = ~new_E7379_ & ~new_E7393_;
  assign new_E7438_ = new_E7379_ & ~new_E7393_;
  assign new_E7439_ = new_E7379_ & ~new_E7393_;
  assign new_E7440_ = ~new_E7379_ & new_E7393_;
  assign new_E7441_ = new_F6296_;
  assign new_E7442_ = new_F6363_;
  assign new_E7443_ = new_F6430_;
  assign new_E7444_ = new_F6497_;
  assign new_E7445_ = new_F6564_;
  assign new_E7446_ = new_F6631_;
  assign new_E7447_ = new_E7454_ & new_E7453_;
  assign new_E7448_ = new_E7456_ | new_E7455_;
  assign new_E7449_ = new_E7458_ | new_E7457_;
  assign new_E7450_ = new_E7460_ & new_E7459_;
  assign new_E7451_ = new_E7460_ & new_E7461_;
  assign new_E7452_ = new_E7453_ | new_E7462_;
  assign new_E7453_ = new_E7442_ | new_E7465_;
  assign new_E7454_ = new_E7464_ | new_E7463_;
  assign new_E7455_ = new_E7469_ & new_E7468_;
  assign new_E7456_ = new_E7467_ & new_E7466_;
  assign new_E7457_ = new_E7472_ | new_E7471_;
  assign new_E7458_ = new_E7467_ & new_E7470_;
  assign new_E7459_ = new_E7442_ | new_E7475_;
  assign new_E7460_ = new_E7474_ | new_E7473_;
  assign new_E7461_ = new_E7477_ | new_E7476_;
  assign new_E7462_ = ~new_E7453_ & new_E7479_;
  assign new_E7463_ = ~new_E7455_ & new_E7467_;
  assign new_E7464_ = new_E7455_ & ~new_E7467_;
  assign new_E7465_ = new_E7441_ & ~new_E7442_;
  assign new_E7466_ = ~new_E7488_ | ~new_E7489_;
  assign new_E7467_ = new_E7481_ | new_E7483_;
  assign new_E7468_ = new_E7491_ | new_E7490_;
  assign new_E7469_ = new_E7485_ | new_E7484_;
  assign new_E7470_ = ~new_E7493_ | ~new_E7492_;
  assign new_E7471_ = ~new_E7494_ & new_E7495_;
  assign new_E7472_ = new_E7494_ & ~new_E7495_;
  assign new_E7473_ = ~new_E7441_ & new_E7442_;
  assign new_E7474_ = new_E7441_ & ~new_E7442_;
  assign new_E7475_ = ~new_E7457_ | new_E7467_;
  assign new_E7476_ = new_E7457_ & new_E7467_;
  assign new_E7477_ = ~new_E7457_ & ~new_E7467_;
  assign new_E7478_ = new_E7499_ | new_E7498_;
  assign new_E7479_ = new_E7445_ | new_E7478_;
  assign new_E7480_ = new_E7503_ | new_E7502_;
  assign new_E7481_ = ~new_E7445_ & new_E7480_;
  assign new_E7482_ = new_E7501_ | new_E7500_;
  assign new_E7483_ = new_E7445_ & new_E7482_;
  assign new_E7484_ = new_E7443_ & ~new_E7453_;
  assign new_E7485_ = ~new_E7443_ & new_E7453_;
  assign new_E7486_ = ~new_E7442_ | ~new_E7467_;
  assign new_E7487_ = new_E7453_ & new_E7486_;
  assign new_E7488_ = ~new_E7453_ & ~new_E7487_;
  assign new_E7489_ = new_E7453_ | new_E7486_;
  assign new_E7490_ = ~new_E7443_ & new_E7444_;
  assign new_E7491_ = new_E7443_ & ~new_E7444_;
  assign new_E7492_ = new_E7460_ | new_E7497_;
  assign new_E7493_ = ~new_E7460_ & ~new_E7496_;
  assign new_E7494_ = new_E7443_ | new_E7460_;
  assign new_E7495_ = new_E7443_ | new_E7444_;
  assign new_E7496_ = new_E7460_ & new_E7497_;
  assign new_E7497_ = ~new_E7442_ | ~new_E7467_;
  assign new_E7498_ = new_E7475_ & new_E7495_;
  assign new_E7499_ = ~new_E7475_ & ~new_E7495_;
  assign new_E7500_ = new_E7504_ | new_E7505_;
  assign new_E7501_ = ~new_E7446_ & new_E7460_;
  assign new_E7502_ = new_E7506_ | new_E7507_;
  assign new_E7503_ = new_E7446_ & new_E7460_;
  assign new_E7504_ = ~new_E7446_ & ~new_E7460_;
  assign new_E7505_ = new_E7446_ & ~new_E7460_;
  assign new_E7506_ = new_E7446_ & ~new_E7460_;
  assign new_E7507_ = ~new_E7446_ & new_E7460_;
  assign new_E7508_ = new_F6698_;
  assign new_E7509_ = new_F6765_;
  assign new_E7510_ = new_F6832_;
  assign new_E7511_ = new_F6899_;
  assign new_E7512_ = new_F6966_;
  assign new_E7513_ = new_F7033_;
  assign new_E7514_ = new_E7521_ & new_E7520_;
  assign new_E7515_ = new_E7523_ | new_E7522_;
  assign new_E7516_ = new_E7525_ | new_E7524_;
  assign new_E7517_ = new_E7527_ & new_E7526_;
  assign new_E7518_ = new_E7527_ & new_E7528_;
  assign new_E7519_ = new_E7520_ | new_E7529_;
  assign new_E7520_ = new_E7509_ | new_E7532_;
  assign new_E7521_ = new_E7531_ | new_E7530_;
  assign new_E7522_ = new_E7536_ & new_E7535_;
  assign new_E7523_ = new_E7534_ & new_E7533_;
  assign new_E7524_ = new_E7539_ | new_E7538_;
  assign new_E7525_ = new_E7534_ & new_E7537_;
  assign new_E7526_ = new_E7509_ | new_E7542_;
  assign new_E7527_ = new_E7541_ | new_E7540_;
  assign new_E7528_ = new_E7544_ | new_E7543_;
  assign new_E7529_ = ~new_E7520_ & new_E7546_;
  assign new_E7530_ = ~new_E7522_ & new_E7534_;
  assign new_E7531_ = new_E7522_ & ~new_E7534_;
  assign new_E7532_ = new_E7508_ & ~new_E7509_;
  assign new_E7533_ = ~new_E7555_ | ~new_E7556_;
  assign new_E7534_ = new_E7548_ | new_E7550_;
  assign new_E7535_ = new_E7558_ | new_E7557_;
  assign new_E7536_ = new_E7552_ | new_E7551_;
  assign new_E7537_ = ~new_E7560_ | ~new_E7559_;
  assign new_E7538_ = ~new_E7561_ & new_E7562_;
  assign new_E7539_ = new_E7561_ & ~new_E7562_;
  assign new_E7540_ = ~new_E7508_ & new_E7509_;
  assign new_E7541_ = new_E7508_ & ~new_E7509_;
  assign new_E7542_ = ~new_E7524_ | new_E7534_;
  assign new_E7543_ = new_E7524_ & new_E7534_;
  assign new_E7544_ = ~new_E7524_ & ~new_E7534_;
  assign new_E7545_ = new_E7566_ | new_E7565_;
  assign new_E7546_ = new_E7512_ | new_E7545_;
  assign new_E7547_ = new_E7570_ | new_E7569_;
  assign new_E7548_ = ~new_E7512_ & new_E7547_;
  assign new_E7549_ = new_E7568_ | new_E7567_;
  assign new_E7550_ = new_E7512_ & new_E7549_;
  assign new_E7551_ = new_E7510_ & ~new_E7520_;
  assign new_E7552_ = ~new_E7510_ & new_E7520_;
  assign new_E7553_ = ~new_E7509_ | ~new_E7534_;
  assign new_E7554_ = new_E7520_ & new_E7553_;
  assign new_E7555_ = ~new_E7520_ & ~new_E7554_;
  assign new_E7556_ = new_E7520_ | new_E7553_;
  assign new_E7557_ = ~new_E7510_ & new_E7511_;
  assign new_E7558_ = new_E7510_ & ~new_E7511_;
  assign new_E7559_ = new_E7527_ | new_E7564_;
  assign new_E7560_ = ~new_E7527_ & ~new_E7563_;
  assign new_E7561_ = new_E7510_ | new_E7527_;
  assign new_E7562_ = new_E7510_ | new_E7511_;
  assign new_E7563_ = new_E7527_ & new_E7564_;
  assign new_E7564_ = ~new_E7509_ | ~new_E7534_;
  assign new_E7565_ = new_E7542_ & new_E7562_;
  assign new_E7566_ = ~new_E7542_ & ~new_E7562_;
  assign new_E7567_ = new_E7571_ | new_E7572_;
  assign new_E7568_ = ~new_E7513_ & new_E7527_;
  assign new_E7569_ = new_E7573_ | new_E7574_;
  assign new_E7570_ = new_E7513_ & new_E7527_;
  assign new_E7571_ = ~new_E7513_ & ~new_E7527_;
  assign new_E7572_ = new_E7513_ & ~new_E7527_;
  assign new_E7573_ = new_E7513_ & ~new_E7527_;
  assign new_E7574_ = ~new_E7513_ & new_E7527_;
  assign new_E7575_ = new_F7100_;
  assign new_E7576_ = new_F7167_;
  assign new_E7577_ = new_F7234_;
  assign new_E7578_ = new_F7301_;
  assign new_E7579_ = new_F7368_;
  assign new_E7580_ = new_F7435_;
  assign new_E7581_ = new_E7588_ & new_E7587_;
  assign new_E7582_ = new_E7590_ | new_E7589_;
  assign new_E7583_ = new_E7592_ | new_E7591_;
  assign new_E7584_ = new_E7594_ & new_E7593_;
  assign new_E7585_ = new_E7594_ & new_E7595_;
  assign new_E7586_ = new_E7587_ | new_E7596_;
  assign new_E7587_ = new_E7576_ | new_E7599_;
  assign new_E7588_ = new_E7598_ | new_E7597_;
  assign new_E7589_ = new_E7603_ & new_E7602_;
  assign new_E7590_ = new_E7601_ & new_E7600_;
  assign new_E7591_ = new_E7606_ | new_E7605_;
  assign new_E7592_ = new_E7601_ & new_E7604_;
  assign new_E7593_ = new_E7576_ | new_E7609_;
  assign new_E7594_ = new_E7608_ | new_E7607_;
  assign new_E7595_ = new_E7611_ | new_E7610_;
  assign new_E7596_ = ~new_E7587_ & new_E7613_;
  assign new_E7597_ = ~new_E7589_ & new_E7601_;
  assign new_E7598_ = new_E7589_ & ~new_E7601_;
  assign new_E7599_ = new_E7575_ & ~new_E7576_;
  assign new_E7600_ = ~new_E7622_ | ~new_E7623_;
  assign new_E7601_ = new_E7615_ | new_E7617_;
  assign new_E7602_ = new_E7625_ | new_E7624_;
  assign new_E7603_ = new_E7619_ | new_E7618_;
  assign new_E7604_ = ~new_E7627_ | ~new_E7626_;
  assign new_E7605_ = ~new_E7628_ & new_E7629_;
  assign new_E7606_ = new_E7628_ & ~new_E7629_;
  assign new_E7607_ = ~new_E7575_ & new_E7576_;
  assign new_E7608_ = new_E7575_ & ~new_E7576_;
  assign new_E7609_ = ~new_E7591_ | new_E7601_;
  assign new_E7610_ = new_E7591_ & new_E7601_;
  assign new_E7611_ = ~new_E7591_ & ~new_E7601_;
  assign new_E7612_ = new_E7633_ | new_E7632_;
  assign new_E7613_ = new_E7579_ | new_E7612_;
  assign new_E7614_ = new_E7637_ | new_E7636_;
  assign new_E7615_ = ~new_E7579_ & new_E7614_;
  assign new_E7616_ = new_E7635_ | new_E7634_;
  assign new_E7617_ = new_E7579_ & new_E7616_;
  assign new_E7618_ = new_E7577_ & ~new_E7587_;
  assign new_E7619_ = ~new_E7577_ & new_E7587_;
  assign new_E7620_ = ~new_E7576_ | ~new_E7601_;
  assign new_E7621_ = new_E7587_ & new_E7620_;
  assign new_E7622_ = ~new_E7587_ & ~new_E7621_;
  assign new_E7623_ = new_E7587_ | new_E7620_;
  assign new_E7624_ = ~new_E7577_ & new_E7578_;
  assign new_E7625_ = new_E7577_ & ~new_E7578_;
  assign new_E7626_ = new_E7594_ | new_E7631_;
  assign new_E7627_ = ~new_E7594_ & ~new_E7630_;
  assign new_E7628_ = new_E7577_ | new_E7594_;
  assign new_E7629_ = new_E7577_ | new_E7578_;
  assign new_E7630_ = new_E7594_ & new_E7631_;
  assign new_E7631_ = ~new_E7576_ | ~new_E7601_;
  assign new_E7632_ = new_E7609_ & new_E7629_;
  assign new_E7633_ = ~new_E7609_ & ~new_E7629_;
  assign new_E7634_ = new_E7638_ | new_E7639_;
  assign new_E7635_ = ~new_E7580_ & new_E7594_;
  assign new_E7636_ = new_E7640_ | new_E7641_;
  assign new_E7637_ = new_E7580_ & new_E7594_;
  assign new_E7638_ = ~new_E7580_ & ~new_E7594_;
  assign new_E7639_ = new_E7580_ & ~new_E7594_;
  assign new_E7640_ = new_E7580_ & ~new_E7594_;
  assign new_E7641_ = ~new_E7580_ & new_E7594_;
  assign new_E7642_ = new_F7502_;
  assign new_E7643_ = new_F7569_;
  assign new_E7644_ = new_F7636_;
  assign new_E7645_ = new_F7703_;
  assign new_E7646_ = new_F7770_;
  assign new_E7647_ = new_F7837_;
  assign new_E7648_ = new_E7655_ & new_E7654_;
  assign new_E7649_ = new_E7657_ | new_E7656_;
  assign new_E7650_ = new_E7659_ | new_E7658_;
  assign new_E7651_ = new_E7661_ & new_E7660_;
  assign new_E7652_ = new_E7661_ & new_E7662_;
  assign new_E7653_ = new_E7654_ | new_E7663_;
  assign new_E7654_ = new_E7643_ | new_E7666_;
  assign new_E7655_ = new_E7665_ | new_E7664_;
  assign new_E7656_ = new_E7670_ & new_E7669_;
  assign new_E7657_ = new_E7668_ & new_E7667_;
  assign new_E7658_ = new_E7673_ | new_E7672_;
  assign new_E7659_ = new_E7668_ & new_E7671_;
  assign new_E7660_ = new_E7643_ | new_E7676_;
  assign new_E7661_ = new_E7675_ | new_E7674_;
  assign new_E7662_ = new_E7678_ | new_E7677_;
  assign new_E7663_ = ~new_E7654_ & new_E7680_;
  assign new_E7664_ = ~new_E7656_ & new_E7668_;
  assign new_E7665_ = new_E7656_ & ~new_E7668_;
  assign new_E7666_ = new_E7642_ & ~new_E7643_;
  assign new_E7667_ = ~new_E7689_ | ~new_E7690_;
  assign new_E7668_ = new_E7682_ | new_E7684_;
  assign new_E7669_ = new_E7692_ | new_E7691_;
  assign new_E7670_ = new_E7686_ | new_E7685_;
  assign new_E7671_ = ~new_E7694_ | ~new_E7693_;
  assign new_E7672_ = ~new_E7695_ & new_E7696_;
  assign new_E7673_ = new_E7695_ & ~new_E7696_;
  assign new_E7674_ = ~new_E7642_ & new_E7643_;
  assign new_E7675_ = new_E7642_ & ~new_E7643_;
  assign new_E7676_ = ~new_E7658_ | new_E7668_;
  assign new_E7677_ = new_E7658_ & new_E7668_;
  assign new_E7678_ = ~new_E7658_ & ~new_E7668_;
  assign new_E7679_ = new_E7700_ | new_E7699_;
  assign new_E7680_ = new_E7646_ | new_E7679_;
  assign new_E7681_ = new_E7704_ | new_E7703_;
  assign new_E7682_ = ~new_E7646_ & new_E7681_;
  assign new_E7683_ = new_E7702_ | new_E7701_;
  assign new_E7684_ = new_E7646_ & new_E7683_;
  assign new_E7685_ = new_E7644_ & ~new_E7654_;
  assign new_E7686_ = ~new_E7644_ & new_E7654_;
  assign new_E7687_ = ~new_E7643_ | ~new_E7668_;
  assign new_E7688_ = new_E7654_ & new_E7687_;
  assign new_E7689_ = ~new_E7654_ & ~new_E7688_;
  assign new_E7690_ = new_E7654_ | new_E7687_;
  assign new_E7691_ = ~new_E7644_ & new_E7645_;
  assign new_E7692_ = new_E7644_ & ~new_E7645_;
  assign new_E7693_ = new_E7661_ | new_E7698_;
  assign new_E7694_ = ~new_E7661_ & ~new_E7697_;
  assign new_E7695_ = new_E7644_ | new_E7661_;
  assign new_E7696_ = new_E7644_ | new_E7645_;
  assign new_E7697_ = new_E7661_ & new_E7698_;
  assign new_E7698_ = ~new_E7643_ | ~new_E7668_;
  assign new_E7699_ = new_E7676_ & new_E7696_;
  assign new_E7700_ = ~new_E7676_ & ~new_E7696_;
  assign new_E7701_ = new_E7705_ | new_E7706_;
  assign new_E7702_ = ~new_E7647_ & new_E7661_;
  assign new_E7703_ = new_E7707_ | new_E7708_;
  assign new_E7704_ = new_E7647_ & new_E7661_;
  assign new_E7705_ = ~new_E7647_ & ~new_E7661_;
  assign new_E7706_ = new_E7647_ & ~new_E7661_;
  assign new_E7707_ = new_E7647_ & ~new_E7661_;
  assign new_E7708_ = ~new_E7647_ & new_E7661_;
  assign new_E7709_ = new_F7904_;
  assign new_E7710_ = new_F7971_;
  assign new_E7711_ = new_F8038_;
  assign new_E7712_ = new_F8105_;
  assign new_E7713_ = new_F8172_;
  assign new_E7714_ = new_F8239_;
  assign new_E7715_ = new_E7722_ & new_E7721_;
  assign new_E7716_ = new_E7724_ | new_E7723_;
  assign new_E7717_ = new_E7726_ | new_E7725_;
  assign new_E7718_ = new_E7728_ & new_E7727_;
  assign new_E7719_ = new_E7728_ & new_E7729_;
  assign new_E7720_ = new_E7721_ | new_E7730_;
  assign new_E7721_ = new_E7710_ | new_E7733_;
  assign new_E7722_ = new_E7732_ | new_E7731_;
  assign new_E7723_ = new_E7737_ & new_E7736_;
  assign new_E7724_ = new_E7735_ & new_E7734_;
  assign new_E7725_ = new_E7740_ | new_E7739_;
  assign new_E7726_ = new_E7735_ & new_E7738_;
  assign new_E7727_ = new_E7710_ | new_E7743_;
  assign new_E7728_ = new_E7742_ | new_E7741_;
  assign new_E7729_ = new_E7745_ | new_E7744_;
  assign new_E7730_ = ~new_E7721_ & new_E7747_;
  assign new_E7731_ = ~new_E7723_ & new_E7735_;
  assign new_E7732_ = new_E7723_ & ~new_E7735_;
  assign new_E7733_ = new_E7709_ & ~new_E7710_;
  assign new_E7734_ = ~new_E7756_ | ~new_E7757_;
  assign new_E7735_ = new_E7749_ | new_E7751_;
  assign new_E7736_ = new_E7759_ | new_E7758_;
  assign new_E7737_ = new_E7753_ | new_E7752_;
  assign new_E7738_ = ~new_E7761_ | ~new_E7760_;
  assign new_E7739_ = ~new_E7762_ & new_E7763_;
  assign new_E7740_ = new_E7762_ & ~new_E7763_;
  assign new_E7741_ = ~new_E7709_ & new_E7710_;
  assign new_E7742_ = new_E7709_ & ~new_E7710_;
  assign new_E7743_ = ~new_E7725_ | new_E7735_;
  assign new_E7744_ = new_E7725_ & new_E7735_;
  assign new_E7745_ = ~new_E7725_ & ~new_E7735_;
  assign new_E7746_ = new_E7767_ | new_E7766_;
  assign new_E7747_ = new_E7713_ | new_E7746_;
  assign new_E7748_ = new_E7771_ | new_E7770_;
  assign new_E7749_ = ~new_E7713_ & new_E7748_;
  assign new_E7750_ = new_E7769_ | new_E7768_;
  assign new_E7751_ = new_E7713_ & new_E7750_;
  assign new_E7752_ = new_E7711_ & ~new_E7721_;
  assign new_E7753_ = ~new_E7711_ & new_E7721_;
  assign new_E7754_ = ~new_E7710_ | ~new_E7735_;
  assign new_E7755_ = new_E7721_ & new_E7754_;
  assign new_E7756_ = ~new_E7721_ & ~new_E7755_;
  assign new_E7757_ = new_E7721_ | new_E7754_;
  assign new_E7758_ = ~new_E7711_ & new_E7712_;
  assign new_E7759_ = new_E7711_ & ~new_E7712_;
  assign new_E7760_ = new_E7728_ | new_E7765_;
  assign new_E7761_ = ~new_E7728_ & ~new_E7764_;
  assign new_E7762_ = new_E7711_ | new_E7728_;
  assign new_E7763_ = new_E7711_ | new_E7712_;
  assign new_E7764_ = new_E7728_ & new_E7765_;
  assign new_E7765_ = ~new_E7710_ | ~new_E7735_;
  assign new_E7766_ = new_E7743_ & new_E7763_;
  assign new_E7767_ = ~new_E7743_ & ~new_E7763_;
  assign new_E7768_ = new_E7772_ | new_E7773_;
  assign new_E7769_ = ~new_E7714_ & new_E7728_;
  assign new_E7770_ = new_E7774_ | new_E7775_;
  assign new_E7771_ = new_E7714_ & new_E7728_;
  assign new_E7772_ = ~new_E7714_ & ~new_E7728_;
  assign new_E7773_ = new_E7714_ & ~new_E7728_;
  assign new_E7774_ = new_E7714_ & ~new_E7728_;
  assign new_E7775_ = ~new_E7714_ & new_E7728_;
  assign new_E7776_ = new_F8306_;
  assign new_E7777_ = new_F8373_;
  assign new_E7778_ = new_F8440_;
  assign new_E7779_ = new_F8507_;
  assign new_E7780_ = new_F8574_;
  assign new_E7781_ = new_F8641_;
  assign new_E7782_ = new_E7789_ & new_E7788_;
  assign new_E7783_ = new_E7791_ | new_E7790_;
  assign new_E7784_ = new_E7793_ | new_E7792_;
  assign new_E7785_ = new_E7795_ & new_E7794_;
  assign new_E7786_ = new_E7795_ & new_E7796_;
  assign new_E7787_ = new_E7788_ | new_E7797_;
  assign new_E7788_ = new_E7777_ | new_E7800_;
  assign new_E7789_ = new_E7799_ | new_E7798_;
  assign new_E7790_ = new_E7804_ & new_E7803_;
  assign new_E7791_ = new_E7802_ & new_E7801_;
  assign new_E7792_ = new_E7807_ | new_E7806_;
  assign new_E7793_ = new_E7802_ & new_E7805_;
  assign new_E7794_ = new_E7777_ | new_E7810_;
  assign new_E7795_ = new_E7809_ | new_E7808_;
  assign new_E7796_ = new_E7812_ | new_E7811_;
  assign new_E7797_ = ~new_E7788_ & new_E7814_;
  assign new_E7798_ = ~new_E7790_ & new_E7802_;
  assign new_E7799_ = new_E7790_ & ~new_E7802_;
  assign new_E7800_ = new_E7776_ & ~new_E7777_;
  assign new_E7801_ = ~new_E7823_ | ~new_E7824_;
  assign new_E7802_ = new_E7816_ | new_E7818_;
  assign new_E7803_ = new_E7826_ | new_E7825_;
  assign new_E7804_ = new_E7820_ | new_E7819_;
  assign new_E7805_ = ~new_E7828_ | ~new_E7827_;
  assign new_E7806_ = ~new_E7829_ & new_E7830_;
  assign new_E7807_ = new_E7829_ & ~new_E7830_;
  assign new_E7808_ = ~new_E7776_ & new_E7777_;
  assign new_E7809_ = new_E7776_ & ~new_E7777_;
  assign new_E7810_ = ~new_E7792_ | new_E7802_;
  assign new_E7811_ = new_E7792_ & new_E7802_;
  assign new_E7812_ = ~new_E7792_ & ~new_E7802_;
  assign new_E7813_ = new_E7834_ | new_E7833_;
  assign new_E7814_ = new_E7780_ | new_E7813_;
  assign new_E7815_ = new_E7838_ | new_E7837_;
  assign new_E7816_ = ~new_E7780_ & new_E7815_;
  assign new_E7817_ = new_E7836_ | new_E7835_;
  assign new_E7818_ = new_E7780_ & new_E7817_;
  assign new_E7819_ = new_E7778_ & ~new_E7788_;
  assign new_E7820_ = ~new_E7778_ & new_E7788_;
  assign new_E7821_ = ~new_E7777_ | ~new_E7802_;
  assign new_E7822_ = new_E7788_ & new_E7821_;
  assign new_E7823_ = ~new_E7788_ & ~new_E7822_;
  assign new_E7824_ = new_E7788_ | new_E7821_;
  assign new_E7825_ = ~new_E7778_ & new_E7779_;
  assign new_E7826_ = new_E7778_ & ~new_E7779_;
  assign new_E7827_ = new_E7795_ | new_E7832_;
  assign new_E7828_ = ~new_E7795_ & ~new_E7831_;
  assign new_E7829_ = new_E7778_ | new_E7795_;
  assign new_E7830_ = new_E7778_ | new_E7779_;
  assign new_E7831_ = new_E7795_ & new_E7832_;
  assign new_E7832_ = ~new_E7777_ | ~new_E7802_;
  assign new_E7833_ = new_E7810_ & new_E7830_;
  assign new_E7834_ = ~new_E7810_ & ~new_E7830_;
  assign new_E7835_ = new_E7839_ | new_E7840_;
  assign new_E7836_ = ~new_E7781_ & new_E7795_;
  assign new_E7837_ = new_E7841_ | new_E7842_;
  assign new_E7838_ = new_E7781_ & new_E7795_;
  assign new_E7839_ = ~new_E7781_ & ~new_E7795_;
  assign new_E7840_ = new_E7781_ & ~new_E7795_;
  assign new_E7841_ = new_E7781_ & ~new_E7795_;
  assign new_E7842_ = ~new_E7781_ & new_E7795_;
  assign new_E7843_ = new_F8708_;
  assign new_E7844_ = new_F8775_;
  assign new_E7845_ = new_F8842_;
  assign new_E7846_ = new_F8909_;
  assign new_E7847_ = new_F8976_;
  assign new_E7848_ = new_F9043_;
  assign new_E7849_ = new_E7856_ & new_E7855_;
  assign new_E7850_ = new_E7858_ | new_E7857_;
  assign new_E7851_ = new_E7860_ | new_E7859_;
  assign new_E7852_ = new_E7862_ & new_E7861_;
  assign new_E7853_ = new_E7862_ & new_E7863_;
  assign new_E7854_ = new_E7855_ | new_E7864_;
  assign new_E7855_ = new_E7844_ | new_E7867_;
  assign new_E7856_ = new_E7866_ | new_E7865_;
  assign new_E7857_ = new_E7871_ & new_E7870_;
  assign new_E7858_ = new_E7869_ & new_E7868_;
  assign new_E7859_ = new_E7874_ | new_E7873_;
  assign new_E7860_ = new_E7869_ & new_E7872_;
  assign new_E7861_ = new_E7844_ | new_E7877_;
  assign new_E7862_ = new_E7876_ | new_E7875_;
  assign new_E7863_ = new_E7879_ | new_E7878_;
  assign new_E7864_ = ~new_E7855_ & new_E7881_;
  assign new_E7865_ = ~new_E7857_ & new_E7869_;
  assign new_E7866_ = new_E7857_ & ~new_E7869_;
  assign new_E7867_ = new_E7843_ & ~new_E7844_;
  assign new_E7868_ = ~new_E7890_ | ~new_E7891_;
  assign new_E7869_ = new_E7883_ | new_E7885_;
  assign new_E7870_ = new_E7893_ | new_E7892_;
  assign new_E7871_ = new_E7887_ | new_E7886_;
  assign new_E7872_ = ~new_E7895_ | ~new_E7894_;
  assign new_E7873_ = ~new_E7896_ & new_E7897_;
  assign new_E7874_ = new_E7896_ & ~new_E7897_;
  assign new_E7875_ = ~new_E7843_ & new_E7844_;
  assign new_E7876_ = new_E7843_ & ~new_E7844_;
  assign new_E7877_ = ~new_E7859_ | new_E7869_;
  assign new_E7878_ = new_E7859_ & new_E7869_;
  assign new_E7879_ = ~new_E7859_ & ~new_E7869_;
  assign new_E7880_ = new_E7901_ | new_E7900_;
  assign new_E7881_ = new_E7847_ | new_E7880_;
  assign new_E7882_ = new_E7905_ | new_E7904_;
  assign new_E7883_ = ~new_E7847_ & new_E7882_;
  assign new_E7884_ = new_E7903_ | new_E7902_;
  assign new_E7885_ = new_E7847_ & new_E7884_;
  assign new_E7886_ = new_E7845_ & ~new_E7855_;
  assign new_E7887_ = ~new_E7845_ & new_E7855_;
  assign new_E7888_ = ~new_E7844_ | ~new_E7869_;
  assign new_E7889_ = new_E7855_ & new_E7888_;
  assign new_E7890_ = ~new_E7855_ & ~new_E7889_;
  assign new_E7891_ = new_E7855_ | new_E7888_;
  assign new_E7892_ = ~new_E7845_ & new_E7846_;
  assign new_E7893_ = new_E7845_ & ~new_E7846_;
  assign new_E7894_ = new_E7862_ | new_E7899_;
  assign new_E7895_ = ~new_E7862_ & ~new_E7898_;
  assign new_E7896_ = new_E7845_ | new_E7862_;
  assign new_E7897_ = new_E7845_ | new_E7846_;
  assign new_E7898_ = new_E7862_ & new_E7899_;
  assign new_E7899_ = ~new_E7844_ | ~new_E7869_;
  assign new_E7900_ = new_E7877_ & new_E7897_;
  assign new_E7901_ = ~new_E7877_ & ~new_E7897_;
  assign new_E7902_ = new_E7906_ | new_E7907_;
  assign new_E7903_ = ~new_E7848_ & new_E7862_;
  assign new_E7904_ = new_E7908_ | new_E7909_;
  assign new_E7905_ = new_E7848_ & new_E7862_;
  assign new_E7906_ = ~new_E7848_ & ~new_E7862_;
  assign new_E7907_ = new_E7848_ & ~new_E7862_;
  assign new_E7908_ = new_E7848_ & ~new_E7862_;
  assign new_E7909_ = ~new_E7848_ & new_E7862_;
  assign new_E7910_ = new_F9110_;
  assign new_E7911_ = new_F9177_;
  assign new_E7912_ = new_F9244_;
  assign new_E7913_ = new_F9311_;
  assign new_E7914_ = new_F9378_;
  assign new_E7915_ = new_F9445_;
  assign new_E7916_ = new_E7923_ & new_E7922_;
  assign new_E7917_ = new_E7925_ | new_E7924_;
  assign new_E7918_ = new_E7927_ | new_E7926_;
  assign new_E7919_ = new_E7929_ & new_E7928_;
  assign new_E7920_ = new_E7929_ & new_E7930_;
  assign new_E7921_ = new_E7922_ | new_E7931_;
  assign new_E7922_ = new_E7911_ | new_E7934_;
  assign new_E7923_ = new_E7933_ | new_E7932_;
  assign new_E7924_ = new_E7938_ & new_E7937_;
  assign new_E7925_ = new_E7936_ & new_E7935_;
  assign new_E7926_ = new_E7941_ | new_E7940_;
  assign new_E7927_ = new_E7936_ & new_E7939_;
  assign new_E7928_ = new_E7911_ | new_E7944_;
  assign new_E7929_ = new_E7943_ | new_E7942_;
  assign new_E7930_ = new_E7946_ | new_E7945_;
  assign new_E7931_ = ~new_E7922_ & new_E7948_;
  assign new_E7932_ = ~new_E7924_ & new_E7936_;
  assign new_E7933_ = new_E7924_ & ~new_E7936_;
  assign new_E7934_ = new_E7910_ & ~new_E7911_;
  assign new_E7935_ = ~new_E7957_ | ~new_E7958_;
  assign new_E7936_ = new_E7950_ | new_E7952_;
  assign new_E7937_ = new_E7960_ | new_E7959_;
  assign new_E7938_ = new_E7954_ | new_E7953_;
  assign new_E7939_ = ~new_E7962_ | ~new_E7961_;
  assign new_E7940_ = ~new_E7963_ & new_E7964_;
  assign new_E7941_ = new_E7963_ & ~new_E7964_;
  assign new_E7942_ = ~new_E7910_ & new_E7911_;
  assign new_E7943_ = new_E7910_ & ~new_E7911_;
  assign new_E7944_ = ~new_E7926_ | new_E7936_;
  assign new_E7945_ = new_E7926_ & new_E7936_;
  assign new_E7946_ = ~new_E7926_ & ~new_E7936_;
  assign new_E7947_ = new_E7968_ | new_E7967_;
  assign new_E7948_ = new_E7914_ | new_E7947_;
  assign new_E7949_ = new_E7972_ | new_E7971_;
  assign new_E7950_ = ~new_E7914_ & new_E7949_;
  assign new_E7951_ = new_E7970_ | new_E7969_;
  assign new_E7952_ = new_E7914_ & new_E7951_;
  assign new_E7953_ = new_E7912_ & ~new_E7922_;
  assign new_E7954_ = ~new_E7912_ & new_E7922_;
  assign new_E7955_ = ~new_E7911_ | ~new_E7936_;
  assign new_E7956_ = new_E7922_ & new_E7955_;
  assign new_E7957_ = ~new_E7922_ & ~new_E7956_;
  assign new_E7958_ = new_E7922_ | new_E7955_;
  assign new_E7959_ = ~new_E7912_ & new_E7913_;
  assign new_E7960_ = new_E7912_ & ~new_E7913_;
  assign new_E7961_ = new_E7929_ | new_E7966_;
  assign new_E7962_ = ~new_E7929_ & ~new_E7965_;
  assign new_E7963_ = new_E7912_ | new_E7929_;
  assign new_E7964_ = new_E7912_ | new_E7913_;
  assign new_E7965_ = new_E7929_ & new_E7966_;
  assign new_E7966_ = ~new_E7911_ | ~new_E7936_;
  assign new_E7967_ = new_E7944_ & new_E7964_;
  assign new_E7968_ = ~new_E7944_ & ~new_E7964_;
  assign new_E7969_ = new_E7973_ | new_E7974_;
  assign new_E7970_ = ~new_E7915_ & new_E7929_;
  assign new_E7971_ = new_E7975_ | new_E7976_;
  assign new_E7972_ = new_E7915_ & new_E7929_;
  assign new_E7973_ = ~new_E7915_ & ~new_E7929_;
  assign new_E7974_ = new_E7915_ & ~new_E7929_;
  assign new_E7975_ = new_E7915_ & ~new_E7929_;
  assign new_E7976_ = ~new_E7915_ & new_E7929_;
  assign new_E7977_ = new_F9512_;
  assign new_E7978_ = new_F9579_;
  assign new_E7979_ = new_F9646_;
  assign new_E7980_ = new_F9713_;
  assign new_E7981_ = new_F9780_;
  assign new_E7982_ = new_F9847_;
  assign new_E7983_ = new_E7990_ & new_E7989_;
  assign new_E7984_ = new_E7992_ | new_E7991_;
  assign new_E7985_ = new_E7994_ | new_E7993_;
  assign new_E7986_ = new_E7996_ & new_E7995_;
  assign new_E7987_ = new_E7996_ & new_E7997_;
  assign new_E7988_ = new_E7989_ | new_E7998_;
  assign new_E7989_ = new_E7978_ | new_E8001_;
  assign new_E7990_ = new_E8000_ | new_E7999_;
  assign new_E7991_ = new_E8005_ & new_E8004_;
  assign new_E7992_ = new_E8003_ & new_E8002_;
  assign new_E7993_ = new_E8008_ | new_E8007_;
  assign new_E7994_ = new_E8003_ & new_E8006_;
  assign new_E7995_ = new_E7978_ | new_E8011_;
  assign new_E7996_ = new_E8010_ | new_E8009_;
  assign new_E7997_ = new_E8013_ | new_E8012_;
  assign new_E7998_ = ~new_E7989_ & new_E8015_;
  assign new_E7999_ = ~new_E7991_ & new_E8003_;
  assign new_E8000_ = new_E7991_ & ~new_E8003_;
  assign new_E8001_ = new_E7977_ & ~new_E7978_;
  assign new_E8002_ = ~new_E8024_ | ~new_E8025_;
  assign new_E8003_ = new_E8017_ | new_E8019_;
  assign new_E8004_ = new_E8027_ | new_E8026_;
  assign new_E8005_ = new_E8021_ | new_E8020_;
  assign new_E8006_ = ~new_E8029_ | ~new_E8028_;
  assign new_E8007_ = ~new_E8030_ & new_E8031_;
  assign new_E8008_ = new_E8030_ & ~new_E8031_;
  assign new_E8009_ = ~new_E7977_ & new_E7978_;
  assign new_E8010_ = new_E7977_ & ~new_E7978_;
  assign new_E8011_ = ~new_E7993_ | new_E8003_;
  assign new_E8012_ = new_E7993_ & new_E8003_;
  assign new_E8013_ = ~new_E7993_ & ~new_E8003_;
  assign new_E8014_ = new_E8035_ | new_E8034_;
  assign new_E8015_ = new_E7981_ | new_E8014_;
  assign new_E8016_ = new_E8039_ | new_E8038_;
  assign new_E8017_ = ~new_E7981_ & new_E8016_;
  assign new_E8018_ = new_E8037_ | new_E8036_;
  assign new_E8019_ = new_E7981_ & new_E8018_;
  assign new_E8020_ = new_E7979_ & ~new_E7989_;
  assign new_E8021_ = ~new_E7979_ & new_E7989_;
  assign new_E8022_ = ~new_E7978_ | ~new_E8003_;
  assign new_E8023_ = new_E7989_ & new_E8022_;
  assign new_E8024_ = ~new_E7989_ & ~new_E8023_;
  assign new_E8025_ = new_E7989_ | new_E8022_;
  assign new_E8026_ = ~new_E7979_ & new_E7980_;
  assign new_E8027_ = new_E7979_ & ~new_E7980_;
  assign new_E8028_ = new_E7996_ | new_E8033_;
  assign new_E8029_ = ~new_E7996_ & ~new_E8032_;
  assign new_E8030_ = new_E7979_ | new_E7996_;
  assign new_E8031_ = new_E7979_ | new_E7980_;
  assign new_E8032_ = new_E7996_ & new_E8033_;
  assign new_E8033_ = ~new_E7978_ | ~new_E8003_;
  assign new_E8034_ = new_E8011_ & new_E8031_;
  assign new_E8035_ = ~new_E8011_ & ~new_E8031_;
  assign new_E8036_ = new_E8040_ | new_E8041_;
  assign new_E8037_ = ~new_E7982_ & new_E7996_;
  assign new_E8038_ = new_E8042_ | new_E8043_;
  assign new_E8039_ = new_E7982_ & new_E7996_;
  assign new_E8040_ = ~new_E7982_ & ~new_E7996_;
  assign new_E8041_ = new_E7982_ & ~new_E7996_;
  assign new_E8042_ = new_E7982_ & ~new_E7996_;
  assign new_E8043_ = ~new_E7982_ & new_E7996_;
  assign new_E8044_ = new_F9914_;
  assign new_E8045_ = new_F9981_;
  assign new_E8046_ = new_G49_;
  assign new_E8047_ = new_G116_;
  assign new_E8048_ = new_G183_;
  assign new_E8049_ = new_G250_;
  assign new_E8050_ = new_E8057_ & new_E8056_;
  assign new_E8051_ = new_E8059_ | new_E8058_;
  assign new_E8052_ = new_E8061_ | new_E8060_;
  assign new_E8053_ = new_E8063_ & new_E8062_;
  assign new_E8054_ = new_E8063_ & new_E8064_;
  assign new_E8055_ = new_E8056_ | new_E8065_;
  assign new_E8056_ = new_E8045_ | new_E8068_;
  assign new_E8057_ = new_E8067_ | new_E8066_;
  assign new_E8058_ = new_E8072_ & new_E8071_;
  assign new_E8059_ = new_E8070_ & new_E8069_;
  assign new_E8060_ = new_E8075_ | new_E8074_;
  assign new_E8061_ = new_E8070_ & new_E8073_;
  assign new_E8062_ = new_E8045_ | new_E8078_;
  assign new_E8063_ = new_E8077_ | new_E8076_;
  assign new_E8064_ = new_E8080_ | new_E8079_;
  assign new_E8065_ = ~new_E8056_ & new_E8082_;
  assign new_E8066_ = ~new_E8058_ & new_E8070_;
  assign new_E8067_ = new_E8058_ & ~new_E8070_;
  assign new_E8068_ = new_E8044_ & ~new_E8045_;
  assign new_E8069_ = ~new_E8091_ | ~new_E8092_;
  assign new_E8070_ = new_E8084_ | new_E8086_;
  assign new_E8071_ = new_E8094_ | new_E8093_;
  assign new_E8072_ = new_E8088_ | new_E8087_;
  assign new_E8073_ = ~new_E8096_ | ~new_E8095_;
  assign new_E8074_ = ~new_E8097_ & new_E8098_;
  assign new_E8075_ = new_E8097_ & ~new_E8098_;
  assign new_E8076_ = ~new_E8044_ & new_E8045_;
  assign new_E8077_ = new_E8044_ & ~new_E8045_;
  assign new_E8078_ = ~new_E8060_ | new_E8070_;
  assign new_E8079_ = new_E8060_ & new_E8070_;
  assign new_E8080_ = ~new_E8060_ & ~new_E8070_;
  assign new_E8081_ = new_E8102_ | new_E8101_;
  assign new_E8082_ = new_E8048_ | new_E8081_;
  assign new_E8083_ = new_E8106_ | new_E8105_;
  assign new_E8084_ = ~new_E8048_ & new_E8083_;
  assign new_E8085_ = new_E8104_ | new_E8103_;
  assign new_E8086_ = new_E8048_ & new_E8085_;
  assign new_E8087_ = new_E8046_ & ~new_E8056_;
  assign new_E8088_ = ~new_E8046_ & new_E8056_;
  assign new_E8089_ = ~new_E8045_ | ~new_E8070_;
  assign new_E8090_ = new_E8056_ & new_E8089_;
  assign new_E8091_ = ~new_E8056_ & ~new_E8090_;
  assign new_E8092_ = new_E8056_ | new_E8089_;
  assign new_E8093_ = ~new_E8046_ & new_E8047_;
  assign new_E8094_ = new_E8046_ & ~new_E8047_;
  assign new_E8095_ = new_E8063_ | new_E8100_;
  assign new_E8096_ = ~new_E8063_ & ~new_E8099_;
  assign new_E8097_ = new_E8046_ | new_E8063_;
  assign new_E8098_ = new_E8046_ | new_E8047_;
  assign new_E8099_ = new_E8063_ & new_E8100_;
  assign new_E8100_ = ~new_E8045_ | ~new_E8070_;
  assign new_E8101_ = new_E8078_ & new_E8098_;
  assign new_E8102_ = ~new_E8078_ & ~new_E8098_;
  assign new_E8103_ = new_E8107_ | new_E8108_;
  assign new_E8104_ = ~new_E8049_ & new_E8063_;
  assign new_E8105_ = new_E8109_ | new_E8110_;
  assign new_E8106_ = new_E8049_ & new_E8063_;
  assign new_E8107_ = ~new_E8049_ & ~new_E8063_;
  assign new_E8108_ = new_E8049_ & ~new_E8063_;
  assign new_E8109_ = new_E8049_ & ~new_E8063_;
  assign new_E8110_ = ~new_E8049_ & new_E8063_;
  assign new_E8111_ = new_G317_;
  assign new_E8112_ = new_G384_;
  assign new_E8113_ = new_G451_;
  assign new_E8114_ = new_G518_;
  assign new_E8115_ = new_G585_;
  assign new_E8116_ = new_G652_;
  assign new_E8117_ = new_E8124_ & new_E8123_;
  assign new_E8118_ = new_E8126_ | new_E8125_;
  assign new_E8119_ = new_E8128_ | new_E8127_;
  assign new_E8120_ = new_E8130_ & new_E8129_;
  assign new_E8121_ = new_E8130_ & new_E8131_;
  assign new_E8122_ = new_E8123_ | new_E8132_;
  assign new_E8123_ = new_E8112_ | new_E8135_;
  assign new_E8124_ = new_E8134_ | new_E8133_;
  assign new_E8125_ = new_E8139_ & new_E8138_;
  assign new_E8126_ = new_E8137_ & new_E8136_;
  assign new_E8127_ = new_E8142_ | new_E8141_;
  assign new_E8128_ = new_E8137_ & new_E8140_;
  assign new_E8129_ = new_E8112_ | new_E8145_;
  assign new_E8130_ = new_E8144_ | new_E8143_;
  assign new_E8131_ = new_E8147_ | new_E8146_;
  assign new_E8132_ = ~new_E8123_ & new_E8149_;
  assign new_E8133_ = ~new_E8125_ & new_E8137_;
  assign new_E8134_ = new_E8125_ & ~new_E8137_;
  assign new_E8135_ = new_E8111_ & ~new_E8112_;
  assign new_E8136_ = ~new_E8158_ | ~new_E8159_;
  assign new_E8137_ = new_E8151_ | new_E8153_;
  assign new_E8138_ = new_E8161_ | new_E8160_;
  assign new_E8139_ = new_E8155_ | new_E8154_;
  assign new_E8140_ = ~new_E8163_ | ~new_E8162_;
  assign new_E8141_ = ~new_E8164_ & new_E8165_;
  assign new_E8142_ = new_E8164_ & ~new_E8165_;
  assign new_E8143_ = ~new_E8111_ & new_E8112_;
  assign new_E8144_ = new_E8111_ & ~new_E8112_;
  assign new_E8145_ = ~new_E8127_ | new_E8137_;
  assign new_E8146_ = new_E8127_ & new_E8137_;
  assign new_E8147_ = ~new_E8127_ & ~new_E8137_;
  assign new_E8148_ = new_E8169_ | new_E8168_;
  assign new_E8149_ = new_E8115_ | new_E8148_;
  assign new_E8150_ = new_E8173_ | new_E8172_;
  assign new_E8151_ = ~new_E8115_ & new_E8150_;
  assign new_E8152_ = new_E8171_ | new_E8170_;
  assign new_E8153_ = new_E8115_ & new_E8152_;
  assign new_E8154_ = new_E8113_ & ~new_E8123_;
  assign new_E8155_ = ~new_E8113_ & new_E8123_;
  assign new_E8156_ = ~new_E8112_ | ~new_E8137_;
  assign new_E8157_ = new_E8123_ & new_E8156_;
  assign new_E8158_ = ~new_E8123_ & ~new_E8157_;
  assign new_E8159_ = new_E8123_ | new_E8156_;
  assign new_E8160_ = ~new_E8113_ & new_E8114_;
  assign new_E8161_ = new_E8113_ & ~new_E8114_;
  assign new_E8162_ = new_E8130_ | new_E8167_;
  assign new_E8163_ = ~new_E8130_ & ~new_E8166_;
  assign new_E8164_ = new_E8113_ | new_E8130_;
  assign new_E8165_ = new_E8113_ | new_E8114_;
  assign new_E8166_ = new_E8130_ & new_E8167_;
  assign new_E8167_ = ~new_E8112_ | ~new_E8137_;
  assign new_E8168_ = new_E8145_ & new_E8165_;
  assign new_E8169_ = ~new_E8145_ & ~new_E8165_;
  assign new_E8170_ = new_E8174_ | new_E8175_;
  assign new_E8171_ = ~new_E8116_ & new_E8130_;
  assign new_E8172_ = new_E8176_ | new_E8177_;
  assign new_E8173_ = new_E8116_ & new_E8130_;
  assign new_E8174_ = ~new_E8116_ & ~new_E8130_;
  assign new_E8175_ = new_E8116_ & ~new_E8130_;
  assign new_E8176_ = new_E8116_ & ~new_E8130_;
  assign new_E8177_ = ~new_E8116_ & new_E8130_;
  assign new_E8178_ = new_G719_;
  assign new_E8179_ = new_G786_;
  assign new_E8180_ = new_G853_;
  assign new_E8181_ = new_G920_;
  assign new_E8182_ = new_G987_;
  assign new_E8183_ = new_G1054_;
  assign new_E8184_ = new_E8191_ & new_E8190_;
  assign new_E8185_ = new_E8193_ | new_E8192_;
  assign new_E8186_ = new_E8195_ | new_E8194_;
  assign new_E8187_ = new_E8197_ & new_E8196_;
  assign new_E8188_ = new_E8197_ & new_E8198_;
  assign new_E8189_ = new_E8190_ | new_E8199_;
  assign new_E8190_ = new_E8179_ | new_E8202_;
  assign new_E8191_ = new_E8201_ | new_E8200_;
  assign new_E8192_ = new_E8206_ & new_E8205_;
  assign new_E8193_ = new_E8204_ & new_E8203_;
  assign new_E8194_ = new_E8209_ | new_E8208_;
  assign new_E8195_ = new_E8204_ & new_E8207_;
  assign new_E8196_ = new_E8179_ | new_E8212_;
  assign new_E8197_ = new_E8211_ | new_E8210_;
  assign new_E8198_ = new_E8214_ | new_E8213_;
  assign new_E8199_ = ~new_E8190_ & new_E8216_;
  assign new_E8200_ = ~new_E8192_ & new_E8204_;
  assign new_E8201_ = new_E8192_ & ~new_E8204_;
  assign new_E8202_ = new_E8178_ & ~new_E8179_;
  assign new_E8203_ = ~new_E8225_ | ~new_E8226_;
  assign new_E8204_ = new_E8218_ | new_E8220_;
  assign new_E8205_ = new_E8228_ | new_E8227_;
  assign new_E8206_ = new_E8222_ | new_E8221_;
  assign new_E8207_ = ~new_E8230_ | ~new_E8229_;
  assign new_E8208_ = ~new_E8231_ & new_E8232_;
  assign new_E8209_ = new_E8231_ & ~new_E8232_;
  assign new_E8210_ = ~new_E8178_ & new_E8179_;
  assign new_E8211_ = new_E8178_ & ~new_E8179_;
  assign new_E8212_ = ~new_E8194_ | new_E8204_;
  assign new_E8213_ = new_E8194_ & new_E8204_;
  assign new_E8214_ = ~new_E8194_ & ~new_E8204_;
  assign new_E8215_ = new_E8236_ | new_E8235_;
  assign new_E8216_ = new_E8182_ | new_E8215_;
  assign new_E8217_ = new_E8240_ | new_E8239_;
  assign new_E8218_ = ~new_E8182_ & new_E8217_;
  assign new_E8219_ = new_E8238_ | new_E8237_;
  assign new_E8220_ = new_E8182_ & new_E8219_;
  assign new_E8221_ = new_E8180_ & ~new_E8190_;
  assign new_E8222_ = ~new_E8180_ & new_E8190_;
  assign new_E8223_ = ~new_E8179_ | ~new_E8204_;
  assign new_E8224_ = new_E8190_ & new_E8223_;
  assign new_E8225_ = ~new_E8190_ & ~new_E8224_;
  assign new_E8226_ = new_E8190_ | new_E8223_;
  assign new_E8227_ = ~new_E8180_ & new_E8181_;
  assign new_E8228_ = new_E8180_ & ~new_E8181_;
  assign new_E8229_ = new_E8197_ | new_E8234_;
  assign new_E8230_ = ~new_E8197_ & ~new_E8233_;
  assign new_E8231_ = new_E8180_ | new_E8197_;
  assign new_E8232_ = new_E8180_ | new_E8181_;
  assign new_E8233_ = new_E8197_ & new_E8234_;
  assign new_E8234_ = ~new_E8179_ | ~new_E8204_;
  assign new_E8235_ = new_E8212_ & new_E8232_;
  assign new_E8236_ = ~new_E8212_ & ~new_E8232_;
  assign new_E8237_ = new_E8241_ | new_E8242_;
  assign new_E8238_ = ~new_E8183_ & new_E8197_;
  assign new_E8239_ = new_E8243_ | new_E8244_;
  assign new_E8240_ = new_E8183_ & new_E8197_;
  assign new_E8241_ = ~new_E8183_ & ~new_E8197_;
  assign new_E8242_ = new_E8183_ & ~new_E8197_;
  assign new_E8243_ = new_E8183_ & ~new_E8197_;
  assign new_E8244_ = ~new_E8183_ & new_E8197_;
  assign new_E8245_ = new_G1121_;
  assign new_E8246_ = new_G1188_;
  assign new_E8247_ = new_G1255_;
  assign new_E8248_ = new_G1322_;
  assign new_E8249_ = new_G1389_;
  assign new_E8250_ = new_G1456_;
  assign new_E8251_ = new_E8258_ & new_E8257_;
  assign new_E8252_ = new_E8260_ | new_E8259_;
  assign new_E8253_ = new_E8262_ | new_E8261_;
  assign new_E8254_ = new_E8264_ & new_E8263_;
  assign new_E8255_ = new_E8264_ & new_E8265_;
  assign new_E8256_ = new_E8257_ | new_E8266_;
  assign new_E8257_ = new_E8246_ | new_E8269_;
  assign new_E8258_ = new_E8268_ | new_E8267_;
  assign new_E8259_ = new_E8273_ & new_E8272_;
  assign new_E8260_ = new_E8271_ & new_E8270_;
  assign new_E8261_ = new_E8276_ | new_E8275_;
  assign new_E8262_ = new_E8271_ & new_E8274_;
  assign new_E8263_ = new_E8246_ | new_E8279_;
  assign new_E8264_ = new_E8278_ | new_E8277_;
  assign new_E8265_ = new_E8281_ | new_E8280_;
  assign new_E8266_ = ~new_E8257_ & new_E8283_;
  assign new_E8267_ = ~new_E8259_ & new_E8271_;
  assign new_E8268_ = new_E8259_ & ~new_E8271_;
  assign new_E8269_ = new_E8245_ & ~new_E8246_;
  assign new_E8270_ = ~new_E8292_ | ~new_E8293_;
  assign new_E8271_ = new_E8285_ | new_E8287_;
  assign new_E8272_ = new_E8295_ | new_E8294_;
  assign new_E8273_ = new_E8289_ | new_E8288_;
  assign new_E8274_ = ~new_E8297_ | ~new_E8296_;
  assign new_E8275_ = ~new_E8298_ & new_E8299_;
  assign new_E8276_ = new_E8298_ & ~new_E8299_;
  assign new_E8277_ = ~new_E8245_ & new_E8246_;
  assign new_E8278_ = new_E8245_ & ~new_E8246_;
  assign new_E8279_ = ~new_E8261_ | new_E8271_;
  assign new_E8280_ = new_E8261_ & new_E8271_;
  assign new_E8281_ = ~new_E8261_ & ~new_E8271_;
  assign new_E8282_ = new_E8303_ | new_E8302_;
  assign new_E8283_ = new_E8249_ | new_E8282_;
  assign new_E8284_ = new_E8307_ | new_E8306_;
  assign new_E8285_ = ~new_E8249_ & new_E8284_;
  assign new_E8286_ = new_E8305_ | new_E8304_;
  assign new_E8287_ = new_E8249_ & new_E8286_;
  assign new_E8288_ = new_E8247_ & ~new_E8257_;
  assign new_E8289_ = ~new_E8247_ & new_E8257_;
  assign new_E8290_ = ~new_E8246_ | ~new_E8271_;
  assign new_E8291_ = new_E8257_ & new_E8290_;
  assign new_E8292_ = ~new_E8257_ & ~new_E8291_;
  assign new_E8293_ = new_E8257_ | new_E8290_;
  assign new_E8294_ = ~new_E8247_ & new_E8248_;
  assign new_E8295_ = new_E8247_ & ~new_E8248_;
  assign new_E8296_ = new_E8264_ | new_E8301_;
  assign new_E8297_ = ~new_E8264_ & ~new_E8300_;
  assign new_E8298_ = new_E8247_ | new_E8264_;
  assign new_E8299_ = new_E8247_ | new_E8248_;
  assign new_E8300_ = new_E8264_ & new_E8301_;
  assign new_E8301_ = ~new_E8246_ | ~new_E8271_;
  assign new_E8302_ = new_E8279_ & new_E8299_;
  assign new_E8303_ = ~new_E8279_ & ~new_E8299_;
  assign new_E8304_ = new_E8308_ | new_E8309_;
  assign new_E8305_ = ~new_E8250_ & new_E8264_;
  assign new_E8306_ = new_E8310_ | new_E8311_;
  assign new_E8307_ = new_E8250_ & new_E8264_;
  assign new_E8308_ = ~new_E8250_ & ~new_E8264_;
  assign new_E8309_ = new_E8250_ & ~new_E8264_;
  assign new_E8310_ = new_E8250_ & ~new_E8264_;
  assign new_E8311_ = ~new_E8250_ & new_E8264_;
  assign new_E8312_ = new_G1523_;
  assign new_E8313_ = new_G1590_;
  assign new_E8314_ = new_G1657_;
  assign new_E8315_ = new_G1724_;
  assign new_E8316_ = new_G1791_;
  assign new_E8317_ = new_G1858_;
  assign new_E8318_ = new_E8325_ & new_E8324_;
  assign new_E8319_ = new_E8327_ | new_E8326_;
  assign new_E8320_ = new_E8329_ | new_E8328_;
  assign new_E8321_ = new_E8331_ & new_E8330_;
  assign new_E8322_ = new_E8331_ & new_E8332_;
  assign new_E8323_ = new_E8324_ | new_E8333_;
  assign new_E8324_ = new_E8313_ | new_E8336_;
  assign new_E8325_ = new_E8335_ | new_E8334_;
  assign new_E8326_ = new_E8340_ & new_E8339_;
  assign new_E8327_ = new_E8338_ & new_E8337_;
  assign new_E8328_ = new_E8343_ | new_E8342_;
  assign new_E8329_ = new_E8338_ & new_E8341_;
  assign new_E8330_ = new_E8313_ | new_E8346_;
  assign new_E8331_ = new_E8345_ | new_E8344_;
  assign new_E8332_ = new_E8348_ | new_E8347_;
  assign new_E8333_ = ~new_E8324_ & new_E8350_;
  assign new_E8334_ = ~new_E8326_ & new_E8338_;
  assign new_E8335_ = new_E8326_ & ~new_E8338_;
  assign new_E8336_ = new_E8312_ & ~new_E8313_;
  assign new_E8337_ = ~new_E8359_ | ~new_E8360_;
  assign new_E8338_ = new_E8352_ | new_E8354_;
  assign new_E8339_ = new_E8362_ | new_E8361_;
  assign new_E8340_ = new_E8356_ | new_E8355_;
  assign new_E8341_ = ~new_E8364_ | ~new_E8363_;
  assign new_E8342_ = ~new_E8365_ & new_E8366_;
  assign new_E8343_ = new_E8365_ & ~new_E8366_;
  assign new_E8344_ = ~new_E8312_ & new_E8313_;
  assign new_E8345_ = new_E8312_ & ~new_E8313_;
  assign new_E8346_ = ~new_E8328_ | new_E8338_;
  assign new_E8347_ = new_E8328_ & new_E8338_;
  assign new_E8348_ = ~new_E8328_ & ~new_E8338_;
  assign new_E8349_ = new_E8370_ | new_E8369_;
  assign new_E8350_ = new_E8316_ | new_E8349_;
  assign new_E8351_ = new_E8374_ | new_E8373_;
  assign new_E8352_ = ~new_E8316_ & new_E8351_;
  assign new_E8353_ = new_E8372_ | new_E8371_;
  assign new_E8354_ = new_E8316_ & new_E8353_;
  assign new_E8355_ = new_E8314_ & ~new_E8324_;
  assign new_E8356_ = ~new_E8314_ & new_E8324_;
  assign new_E8357_ = ~new_E8313_ | ~new_E8338_;
  assign new_E8358_ = new_E8324_ & new_E8357_;
  assign new_E8359_ = ~new_E8324_ & ~new_E8358_;
  assign new_E8360_ = new_E8324_ | new_E8357_;
  assign new_E8361_ = ~new_E8314_ & new_E8315_;
  assign new_E8362_ = new_E8314_ & ~new_E8315_;
  assign new_E8363_ = new_E8331_ | new_E8368_;
  assign new_E8364_ = ~new_E8331_ & ~new_E8367_;
  assign new_E8365_ = new_E8314_ | new_E8331_;
  assign new_E8366_ = new_E8314_ | new_E8315_;
  assign new_E8367_ = new_E8331_ & new_E8368_;
  assign new_E8368_ = ~new_E8313_ | ~new_E8338_;
  assign new_E8369_ = new_E8346_ & new_E8366_;
  assign new_E8370_ = ~new_E8346_ & ~new_E8366_;
  assign new_E8371_ = new_E8375_ | new_E8376_;
  assign new_E8372_ = ~new_E8317_ & new_E8331_;
  assign new_E8373_ = new_E8377_ | new_E8378_;
  assign new_E8374_ = new_E8317_ & new_E8331_;
  assign new_E8375_ = ~new_E8317_ & ~new_E8331_;
  assign new_E8376_ = new_E8317_ & ~new_E8331_;
  assign new_E8377_ = new_E8317_ & ~new_E8331_;
  assign new_E8378_ = ~new_E8317_ & new_E8331_;
  assign new_E8379_ = new_G1925_;
  assign new_E8380_ = new_G1992_;
  assign new_E8381_ = new_G2059_;
  assign new_E8382_ = new_G2126_;
  assign new_E8383_ = new_G2193_;
  assign new_E8384_ = new_G2260_;
  assign new_E8385_ = new_E8392_ & new_E8391_;
  assign new_E8386_ = new_E8394_ | new_E8393_;
  assign new_E8387_ = new_E8396_ | new_E8395_;
  assign new_E8388_ = new_E8398_ & new_E8397_;
  assign new_E8389_ = new_E8398_ & new_E8399_;
  assign new_E8390_ = new_E8391_ | new_E8400_;
  assign new_E8391_ = new_E8380_ | new_E8403_;
  assign new_E8392_ = new_E8402_ | new_E8401_;
  assign new_E8393_ = new_E8407_ & new_E8406_;
  assign new_E8394_ = new_E8405_ & new_E8404_;
  assign new_E8395_ = new_E8410_ | new_E8409_;
  assign new_E8396_ = new_E8405_ & new_E8408_;
  assign new_E8397_ = new_E8380_ | new_E8413_;
  assign new_E8398_ = new_E8412_ | new_E8411_;
  assign new_E8399_ = new_E8415_ | new_E8414_;
  assign new_E8400_ = ~new_E8391_ & new_E8417_;
  assign new_E8401_ = ~new_E8393_ & new_E8405_;
  assign new_E8402_ = new_E8393_ & ~new_E8405_;
  assign new_E8403_ = new_E8379_ & ~new_E8380_;
  assign new_E8404_ = ~new_E8426_ | ~new_E8427_;
  assign new_E8405_ = new_E8419_ | new_E8421_;
  assign new_E8406_ = new_E8429_ | new_E8428_;
  assign new_E8407_ = new_E8423_ | new_E8422_;
  assign new_E8408_ = ~new_E8431_ | ~new_E8430_;
  assign new_E8409_ = ~new_E8432_ & new_E8433_;
  assign new_E8410_ = new_E8432_ & ~new_E8433_;
  assign new_E8411_ = ~new_E8379_ & new_E8380_;
  assign new_E8412_ = new_E8379_ & ~new_E8380_;
  assign new_E8413_ = ~new_E8395_ | new_E8405_;
  assign new_E8414_ = new_E8395_ & new_E8405_;
  assign new_E8415_ = ~new_E8395_ & ~new_E8405_;
  assign new_E8416_ = new_E8437_ | new_E8436_;
  assign new_E8417_ = new_E8383_ | new_E8416_;
  assign new_E8418_ = new_E8441_ | new_E8440_;
  assign new_E8419_ = ~new_E8383_ & new_E8418_;
  assign new_E8420_ = new_E8439_ | new_E8438_;
  assign new_E8421_ = new_E8383_ & new_E8420_;
  assign new_E8422_ = new_E8381_ & ~new_E8391_;
  assign new_E8423_ = ~new_E8381_ & new_E8391_;
  assign new_E8424_ = ~new_E8380_ | ~new_E8405_;
  assign new_E8425_ = new_E8391_ & new_E8424_;
  assign new_E8426_ = ~new_E8391_ & ~new_E8425_;
  assign new_E8427_ = new_E8391_ | new_E8424_;
  assign new_E8428_ = ~new_E8381_ & new_E8382_;
  assign new_E8429_ = new_E8381_ & ~new_E8382_;
  assign new_E8430_ = new_E8398_ | new_E8435_;
  assign new_E8431_ = ~new_E8398_ & ~new_E8434_;
  assign new_E8432_ = new_E8381_ | new_E8398_;
  assign new_E8433_ = new_E8381_ | new_E8382_;
  assign new_E8434_ = new_E8398_ & new_E8435_;
  assign new_E8435_ = ~new_E8380_ | ~new_E8405_;
  assign new_E8436_ = new_E8413_ & new_E8433_;
  assign new_E8437_ = ~new_E8413_ & ~new_E8433_;
  assign new_E8438_ = new_E8442_ | new_E8443_;
  assign new_E8439_ = ~new_E8384_ & new_E8398_;
  assign new_E8440_ = new_E8444_ | new_E8445_;
  assign new_E8441_ = new_E8384_ & new_E8398_;
  assign new_E8442_ = ~new_E8384_ & ~new_E8398_;
  assign new_E8443_ = new_E8384_ & ~new_E8398_;
  assign new_E8444_ = new_E8384_ & ~new_E8398_;
  assign new_E8445_ = ~new_E8384_ & new_E8398_;
  assign new_E8446_ = new_G2327_;
  assign new_E8447_ = new_G2394_;
  assign new_E8448_ = new_G2461_;
  assign new_E8449_ = new_G2528_;
  assign new_E8450_ = new_G2595_;
  assign new_E8451_ = new_G2662_;
  assign new_E8452_ = new_E8459_ & new_E8458_;
  assign new_E8453_ = new_E8461_ | new_E8460_;
  assign new_E8454_ = new_E8463_ | new_E8462_;
  assign new_E8455_ = new_E8465_ & new_E8464_;
  assign new_E8456_ = new_E8465_ & new_E8466_;
  assign new_E8457_ = new_E8458_ | new_E8467_;
  assign new_E8458_ = new_E8447_ | new_E8470_;
  assign new_E8459_ = new_E8469_ | new_E8468_;
  assign new_E8460_ = new_E8474_ & new_E8473_;
  assign new_E8461_ = new_E8472_ & new_E8471_;
  assign new_E8462_ = new_E8477_ | new_E8476_;
  assign new_E8463_ = new_E8472_ & new_E8475_;
  assign new_E8464_ = new_E8447_ | new_E8480_;
  assign new_E8465_ = new_E8479_ | new_E8478_;
  assign new_E8466_ = new_E8482_ | new_E8481_;
  assign new_E8467_ = ~new_E8458_ & new_E8484_;
  assign new_E8468_ = ~new_E8460_ & new_E8472_;
  assign new_E8469_ = new_E8460_ & ~new_E8472_;
  assign new_E8470_ = new_E8446_ & ~new_E8447_;
  assign new_E8471_ = ~new_E8493_ | ~new_E8494_;
  assign new_E8472_ = new_E8486_ | new_E8488_;
  assign new_E8473_ = new_E8496_ | new_E8495_;
  assign new_E8474_ = new_E8490_ | new_E8489_;
  assign new_E8475_ = ~new_E8498_ | ~new_E8497_;
  assign new_E8476_ = ~new_E8499_ & new_E8500_;
  assign new_E8477_ = new_E8499_ & ~new_E8500_;
  assign new_E8478_ = ~new_E8446_ & new_E8447_;
  assign new_E8479_ = new_E8446_ & ~new_E8447_;
  assign new_E8480_ = ~new_E8462_ | new_E8472_;
  assign new_E8481_ = new_E8462_ & new_E8472_;
  assign new_E8482_ = ~new_E8462_ & ~new_E8472_;
  assign new_E8483_ = new_E8504_ | new_E8503_;
  assign new_E8484_ = new_E8450_ | new_E8483_;
  assign new_E8485_ = new_E8508_ | new_E8507_;
  assign new_E8486_ = ~new_E8450_ & new_E8485_;
  assign new_E8487_ = new_E8506_ | new_E8505_;
  assign new_E8488_ = new_E8450_ & new_E8487_;
  assign new_E8489_ = new_E8448_ & ~new_E8458_;
  assign new_E8490_ = ~new_E8448_ & new_E8458_;
  assign new_E8491_ = ~new_E8447_ | ~new_E8472_;
  assign new_E8492_ = new_E8458_ & new_E8491_;
  assign new_E8493_ = ~new_E8458_ & ~new_E8492_;
  assign new_E8494_ = new_E8458_ | new_E8491_;
  assign new_E8495_ = ~new_E8448_ & new_E8449_;
  assign new_E8496_ = new_E8448_ & ~new_E8449_;
  assign new_E8497_ = new_E8465_ | new_E8502_;
  assign new_E8498_ = ~new_E8465_ & ~new_E8501_;
  assign new_E8499_ = new_E8448_ | new_E8465_;
  assign new_E8500_ = new_E8448_ | new_E8449_;
  assign new_E8501_ = new_E8465_ & new_E8502_;
  assign new_E8502_ = ~new_E8447_ | ~new_E8472_;
  assign new_E8503_ = new_E8480_ & new_E8500_;
  assign new_E8504_ = ~new_E8480_ & ~new_E8500_;
  assign new_E8505_ = new_E8509_ | new_E8510_;
  assign new_E8506_ = ~new_E8451_ & new_E8465_;
  assign new_E8507_ = new_E8511_ | new_E8512_;
  assign new_E8508_ = new_E8451_ & new_E8465_;
  assign new_E8509_ = ~new_E8451_ & ~new_E8465_;
  assign new_E8510_ = new_E8451_ & ~new_E8465_;
  assign new_E8511_ = new_E8451_ & ~new_E8465_;
  assign new_E8512_ = ~new_E8451_ & new_E8465_;
  assign new_E8513_ = new_G2729_;
  assign new_E8514_ = new_G2796_;
  assign new_E8515_ = new_G2863_;
  assign new_E8516_ = new_G2930_;
  assign new_E8517_ = new_G2997_;
  assign new_E8518_ = new_G3064_;
  assign new_E8519_ = new_E8526_ & new_E8525_;
  assign new_E8520_ = new_E8528_ | new_E8527_;
  assign new_E8521_ = new_E8530_ | new_E8529_;
  assign new_E8522_ = new_E8532_ & new_E8531_;
  assign new_E8523_ = new_E8532_ & new_E8533_;
  assign new_E8524_ = new_E8525_ | new_E8534_;
  assign new_E8525_ = new_E8514_ | new_E8537_;
  assign new_E8526_ = new_E8536_ | new_E8535_;
  assign new_E8527_ = new_E8541_ & new_E8540_;
  assign new_E8528_ = new_E8539_ & new_E8538_;
  assign new_E8529_ = new_E8544_ | new_E8543_;
  assign new_E8530_ = new_E8539_ & new_E8542_;
  assign new_E8531_ = new_E8514_ | new_E8547_;
  assign new_E8532_ = new_E8546_ | new_E8545_;
  assign new_E8533_ = new_E8549_ | new_E8548_;
  assign new_E8534_ = ~new_E8525_ & new_E8551_;
  assign new_E8535_ = ~new_E8527_ & new_E8539_;
  assign new_E8536_ = new_E8527_ & ~new_E8539_;
  assign new_E8537_ = new_E8513_ & ~new_E8514_;
  assign new_E8538_ = ~new_E8560_ | ~new_E8561_;
  assign new_E8539_ = new_E8553_ | new_E8555_;
  assign new_E8540_ = new_E8563_ | new_E8562_;
  assign new_E8541_ = new_E8557_ | new_E8556_;
  assign new_E8542_ = ~new_E8565_ | ~new_E8564_;
  assign new_E8543_ = ~new_E8566_ & new_E8567_;
  assign new_E8544_ = new_E8566_ & ~new_E8567_;
  assign new_E8545_ = ~new_E8513_ & new_E8514_;
  assign new_E8546_ = new_E8513_ & ~new_E8514_;
  assign new_E8547_ = ~new_E8529_ | new_E8539_;
  assign new_E8548_ = new_E8529_ & new_E8539_;
  assign new_E8549_ = ~new_E8529_ & ~new_E8539_;
  assign new_E8550_ = new_E8571_ | new_E8570_;
  assign new_E8551_ = new_E8517_ | new_E8550_;
  assign new_E8552_ = new_E8575_ | new_E8574_;
  assign new_E8553_ = ~new_E8517_ & new_E8552_;
  assign new_E8554_ = new_E8573_ | new_E8572_;
  assign new_E8555_ = new_E8517_ & new_E8554_;
  assign new_E8556_ = new_E8515_ & ~new_E8525_;
  assign new_E8557_ = ~new_E8515_ & new_E8525_;
  assign new_E8558_ = ~new_E8514_ | ~new_E8539_;
  assign new_E8559_ = new_E8525_ & new_E8558_;
  assign new_E8560_ = ~new_E8525_ & ~new_E8559_;
  assign new_E8561_ = new_E8525_ | new_E8558_;
  assign new_E8562_ = ~new_E8515_ & new_E8516_;
  assign new_E8563_ = new_E8515_ & ~new_E8516_;
  assign new_E8564_ = new_E8532_ | new_E8569_;
  assign new_E8565_ = ~new_E8532_ & ~new_E8568_;
  assign new_E8566_ = new_E8515_ | new_E8532_;
  assign new_E8567_ = new_E8515_ | new_E8516_;
  assign new_E8568_ = new_E8532_ & new_E8569_;
  assign new_E8569_ = ~new_E8514_ | ~new_E8539_;
  assign new_E8570_ = new_E8547_ & new_E8567_;
  assign new_E8571_ = ~new_E8547_ & ~new_E8567_;
  assign new_E8572_ = new_E8576_ | new_E8577_;
  assign new_E8573_ = ~new_E8518_ & new_E8532_;
  assign new_E8574_ = new_E8578_ | new_E8579_;
  assign new_E8575_ = new_E8518_ & new_E8532_;
  assign new_E8576_ = ~new_E8518_ & ~new_E8532_;
  assign new_E8577_ = new_E8518_ & ~new_E8532_;
  assign new_E8578_ = new_E8518_ & ~new_E8532_;
  assign new_E8579_ = ~new_E8518_ & new_E8532_;
  assign new_E8580_ = new_G3131_;
  assign new_E8581_ = new_G3198_;
  assign new_E8582_ = new_G3265_;
  assign new_E8583_ = new_G3332_;
  assign new_E8584_ = new_G3399_;
  assign new_E8585_ = new_G3466_;
  assign new_E8586_ = new_E8593_ & new_E8592_;
  assign new_E8587_ = new_E8595_ | new_E8594_;
  assign new_E8588_ = new_E8597_ | new_E8596_;
  assign new_E8589_ = new_E8599_ & new_E8598_;
  assign new_E8590_ = new_E8599_ & new_E8600_;
  assign new_E8591_ = new_E8592_ | new_E8601_;
  assign new_E8592_ = new_E8581_ | new_E8604_;
  assign new_E8593_ = new_E8603_ | new_E8602_;
  assign new_E8594_ = new_E8608_ & new_E8607_;
  assign new_E8595_ = new_E8606_ & new_E8605_;
  assign new_E8596_ = new_E8611_ | new_E8610_;
  assign new_E8597_ = new_E8606_ & new_E8609_;
  assign new_E8598_ = new_E8581_ | new_E8614_;
  assign new_E8599_ = new_E8613_ | new_E8612_;
  assign new_E8600_ = new_E8616_ | new_E8615_;
  assign new_E8601_ = ~new_E8592_ & new_E8618_;
  assign new_E8602_ = ~new_E8594_ & new_E8606_;
  assign new_E8603_ = new_E8594_ & ~new_E8606_;
  assign new_E8604_ = new_E8580_ & ~new_E8581_;
  assign new_E8605_ = ~new_E8627_ | ~new_E8628_;
  assign new_E8606_ = new_E8620_ | new_E8622_;
  assign new_E8607_ = new_E8630_ | new_E8629_;
  assign new_E8608_ = new_E8624_ | new_E8623_;
  assign new_E8609_ = ~new_E8632_ | ~new_E8631_;
  assign new_E8610_ = ~new_E8633_ & new_E8634_;
  assign new_E8611_ = new_E8633_ & ~new_E8634_;
  assign new_E8612_ = ~new_E8580_ & new_E8581_;
  assign new_E8613_ = new_E8580_ & ~new_E8581_;
  assign new_E8614_ = ~new_E8596_ | new_E8606_;
  assign new_E8615_ = new_E8596_ & new_E8606_;
  assign new_E8616_ = ~new_E8596_ & ~new_E8606_;
  assign new_E8617_ = new_E8638_ | new_E8637_;
  assign new_E8618_ = new_E8584_ | new_E8617_;
  assign new_E8619_ = new_E8642_ | new_E8641_;
  assign new_E8620_ = ~new_E8584_ & new_E8619_;
  assign new_E8621_ = new_E8640_ | new_E8639_;
  assign new_E8622_ = new_E8584_ & new_E8621_;
  assign new_E8623_ = new_E8582_ & ~new_E8592_;
  assign new_E8624_ = ~new_E8582_ & new_E8592_;
  assign new_E8625_ = ~new_E8581_ | ~new_E8606_;
  assign new_E8626_ = new_E8592_ & new_E8625_;
  assign new_E8627_ = ~new_E8592_ & ~new_E8626_;
  assign new_E8628_ = new_E8592_ | new_E8625_;
  assign new_E8629_ = ~new_E8582_ & new_E8583_;
  assign new_E8630_ = new_E8582_ & ~new_E8583_;
  assign new_E8631_ = new_E8599_ | new_E8636_;
  assign new_E8632_ = ~new_E8599_ & ~new_E8635_;
  assign new_E8633_ = new_E8582_ | new_E8599_;
  assign new_E8634_ = new_E8582_ | new_E8583_;
  assign new_E8635_ = new_E8599_ & new_E8636_;
  assign new_E8636_ = ~new_E8581_ | ~new_E8606_;
  assign new_E8637_ = new_E8614_ & new_E8634_;
  assign new_E8638_ = ~new_E8614_ & ~new_E8634_;
  assign new_E8639_ = new_E8643_ | new_E8644_;
  assign new_E8640_ = ~new_E8585_ & new_E8599_;
  assign new_E8641_ = new_E8645_ | new_E8646_;
  assign new_E8642_ = new_E8585_ & new_E8599_;
  assign new_E8643_ = ~new_E8585_ & ~new_E8599_;
  assign new_E8644_ = new_E8585_ & ~new_E8599_;
  assign new_E8645_ = new_E8585_ & ~new_E8599_;
  assign new_E8646_ = ~new_E8585_ & new_E8599_;
  assign new_E8647_ = new_G3533_;
  assign new_E8648_ = new_G3600_;
  assign new_E8649_ = new_G3667_;
  assign new_E8650_ = new_G3734_;
  assign new_E8651_ = new_G3801_;
  assign new_E8652_ = new_G3868_;
  assign new_E8653_ = new_E8660_ & new_E8659_;
  assign new_E8654_ = new_E8662_ | new_E8661_;
  assign new_E8655_ = new_E8664_ | new_E8663_;
  assign new_E8656_ = new_E8666_ & new_E8665_;
  assign new_E8657_ = new_E8666_ & new_E8667_;
  assign new_E8658_ = new_E8659_ | new_E8668_;
  assign new_E8659_ = new_E8648_ | new_E8671_;
  assign new_E8660_ = new_E8670_ | new_E8669_;
  assign new_E8661_ = new_E8675_ & new_E8674_;
  assign new_E8662_ = new_E8673_ & new_E8672_;
  assign new_E8663_ = new_E8678_ | new_E8677_;
  assign new_E8664_ = new_E8673_ & new_E8676_;
  assign new_E8665_ = new_E8648_ | new_E8681_;
  assign new_E8666_ = new_E8680_ | new_E8679_;
  assign new_E8667_ = new_E8683_ | new_E8682_;
  assign new_E8668_ = ~new_E8659_ & new_E8685_;
  assign new_E8669_ = ~new_E8661_ & new_E8673_;
  assign new_E8670_ = new_E8661_ & ~new_E8673_;
  assign new_E8671_ = new_E8647_ & ~new_E8648_;
  assign new_E8672_ = ~new_E8694_ | ~new_E8695_;
  assign new_E8673_ = new_E8687_ | new_E8689_;
  assign new_E8674_ = new_E8697_ | new_E8696_;
  assign new_E8675_ = new_E8691_ | new_E8690_;
  assign new_E8676_ = ~new_E8699_ | ~new_E8698_;
  assign new_E8677_ = ~new_E8700_ & new_E8701_;
  assign new_E8678_ = new_E8700_ & ~new_E8701_;
  assign new_E8679_ = ~new_E8647_ & new_E8648_;
  assign new_E8680_ = new_E8647_ & ~new_E8648_;
  assign new_E8681_ = ~new_E8663_ | new_E8673_;
  assign new_E8682_ = new_E8663_ & new_E8673_;
  assign new_E8683_ = ~new_E8663_ & ~new_E8673_;
  assign new_E8684_ = new_E8705_ | new_E8704_;
  assign new_E8685_ = new_E8651_ | new_E8684_;
  assign new_E8686_ = new_E8709_ | new_E8708_;
  assign new_E8687_ = ~new_E8651_ & new_E8686_;
  assign new_E8688_ = new_E8707_ | new_E8706_;
  assign new_E8689_ = new_E8651_ & new_E8688_;
  assign new_E8690_ = new_E8649_ & ~new_E8659_;
  assign new_E8691_ = ~new_E8649_ & new_E8659_;
  assign new_E8692_ = ~new_E8648_ | ~new_E8673_;
  assign new_E8693_ = new_E8659_ & new_E8692_;
  assign new_E8694_ = ~new_E8659_ & ~new_E8693_;
  assign new_E8695_ = new_E8659_ | new_E8692_;
  assign new_E8696_ = ~new_E8649_ & new_E8650_;
  assign new_E8697_ = new_E8649_ & ~new_E8650_;
  assign new_E8698_ = new_E8666_ | new_E8703_;
  assign new_E8699_ = ~new_E8666_ & ~new_E8702_;
  assign new_E8700_ = new_E8649_ | new_E8666_;
  assign new_E8701_ = new_E8649_ | new_E8650_;
  assign new_E8702_ = new_E8666_ & new_E8703_;
  assign new_E8703_ = ~new_E8648_ | ~new_E8673_;
  assign new_E8704_ = new_E8681_ & new_E8701_;
  assign new_E8705_ = ~new_E8681_ & ~new_E8701_;
  assign new_E8706_ = new_E8710_ | new_E8711_;
  assign new_E8707_ = ~new_E8652_ & new_E8666_;
  assign new_E8708_ = new_E8712_ | new_E8713_;
  assign new_E8709_ = new_E8652_ & new_E8666_;
  assign new_E8710_ = ~new_E8652_ & ~new_E8666_;
  assign new_E8711_ = new_E8652_ & ~new_E8666_;
  assign new_E8712_ = new_E8652_ & ~new_E8666_;
  assign new_E8713_ = ~new_E8652_ & new_E8666_;
  assign new_E8714_ = new_G3935_;
  assign new_E8715_ = new_G4002_;
  assign new_E8716_ = new_G4069_;
  assign new_E8717_ = new_G4136_;
  assign new_E8718_ = new_G4203_;
  assign new_E8719_ = new_G4270_;
  assign new_E8720_ = new_E8727_ & new_E8726_;
  assign new_E8721_ = new_E8729_ | new_E8728_;
  assign new_E8722_ = new_E8731_ | new_E8730_;
  assign new_E8723_ = new_E8733_ & new_E8732_;
  assign new_E8724_ = new_E8733_ & new_E8734_;
  assign new_E8725_ = new_E8726_ | new_E8735_;
  assign new_E8726_ = new_E8715_ | new_E8738_;
  assign new_E8727_ = new_E8737_ | new_E8736_;
  assign new_E8728_ = new_E8742_ & new_E8741_;
  assign new_E8729_ = new_E8740_ & new_E8739_;
  assign new_E8730_ = new_E8745_ | new_E8744_;
  assign new_E8731_ = new_E8740_ & new_E8743_;
  assign new_E8732_ = new_E8715_ | new_E8748_;
  assign new_E8733_ = new_E8747_ | new_E8746_;
  assign new_E8734_ = new_E8750_ | new_E8749_;
  assign new_E8735_ = ~new_E8726_ & new_E8752_;
  assign new_E8736_ = ~new_E8728_ & new_E8740_;
  assign new_E8737_ = new_E8728_ & ~new_E8740_;
  assign new_E8738_ = new_E8714_ & ~new_E8715_;
  assign new_E8739_ = ~new_E8761_ | ~new_E8762_;
  assign new_E8740_ = new_E8754_ | new_E8756_;
  assign new_E8741_ = new_E8764_ | new_E8763_;
  assign new_E8742_ = new_E8758_ | new_E8757_;
  assign new_E8743_ = ~new_E8766_ | ~new_E8765_;
  assign new_E8744_ = ~new_E8767_ & new_E8768_;
  assign new_E8745_ = new_E8767_ & ~new_E8768_;
  assign new_E8746_ = ~new_E8714_ & new_E8715_;
  assign new_E8747_ = new_E8714_ & ~new_E8715_;
  assign new_E8748_ = ~new_E8730_ | new_E8740_;
  assign new_E8749_ = new_E8730_ & new_E8740_;
  assign new_E8750_ = ~new_E8730_ & ~new_E8740_;
  assign new_E8751_ = new_E8772_ | new_E8771_;
  assign new_E8752_ = new_E8718_ | new_E8751_;
  assign new_E8753_ = new_E8776_ | new_E8775_;
  assign new_E8754_ = ~new_E8718_ & new_E8753_;
  assign new_E8755_ = new_E8774_ | new_E8773_;
  assign new_E8756_ = new_E8718_ & new_E8755_;
  assign new_E8757_ = new_E8716_ & ~new_E8726_;
  assign new_E8758_ = ~new_E8716_ & new_E8726_;
  assign new_E8759_ = ~new_E8715_ | ~new_E8740_;
  assign new_E8760_ = new_E8726_ & new_E8759_;
  assign new_E8761_ = ~new_E8726_ & ~new_E8760_;
  assign new_E8762_ = new_E8726_ | new_E8759_;
  assign new_E8763_ = ~new_E8716_ & new_E8717_;
  assign new_E8764_ = new_E8716_ & ~new_E8717_;
  assign new_E8765_ = new_E8733_ | new_E8770_;
  assign new_E8766_ = ~new_E8733_ & ~new_E8769_;
  assign new_E8767_ = new_E8716_ | new_E8733_;
  assign new_E8768_ = new_E8716_ | new_E8717_;
  assign new_E8769_ = new_E8733_ & new_E8770_;
  assign new_E8770_ = ~new_E8715_ | ~new_E8740_;
  assign new_E8771_ = new_E8748_ & new_E8768_;
  assign new_E8772_ = ~new_E8748_ & ~new_E8768_;
  assign new_E8773_ = new_E8777_ | new_E8778_;
  assign new_E8774_ = ~new_E8719_ & new_E8733_;
  assign new_E8775_ = new_E8779_ | new_E8780_;
  assign new_E8776_ = new_E8719_ & new_E8733_;
  assign new_E8777_ = ~new_E8719_ & ~new_E8733_;
  assign new_E8778_ = new_E8719_ & ~new_E8733_;
  assign new_E8779_ = new_E8719_ & ~new_E8733_;
  assign new_E8780_ = ~new_E8719_ & new_E8733_;
  assign new_E8781_ = new_G4337_;
  assign new_E8782_ = new_G4404_;
  assign new_E8783_ = new_G4471_;
  assign new_E8784_ = new_G4538_;
  assign new_E8785_ = new_G4605_;
  assign new_E8786_ = new_G4672_;
  assign new_E8787_ = new_E8794_ & new_E8793_;
  assign new_E8788_ = new_E8796_ | new_E8795_;
  assign new_E8789_ = new_E8798_ | new_E8797_;
  assign new_E8790_ = new_E8800_ & new_E8799_;
  assign new_E8791_ = new_E8800_ & new_E8801_;
  assign new_E8792_ = new_E8793_ | new_E8802_;
  assign new_E8793_ = new_E8782_ | new_E8805_;
  assign new_E8794_ = new_E8804_ | new_E8803_;
  assign new_E8795_ = new_E8809_ & new_E8808_;
  assign new_E8796_ = new_E8807_ & new_E8806_;
  assign new_E8797_ = new_E8812_ | new_E8811_;
  assign new_E8798_ = new_E8807_ & new_E8810_;
  assign new_E8799_ = new_E8782_ | new_E8815_;
  assign new_E8800_ = new_E8814_ | new_E8813_;
  assign new_E8801_ = new_E8817_ | new_E8816_;
  assign new_E8802_ = ~new_E8793_ & new_E8819_;
  assign new_E8803_ = ~new_E8795_ & new_E8807_;
  assign new_E8804_ = new_E8795_ & ~new_E8807_;
  assign new_E8805_ = new_E8781_ & ~new_E8782_;
  assign new_E8806_ = ~new_E8828_ | ~new_E8829_;
  assign new_E8807_ = new_E8821_ | new_E8823_;
  assign new_E8808_ = new_E8831_ | new_E8830_;
  assign new_E8809_ = new_E8825_ | new_E8824_;
  assign new_E8810_ = ~new_E8833_ | ~new_E8832_;
  assign new_E8811_ = ~new_E8834_ & new_E8835_;
  assign new_E8812_ = new_E8834_ & ~new_E8835_;
  assign new_E8813_ = ~new_E8781_ & new_E8782_;
  assign new_E8814_ = new_E8781_ & ~new_E8782_;
  assign new_E8815_ = ~new_E8797_ | new_E8807_;
  assign new_E8816_ = new_E8797_ & new_E8807_;
  assign new_E8817_ = ~new_E8797_ & ~new_E8807_;
  assign new_E8818_ = new_E8839_ | new_E8838_;
  assign new_E8819_ = new_E8785_ | new_E8818_;
  assign new_E8820_ = new_E8843_ | new_E8842_;
  assign new_E8821_ = ~new_E8785_ & new_E8820_;
  assign new_E8822_ = new_E8841_ | new_E8840_;
  assign new_E8823_ = new_E8785_ & new_E8822_;
  assign new_E8824_ = new_E8783_ & ~new_E8793_;
  assign new_E8825_ = ~new_E8783_ & new_E8793_;
  assign new_E8826_ = ~new_E8782_ | ~new_E8807_;
  assign new_E8827_ = new_E8793_ & new_E8826_;
  assign new_E8828_ = ~new_E8793_ & ~new_E8827_;
  assign new_E8829_ = new_E8793_ | new_E8826_;
  assign new_E8830_ = ~new_E8783_ & new_E8784_;
  assign new_E8831_ = new_E8783_ & ~new_E8784_;
  assign new_E8832_ = new_E8800_ | new_E8837_;
  assign new_E8833_ = ~new_E8800_ & ~new_E8836_;
  assign new_E8834_ = new_E8783_ | new_E8800_;
  assign new_E8835_ = new_E8783_ | new_E8784_;
  assign new_E8836_ = new_E8800_ & new_E8837_;
  assign new_E8837_ = ~new_E8782_ | ~new_E8807_;
  assign new_E8838_ = new_E8815_ & new_E8835_;
  assign new_E8839_ = ~new_E8815_ & ~new_E8835_;
  assign new_E8840_ = new_E8844_ | new_E8845_;
  assign new_E8841_ = ~new_E8786_ & new_E8800_;
  assign new_E8842_ = new_E8846_ | new_E8847_;
  assign new_E8843_ = new_E8786_ & new_E8800_;
  assign new_E8844_ = ~new_E8786_ & ~new_E8800_;
  assign new_E8845_ = new_E8786_ & ~new_E8800_;
  assign new_E8846_ = new_E8786_ & ~new_E8800_;
  assign new_E8847_ = ~new_E8786_ & new_E8800_;
  assign new_E8848_ = new_G4739_;
  assign new_E8849_ = new_G4806_;
  assign new_E8850_ = new_G4873_;
  assign new_E8851_ = new_G4940_;
  assign new_E8852_ = new_G5007_;
  assign new_E8853_ = new_G5074_;
  assign new_E8854_ = new_E8861_ & new_E8860_;
  assign new_E8855_ = new_E8863_ | new_E8862_;
  assign new_E8856_ = new_E8865_ | new_E8864_;
  assign new_E8857_ = new_E8867_ & new_E8866_;
  assign new_E8858_ = new_E8867_ & new_E8868_;
  assign new_E8859_ = new_E8860_ | new_E8869_;
  assign new_E8860_ = new_E8849_ | new_E8872_;
  assign new_E8861_ = new_E8871_ | new_E8870_;
  assign new_E8862_ = new_E8876_ & new_E8875_;
  assign new_E8863_ = new_E8874_ & new_E8873_;
  assign new_E8864_ = new_E8879_ | new_E8878_;
  assign new_E8865_ = new_E8874_ & new_E8877_;
  assign new_E8866_ = new_E8849_ | new_E8882_;
  assign new_E8867_ = new_E8881_ | new_E8880_;
  assign new_E8868_ = new_E8884_ | new_E8883_;
  assign new_E8869_ = ~new_E8860_ & new_E8886_;
  assign new_E8870_ = ~new_E8862_ & new_E8874_;
  assign new_E8871_ = new_E8862_ & ~new_E8874_;
  assign new_E8872_ = new_E8848_ & ~new_E8849_;
  assign new_E8873_ = ~new_E8895_ | ~new_E8896_;
  assign new_E8874_ = new_E8888_ | new_E8890_;
  assign new_E8875_ = new_E8898_ | new_E8897_;
  assign new_E8876_ = new_E8892_ | new_E8891_;
  assign new_E8877_ = ~new_E8900_ | ~new_E8899_;
  assign new_E8878_ = ~new_E8901_ & new_E8902_;
  assign new_E8879_ = new_E8901_ & ~new_E8902_;
  assign new_E8880_ = ~new_E8848_ & new_E8849_;
  assign new_E8881_ = new_E8848_ & ~new_E8849_;
  assign new_E8882_ = ~new_E8864_ | new_E8874_;
  assign new_E8883_ = new_E8864_ & new_E8874_;
  assign new_E8884_ = ~new_E8864_ & ~new_E8874_;
  assign new_E8885_ = new_E8906_ | new_E8905_;
  assign new_E8886_ = new_E8852_ | new_E8885_;
  assign new_E8887_ = new_E8910_ | new_E8909_;
  assign new_E8888_ = ~new_E8852_ & new_E8887_;
  assign new_E8889_ = new_E8908_ | new_E8907_;
  assign new_E8890_ = new_E8852_ & new_E8889_;
  assign new_E8891_ = new_E8850_ & ~new_E8860_;
  assign new_E8892_ = ~new_E8850_ & new_E8860_;
  assign new_E8893_ = ~new_E8849_ | ~new_E8874_;
  assign new_E8894_ = new_E8860_ & new_E8893_;
  assign new_E8895_ = ~new_E8860_ & ~new_E8894_;
  assign new_E8896_ = new_E8860_ | new_E8893_;
  assign new_E8897_ = ~new_E8850_ & new_E8851_;
  assign new_E8898_ = new_E8850_ & ~new_E8851_;
  assign new_E8899_ = new_E8867_ | new_E8904_;
  assign new_E8900_ = ~new_E8867_ & ~new_E8903_;
  assign new_E8901_ = new_E8850_ | new_E8867_;
  assign new_E8902_ = new_E8850_ | new_E8851_;
  assign new_E8903_ = new_E8867_ & new_E8904_;
  assign new_E8904_ = ~new_E8849_ | ~new_E8874_;
  assign new_E8905_ = new_E8882_ & new_E8902_;
  assign new_E8906_ = ~new_E8882_ & ~new_E8902_;
  assign new_E8907_ = new_E8911_ | new_E8912_;
  assign new_E8908_ = ~new_E8853_ & new_E8867_;
  assign new_E8909_ = new_E8913_ | new_E8914_;
  assign new_E8910_ = new_E8853_ & new_E8867_;
  assign new_E8911_ = ~new_E8853_ & ~new_E8867_;
  assign new_E8912_ = new_E8853_ & ~new_E8867_;
  assign new_E8913_ = new_E8853_ & ~new_E8867_;
  assign new_E8914_ = ~new_E8853_ & new_E8867_;
  assign new_E8915_ = new_G5141_;
  assign new_E8916_ = new_G5208_;
  assign new_E8917_ = new_G5275_;
  assign new_E8918_ = new_G5342_;
  assign new_E8919_ = new_G5409_;
  assign new_E8920_ = new_G5476_;
  assign new_E8921_ = new_E8928_ & new_E8927_;
  assign new_E8922_ = new_E8930_ | new_E8929_;
  assign new_E8923_ = new_E8932_ | new_E8931_;
  assign new_E8924_ = new_E8934_ & new_E8933_;
  assign new_E8925_ = new_E8934_ & new_E8935_;
  assign new_E8926_ = new_E8927_ | new_E8936_;
  assign new_E8927_ = new_E8916_ | new_E8939_;
  assign new_E8928_ = new_E8938_ | new_E8937_;
  assign new_E8929_ = new_E8943_ & new_E8942_;
  assign new_E8930_ = new_E8941_ & new_E8940_;
  assign new_E8931_ = new_E8946_ | new_E8945_;
  assign new_E8932_ = new_E8941_ & new_E8944_;
  assign new_E8933_ = new_E8916_ | new_E8949_;
  assign new_E8934_ = new_E8948_ | new_E8947_;
  assign new_E8935_ = new_E8951_ | new_E8950_;
  assign new_E8936_ = ~new_E8927_ & new_E8953_;
  assign new_E8937_ = ~new_E8929_ & new_E8941_;
  assign new_E8938_ = new_E8929_ & ~new_E8941_;
  assign new_E8939_ = new_E8915_ & ~new_E8916_;
  assign new_E8940_ = ~new_E8962_ | ~new_E8963_;
  assign new_E8941_ = new_E8955_ | new_E8957_;
  assign new_E8942_ = new_E8965_ | new_E8964_;
  assign new_E8943_ = new_E8959_ | new_E8958_;
  assign new_E8944_ = ~new_E8967_ | ~new_E8966_;
  assign new_E8945_ = ~new_E8968_ & new_E8969_;
  assign new_E8946_ = new_E8968_ & ~new_E8969_;
  assign new_E8947_ = ~new_E8915_ & new_E8916_;
  assign new_E8948_ = new_E8915_ & ~new_E8916_;
  assign new_E8949_ = ~new_E8931_ | new_E8941_;
  assign new_E8950_ = new_E8931_ & new_E8941_;
  assign new_E8951_ = ~new_E8931_ & ~new_E8941_;
  assign new_E8952_ = new_E8973_ | new_E8972_;
  assign new_E8953_ = new_E8919_ | new_E8952_;
  assign new_E8954_ = new_E8977_ | new_E8976_;
  assign new_E8955_ = ~new_E8919_ & new_E8954_;
  assign new_E8956_ = new_E8975_ | new_E8974_;
  assign new_E8957_ = new_E8919_ & new_E8956_;
  assign new_E8958_ = new_E8917_ & ~new_E8927_;
  assign new_E8959_ = ~new_E8917_ & new_E8927_;
  assign new_E8960_ = ~new_E8916_ | ~new_E8941_;
  assign new_E8961_ = new_E8927_ & new_E8960_;
  assign new_E8962_ = ~new_E8927_ & ~new_E8961_;
  assign new_E8963_ = new_E8927_ | new_E8960_;
  assign new_E8964_ = ~new_E8917_ & new_E8918_;
  assign new_E8965_ = new_E8917_ & ~new_E8918_;
  assign new_E8966_ = new_E8934_ | new_E8971_;
  assign new_E8967_ = ~new_E8934_ & ~new_E8970_;
  assign new_E8968_ = new_E8917_ | new_E8934_;
  assign new_E8969_ = new_E8917_ | new_E8918_;
  assign new_E8970_ = new_E8934_ & new_E8971_;
  assign new_E8971_ = ~new_E8916_ | ~new_E8941_;
  assign new_E8972_ = new_E8949_ & new_E8969_;
  assign new_E8973_ = ~new_E8949_ & ~new_E8969_;
  assign new_E8974_ = new_E8978_ | new_E8979_;
  assign new_E8975_ = ~new_E8920_ & new_E8934_;
  assign new_E8976_ = new_E8980_ | new_E8981_;
  assign new_E8977_ = new_E8920_ & new_E8934_;
  assign new_E8978_ = ~new_E8920_ & ~new_E8934_;
  assign new_E8979_ = new_E8920_ & ~new_E8934_;
  assign new_E8980_ = new_E8920_ & ~new_E8934_;
  assign new_E8981_ = ~new_E8920_ & new_E8934_;
  assign new_E8982_ = new_G5543_;
  assign new_E8983_ = new_G5610_;
  assign new_E8984_ = new_G5677_;
  assign new_E8985_ = new_G5744_;
  assign new_E8986_ = new_G5811_;
  assign new_E8987_ = new_G5878_;
  assign new_E8988_ = new_E8995_ & new_E8994_;
  assign new_E8989_ = new_E8997_ | new_E8996_;
  assign new_E8990_ = new_E8999_ | new_E8998_;
  assign new_E8991_ = new_E9001_ & new_E9000_;
  assign new_E8992_ = new_E9001_ & new_E9002_;
  assign new_E8993_ = new_E8994_ | new_E9003_;
  assign new_E8994_ = new_E8983_ | new_E9006_;
  assign new_E8995_ = new_E9005_ | new_E9004_;
  assign new_E8996_ = new_E9010_ & new_E9009_;
  assign new_E8997_ = new_E9008_ & new_E9007_;
  assign new_E8998_ = new_E9013_ | new_E9012_;
  assign new_E8999_ = new_E9008_ & new_E9011_;
  assign new_E9000_ = new_E8983_ | new_E9016_;
  assign new_E9001_ = new_E9015_ | new_E9014_;
  assign new_E9002_ = new_E9018_ | new_E9017_;
  assign new_E9003_ = ~new_E8994_ & new_E9020_;
  assign new_E9004_ = ~new_E8996_ & new_E9008_;
  assign new_E9005_ = new_E8996_ & ~new_E9008_;
  assign new_E9006_ = new_E8982_ & ~new_E8983_;
  assign new_E9007_ = ~new_E9029_ | ~new_E9030_;
  assign new_E9008_ = new_E9022_ | new_E9024_;
  assign new_E9009_ = new_E9032_ | new_E9031_;
  assign new_E9010_ = new_E9026_ | new_E9025_;
  assign new_E9011_ = ~new_E9034_ | ~new_E9033_;
  assign new_E9012_ = ~new_E9035_ & new_E9036_;
  assign new_E9013_ = new_E9035_ & ~new_E9036_;
  assign new_E9014_ = ~new_E8982_ & new_E8983_;
  assign new_E9015_ = new_E8982_ & ~new_E8983_;
  assign new_E9016_ = ~new_E8998_ | new_E9008_;
  assign new_E9017_ = new_E8998_ & new_E9008_;
  assign new_E9018_ = ~new_E8998_ & ~new_E9008_;
  assign new_E9019_ = new_E9040_ | new_E9039_;
  assign new_E9020_ = new_E8986_ | new_E9019_;
  assign new_E9021_ = new_E9044_ | new_E9043_;
  assign new_E9022_ = ~new_E8986_ & new_E9021_;
  assign new_E9023_ = new_E9042_ | new_E9041_;
  assign new_E9024_ = new_E8986_ & new_E9023_;
  assign new_E9025_ = new_E8984_ & ~new_E8994_;
  assign new_E9026_ = ~new_E8984_ & new_E8994_;
  assign new_E9027_ = ~new_E8983_ | ~new_E9008_;
  assign new_E9028_ = new_E8994_ & new_E9027_;
  assign new_E9029_ = ~new_E8994_ & ~new_E9028_;
  assign new_E9030_ = new_E8994_ | new_E9027_;
  assign new_E9031_ = ~new_E8984_ & new_E8985_;
  assign new_E9032_ = new_E8984_ & ~new_E8985_;
  assign new_E9033_ = new_E9001_ | new_E9038_;
  assign new_E9034_ = ~new_E9001_ & ~new_E9037_;
  assign new_E9035_ = new_E8984_ | new_E9001_;
  assign new_E9036_ = new_E8984_ | new_E8985_;
  assign new_E9037_ = new_E9001_ & new_E9038_;
  assign new_E9038_ = ~new_E8983_ | ~new_E9008_;
  assign new_E9039_ = new_E9016_ & new_E9036_;
  assign new_E9040_ = ~new_E9016_ & ~new_E9036_;
  assign new_E9041_ = new_E9045_ | new_E9046_;
  assign new_E9042_ = ~new_E8987_ & new_E9001_;
  assign new_E9043_ = new_E9047_ | new_E9048_;
  assign new_E9044_ = new_E8987_ & new_E9001_;
  assign new_E9045_ = ~new_E8987_ & ~new_E9001_;
  assign new_E9046_ = new_E8987_ & ~new_E9001_;
  assign new_E9047_ = new_E8987_ & ~new_E9001_;
  assign new_E9048_ = ~new_E8987_ & new_E9001_;
  assign new_E9049_ = new_F1468_;
  assign new_E9050_ = new_F1540_;
  assign new_E9051_ = new_F1607_;
  assign new_E9052_ = new_F1674_;
  assign new_E9053_ = new_F1741_;
  assign new_E9054_ = new_F1808_;
  assign new_E9055_ = new_E9062_ & new_E9061_;
  assign new_E9056_ = new_E9064_ | new_E9063_;
  assign new_E9057_ = new_E9066_ | new_E9065_;
  assign new_E9058_ = new_E9068_ & new_E9067_;
  assign new_E9059_ = new_E9068_ & new_E9069_;
  assign new_E9060_ = new_E9061_ | new_E9070_;
  assign new_E9061_ = new_E9050_ | new_E9073_;
  assign new_E9062_ = new_E9072_ | new_E9071_;
  assign new_E9063_ = new_E9077_ & new_E9076_;
  assign new_E9064_ = new_E9075_ & new_E9074_;
  assign new_E9065_ = new_E9080_ | new_E9079_;
  assign new_E9066_ = new_E9075_ & new_E9078_;
  assign new_E9067_ = new_E9050_ | new_E9083_;
  assign new_E9068_ = new_E9082_ | new_E9081_;
  assign new_E9069_ = new_E9085_ | new_E9084_;
  assign new_E9070_ = ~new_E9061_ & new_E9087_;
  assign new_E9071_ = ~new_E9063_ & new_E9075_;
  assign new_E9072_ = new_E9063_ & ~new_E9075_;
  assign new_E9073_ = new_E9049_ & ~new_E9050_;
  assign new_E9074_ = ~new_E9096_ | ~new_E9097_;
  assign new_E9075_ = new_E9089_ | new_E9091_;
  assign new_E9076_ = new_E9099_ | new_E9098_;
  assign new_E9077_ = new_E9093_ | new_E9092_;
  assign new_E9078_ = ~new_E9101_ | ~new_E9100_;
  assign new_E9079_ = ~new_E9102_ & new_E9103_;
  assign new_E9080_ = new_E9102_ & ~new_E9103_;
  assign new_E9081_ = ~new_E9049_ & new_E9050_;
  assign new_E9082_ = new_E9049_ & ~new_E9050_;
  assign new_E9083_ = ~new_E9065_ | new_E9075_;
  assign new_E9084_ = new_E9065_ & new_E9075_;
  assign new_E9085_ = ~new_E9065_ & ~new_E9075_;
  assign new_E9086_ = new_E9107_ | new_E9106_;
  assign new_E9087_ = new_E9053_ | new_E9086_;
  assign new_E9088_ = new_E9111_ | new_E9110_;
  assign new_E9089_ = ~new_E9053_ & new_E9088_;
  assign new_E9090_ = new_E9109_ | new_E9108_;
  assign new_E9091_ = new_E9053_ & new_E9090_;
  assign new_E9092_ = new_E9051_ & ~new_E9061_;
  assign new_E9093_ = ~new_E9051_ & new_E9061_;
  assign new_E9094_ = ~new_E9050_ | ~new_E9075_;
  assign new_E9095_ = new_E9061_ & new_E9094_;
  assign new_E9096_ = ~new_E9061_ & ~new_E9095_;
  assign new_E9097_ = new_E9061_ | new_E9094_;
  assign new_E9098_ = ~new_E9051_ & new_E9052_;
  assign new_E9099_ = new_E9051_ & ~new_E9052_;
  assign new_E9100_ = new_E9068_ | new_E9105_;
  assign new_E9101_ = ~new_E9068_ & ~new_E9104_;
  assign new_E9102_ = new_E9051_ | new_E9068_;
  assign new_E9103_ = new_E9051_ | new_E9052_;
  assign new_E9104_ = new_E9068_ & new_E9105_;
  assign new_E9105_ = ~new_E9050_ | ~new_E9075_;
  assign new_E9106_ = new_E9083_ & new_E9103_;
  assign new_E9107_ = ~new_E9083_ & ~new_E9103_;
  assign new_E9108_ = new_E9112_ | new_E9113_;
  assign new_E9109_ = ~new_E9054_ & new_E9068_;
  assign new_E9110_ = new_E9114_ | new_E9115_;
  assign new_E9111_ = new_E9054_ & new_E9068_;
  assign new_E9112_ = ~new_E9054_ & ~new_E9068_;
  assign new_E9113_ = new_E9054_ & ~new_E9068_;
  assign new_E9114_ = new_E9054_ & ~new_E9068_;
  assign new_E9115_ = ~new_E9054_ & new_E9068_;
  assign new_E9116_ = new_F1875_;
  assign new_E9117_ = new_F1942_;
  assign new_E9118_ = new_F2009_;
  assign new_E9119_ = new_F2076_;
  assign new_E9120_ = new_F2143_;
  assign new_E9121_ = new_F2210_;
  assign new_E9122_ = new_E9129_ & new_E9128_;
  assign new_E9123_ = new_E9131_ | new_E9130_;
  assign new_E9124_ = new_E9133_ | new_E9132_;
  assign new_E9125_ = new_E9135_ & new_E9134_;
  assign new_E9126_ = new_E9135_ & new_E9136_;
  assign new_E9127_ = new_E9128_ | new_E9137_;
  assign new_E9128_ = new_E9117_ | new_E9140_;
  assign new_E9129_ = new_E9139_ | new_E9138_;
  assign new_E9130_ = new_E9144_ & new_E9143_;
  assign new_E9131_ = new_E9142_ & new_E9141_;
  assign new_E9132_ = new_E9147_ | new_E9146_;
  assign new_E9133_ = new_E9142_ & new_E9145_;
  assign new_E9134_ = new_E9117_ | new_E9150_;
  assign new_E9135_ = new_E9149_ | new_E9148_;
  assign new_E9136_ = new_E9152_ | new_E9151_;
  assign new_E9137_ = ~new_E9128_ & new_E9154_;
  assign new_E9138_ = ~new_E9130_ & new_E9142_;
  assign new_E9139_ = new_E9130_ & ~new_E9142_;
  assign new_E9140_ = new_E9116_ & ~new_E9117_;
  assign new_E9141_ = ~new_E9163_ | ~new_E9164_;
  assign new_E9142_ = new_E9156_ | new_E9158_;
  assign new_E9143_ = new_E9166_ | new_E9165_;
  assign new_E9144_ = new_E9160_ | new_E9159_;
  assign new_E9145_ = ~new_E9168_ | ~new_E9167_;
  assign new_E9146_ = ~new_E9169_ & new_E9170_;
  assign new_E9147_ = new_E9169_ & ~new_E9170_;
  assign new_E9148_ = ~new_E9116_ & new_E9117_;
  assign new_E9149_ = new_E9116_ & ~new_E9117_;
  assign new_E9150_ = ~new_E9132_ | new_E9142_;
  assign new_E9151_ = new_E9132_ & new_E9142_;
  assign new_E9152_ = ~new_E9132_ & ~new_E9142_;
  assign new_E9153_ = new_E9174_ | new_E9173_;
  assign new_E9154_ = new_E9120_ | new_E9153_;
  assign new_E9155_ = new_E9178_ | new_E9177_;
  assign new_E9156_ = ~new_E9120_ & new_E9155_;
  assign new_E9157_ = new_E9176_ | new_E9175_;
  assign new_E9158_ = new_E9120_ & new_E9157_;
  assign new_E9159_ = new_E9118_ & ~new_E9128_;
  assign new_E9160_ = ~new_E9118_ & new_E9128_;
  assign new_E9161_ = ~new_E9117_ | ~new_E9142_;
  assign new_E9162_ = new_E9128_ & new_E9161_;
  assign new_E9163_ = ~new_E9128_ & ~new_E9162_;
  assign new_E9164_ = new_E9128_ | new_E9161_;
  assign new_E9165_ = ~new_E9118_ & new_E9119_;
  assign new_E9166_ = new_E9118_ & ~new_E9119_;
  assign new_E9167_ = new_E9135_ | new_E9172_;
  assign new_E9168_ = ~new_E9135_ & ~new_E9171_;
  assign new_E9169_ = new_E9118_ | new_E9135_;
  assign new_E9170_ = new_E9118_ | new_E9119_;
  assign new_E9171_ = new_E9135_ & new_E9172_;
  assign new_E9172_ = ~new_E9117_ | ~new_E9142_;
  assign new_E9173_ = new_E9150_ & new_E9170_;
  assign new_E9174_ = ~new_E9150_ & ~new_E9170_;
  assign new_E9175_ = new_E9179_ | new_E9180_;
  assign new_E9176_ = ~new_E9121_ & new_E9135_;
  assign new_E9177_ = new_E9181_ | new_E9182_;
  assign new_E9178_ = new_E9121_ & new_E9135_;
  assign new_E9179_ = ~new_E9121_ & ~new_E9135_;
  assign new_E9180_ = new_E9121_ & ~new_E9135_;
  assign new_E9181_ = new_E9121_ & ~new_E9135_;
  assign new_E9182_ = ~new_E9121_ & new_E9135_;
  assign new_E9183_ = new_F2277_;
  assign new_E9184_ = new_F2344_;
  assign new_E9185_ = new_F2411_;
  assign new_E9186_ = new_F2478_;
  assign new_E9187_ = new_F2545_;
  assign new_E9188_ = new_F2612_;
  assign new_E9189_ = new_E9196_ & new_E9195_;
  assign new_E9190_ = new_E9198_ | new_E9197_;
  assign new_E9191_ = new_E9200_ | new_E9199_;
  assign new_E9192_ = new_E9202_ & new_E9201_;
  assign new_E9193_ = new_E9202_ & new_E9203_;
  assign new_E9194_ = new_E9195_ | new_E9204_;
  assign new_E9195_ = new_E9184_ | new_E9207_;
  assign new_E9196_ = new_E9206_ | new_E9205_;
  assign new_E9197_ = new_E9211_ & new_E9210_;
  assign new_E9198_ = new_E9209_ & new_E9208_;
  assign new_E9199_ = new_E9214_ | new_E9213_;
  assign new_E9200_ = new_E9209_ & new_E9212_;
  assign new_E9201_ = new_E9184_ | new_E9217_;
  assign new_E9202_ = new_E9216_ | new_E9215_;
  assign new_E9203_ = new_E9219_ | new_E9218_;
  assign new_E9204_ = ~new_E9195_ & new_E9221_;
  assign new_E9205_ = ~new_E9197_ & new_E9209_;
  assign new_E9206_ = new_E9197_ & ~new_E9209_;
  assign new_E9207_ = new_E9183_ & ~new_E9184_;
  assign new_E9208_ = ~new_E9230_ | ~new_E9231_;
  assign new_E9209_ = new_E9223_ | new_E9225_;
  assign new_E9210_ = new_E9233_ | new_E9232_;
  assign new_E9211_ = new_E9227_ | new_E9226_;
  assign new_E9212_ = ~new_E9235_ | ~new_E9234_;
  assign new_E9213_ = ~new_E9236_ & new_E9237_;
  assign new_E9214_ = new_E9236_ & ~new_E9237_;
  assign new_E9215_ = ~new_E9183_ & new_E9184_;
  assign new_E9216_ = new_E9183_ & ~new_E9184_;
  assign new_E9217_ = ~new_E9199_ | new_E9209_;
  assign new_E9218_ = new_E9199_ & new_E9209_;
  assign new_E9219_ = ~new_E9199_ & ~new_E9209_;
  assign new_E9220_ = new_E9241_ | new_E9240_;
  assign new_E9221_ = new_E9187_ | new_E9220_;
  assign new_E9222_ = new_E9245_ | new_E9244_;
  assign new_E9223_ = ~new_E9187_ & new_E9222_;
  assign new_E9224_ = new_E9243_ | new_E9242_;
  assign new_E9225_ = new_E9187_ & new_E9224_;
  assign new_E9226_ = new_E9185_ & ~new_E9195_;
  assign new_E9227_ = ~new_E9185_ & new_E9195_;
  assign new_E9228_ = ~new_E9184_ | ~new_E9209_;
  assign new_E9229_ = new_E9195_ & new_E9228_;
  assign new_E9230_ = ~new_E9195_ & ~new_E9229_;
  assign new_E9231_ = new_E9195_ | new_E9228_;
  assign new_E9232_ = ~new_E9185_ & new_E9186_;
  assign new_E9233_ = new_E9185_ & ~new_E9186_;
  assign new_E9234_ = new_E9202_ | new_E9239_;
  assign new_E9235_ = ~new_E9202_ & ~new_E9238_;
  assign new_E9236_ = new_E9185_ | new_E9202_;
  assign new_E9237_ = new_E9185_ | new_E9186_;
  assign new_E9238_ = new_E9202_ & new_E9239_;
  assign new_E9239_ = ~new_E9184_ | ~new_E9209_;
  assign new_E9240_ = new_E9217_ & new_E9237_;
  assign new_E9241_ = ~new_E9217_ & ~new_E9237_;
  assign new_E9242_ = new_E9246_ | new_E9247_;
  assign new_E9243_ = ~new_E9188_ & new_E9202_;
  assign new_E9244_ = new_E9248_ | new_E9249_;
  assign new_E9245_ = new_E9188_ & new_E9202_;
  assign new_E9246_ = ~new_E9188_ & ~new_E9202_;
  assign new_E9247_ = new_E9188_ & ~new_E9202_;
  assign new_E9248_ = new_E9188_ & ~new_E9202_;
  assign new_E9249_ = ~new_E9188_ & new_E9202_;
  assign new_E9250_ = new_F2679_;
  assign new_E9251_ = new_F2746_;
  assign new_E9252_ = new_F2813_;
  assign new_E9253_ = new_F2880_;
  assign new_E9254_ = new_F2947_;
  assign new_E9255_ = new_F3014_;
  assign new_E9256_ = new_E9263_ & new_E9262_;
  assign new_E9257_ = new_E9265_ | new_E9264_;
  assign new_E9258_ = new_E9267_ | new_E9266_;
  assign new_E9259_ = new_E9269_ & new_E9268_;
  assign new_E9260_ = new_E9269_ & new_E9270_;
  assign new_E9261_ = new_E9262_ | new_E9271_;
  assign new_E9262_ = new_E9251_ | new_E9274_;
  assign new_E9263_ = new_E9273_ | new_E9272_;
  assign new_E9264_ = new_E9278_ & new_E9277_;
  assign new_E9265_ = new_E9276_ & new_E9275_;
  assign new_E9266_ = new_E9281_ | new_E9280_;
  assign new_E9267_ = new_E9276_ & new_E9279_;
  assign new_E9268_ = new_E9251_ | new_E9284_;
  assign new_E9269_ = new_E9283_ | new_E9282_;
  assign new_E9270_ = new_E9286_ | new_E9285_;
  assign new_E9271_ = ~new_E9262_ & new_E9288_;
  assign new_E9272_ = ~new_E9264_ & new_E9276_;
  assign new_E9273_ = new_E9264_ & ~new_E9276_;
  assign new_E9274_ = new_E9250_ & ~new_E9251_;
  assign new_E9275_ = ~new_E9297_ | ~new_E9298_;
  assign new_E9276_ = new_E9290_ | new_E9292_;
  assign new_E9277_ = new_E9300_ | new_E9299_;
  assign new_E9278_ = new_E9294_ | new_E9293_;
  assign new_E9279_ = ~new_E9302_ | ~new_E9301_;
  assign new_E9280_ = ~new_E9303_ & new_E9304_;
  assign new_E9281_ = new_E9303_ & ~new_E9304_;
  assign new_E9282_ = ~new_E9250_ & new_E9251_;
  assign new_E9283_ = new_E9250_ & ~new_E9251_;
  assign new_E9284_ = ~new_E9266_ | new_E9276_;
  assign new_E9285_ = new_E9266_ & new_E9276_;
  assign new_E9286_ = ~new_E9266_ & ~new_E9276_;
  assign new_E9287_ = new_E9308_ | new_E9307_;
  assign new_E9288_ = new_E9254_ | new_E9287_;
  assign new_E9289_ = new_E9312_ | new_E9311_;
  assign new_E9290_ = ~new_E9254_ & new_E9289_;
  assign new_E9291_ = new_E9310_ | new_E9309_;
  assign new_E9292_ = new_E9254_ & new_E9291_;
  assign new_E9293_ = new_E9252_ & ~new_E9262_;
  assign new_E9294_ = ~new_E9252_ & new_E9262_;
  assign new_E9295_ = ~new_E9251_ | ~new_E9276_;
  assign new_E9296_ = new_E9262_ & new_E9295_;
  assign new_E9297_ = ~new_E9262_ & ~new_E9296_;
  assign new_E9298_ = new_E9262_ | new_E9295_;
  assign new_E9299_ = ~new_E9252_ & new_E9253_;
  assign new_E9300_ = new_E9252_ & ~new_E9253_;
  assign new_E9301_ = new_E9269_ | new_E9306_;
  assign new_E9302_ = ~new_E9269_ & ~new_E9305_;
  assign new_E9303_ = new_E9252_ | new_E9269_;
  assign new_E9304_ = new_E9252_ | new_E9253_;
  assign new_E9305_ = new_E9269_ & new_E9306_;
  assign new_E9306_ = ~new_E9251_ | ~new_E9276_;
  assign new_E9307_ = new_E9284_ & new_E9304_;
  assign new_E9308_ = ~new_E9284_ & ~new_E9304_;
  assign new_E9309_ = new_E9313_ | new_E9314_;
  assign new_E9310_ = ~new_E9255_ & new_E9269_;
  assign new_E9311_ = new_E9315_ | new_E9316_;
  assign new_E9312_ = new_E9255_ & new_E9269_;
  assign new_E9313_ = ~new_E9255_ & ~new_E9269_;
  assign new_E9314_ = new_E9255_ & ~new_E9269_;
  assign new_E9315_ = new_E9255_ & ~new_E9269_;
  assign new_E9316_ = ~new_E9255_ & new_E9269_;
  assign new_E9317_ = new_F3081_;
  assign new_E9318_ = new_F3148_;
  assign new_E9319_ = new_F3215_;
  assign new_E9320_ = new_F3282_;
  assign new_E9321_ = new_F3349_;
  assign new_E9322_ = new_F3416_;
  assign new_E9323_ = new_E9330_ & new_E9329_;
  assign new_E9324_ = new_E9332_ | new_E9331_;
  assign new_E9325_ = new_E9334_ | new_E9333_;
  assign new_E9326_ = new_E9336_ & new_E9335_;
  assign new_E9327_ = new_E9336_ & new_E9337_;
  assign new_E9328_ = new_E9329_ | new_E9338_;
  assign new_E9329_ = new_E9318_ | new_E9341_;
  assign new_E9330_ = new_E9340_ | new_E9339_;
  assign new_E9331_ = new_E9345_ & new_E9344_;
  assign new_E9332_ = new_E9343_ & new_E9342_;
  assign new_E9333_ = new_E9348_ | new_E9347_;
  assign new_E9334_ = new_E9343_ & new_E9346_;
  assign new_E9335_ = new_E9318_ | new_E9351_;
  assign new_E9336_ = new_E9350_ | new_E9349_;
  assign new_E9337_ = new_E9353_ | new_E9352_;
  assign new_E9338_ = ~new_E9329_ & new_E9355_;
  assign new_E9339_ = ~new_E9331_ & new_E9343_;
  assign new_E9340_ = new_E9331_ & ~new_E9343_;
  assign new_E9341_ = new_E9317_ & ~new_E9318_;
  assign new_E9342_ = ~new_E9364_ | ~new_E9365_;
  assign new_E9343_ = new_E9357_ | new_E9359_;
  assign new_E9344_ = new_E9367_ | new_E9366_;
  assign new_E9345_ = new_E9361_ | new_E9360_;
  assign new_E9346_ = ~new_E9369_ | ~new_E9368_;
  assign new_E9347_ = ~new_E9370_ & new_E9371_;
  assign new_E9348_ = new_E9370_ & ~new_E9371_;
  assign new_E9349_ = ~new_E9317_ & new_E9318_;
  assign new_E9350_ = new_E9317_ & ~new_E9318_;
  assign new_E9351_ = ~new_E9333_ | new_E9343_;
  assign new_E9352_ = new_E9333_ & new_E9343_;
  assign new_E9353_ = ~new_E9333_ & ~new_E9343_;
  assign new_E9354_ = new_E9375_ | new_E9374_;
  assign new_E9355_ = new_E9321_ | new_E9354_;
  assign new_E9356_ = new_E9379_ | new_E9378_;
  assign new_E9357_ = ~new_E9321_ & new_E9356_;
  assign new_E9358_ = new_E9377_ | new_E9376_;
  assign new_E9359_ = new_E9321_ & new_E9358_;
  assign new_E9360_ = new_E9319_ & ~new_E9329_;
  assign new_E9361_ = ~new_E9319_ & new_E9329_;
  assign new_E9362_ = ~new_E9318_ | ~new_E9343_;
  assign new_E9363_ = new_E9329_ & new_E9362_;
  assign new_E9364_ = ~new_E9329_ & ~new_E9363_;
  assign new_E9365_ = new_E9329_ | new_E9362_;
  assign new_E9366_ = ~new_E9319_ & new_E9320_;
  assign new_E9367_ = new_E9319_ & ~new_E9320_;
  assign new_E9368_ = new_E9336_ | new_E9373_;
  assign new_E9369_ = ~new_E9336_ & ~new_E9372_;
  assign new_E9370_ = new_E9319_ | new_E9336_;
  assign new_E9371_ = new_E9319_ | new_E9320_;
  assign new_E9372_ = new_E9336_ & new_E9373_;
  assign new_E9373_ = ~new_E9318_ | ~new_E9343_;
  assign new_E9374_ = new_E9351_ & new_E9371_;
  assign new_E9375_ = ~new_E9351_ & ~new_E9371_;
  assign new_E9376_ = new_E9380_ | new_E9381_;
  assign new_E9377_ = ~new_E9322_ & new_E9336_;
  assign new_E9378_ = new_E9382_ | new_E9383_;
  assign new_E9379_ = new_E9322_ & new_E9336_;
  assign new_E9380_ = ~new_E9322_ & ~new_E9336_;
  assign new_E9381_ = new_E9322_ & ~new_E9336_;
  assign new_E9382_ = new_E9322_ & ~new_E9336_;
  assign new_E9383_ = ~new_E9322_ & new_E9336_;
  assign new_E9384_ = new_F3483_;
  assign new_E9385_ = new_F3550_;
  assign new_E9386_ = new_F3617_;
  assign new_E9387_ = new_F3684_;
  assign new_E9388_ = new_F3751_;
  assign new_E9389_ = new_F3818_;
  assign new_E9390_ = new_E9397_ & new_E9396_;
  assign new_E9391_ = new_E9399_ | new_E9398_;
  assign new_E9392_ = new_E9401_ | new_E9400_;
  assign new_E9393_ = new_E9403_ & new_E9402_;
  assign new_E9394_ = new_E9403_ & new_E9404_;
  assign new_E9395_ = new_E9396_ | new_E9405_;
  assign new_E9396_ = new_E9385_ | new_E9408_;
  assign new_E9397_ = new_E9407_ | new_E9406_;
  assign new_E9398_ = new_E9412_ & new_E9411_;
  assign new_E9399_ = new_E9410_ & new_E9409_;
  assign new_E9400_ = new_E9415_ | new_E9414_;
  assign new_E9401_ = new_E9410_ & new_E9413_;
  assign new_E9402_ = new_E9385_ | new_E9418_;
  assign new_E9403_ = new_E9417_ | new_E9416_;
  assign new_E9404_ = new_E9420_ | new_E9419_;
  assign new_E9405_ = ~new_E9396_ & new_E9422_;
  assign new_E9406_ = ~new_E9398_ & new_E9410_;
  assign new_E9407_ = new_E9398_ & ~new_E9410_;
  assign new_E9408_ = new_E9384_ & ~new_E9385_;
  assign new_E9409_ = ~new_E9431_ | ~new_E9432_;
  assign new_E9410_ = new_E9424_ | new_E9426_;
  assign new_E9411_ = new_E9434_ | new_E9433_;
  assign new_E9412_ = new_E9428_ | new_E9427_;
  assign new_E9413_ = ~new_E9436_ | ~new_E9435_;
  assign new_E9414_ = ~new_E9437_ & new_E9438_;
  assign new_E9415_ = new_E9437_ & ~new_E9438_;
  assign new_E9416_ = ~new_E9384_ & new_E9385_;
  assign new_E9417_ = new_E9384_ & ~new_E9385_;
  assign new_E9418_ = ~new_E9400_ | new_E9410_;
  assign new_E9419_ = new_E9400_ & new_E9410_;
  assign new_E9420_ = ~new_E9400_ & ~new_E9410_;
  assign new_E9421_ = new_E9442_ | new_E9441_;
  assign new_E9422_ = new_E9388_ | new_E9421_;
  assign new_E9423_ = new_E9446_ | new_E9445_;
  assign new_E9424_ = ~new_E9388_ & new_E9423_;
  assign new_E9425_ = new_E9444_ | new_E9443_;
  assign new_E9426_ = new_E9388_ & new_E9425_;
  assign new_E9427_ = new_E9386_ & ~new_E9396_;
  assign new_E9428_ = ~new_E9386_ & new_E9396_;
  assign new_E9429_ = ~new_E9385_ | ~new_E9410_;
  assign new_E9430_ = new_E9396_ & new_E9429_;
  assign new_E9431_ = ~new_E9396_ & ~new_E9430_;
  assign new_E9432_ = new_E9396_ | new_E9429_;
  assign new_E9433_ = ~new_E9386_ & new_E9387_;
  assign new_E9434_ = new_E9386_ & ~new_E9387_;
  assign new_E9435_ = new_E9403_ | new_E9440_;
  assign new_E9436_ = ~new_E9403_ & ~new_E9439_;
  assign new_E9437_ = new_E9386_ | new_E9403_;
  assign new_E9438_ = new_E9386_ | new_E9387_;
  assign new_E9439_ = new_E9403_ & new_E9440_;
  assign new_E9440_ = ~new_E9385_ | ~new_E9410_;
  assign new_E9441_ = new_E9418_ & new_E9438_;
  assign new_E9442_ = ~new_E9418_ & ~new_E9438_;
  assign new_E9443_ = new_E9447_ | new_E9448_;
  assign new_E9444_ = ~new_E9389_ & new_E9403_;
  assign new_E9445_ = new_E9449_ | new_E9450_;
  assign new_E9446_ = new_E9389_ & new_E9403_;
  assign new_E9447_ = ~new_E9389_ & ~new_E9403_;
  assign new_E9448_ = new_E9389_ & ~new_E9403_;
  assign new_E9449_ = new_E9389_ & ~new_E9403_;
  assign new_E9450_ = ~new_E9389_ & new_E9403_;
  assign new_E9451_ = new_F3885_;
  assign new_E9452_ = new_F3952_;
  assign new_E9453_ = new_F4019_;
  assign new_E9454_ = new_F4086_;
  assign new_E9455_ = new_F4153_;
  assign new_E9456_ = new_F4220_;
  assign new_E9457_ = new_E9464_ & new_E9463_;
  assign new_E9458_ = new_E9466_ | new_E9465_;
  assign new_E9459_ = new_E9468_ | new_E9467_;
  assign new_E9460_ = new_E9470_ & new_E9469_;
  assign new_E9461_ = new_E9470_ & new_E9471_;
  assign new_E9462_ = new_E9463_ | new_E9472_;
  assign new_E9463_ = new_E9452_ | new_E9475_;
  assign new_E9464_ = new_E9474_ | new_E9473_;
  assign new_E9465_ = new_E9479_ & new_E9478_;
  assign new_E9466_ = new_E9477_ & new_E9476_;
  assign new_E9467_ = new_E9482_ | new_E9481_;
  assign new_E9468_ = new_E9477_ & new_E9480_;
  assign new_E9469_ = new_E9452_ | new_E9485_;
  assign new_E9470_ = new_E9484_ | new_E9483_;
  assign new_E9471_ = new_E9487_ | new_E9486_;
  assign new_E9472_ = ~new_E9463_ & new_E9489_;
  assign new_E9473_ = ~new_E9465_ & new_E9477_;
  assign new_E9474_ = new_E9465_ & ~new_E9477_;
  assign new_E9475_ = new_E9451_ & ~new_E9452_;
  assign new_E9476_ = ~new_E9498_ | ~new_E9499_;
  assign new_E9477_ = new_E9491_ | new_E9493_;
  assign new_E9478_ = new_E9501_ | new_E9500_;
  assign new_E9479_ = new_E9495_ | new_E9494_;
  assign new_E9480_ = ~new_E9503_ | ~new_E9502_;
  assign new_E9481_ = ~new_E9504_ & new_E9505_;
  assign new_E9482_ = new_E9504_ & ~new_E9505_;
  assign new_E9483_ = ~new_E9451_ & new_E9452_;
  assign new_E9484_ = new_E9451_ & ~new_E9452_;
  assign new_E9485_ = ~new_E9467_ | new_E9477_;
  assign new_E9486_ = new_E9467_ & new_E9477_;
  assign new_E9487_ = ~new_E9467_ & ~new_E9477_;
  assign new_E9488_ = new_E9509_ | new_E9508_;
  assign new_E9489_ = new_E9455_ | new_E9488_;
  assign new_E9490_ = new_E9513_ | new_E9512_;
  assign new_E9491_ = ~new_E9455_ & new_E9490_;
  assign new_E9492_ = new_E9511_ | new_E9510_;
  assign new_E9493_ = new_E9455_ & new_E9492_;
  assign new_E9494_ = new_E9453_ & ~new_E9463_;
  assign new_E9495_ = ~new_E9453_ & new_E9463_;
  assign new_E9496_ = ~new_E9452_ | ~new_E9477_;
  assign new_E9497_ = new_E9463_ & new_E9496_;
  assign new_E9498_ = ~new_E9463_ & ~new_E9497_;
  assign new_E9499_ = new_E9463_ | new_E9496_;
  assign new_E9500_ = ~new_E9453_ & new_E9454_;
  assign new_E9501_ = new_E9453_ & ~new_E9454_;
  assign new_E9502_ = new_E9470_ | new_E9507_;
  assign new_E9503_ = ~new_E9470_ & ~new_E9506_;
  assign new_E9504_ = new_E9453_ | new_E9470_;
  assign new_E9505_ = new_E9453_ | new_E9454_;
  assign new_E9506_ = new_E9470_ & new_E9507_;
  assign new_E9507_ = ~new_E9452_ | ~new_E9477_;
  assign new_E9508_ = new_E9485_ & new_E9505_;
  assign new_E9509_ = ~new_E9485_ & ~new_E9505_;
  assign new_E9510_ = new_E9514_ | new_E9515_;
  assign new_E9511_ = ~new_E9456_ & new_E9470_;
  assign new_E9512_ = new_E9516_ | new_E9517_;
  assign new_E9513_ = new_E9456_ & new_E9470_;
  assign new_E9514_ = ~new_E9456_ & ~new_E9470_;
  assign new_E9515_ = new_E9456_ & ~new_E9470_;
  assign new_E9516_ = new_E9456_ & ~new_E9470_;
  assign new_E9517_ = ~new_E9456_ & new_E9470_;
  assign new_E9518_ = new_F4287_;
  assign new_E9519_ = new_F4354_;
  assign new_E9520_ = new_F4421_;
  assign new_E9521_ = new_F4488_;
  assign new_E9522_ = new_F4555_;
  assign new_E9523_ = new_F4622_;
  assign new_E9524_ = new_E9531_ & new_E9530_;
  assign new_E9525_ = new_E9533_ | new_E9532_;
  assign new_E9526_ = new_E9535_ | new_E9534_;
  assign new_E9527_ = new_E9537_ & new_E9536_;
  assign new_E9528_ = new_E9537_ & new_E9538_;
  assign new_E9529_ = new_E9530_ | new_E9539_;
  assign new_E9530_ = new_E9519_ | new_E9542_;
  assign new_E9531_ = new_E9541_ | new_E9540_;
  assign new_E9532_ = new_E9546_ & new_E9545_;
  assign new_E9533_ = new_E9544_ & new_E9543_;
  assign new_E9534_ = new_E9549_ | new_E9548_;
  assign new_E9535_ = new_E9544_ & new_E9547_;
  assign new_E9536_ = new_E9519_ | new_E9552_;
  assign new_E9537_ = new_E9551_ | new_E9550_;
  assign new_E9538_ = new_E9554_ | new_E9553_;
  assign new_E9539_ = ~new_E9530_ & new_E9556_;
  assign new_E9540_ = ~new_E9532_ & new_E9544_;
  assign new_E9541_ = new_E9532_ & ~new_E9544_;
  assign new_E9542_ = new_E9518_ & ~new_E9519_;
  assign new_E9543_ = ~new_E9565_ | ~new_E9566_;
  assign new_E9544_ = new_E9558_ | new_E9560_;
  assign new_E9545_ = new_E9568_ | new_E9567_;
  assign new_E9546_ = new_E9562_ | new_E9561_;
  assign new_E9547_ = ~new_E9570_ | ~new_E9569_;
  assign new_E9548_ = ~new_E9571_ & new_E9572_;
  assign new_E9549_ = new_E9571_ & ~new_E9572_;
  assign new_E9550_ = ~new_E9518_ & new_E9519_;
  assign new_E9551_ = new_E9518_ & ~new_E9519_;
  assign new_E9552_ = ~new_E9534_ | new_E9544_;
  assign new_E9553_ = new_E9534_ & new_E9544_;
  assign new_E9554_ = ~new_E9534_ & ~new_E9544_;
  assign new_E9555_ = new_E9576_ | new_E9575_;
  assign new_E9556_ = new_E9522_ | new_E9555_;
  assign new_E9557_ = new_E9580_ | new_E9579_;
  assign new_E9558_ = ~new_E9522_ & new_E9557_;
  assign new_E9559_ = new_E9578_ | new_E9577_;
  assign new_E9560_ = new_E9522_ & new_E9559_;
  assign new_E9561_ = new_E9520_ & ~new_E9530_;
  assign new_E9562_ = ~new_E9520_ & new_E9530_;
  assign new_E9563_ = ~new_E9519_ | ~new_E9544_;
  assign new_E9564_ = new_E9530_ & new_E9563_;
  assign new_E9565_ = ~new_E9530_ & ~new_E9564_;
  assign new_E9566_ = new_E9530_ | new_E9563_;
  assign new_E9567_ = ~new_E9520_ & new_E9521_;
  assign new_E9568_ = new_E9520_ & ~new_E9521_;
  assign new_E9569_ = new_E9537_ | new_E9574_;
  assign new_E9570_ = ~new_E9537_ & ~new_E9573_;
  assign new_E9571_ = new_E9520_ | new_E9537_;
  assign new_E9572_ = new_E9520_ | new_E9521_;
  assign new_E9573_ = new_E9537_ & new_E9574_;
  assign new_E9574_ = ~new_E9519_ | ~new_E9544_;
  assign new_E9575_ = new_E9552_ & new_E9572_;
  assign new_E9576_ = ~new_E9552_ & ~new_E9572_;
  assign new_E9577_ = new_E9581_ | new_E9582_;
  assign new_E9578_ = ~new_E9523_ & new_E9537_;
  assign new_E9579_ = new_E9583_ | new_E9584_;
  assign new_E9580_ = new_E9523_ & new_E9537_;
  assign new_E9581_ = ~new_E9523_ & ~new_E9537_;
  assign new_E9582_ = new_E9523_ & ~new_E9537_;
  assign new_E9583_ = new_E9523_ & ~new_E9537_;
  assign new_E9584_ = ~new_E9523_ & new_E9537_;
  assign new_E9585_ = new_F4689_;
  assign new_E9586_ = new_F4756_;
  assign new_E9587_ = new_F4823_;
  assign new_E9588_ = new_F4890_;
  assign new_E9589_ = new_F4957_;
  assign new_E9590_ = new_F5024_;
  assign new_E9591_ = new_E9598_ & new_E9597_;
  assign new_E9592_ = new_E9600_ | new_E9599_;
  assign new_E9593_ = new_E9602_ | new_E9601_;
  assign new_E9594_ = new_E9604_ & new_E9603_;
  assign new_E9595_ = new_E9604_ & new_E9605_;
  assign new_E9596_ = new_E9597_ | new_E9606_;
  assign new_E9597_ = new_E9586_ | new_E9609_;
  assign new_E9598_ = new_E9608_ | new_E9607_;
  assign new_E9599_ = new_E9613_ & new_E9612_;
  assign new_E9600_ = new_E9611_ & new_E9610_;
  assign new_E9601_ = new_E9616_ | new_E9615_;
  assign new_E9602_ = new_E9611_ & new_E9614_;
  assign new_E9603_ = new_E9586_ | new_E9619_;
  assign new_E9604_ = new_E9618_ | new_E9617_;
  assign new_E9605_ = new_E9621_ | new_E9620_;
  assign new_E9606_ = ~new_E9597_ & new_E9623_;
  assign new_E9607_ = ~new_E9599_ & new_E9611_;
  assign new_E9608_ = new_E9599_ & ~new_E9611_;
  assign new_E9609_ = new_E9585_ & ~new_E9586_;
  assign new_E9610_ = ~new_E9632_ | ~new_E9633_;
  assign new_E9611_ = new_E9625_ | new_E9627_;
  assign new_E9612_ = new_E9635_ | new_E9634_;
  assign new_E9613_ = new_E9629_ | new_E9628_;
  assign new_E9614_ = ~new_E9637_ | ~new_E9636_;
  assign new_E9615_ = ~new_E9638_ & new_E9639_;
  assign new_E9616_ = new_E9638_ & ~new_E9639_;
  assign new_E9617_ = ~new_E9585_ & new_E9586_;
  assign new_E9618_ = new_E9585_ & ~new_E9586_;
  assign new_E9619_ = ~new_E9601_ | new_E9611_;
  assign new_E9620_ = new_E9601_ & new_E9611_;
  assign new_E9621_ = ~new_E9601_ & ~new_E9611_;
  assign new_E9622_ = new_E9643_ | new_E9642_;
  assign new_E9623_ = new_E9589_ | new_E9622_;
  assign new_E9624_ = new_E9647_ | new_E9646_;
  assign new_E9625_ = ~new_E9589_ & new_E9624_;
  assign new_E9626_ = new_E9645_ | new_E9644_;
  assign new_E9627_ = new_E9589_ & new_E9626_;
  assign new_E9628_ = new_E9587_ & ~new_E9597_;
  assign new_E9629_ = ~new_E9587_ & new_E9597_;
  assign new_E9630_ = ~new_E9586_ | ~new_E9611_;
  assign new_E9631_ = new_E9597_ & new_E9630_;
  assign new_E9632_ = ~new_E9597_ & ~new_E9631_;
  assign new_E9633_ = new_E9597_ | new_E9630_;
  assign new_E9634_ = ~new_E9587_ & new_E9588_;
  assign new_E9635_ = new_E9587_ & ~new_E9588_;
  assign new_E9636_ = new_E9604_ | new_E9641_;
  assign new_E9637_ = ~new_E9604_ & ~new_E9640_;
  assign new_E9638_ = new_E9587_ | new_E9604_;
  assign new_E9639_ = new_E9587_ | new_E9588_;
  assign new_E9640_ = new_E9604_ & new_E9641_;
  assign new_E9641_ = ~new_E9586_ | ~new_E9611_;
  assign new_E9642_ = new_E9619_ & new_E9639_;
  assign new_E9643_ = ~new_E9619_ & ~new_E9639_;
  assign new_E9644_ = new_E9648_ | new_E9649_;
  assign new_E9645_ = ~new_E9590_ & new_E9604_;
  assign new_E9646_ = new_E9650_ | new_E9651_;
  assign new_E9647_ = new_E9590_ & new_E9604_;
  assign new_E9648_ = ~new_E9590_ & ~new_E9604_;
  assign new_E9649_ = new_E9590_ & ~new_E9604_;
  assign new_E9650_ = new_E9590_ & ~new_E9604_;
  assign new_E9651_ = ~new_E9590_ & new_E9604_;
  assign new_E9652_ = new_F5091_;
  assign new_E9653_ = new_F5158_;
  assign new_E9654_ = new_F5225_;
  assign new_E9655_ = new_F5292_;
  assign new_E9656_ = new_F5359_;
  assign new_E9657_ = new_F5426_;
  assign new_E9658_ = new_E9665_ & new_E9664_;
  assign new_E9659_ = new_E9667_ | new_E9666_;
  assign new_E9660_ = new_E9669_ | new_E9668_;
  assign new_E9661_ = new_E9671_ & new_E9670_;
  assign new_E9662_ = new_E9671_ & new_E9672_;
  assign new_E9663_ = new_E9664_ | new_E9673_;
  assign new_E9664_ = new_E9653_ | new_E9676_;
  assign new_E9665_ = new_E9675_ | new_E9674_;
  assign new_E9666_ = new_E9680_ & new_E9679_;
  assign new_E9667_ = new_E9678_ & new_E9677_;
  assign new_E9668_ = new_E9683_ | new_E9682_;
  assign new_E9669_ = new_E9678_ & new_E9681_;
  assign new_E9670_ = new_E9653_ | new_E9686_;
  assign new_E9671_ = new_E9685_ | new_E9684_;
  assign new_E9672_ = new_E9688_ | new_E9687_;
  assign new_E9673_ = ~new_E9664_ & new_E9690_;
  assign new_E9674_ = ~new_E9666_ & new_E9678_;
  assign new_E9675_ = new_E9666_ & ~new_E9678_;
  assign new_E9676_ = new_E9652_ & ~new_E9653_;
  assign new_E9677_ = ~new_E9699_ | ~new_E9700_;
  assign new_E9678_ = new_E9692_ | new_E9694_;
  assign new_E9679_ = new_E9702_ | new_E9701_;
  assign new_E9680_ = new_E9696_ | new_E9695_;
  assign new_E9681_ = ~new_E9704_ | ~new_E9703_;
  assign new_E9682_ = ~new_E9705_ & new_E9706_;
  assign new_E9683_ = new_E9705_ & ~new_E9706_;
  assign new_E9684_ = ~new_E9652_ & new_E9653_;
  assign new_E9685_ = new_E9652_ & ~new_E9653_;
  assign new_E9686_ = ~new_E9668_ | new_E9678_;
  assign new_E9687_ = new_E9668_ & new_E9678_;
  assign new_E9688_ = ~new_E9668_ & ~new_E9678_;
  assign new_E9689_ = new_E9710_ | new_E9709_;
  assign new_E9690_ = new_E9656_ | new_E9689_;
  assign new_E9691_ = new_E9714_ | new_E9713_;
  assign new_E9692_ = ~new_E9656_ & new_E9691_;
  assign new_E9693_ = new_E9712_ | new_E9711_;
  assign new_E9694_ = new_E9656_ & new_E9693_;
  assign new_E9695_ = new_E9654_ & ~new_E9664_;
  assign new_E9696_ = ~new_E9654_ & new_E9664_;
  assign new_E9697_ = ~new_E9653_ | ~new_E9678_;
  assign new_E9698_ = new_E9664_ & new_E9697_;
  assign new_E9699_ = ~new_E9664_ & ~new_E9698_;
  assign new_E9700_ = new_E9664_ | new_E9697_;
  assign new_E9701_ = ~new_E9654_ & new_E9655_;
  assign new_E9702_ = new_E9654_ & ~new_E9655_;
  assign new_E9703_ = new_E9671_ | new_E9708_;
  assign new_E9704_ = ~new_E9671_ & ~new_E9707_;
  assign new_E9705_ = new_E9654_ | new_E9671_;
  assign new_E9706_ = new_E9654_ | new_E9655_;
  assign new_E9707_ = new_E9671_ & new_E9708_;
  assign new_E9708_ = ~new_E9653_ | ~new_E9678_;
  assign new_E9709_ = new_E9686_ & new_E9706_;
  assign new_E9710_ = ~new_E9686_ & ~new_E9706_;
  assign new_E9711_ = new_E9715_ | new_E9716_;
  assign new_E9712_ = ~new_E9657_ & new_E9671_;
  assign new_E9713_ = new_E9717_ | new_E9718_;
  assign new_E9714_ = new_E9657_ & new_E9671_;
  assign new_E9715_ = ~new_E9657_ & ~new_E9671_;
  assign new_E9716_ = new_E9657_ & ~new_E9671_;
  assign new_E9717_ = new_E9657_ & ~new_E9671_;
  assign new_E9718_ = ~new_E9657_ & new_E9671_;
  assign new_E9719_ = new_F5493_;
  assign new_E9720_ = new_F5560_;
  assign new_E9721_ = new_F5627_;
  assign new_E9722_ = new_F5694_;
  assign new_E9723_ = new_F5761_;
  assign new_E9724_ = new_F5828_;
  assign new_E9725_ = new_E9732_ & new_E9731_;
  assign new_E9726_ = new_E9734_ | new_E9733_;
  assign new_E9727_ = new_E9736_ | new_E9735_;
  assign new_E9728_ = new_E9738_ & new_E9737_;
  assign new_E9729_ = new_E9738_ & new_E9739_;
  assign new_E9730_ = new_E9731_ | new_E9740_;
  assign new_E9731_ = new_E9720_ | new_E9743_;
  assign new_E9732_ = new_E9742_ | new_E9741_;
  assign new_E9733_ = new_E9747_ & new_E9746_;
  assign new_E9734_ = new_E9745_ & new_E9744_;
  assign new_E9735_ = new_E9750_ | new_E9749_;
  assign new_E9736_ = new_E9745_ & new_E9748_;
  assign new_E9737_ = new_E9720_ | new_E9753_;
  assign new_E9738_ = new_E9752_ | new_E9751_;
  assign new_E9739_ = new_E9755_ | new_E9754_;
  assign new_E9740_ = ~new_E9731_ & new_E9757_;
  assign new_E9741_ = ~new_E9733_ & new_E9745_;
  assign new_E9742_ = new_E9733_ & ~new_E9745_;
  assign new_E9743_ = new_E9719_ & ~new_E9720_;
  assign new_E9744_ = ~new_E9766_ | ~new_E9767_;
  assign new_E9745_ = new_E9759_ | new_E9761_;
  assign new_E9746_ = new_E9769_ | new_E9768_;
  assign new_E9747_ = new_E9763_ | new_E9762_;
  assign new_E9748_ = ~new_E9771_ | ~new_E9770_;
  assign new_E9749_ = ~new_E9772_ & new_E9773_;
  assign new_E9750_ = new_E9772_ & ~new_E9773_;
  assign new_E9751_ = ~new_E9719_ & new_E9720_;
  assign new_E9752_ = new_E9719_ & ~new_E9720_;
  assign new_E9753_ = ~new_E9735_ | new_E9745_;
  assign new_E9754_ = new_E9735_ & new_E9745_;
  assign new_E9755_ = ~new_E9735_ & ~new_E9745_;
  assign new_E9756_ = new_E9777_ | new_E9776_;
  assign new_E9757_ = new_E9723_ | new_E9756_;
  assign new_E9758_ = new_E9781_ | new_E9780_;
  assign new_E9759_ = ~new_E9723_ & new_E9758_;
  assign new_E9760_ = new_E9779_ | new_E9778_;
  assign new_E9761_ = new_E9723_ & new_E9760_;
  assign new_E9762_ = new_E9721_ & ~new_E9731_;
  assign new_E9763_ = ~new_E9721_ & new_E9731_;
  assign new_E9764_ = ~new_E9720_ | ~new_E9745_;
  assign new_E9765_ = new_E9731_ & new_E9764_;
  assign new_E9766_ = ~new_E9731_ & ~new_E9765_;
  assign new_E9767_ = new_E9731_ | new_E9764_;
  assign new_E9768_ = ~new_E9721_ & new_E9722_;
  assign new_E9769_ = new_E9721_ & ~new_E9722_;
  assign new_E9770_ = new_E9738_ | new_E9775_;
  assign new_E9771_ = ~new_E9738_ & ~new_E9774_;
  assign new_E9772_ = new_E9721_ | new_E9738_;
  assign new_E9773_ = new_E9721_ | new_E9722_;
  assign new_E9774_ = new_E9738_ & new_E9775_;
  assign new_E9775_ = ~new_E9720_ | ~new_E9745_;
  assign new_E9776_ = new_E9753_ & new_E9773_;
  assign new_E9777_ = ~new_E9753_ & ~new_E9773_;
  assign new_E9778_ = new_E9782_ | new_E9783_;
  assign new_E9779_ = ~new_E9724_ & new_E9738_;
  assign new_E9780_ = new_E9784_ | new_E9785_;
  assign new_E9781_ = new_E9724_ & new_E9738_;
  assign new_E9782_ = ~new_E9724_ & ~new_E9738_;
  assign new_E9783_ = new_E9724_ & ~new_E9738_;
  assign new_E9784_ = new_E9724_ & ~new_E9738_;
  assign new_E9785_ = ~new_E9724_ & new_E9738_;
  assign new_E9786_ = new_F5895_;
  assign new_E9787_ = new_F5962_;
  assign new_E9788_ = new_F6029_;
  assign new_E9789_ = new_F6096_;
  assign new_E9790_ = new_F6163_;
  assign new_E9791_ = new_F6230_;
  assign new_E9792_ = new_E9799_ & new_E9798_;
  assign new_E9793_ = new_E9801_ | new_E9800_;
  assign new_E9794_ = new_E9803_ | new_E9802_;
  assign new_E9795_ = new_E9805_ & new_E9804_;
  assign new_E9796_ = new_E9805_ & new_E9806_;
  assign new_E9797_ = new_E9798_ | new_E9807_;
  assign new_E9798_ = new_E9787_ | new_E9810_;
  assign new_E9799_ = new_E9809_ | new_E9808_;
  assign new_E9800_ = new_E9814_ & new_E9813_;
  assign new_E9801_ = new_E9812_ & new_E9811_;
  assign new_E9802_ = new_E9817_ | new_E9816_;
  assign new_E9803_ = new_E9812_ & new_E9815_;
  assign new_E9804_ = new_E9787_ | new_E9820_;
  assign new_E9805_ = new_E9819_ | new_E9818_;
  assign new_E9806_ = new_E9822_ | new_E9821_;
  assign new_E9807_ = ~new_E9798_ & new_E9824_;
  assign new_E9808_ = ~new_E9800_ & new_E9812_;
  assign new_E9809_ = new_E9800_ & ~new_E9812_;
  assign new_E9810_ = new_E9786_ & ~new_E9787_;
  assign new_E9811_ = ~new_E9833_ | ~new_E9834_;
  assign new_E9812_ = new_E9826_ | new_E9828_;
  assign new_E9813_ = new_E9836_ | new_E9835_;
  assign new_E9814_ = new_E9830_ | new_E9829_;
  assign new_E9815_ = ~new_E9838_ | ~new_E9837_;
  assign new_E9816_ = ~new_E9839_ & new_E9840_;
  assign new_E9817_ = new_E9839_ & ~new_E9840_;
  assign new_E9818_ = ~new_E9786_ & new_E9787_;
  assign new_E9819_ = new_E9786_ & ~new_E9787_;
  assign new_E9820_ = ~new_E9802_ | new_E9812_;
  assign new_E9821_ = new_E9802_ & new_E9812_;
  assign new_E9822_ = ~new_E9802_ & ~new_E9812_;
  assign new_E9823_ = new_E9844_ | new_E9843_;
  assign new_E9824_ = new_E9790_ | new_E9823_;
  assign new_E9825_ = new_E9848_ | new_E9847_;
  assign new_E9826_ = ~new_E9790_ & new_E9825_;
  assign new_E9827_ = new_E9846_ | new_E9845_;
  assign new_E9828_ = new_E9790_ & new_E9827_;
  assign new_E9829_ = new_E9788_ & ~new_E9798_;
  assign new_E9830_ = ~new_E9788_ & new_E9798_;
  assign new_E9831_ = ~new_E9787_ | ~new_E9812_;
  assign new_E9832_ = new_E9798_ & new_E9831_;
  assign new_E9833_ = ~new_E9798_ & ~new_E9832_;
  assign new_E9834_ = new_E9798_ | new_E9831_;
  assign new_E9835_ = ~new_E9788_ & new_E9789_;
  assign new_E9836_ = new_E9788_ & ~new_E9789_;
  assign new_E9837_ = new_E9805_ | new_E9842_;
  assign new_E9838_ = ~new_E9805_ & ~new_E9841_;
  assign new_E9839_ = new_E9788_ | new_E9805_;
  assign new_E9840_ = new_E9788_ | new_E9789_;
  assign new_E9841_ = new_E9805_ & new_E9842_;
  assign new_E9842_ = ~new_E9787_ | ~new_E9812_;
  assign new_E9843_ = new_E9820_ & new_E9840_;
  assign new_E9844_ = ~new_E9820_ & ~new_E9840_;
  assign new_E9845_ = new_E9849_ | new_E9850_;
  assign new_E9846_ = ~new_E9791_ & new_E9805_;
  assign new_E9847_ = new_E9851_ | new_E9852_;
  assign new_E9848_ = new_E9791_ & new_E9805_;
  assign new_E9849_ = ~new_E9791_ & ~new_E9805_;
  assign new_E9850_ = new_E9791_ & ~new_E9805_;
  assign new_E9851_ = new_E9791_ & ~new_E9805_;
  assign new_E9852_ = ~new_E9791_ & new_E9805_;
  assign new_E9853_ = new_F6297_;
  assign new_E9854_ = new_F6364_;
  assign new_E9855_ = new_F6431_;
  assign new_E9856_ = new_F6498_;
  assign new_E9857_ = new_F6565_;
  assign new_E9858_ = new_F6632_;
  assign new_E9859_ = new_E9866_ & new_E9865_;
  assign new_E9860_ = new_E9868_ | new_E9867_;
  assign new_E9861_ = new_E9870_ | new_E9869_;
  assign new_E9862_ = new_E9872_ & new_E9871_;
  assign new_E9863_ = new_E9872_ & new_E9873_;
  assign new_E9864_ = new_E9865_ | new_E9874_;
  assign new_E9865_ = new_E9854_ | new_E9877_;
  assign new_E9866_ = new_E9876_ | new_E9875_;
  assign new_E9867_ = new_E9881_ & new_E9880_;
  assign new_E9868_ = new_E9879_ & new_E9878_;
  assign new_E9869_ = new_E9884_ | new_E9883_;
  assign new_E9870_ = new_E9879_ & new_E9882_;
  assign new_E9871_ = new_E9854_ | new_E9887_;
  assign new_E9872_ = new_E9886_ | new_E9885_;
  assign new_E9873_ = new_E9889_ | new_E9888_;
  assign new_E9874_ = ~new_E9865_ & new_E9891_;
  assign new_E9875_ = ~new_E9867_ & new_E9879_;
  assign new_E9876_ = new_E9867_ & ~new_E9879_;
  assign new_E9877_ = new_E9853_ & ~new_E9854_;
  assign new_E9878_ = ~new_E9900_ | ~new_E9901_;
  assign new_E9879_ = new_E9893_ | new_E9895_;
  assign new_E9880_ = new_E9903_ | new_E9902_;
  assign new_E9881_ = new_E9897_ | new_E9896_;
  assign new_E9882_ = ~new_E9905_ | ~new_E9904_;
  assign new_E9883_ = ~new_E9906_ & new_E9907_;
  assign new_E9884_ = new_E9906_ & ~new_E9907_;
  assign new_E9885_ = ~new_E9853_ & new_E9854_;
  assign new_E9886_ = new_E9853_ & ~new_E9854_;
  assign new_E9887_ = ~new_E9869_ | new_E9879_;
  assign new_E9888_ = new_E9869_ & new_E9879_;
  assign new_E9889_ = ~new_E9869_ & ~new_E9879_;
  assign new_E9890_ = new_E9911_ | new_E9910_;
  assign new_E9891_ = new_E9857_ | new_E9890_;
  assign new_E9892_ = new_E9915_ | new_E9914_;
  assign new_E9893_ = ~new_E9857_ & new_E9892_;
  assign new_E9894_ = new_E9913_ | new_E9912_;
  assign new_E9895_ = new_E9857_ & new_E9894_;
  assign new_E9896_ = new_E9855_ & ~new_E9865_;
  assign new_E9897_ = ~new_E9855_ & new_E9865_;
  assign new_E9898_ = ~new_E9854_ | ~new_E9879_;
  assign new_E9899_ = new_E9865_ & new_E9898_;
  assign new_E9900_ = ~new_E9865_ & ~new_E9899_;
  assign new_E9901_ = new_E9865_ | new_E9898_;
  assign new_E9902_ = ~new_E9855_ & new_E9856_;
  assign new_E9903_ = new_E9855_ & ~new_E9856_;
  assign new_E9904_ = new_E9872_ | new_E9909_;
  assign new_E9905_ = ~new_E9872_ & ~new_E9908_;
  assign new_E9906_ = new_E9855_ | new_E9872_;
  assign new_E9907_ = new_E9855_ | new_E9856_;
  assign new_E9908_ = new_E9872_ & new_E9909_;
  assign new_E9909_ = ~new_E9854_ | ~new_E9879_;
  assign new_E9910_ = new_E9887_ & new_E9907_;
  assign new_E9911_ = ~new_E9887_ & ~new_E9907_;
  assign new_E9912_ = new_E9916_ | new_E9917_;
  assign new_E9913_ = ~new_E9858_ & new_E9872_;
  assign new_E9914_ = new_E9918_ | new_E9919_;
  assign new_E9915_ = new_E9858_ & new_E9872_;
  assign new_E9916_ = ~new_E9858_ & ~new_E9872_;
  assign new_E9917_ = new_E9858_ & ~new_E9872_;
  assign new_E9918_ = new_E9858_ & ~new_E9872_;
  assign new_E9919_ = ~new_E9858_ & new_E9872_;
  assign new_E9920_ = new_F6699_;
  assign new_E9921_ = new_F6766_;
  assign new_E9922_ = new_F6833_;
  assign new_E9923_ = new_F6900_;
  assign new_E9924_ = new_F6967_;
  assign new_E9925_ = new_F7034_;
  assign new_E9926_ = new_E9933_ & new_E9932_;
  assign new_E9927_ = new_E9935_ | new_E9934_;
  assign new_E9928_ = new_E9937_ | new_E9936_;
  assign new_E9929_ = new_E9939_ & new_E9938_;
  assign new_E9930_ = new_E9939_ & new_E9940_;
  assign new_E9931_ = new_E9932_ | new_E9941_;
  assign new_E9932_ = new_E9921_ | new_E9944_;
  assign new_E9933_ = new_E9943_ | new_E9942_;
  assign new_E9934_ = new_E9948_ & new_E9947_;
  assign new_E9935_ = new_E9946_ & new_E9945_;
  assign new_E9936_ = new_E9951_ | new_E9950_;
  assign new_E9937_ = new_E9946_ & new_E9949_;
  assign new_E9938_ = new_E9921_ | new_E9954_;
  assign new_E9939_ = new_E9953_ | new_E9952_;
  assign new_E9940_ = new_E9956_ | new_E9955_;
  assign new_E9941_ = ~new_E9932_ & new_E9958_;
  assign new_E9942_ = ~new_E9934_ & new_E9946_;
  assign new_E9943_ = new_E9934_ & ~new_E9946_;
  assign new_E9944_ = new_E9920_ & ~new_E9921_;
  assign new_E9945_ = ~new_E9967_ | ~new_E9968_;
  assign new_E9946_ = new_E9960_ | new_E9962_;
  assign new_E9947_ = new_E9970_ | new_E9969_;
  assign new_E9948_ = new_E9964_ | new_E9963_;
  assign new_E9949_ = ~new_E9972_ | ~new_E9971_;
  assign new_E9950_ = ~new_E9973_ & new_E9974_;
  assign new_E9951_ = new_E9973_ & ~new_E9974_;
  assign new_E9952_ = ~new_E9920_ & new_E9921_;
  assign new_E9953_ = new_E9920_ & ~new_E9921_;
  assign new_E9954_ = ~new_E9936_ | new_E9946_;
  assign new_E9955_ = new_E9936_ & new_E9946_;
  assign new_E9956_ = ~new_E9936_ & ~new_E9946_;
  assign new_E9957_ = new_E9978_ | new_E9977_;
  assign new_E9958_ = new_E9924_ | new_E9957_;
  assign new_E9959_ = new_E9982_ | new_E9981_;
  assign new_E9960_ = ~new_E9924_ & new_E9959_;
  assign new_E9961_ = new_E9980_ | new_E9979_;
  assign new_E9962_ = new_E9924_ & new_E9961_;
  assign new_E9963_ = new_E9922_ & ~new_E9932_;
  assign new_E9964_ = ~new_E9922_ & new_E9932_;
  assign new_E9965_ = ~new_E9921_ | ~new_E9946_;
  assign new_E9966_ = new_E9932_ & new_E9965_;
  assign new_E9967_ = ~new_E9932_ & ~new_E9966_;
  assign new_E9968_ = new_E9932_ | new_E9965_;
  assign new_E9969_ = ~new_E9922_ & new_E9923_;
  assign new_E9970_ = new_E9922_ & ~new_E9923_;
  assign new_E9971_ = new_E9939_ | new_E9976_;
  assign new_E9972_ = ~new_E9939_ & ~new_E9975_;
  assign new_E9973_ = new_E9922_ | new_E9939_;
  assign new_E9974_ = new_E9922_ | new_E9923_;
  assign new_E9975_ = new_E9939_ & new_E9976_;
  assign new_E9976_ = ~new_E9921_ | ~new_E9946_;
  assign new_E9977_ = new_E9954_ & new_E9974_;
  assign new_E9978_ = ~new_E9954_ & ~new_E9974_;
  assign new_E9979_ = new_E9983_ | new_E9984_;
  assign new_E9980_ = ~new_E9925_ & new_E9939_;
  assign new_E9981_ = new_E9985_ | new_E9986_;
  assign new_E9982_ = new_E9925_ & new_E9939_;
  assign new_E9983_ = ~new_E9925_ & ~new_E9939_;
  assign new_E9984_ = new_E9925_ & ~new_E9939_;
  assign new_E9985_ = new_E9925_ & ~new_E9939_;
  assign new_E9986_ = ~new_E9925_ & new_E9939_;
  assign new_E9987_ = new_F7101_;
  assign new_E9988_ = new_F7168_;
  assign new_E9989_ = new_F7235_;
  assign new_E9990_ = new_F7302_;
  assign new_E9991_ = new_F7369_;
  assign new_E9992_ = new_F7436_;
  assign new_E9993_ = new_F1_ & new_E9999_;
  assign new_E9994_ = new_F3_ | new_F2_;
  assign new_E9995_ = new_F5_ | new_F4_;
  assign new_E9996_ = new_F7_ & new_F6_;
  assign new_E9997_ = new_F7_ & new_F8_;
  assign new_E9998_ = new_E9999_ | new_F9_;
  assign new_E9999_ = new_E9988_ | new_F12_;
  assign new_F1_ = new_F11_ | new_F10_;
  assign new_F2_ = new_F16_ & new_F15_;
  assign new_F3_ = new_F14_ & new_F13_;
  assign new_F4_ = new_F19_ | new_F18_;
  assign new_F5_ = new_F14_ & new_F17_;
  assign new_F6_ = new_E9988_ | new_F22_;
  assign new_F7_ = new_F21_ | new_F20_;
  assign new_F8_ = new_F24_ | new_F23_;
  assign new_F9_ = ~new_E9999_ & new_F26_;
  assign new_F10_ = ~new_F2_ & new_F14_;
  assign new_F11_ = new_F2_ & ~new_F14_;
  assign new_F12_ = new_E9987_ & ~new_E9988_;
  assign new_F13_ = ~new_F35_ | ~new_F36_;
  assign new_F14_ = new_F28_ | new_F30_;
  assign new_F15_ = new_F38_ | new_F37_;
  assign new_F16_ = new_F32_ | new_F31_;
  assign new_F17_ = ~new_F40_ | ~new_F39_;
  assign new_F18_ = ~new_F41_ & new_F42_;
  assign new_F19_ = new_F41_ & ~new_F42_;
  assign new_F20_ = ~new_E9987_ & new_E9988_;
  assign new_F21_ = new_E9987_ & ~new_E9988_;
  assign new_F22_ = ~new_F4_ | new_F14_;
  assign new_F23_ = new_F4_ & new_F14_;
  assign new_F24_ = ~new_F4_ & ~new_F14_;
  assign new_F25_ = new_F46_ | new_F45_;
  assign new_F26_ = new_E9991_ | new_F25_;
  assign new_F27_ = new_F50_ | new_F49_;
  assign new_F28_ = ~new_E9991_ & new_F27_;
  assign new_F29_ = new_F48_ | new_F47_;
  assign new_F30_ = new_E9991_ & new_F29_;
  assign new_F31_ = new_E9989_ & ~new_E9999_;
  assign new_F32_ = ~new_E9989_ & new_E9999_;
  assign new_F33_ = ~new_E9988_ | ~new_F14_;
  assign new_F34_ = new_E9999_ & new_F33_;
  assign new_F35_ = ~new_E9999_ & ~new_F34_;
  assign new_F36_ = new_E9999_ | new_F33_;
  assign new_F37_ = ~new_E9989_ & new_E9990_;
  assign new_F38_ = new_E9989_ & ~new_E9990_;
  assign new_F39_ = new_F7_ | new_F44_;
  assign new_F40_ = ~new_F7_ & ~new_F43_;
  assign new_F41_ = new_E9989_ | new_F7_;
  assign new_F42_ = new_E9989_ | new_E9990_;
  assign new_F43_ = new_F7_ & new_F44_;
  assign new_F44_ = ~new_E9988_ | ~new_F14_;
  assign new_F45_ = new_F22_ & new_F42_;
  assign new_F46_ = ~new_F22_ & ~new_F42_;
  assign new_F47_ = new_F51_ | new_F52_;
  assign new_F48_ = ~new_E9992_ & new_F7_;
  assign new_F49_ = new_F53_ | new_F54_;
  assign new_F50_ = new_E9992_ & new_F7_;
  assign new_F51_ = ~new_E9992_ & ~new_F7_;
  assign new_F52_ = new_E9992_ & ~new_F7_;
  assign new_F53_ = new_E9992_ & ~new_F7_;
  assign new_F54_ = ~new_E9992_ & new_F7_;
  assign new_F55_ = new_F7503_;
  assign new_F56_ = new_F7570_;
  assign new_F57_ = new_F7637_;
  assign new_F58_ = new_F7704_;
  assign new_F59_ = new_F7771_;
  assign new_F60_ = new_F7838_;
  assign new_F61_ = new_F68_ & new_F67_;
  assign new_F62_ = new_F70_ | new_F69_;
  assign new_F63_ = new_F72_ | new_F71_;
  assign new_F64_ = new_F74_ & new_F73_;
  assign new_F65_ = new_F74_ & new_F75_;
  assign new_F66_ = new_F67_ | new_F76_;
  assign new_F67_ = new_F56_ | new_F79_;
  assign new_F68_ = new_F78_ | new_F77_;
  assign new_F69_ = new_F83_ & new_F82_;
  assign new_F70_ = new_F81_ & new_F80_;
  assign new_F71_ = new_F86_ | new_F85_;
  assign new_F72_ = new_F81_ & new_F84_;
  assign new_F73_ = new_F56_ | new_F89_;
  assign new_F74_ = new_F88_ | new_F87_;
  assign new_F75_ = new_F91_ | new_F90_;
  assign new_F76_ = ~new_F67_ & new_F93_;
  assign new_F77_ = ~new_F69_ & new_F81_;
  assign new_F78_ = new_F69_ & ~new_F81_;
  assign new_F79_ = new_F55_ & ~new_F56_;
  assign new_F80_ = ~new_F102_ | ~new_F103_;
  assign new_F81_ = new_F95_ | new_F97_;
  assign new_F82_ = new_F105_ | new_F104_;
  assign new_F83_ = new_F99_ | new_F98_;
  assign new_F84_ = ~new_F107_ | ~new_F106_;
  assign new_F85_ = ~new_F108_ & new_F109_;
  assign new_F86_ = new_F108_ & ~new_F109_;
  assign new_F87_ = ~new_F55_ & new_F56_;
  assign new_F88_ = new_F55_ & ~new_F56_;
  assign new_F89_ = ~new_F71_ | new_F81_;
  assign new_F90_ = new_F71_ & new_F81_;
  assign new_F91_ = ~new_F71_ & ~new_F81_;
  assign new_F92_ = new_F113_ | new_F112_;
  assign new_F93_ = new_F59_ | new_F92_;
  assign new_F94_ = new_F117_ | new_F116_;
  assign new_F95_ = ~new_F59_ & new_F94_;
  assign new_F96_ = new_F115_ | new_F114_;
  assign new_F97_ = new_F59_ & new_F96_;
  assign new_F98_ = new_F57_ & ~new_F67_;
  assign new_F99_ = ~new_F57_ & new_F67_;
  assign new_F100_ = ~new_F56_ | ~new_F81_;
  assign new_F101_ = new_F67_ & new_F100_;
  assign new_F102_ = ~new_F67_ & ~new_F101_;
  assign new_F103_ = new_F67_ | new_F100_;
  assign new_F104_ = ~new_F57_ & new_F58_;
  assign new_F105_ = new_F57_ & ~new_F58_;
  assign new_F106_ = new_F74_ | new_F111_;
  assign new_F107_ = ~new_F74_ & ~new_F110_;
  assign new_F108_ = new_F57_ | new_F74_;
  assign new_F109_ = new_F57_ | new_F58_;
  assign new_F110_ = new_F74_ & new_F111_;
  assign new_F111_ = ~new_F56_ | ~new_F81_;
  assign new_F112_ = new_F89_ & new_F109_;
  assign new_F113_ = ~new_F89_ & ~new_F109_;
  assign new_F114_ = new_F118_ | new_F119_;
  assign new_F115_ = ~new_F60_ & new_F74_;
  assign new_F116_ = new_F120_ | new_F121_;
  assign new_F117_ = new_F60_ & new_F74_;
  assign new_F118_ = ~new_F60_ & ~new_F74_;
  assign new_F119_ = new_F60_ & ~new_F74_;
  assign new_F120_ = new_F60_ & ~new_F74_;
  assign new_F121_ = ~new_F60_ & new_F74_;
  assign new_F122_ = new_F7905_;
  assign new_F123_ = new_F7972_;
  assign new_F124_ = new_F8039_;
  assign new_F125_ = new_F8106_;
  assign new_F126_ = new_F8173_;
  assign new_F127_ = new_F8240_;
  assign new_F128_ = new_F135_ & new_F134_;
  assign new_F129_ = new_F137_ | new_F136_;
  assign new_F130_ = new_F139_ | new_F138_;
  assign new_F131_ = new_F141_ & new_F140_;
  assign new_F132_ = new_F141_ & new_F142_;
  assign new_F133_ = new_F134_ | new_F143_;
  assign new_F134_ = new_F123_ | new_F146_;
  assign new_F135_ = new_F145_ | new_F144_;
  assign new_F136_ = new_F150_ & new_F149_;
  assign new_F137_ = new_F148_ & new_F147_;
  assign new_F138_ = new_F153_ | new_F152_;
  assign new_F139_ = new_F148_ & new_F151_;
  assign new_F140_ = new_F123_ | new_F156_;
  assign new_F141_ = new_F155_ | new_F154_;
  assign new_F142_ = new_F158_ | new_F157_;
  assign new_F143_ = ~new_F134_ & new_F160_;
  assign new_F144_ = ~new_F136_ & new_F148_;
  assign new_F145_ = new_F136_ & ~new_F148_;
  assign new_F146_ = new_F122_ & ~new_F123_;
  assign new_F147_ = ~new_F169_ | ~new_F170_;
  assign new_F148_ = new_F162_ | new_F164_;
  assign new_F149_ = new_F172_ | new_F171_;
  assign new_F150_ = new_F166_ | new_F165_;
  assign new_F151_ = ~new_F174_ | ~new_F173_;
  assign new_F152_ = ~new_F175_ & new_F176_;
  assign new_F153_ = new_F175_ & ~new_F176_;
  assign new_F154_ = ~new_F122_ & new_F123_;
  assign new_F155_ = new_F122_ & ~new_F123_;
  assign new_F156_ = ~new_F138_ | new_F148_;
  assign new_F157_ = new_F138_ & new_F148_;
  assign new_F158_ = ~new_F138_ & ~new_F148_;
  assign new_F159_ = new_F180_ | new_F179_;
  assign new_F160_ = new_F126_ | new_F159_;
  assign new_F161_ = new_F184_ | new_F183_;
  assign new_F162_ = ~new_F126_ & new_F161_;
  assign new_F163_ = new_F182_ | new_F181_;
  assign new_F164_ = new_F126_ & new_F163_;
  assign new_F165_ = new_F124_ & ~new_F134_;
  assign new_F166_ = ~new_F124_ & new_F134_;
  assign new_F167_ = ~new_F123_ | ~new_F148_;
  assign new_F168_ = new_F134_ & new_F167_;
  assign new_F169_ = ~new_F134_ & ~new_F168_;
  assign new_F170_ = new_F134_ | new_F167_;
  assign new_F171_ = ~new_F124_ & new_F125_;
  assign new_F172_ = new_F124_ & ~new_F125_;
  assign new_F173_ = new_F141_ | new_F178_;
  assign new_F174_ = ~new_F141_ & ~new_F177_;
  assign new_F175_ = new_F124_ | new_F141_;
  assign new_F176_ = new_F124_ | new_F125_;
  assign new_F177_ = new_F141_ & new_F178_;
  assign new_F178_ = ~new_F123_ | ~new_F148_;
  assign new_F179_ = new_F156_ & new_F176_;
  assign new_F180_ = ~new_F156_ & ~new_F176_;
  assign new_F181_ = new_F185_ | new_F186_;
  assign new_F182_ = ~new_F127_ & new_F141_;
  assign new_F183_ = new_F187_ | new_F188_;
  assign new_F184_ = new_F127_ & new_F141_;
  assign new_F185_ = ~new_F127_ & ~new_F141_;
  assign new_F186_ = new_F127_ & ~new_F141_;
  assign new_F187_ = new_F127_ & ~new_F141_;
  assign new_F188_ = ~new_F127_ & new_F141_;
  assign new_F189_ = new_F8307_;
  assign new_F190_ = new_F8374_;
  assign new_F191_ = new_F8441_;
  assign new_F192_ = new_F8508_;
  assign new_F193_ = new_F8575_;
  assign new_F194_ = new_F8642_;
  assign new_F195_ = new_F202_ & new_F201_;
  assign new_F196_ = new_F204_ | new_F203_;
  assign new_F197_ = new_F206_ | new_F205_;
  assign new_F198_ = new_F208_ & new_F207_;
  assign new_F199_ = new_F208_ & new_F209_;
  assign new_F200_ = new_F201_ | new_F210_;
  assign new_F201_ = new_F190_ | new_F213_;
  assign new_F202_ = new_F212_ | new_F211_;
  assign new_F203_ = new_F217_ & new_F216_;
  assign new_F204_ = new_F215_ & new_F214_;
  assign new_F205_ = new_F220_ | new_F219_;
  assign new_F206_ = new_F215_ & new_F218_;
  assign new_F207_ = new_F190_ | new_F223_;
  assign new_F208_ = new_F222_ | new_F221_;
  assign new_F209_ = new_F225_ | new_F224_;
  assign new_F210_ = ~new_F201_ & new_F227_;
  assign new_F211_ = ~new_F203_ & new_F215_;
  assign new_F212_ = new_F203_ & ~new_F215_;
  assign new_F213_ = new_F189_ & ~new_F190_;
  assign new_F214_ = ~new_F236_ | ~new_F237_;
  assign new_F215_ = new_F229_ | new_F231_;
  assign new_F216_ = new_F239_ | new_F238_;
  assign new_F217_ = new_F233_ | new_F232_;
  assign new_F218_ = ~new_F241_ | ~new_F240_;
  assign new_F219_ = ~new_F242_ & new_F243_;
  assign new_F220_ = new_F242_ & ~new_F243_;
  assign new_F221_ = ~new_F189_ & new_F190_;
  assign new_F222_ = new_F189_ & ~new_F190_;
  assign new_F223_ = ~new_F205_ | new_F215_;
  assign new_F224_ = new_F205_ & new_F215_;
  assign new_F225_ = ~new_F205_ & ~new_F215_;
  assign new_F226_ = new_F247_ | new_F246_;
  assign new_F227_ = new_F193_ | new_F226_;
  assign new_F228_ = new_F251_ | new_F250_;
  assign new_F229_ = ~new_F193_ & new_F228_;
  assign new_F230_ = new_F249_ | new_F248_;
  assign new_F231_ = new_F193_ & new_F230_;
  assign new_F232_ = new_F191_ & ~new_F201_;
  assign new_F233_ = ~new_F191_ & new_F201_;
  assign new_F234_ = ~new_F190_ | ~new_F215_;
  assign new_F235_ = new_F201_ & new_F234_;
  assign new_F236_ = ~new_F201_ & ~new_F235_;
  assign new_F237_ = new_F201_ | new_F234_;
  assign new_F238_ = ~new_F191_ & new_F192_;
  assign new_F239_ = new_F191_ & ~new_F192_;
  assign new_F240_ = new_F208_ | new_F245_;
  assign new_F241_ = ~new_F208_ & ~new_F244_;
  assign new_F242_ = new_F191_ | new_F208_;
  assign new_F243_ = new_F191_ | new_F192_;
  assign new_F244_ = new_F208_ & new_F245_;
  assign new_F245_ = ~new_F190_ | ~new_F215_;
  assign new_F246_ = new_F223_ & new_F243_;
  assign new_F247_ = ~new_F223_ & ~new_F243_;
  assign new_F248_ = new_F252_ | new_F253_;
  assign new_F249_ = ~new_F194_ & new_F208_;
  assign new_F250_ = new_F254_ | new_F255_;
  assign new_F251_ = new_F194_ & new_F208_;
  assign new_F252_ = ~new_F194_ & ~new_F208_;
  assign new_F253_ = new_F194_ & ~new_F208_;
  assign new_F254_ = new_F194_ & ~new_F208_;
  assign new_F255_ = ~new_F194_ & new_F208_;
  assign new_F256_ = new_F8709_;
  assign new_F257_ = new_F8776_;
  assign new_F258_ = new_F8843_;
  assign new_F259_ = new_F8910_;
  assign new_F260_ = new_F8977_;
  assign new_F261_ = new_F9044_;
  assign new_F262_ = new_F269_ & new_F268_;
  assign new_F263_ = new_F271_ | new_F270_;
  assign new_F264_ = new_F273_ | new_F272_;
  assign new_F265_ = new_F275_ & new_F274_;
  assign new_F266_ = new_F275_ & new_F276_;
  assign new_F267_ = new_F268_ | new_F277_;
  assign new_F268_ = new_F257_ | new_F280_;
  assign new_F269_ = new_F279_ | new_F278_;
  assign new_F270_ = new_F284_ & new_F283_;
  assign new_F271_ = new_F282_ & new_F281_;
  assign new_F272_ = new_F287_ | new_F286_;
  assign new_F273_ = new_F282_ & new_F285_;
  assign new_F274_ = new_F257_ | new_F290_;
  assign new_F275_ = new_F289_ | new_F288_;
  assign new_F276_ = new_F292_ | new_F291_;
  assign new_F277_ = ~new_F268_ & new_F294_;
  assign new_F278_ = ~new_F270_ & new_F282_;
  assign new_F279_ = new_F270_ & ~new_F282_;
  assign new_F280_ = new_F256_ & ~new_F257_;
  assign new_F281_ = ~new_F303_ | ~new_F304_;
  assign new_F282_ = new_F296_ | new_F298_;
  assign new_F283_ = new_F306_ | new_F305_;
  assign new_F284_ = new_F300_ | new_F299_;
  assign new_F285_ = ~new_F308_ | ~new_F307_;
  assign new_F286_ = ~new_F309_ & new_F310_;
  assign new_F287_ = new_F309_ & ~new_F310_;
  assign new_F288_ = ~new_F256_ & new_F257_;
  assign new_F289_ = new_F256_ & ~new_F257_;
  assign new_F290_ = ~new_F272_ | new_F282_;
  assign new_F291_ = new_F272_ & new_F282_;
  assign new_F292_ = ~new_F272_ & ~new_F282_;
  assign new_F293_ = new_F314_ | new_F313_;
  assign new_F294_ = new_F260_ | new_F293_;
  assign new_F295_ = new_F318_ | new_F317_;
  assign new_F296_ = ~new_F260_ & new_F295_;
  assign new_F297_ = new_F316_ | new_F315_;
  assign new_F298_ = new_F260_ & new_F297_;
  assign new_F299_ = new_F258_ & ~new_F268_;
  assign new_F300_ = ~new_F258_ & new_F268_;
  assign new_F301_ = ~new_F257_ | ~new_F282_;
  assign new_F302_ = new_F268_ & new_F301_;
  assign new_F303_ = ~new_F268_ & ~new_F302_;
  assign new_F304_ = new_F268_ | new_F301_;
  assign new_F305_ = ~new_F258_ & new_F259_;
  assign new_F306_ = new_F258_ & ~new_F259_;
  assign new_F307_ = new_F275_ | new_F312_;
  assign new_F308_ = ~new_F275_ & ~new_F311_;
  assign new_F309_ = new_F258_ | new_F275_;
  assign new_F310_ = new_F258_ | new_F259_;
  assign new_F311_ = new_F275_ & new_F312_;
  assign new_F312_ = ~new_F257_ | ~new_F282_;
  assign new_F313_ = new_F290_ & new_F310_;
  assign new_F314_ = ~new_F290_ & ~new_F310_;
  assign new_F315_ = new_F319_ | new_F320_;
  assign new_F316_ = ~new_F261_ & new_F275_;
  assign new_F317_ = new_F321_ | new_F322_;
  assign new_F318_ = new_F261_ & new_F275_;
  assign new_F319_ = ~new_F261_ & ~new_F275_;
  assign new_F320_ = new_F261_ & ~new_F275_;
  assign new_F321_ = new_F261_ & ~new_F275_;
  assign new_F322_ = ~new_F261_ & new_F275_;
  assign new_F323_ = new_F9111_;
  assign new_F324_ = new_F9178_;
  assign new_F325_ = new_F9245_;
  assign new_F326_ = new_F9312_;
  assign new_F327_ = new_F9379_;
  assign new_F328_ = new_F9446_;
  assign new_F329_ = new_F336_ & new_F335_;
  assign new_F330_ = new_F338_ | new_F337_;
  assign new_F331_ = new_F340_ | new_F339_;
  assign new_F332_ = new_F342_ & new_F341_;
  assign new_F333_ = new_F342_ & new_F343_;
  assign new_F334_ = new_F335_ | new_F344_;
  assign new_F335_ = new_F324_ | new_F347_;
  assign new_F336_ = new_F346_ | new_F345_;
  assign new_F337_ = new_F351_ & new_F350_;
  assign new_F338_ = new_F349_ & new_F348_;
  assign new_F339_ = new_F354_ | new_F353_;
  assign new_F340_ = new_F349_ & new_F352_;
  assign new_F341_ = new_F324_ | new_F357_;
  assign new_F342_ = new_F356_ | new_F355_;
  assign new_F343_ = new_F359_ | new_F358_;
  assign new_F344_ = ~new_F335_ & new_F361_;
  assign new_F345_ = ~new_F337_ & new_F349_;
  assign new_F346_ = new_F337_ & ~new_F349_;
  assign new_F347_ = new_F323_ & ~new_F324_;
  assign new_F348_ = ~new_F370_ | ~new_F371_;
  assign new_F349_ = new_F363_ | new_F365_;
  assign new_F350_ = new_F373_ | new_F372_;
  assign new_F351_ = new_F367_ | new_F366_;
  assign new_F352_ = ~new_F375_ | ~new_F374_;
  assign new_F353_ = ~new_F376_ & new_F377_;
  assign new_F354_ = new_F376_ & ~new_F377_;
  assign new_F355_ = ~new_F323_ & new_F324_;
  assign new_F356_ = new_F323_ & ~new_F324_;
  assign new_F357_ = ~new_F339_ | new_F349_;
  assign new_F358_ = new_F339_ & new_F349_;
  assign new_F359_ = ~new_F339_ & ~new_F349_;
  assign new_F360_ = new_F381_ | new_F380_;
  assign new_F361_ = new_F327_ | new_F360_;
  assign new_F362_ = new_F385_ | new_F384_;
  assign new_F363_ = ~new_F327_ & new_F362_;
  assign new_F364_ = new_F383_ | new_F382_;
  assign new_F365_ = new_F327_ & new_F364_;
  assign new_F366_ = new_F325_ & ~new_F335_;
  assign new_F367_ = ~new_F325_ & new_F335_;
  assign new_F368_ = ~new_F324_ | ~new_F349_;
  assign new_F369_ = new_F335_ & new_F368_;
  assign new_F370_ = ~new_F335_ & ~new_F369_;
  assign new_F371_ = new_F335_ | new_F368_;
  assign new_F372_ = ~new_F325_ & new_F326_;
  assign new_F373_ = new_F325_ & ~new_F326_;
  assign new_F374_ = new_F342_ | new_F379_;
  assign new_F375_ = ~new_F342_ & ~new_F378_;
  assign new_F376_ = new_F325_ | new_F342_;
  assign new_F377_ = new_F325_ | new_F326_;
  assign new_F378_ = new_F342_ & new_F379_;
  assign new_F379_ = ~new_F324_ | ~new_F349_;
  assign new_F380_ = new_F357_ & new_F377_;
  assign new_F381_ = ~new_F357_ & ~new_F377_;
  assign new_F382_ = new_F386_ | new_F387_;
  assign new_F383_ = ~new_F328_ & new_F342_;
  assign new_F384_ = new_F388_ | new_F389_;
  assign new_F385_ = new_F328_ & new_F342_;
  assign new_F386_ = ~new_F328_ & ~new_F342_;
  assign new_F387_ = new_F328_ & ~new_F342_;
  assign new_F388_ = new_F328_ & ~new_F342_;
  assign new_F389_ = ~new_F328_ & new_F342_;
  assign new_F390_ = new_F9513_;
  assign new_F391_ = new_F9580_;
  assign new_F392_ = new_F9647_;
  assign new_F393_ = new_F9714_;
  assign new_F394_ = new_F9781_;
  assign new_F395_ = new_F9848_;
  assign new_F396_ = new_F403_ & new_F402_;
  assign new_F397_ = new_F405_ | new_F404_;
  assign new_F398_ = new_F407_ | new_F406_;
  assign new_F399_ = new_F409_ & new_F408_;
  assign new_F400_ = new_F409_ & new_F410_;
  assign new_F401_ = new_F402_ | new_F411_;
  assign new_F402_ = new_F391_ | new_F414_;
  assign new_F403_ = new_F413_ | new_F412_;
  assign new_F404_ = new_F418_ & new_F417_;
  assign new_F405_ = new_F416_ & new_F415_;
  assign new_F406_ = new_F421_ | new_F420_;
  assign new_F407_ = new_F416_ & new_F419_;
  assign new_F408_ = new_F391_ | new_F424_;
  assign new_F409_ = new_F423_ | new_F422_;
  assign new_F410_ = new_F426_ | new_F425_;
  assign new_F411_ = ~new_F402_ & new_F428_;
  assign new_F412_ = ~new_F404_ & new_F416_;
  assign new_F413_ = new_F404_ & ~new_F416_;
  assign new_F414_ = new_F390_ & ~new_F391_;
  assign new_F415_ = ~new_F437_ | ~new_F438_;
  assign new_F416_ = new_F430_ | new_F432_;
  assign new_F417_ = new_F440_ | new_F439_;
  assign new_F418_ = new_F434_ | new_F433_;
  assign new_F419_ = ~new_F442_ | ~new_F441_;
  assign new_F420_ = ~new_F443_ & new_F444_;
  assign new_F421_ = new_F443_ & ~new_F444_;
  assign new_F422_ = ~new_F390_ & new_F391_;
  assign new_F423_ = new_F390_ & ~new_F391_;
  assign new_F424_ = ~new_F406_ | new_F416_;
  assign new_F425_ = new_F406_ & new_F416_;
  assign new_F426_ = ~new_F406_ & ~new_F416_;
  assign new_F427_ = new_F448_ | new_F447_;
  assign new_F428_ = new_F394_ | new_F427_;
  assign new_F429_ = new_F452_ | new_F451_;
  assign new_F430_ = ~new_F394_ & new_F429_;
  assign new_F431_ = new_F450_ | new_F449_;
  assign new_F432_ = new_F394_ & new_F431_;
  assign new_F433_ = new_F392_ & ~new_F402_;
  assign new_F434_ = ~new_F392_ & new_F402_;
  assign new_F435_ = ~new_F391_ | ~new_F416_;
  assign new_F436_ = new_F402_ & new_F435_;
  assign new_F437_ = ~new_F402_ & ~new_F436_;
  assign new_F438_ = new_F402_ | new_F435_;
  assign new_F439_ = ~new_F392_ & new_F393_;
  assign new_F440_ = new_F392_ & ~new_F393_;
  assign new_F441_ = new_F409_ | new_F446_;
  assign new_F442_ = ~new_F409_ & ~new_F445_;
  assign new_F443_ = new_F392_ | new_F409_;
  assign new_F444_ = new_F392_ | new_F393_;
  assign new_F445_ = new_F409_ & new_F446_;
  assign new_F446_ = ~new_F391_ | ~new_F416_;
  assign new_F447_ = new_F424_ & new_F444_;
  assign new_F448_ = ~new_F424_ & ~new_F444_;
  assign new_F449_ = new_F453_ | new_F454_;
  assign new_F450_ = ~new_F395_ & new_F409_;
  assign new_F451_ = new_F455_ | new_F456_;
  assign new_F452_ = new_F395_ & new_F409_;
  assign new_F453_ = ~new_F395_ & ~new_F409_;
  assign new_F454_ = new_F395_ & ~new_F409_;
  assign new_F455_ = new_F395_ & ~new_F409_;
  assign new_F456_ = ~new_F395_ & new_F409_;
  assign new_F457_ = new_F9915_;
  assign new_F458_ = new_F9982_;
  assign new_F459_ = new_G50_;
  assign new_F460_ = new_G117_;
  assign new_F461_ = new_G184_;
  assign new_F462_ = new_G251_;
  assign new_F463_ = new_F470_ & new_F469_;
  assign new_F464_ = new_F472_ | new_F471_;
  assign new_F465_ = new_F474_ | new_F473_;
  assign new_F466_ = new_F476_ & new_F475_;
  assign new_F467_ = new_F476_ & new_F477_;
  assign new_F468_ = new_F469_ | new_F478_;
  assign new_F469_ = new_F458_ | new_F481_;
  assign new_F470_ = new_F480_ | new_F479_;
  assign new_F471_ = new_F485_ & new_F484_;
  assign new_F472_ = new_F483_ & new_F482_;
  assign new_F473_ = new_F488_ | new_F487_;
  assign new_F474_ = new_F483_ & new_F486_;
  assign new_F475_ = new_F458_ | new_F491_;
  assign new_F476_ = new_F490_ | new_F489_;
  assign new_F477_ = new_F493_ | new_F492_;
  assign new_F478_ = ~new_F469_ & new_F495_;
  assign new_F479_ = ~new_F471_ & new_F483_;
  assign new_F480_ = new_F471_ & ~new_F483_;
  assign new_F481_ = new_F457_ & ~new_F458_;
  assign new_F482_ = ~new_F504_ | ~new_F505_;
  assign new_F483_ = new_F497_ | new_F499_;
  assign new_F484_ = new_F507_ | new_F506_;
  assign new_F485_ = new_F501_ | new_F500_;
  assign new_F486_ = ~new_F509_ | ~new_F508_;
  assign new_F487_ = ~new_F510_ & new_F511_;
  assign new_F488_ = new_F510_ & ~new_F511_;
  assign new_F489_ = ~new_F457_ & new_F458_;
  assign new_F490_ = new_F457_ & ~new_F458_;
  assign new_F491_ = ~new_F473_ | new_F483_;
  assign new_F492_ = new_F473_ & new_F483_;
  assign new_F493_ = ~new_F473_ & ~new_F483_;
  assign new_F494_ = new_F515_ | new_F514_;
  assign new_F495_ = new_F461_ | new_F494_;
  assign new_F496_ = new_F519_ | new_F518_;
  assign new_F497_ = ~new_F461_ & new_F496_;
  assign new_F498_ = new_F517_ | new_F516_;
  assign new_F499_ = new_F461_ & new_F498_;
  assign new_F500_ = new_F459_ & ~new_F469_;
  assign new_F501_ = ~new_F459_ & new_F469_;
  assign new_F502_ = ~new_F458_ | ~new_F483_;
  assign new_F503_ = new_F469_ & new_F502_;
  assign new_F504_ = ~new_F469_ & ~new_F503_;
  assign new_F505_ = new_F469_ | new_F502_;
  assign new_F506_ = ~new_F459_ & new_F460_;
  assign new_F507_ = new_F459_ & ~new_F460_;
  assign new_F508_ = new_F476_ | new_F513_;
  assign new_F509_ = ~new_F476_ & ~new_F512_;
  assign new_F510_ = new_F459_ | new_F476_;
  assign new_F511_ = new_F459_ | new_F460_;
  assign new_F512_ = new_F476_ & new_F513_;
  assign new_F513_ = ~new_F458_ | ~new_F483_;
  assign new_F514_ = new_F491_ & new_F511_;
  assign new_F515_ = ~new_F491_ & ~new_F511_;
  assign new_F516_ = new_F520_ | new_F521_;
  assign new_F517_ = ~new_F462_ & new_F476_;
  assign new_F518_ = new_F522_ | new_F523_;
  assign new_F519_ = new_F462_ & new_F476_;
  assign new_F520_ = ~new_F462_ & ~new_F476_;
  assign new_F521_ = new_F462_ & ~new_F476_;
  assign new_F522_ = new_F462_ & ~new_F476_;
  assign new_F523_ = ~new_F462_ & new_F476_;
  assign new_F524_ = new_G318_;
  assign new_F525_ = new_G385_;
  assign new_F526_ = new_G452_;
  assign new_F527_ = new_G519_;
  assign new_F528_ = new_G586_;
  assign new_F529_ = new_G653_;
  assign new_F530_ = new_F537_ & new_F536_;
  assign new_F531_ = new_F539_ | new_F538_;
  assign new_F532_ = new_F541_ | new_F540_;
  assign new_F533_ = new_F543_ & new_F542_;
  assign new_F534_ = new_F543_ & new_F544_;
  assign new_F535_ = new_F536_ | new_F545_;
  assign new_F536_ = new_F525_ | new_F548_;
  assign new_F537_ = new_F547_ | new_F546_;
  assign new_F538_ = new_F552_ & new_F551_;
  assign new_F539_ = new_F550_ & new_F549_;
  assign new_F540_ = new_F555_ | new_F554_;
  assign new_F541_ = new_F550_ & new_F553_;
  assign new_F542_ = new_F525_ | new_F558_;
  assign new_F543_ = new_F557_ | new_F556_;
  assign new_F544_ = new_F560_ | new_F559_;
  assign new_F545_ = ~new_F536_ & new_F562_;
  assign new_F546_ = ~new_F538_ & new_F550_;
  assign new_F547_ = new_F538_ & ~new_F550_;
  assign new_F548_ = new_F524_ & ~new_F525_;
  assign new_F549_ = ~new_F571_ | ~new_F572_;
  assign new_F550_ = new_F564_ | new_F566_;
  assign new_F551_ = new_F574_ | new_F573_;
  assign new_F552_ = new_F568_ | new_F567_;
  assign new_F553_ = ~new_F576_ | ~new_F575_;
  assign new_F554_ = ~new_F577_ & new_F578_;
  assign new_F555_ = new_F577_ & ~new_F578_;
  assign new_F556_ = ~new_F524_ & new_F525_;
  assign new_F557_ = new_F524_ & ~new_F525_;
  assign new_F558_ = ~new_F540_ | new_F550_;
  assign new_F559_ = new_F540_ & new_F550_;
  assign new_F560_ = ~new_F540_ & ~new_F550_;
  assign new_F561_ = new_F582_ | new_F581_;
  assign new_F562_ = new_F528_ | new_F561_;
  assign new_F563_ = new_F586_ | new_F585_;
  assign new_F564_ = ~new_F528_ & new_F563_;
  assign new_F565_ = new_F584_ | new_F583_;
  assign new_F566_ = new_F528_ & new_F565_;
  assign new_F567_ = new_F526_ & ~new_F536_;
  assign new_F568_ = ~new_F526_ & new_F536_;
  assign new_F569_ = ~new_F525_ | ~new_F550_;
  assign new_F570_ = new_F536_ & new_F569_;
  assign new_F571_ = ~new_F536_ & ~new_F570_;
  assign new_F572_ = new_F536_ | new_F569_;
  assign new_F573_ = ~new_F526_ & new_F527_;
  assign new_F574_ = new_F526_ & ~new_F527_;
  assign new_F575_ = new_F543_ | new_F580_;
  assign new_F576_ = ~new_F543_ & ~new_F579_;
  assign new_F577_ = new_F526_ | new_F543_;
  assign new_F578_ = new_F526_ | new_F527_;
  assign new_F579_ = new_F543_ & new_F580_;
  assign new_F580_ = ~new_F525_ | ~new_F550_;
  assign new_F581_ = new_F558_ & new_F578_;
  assign new_F582_ = ~new_F558_ & ~new_F578_;
  assign new_F583_ = new_F587_ | new_F588_;
  assign new_F584_ = ~new_F529_ & new_F543_;
  assign new_F585_ = new_F589_ | new_F590_;
  assign new_F586_ = new_F529_ & new_F543_;
  assign new_F587_ = ~new_F529_ & ~new_F543_;
  assign new_F588_ = new_F529_ & ~new_F543_;
  assign new_F589_ = new_F529_ & ~new_F543_;
  assign new_F590_ = ~new_F529_ & new_F543_;
  assign new_F591_ = new_G720_;
  assign new_F592_ = new_G787_;
  assign new_F593_ = new_G854_;
  assign new_F594_ = new_G921_;
  assign new_F595_ = new_G988_;
  assign new_F596_ = new_G1055_;
  assign new_F597_ = new_F604_ & new_F603_;
  assign new_F598_ = new_F606_ | new_F605_;
  assign new_F599_ = new_F608_ | new_F607_;
  assign new_F600_ = new_F610_ & new_F609_;
  assign new_F601_ = new_F610_ & new_F611_;
  assign new_F602_ = new_F603_ | new_F612_;
  assign new_F603_ = new_F592_ | new_F615_;
  assign new_F604_ = new_F614_ | new_F613_;
  assign new_F605_ = new_F619_ & new_F618_;
  assign new_F606_ = new_F617_ & new_F616_;
  assign new_F607_ = new_F622_ | new_F621_;
  assign new_F608_ = new_F617_ & new_F620_;
  assign new_F609_ = new_F592_ | new_F625_;
  assign new_F610_ = new_F624_ | new_F623_;
  assign new_F611_ = new_F627_ | new_F626_;
  assign new_F612_ = ~new_F603_ & new_F629_;
  assign new_F613_ = ~new_F605_ & new_F617_;
  assign new_F614_ = new_F605_ & ~new_F617_;
  assign new_F615_ = new_F591_ & ~new_F592_;
  assign new_F616_ = ~new_F638_ | ~new_F639_;
  assign new_F617_ = new_F631_ | new_F633_;
  assign new_F618_ = new_F641_ | new_F640_;
  assign new_F619_ = new_F635_ | new_F634_;
  assign new_F620_ = ~new_F643_ | ~new_F642_;
  assign new_F621_ = ~new_F644_ & new_F645_;
  assign new_F622_ = new_F644_ & ~new_F645_;
  assign new_F623_ = ~new_F591_ & new_F592_;
  assign new_F624_ = new_F591_ & ~new_F592_;
  assign new_F625_ = ~new_F607_ | new_F617_;
  assign new_F626_ = new_F607_ & new_F617_;
  assign new_F627_ = ~new_F607_ & ~new_F617_;
  assign new_F628_ = new_F649_ | new_F648_;
  assign new_F629_ = new_F595_ | new_F628_;
  assign new_F630_ = new_F653_ | new_F652_;
  assign new_F631_ = ~new_F595_ & new_F630_;
  assign new_F632_ = new_F651_ | new_F650_;
  assign new_F633_ = new_F595_ & new_F632_;
  assign new_F634_ = new_F593_ & ~new_F603_;
  assign new_F635_ = ~new_F593_ & new_F603_;
  assign new_F636_ = ~new_F592_ | ~new_F617_;
  assign new_F637_ = new_F603_ & new_F636_;
  assign new_F638_ = ~new_F603_ & ~new_F637_;
  assign new_F639_ = new_F603_ | new_F636_;
  assign new_F640_ = ~new_F593_ & new_F594_;
  assign new_F641_ = new_F593_ & ~new_F594_;
  assign new_F642_ = new_F610_ | new_F647_;
  assign new_F643_ = ~new_F610_ & ~new_F646_;
  assign new_F644_ = new_F593_ | new_F610_;
  assign new_F645_ = new_F593_ | new_F594_;
  assign new_F646_ = new_F610_ & new_F647_;
  assign new_F647_ = ~new_F592_ | ~new_F617_;
  assign new_F648_ = new_F625_ & new_F645_;
  assign new_F649_ = ~new_F625_ & ~new_F645_;
  assign new_F650_ = new_F654_ | new_F655_;
  assign new_F651_ = ~new_F596_ & new_F610_;
  assign new_F652_ = new_F656_ | new_F657_;
  assign new_F653_ = new_F596_ & new_F610_;
  assign new_F654_ = ~new_F596_ & ~new_F610_;
  assign new_F655_ = new_F596_ & ~new_F610_;
  assign new_F656_ = new_F596_ & ~new_F610_;
  assign new_F657_ = ~new_F596_ & new_F610_;
  assign new_F658_ = new_G1122_;
  assign new_F659_ = new_G1189_;
  assign new_F660_ = new_G1256_;
  assign new_F661_ = new_G1323_;
  assign new_F662_ = new_G1390_;
  assign new_F663_ = new_G1457_;
  assign new_F664_ = new_F671_ & new_F670_;
  assign new_F665_ = new_F673_ | new_F672_;
  assign new_F666_ = new_F675_ | new_F674_;
  assign new_F667_ = new_F677_ & new_F676_;
  assign new_F668_ = new_F677_ & new_F678_;
  assign new_F669_ = new_F670_ | new_F679_;
  assign new_F670_ = new_F659_ | new_F682_;
  assign new_F671_ = new_F681_ | new_F680_;
  assign new_F672_ = new_F686_ & new_F685_;
  assign new_F673_ = new_F684_ & new_F683_;
  assign new_F674_ = new_F689_ | new_F688_;
  assign new_F675_ = new_F684_ & new_F687_;
  assign new_F676_ = new_F659_ | new_F692_;
  assign new_F677_ = new_F691_ | new_F690_;
  assign new_F678_ = new_F694_ | new_F693_;
  assign new_F679_ = ~new_F670_ & new_F696_;
  assign new_F680_ = ~new_F672_ & new_F684_;
  assign new_F681_ = new_F672_ & ~new_F684_;
  assign new_F682_ = new_F658_ & ~new_F659_;
  assign new_F683_ = ~new_F705_ | ~new_F706_;
  assign new_F684_ = new_F698_ | new_F700_;
  assign new_F685_ = new_F708_ | new_F707_;
  assign new_F686_ = new_F702_ | new_F701_;
  assign new_F687_ = ~new_F710_ | ~new_F709_;
  assign new_F688_ = ~new_F711_ & new_F712_;
  assign new_F689_ = new_F711_ & ~new_F712_;
  assign new_F690_ = ~new_F658_ & new_F659_;
  assign new_F691_ = new_F658_ & ~new_F659_;
  assign new_F692_ = ~new_F674_ | new_F684_;
  assign new_F693_ = new_F674_ & new_F684_;
  assign new_F694_ = ~new_F674_ & ~new_F684_;
  assign new_F695_ = new_F716_ | new_F715_;
  assign new_F696_ = new_F662_ | new_F695_;
  assign new_F697_ = new_F720_ | new_F719_;
  assign new_F698_ = ~new_F662_ & new_F697_;
  assign new_F699_ = new_F718_ | new_F717_;
  assign new_F700_ = new_F662_ & new_F699_;
  assign new_F701_ = new_F660_ & ~new_F670_;
  assign new_F702_ = ~new_F660_ & new_F670_;
  assign new_F703_ = ~new_F659_ | ~new_F684_;
  assign new_F704_ = new_F670_ & new_F703_;
  assign new_F705_ = ~new_F670_ & ~new_F704_;
  assign new_F706_ = new_F670_ | new_F703_;
  assign new_F707_ = ~new_F660_ & new_F661_;
  assign new_F708_ = new_F660_ & ~new_F661_;
  assign new_F709_ = new_F677_ | new_F714_;
  assign new_F710_ = ~new_F677_ & ~new_F713_;
  assign new_F711_ = new_F660_ | new_F677_;
  assign new_F712_ = new_F660_ | new_F661_;
  assign new_F713_ = new_F677_ & new_F714_;
  assign new_F714_ = ~new_F659_ | ~new_F684_;
  assign new_F715_ = new_F692_ & new_F712_;
  assign new_F716_ = ~new_F692_ & ~new_F712_;
  assign new_F717_ = new_F721_ | new_F722_;
  assign new_F718_ = ~new_F663_ & new_F677_;
  assign new_F719_ = new_F723_ | new_F724_;
  assign new_F720_ = new_F663_ & new_F677_;
  assign new_F721_ = ~new_F663_ & ~new_F677_;
  assign new_F722_ = new_F663_ & ~new_F677_;
  assign new_F723_ = new_F663_ & ~new_F677_;
  assign new_F724_ = ~new_F663_ & new_F677_;
  assign new_F725_ = new_G1524_;
  assign new_F726_ = new_G1591_;
  assign new_F727_ = new_G1658_;
  assign new_F728_ = new_G1725_;
  assign new_F729_ = new_G1792_;
  assign new_F730_ = new_G1859_;
  assign new_F731_ = new_F738_ & new_F737_;
  assign new_F732_ = new_F740_ | new_F739_;
  assign new_F733_ = new_F742_ | new_F741_;
  assign new_F734_ = new_F744_ & new_F743_;
  assign new_F735_ = new_F744_ & new_F745_;
  assign new_F736_ = new_F737_ | new_F746_;
  assign new_F737_ = new_F726_ | new_F749_;
  assign new_F738_ = new_F748_ | new_F747_;
  assign new_F739_ = new_F753_ & new_F752_;
  assign new_F740_ = new_F751_ & new_F750_;
  assign new_F741_ = new_F756_ | new_F755_;
  assign new_F742_ = new_F751_ & new_F754_;
  assign new_F743_ = new_F726_ | new_F759_;
  assign new_F744_ = new_F758_ | new_F757_;
  assign new_F745_ = new_F761_ | new_F760_;
  assign new_F746_ = ~new_F737_ & new_F763_;
  assign new_F747_ = ~new_F739_ & new_F751_;
  assign new_F748_ = new_F739_ & ~new_F751_;
  assign new_F749_ = new_F725_ & ~new_F726_;
  assign new_F750_ = ~new_F772_ | ~new_F773_;
  assign new_F751_ = new_F765_ | new_F767_;
  assign new_F752_ = new_F775_ | new_F774_;
  assign new_F753_ = new_F769_ | new_F768_;
  assign new_F754_ = ~new_F777_ | ~new_F776_;
  assign new_F755_ = ~new_F778_ & new_F779_;
  assign new_F756_ = new_F778_ & ~new_F779_;
  assign new_F757_ = ~new_F725_ & new_F726_;
  assign new_F758_ = new_F725_ & ~new_F726_;
  assign new_F759_ = ~new_F741_ | new_F751_;
  assign new_F760_ = new_F741_ & new_F751_;
  assign new_F761_ = ~new_F741_ & ~new_F751_;
  assign new_F762_ = new_F783_ | new_F782_;
  assign new_F763_ = new_F729_ | new_F762_;
  assign new_F764_ = new_F787_ | new_F786_;
  assign new_F765_ = ~new_F729_ & new_F764_;
  assign new_F766_ = new_F785_ | new_F784_;
  assign new_F767_ = new_F729_ & new_F766_;
  assign new_F768_ = new_F727_ & ~new_F737_;
  assign new_F769_ = ~new_F727_ & new_F737_;
  assign new_F770_ = ~new_F726_ | ~new_F751_;
  assign new_F771_ = new_F737_ & new_F770_;
  assign new_F772_ = ~new_F737_ & ~new_F771_;
  assign new_F773_ = new_F737_ | new_F770_;
  assign new_F774_ = ~new_F727_ & new_F728_;
  assign new_F775_ = new_F727_ & ~new_F728_;
  assign new_F776_ = new_F744_ | new_F781_;
  assign new_F777_ = ~new_F744_ & ~new_F780_;
  assign new_F778_ = new_F727_ | new_F744_;
  assign new_F779_ = new_F727_ | new_F728_;
  assign new_F780_ = new_F744_ & new_F781_;
  assign new_F781_ = ~new_F726_ | ~new_F751_;
  assign new_F782_ = new_F759_ & new_F779_;
  assign new_F783_ = ~new_F759_ & ~new_F779_;
  assign new_F784_ = new_F788_ | new_F789_;
  assign new_F785_ = ~new_F730_ & new_F744_;
  assign new_F786_ = new_F790_ | new_F791_;
  assign new_F787_ = new_F730_ & new_F744_;
  assign new_F788_ = ~new_F730_ & ~new_F744_;
  assign new_F789_ = new_F730_ & ~new_F744_;
  assign new_F790_ = new_F730_ & ~new_F744_;
  assign new_F791_ = ~new_F730_ & new_F744_;
  assign new_F792_ = new_G1926_;
  assign new_F793_ = new_G1993_;
  assign new_F794_ = new_G2060_;
  assign new_F795_ = new_G2127_;
  assign new_F796_ = new_G2194_;
  assign new_F797_ = new_G2261_;
  assign new_F798_ = new_F805_ & new_F804_;
  assign new_F799_ = new_F807_ | new_F806_;
  assign new_F800_ = new_F809_ | new_F808_;
  assign new_F801_ = new_F811_ & new_F810_;
  assign new_F802_ = new_F811_ & new_F812_;
  assign new_F803_ = new_F804_ | new_F813_;
  assign new_F804_ = new_F793_ | new_F816_;
  assign new_F805_ = new_F815_ | new_F814_;
  assign new_F806_ = new_F820_ & new_F819_;
  assign new_F807_ = new_F818_ & new_F817_;
  assign new_F808_ = new_F823_ | new_F822_;
  assign new_F809_ = new_F818_ & new_F821_;
  assign new_F810_ = new_F793_ | new_F826_;
  assign new_F811_ = new_F825_ | new_F824_;
  assign new_F812_ = new_F828_ | new_F827_;
  assign new_F813_ = ~new_F804_ & new_F830_;
  assign new_F814_ = ~new_F806_ & new_F818_;
  assign new_F815_ = new_F806_ & ~new_F818_;
  assign new_F816_ = new_F792_ & ~new_F793_;
  assign new_F817_ = ~new_F839_ | ~new_F840_;
  assign new_F818_ = new_F832_ | new_F834_;
  assign new_F819_ = new_F842_ | new_F841_;
  assign new_F820_ = new_F836_ | new_F835_;
  assign new_F821_ = ~new_F844_ | ~new_F843_;
  assign new_F822_ = ~new_F845_ & new_F846_;
  assign new_F823_ = new_F845_ & ~new_F846_;
  assign new_F824_ = ~new_F792_ & new_F793_;
  assign new_F825_ = new_F792_ & ~new_F793_;
  assign new_F826_ = ~new_F808_ | new_F818_;
  assign new_F827_ = new_F808_ & new_F818_;
  assign new_F828_ = ~new_F808_ & ~new_F818_;
  assign new_F829_ = new_F850_ | new_F849_;
  assign new_F830_ = new_F796_ | new_F829_;
  assign new_F831_ = new_F854_ | new_F853_;
  assign new_F832_ = ~new_F796_ & new_F831_;
  assign new_F833_ = new_F852_ | new_F851_;
  assign new_F834_ = new_F796_ & new_F833_;
  assign new_F835_ = new_F794_ & ~new_F804_;
  assign new_F836_ = ~new_F794_ & new_F804_;
  assign new_F837_ = ~new_F793_ | ~new_F818_;
  assign new_F838_ = new_F804_ & new_F837_;
  assign new_F839_ = ~new_F804_ & ~new_F838_;
  assign new_F840_ = new_F804_ | new_F837_;
  assign new_F841_ = ~new_F794_ & new_F795_;
  assign new_F842_ = new_F794_ & ~new_F795_;
  assign new_F843_ = new_F811_ | new_F848_;
  assign new_F844_ = ~new_F811_ & ~new_F847_;
  assign new_F845_ = new_F794_ | new_F811_;
  assign new_F846_ = new_F794_ | new_F795_;
  assign new_F847_ = new_F811_ & new_F848_;
  assign new_F848_ = ~new_F793_ | ~new_F818_;
  assign new_F849_ = new_F826_ & new_F846_;
  assign new_F850_ = ~new_F826_ & ~new_F846_;
  assign new_F851_ = new_F855_ | new_F856_;
  assign new_F852_ = ~new_F797_ & new_F811_;
  assign new_F853_ = new_F857_ | new_F858_;
  assign new_F854_ = new_F797_ & new_F811_;
  assign new_F855_ = ~new_F797_ & ~new_F811_;
  assign new_F856_ = new_F797_ & ~new_F811_;
  assign new_F857_ = new_F797_ & ~new_F811_;
  assign new_F858_ = ~new_F797_ & new_F811_;
  assign new_F859_ = new_G2328_;
  assign new_F860_ = new_G2395_;
  assign new_F861_ = new_G2462_;
  assign new_F862_ = new_G2529_;
  assign new_F863_ = new_G2596_;
  assign new_F864_ = new_G2663_;
  assign new_F865_ = new_F872_ & new_F871_;
  assign new_F866_ = new_F874_ | new_F873_;
  assign new_F867_ = new_F876_ | new_F875_;
  assign new_F868_ = new_F878_ & new_F877_;
  assign new_F869_ = new_F878_ & new_F879_;
  assign new_F870_ = new_F871_ | new_F880_;
  assign new_F871_ = new_F860_ | new_F883_;
  assign new_F872_ = new_F882_ | new_F881_;
  assign new_F873_ = new_F887_ & new_F886_;
  assign new_F874_ = new_F885_ & new_F884_;
  assign new_F875_ = new_F890_ | new_F889_;
  assign new_F876_ = new_F885_ & new_F888_;
  assign new_F877_ = new_F860_ | new_F893_;
  assign new_F878_ = new_F892_ | new_F891_;
  assign new_F879_ = new_F895_ | new_F894_;
  assign new_F880_ = ~new_F871_ & new_F897_;
  assign new_F881_ = ~new_F873_ & new_F885_;
  assign new_F882_ = new_F873_ & ~new_F885_;
  assign new_F883_ = new_F859_ & ~new_F860_;
  assign new_F884_ = ~new_F906_ | ~new_F907_;
  assign new_F885_ = new_F899_ | new_F901_;
  assign new_F886_ = new_F909_ | new_F908_;
  assign new_F887_ = new_F903_ | new_F902_;
  assign new_F888_ = ~new_F911_ | ~new_F910_;
  assign new_F889_ = ~new_F912_ & new_F913_;
  assign new_F890_ = new_F912_ & ~new_F913_;
  assign new_F891_ = ~new_F859_ & new_F860_;
  assign new_F892_ = new_F859_ & ~new_F860_;
  assign new_F893_ = ~new_F875_ | new_F885_;
  assign new_F894_ = new_F875_ & new_F885_;
  assign new_F895_ = ~new_F875_ & ~new_F885_;
  assign new_F896_ = new_F917_ | new_F916_;
  assign new_F897_ = new_F863_ | new_F896_;
  assign new_F898_ = new_F921_ | new_F920_;
  assign new_F899_ = ~new_F863_ & new_F898_;
  assign new_F900_ = new_F919_ | new_F918_;
  assign new_F901_ = new_F863_ & new_F900_;
  assign new_F902_ = new_F861_ & ~new_F871_;
  assign new_F903_ = ~new_F861_ & new_F871_;
  assign new_F904_ = ~new_F860_ | ~new_F885_;
  assign new_F905_ = new_F871_ & new_F904_;
  assign new_F906_ = ~new_F871_ & ~new_F905_;
  assign new_F907_ = new_F871_ | new_F904_;
  assign new_F908_ = ~new_F861_ & new_F862_;
  assign new_F909_ = new_F861_ & ~new_F862_;
  assign new_F910_ = new_F878_ | new_F915_;
  assign new_F911_ = ~new_F878_ & ~new_F914_;
  assign new_F912_ = new_F861_ | new_F878_;
  assign new_F913_ = new_F861_ | new_F862_;
  assign new_F914_ = new_F878_ & new_F915_;
  assign new_F915_ = ~new_F860_ | ~new_F885_;
  assign new_F916_ = new_F893_ & new_F913_;
  assign new_F917_ = ~new_F893_ & ~new_F913_;
  assign new_F918_ = new_F922_ | new_F923_;
  assign new_F919_ = ~new_F864_ & new_F878_;
  assign new_F920_ = new_F924_ | new_F925_;
  assign new_F921_ = new_F864_ & new_F878_;
  assign new_F922_ = ~new_F864_ & ~new_F878_;
  assign new_F923_ = new_F864_ & ~new_F878_;
  assign new_F924_ = new_F864_ & ~new_F878_;
  assign new_F925_ = ~new_F864_ & new_F878_;
  assign new_F926_ = new_G2730_;
  assign new_F927_ = new_G2797_;
  assign new_F928_ = new_G2864_;
  assign new_F929_ = new_G2931_;
  assign new_F930_ = new_G2998_;
  assign new_F931_ = new_G3065_;
  assign new_F932_ = new_F939_ & new_F938_;
  assign new_F933_ = new_F941_ | new_F940_;
  assign new_F934_ = new_F943_ | new_F942_;
  assign new_F935_ = new_F945_ & new_F944_;
  assign new_F936_ = new_F945_ & new_F946_;
  assign new_F937_ = new_F938_ | new_F947_;
  assign new_F938_ = new_F927_ | new_F950_;
  assign new_F939_ = new_F949_ | new_F948_;
  assign new_F940_ = new_F954_ & new_F953_;
  assign new_F941_ = new_F952_ & new_F951_;
  assign new_F942_ = new_F957_ | new_F956_;
  assign new_F943_ = new_F952_ & new_F955_;
  assign new_F944_ = new_F927_ | new_F960_;
  assign new_F945_ = new_F959_ | new_F958_;
  assign new_F946_ = new_F962_ | new_F961_;
  assign new_F947_ = ~new_F938_ & new_F964_;
  assign new_F948_ = ~new_F940_ & new_F952_;
  assign new_F949_ = new_F940_ & ~new_F952_;
  assign new_F950_ = new_F926_ & ~new_F927_;
  assign new_F951_ = ~new_F973_ | ~new_F974_;
  assign new_F952_ = new_F966_ | new_F968_;
  assign new_F953_ = new_F976_ | new_F975_;
  assign new_F954_ = new_F970_ | new_F969_;
  assign new_F955_ = ~new_F978_ | ~new_F977_;
  assign new_F956_ = ~new_F979_ & new_F980_;
  assign new_F957_ = new_F979_ & ~new_F980_;
  assign new_F958_ = ~new_F926_ & new_F927_;
  assign new_F959_ = new_F926_ & ~new_F927_;
  assign new_F960_ = ~new_F942_ | new_F952_;
  assign new_F961_ = new_F942_ & new_F952_;
  assign new_F962_ = ~new_F942_ & ~new_F952_;
  assign new_F963_ = new_F984_ | new_F983_;
  assign new_F964_ = new_F930_ | new_F963_;
  assign new_F965_ = new_F988_ | new_F987_;
  assign new_F966_ = ~new_F930_ & new_F965_;
  assign new_F967_ = new_F986_ | new_F985_;
  assign new_F968_ = new_F930_ & new_F967_;
  assign new_F969_ = new_F928_ & ~new_F938_;
  assign new_F970_ = ~new_F928_ & new_F938_;
  assign new_F971_ = ~new_F927_ | ~new_F952_;
  assign new_F972_ = new_F938_ & new_F971_;
  assign new_F973_ = ~new_F938_ & ~new_F972_;
  assign new_F974_ = new_F938_ | new_F971_;
  assign new_F975_ = ~new_F928_ & new_F929_;
  assign new_F976_ = new_F928_ & ~new_F929_;
  assign new_F977_ = new_F945_ | new_F982_;
  assign new_F978_ = ~new_F945_ & ~new_F981_;
  assign new_F979_ = new_F928_ | new_F945_;
  assign new_F980_ = new_F928_ | new_F929_;
  assign new_F981_ = new_F945_ & new_F982_;
  assign new_F982_ = ~new_F927_ | ~new_F952_;
  assign new_F983_ = new_F960_ & new_F980_;
  assign new_F984_ = ~new_F960_ & ~new_F980_;
  assign new_F985_ = new_F989_ | new_F990_;
  assign new_F986_ = ~new_F931_ & new_F945_;
  assign new_F987_ = new_F991_ | new_F992_;
  assign new_F988_ = new_F931_ & new_F945_;
  assign new_F989_ = ~new_F931_ & ~new_F945_;
  assign new_F990_ = new_F931_ & ~new_F945_;
  assign new_F991_ = new_F931_ & ~new_F945_;
  assign new_F992_ = ~new_F931_ & new_F945_;
  assign new_F993_ = new_G3132_;
  assign new_F994_ = new_G3199_;
  assign new_F995_ = new_G3266_;
  assign new_F996_ = new_G3333_;
  assign new_F997_ = new_G3400_;
  assign new_F998_ = new_G3467_;
  assign new_F999_ = new_F1006_ & new_F1005_;
  assign new_F1000_ = new_F1008_ | new_F1007_;
  assign new_F1001_ = new_F1010_ | new_F1009_;
  assign new_F1002_ = new_F1012_ & new_F1011_;
  assign new_F1003_ = new_F1012_ & new_F1013_;
  assign new_F1004_ = new_F1005_ | new_F1014_;
  assign new_F1005_ = new_F994_ | new_F1017_;
  assign new_F1006_ = new_F1016_ | new_F1015_;
  assign new_F1007_ = new_F1021_ & new_F1020_;
  assign new_F1008_ = new_F1019_ & new_F1018_;
  assign new_F1009_ = new_F1024_ | new_F1023_;
  assign new_F1010_ = new_F1019_ & new_F1022_;
  assign new_F1011_ = new_F994_ | new_F1027_;
  assign new_F1012_ = new_F1026_ | new_F1025_;
  assign new_F1013_ = new_F1029_ | new_F1028_;
  assign new_F1014_ = ~new_F1005_ & new_F1031_;
  assign new_F1015_ = ~new_F1007_ & new_F1019_;
  assign new_F1016_ = new_F1007_ & ~new_F1019_;
  assign new_F1017_ = new_F993_ & ~new_F994_;
  assign new_F1018_ = ~new_F1040_ | ~new_F1041_;
  assign new_F1019_ = new_F1033_ | new_F1035_;
  assign new_F1020_ = new_F1043_ | new_F1042_;
  assign new_F1021_ = new_F1037_ | new_F1036_;
  assign new_F1022_ = ~new_F1045_ | ~new_F1044_;
  assign new_F1023_ = ~new_F1046_ & new_F1047_;
  assign new_F1024_ = new_F1046_ & ~new_F1047_;
  assign new_F1025_ = ~new_F993_ & new_F994_;
  assign new_F1026_ = new_F993_ & ~new_F994_;
  assign new_F1027_ = ~new_F1009_ | new_F1019_;
  assign new_F1028_ = new_F1009_ & new_F1019_;
  assign new_F1029_ = ~new_F1009_ & ~new_F1019_;
  assign new_F1030_ = new_F1051_ | new_F1050_;
  assign new_F1031_ = new_F997_ | new_F1030_;
  assign new_F1032_ = new_F1055_ | new_F1054_;
  assign new_F1033_ = ~new_F997_ & new_F1032_;
  assign new_F1034_ = new_F1053_ | new_F1052_;
  assign new_F1035_ = new_F997_ & new_F1034_;
  assign new_F1036_ = new_F995_ & ~new_F1005_;
  assign new_F1037_ = ~new_F995_ & new_F1005_;
  assign new_F1038_ = ~new_F994_ | ~new_F1019_;
  assign new_F1039_ = new_F1005_ & new_F1038_;
  assign new_F1040_ = ~new_F1005_ & ~new_F1039_;
  assign new_F1041_ = new_F1005_ | new_F1038_;
  assign new_F1042_ = ~new_F995_ & new_F996_;
  assign new_F1043_ = new_F995_ & ~new_F996_;
  assign new_F1044_ = new_F1012_ | new_F1049_;
  assign new_F1045_ = ~new_F1012_ & ~new_F1048_;
  assign new_F1046_ = new_F995_ | new_F1012_;
  assign new_F1047_ = new_F995_ | new_F996_;
  assign new_F1048_ = new_F1012_ & new_F1049_;
  assign new_F1049_ = ~new_F994_ | ~new_F1019_;
  assign new_F1050_ = new_F1027_ & new_F1047_;
  assign new_F1051_ = ~new_F1027_ & ~new_F1047_;
  assign new_F1052_ = new_F1056_ | new_F1057_;
  assign new_F1053_ = ~new_F998_ & new_F1012_;
  assign new_F1054_ = new_F1058_ | new_F1059_;
  assign new_F1055_ = new_F998_ & new_F1012_;
  assign new_F1056_ = ~new_F998_ & ~new_F1012_;
  assign new_F1057_ = new_F998_ & ~new_F1012_;
  assign new_F1058_ = new_F998_ & ~new_F1012_;
  assign new_F1059_ = ~new_F998_ & new_F1012_;
  assign new_F1060_ = new_G3534_;
  assign new_F1061_ = new_G3601_;
  assign new_F1062_ = new_G3668_;
  assign new_F1063_ = new_G3735_;
  assign new_F1064_ = new_G3802_;
  assign new_F1065_ = new_G3869_;
  assign new_F1066_ = new_F1073_ & new_F1072_;
  assign new_F1067_ = new_F1075_ | new_F1074_;
  assign new_F1068_ = new_F1077_ | new_F1076_;
  assign new_F1069_ = new_F1079_ & new_F1078_;
  assign new_F1070_ = new_F1079_ & new_F1080_;
  assign new_F1071_ = new_F1072_ | new_F1081_;
  assign new_F1072_ = new_F1061_ | new_F1084_;
  assign new_F1073_ = new_F1083_ | new_F1082_;
  assign new_F1074_ = new_F1088_ & new_F1087_;
  assign new_F1075_ = new_F1086_ & new_F1085_;
  assign new_F1076_ = new_F1091_ | new_F1090_;
  assign new_F1077_ = new_F1086_ & new_F1089_;
  assign new_F1078_ = new_F1061_ | new_F1094_;
  assign new_F1079_ = new_F1093_ | new_F1092_;
  assign new_F1080_ = new_F1096_ | new_F1095_;
  assign new_F1081_ = ~new_F1072_ & new_F1098_;
  assign new_F1082_ = ~new_F1074_ & new_F1086_;
  assign new_F1083_ = new_F1074_ & ~new_F1086_;
  assign new_F1084_ = new_F1060_ & ~new_F1061_;
  assign new_F1085_ = ~new_F1107_ | ~new_F1108_;
  assign new_F1086_ = new_F1100_ | new_F1102_;
  assign new_F1087_ = new_F1110_ | new_F1109_;
  assign new_F1088_ = new_F1104_ | new_F1103_;
  assign new_F1089_ = ~new_F1112_ | ~new_F1111_;
  assign new_F1090_ = ~new_F1113_ & new_F1114_;
  assign new_F1091_ = new_F1113_ & ~new_F1114_;
  assign new_F1092_ = ~new_F1060_ & new_F1061_;
  assign new_F1093_ = new_F1060_ & ~new_F1061_;
  assign new_F1094_ = ~new_F1076_ | new_F1086_;
  assign new_F1095_ = new_F1076_ & new_F1086_;
  assign new_F1096_ = ~new_F1076_ & ~new_F1086_;
  assign new_F1097_ = new_F1118_ | new_F1117_;
  assign new_F1098_ = new_F1064_ | new_F1097_;
  assign new_F1099_ = new_F1122_ | new_F1121_;
  assign new_F1100_ = ~new_F1064_ & new_F1099_;
  assign new_F1101_ = new_F1120_ | new_F1119_;
  assign new_F1102_ = new_F1064_ & new_F1101_;
  assign new_F1103_ = new_F1062_ & ~new_F1072_;
  assign new_F1104_ = ~new_F1062_ & new_F1072_;
  assign new_F1105_ = ~new_F1061_ | ~new_F1086_;
  assign new_F1106_ = new_F1072_ & new_F1105_;
  assign new_F1107_ = ~new_F1072_ & ~new_F1106_;
  assign new_F1108_ = new_F1072_ | new_F1105_;
  assign new_F1109_ = ~new_F1062_ & new_F1063_;
  assign new_F1110_ = new_F1062_ & ~new_F1063_;
  assign new_F1111_ = new_F1079_ | new_F1116_;
  assign new_F1112_ = ~new_F1079_ & ~new_F1115_;
  assign new_F1113_ = new_F1062_ | new_F1079_;
  assign new_F1114_ = new_F1062_ | new_F1063_;
  assign new_F1115_ = new_F1079_ & new_F1116_;
  assign new_F1116_ = ~new_F1061_ | ~new_F1086_;
  assign new_F1117_ = new_F1094_ & new_F1114_;
  assign new_F1118_ = ~new_F1094_ & ~new_F1114_;
  assign new_F1119_ = new_F1123_ | new_F1124_;
  assign new_F1120_ = ~new_F1065_ & new_F1079_;
  assign new_F1121_ = new_F1125_ | new_F1126_;
  assign new_F1122_ = new_F1065_ & new_F1079_;
  assign new_F1123_ = ~new_F1065_ & ~new_F1079_;
  assign new_F1124_ = new_F1065_ & ~new_F1079_;
  assign new_F1125_ = new_F1065_ & ~new_F1079_;
  assign new_F1126_ = ~new_F1065_ & new_F1079_;
  assign new_F1127_ = new_G3936_;
  assign new_F1128_ = new_G4003_;
  assign new_F1129_ = new_G4070_;
  assign new_F1130_ = new_G4137_;
  assign new_F1131_ = new_G4204_;
  assign new_F1132_ = new_G4271_;
  assign new_F1133_ = new_F1140_ & new_F1139_;
  assign new_F1134_ = new_F1142_ | new_F1141_;
  assign new_F1135_ = new_F1144_ | new_F1143_;
  assign new_F1136_ = new_F1146_ & new_F1145_;
  assign new_F1137_ = new_F1146_ & new_F1147_;
  assign new_F1138_ = new_F1139_ | new_F1148_;
  assign new_F1139_ = new_F1128_ | new_F1151_;
  assign new_F1140_ = new_F1150_ | new_F1149_;
  assign new_F1141_ = new_F1155_ & new_F1154_;
  assign new_F1142_ = new_F1153_ & new_F1152_;
  assign new_F1143_ = new_F1158_ | new_F1157_;
  assign new_F1144_ = new_F1153_ & new_F1156_;
  assign new_F1145_ = new_F1128_ | new_F1161_;
  assign new_F1146_ = new_F1160_ | new_F1159_;
  assign new_F1147_ = new_F1163_ | new_F1162_;
  assign new_F1148_ = ~new_F1139_ & new_F1165_;
  assign new_F1149_ = ~new_F1141_ & new_F1153_;
  assign new_F1150_ = new_F1141_ & ~new_F1153_;
  assign new_F1151_ = new_F1127_ & ~new_F1128_;
  assign new_F1152_ = ~new_F1174_ | ~new_F1175_;
  assign new_F1153_ = new_F1167_ | new_F1169_;
  assign new_F1154_ = new_F1177_ | new_F1176_;
  assign new_F1155_ = new_F1171_ | new_F1170_;
  assign new_F1156_ = ~new_F1179_ | ~new_F1178_;
  assign new_F1157_ = ~new_F1180_ & new_F1181_;
  assign new_F1158_ = new_F1180_ & ~new_F1181_;
  assign new_F1159_ = ~new_F1127_ & new_F1128_;
  assign new_F1160_ = new_F1127_ & ~new_F1128_;
  assign new_F1161_ = ~new_F1143_ | new_F1153_;
  assign new_F1162_ = new_F1143_ & new_F1153_;
  assign new_F1163_ = ~new_F1143_ & ~new_F1153_;
  assign new_F1164_ = new_F1185_ | new_F1184_;
  assign new_F1165_ = new_F1131_ | new_F1164_;
  assign new_F1166_ = new_F1189_ | new_F1188_;
  assign new_F1167_ = ~new_F1131_ & new_F1166_;
  assign new_F1168_ = new_F1187_ | new_F1186_;
  assign new_F1169_ = new_F1131_ & new_F1168_;
  assign new_F1170_ = new_F1129_ & ~new_F1139_;
  assign new_F1171_ = ~new_F1129_ & new_F1139_;
  assign new_F1172_ = ~new_F1128_ | ~new_F1153_;
  assign new_F1173_ = new_F1139_ & new_F1172_;
  assign new_F1174_ = ~new_F1139_ & ~new_F1173_;
  assign new_F1175_ = new_F1139_ | new_F1172_;
  assign new_F1176_ = ~new_F1129_ & new_F1130_;
  assign new_F1177_ = new_F1129_ & ~new_F1130_;
  assign new_F1178_ = new_F1146_ | new_F1183_;
  assign new_F1179_ = ~new_F1146_ & ~new_F1182_;
  assign new_F1180_ = new_F1129_ | new_F1146_;
  assign new_F1181_ = new_F1129_ | new_F1130_;
  assign new_F1182_ = new_F1146_ & new_F1183_;
  assign new_F1183_ = ~new_F1128_ | ~new_F1153_;
  assign new_F1184_ = new_F1161_ & new_F1181_;
  assign new_F1185_ = ~new_F1161_ & ~new_F1181_;
  assign new_F1186_ = new_F1190_ | new_F1191_;
  assign new_F1187_ = ~new_F1132_ & new_F1146_;
  assign new_F1188_ = new_F1192_ | new_F1193_;
  assign new_F1189_ = new_F1132_ & new_F1146_;
  assign new_F1190_ = ~new_F1132_ & ~new_F1146_;
  assign new_F1191_ = new_F1132_ & ~new_F1146_;
  assign new_F1192_ = new_F1132_ & ~new_F1146_;
  assign new_F1193_ = ~new_F1132_ & new_F1146_;
  assign new_F1194_ = new_G4338_;
  assign new_F1195_ = new_G4405_;
  assign new_F1196_ = new_G4472_;
  assign new_F1197_ = new_G4539_;
  assign new_F1198_ = new_G4606_;
  assign new_F1199_ = new_G4673_;
  assign new_F1200_ = new_F1207_ & new_F1206_;
  assign new_F1201_ = new_F1209_ | new_F1208_;
  assign new_F1202_ = new_F1211_ | new_F1210_;
  assign new_F1203_ = new_F1213_ & new_F1212_;
  assign new_F1204_ = new_F1213_ & new_F1214_;
  assign new_F1205_ = new_F1206_ | new_F1215_;
  assign new_F1206_ = new_F1195_ | new_F1218_;
  assign new_F1207_ = new_F1217_ | new_F1216_;
  assign new_F1208_ = new_F1222_ & new_F1221_;
  assign new_F1209_ = new_F1220_ & new_F1219_;
  assign new_F1210_ = new_F1225_ | new_F1224_;
  assign new_F1211_ = new_F1220_ & new_F1223_;
  assign new_F1212_ = new_F1195_ | new_F1228_;
  assign new_F1213_ = new_F1227_ | new_F1226_;
  assign new_F1214_ = new_F1230_ | new_F1229_;
  assign new_F1215_ = ~new_F1206_ & new_F1232_;
  assign new_F1216_ = ~new_F1208_ & new_F1220_;
  assign new_F1217_ = new_F1208_ & ~new_F1220_;
  assign new_F1218_ = new_F1194_ & ~new_F1195_;
  assign new_F1219_ = ~new_F1241_ | ~new_F1242_;
  assign new_F1220_ = new_F1234_ | new_F1236_;
  assign new_F1221_ = new_F1244_ | new_F1243_;
  assign new_F1222_ = new_F1238_ | new_F1237_;
  assign new_F1223_ = ~new_F1246_ | ~new_F1245_;
  assign new_F1224_ = ~new_F1247_ & new_F1248_;
  assign new_F1225_ = new_F1247_ & ~new_F1248_;
  assign new_F1226_ = ~new_F1194_ & new_F1195_;
  assign new_F1227_ = new_F1194_ & ~new_F1195_;
  assign new_F1228_ = ~new_F1210_ | new_F1220_;
  assign new_F1229_ = new_F1210_ & new_F1220_;
  assign new_F1230_ = ~new_F1210_ & ~new_F1220_;
  assign new_F1231_ = new_F1252_ | new_F1251_;
  assign new_F1232_ = new_F1198_ | new_F1231_;
  assign new_F1233_ = new_F1256_ | new_F1255_;
  assign new_F1234_ = ~new_F1198_ & new_F1233_;
  assign new_F1235_ = new_F1254_ | new_F1253_;
  assign new_F1236_ = new_F1198_ & new_F1235_;
  assign new_F1237_ = new_F1196_ & ~new_F1206_;
  assign new_F1238_ = ~new_F1196_ & new_F1206_;
  assign new_F1239_ = ~new_F1195_ | ~new_F1220_;
  assign new_F1240_ = new_F1206_ & new_F1239_;
  assign new_F1241_ = ~new_F1206_ & ~new_F1240_;
  assign new_F1242_ = new_F1206_ | new_F1239_;
  assign new_F1243_ = ~new_F1196_ & new_F1197_;
  assign new_F1244_ = new_F1196_ & ~new_F1197_;
  assign new_F1245_ = new_F1213_ | new_F1250_;
  assign new_F1246_ = ~new_F1213_ & ~new_F1249_;
  assign new_F1247_ = new_F1196_ | new_F1213_;
  assign new_F1248_ = new_F1196_ | new_F1197_;
  assign new_F1249_ = new_F1213_ & new_F1250_;
  assign new_F1250_ = ~new_F1195_ | ~new_F1220_;
  assign new_F1251_ = new_F1228_ & new_F1248_;
  assign new_F1252_ = ~new_F1228_ & ~new_F1248_;
  assign new_F1253_ = new_F1257_ | new_F1258_;
  assign new_F1254_ = ~new_F1199_ & new_F1213_;
  assign new_F1255_ = new_F1259_ | new_F1260_;
  assign new_F1256_ = new_F1199_ & new_F1213_;
  assign new_F1257_ = ~new_F1199_ & ~new_F1213_;
  assign new_F1258_ = new_F1199_ & ~new_F1213_;
  assign new_F1259_ = new_F1199_ & ~new_F1213_;
  assign new_F1260_ = ~new_F1199_ & new_F1213_;
  assign new_F1261_ = new_G4740_;
  assign new_F1262_ = new_G4807_;
  assign new_F1263_ = new_G4874_;
  assign new_F1264_ = new_G4941_;
  assign new_F1265_ = new_G5008_;
  assign new_F1266_ = new_G5075_;
  assign new_F1267_ = new_F1274_ & new_F1273_;
  assign new_F1268_ = new_F1276_ | new_F1275_;
  assign new_F1269_ = new_F1278_ | new_F1277_;
  assign new_F1270_ = new_F1280_ & new_F1279_;
  assign new_F1271_ = new_F1280_ & new_F1281_;
  assign new_F1272_ = new_F1273_ | new_F1282_;
  assign new_F1273_ = new_F1262_ | new_F1285_;
  assign new_F1274_ = new_F1284_ | new_F1283_;
  assign new_F1275_ = new_F1289_ & new_F1288_;
  assign new_F1276_ = new_F1287_ & new_F1286_;
  assign new_F1277_ = new_F1292_ | new_F1291_;
  assign new_F1278_ = new_F1287_ & new_F1290_;
  assign new_F1279_ = new_F1262_ | new_F1295_;
  assign new_F1280_ = new_F1294_ | new_F1293_;
  assign new_F1281_ = new_F1297_ | new_F1296_;
  assign new_F1282_ = ~new_F1273_ & new_F1299_;
  assign new_F1283_ = ~new_F1275_ & new_F1287_;
  assign new_F1284_ = new_F1275_ & ~new_F1287_;
  assign new_F1285_ = new_F1261_ & ~new_F1262_;
  assign new_F1286_ = ~new_F1308_ | ~new_F1309_;
  assign new_F1287_ = new_F1301_ | new_F1303_;
  assign new_F1288_ = new_F1311_ | new_F1310_;
  assign new_F1289_ = new_F1305_ | new_F1304_;
  assign new_F1290_ = ~new_F1313_ | ~new_F1312_;
  assign new_F1291_ = ~new_F1314_ & new_F1315_;
  assign new_F1292_ = new_F1314_ & ~new_F1315_;
  assign new_F1293_ = ~new_F1261_ & new_F1262_;
  assign new_F1294_ = new_F1261_ & ~new_F1262_;
  assign new_F1295_ = ~new_F1277_ | new_F1287_;
  assign new_F1296_ = new_F1277_ & new_F1287_;
  assign new_F1297_ = ~new_F1277_ & ~new_F1287_;
  assign new_F1298_ = new_F1319_ | new_F1318_;
  assign new_F1299_ = new_F1265_ | new_F1298_;
  assign new_F1300_ = new_F1323_ | new_F1322_;
  assign new_F1301_ = ~new_F1265_ & new_F1300_;
  assign new_F1302_ = new_F1321_ | new_F1320_;
  assign new_F1303_ = new_F1265_ & new_F1302_;
  assign new_F1304_ = new_F1263_ & ~new_F1273_;
  assign new_F1305_ = ~new_F1263_ & new_F1273_;
  assign new_F1306_ = ~new_F1262_ | ~new_F1287_;
  assign new_F1307_ = new_F1273_ & new_F1306_;
  assign new_F1308_ = ~new_F1273_ & ~new_F1307_;
  assign new_F1309_ = new_F1273_ | new_F1306_;
  assign new_F1310_ = ~new_F1263_ & new_F1264_;
  assign new_F1311_ = new_F1263_ & ~new_F1264_;
  assign new_F1312_ = new_F1280_ | new_F1317_;
  assign new_F1313_ = ~new_F1280_ & ~new_F1316_;
  assign new_F1314_ = new_F1263_ | new_F1280_;
  assign new_F1315_ = new_F1263_ | new_F1264_;
  assign new_F1316_ = new_F1280_ & new_F1317_;
  assign new_F1317_ = ~new_F1262_ | ~new_F1287_;
  assign new_F1318_ = new_F1295_ & new_F1315_;
  assign new_F1319_ = ~new_F1295_ & ~new_F1315_;
  assign new_F1320_ = new_F1324_ | new_F1325_;
  assign new_F1321_ = ~new_F1266_ & new_F1280_;
  assign new_F1322_ = new_F1326_ | new_F1327_;
  assign new_F1323_ = new_F1266_ & new_F1280_;
  assign new_F1324_ = ~new_F1266_ & ~new_F1280_;
  assign new_F1325_ = new_F1266_ & ~new_F1280_;
  assign new_F1326_ = new_F1266_ & ~new_F1280_;
  assign new_F1327_ = ~new_F1266_ & new_F1280_;
  assign new_F1328_ = new_G5142_;
  assign new_F1329_ = new_G5209_;
  assign new_F1330_ = new_G5276_;
  assign new_F1331_ = new_G5343_;
  assign new_F1332_ = new_G5410_;
  assign new_F1333_ = new_G5477_;
  assign new_F1334_ = new_F1341_ & new_F1340_;
  assign new_F1335_ = new_F1343_ | new_F1342_;
  assign new_F1336_ = new_F1345_ | new_F1344_;
  assign new_F1337_ = new_F1347_ & new_F1346_;
  assign new_F1338_ = new_F1347_ & new_F1348_;
  assign new_F1339_ = new_F1340_ | new_F1349_;
  assign new_F1340_ = new_F1329_ | new_F1352_;
  assign new_F1341_ = new_F1351_ | new_F1350_;
  assign new_F1342_ = new_F1356_ & new_F1355_;
  assign new_F1343_ = new_F1354_ & new_F1353_;
  assign new_F1344_ = new_F1359_ | new_F1358_;
  assign new_F1345_ = new_F1354_ & new_F1357_;
  assign new_F1346_ = new_F1329_ | new_F1362_;
  assign new_F1347_ = new_F1361_ | new_F1360_;
  assign new_F1348_ = new_F1364_ | new_F1363_;
  assign new_F1349_ = ~new_F1340_ & new_F1366_;
  assign new_F1350_ = ~new_F1342_ & new_F1354_;
  assign new_F1351_ = new_F1342_ & ~new_F1354_;
  assign new_F1352_ = new_F1328_ & ~new_F1329_;
  assign new_F1353_ = ~new_F1375_ | ~new_F1376_;
  assign new_F1354_ = new_F1368_ | new_F1370_;
  assign new_F1355_ = new_F1378_ | new_F1377_;
  assign new_F1356_ = new_F1372_ | new_F1371_;
  assign new_F1357_ = ~new_F1380_ | ~new_F1379_;
  assign new_F1358_ = ~new_F1381_ & new_F1382_;
  assign new_F1359_ = new_F1381_ & ~new_F1382_;
  assign new_F1360_ = ~new_F1328_ & new_F1329_;
  assign new_F1361_ = new_F1328_ & ~new_F1329_;
  assign new_F1362_ = ~new_F1344_ | new_F1354_;
  assign new_F1363_ = new_F1344_ & new_F1354_;
  assign new_F1364_ = ~new_F1344_ & ~new_F1354_;
  assign new_F1365_ = new_F1386_ | new_F1385_;
  assign new_F1366_ = new_F1332_ | new_F1365_;
  assign new_F1367_ = new_F1390_ | new_F1389_;
  assign new_F1368_ = ~new_F1332_ & new_F1367_;
  assign new_F1369_ = new_F1388_ | new_F1387_;
  assign new_F1370_ = new_F1332_ & new_F1369_;
  assign new_F1371_ = new_F1330_ & ~new_F1340_;
  assign new_F1372_ = ~new_F1330_ & new_F1340_;
  assign new_F1373_ = ~new_F1329_ | ~new_F1354_;
  assign new_F1374_ = new_F1340_ & new_F1373_;
  assign new_F1375_ = ~new_F1340_ & ~new_F1374_;
  assign new_F1376_ = new_F1340_ | new_F1373_;
  assign new_F1377_ = ~new_F1330_ & new_F1331_;
  assign new_F1378_ = new_F1330_ & ~new_F1331_;
  assign new_F1379_ = new_F1347_ | new_F1384_;
  assign new_F1380_ = ~new_F1347_ & ~new_F1383_;
  assign new_F1381_ = new_F1330_ | new_F1347_;
  assign new_F1382_ = new_F1330_ | new_F1331_;
  assign new_F1383_ = new_F1347_ & new_F1384_;
  assign new_F1384_ = ~new_F1329_ | ~new_F1354_;
  assign new_F1385_ = new_F1362_ & new_F1382_;
  assign new_F1386_ = ~new_F1362_ & ~new_F1382_;
  assign new_F1387_ = new_F1391_ | new_F1392_;
  assign new_F1388_ = ~new_F1333_ & new_F1347_;
  assign new_F1389_ = new_F1393_ | new_F1394_;
  assign new_F1390_ = new_F1333_ & new_F1347_;
  assign new_F1391_ = ~new_F1333_ & ~new_F1347_;
  assign new_F1392_ = new_F1333_ & ~new_F1347_;
  assign new_F1393_ = new_F1333_ & ~new_F1347_;
  assign new_F1394_ = ~new_F1333_ & new_F1347_;
  assign new_F1395_ = new_G5544_;
  assign new_F1396_ = new_G5611_;
  assign new_F1397_ = new_G5678_;
  assign new_F1398_ = new_G5745_;
  assign new_F1399_ = new_G5812_;
  assign new_F1400_ = new_G5879_;
  assign new_F1401_ = new_F1408_ & new_F1407_;
  assign new_F1402_ = new_F1410_ | new_F1409_;
  assign new_F1403_ = new_F1412_ | new_F1411_;
  assign new_F1404_ = new_F1414_ & new_F1413_;
  assign new_F1405_ = new_F1414_ & new_F1415_;
  assign new_F1406_ = new_F1407_ | new_F1416_;
  assign new_F1407_ = new_F1396_ | new_F1419_;
  assign new_F1408_ = new_F1418_ | new_F1417_;
  assign new_F1409_ = new_F1423_ & new_F1422_;
  assign new_F1410_ = new_F1421_ & new_F1420_;
  assign new_F1411_ = new_F1426_ | new_F1425_;
  assign new_F1412_ = new_F1421_ & new_F1424_;
  assign new_F1413_ = new_F1396_ | new_F1429_;
  assign new_F1414_ = new_F1428_ | new_F1427_;
  assign new_F1415_ = new_F1431_ | new_F1430_;
  assign new_F1416_ = ~new_F1407_ & new_F1433_;
  assign new_F1417_ = ~new_F1409_ & new_F1421_;
  assign new_F1418_ = new_F1409_ & ~new_F1421_;
  assign new_F1419_ = new_F1395_ & ~new_F1396_;
  assign new_F1420_ = ~new_F1442_ | ~new_F1443_;
  assign new_F1421_ = new_F1435_ | new_F1437_;
  assign new_F1422_ = new_F1445_ | new_F1444_;
  assign new_F1423_ = new_F1439_ | new_F1438_;
  assign new_F1424_ = ~new_F1447_ | ~new_F1446_;
  assign new_F1425_ = ~new_F1448_ & new_F1449_;
  assign new_F1426_ = new_F1448_ & ~new_F1449_;
  assign new_F1427_ = ~new_F1395_ & new_F1396_;
  assign new_F1428_ = new_F1395_ & ~new_F1396_;
  assign new_F1429_ = ~new_F1411_ | new_F1421_;
  assign new_F1430_ = new_F1411_ & new_F1421_;
  assign new_F1431_ = ~new_F1411_ & ~new_F1421_;
  assign new_F1432_ = new_F1453_ | new_F1452_;
  assign new_F1433_ = new_F1399_ | new_F1432_;
  assign new_F1434_ = new_F1457_ | new_F1456_;
  assign new_F1435_ = ~new_F1399_ & new_F1434_;
  assign new_F1436_ = new_F1455_ | new_F1454_;
  assign new_F1437_ = new_F1399_ & new_F1436_;
  assign new_F1438_ = new_F1397_ & ~new_F1407_;
  assign new_F1439_ = ~new_F1397_ & new_F1407_;
  assign new_F1440_ = ~new_F1396_ | ~new_F1421_;
  assign new_F1441_ = new_F1407_ & new_F1440_;
  assign new_F1442_ = ~new_F1407_ & ~new_F1441_;
  assign new_F1443_ = new_F1407_ | new_F1440_;
  assign new_F1444_ = ~new_F1397_ & new_F1398_;
  assign new_F1445_ = new_F1397_ & ~new_F1398_;
  assign new_F1446_ = new_F1414_ | new_F1451_;
  assign new_F1447_ = ~new_F1414_ & ~new_F1450_;
  assign new_F1448_ = new_F1397_ | new_F1414_;
  assign new_F1449_ = new_F1397_ | new_F1398_;
  assign new_F1450_ = new_F1414_ & new_F1451_;
  assign new_F1451_ = ~new_F1396_ | ~new_F1421_;
  assign new_F1452_ = new_F1429_ & new_F1449_;
  assign new_F1453_ = ~new_F1429_ & ~new_F1449_;
  assign new_F1454_ = new_F1458_ | new_F1459_;
  assign new_F1455_ = ~new_F1400_ & new_F1414_;
  assign new_F1456_ = new_F1460_ | new_F1461_;
  assign new_F1457_ = new_F1400_ & new_F1414_;
  assign new_F1458_ = ~new_F1400_ & ~new_F1414_;
  assign new_F1459_ = new_F1400_ & ~new_F1414_;
  assign new_F1460_ = new_F1400_ & ~new_F1414_;
  assign new_F1461_ = ~new_F1400_ & new_F1414_;
  assign new_C2581_ = ~new_C2520_ & new_C2534_;
  assign new_C2580_ = new_C2520_ & ~new_C2534_;
  assign new_C2579_ = new_C2520_ & ~new_C2534_;
  assign new_C2578_ = ~new_C2520_ & ~new_C2534_;
  assign new_C2577_ = new_C2520_ & new_C2534_;
  assign new_C2576_ = new_C2580_ | new_C2581_;
  assign new_C2575_ = ~new_C2520_ & new_C2534_;
  assign new_C2574_ = new_C2578_ | new_C2579_;
  assign new_C2573_ = ~new_C2549_ & ~new_C2569_;
  assign new_C2572_ = new_C2549_ & new_C2569_;
  assign new_C2571_ = ~new_C2516_ | ~new_C2541_;
  assign new_C2570_ = new_C2534_ & new_C2571_;
  assign new_C2569_ = new_C2517_ | new_C2518_;
  assign new_C2568_ = new_C2517_ | new_C2534_;
  assign new_C2567_ = ~new_C2534_ & ~new_C2570_;
  assign new_C2566_ = new_C2534_ | new_C2571_;
  assign new_C2565_ = new_C2517_ & ~new_C2518_;
  assign new_C2564_ = ~new_C2517_ & new_C2518_;
  assign new_C2563_ = new_C2527_ | new_C2560_;
  assign new_C2562_ = ~new_C2527_ & ~new_C2561_;
  assign new_C2561_ = new_C2527_ & new_C2560_;
  assign new_C2560_ = ~new_C2516_ | ~new_C2541_;
  assign new_C2559_ = ~new_C2517_ & new_C2527_;
  assign new_C2558_ = new_C2517_ & ~new_C2527_;
  assign new_C2557_ = new_C2519_ & new_C2556_;
  assign new_C2556_ = new_C2575_ | new_C2574_;
  assign new_C2555_ = ~new_C2519_ & new_C2554_;
  assign new_C2554_ = new_C2577_ | new_C2576_;
  assign new_C2553_ = new_C2519_ | new_C2552_;
  assign new_C2552_ = new_C2573_ | new_C2572_;
  assign new_C2551_ = ~new_C2531_ & ~new_C2541_;
  assign new_C2550_ = new_C2531_ & new_C2541_;
  assign new_C2549_ = ~new_C2531_ | new_C2541_;
  assign new_C2548_ = new_C2515_ & ~new_C2516_;
  assign new_C2547_ = ~new_C2515_ & new_C2516_;
  assign new_C2546_ = new_C2568_ & ~new_C2569_;
  assign new_C2545_ = ~new_C2568_ & new_C2569_;
  assign new_C2544_ = ~new_C2567_ | ~new_C2566_;
  assign new_C2543_ = new_C2559_ | new_C2558_;
  assign new_C2542_ = new_C2565_ | new_C2564_;
  assign new_C2541_ = new_C2555_ | new_C2557_;
  assign new_C2540_ = ~new_C2562_ | ~new_C2563_;
  assign new_C2539_ = new_C2515_ & ~new_C2516_;
  assign new_C2538_ = new_C2529_ & ~new_C2541_;
  assign new_C2537_ = ~new_C2529_ & new_C2541_;
  assign new_C2536_ = ~new_C2527_ & new_C2553_;
  assign new_C2535_ = new_C2551_ | new_C2550_;
  assign new_C2534_ = new_C2548_ | new_C2547_;
  assign new_C2533_ = new_C2516_ | new_C2549_;
  assign new_C2532_ = new_C2541_ & new_C2544_;
  assign new_C2531_ = new_C2546_ | new_C2545_;
  assign new_C2530_ = new_C2541_ & new_C2540_;
  assign new_C2529_ = new_C2543_ & new_C2542_;
  assign new_C2528_ = new_C2538_ | new_C2537_;
  assign new_C2527_ = new_C2516_ | new_C2539_;
  assign new_C2526_ = new_C2527_ | new_C2536_;
  assign new_C2525_ = new_C2534_ & new_C2535_;
  assign new_C2524_ = new_C2534_ & new_C2533_;
  assign new_C2523_ = new_C2532_ | new_C2531_;
  assign new_C2522_ = new_C2530_ | new_C2529_;
  assign new_C2521_ = new_C2528_ & new_C2527_;
  assign new_C2520_ = new_D6999_;
  assign new_C2519_ = new_D7061_;
  assign new_C2518_ = new_D7128_;
  assign new_C2517_ = new_D7195_;
  assign new_C2516_ = new_D7262_;
  assign new_C2515_ = new_D7329_;
  assign new_C2582_ = new_D7396_;
  assign new_C2583_ = new_D7463_;
  assign new_C2584_ = new_D7530_;
  assign new_C2585_ = new_D7597_;
  assign new_C2586_ = new_D7664_;
  assign new_C2587_ = new_D7731_;
  assign new_C2588_ = new_C2595_ & new_C2594_;
  assign new_C2589_ = new_C2597_ | new_C2596_;
  assign new_C2590_ = new_C2599_ | new_C2598_;
  assign new_C2591_ = new_C2601_ & new_C2600_;
  assign new_C2592_ = new_C2601_ & new_C2602_;
  assign new_C2593_ = new_C2594_ | new_C2603_;
  assign new_C2594_ = new_C2583_ | new_C2606_;
  assign new_C2595_ = new_C2605_ | new_C2604_;
  assign new_C2596_ = new_C2610_ & new_C2609_;
  assign new_C2597_ = new_C2608_ & new_C2607_;
  assign new_C2598_ = new_C2613_ | new_C2612_;
  assign new_C2599_ = new_C2608_ & new_C2611_;
  assign new_C2600_ = new_C2583_ | new_C2616_;
  assign new_C2601_ = new_C2615_ | new_C2614_;
  assign new_C2602_ = new_C2618_ | new_C2617_;
  assign new_C2603_ = ~new_C2594_ & new_C2620_;
  assign new_C2604_ = ~new_C2596_ & new_C2608_;
  assign new_C2605_ = new_C2596_ & ~new_C2608_;
  assign new_C2606_ = new_C2582_ & ~new_C2583_;
  assign new_C2607_ = ~new_C2629_ | ~new_C2630_;
  assign new_C2608_ = new_C2622_ | new_C2624_;
  assign new_C2609_ = new_C2632_ | new_C2631_;
  assign new_C2610_ = new_C2626_ | new_C2625_;
  assign new_C2611_ = ~new_C2634_ | ~new_C2633_;
  assign new_C2612_ = ~new_C2635_ & new_C2636_;
  assign new_C2613_ = new_C2635_ & ~new_C2636_;
  assign new_C2614_ = ~new_C2582_ & new_C2583_;
  assign new_C2615_ = new_C2582_ & ~new_C2583_;
  assign new_C2616_ = ~new_C2598_ | new_C2608_;
  assign new_C2617_ = new_C2598_ & new_C2608_;
  assign new_C2618_ = ~new_C2598_ & ~new_C2608_;
  assign new_C2619_ = new_C2640_ | new_C2639_;
  assign new_C2620_ = new_C2586_ | new_C2619_;
  assign new_C2621_ = new_C2644_ | new_C2643_;
  assign new_C2622_ = ~new_C2586_ & new_C2621_;
  assign new_C2623_ = new_C2642_ | new_C2641_;
  assign new_C2624_ = new_C2586_ & new_C2623_;
  assign new_C2625_ = new_C2584_ & ~new_C2594_;
  assign new_C2626_ = ~new_C2584_ & new_C2594_;
  assign new_C2627_ = ~new_C2583_ | ~new_C2608_;
  assign new_C2628_ = new_C2594_ & new_C2627_;
  assign new_C2629_ = ~new_C2594_ & ~new_C2628_;
  assign new_C2630_ = new_C2594_ | new_C2627_;
  assign new_C2631_ = ~new_C2584_ & new_C2585_;
  assign new_C2632_ = new_C2584_ & ~new_C2585_;
  assign new_C2633_ = new_C2601_ | new_C2638_;
  assign new_C2634_ = ~new_C2601_ & ~new_C2637_;
  assign new_C2635_ = new_C2584_ | new_C2601_;
  assign new_C2636_ = new_C2584_ | new_C2585_;
  assign new_C2637_ = new_C2601_ & new_C2638_;
  assign new_C2638_ = ~new_C2583_ | ~new_C2608_;
  assign new_C2639_ = new_C2616_ & new_C2636_;
  assign new_C2640_ = ~new_C2616_ & ~new_C2636_;
  assign new_C2641_ = new_C2645_ | new_C2646_;
  assign new_C2642_ = ~new_C2587_ & new_C2601_;
  assign new_C2643_ = new_C2647_ | new_C2648_;
  assign new_C2644_ = new_C2587_ & new_C2601_;
  assign new_C2645_ = ~new_C2587_ & ~new_C2601_;
  assign new_C2646_ = new_C2587_ & ~new_C2601_;
  assign new_C2647_ = new_C2587_ & ~new_C2601_;
  assign new_C2648_ = ~new_C2587_ & new_C2601_;
  assign new_C2649_ = new_D7798_;
  assign new_C2650_ = new_D7865_;
  assign new_C2651_ = new_D7932_;
  assign new_C2652_ = new_D7999_;
  assign new_C2653_ = new_D8066_;
  assign new_C2654_ = new_D8133_;
  assign new_C2655_ = new_C2662_ & new_C2661_;
  assign new_C2656_ = new_C2664_ | new_C2663_;
  assign new_C2657_ = new_C2666_ | new_C2665_;
  assign new_C2658_ = new_C2668_ & new_C2667_;
  assign new_C2659_ = new_C2668_ & new_C2669_;
  assign new_C2660_ = new_C2661_ | new_C2670_;
  assign new_C2661_ = new_C2650_ | new_C2673_;
  assign new_C2662_ = new_C2672_ | new_C2671_;
  assign new_C2663_ = new_C2677_ & new_C2676_;
  assign new_C2664_ = new_C2675_ & new_C2674_;
  assign new_C2665_ = new_C2680_ | new_C2679_;
  assign new_C2666_ = new_C2675_ & new_C2678_;
  assign new_C2667_ = new_C2650_ | new_C2683_;
  assign new_C2668_ = new_C2682_ | new_C2681_;
  assign new_C2669_ = new_C2685_ | new_C2684_;
  assign new_C2670_ = ~new_C2661_ & new_C2687_;
  assign new_C2671_ = ~new_C2663_ & new_C2675_;
  assign new_C2672_ = new_C2663_ & ~new_C2675_;
  assign new_C2673_ = new_C2649_ & ~new_C2650_;
  assign new_C2674_ = ~new_C2696_ | ~new_C2697_;
  assign new_C2675_ = new_C2689_ | new_C2691_;
  assign new_C2676_ = new_C2699_ | new_C2698_;
  assign new_C2677_ = new_C2693_ | new_C2692_;
  assign new_C2678_ = ~new_C2701_ | ~new_C2700_;
  assign new_C2679_ = ~new_C2702_ & new_C2703_;
  assign new_C2680_ = new_C2702_ & ~new_C2703_;
  assign new_C2681_ = ~new_C2649_ & new_C2650_;
  assign new_C2682_ = new_C2649_ & ~new_C2650_;
  assign new_C2683_ = ~new_C2665_ | new_C2675_;
  assign new_C2684_ = new_C2665_ & new_C2675_;
  assign new_C2685_ = ~new_C2665_ & ~new_C2675_;
  assign new_C2686_ = new_C2707_ | new_C2706_;
  assign new_C2687_ = new_C2653_ | new_C2686_;
  assign new_C2688_ = new_C2711_ | new_C2710_;
  assign new_C2689_ = ~new_C2653_ & new_C2688_;
  assign new_C2690_ = new_C2709_ | new_C2708_;
  assign new_C2691_ = new_C2653_ & new_C2690_;
  assign new_C2692_ = new_C2651_ & ~new_C2661_;
  assign new_C2693_ = ~new_C2651_ & new_C2661_;
  assign new_C2694_ = ~new_C2650_ | ~new_C2675_;
  assign new_C2695_ = new_C2661_ & new_C2694_;
  assign new_C2696_ = ~new_C2661_ & ~new_C2695_;
  assign new_C2697_ = new_C2661_ | new_C2694_;
  assign new_C2698_ = ~new_C2651_ & new_C2652_;
  assign new_C2699_ = new_C2651_ & ~new_C2652_;
  assign new_C2700_ = new_C2668_ | new_C2705_;
  assign new_C2701_ = ~new_C2668_ & ~new_C2704_;
  assign new_C2702_ = new_C2651_ | new_C2668_;
  assign new_C2703_ = new_C2651_ | new_C2652_;
  assign new_C2704_ = new_C2668_ & new_C2705_;
  assign new_C2705_ = ~new_C2650_ | ~new_C2675_;
  assign new_C2706_ = new_C2683_ & new_C2703_;
  assign new_C2707_ = ~new_C2683_ & ~new_C2703_;
  assign new_C2708_ = new_C2712_ | new_C2713_;
  assign new_C2709_ = ~new_C2654_ & new_C2668_;
  assign new_C2710_ = new_C2714_ | new_C2715_;
  assign new_C2711_ = new_C2654_ & new_C2668_;
  assign new_C2712_ = ~new_C2654_ & ~new_C2668_;
  assign new_C2713_ = new_C2654_ & ~new_C2668_;
  assign new_C2714_ = new_C2654_ & ~new_C2668_;
  assign new_C2715_ = ~new_C2654_ & new_C2668_;
  assign new_C2716_ = new_D8200_;
  assign new_C2717_ = new_D8267_;
  assign new_C2718_ = new_D8334_;
  assign new_C2719_ = new_D8401_;
  assign new_C2720_ = new_D8468_;
  assign new_C2721_ = new_D8535_;
  assign new_C2722_ = new_C2729_ & new_C2728_;
  assign new_C2723_ = new_C2731_ | new_C2730_;
  assign new_C2724_ = new_C2733_ | new_C2732_;
  assign new_C2725_ = new_C2735_ & new_C2734_;
  assign new_C2726_ = new_C2735_ & new_C2736_;
  assign new_C2727_ = new_C2728_ | new_C2737_;
  assign new_C2728_ = new_C2717_ | new_C2740_;
  assign new_C2729_ = new_C2739_ | new_C2738_;
  assign new_C2730_ = new_C2744_ & new_C2743_;
  assign new_C2731_ = new_C2742_ & new_C2741_;
  assign new_C2732_ = new_C2747_ | new_C2746_;
  assign new_C2733_ = new_C2742_ & new_C2745_;
  assign new_C2734_ = new_C2717_ | new_C2750_;
  assign new_C2735_ = new_C2749_ | new_C2748_;
  assign new_C2736_ = new_C2752_ | new_C2751_;
  assign new_C2737_ = ~new_C2728_ & new_C2754_;
  assign new_C2738_ = ~new_C2730_ & new_C2742_;
  assign new_C2739_ = new_C2730_ & ~new_C2742_;
  assign new_C2740_ = new_C2716_ & ~new_C2717_;
  assign new_C2741_ = ~new_C2763_ | ~new_C2764_;
  assign new_C2742_ = new_C2756_ | new_C2758_;
  assign new_C2743_ = new_C2766_ | new_C2765_;
  assign new_C2744_ = new_C2760_ | new_C2759_;
  assign new_C2745_ = ~new_C2768_ | ~new_C2767_;
  assign new_C2746_ = ~new_C2769_ & new_C2770_;
  assign new_C2747_ = new_C2769_ & ~new_C2770_;
  assign new_C2748_ = ~new_C2716_ & new_C2717_;
  assign new_C2749_ = new_C2716_ & ~new_C2717_;
  assign new_C2750_ = ~new_C2732_ | new_C2742_;
  assign new_C2751_ = new_C2732_ & new_C2742_;
  assign new_C2752_ = ~new_C2732_ & ~new_C2742_;
  assign new_C2753_ = new_C2774_ | new_C2773_;
  assign new_C2754_ = new_C2720_ | new_C2753_;
  assign new_C2755_ = new_C2778_ | new_C2777_;
  assign new_C2756_ = ~new_C2720_ & new_C2755_;
  assign new_C2757_ = new_C2776_ | new_C2775_;
  assign new_C2758_ = new_C2720_ & new_C2757_;
  assign new_C2759_ = new_C2718_ & ~new_C2728_;
  assign new_C2760_ = ~new_C2718_ & new_C2728_;
  assign new_C2761_ = ~new_C2717_ | ~new_C2742_;
  assign new_C2762_ = new_C2728_ & new_C2761_;
  assign new_C2763_ = ~new_C2728_ & ~new_C2762_;
  assign new_C2764_ = new_C2728_ | new_C2761_;
  assign new_C2765_ = ~new_C2718_ & new_C2719_;
  assign new_C2766_ = new_C2718_ & ~new_C2719_;
  assign new_C2767_ = new_C2735_ | new_C2772_;
  assign new_C2768_ = ~new_C2735_ & ~new_C2771_;
  assign new_C2769_ = new_C2718_ | new_C2735_;
  assign new_C2770_ = new_C2718_ | new_C2719_;
  assign new_C2771_ = new_C2735_ & new_C2772_;
  assign new_C2772_ = ~new_C2717_ | ~new_C2742_;
  assign new_C2773_ = new_C2750_ & new_C2770_;
  assign new_C2774_ = ~new_C2750_ & ~new_C2770_;
  assign new_C2775_ = new_C2779_ | new_C2780_;
  assign new_C2776_ = ~new_C2721_ & new_C2735_;
  assign new_C2777_ = new_C2781_ | new_C2782_;
  assign new_C2778_ = new_C2721_ & new_C2735_;
  assign new_C2779_ = ~new_C2721_ & ~new_C2735_;
  assign new_C2780_ = new_C2721_ & ~new_C2735_;
  assign new_C2781_ = new_C2721_ & ~new_C2735_;
  assign new_C2782_ = ~new_C2721_ & new_C2735_;
  assign new_C2783_ = new_D8602_;
  assign new_C2784_ = new_D8669_;
  assign new_C2785_ = new_D8736_;
  assign new_C2786_ = new_D8803_;
  assign new_C2787_ = new_D8870_;
  assign new_C2788_ = new_D8937_;
  assign new_C2789_ = new_C2796_ & new_C2795_;
  assign new_C2790_ = new_C2798_ | new_C2797_;
  assign new_C2791_ = new_C2800_ | new_C2799_;
  assign new_C2792_ = new_C2802_ & new_C2801_;
  assign new_C2793_ = new_C2802_ & new_C2803_;
  assign new_C2794_ = new_C2795_ | new_C2804_;
  assign new_C2795_ = new_C2784_ | new_C2807_;
  assign new_C2796_ = new_C2806_ | new_C2805_;
  assign new_C2797_ = new_C2811_ & new_C2810_;
  assign new_C2798_ = new_C2809_ & new_C2808_;
  assign new_C2799_ = new_C2814_ | new_C2813_;
  assign new_C2800_ = new_C2809_ & new_C2812_;
  assign new_C2801_ = new_C2784_ | new_C2817_;
  assign new_C2802_ = new_C2816_ | new_C2815_;
  assign new_C2803_ = new_C2819_ | new_C2818_;
  assign new_C2804_ = ~new_C2795_ & new_C2821_;
  assign new_C2805_ = ~new_C2797_ & new_C2809_;
  assign new_C2806_ = new_C2797_ & ~new_C2809_;
  assign new_C2807_ = new_C2783_ & ~new_C2784_;
  assign new_C2808_ = ~new_C2830_ | ~new_C2831_;
  assign new_C2809_ = new_C2823_ | new_C2825_;
  assign new_C2810_ = new_C2833_ | new_C2832_;
  assign new_C2811_ = new_C2827_ | new_C2826_;
  assign new_C2812_ = ~new_C2835_ | ~new_C2834_;
  assign new_C2813_ = ~new_C2836_ & new_C2837_;
  assign new_C2814_ = new_C2836_ & ~new_C2837_;
  assign new_C2815_ = ~new_C2783_ & new_C2784_;
  assign new_C2816_ = new_C2783_ & ~new_C2784_;
  assign new_C2817_ = ~new_C2799_ | new_C2809_;
  assign new_C2818_ = new_C2799_ & new_C2809_;
  assign new_C2819_ = ~new_C2799_ & ~new_C2809_;
  assign new_C2820_ = new_C2841_ | new_C2840_;
  assign new_C2821_ = new_C2787_ | new_C2820_;
  assign new_C2822_ = new_C2845_ | new_C2844_;
  assign new_C2823_ = ~new_C2787_ & new_C2822_;
  assign new_C2824_ = new_C2843_ | new_C2842_;
  assign new_C2825_ = new_C2787_ & new_C2824_;
  assign new_C2826_ = new_C2785_ & ~new_C2795_;
  assign new_C2827_ = ~new_C2785_ & new_C2795_;
  assign new_C2828_ = ~new_C2784_ | ~new_C2809_;
  assign new_C2829_ = new_C2795_ & new_C2828_;
  assign new_C2830_ = ~new_C2795_ & ~new_C2829_;
  assign new_C2831_ = new_C2795_ | new_C2828_;
  assign new_C2832_ = ~new_C2785_ & new_C2786_;
  assign new_C2833_ = new_C2785_ & ~new_C2786_;
  assign new_C2834_ = new_C2802_ | new_C2839_;
  assign new_C2835_ = ~new_C2802_ & ~new_C2838_;
  assign new_C2836_ = new_C2785_ | new_C2802_;
  assign new_C2837_ = new_C2785_ | new_C2786_;
  assign new_C2838_ = new_C2802_ & new_C2839_;
  assign new_C2839_ = ~new_C2784_ | ~new_C2809_;
  assign new_C2840_ = new_C2817_ & new_C2837_;
  assign new_C2841_ = ~new_C2817_ & ~new_C2837_;
  assign new_C2842_ = new_C2846_ | new_C2847_;
  assign new_C2843_ = ~new_C2788_ & new_C2802_;
  assign new_C2844_ = new_C2848_ | new_C2849_;
  assign new_C2845_ = new_C2788_ & new_C2802_;
  assign new_C2846_ = ~new_C2788_ & ~new_C2802_;
  assign new_C2847_ = new_C2788_ & ~new_C2802_;
  assign new_C2848_ = new_C2788_ & ~new_C2802_;
  assign new_C2849_ = ~new_C2788_ & new_C2802_;
  assign new_C2850_ = new_D9004_;
  assign new_C2851_ = new_D9071_;
  assign new_C2852_ = new_D9138_;
  assign new_C2853_ = new_D9205_;
  assign new_C2854_ = new_D9272_;
  assign new_C2855_ = new_D9339_;
  assign new_C2856_ = new_C2863_ & new_C2862_;
  assign new_C2857_ = new_C2865_ | new_C2864_;
  assign new_C2858_ = new_C2867_ | new_C2866_;
  assign new_C2859_ = new_C2869_ & new_C2868_;
  assign new_C2860_ = new_C2869_ & new_C2870_;
  assign new_C2861_ = new_C2862_ | new_C2871_;
  assign new_C2862_ = new_C2851_ | new_C2874_;
  assign new_C2863_ = new_C2873_ | new_C2872_;
  assign new_C2864_ = new_C2878_ & new_C2877_;
  assign new_C2865_ = new_C2876_ & new_C2875_;
  assign new_C2866_ = new_C2881_ | new_C2880_;
  assign new_C2867_ = new_C2876_ & new_C2879_;
  assign new_C2868_ = new_C2851_ | new_C2884_;
  assign new_C2869_ = new_C2883_ | new_C2882_;
  assign new_C2870_ = new_C2886_ | new_C2885_;
  assign new_C2871_ = ~new_C2862_ & new_C2888_;
  assign new_C2872_ = ~new_C2864_ & new_C2876_;
  assign new_C2873_ = new_C2864_ & ~new_C2876_;
  assign new_C2874_ = new_C2850_ & ~new_C2851_;
  assign new_C2875_ = ~new_C2897_ | ~new_C2898_;
  assign new_C2876_ = new_C2890_ | new_C2892_;
  assign new_C2877_ = new_C2900_ | new_C2899_;
  assign new_C2878_ = new_C2894_ | new_C2893_;
  assign new_C2879_ = ~new_C2902_ | ~new_C2901_;
  assign new_C2880_ = ~new_C2903_ & new_C2904_;
  assign new_C2881_ = new_C2903_ & ~new_C2904_;
  assign new_C2882_ = ~new_C2850_ & new_C2851_;
  assign new_C2883_ = new_C2850_ & ~new_C2851_;
  assign new_C2884_ = ~new_C2866_ | new_C2876_;
  assign new_C2885_ = new_C2866_ & new_C2876_;
  assign new_C2886_ = ~new_C2866_ & ~new_C2876_;
  assign new_C2887_ = new_C2908_ | new_C2907_;
  assign new_C2888_ = new_C2854_ | new_C2887_;
  assign new_C2889_ = new_C2912_ | new_C2911_;
  assign new_C2890_ = ~new_C2854_ & new_C2889_;
  assign new_C2891_ = new_C2910_ | new_C2909_;
  assign new_C2892_ = new_C2854_ & new_C2891_;
  assign new_C2893_ = new_C2852_ & ~new_C2862_;
  assign new_C2894_ = ~new_C2852_ & new_C2862_;
  assign new_C2895_ = ~new_C2851_ | ~new_C2876_;
  assign new_C2896_ = new_C2862_ & new_C2895_;
  assign new_C2897_ = ~new_C2862_ & ~new_C2896_;
  assign new_C2898_ = new_C2862_ | new_C2895_;
  assign new_C2899_ = ~new_C2852_ & new_C2853_;
  assign new_C2900_ = new_C2852_ & ~new_C2853_;
  assign new_C2901_ = new_C2869_ | new_C2906_;
  assign new_C2902_ = ~new_C2869_ & ~new_C2905_;
  assign new_C2903_ = new_C2852_ | new_C2869_;
  assign new_C2904_ = new_C2852_ | new_C2853_;
  assign new_C2905_ = new_C2869_ & new_C2906_;
  assign new_C2906_ = ~new_C2851_ | ~new_C2876_;
  assign new_C2907_ = new_C2884_ & new_C2904_;
  assign new_C2908_ = ~new_C2884_ & ~new_C2904_;
  assign new_C2909_ = new_C2913_ | new_C2914_;
  assign new_C2910_ = ~new_C2855_ & new_C2869_;
  assign new_C2911_ = new_C2915_ | new_C2916_;
  assign new_C2912_ = new_C2855_ & new_C2869_;
  assign new_C2913_ = ~new_C2855_ & ~new_C2869_;
  assign new_C2914_ = new_C2855_ & ~new_C2869_;
  assign new_C2915_ = new_C2855_ & ~new_C2869_;
  assign new_C2916_ = ~new_C2855_ & new_C2869_;
  assign new_C2917_ = new_D9406_;
  assign new_C2918_ = new_D9473_;
  assign new_C2919_ = new_D9540_;
  assign new_C2920_ = new_D9607_;
  assign new_C2921_ = new_D9674_;
  assign new_C2922_ = new_D9741_;
  assign new_C2923_ = new_C2930_ & new_C2929_;
  assign new_C2924_ = new_C2932_ | new_C2931_;
  assign new_C2925_ = new_C2934_ | new_C2933_;
  assign new_C2926_ = new_C2936_ & new_C2935_;
  assign new_C2927_ = new_C2936_ & new_C2937_;
  assign new_C2928_ = new_C2929_ | new_C2938_;
  assign new_C2929_ = new_C2918_ | new_C2941_;
  assign new_C2930_ = new_C2940_ | new_C2939_;
  assign new_C2931_ = new_C2945_ & new_C2944_;
  assign new_C2932_ = new_C2943_ & new_C2942_;
  assign new_C2933_ = new_C2948_ | new_C2947_;
  assign new_C2934_ = new_C2943_ & new_C2946_;
  assign new_C2935_ = new_C2918_ | new_C2951_;
  assign new_C2936_ = new_C2950_ | new_C2949_;
  assign new_C2937_ = new_C2953_ | new_C2952_;
  assign new_C2938_ = ~new_C2929_ & new_C2955_;
  assign new_C2939_ = ~new_C2931_ & new_C2943_;
  assign new_C2940_ = new_C2931_ & ~new_C2943_;
  assign new_C2941_ = new_C2917_ & ~new_C2918_;
  assign new_C2942_ = ~new_C2964_ | ~new_C2965_;
  assign new_C2943_ = new_C2957_ | new_C2959_;
  assign new_C2944_ = new_C2967_ | new_C2966_;
  assign new_C2945_ = new_C2961_ | new_C2960_;
  assign new_C2946_ = ~new_C2969_ | ~new_C2968_;
  assign new_C2947_ = ~new_C2970_ & new_C2971_;
  assign new_C2948_ = new_C2970_ & ~new_C2971_;
  assign new_C2949_ = ~new_C2917_ & new_C2918_;
  assign new_C2950_ = new_C2917_ & ~new_C2918_;
  assign new_C2951_ = ~new_C2933_ | new_C2943_;
  assign new_C2952_ = new_C2933_ & new_C2943_;
  assign new_C2953_ = ~new_C2933_ & ~new_C2943_;
  assign new_C2954_ = new_C2975_ | new_C2974_;
  assign new_C2955_ = new_C2921_ | new_C2954_;
  assign new_C2956_ = new_C2979_ | new_C2978_;
  assign new_C2957_ = ~new_C2921_ & new_C2956_;
  assign new_C2958_ = new_C2977_ | new_C2976_;
  assign new_C2959_ = new_C2921_ & new_C2958_;
  assign new_C2960_ = new_C2919_ & ~new_C2929_;
  assign new_C2961_ = ~new_C2919_ & new_C2929_;
  assign new_C2962_ = ~new_C2918_ | ~new_C2943_;
  assign new_C2963_ = new_C2929_ & new_C2962_;
  assign new_C2964_ = ~new_C2929_ & ~new_C2963_;
  assign new_C2965_ = new_C2929_ | new_C2962_;
  assign new_C2966_ = ~new_C2919_ & new_C2920_;
  assign new_C2967_ = new_C2919_ & ~new_C2920_;
  assign new_C2968_ = new_C2936_ | new_C2973_;
  assign new_C2969_ = ~new_C2936_ & ~new_C2972_;
  assign new_C2970_ = new_C2919_ | new_C2936_;
  assign new_C2971_ = new_C2919_ | new_C2920_;
  assign new_C2972_ = new_C2936_ & new_C2973_;
  assign new_C2973_ = ~new_C2918_ | ~new_C2943_;
  assign new_C2974_ = new_C2951_ & new_C2971_;
  assign new_C2975_ = ~new_C2951_ & ~new_C2971_;
  assign new_C2976_ = new_C2980_ | new_C2981_;
  assign new_C2977_ = ~new_C2922_ & new_C2936_;
  assign new_C2978_ = new_C2982_ | new_C2983_;
  assign new_C2979_ = new_C2922_ & new_C2936_;
  assign new_C2980_ = ~new_C2922_ & ~new_C2936_;
  assign new_C2981_ = new_C2922_ & ~new_C2936_;
  assign new_C2982_ = new_C2922_ & ~new_C2936_;
  assign new_C2983_ = ~new_C2922_ & new_C2936_;
  assign new_C2984_ = new_D9808_;
  assign new_C2985_ = new_D9875_;
  assign new_C2986_ = new_D9942_;
  assign new_C2987_ = new_E10_;
  assign new_C2988_ = new_E77_;
  assign new_C2989_ = new_E144_;
  assign new_C2990_ = new_C2997_ & new_C2996_;
  assign new_C2991_ = new_C2999_ | new_C2998_;
  assign new_C2992_ = new_C3001_ | new_C3000_;
  assign new_C2993_ = new_C3003_ & new_C3002_;
  assign new_C2994_ = new_C3003_ & new_C3004_;
  assign new_C2995_ = new_C2996_ | new_C3005_;
  assign new_C2996_ = new_C2985_ | new_C3008_;
  assign new_C2997_ = new_C3007_ | new_C3006_;
  assign new_C2998_ = new_C3012_ & new_C3011_;
  assign new_C2999_ = new_C3010_ & new_C3009_;
  assign new_C3000_ = new_C3015_ | new_C3014_;
  assign new_C3001_ = new_C3010_ & new_C3013_;
  assign new_C3002_ = new_C2985_ | new_C3018_;
  assign new_C3003_ = new_C3017_ | new_C3016_;
  assign new_C3004_ = new_C3020_ | new_C3019_;
  assign new_C3005_ = ~new_C2996_ & new_C3022_;
  assign new_C3006_ = ~new_C2998_ & new_C3010_;
  assign new_C3007_ = new_C2998_ & ~new_C3010_;
  assign new_C3008_ = new_C2984_ & ~new_C2985_;
  assign new_C3009_ = ~new_C3031_ | ~new_C3032_;
  assign new_C3010_ = new_C3024_ | new_C3026_;
  assign new_C3011_ = new_C3034_ | new_C3033_;
  assign new_C3012_ = new_C3028_ | new_C3027_;
  assign new_C3013_ = ~new_C3036_ | ~new_C3035_;
  assign new_C3014_ = ~new_C3037_ & new_C3038_;
  assign new_C3015_ = new_C3037_ & ~new_C3038_;
  assign new_C3016_ = ~new_C2984_ & new_C2985_;
  assign new_C3017_ = new_C2984_ & ~new_C2985_;
  assign new_C3018_ = ~new_C3000_ | new_C3010_;
  assign new_C3019_ = new_C3000_ & new_C3010_;
  assign new_C3020_ = ~new_C3000_ & ~new_C3010_;
  assign new_C3021_ = new_C3042_ | new_C3041_;
  assign new_C3022_ = new_C2988_ | new_C3021_;
  assign new_C3023_ = new_C3046_ | new_C3045_;
  assign new_C3024_ = ~new_C2988_ & new_C3023_;
  assign new_C3025_ = new_C3044_ | new_C3043_;
  assign new_C3026_ = new_C2988_ & new_C3025_;
  assign new_C3027_ = new_C2986_ & ~new_C2996_;
  assign new_C3028_ = ~new_C2986_ & new_C2996_;
  assign new_C3029_ = ~new_C2985_ | ~new_C3010_;
  assign new_C3030_ = new_C2996_ & new_C3029_;
  assign new_C3031_ = ~new_C2996_ & ~new_C3030_;
  assign new_C3032_ = new_C2996_ | new_C3029_;
  assign new_C3033_ = ~new_C2986_ & new_C2987_;
  assign new_C3034_ = new_C2986_ & ~new_C2987_;
  assign new_C3035_ = new_C3003_ | new_C3040_;
  assign new_C3036_ = ~new_C3003_ & ~new_C3039_;
  assign new_C3037_ = new_C2986_ | new_C3003_;
  assign new_C3038_ = new_C2986_ | new_C2987_;
  assign new_C3039_ = new_C3003_ & new_C3040_;
  assign new_C3040_ = ~new_C2985_ | ~new_C3010_;
  assign new_C3041_ = new_C3018_ & new_C3038_;
  assign new_C3042_ = ~new_C3018_ & ~new_C3038_;
  assign new_C3043_ = new_C3047_ | new_C3048_;
  assign new_C3044_ = ~new_C2989_ & new_C3003_;
  assign new_C3045_ = new_C3049_ | new_C3050_;
  assign new_C3046_ = new_C2989_ & new_C3003_;
  assign new_C3047_ = ~new_C2989_ & ~new_C3003_;
  assign new_C3048_ = new_C2989_ & ~new_C3003_;
  assign new_C3049_ = new_C2989_ & ~new_C3003_;
  assign new_C3050_ = ~new_C2989_ & new_C3003_;
  assign new_C3051_ = new_E211_;
  assign new_C3052_ = new_E278_;
  assign new_C3053_ = new_E345_;
  assign new_C3054_ = new_E412_;
  assign new_C3055_ = new_E479_;
  assign new_C3056_ = new_E546_;
  assign new_C3057_ = new_C3064_ & new_C3063_;
  assign new_C3058_ = new_C3066_ | new_C3065_;
  assign new_C3059_ = new_C3068_ | new_C3067_;
  assign new_C3060_ = new_C3070_ & new_C3069_;
  assign new_C3061_ = new_C3070_ & new_C3071_;
  assign new_C3062_ = new_C3063_ | new_C3072_;
  assign new_C3063_ = new_C3052_ | new_C3075_;
  assign new_C3064_ = new_C3074_ | new_C3073_;
  assign new_C3065_ = new_C3079_ & new_C3078_;
  assign new_C3066_ = new_C3077_ & new_C3076_;
  assign new_C3067_ = new_C3082_ | new_C3081_;
  assign new_C3068_ = new_C3077_ & new_C3080_;
  assign new_C3069_ = new_C3052_ | new_C3085_;
  assign new_C3070_ = new_C3084_ | new_C3083_;
  assign new_C3071_ = new_C3087_ | new_C3086_;
  assign new_C3072_ = ~new_C3063_ & new_C3089_;
  assign new_C3073_ = ~new_C3065_ & new_C3077_;
  assign new_C3074_ = new_C3065_ & ~new_C3077_;
  assign new_C3075_ = new_C3051_ & ~new_C3052_;
  assign new_C3076_ = ~new_C3098_ | ~new_C3099_;
  assign new_C3077_ = new_C3091_ | new_C3093_;
  assign new_C3078_ = new_C3101_ | new_C3100_;
  assign new_C3079_ = new_C3095_ | new_C3094_;
  assign new_C3080_ = ~new_C3103_ | ~new_C3102_;
  assign new_C3081_ = ~new_C3104_ & new_C3105_;
  assign new_C3082_ = new_C3104_ & ~new_C3105_;
  assign new_C3083_ = ~new_C3051_ & new_C3052_;
  assign new_C3084_ = new_C3051_ & ~new_C3052_;
  assign new_C3085_ = ~new_C3067_ | new_C3077_;
  assign new_C3086_ = new_C3067_ & new_C3077_;
  assign new_C3087_ = ~new_C3067_ & ~new_C3077_;
  assign new_C3088_ = new_C3109_ | new_C3108_;
  assign new_C3089_ = new_C3055_ | new_C3088_;
  assign new_C3090_ = new_C3113_ | new_C3112_;
  assign new_C3091_ = ~new_C3055_ & new_C3090_;
  assign new_C3092_ = new_C3111_ | new_C3110_;
  assign new_C3093_ = new_C3055_ & new_C3092_;
  assign new_C3094_ = new_C3053_ & ~new_C3063_;
  assign new_C3095_ = ~new_C3053_ & new_C3063_;
  assign new_C3096_ = ~new_C3052_ | ~new_C3077_;
  assign new_C3097_ = new_C3063_ & new_C3096_;
  assign new_C3098_ = ~new_C3063_ & ~new_C3097_;
  assign new_C3099_ = new_C3063_ | new_C3096_;
  assign new_C3100_ = ~new_C3053_ & new_C3054_;
  assign new_C3101_ = new_C3053_ & ~new_C3054_;
  assign new_C3102_ = new_C3070_ | new_C3107_;
  assign new_C3103_ = ~new_C3070_ & ~new_C3106_;
  assign new_C3104_ = new_C3053_ | new_C3070_;
  assign new_C3105_ = new_C3053_ | new_C3054_;
  assign new_C3106_ = new_C3070_ & new_C3107_;
  assign new_C3107_ = ~new_C3052_ | ~new_C3077_;
  assign new_C3108_ = new_C3085_ & new_C3105_;
  assign new_C3109_ = ~new_C3085_ & ~new_C3105_;
  assign new_C3110_ = new_C3114_ | new_C3115_;
  assign new_C3111_ = ~new_C3056_ & new_C3070_;
  assign new_C3112_ = new_C3116_ | new_C3117_;
  assign new_C3113_ = new_C3056_ & new_C3070_;
  assign new_C3114_ = ~new_C3056_ & ~new_C3070_;
  assign new_C3115_ = new_C3056_ & ~new_C3070_;
  assign new_C3116_ = new_C3056_ & ~new_C3070_;
  assign new_C3117_ = ~new_C3056_ & new_C3070_;
  assign new_C3118_ = new_E613_;
  assign new_C3119_ = new_E680_;
  assign new_C3120_ = new_E747_;
  assign new_C3121_ = new_E814_;
  assign new_C3122_ = new_E881_;
  assign new_C3123_ = new_E948_;
  assign new_C3124_ = new_C3131_ & new_C3130_;
  assign new_C3125_ = new_C3133_ | new_C3132_;
  assign new_C3126_ = new_C3135_ | new_C3134_;
  assign new_C3127_ = new_C3137_ & new_C3136_;
  assign new_C3128_ = new_C3137_ & new_C3138_;
  assign new_C3129_ = new_C3130_ | new_C3139_;
  assign new_C3130_ = new_C3119_ | new_C3142_;
  assign new_C3131_ = new_C3141_ | new_C3140_;
  assign new_C3132_ = new_C3146_ & new_C3145_;
  assign new_C3133_ = new_C3144_ & new_C3143_;
  assign new_C3134_ = new_C3149_ | new_C3148_;
  assign new_C3135_ = new_C3144_ & new_C3147_;
  assign new_C3136_ = new_C3119_ | new_C3152_;
  assign new_C3137_ = new_C3151_ | new_C3150_;
  assign new_C3138_ = new_C3154_ | new_C3153_;
  assign new_C3139_ = ~new_C3130_ & new_C3156_;
  assign new_C3140_ = ~new_C3132_ & new_C3144_;
  assign new_C3141_ = new_C3132_ & ~new_C3144_;
  assign new_C3142_ = new_C3118_ & ~new_C3119_;
  assign new_C3143_ = ~new_C3165_ | ~new_C3166_;
  assign new_C3144_ = new_C3158_ | new_C3160_;
  assign new_C3145_ = new_C3168_ | new_C3167_;
  assign new_C3146_ = new_C3162_ | new_C3161_;
  assign new_C3147_ = ~new_C3170_ | ~new_C3169_;
  assign new_C3148_ = ~new_C3171_ & new_C3172_;
  assign new_C3149_ = new_C3171_ & ~new_C3172_;
  assign new_C3150_ = ~new_C3118_ & new_C3119_;
  assign new_C3151_ = new_C3118_ & ~new_C3119_;
  assign new_C3152_ = ~new_C3134_ | new_C3144_;
  assign new_C3153_ = new_C3134_ & new_C3144_;
  assign new_C3154_ = ~new_C3134_ & ~new_C3144_;
  assign new_C3155_ = new_C3176_ | new_C3175_;
  assign new_C3156_ = new_C3122_ | new_C3155_;
  assign new_C3157_ = new_C3180_ | new_C3179_;
  assign new_C3158_ = ~new_C3122_ & new_C3157_;
  assign new_C3159_ = new_C3178_ | new_C3177_;
  assign new_C3160_ = new_C3122_ & new_C3159_;
  assign new_C3161_ = new_C3120_ & ~new_C3130_;
  assign new_C3162_ = ~new_C3120_ & new_C3130_;
  assign new_C3163_ = ~new_C3119_ | ~new_C3144_;
  assign new_C3164_ = new_C3130_ & new_C3163_;
  assign new_C3165_ = ~new_C3130_ & ~new_C3164_;
  assign new_C3166_ = new_C3130_ | new_C3163_;
  assign new_C3167_ = ~new_C3120_ & new_C3121_;
  assign new_C3168_ = new_C3120_ & ~new_C3121_;
  assign new_C3169_ = new_C3137_ | new_C3174_;
  assign new_C3170_ = ~new_C3137_ & ~new_C3173_;
  assign new_C3171_ = new_C3120_ | new_C3137_;
  assign new_C3172_ = new_C3120_ | new_C3121_;
  assign new_C3173_ = new_C3137_ & new_C3174_;
  assign new_C3174_ = ~new_C3119_ | ~new_C3144_;
  assign new_C3175_ = new_C3152_ & new_C3172_;
  assign new_C3176_ = ~new_C3152_ & ~new_C3172_;
  assign new_C3177_ = new_C3181_ | new_C3182_;
  assign new_C3178_ = ~new_C3123_ & new_C3137_;
  assign new_C3179_ = new_C3183_ | new_C3184_;
  assign new_C3180_ = new_C3123_ & new_C3137_;
  assign new_C3181_ = ~new_C3123_ & ~new_C3137_;
  assign new_C3182_ = new_C3123_ & ~new_C3137_;
  assign new_C3183_ = new_C3123_ & ~new_C3137_;
  assign new_C3184_ = ~new_C3123_ & new_C3137_;
  assign new_C3185_ = new_E1015_;
  assign new_C3186_ = new_E1082_;
  assign new_C3187_ = new_E1149_;
  assign new_C3188_ = new_E1216_;
  assign new_C3189_ = new_E1283_;
  assign new_C3190_ = new_E1350_;
  assign new_C3191_ = new_C3198_ & new_C3197_;
  assign new_C3192_ = new_C3200_ | new_C3199_;
  assign new_C3193_ = new_C3202_ | new_C3201_;
  assign new_C3194_ = new_C3204_ & new_C3203_;
  assign new_C3195_ = new_C3204_ & new_C3205_;
  assign new_C3196_ = new_C3197_ | new_C3206_;
  assign new_C3197_ = new_C3186_ | new_C3209_;
  assign new_C3198_ = new_C3208_ | new_C3207_;
  assign new_C3199_ = new_C3213_ & new_C3212_;
  assign new_C3200_ = new_C3211_ & new_C3210_;
  assign new_C3201_ = new_C3216_ | new_C3215_;
  assign new_C3202_ = new_C3211_ & new_C3214_;
  assign new_C3203_ = new_C3186_ | new_C3219_;
  assign new_C3204_ = new_C3218_ | new_C3217_;
  assign new_C3205_ = new_C3221_ | new_C3220_;
  assign new_C3206_ = ~new_C3197_ & new_C3223_;
  assign new_C3207_ = ~new_C3199_ & new_C3211_;
  assign new_C3208_ = new_C3199_ & ~new_C3211_;
  assign new_C3209_ = new_C3185_ & ~new_C3186_;
  assign new_C3210_ = ~new_C3232_ | ~new_C3233_;
  assign new_C3211_ = new_C3225_ | new_C3227_;
  assign new_C3212_ = new_C3235_ | new_C3234_;
  assign new_C3213_ = new_C3229_ | new_C3228_;
  assign new_C3214_ = ~new_C3237_ | ~new_C3236_;
  assign new_C3215_ = ~new_C3238_ & new_C3239_;
  assign new_C3216_ = new_C3238_ & ~new_C3239_;
  assign new_C3217_ = ~new_C3185_ & new_C3186_;
  assign new_C3218_ = new_C3185_ & ~new_C3186_;
  assign new_C3219_ = ~new_C3201_ | new_C3211_;
  assign new_C3220_ = new_C3201_ & new_C3211_;
  assign new_C3221_ = ~new_C3201_ & ~new_C3211_;
  assign new_C3222_ = new_C3243_ | new_C3242_;
  assign new_C3223_ = new_C3189_ | new_C3222_;
  assign new_C3224_ = new_C3247_ | new_C3246_;
  assign new_C3225_ = ~new_C3189_ & new_C3224_;
  assign new_C3226_ = new_C3245_ | new_C3244_;
  assign new_C3227_ = new_C3189_ & new_C3226_;
  assign new_C3228_ = new_C3187_ & ~new_C3197_;
  assign new_C3229_ = ~new_C3187_ & new_C3197_;
  assign new_C3230_ = ~new_C3186_ | ~new_C3211_;
  assign new_C3231_ = new_C3197_ & new_C3230_;
  assign new_C3232_ = ~new_C3197_ & ~new_C3231_;
  assign new_C3233_ = new_C3197_ | new_C3230_;
  assign new_C3234_ = ~new_C3187_ & new_C3188_;
  assign new_C3235_ = new_C3187_ & ~new_C3188_;
  assign new_C3236_ = new_C3204_ | new_C3241_;
  assign new_C3237_ = ~new_C3204_ & ~new_C3240_;
  assign new_C3238_ = new_C3187_ | new_C3204_;
  assign new_C3239_ = new_C3187_ | new_C3188_;
  assign new_C3240_ = new_C3204_ & new_C3241_;
  assign new_C3241_ = ~new_C3186_ | ~new_C3211_;
  assign new_C3242_ = new_C3219_ & new_C3239_;
  assign new_C3243_ = ~new_C3219_ & ~new_C3239_;
  assign new_C3244_ = new_C3248_ | new_C3249_;
  assign new_C3245_ = ~new_C3190_ & new_C3204_;
  assign new_C3246_ = new_C3250_ | new_C3251_;
  assign new_C3247_ = new_C3190_ & new_C3204_;
  assign new_C3248_ = ~new_C3190_ & ~new_C3204_;
  assign new_C3249_ = new_C3190_ & ~new_C3204_;
  assign new_C3250_ = new_C3190_ & ~new_C3204_;
  assign new_C3251_ = ~new_C3190_ & new_C3204_;
  assign new_C3252_ = new_E1417_;
  assign new_C3253_ = new_E1484_;
  assign new_C3254_ = new_E1551_;
  assign new_C3255_ = new_E1618_;
  assign new_C3256_ = new_E1685_;
  assign new_C3257_ = new_E1752_;
  assign new_C3258_ = new_C3265_ & new_C3264_;
  assign new_C3259_ = new_C3267_ | new_C3266_;
  assign new_C3260_ = new_C3269_ | new_C3268_;
  assign new_C3261_ = new_C3271_ & new_C3270_;
  assign new_C3262_ = new_C3271_ & new_C3272_;
  assign new_C3263_ = new_C3264_ | new_C3273_;
  assign new_C3264_ = new_C3253_ | new_C3276_;
  assign new_C3265_ = new_C3275_ | new_C3274_;
  assign new_C3266_ = new_C3280_ & new_C3279_;
  assign new_C3267_ = new_C3278_ & new_C3277_;
  assign new_C3268_ = new_C3283_ | new_C3282_;
  assign new_C3269_ = new_C3278_ & new_C3281_;
  assign new_C3270_ = new_C3253_ | new_C3286_;
  assign new_C3271_ = new_C3285_ | new_C3284_;
  assign new_C3272_ = new_C3288_ | new_C3287_;
  assign new_C3273_ = ~new_C3264_ & new_C3290_;
  assign new_C3274_ = ~new_C3266_ & new_C3278_;
  assign new_C3275_ = new_C3266_ & ~new_C3278_;
  assign new_C3276_ = new_C3252_ & ~new_C3253_;
  assign new_C3277_ = ~new_C3299_ | ~new_C3300_;
  assign new_C3278_ = new_C3292_ | new_C3294_;
  assign new_C3279_ = new_C3302_ | new_C3301_;
  assign new_C3280_ = new_C3296_ | new_C3295_;
  assign new_C3281_ = ~new_C3304_ | ~new_C3303_;
  assign new_C3282_ = ~new_C3305_ & new_C3306_;
  assign new_C3283_ = new_C3305_ & ~new_C3306_;
  assign new_C3284_ = ~new_C3252_ & new_C3253_;
  assign new_C3285_ = new_C3252_ & ~new_C3253_;
  assign new_C3286_ = ~new_C3268_ | new_C3278_;
  assign new_C3287_ = new_C3268_ & new_C3278_;
  assign new_C3288_ = ~new_C3268_ & ~new_C3278_;
  assign new_C3289_ = new_C3310_ | new_C3309_;
  assign new_C3290_ = new_C3256_ | new_C3289_;
  assign new_C3291_ = new_C3314_ | new_C3313_;
  assign new_C3292_ = ~new_C3256_ & new_C3291_;
  assign new_C3293_ = new_C3312_ | new_C3311_;
  assign new_C3294_ = new_C3256_ & new_C3293_;
  assign new_C3295_ = new_C3254_ & ~new_C3264_;
  assign new_C3296_ = ~new_C3254_ & new_C3264_;
  assign new_C3297_ = ~new_C3253_ | ~new_C3278_;
  assign new_C3298_ = new_C3264_ & new_C3297_;
  assign new_C3299_ = ~new_C3264_ & ~new_C3298_;
  assign new_C3300_ = new_C3264_ | new_C3297_;
  assign new_C3301_ = ~new_C3254_ & new_C3255_;
  assign new_C3302_ = new_C3254_ & ~new_C3255_;
  assign new_C3303_ = new_C3271_ | new_C3308_;
  assign new_C3304_ = ~new_C3271_ & ~new_C3307_;
  assign new_C3305_ = new_C3254_ | new_C3271_;
  assign new_C3306_ = new_C3254_ | new_C3255_;
  assign new_C3307_ = new_C3271_ & new_C3308_;
  assign new_C3308_ = ~new_C3253_ | ~new_C3278_;
  assign new_C3309_ = new_C3286_ & new_C3306_;
  assign new_C3310_ = ~new_C3286_ & ~new_C3306_;
  assign new_C3311_ = new_C3315_ | new_C3316_;
  assign new_C3312_ = ~new_C3257_ & new_C3271_;
  assign new_C3313_ = new_C3317_ | new_C3318_;
  assign new_C3314_ = new_C3257_ & new_C3271_;
  assign new_C3315_ = ~new_C3257_ & ~new_C3271_;
  assign new_C3316_ = new_C3257_ & ~new_C3271_;
  assign new_C3317_ = new_C3257_ & ~new_C3271_;
  assign new_C3318_ = ~new_C3257_ & new_C3271_;
  assign new_C3319_ = new_E1819_;
  assign new_C3320_ = new_E1886_;
  assign new_C3321_ = new_E1953_;
  assign new_C3322_ = new_E2020_;
  assign new_C3323_ = new_E2087_;
  assign new_C3324_ = new_E2154_;
  assign new_C3325_ = new_C3332_ & new_C3331_;
  assign new_C3326_ = new_C3334_ | new_C3333_;
  assign new_C3327_ = new_C3336_ | new_C3335_;
  assign new_C3328_ = new_C3338_ & new_C3337_;
  assign new_C3329_ = new_C3338_ & new_C3339_;
  assign new_C3330_ = new_C3331_ | new_C3340_;
  assign new_C3331_ = new_C3320_ | new_C3343_;
  assign new_C3332_ = new_C3342_ | new_C3341_;
  assign new_C3333_ = new_C3347_ & new_C3346_;
  assign new_C3334_ = new_C3345_ & new_C3344_;
  assign new_C3335_ = new_C3350_ | new_C3349_;
  assign new_C3336_ = new_C3345_ & new_C3348_;
  assign new_C3337_ = new_C3320_ | new_C3353_;
  assign new_C3338_ = new_C3352_ | new_C3351_;
  assign new_C3339_ = new_C3355_ | new_C3354_;
  assign new_C3340_ = ~new_C3331_ & new_C3357_;
  assign new_C3341_ = ~new_C3333_ & new_C3345_;
  assign new_C3342_ = new_C3333_ & ~new_C3345_;
  assign new_C3343_ = new_C3319_ & ~new_C3320_;
  assign new_C3344_ = ~new_C3366_ | ~new_C3367_;
  assign new_C3345_ = new_C3359_ | new_C3361_;
  assign new_C3346_ = new_C3369_ | new_C3368_;
  assign new_C3347_ = new_C3363_ | new_C3362_;
  assign new_C3348_ = ~new_C3371_ | ~new_C3370_;
  assign new_C3349_ = ~new_C3372_ & new_C3373_;
  assign new_C3350_ = new_C3372_ & ~new_C3373_;
  assign new_C3351_ = ~new_C3319_ & new_C3320_;
  assign new_C3352_ = new_C3319_ & ~new_C3320_;
  assign new_C3353_ = ~new_C3335_ | new_C3345_;
  assign new_C3354_ = new_C3335_ & new_C3345_;
  assign new_C3355_ = ~new_C3335_ & ~new_C3345_;
  assign new_C3356_ = new_C3377_ | new_C3376_;
  assign new_C3357_ = new_C3323_ | new_C3356_;
  assign new_C3358_ = new_C3381_ | new_C3380_;
  assign new_C3359_ = ~new_C3323_ & new_C3358_;
  assign new_C3360_ = new_C3379_ | new_C3378_;
  assign new_C3361_ = new_C3323_ & new_C3360_;
  assign new_C3362_ = new_C3321_ & ~new_C3331_;
  assign new_C3363_ = ~new_C3321_ & new_C3331_;
  assign new_C3364_ = ~new_C3320_ | ~new_C3345_;
  assign new_C3365_ = new_C3331_ & new_C3364_;
  assign new_C3366_ = ~new_C3331_ & ~new_C3365_;
  assign new_C3367_ = new_C3331_ | new_C3364_;
  assign new_C3368_ = ~new_C3321_ & new_C3322_;
  assign new_C3369_ = new_C3321_ & ~new_C3322_;
  assign new_C3370_ = new_C3338_ | new_C3375_;
  assign new_C3371_ = ~new_C3338_ & ~new_C3374_;
  assign new_C3372_ = new_C3321_ | new_C3338_;
  assign new_C3373_ = new_C3321_ | new_C3322_;
  assign new_C3374_ = new_C3338_ & new_C3375_;
  assign new_C3375_ = ~new_C3320_ | ~new_C3345_;
  assign new_C3376_ = new_C3353_ & new_C3373_;
  assign new_C3377_ = ~new_C3353_ & ~new_C3373_;
  assign new_C3378_ = new_C3382_ | new_C3383_;
  assign new_C3379_ = ~new_C3324_ & new_C3338_;
  assign new_C3380_ = new_C3384_ | new_C3385_;
  assign new_C3381_ = new_C3324_ & new_C3338_;
  assign new_C3382_ = ~new_C3324_ & ~new_C3338_;
  assign new_C3383_ = new_C3324_ & ~new_C3338_;
  assign new_C3384_ = new_C3324_ & ~new_C3338_;
  assign new_C3385_ = ~new_C3324_ & new_C3338_;
  assign new_C3386_ = new_E2221_;
  assign new_C3387_ = new_E2288_;
  assign new_C3388_ = new_E2355_;
  assign new_C3389_ = new_E2422_;
  assign new_C3390_ = new_E2489_;
  assign new_C3391_ = new_E2556_;
  assign new_C3392_ = new_C3399_ & new_C3398_;
  assign new_C3393_ = new_C3401_ | new_C3400_;
  assign new_C3394_ = new_C3403_ | new_C3402_;
  assign new_C3395_ = new_C3405_ & new_C3404_;
  assign new_C3396_ = new_C3405_ & new_C3406_;
  assign new_C3397_ = new_C3398_ | new_C3407_;
  assign new_C3398_ = new_C3387_ | new_C3410_;
  assign new_C3399_ = new_C3409_ | new_C3408_;
  assign new_C3400_ = new_C3414_ & new_C3413_;
  assign new_C3401_ = new_C3412_ & new_C3411_;
  assign new_C3402_ = new_C3417_ | new_C3416_;
  assign new_C3403_ = new_C3412_ & new_C3415_;
  assign new_C3404_ = new_C3387_ | new_C3420_;
  assign new_C3405_ = new_C3419_ | new_C3418_;
  assign new_C3406_ = new_C3422_ | new_C3421_;
  assign new_C3407_ = ~new_C3398_ & new_C3424_;
  assign new_C3408_ = ~new_C3400_ & new_C3412_;
  assign new_C3409_ = new_C3400_ & ~new_C3412_;
  assign new_C3410_ = new_C3386_ & ~new_C3387_;
  assign new_C3411_ = ~new_C3433_ | ~new_C3434_;
  assign new_C3412_ = new_C3426_ | new_C3428_;
  assign new_C3413_ = new_C3436_ | new_C3435_;
  assign new_C3414_ = new_C3430_ | new_C3429_;
  assign new_C3415_ = ~new_C3438_ | ~new_C3437_;
  assign new_C3416_ = ~new_C3439_ & new_C3440_;
  assign new_C3417_ = new_C3439_ & ~new_C3440_;
  assign new_C3418_ = ~new_C3386_ & new_C3387_;
  assign new_C3419_ = new_C3386_ & ~new_C3387_;
  assign new_C3420_ = ~new_C3402_ | new_C3412_;
  assign new_C3421_ = new_C3402_ & new_C3412_;
  assign new_C3422_ = ~new_C3402_ & ~new_C3412_;
  assign new_C3423_ = new_C3444_ | new_C3443_;
  assign new_C3424_ = new_C3390_ | new_C3423_;
  assign new_C3425_ = new_C3448_ | new_C3447_;
  assign new_C3426_ = ~new_C3390_ & new_C3425_;
  assign new_C3427_ = new_C3446_ | new_C3445_;
  assign new_C3428_ = new_C3390_ & new_C3427_;
  assign new_C3429_ = new_C3388_ & ~new_C3398_;
  assign new_C3430_ = ~new_C3388_ & new_C3398_;
  assign new_C3431_ = ~new_C3387_ | ~new_C3412_;
  assign new_C3432_ = new_C3398_ & new_C3431_;
  assign new_C3433_ = ~new_C3398_ & ~new_C3432_;
  assign new_C3434_ = new_C3398_ | new_C3431_;
  assign new_C3435_ = ~new_C3388_ & new_C3389_;
  assign new_C3436_ = new_C3388_ & ~new_C3389_;
  assign new_C3437_ = new_C3405_ | new_C3442_;
  assign new_C3438_ = ~new_C3405_ & ~new_C3441_;
  assign new_C3439_ = new_C3388_ | new_C3405_;
  assign new_C3440_ = new_C3388_ | new_C3389_;
  assign new_C3441_ = new_C3405_ & new_C3442_;
  assign new_C3442_ = ~new_C3387_ | ~new_C3412_;
  assign new_C3443_ = new_C3420_ & new_C3440_;
  assign new_C3444_ = ~new_C3420_ & ~new_C3440_;
  assign new_C3445_ = new_C3449_ | new_C3450_;
  assign new_C3446_ = ~new_C3391_ & new_C3405_;
  assign new_C3447_ = new_C3451_ | new_C3452_;
  assign new_C3448_ = new_C3391_ & new_C3405_;
  assign new_C3449_ = ~new_C3391_ & ~new_C3405_;
  assign new_C3450_ = new_C3391_ & ~new_C3405_;
  assign new_C3451_ = new_C3391_ & ~new_C3405_;
  assign new_C3452_ = ~new_C3391_ & new_C3405_;
  assign new_C3453_ = new_E2623_;
  assign new_C3454_ = new_E2690_;
  assign new_C3455_ = new_E2757_;
  assign new_C3456_ = new_E2824_;
  assign new_C3457_ = new_E2891_;
  assign new_C3458_ = new_E2958_;
  assign new_C3459_ = new_C3466_ & new_C3465_;
  assign new_C3460_ = new_C3468_ | new_C3467_;
  assign new_C3461_ = new_C3470_ | new_C3469_;
  assign new_C3462_ = new_C3472_ & new_C3471_;
  assign new_C3463_ = new_C3472_ & new_C3473_;
  assign new_C3464_ = new_C3465_ | new_C3474_;
  assign new_C3465_ = new_C3454_ | new_C3477_;
  assign new_C3466_ = new_C3476_ | new_C3475_;
  assign new_C3467_ = new_C3481_ & new_C3480_;
  assign new_C3468_ = new_C3479_ & new_C3478_;
  assign new_C3469_ = new_C3484_ | new_C3483_;
  assign new_C3470_ = new_C3479_ & new_C3482_;
  assign new_C3471_ = new_C3454_ | new_C3487_;
  assign new_C3472_ = new_C3486_ | new_C3485_;
  assign new_C3473_ = new_C3489_ | new_C3488_;
  assign new_C3474_ = ~new_C3465_ & new_C3491_;
  assign new_C3475_ = ~new_C3467_ & new_C3479_;
  assign new_C3476_ = new_C3467_ & ~new_C3479_;
  assign new_C3477_ = new_C3453_ & ~new_C3454_;
  assign new_C3478_ = ~new_C3500_ | ~new_C3501_;
  assign new_C3479_ = new_C3493_ | new_C3495_;
  assign new_C3480_ = new_C3503_ | new_C3502_;
  assign new_C3481_ = new_C3497_ | new_C3496_;
  assign new_C3482_ = ~new_C3505_ | ~new_C3504_;
  assign new_C3483_ = ~new_C3506_ & new_C3507_;
  assign new_C3484_ = new_C3506_ & ~new_C3507_;
  assign new_C3485_ = ~new_C3453_ & new_C3454_;
  assign new_C3486_ = new_C3453_ & ~new_C3454_;
  assign new_C3487_ = ~new_C3469_ | new_C3479_;
  assign new_C3488_ = new_C3469_ & new_C3479_;
  assign new_C3489_ = ~new_C3469_ & ~new_C3479_;
  assign new_C3490_ = new_C3511_ | new_C3510_;
  assign new_C3491_ = new_C3457_ | new_C3490_;
  assign new_C3492_ = new_C3515_ | new_C3514_;
  assign new_C3493_ = ~new_C3457_ & new_C3492_;
  assign new_C3494_ = new_C3513_ | new_C3512_;
  assign new_C3495_ = new_C3457_ & new_C3494_;
  assign new_C3496_ = new_C3455_ & ~new_C3465_;
  assign new_C3497_ = ~new_C3455_ & new_C3465_;
  assign new_C3498_ = ~new_C3454_ | ~new_C3479_;
  assign new_C3499_ = new_C3465_ & new_C3498_;
  assign new_C3500_ = ~new_C3465_ & ~new_C3499_;
  assign new_C3501_ = new_C3465_ | new_C3498_;
  assign new_C3502_ = ~new_C3455_ & new_C3456_;
  assign new_C3503_ = new_C3455_ & ~new_C3456_;
  assign new_C3504_ = new_C3472_ | new_C3509_;
  assign new_C3505_ = ~new_C3472_ & ~new_C3508_;
  assign new_C3506_ = new_C3455_ | new_C3472_;
  assign new_C3507_ = new_C3455_ | new_C3456_;
  assign new_C3508_ = new_C3472_ & new_C3509_;
  assign new_C3509_ = ~new_C3454_ | ~new_C3479_;
  assign new_C3510_ = new_C3487_ & new_C3507_;
  assign new_C3511_ = ~new_C3487_ & ~new_C3507_;
  assign new_C3512_ = new_C3516_ | new_C3517_;
  assign new_C3513_ = ~new_C3458_ & new_C3472_;
  assign new_C3514_ = new_C3518_ | new_C3519_;
  assign new_C3515_ = new_C3458_ & new_C3472_;
  assign new_C3516_ = ~new_C3458_ & ~new_C3472_;
  assign new_C3517_ = new_C3458_ & ~new_C3472_;
  assign new_C3518_ = new_C3458_ & ~new_C3472_;
  assign new_C3519_ = ~new_C3458_ & new_C3472_;
  assign new_C3520_ = new_E3025_;
  assign new_C3521_ = new_E3092_;
  assign new_C3522_ = new_E3159_;
  assign new_C3523_ = new_E3226_;
  assign new_C3524_ = new_E3293_;
  assign new_C3525_ = new_E3360_;
  assign new_C3526_ = new_C3533_ & new_C3532_;
  assign new_C3527_ = new_C3535_ | new_C3534_;
  assign new_C3528_ = new_C3537_ | new_C3536_;
  assign new_C3529_ = new_C3539_ & new_C3538_;
  assign new_C3530_ = new_C3539_ & new_C3540_;
  assign new_C3531_ = new_C3532_ | new_C3541_;
  assign new_C3532_ = new_C3521_ | new_C3544_;
  assign new_C3533_ = new_C3543_ | new_C3542_;
  assign new_C3534_ = new_C3548_ & new_C3547_;
  assign new_C3535_ = new_C3546_ & new_C3545_;
  assign new_C3536_ = new_C3551_ | new_C3550_;
  assign new_C3537_ = new_C3546_ & new_C3549_;
  assign new_C3538_ = new_C3521_ | new_C3554_;
  assign new_C3539_ = new_C3553_ | new_C3552_;
  assign new_C3540_ = new_C3556_ | new_C3555_;
  assign new_C3541_ = ~new_C3532_ & new_C3558_;
  assign new_C3542_ = ~new_C3534_ & new_C3546_;
  assign new_C3543_ = new_C3534_ & ~new_C3546_;
  assign new_C3544_ = new_C3520_ & ~new_C3521_;
  assign new_C3545_ = ~new_C3567_ | ~new_C3568_;
  assign new_C3546_ = new_C3560_ | new_C3562_;
  assign new_C3547_ = new_C3570_ | new_C3569_;
  assign new_C3548_ = new_C3564_ | new_C3563_;
  assign new_C3549_ = ~new_C3572_ | ~new_C3571_;
  assign new_C3550_ = ~new_C3573_ & new_C3574_;
  assign new_C3551_ = new_C3573_ & ~new_C3574_;
  assign new_C3552_ = ~new_C3520_ & new_C3521_;
  assign new_C3553_ = new_C3520_ & ~new_C3521_;
  assign new_C3554_ = ~new_C3536_ | new_C3546_;
  assign new_C3555_ = new_C3536_ & new_C3546_;
  assign new_C3556_ = ~new_C3536_ & ~new_C3546_;
  assign new_C3557_ = new_C3578_ | new_C3577_;
  assign new_C3558_ = new_C3524_ | new_C3557_;
  assign new_C3559_ = new_C3582_ | new_C3581_;
  assign new_C3560_ = ~new_C3524_ & new_C3559_;
  assign new_C3561_ = new_C3580_ | new_C3579_;
  assign new_C3562_ = new_C3524_ & new_C3561_;
  assign new_C3563_ = new_C3522_ & ~new_C3532_;
  assign new_C3564_ = ~new_C3522_ & new_C3532_;
  assign new_C3565_ = ~new_C3521_ | ~new_C3546_;
  assign new_C3566_ = new_C3532_ & new_C3565_;
  assign new_C3567_ = ~new_C3532_ & ~new_C3566_;
  assign new_C3568_ = new_C3532_ | new_C3565_;
  assign new_C3569_ = ~new_C3522_ & new_C3523_;
  assign new_C3570_ = new_C3522_ & ~new_C3523_;
  assign new_C3571_ = new_C3539_ | new_C3576_;
  assign new_C3572_ = ~new_C3539_ & ~new_C3575_;
  assign new_C3573_ = new_C3522_ | new_C3539_;
  assign new_C3574_ = new_C3522_ | new_C3523_;
  assign new_C3575_ = new_C3539_ & new_C3576_;
  assign new_C3576_ = ~new_C3521_ | ~new_C3546_;
  assign new_C3577_ = new_C3554_ & new_C3574_;
  assign new_C3578_ = ~new_C3554_ & ~new_C3574_;
  assign new_C3579_ = new_C3583_ | new_C3584_;
  assign new_C3580_ = ~new_C3525_ & new_C3539_;
  assign new_C3581_ = new_C3585_ | new_C3586_;
  assign new_C3582_ = new_C3525_ & new_C3539_;
  assign new_C3583_ = ~new_C3525_ & ~new_C3539_;
  assign new_C3584_ = new_C3525_ & ~new_C3539_;
  assign new_C3585_ = new_C3525_ & ~new_C3539_;
  assign new_C3586_ = ~new_C3525_ & new_C3539_;
  assign new_C3587_ = new_E3427_;
  assign new_C3588_ = new_E3494_;
  assign new_C3589_ = new_E3561_;
  assign new_C3590_ = new_E3628_;
  assign new_C3591_ = new_E3695_;
  assign new_C3592_ = new_E3762_;
  assign new_C3593_ = new_C3600_ & new_C3599_;
  assign new_C3594_ = new_C3602_ | new_C3601_;
  assign new_C3595_ = new_C3604_ | new_C3603_;
  assign new_C3596_ = new_C3606_ & new_C3605_;
  assign new_C3597_ = new_C3606_ & new_C3607_;
  assign new_C3598_ = new_C3599_ | new_C3608_;
  assign new_C3599_ = new_C3588_ | new_C3611_;
  assign new_C3600_ = new_C3610_ | new_C3609_;
  assign new_C3601_ = new_C3615_ & new_C3614_;
  assign new_C3602_ = new_C3613_ & new_C3612_;
  assign new_C3603_ = new_C3618_ | new_C3617_;
  assign new_C3604_ = new_C3613_ & new_C3616_;
  assign new_C3605_ = new_C3588_ | new_C3621_;
  assign new_C3606_ = new_C3620_ | new_C3619_;
  assign new_C3607_ = new_C3623_ | new_C3622_;
  assign new_C3608_ = ~new_C3599_ & new_C3625_;
  assign new_C3609_ = ~new_C3601_ & new_C3613_;
  assign new_C3610_ = new_C3601_ & ~new_C3613_;
  assign new_C3611_ = new_C3587_ & ~new_C3588_;
  assign new_C3612_ = ~new_C3634_ | ~new_C3635_;
  assign new_C3613_ = new_C3627_ | new_C3629_;
  assign new_C3614_ = new_C3637_ | new_C3636_;
  assign new_C3615_ = new_C3631_ | new_C3630_;
  assign new_C3616_ = ~new_C3639_ | ~new_C3638_;
  assign new_C3617_ = ~new_C3640_ & new_C3641_;
  assign new_C3618_ = new_C3640_ & ~new_C3641_;
  assign new_C3619_ = ~new_C3587_ & new_C3588_;
  assign new_C3620_ = new_C3587_ & ~new_C3588_;
  assign new_C3621_ = ~new_C3603_ | new_C3613_;
  assign new_C3622_ = new_C3603_ & new_C3613_;
  assign new_C3623_ = ~new_C3603_ & ~new_C3613_;
  assign new_C3624_ = new_C3645_ | new_C3644_;
  assign new_C3625_ = new_C3591_ | new_C3624_;
  assign new_C3626_ = new_C3649_ | new_C3648_;
  assign new_C3627_ = ~new_C3591_ & new_C3626_;
  assign new_C3628_ = new_C3647_ | new_C3646_;
  assign new_C3629_ = new_C3591_ & new_C3628_;
  assign new_C3630_ = new_C3589_ & ~new_C3599_;
  assign new_C3631_ = ~new_C3589_ & new_C3599_;
  assign new_C3632_ = ~new_C3588_ | ~new_C3613_;
  assign new_C3633_ = new_C3599_ & new_C3632_;
  assign new_C3634_ = ~new_C3599_ & ~new_C3633_;
  assign new_C3635_ = new_C3599_ | new_C3632_;
  assign new_C3636_ = ~new_C3589_ & new_C3590_;
  assign new_C3637_ = new_C3589_ & ~new_C3590_;
  assign new_C3638_ = new_C3606_ | new_C3643_;
  assign new_C3639_ = ~new_C3606_ & ~new_C3642_;
  assign new_C3640_ = new_C3589_ | new_C3606_;
  assign new_C3641_ = new_C3589_ | new_C3590_;
  assign new_C3642_ = new_C3606_ & new_C3643_;
  assign new_C3643_ = ~new_C3588_ | ~new_C3613_;
  assign new_C3644_ = new_C3621_ & new_C3641_;
  assign new_C3645_ = ~new_C3621_ & ~new_C3641_;
  assign new_C3646_ = new_C3650_ | new_C3651_;
  assign new_C3647_ = ~new_C3592_ & new_C3606_;
  assign new_C3648_ = new_C3652_ | new_C3653_;
  assign new_C3649_ = new_C3592_ & new_C3606_;
  assign new_C3650_ = ~new_C3592_ & ~new_C3606_;
  assign new_C3651_ = new_C3592_ & ~new_C3606_;
  assign new_C3652_ = new_C3592_ & ~new_C3606_;
  assign new_C3653_ = ~new_C3592_ & new_C3606_;
  assign new_C3654_ = new_E3829_;
  assign new_C3655_ = new_E3896_;
  assign new_C3656_ = new_E3963_;
  assign new_C3657_ = new_E4030_;
  assign new_C3658_ = new_E4097_;
  assign new_C3659_ = new_E4164_;
  assign new_C3660_ = new_C3667_ & new_C3666_;
  assign new_C3661_ = new_C3669_ | new_C3668_;
  assign new_C3662_ = new_C3671_ | new_C3670_;
  assign new_C3663_ = new_C3673_ & new_C3672_;
  assign new_C3664_ = new_C3673_ & new_C3674_;
  assign new_C3665_ = new_C3666_ | new_C3675_;
  assign new_C3666_ = new_C3655_ | new_C3678_;
  assign new_C3667_ = new_C3677_ | new_C3676_;
  assign new_C3668_ = new_C3682_ & new_C3681_;
  assign new_C3669_ = new_C3680_ & new_C3679_;
  assign new_C3670_ = new_C3685_ | new_C3684_;
  assign new_C3671_ = new_C3680_ & new_C3683_;
  assign new_C3672_ = new_C3655_ | new_C3688_;
  assign new_C3673_ = new_C3687_ | new_C3686_;
  assign new_C3674_ = new_C3690_ | new_C3689_;
  assign new_C3675_ = ~new_C3666_ & new_C3692_;
  assign new_C3676_ = ~new_C3668_ & new_C3680_;
  assign new_C3677_ = new_C3668_ & ~new_C3680_;
  assign new_C3678_ = new_C3654_ & ~new_C3655_;
  assign new_C3679_ = ~new_C3701_ | ~new_C3702_;
  assign new_C3680_ = new_C3694_ | new_C3696_;
  assign new_C3681_ = new_C3704_ | new_C3703_;
  assign new_C3682_ = new_C3698_ | new_C3697_;
  assign new_C3683_ = ~new_C3706_ | ~new_C3705_;
  assign new_C3684_ = ~new_C3707_ & new_C3708_;
  assign new_C3685_ = new_C3707_ & ~new_C3708_;
  assign new_C3686_ = ~new_C3654_ & new_C3655_;
  assign new_C3687_ = new_C3654_ & ~new_C3655_;
  assign new_C3688_ = ~new_C3670_ | new_C3680_;
  assign new_C3689_ = new_C3670_ & new_C3680_;
  assign new_C3690_ = ~new_C3670_ & ~new_C3680_;
  assign new_C3691_ = new_C3712_ | new_C3711_;
  assign new_C3692_ = new_C3658_ | new_C3691_;
  assign new_C3693_ = new_C3716_ | new_C3715_;
  assign new_C3694_ = ~new_C3658_ & new_C3693_;
  assign new_C3695_ = new_C3714_ | new_C3713_;
  assign new_C3696_ = new_C3658_ & new_C3695_;
  assign new_C3697_ = new_C3656_ & ~new_C3666_;
  assign new_C3698_ = ~new_C3656_ & new_C3666_;
  assign new_C3699_ = ~new_C3655_ | ~new_C3680_;
  assign new_C3700_ = new_C3666_ & new_C3699_;
  assign new_C3701_ = ~new_C3666_ & ~new_C3700_;
  assign new_C3702_ = new_C3666_ | new_C3699_;
  assign new_C3703_ = ~new_C3656_ & new_C3657_;
  assign new_C3704_ = new_C3656_ & ~new_C3657_;
  assign new_C3705_ = new_C3673_ | new_C3710_;
  assign new_C3706_ = ~new_C3673_ & ~new_C3709_;
  assign new_C3707_ = new_C3656_ | new_C3673_;
  assign new_C3708_ = new_C3656_ | new_C3657_;
  assign new_C3709_ = new_C3673_ & new_C3710_;
  assign new_C3710_ = ~new_C3655_ | ~new_C3680_;
  assign new_C3711_ = new_C3688_ & new_C3708_;
  assign new_C3712_ = ~new_C3688_ & ~new_C3708_;
  assign new_C3713_ = new_C3717_ | new_C3718_;
  assign new_C3714_ = ~new_C3659_ & new_C3673_;
  assign new_C3715_ = new_C3719_ | new_C3720_;
  assign new_C3716_ = new_C3659_ & new_C3673_;
  assign new_C3717_ = ~new_C3659_ & ~new_C3673_;
  assign new_C3718_ = new_C3659_ & ~new_C3673_;
  assign new_C3719_ = new_C3659_ & ~new_C3673_;
  assign new_C3720_ = ~new_C3659_ & new_C3673_;
  assign new_C3721_ = new_E4231_;
  assign new_C3722_ = new_E4298_;
  assign new_C3723_ = new_E4365_;
  assign new_C3724_ = new_E4432_;
  assign new_C3725_ = new_E4499_;
  assign new_C3726_ = new_E4566_;
  assign new_C3727_ = new_C3734_ & new_C3733_;
  assign new_C3728_ = new_C3736_ | new_C3735_;
  assign new_C3729_ = new_C3738_ | new_C3737_;
  assign new_C3730_ = new_C3740_ & new_C3739_;
  assign new_C3731_ = new_C3740_ & new_C3741_;
  assign new_C3732_ = new_C3733_ | new_C3742_;
  assign new_C3733_ = new_C3722_ | new_C3745_;
  assign new_C3734_ = new_C3744_ | new_C3743_;
  assign new_C3735_ = new_C3749_ & new_C3748_;
  assign new_C3736_ = new_C3747_ & new_C3746_;
  assign new_C3737_ = new_C3752_ | new_C3751_;
  assign new_C3738_ = new_C3747_ & new_C3750_;
  assign new_C3739_ = new_C3722_ | new_C3755_;
  assign new_C3740_ = new_C3754_ | new_C3753_;
  assign new_C3741_ = new_C3757_ | new_C3756_;
  assign new_C3742_ = ~new_C3733_ & new_C3759_;
  assign new_C3743_ = ~new_C3735_ & new_C3747_;
  assign new_C3744_ = new_C3735_ & ~new_C3747_;
  assign new_C3745_ = new_C3721_ & ~new_C3722_;
  assign new_C3746_ = ~new_C3768_ | ~new_C3769_;
  assign new_C3747_ = new_C3761_ | new_C3763_;
  assign new_C3748_ = new_C3771_ | new_C3770_;
  assign new_C3749_ = new_C3765_ | new_C3764_;
  assign new_C3750_ = ~new_C3773_ | ~new_C3772_;
  assign new_C3751_ = ~new_C3774_ & new_C3775_;
  assign new_C3752_ = new_C3774_ & ~new_C3775_;
  assign new_C3753_ = ~new_C3721_ & new_C3722_;
  assign new_C3754_ = new_C3721_ & ~new_C3722_;
  assign new_C3755_ = ~new_C3737_ | new_C3747_;
  assign new_C3756_ = new_C3737_ & new_C3747_;
  assign new_C3757_ = ~new_C3737_ & ~new_C3747_;
  assign new_C3758_ = new_C3779_ | new_C3778_;
  assign new_C3759_ = new_C3725_ | new_C3758_;
  assign new_C3760_ = new_C3783_ | new_C3782_;
  assign new_C3761_ = ~new_C3725_ & new_C3760_;
  assign new_C3762_ = new_C3781_ | new_C3780_;
  assign new_C3763_ = new_C3725_ & new_C3762_;
  assign new_C3764_ = new_C3723_ & ~new_C3733_;
  assign new_C3765_ = ~new_C3723_ & new_C3733_;
  assign new_C3766_ = ~new_C3722_ | ~new_C3747_;
  assign new_C3767_ = new_C3733_ & new_C3766_;
  assign new_C3768_ = ~new_C3733_ & ~new_C3767_;
  assign new_C3769_ = new_C3733_ | new_C3766_;
  assign new_C3770_ = ~new_C3723_ & new_C3724_;
  assign new_C3771_ = new_C3723_ & ~new_C3724_;
  assign new_C3772_ = new_C3740_ | new_C3777_;
  assign new_C3773_ = ~new_C3740_ & ~new_C3776_;
  assign new_C3774_ = new_C3723_ | new_C3740_;
  assign new_C3775_ = new_C3723_ | new_C3724_;
  assign new_C3776_ = new_C3740_ & new_C3777_;
  assign new_C3777_ = ~new_C3722_ | ~new_C3747_;
  assign new_C3778_ = new_C3755_ & new_C3775_;
  assign new_C3779_ = ~new_C3755_ & ~new_C3775_;
  assign new_C3780_ = new_C3784_ | new_C3785_;
  assign new_C3781_ = ~new_C3726_ & new_C3740_;
  assign new_C3782_ = new_C3786_ | new_C3787_;
  assign new_C3783_ = new_C3726_ & new_C3740_;
  assign new_C3784_ = ~new_C3726_ & ~new_C3740_;
  assign new_C3785_ = new_C3726_ & ~new_C3740_;
  assign new_C3786_ = new_C3726_ & ~new_C3740_;
  assign new_C3787_ = ~new_C3726_ & new_C3740_;
  assign new_C3788_ = new_E4633_;
  assign new_C3789_ = new_E4700_;
  assign new_C3790_ = new_E4767_;
  assign new_C3791_ = new_E4834_;
  assign new_C3792_ = new_E4901_;
  assign new_C3793_ = new_E4968_;
  assign new_C3794_ = new_C3801_ & new_C3800_;
  assign new_C3795_ = new_C3803_ | new_C3802_;
  assign new_C3796_ = new_C3805_ | new_C3804_;
  assign new_C3797_ = new_C3807_ & new_C3806_;
  assign new_C3798_ = new_C3807_ & new_C3808_;
  assign new_C3799_ = new_C3800_ | new_C3809_;
  assign new_C3800_ = new_C3789_ | new_C3812_;
  assign new_C3801_ = new_C3811_ | new_C3810_;
  assign new_C3802_ = new_C3816_ & new_C3815_;
  assign new_C3803_ = new_C3814_ & new_C3813_;
  assign new_C3804_ = new_C3819_ | new_C3818_;
  assign new_C3805_ = new_C3814_ & new_C3817_;
  assign new_C3806_ = new_C3789_ | new_C3822_;
  assign new_C3807_ = new_C3821_ | new_C3820_;
  assign new_C3808_ = new_C3824_ | new_C3823_;
  assign new_C3809_ = ~new_C3800_ & new_C3826_;
  assign new_C3810_ = ~new_C3802_ & new_C3814_;
  assign new_C3811_ = new_C3802_ & ~new_C3814_;
  assign new_C3812_ = new_C3788_ & ~new_C3789_;
  assign new_C3813_ = ~new_C3835_ | ~new_C3836_;
  assign new_C3814_ = new_C3828_ | new_C3830_;
  assign new_C3815_ = new_C3838_ | new_C3837_;
  assign new_C3816_ = new_C3832_ | new_C3831_;
  assign new_C3817_ = ~new_C3840_ | ~new_C3839_;
  assign new_C3818_ = ~new_C3841_ & new_C3842_;
  assign new_C3819_ = new_C3841_ & ~new_C3842_;
  assign new_C3820_ = ~new_C3788_ & new_C3789_;
  assign new_C3821_ = new_C3788_ & ~new_C3789_;
  assign new_C3822_ = ~new_C3804_ | new_C3814_;
  assign new_C3823_ = new_C3804_ & new_C3814_;
  assign new_C3824_ = ~new_C3804_ & ~new_C3814_;
  assign new_C3825_ = new_C3846_ | new_C3845_;
  assign new_C3826_ = new_C3792_ | new_C3825_;
  assign new_C3827_ = new_C3850_ | new_C3849_;
  assign new_C3828_ = ~new_C3792_ & new_C3827_;
  assign new_C3829_ = new_C3848_ | new_C3847_;
  assign new_C3830_ = new_C3792_ & new_C3829_;
  assign new_C3831_ = new_C3790_ & ~new_C3800_;
  assign new_C3832_ = ~new_C3790_ & new_C3800_;
  assign new_C3833_ = ~new_C3789_ | ~new_C3814_;
  assign new_C3834_ = new_C3800_ & new_C3833_;
  assign new_C3835_ = ~new_C3800_ & ~new_C3834_;
  assign new_C3836_ = new_C3800_ | new_C3833_;
  assign new_C3837_ = ~new_C3790_ & new_C3791_;
  assign new_C3838_ = new_C3790_ & ~new_C3791_;
  assign new_C3839_ = new_C3807_ | new_C3844_;
  assign new_C3840_ = ~new_C3807_ & ~new_C3843_;
  assign new_C3841_ = new_C3790_ | new_C3807_;
  assign new_C3842_ = new_C3790_ | new_C3791_;
  assign new_C3843_ = new_C3807_ & new_C3844_;
  assign new_C3844_ = ~new_C3789_ | ~new_C3814_;
  assign new_C3845_ = new_C3822_ & new_C3842_;
  assign new_C3846_ = ~new_C3822_ & ~new_C3842_;
  assign new_C3847_ = new_C3851_ | new_C3852_;
  assign new_C3848_ = ~new_C3793_ & new_C3807_;
  assign new_C3849_ = new_C3853_ | new_C3854_;
  assign new_C3850_ = new_C3793_ & new_C3807_;
  assign new_C3851_ = ~new_C3793_ & ~new_C3807_;
  assign new_C3852_ = new_C3793_ & ~new_C3807_;
  assign new_C3853_ = new_C3793_ & ~new_C3807_;
  assign new_C3854_ = ~new_C3793_ & new_C3807_;
  assign new_C3855_ = new_E5035_;
  assign new_C3856_ = new_E5102_;
  assign new_C3857_ = new_E5169_;
  assign new_C3858_ = new_E5236_;
  assign new_C3859_ = new_E5303_;
  assign new_C3860_ = new_E5370_;
  assign new_C3861_ = new_C3868_ & new_C3867_;
  assign new_C3862_ = new_C3870_ | new_C3869_;
  assign new_C3863_ = new_C3872_ | new_C3871_;
  assign new_C3864_ = new_C3874_ & new_C3873_;
  assign new_C3865_ = new_C3874_ & new_C3875_;
  assign new_C3866_ = new_C3867_ | new_C3876_;
  assign new_C3867_ = new_C3856_ | new_C3879_;
  assign new_C3868_ = new_C3878_ | new_C3877_;
  assign new_C3869_ = new_C3883_ & new_C3882_;
  assign new_C3870_ = new_C3881_ & new_C3880_;
  assign new_C3871_ = new_C3886_ | new_C3885_;
  assign new_C3872_ = new_C3881_ & new_C3884_;
  assign new_C3873_ = new_C3856_ | new_C3889_;
  assign new_C3874_ = new_C3888_ | new_C3887_;
  assign new_C3875_ = new_C3891_ | new_C3890_;
  assign new_C3876_ = ~new_C3867_ & new_C3893_;
  assign new_C3877_ = ~new_C3869_ & new_C3881_;
  assign new_C3878_ = new_C3869_ & ~new_C3881_;
  assign new_C3879_ = new_C3855_ & ~new_C3856_;
  assign new_C3880_ = ~new_C3902_ | ~new_C3903_;
  assign new_C3881_ = new_C3895_ | new_C3897_;
  assign new_C3882_ = new_C3905_ | new_C3904_;
  assign new_C3883_ = new_C3899_ | new_C3898_;
  assign new_C3884_ = ~new_C3907_ | ~new_C3906_;
  assign new_C3885_ = ~new_C3908_ & new_C3909_;
  assign new_C3886_ = new_C3908_ & ~new_C3909_;
  assign new_C3887_ = ~new_C3855_ & new_C3856_;
  assign new_C3888_ = new_C3855_ & ~new_C3856_;
  assign new_C3889_ = ~new_C3871_ | new_C3881_;
  assign new_C3890_ = new_C3871_ & new_C3881_;
  assign new_C3891_ = ~new_C3871_ & ~new_C3881_;
  assign new_C3892_ = new_C3913_ | new_C3912_;
  assign new_C3893_ = new_C3859_ | new_C3892_;
  assign new_C3894_ = new_C3917_ | new_C3916_;
  assign new_C3895_ = ~new_C3859_ & new_C3894_;
  assign new_C3896_ = new_C3915_ | new_C3914_;
  assign new_C3897_ = new_C3859_ & new_C3896_;
  assign new_C3898_ = new_C3857_ & ~new_C3867_;
  assign new_C3899_ = ~new_C3857_ & new_C3867_;
  assign new_C3900_ = ~new_C3856_ | ~new_C3881_;
  assign new_C3901_ = new_C3867_ & new_C3900_;
  assign new_C3902_ = ~new_C3867_ & ~new_C3901_;
  assign new_C3903_ = new_C3867_ | new_C3900_;
  assign new_C3904_ = ~new_C3857_ & new_C3858_;
  assign new_C3905_ = new_C3857_ & ~new_C3858_;
  assign new_C3906_ = new_C3874_ | new_C3911_;
  assign new_C3907_ = ~new_C3874_ & ~new_C3910_;
  assign new_C3908_ = new_C3857_ | new_C3874_;
  assign new_C3909_ = new_C3857_ | new_C3858_;
  assign new_C3910_ = new_C3874_ & new_C3911_;
  assign new_C3911_ = ~new_C3856_ | ~new_C3881_;
  assign new_C3912_ = new_C3889_ & new_C3909_;
  assign new_C3913_ = ~new_C3889_ & ~new_C3909_;
  assign new_C3914_ = new_C3918_ | new_C3919_;
  assign new_C3915_ = ~new_C3860_ & new_C3874_;
  assign new_C3916_ = new_C3920_ | new_C3921_;
  assign new_C3917_ = new_C3860_ & new_C3874_;
  assign new_C3918_ = ~new_C3860_ & ~new_C3874_;
  assign new_C3919_ = new_C3860_ & ~new_C3874_;
  assign new_C3920_ = new_C3860_ & ~new_C3874_;
  assign new_C3921_ = ~new_C3860_ & new_C3874_;
  assign new_C3922_ = new_E5437_;
  assign new_C3923_ = new_E5504_;
  assign new_C3924_ = new_E5571_;
  assign new_C3925_ = new_E5638_;
  assign new_C3926_ = new_E5705_;
  assign new_C3927_ = new_E5772_;
  assign new_C3928_ = new_C3935_ & new_C3934_;
  assign new_C3929_ = new_C3937_ | new_C3936_;
  assign new_C3930_ = new_C3939_ | new_C3938_;
  assign new_C3931_ = new_C3941_ & new_C3940_;
  assign new_C3932_ = new_C3941_ & new_C3942_;
  assign new_C3933_ = new_C3934_ | new_C3943_;
  assign new_C3934_ = new_C3923_ | new_C3946_;
  assign new_C3935_ = new_C3945_ | new_C3944_;
  assign new_C3936_ = new_C3950_ & new_C3949_;
  assign new_C3937_ = new_C3948_ & new_C3947_;
  assign new_C3938_ = new_C3953_ | new_C3952_;
  assign new_C3939_ = new_C3948_ & new_C3951_;
  assign new_C3940_ = new_C3923_ | new_C3956_;
  assign new_C3941_ = new_C3955_ | new_C3954_;
  assign new_C3942_ = new_C3958_ | new_C3957_;
  assign new_C3943_ = ~new_C3934_ & new_C3960_;
  assign new_C3944_ = ~new_C3936_ & new_C3948_;
  assign new_C3945_ = new_C3936_ & ~new_C3948_;
  assign new_C3946_ = new_C3922_ & ~new_C3923_;
  assign new_C3947_ = ~new_C3969_ | ~new_C3970_;
  assign new_C3948_ = new_C3962_ | new_C3964_;
  assign new_C3949_ = new_C3972_ | new_C3971_;
  assign new_C3950_ = new_C3966_ | new_C3965_;
  assign new_C3951_ = ~new_C3974_ | ~new_C3973_;
  assign new_C3952_ = ~new_C3975_ & new_C3976_;
  assign new_C3953_ = new_C3975_ & ~new_C3976_;
  assign new_C3954_ = ~new_C3922_ & new_C3923_;
  assign new_C3955_ = new_C3922_ & ~new_C3923_;
  assign new_C3956_ = ~new_C3938_ | new_C3948_;
  assign new_C3957_ = new_C3938_ & new_C3948_;
  assign new_C3958_ = ~new_C3938_ & ~new_C3948_;
  assign new_C3959_ = new_C3980_ | new_C3979_;
  assign new_C3960_ = new_C3926_ | new_C3959_;
  assign new_C3961_ = new_C3984_ | new_C3983_;
  assign new_C3962_ = ~new_C3926_ & new_C3961_;
  assign new_C3963_ = new_C3982_ | new_C3981_;
  assign new_C3964_ = new_C3926_ & new_C3963_;
  assign new_C3965_ = new_C3924_ & ~new_C3934_;
  assign new_C3966_ = ~new_C3924_ & new_C3934_;
  assign new_C3967_ = ~new_C3923_ | ~new_C3948_;
  assign new_C3968_ = new_C3934_ & new_C3967_;
  assign new_C3969_ = ~new_C3934_ & ~new_C3968_;
  assign new_C3970_ = new_C3934_ | new_C3967_;
  assign new_C3971_ = ~new_C3924_ & new_C3925_;
  assign new_C3972_ = new_C3924_ & ~new_C3925_;
  assign new_C3973_ = new_C3941_ | new_C3978_;
  assign new_C3974_ = ~new_C3941_ & ~new_C3977_;
  assign new_C3975_ = new_C3924_ | new_C3941_;
  assign new_C3976_ = new_C3924_ | new_C3925_;
  assign new_C3977_ = new_C3941_ & new_C3978_;
  assign new_C3978_ = ~new_C3923_ | ~new_C3948_;
  assign new_C3979_ = new_C3956_ & new_C3976_;
  assign new_C3980_ = ~new_C3956_ & ~new_C3976_;
  assign new_C3981_ = new_C3985_ | new_C3986_;
  assign new_C3982_ = ~new_C3927_ & new_C3941_;
  assign new_C3983_ = new_C3987_ | new_C3988_;
  assign new_C3984_ = new_C3927_ & new_C3941_;
  assign new_C3985_ = ~new_C3927_ & ~new_C3941_;
  assign new_C3986_ = new_C3927_ & ~new_C3941_;
  assign new_C3987_ = new_C3927_ & ~new_C3941_;
  assign new_C3988_ = ~new_C3927_ & new_C3941_;
  assign new_C3989_ = new_E5839_;
  assign new_C3990_ = new_E5906_;
  assign new_C3991_ = new_E5973_;
  assign new_C3992_ = new_E6040_;
  assign new_C3993_ = new_E6107_;
  assign new_C3994_ = new_E6174_;
  assign new_C3995_ = new_C4002_ & new_C4001_;
  assign new_C3996_ = new_C4004_ | new_C4003_;
  assign new_C3997_ = new_C4006_ | new_C4005_;
  assign new_C3998_ = new_C4008_ & new_C4007_;
  assign new_C3999_ = new_C4008_ & new_C4009_;
  assign new_C4000_ = new_C4001_ | new_C4010_;
  assign new_C4001_ = new_C3990_ | new_C4013_;
  assign new_C4002_ = new_C4012_ | new_C4011_;
  assign new_C4003_ = new_C4017_ & new_C4016_;
  assign new_C4004_ = new_C4015_ & new_C4014_;
  assign new_C4005_ = new_C4020_ | new_C4019_;
  assign new_C4006_ = new_C4015_ & new_C4018_;
  assign new_C4007_ = new_C3990_ | new_C4023_;
  assign new_C4008_ = new_C4022_ | new_C4021_;
  assign new_C4009_ = new_C4025_ | new_C4024_;
  assign new_C4010_ = ~new_C4001_ & new_C4027_;
  assign new_C4011_ = ~new_C4003_ & new_C4015_;
  assign new_C4012_ = new_C4003_ & ~new_C4015_;
  assign new_C4013_ = new_C3989_ & ~new_C3990_;
  assign new_C4014_ = ~new_C4036_ | ~new_C4037_;
  assign new_C4015_ = new_C4029_ | new_C4031_;
  assign new_C4016_ = new_C4039_ | new_C4038_;
  assign new_C4017_ = new_C4033_ | new_C4032_;
  assign new_C4018_ = ~new_C4041_ | ~new_C4040_;
  assign new_C4019_ = ~new_C4042_ & new_C4043_;
  assign new_C4020_ = new_C4042_ & ~new_C4043_;
  assign new_C4021_ = ~new_C3989_ & new_C3990_;
  assign new_C4022_ = new_C3989_ & ~new_C3990_;
  assign new_C4023_ = ~new_C4005_ | new_C4015_;
  assign new_C4024_ = new_C4005_ & new_C4015_;
  assign new_C4025_ = ~new_C4005_ & ~new_C4015_;
  assign new_C4026_ = new_C4047_ | new_C4046_;
  assign new_C4027_ = new_C3993_ | new_C4026_;
  assign new_C4028_ = new_C4051_ | new_C4050_;
  assign new_C4029_ = ~new_C3993_ & new_C4028_;
  assign new_C4030_ = new_C4049_ | new_C4048_;
  assign new_C4031_ = new_C3993_ & new_C4030_;
  assign new_C4032_ = new_C3991_ & ~new_C4001_;
  assign new_C4033_ = ~new_C3991_ & new_C4001_;
  assign new_C4034_ = ~new_C3990_ | ~new_C4015_;
  assign new_C4035_ = new_C4001_ & new_C4034_;
  assign new_C4036_ = ~new_C4001_ & ~new_C4035_;
  assign new_C4037_ = new_C4001_ | new_C4034_;
  assign new_C4038_ = ~new_C3991_ & new_C3992_;
  assign new_C4039_ = new_C3991_ & ~new_C3992_;
  assign new_C4040_ = new_C4008_ | new_C4045_;
  assign new_C4041_ = ~new_C4008_ & ~new_C4044_;
  assign new_C4042_ = new_C3991_ | new_C4008_;
  assign new_C4043_ = new_C3991_ | new_C3992_;
  assign new_C4044_ = new_C4008_ & new_C4045_;
  assign new_C4045_ = ~new_C3990_ | ~new_C4015_;
  assign new_C4046_ = new_C4023_ & new_C4043_;
  assign new_C4047_ = ~new_C4023_ & ~new_C4043_;
  assign new_C4048_ = new_C4052_ | new_C4053_;
  assign new_C4049_ = ~new_C3994_ & new_C4008_;
  assign new_C4050_ = new_C4054_ | new_C4055_;
  assign new_C4051_ = new_C3994_ & new_C4008_;
  assign new_C4052_ = ~new_C3994_ & ~new_C4008_;
  assign new_C4053_ = new_C3994_ & ~new_C4008_;
  assign new_C4054_ = new_C3994_ & ~new_C4008_;
  assign new_C4055_ = ~new_C3994_ & new_C4008_;
  assign new_C4056_ = new_E6241_;
  assign new_C4057_ = new_E6308_;
  assign new_C4058_ = new_E6375_;
  assign new_C4059_ = new_E6442_;
  assign new_C4060_ = new_E6509_;
  assign new_C4061_ = new_E6576_;
  assign new_C4062_ = new_C4069_ & new_C4068_;
  assign new_C4063_ = new_C4071_ | new_C4070_;
  assign new_C4064_ = new_C4073_ | new_C4072_;
  assign new_C4065_ = new_C4075_ & new_C4074_;
  assign new_C4066_ = new_C4075_ & new_C4076_;
  assign new_C4067_ = new_C4068_ | new_C4077_;
  assign new_C4068_ = new_C4057_ | new_C4080_;
  assign new_C4069_ = new_C4079_ | new_C4078_;
  assign new_C4070_ = new_C4084_ & new_C4083_;
  assign new_C4071_ = new_C4082_ & new_C4081_;
  assign new_C4072_ = new_C4087_ | new_C4086_;
  assign new_C4073_ = new_C4082_ & new_C4085_;
  assign new_C4074_ = new_C4057_ | new_C4090_;
  assign new_C4075_ = new_C4089_ | new_C4088_;
  assign new_C4076_ = new_C4092_ | new_C4091_;
  assign new_C4077_ = ~new_C4068_ & new_C4094_;
  assign new_C4078_ = ~new_C4070_ & new_C4082_;
  assign new_C4079_ = new_C4070_ & ~new_C4082_;
  assign new_C4080_ = new_C4056_ & ~new_C4057_;
  assign new_C4081_ = ~new_C4103_ | ~new_C4104_;
  assign new_C4082_ = new_C4096_ | new_C4098_;
  assign new_C4083_ = new_C4106_ | new_C4105_;
  assign new_C4084_ = new_C4100_ | new_C4099_;
  assign new_C4085_ = ~new_C4108_ | ~new_C4107_;
  assign new_C4086_ = ~new_C4109_ & new_C4110_;
  assign new_C4087_ = new_C4109_ & ~new_C4110_;
  assign new_C4088_ = ~new_C4056_ & new_C4057_;
  assign new_C4089_ = new_C4056_ & ~new_C4057_;
  assign new_C4090_ = ~new_C4072_ | new_C4082_;
  assign new_C4091_ = new_C4072_ & new_C4082_;
  assign new_C4092_ = ~new_C4072_ & ~new_C4082_;
  assign new_C4093_ = new_C4114_ | new_C4113_;
  assign new_C4094_ = new_C4060_ | new_C4093_;
  assign new_C4095_ = new_C4118_ | new_C4117_;
  assign new_C4096_ = ~new_C4060_ & new_C4095_;
  assign new_C4097_ = new_C4116_ | new_C4115_;
  assign new_C4098_ = new_C4060_ & new_C4097_;
  assign new_C4099_ = new_C4058_ & ~new_C4068_;
  assign new_C4100_ = ~new_C4058_ & new_C4068_;
  assign new_C4101_ = ~new_C4057_ | ~new_C4082_;
  assign new_C4102_ = new_C4068_ & new_C4101_;
  assign new_C4103_ = ~new_C4068_ & ~new_C4102_;
  assign new_C4104_ = new_C4068_ | new_C4101_;
  assign new_C4105_ = ~new_C4058_ & new_C4059_;
  assign new_C4106_ = new_C4058_ & ~new_C4059_;
  assign new_C4107_ = new_C4075_ | new_C4112_;
  assign new_C4108_ = ~new_C4075_ & ~new_C4111_;
  assign new_C4109_ = new_C4058_ | new_C4075_;
  assign new_C4110_ = new_C4058_ | new_C4059_;
  assign new_C4111_ = new_C4075_ & new_C4112_;
  assign new_C4112_ = ~new_C4057_ | ~new_C4082_;
  assign new_C4113_ = new_C4090_ & new_C4110_;
  assign new_C4114_ = ~new_C4090_ & ~new_C4110_;
  assign new_C4115_ = new_C4119_ | new_C4120_;
  assign new_C4116_ = ~new_C4061_ & new_C4075_;
  assign new_C4117_ = new_C4121_ | new_C4122_;
  assign new_C4118_ = new_C4061_ & new_C4075_;
  assign new_C4119_ = ~new_C4061_ & ~new_C4075_;
  assign new_C4120_ = new_C4061_ & ~new_C4075_;
  assign new_C4121_ = new_C4061_ & ~new_C4075_;
  assign new_C4122_ = ~new_C4061_ & new_C4075_;
  assign new_C4123_ = new_E6643_;
  assign new_C4124_ = new_E6710_;
  assign new_C4125_ = new_E6777_;
  assign new_C4126_ = new_E6844_;
  assign new_C4127_ = new_E6911_;
  assign new_C4128_ = new_E6978_;
  assign new_C4129_ = new_C4136_ & new_C4135_;
  assign new_C4130_ = new_C4138_ | new_C4137_;
  assign new_C4131_ = new_C4140_ | new_C4139_;
  assign new_C4132_ = new_C4142_ & new_C4141_;
  assign new_C4133_ = new_C4142_ & new_C4143_;
  assign new_C4134_ = new_C4135_ | new_C4144_;
  assign new_C4135_ = new_C4124_ | new_C4147_;
  assign new_C4136_ = new_C4146_ | new_C4145_;
  assign new_C4137_ = new_C4151_ & new_C4150_;
  assign new_C4138_ = new_C4149_ & new_C4148_;
  assign new_C4139_ = new_C4154_ | new_C4153_;
  assign new_C4140_ = new_C4149_ & new_C4152_;
  assign new_C4141_ = new_C4124_ | new_C4157_;
  assign new_C4142_ = new_C4156_ | new_C4155_;
  assign new_C4143_ = new_C4159_ | new_C4158_;
  assign new_C4144_ = ~new_C4135_ & new_C4161_;
  assign new_C4145_ = ~new_C4137_ & new_C4149_;
  assign new_C4146_ = new_C4137_ & ~new_C4149_;
  assign new_C4147_ = new_C4123_ & ~new_C4124_;
  assign new_C4148_ = ~new_C4170_ | ~new_C4171_;
  assign new_C4149_ = new_C4163_ | new_C4165_;
  assign new_C4150_ = new_C4173_ | new_C4172_;
  assign new_C4151_ = new_C4167_ | new_C4166_;
  assign new_C4152_ = ~new_C4175_ | ~new_C4174_;
  assign new_C4153_ = ~new_C4176_ & new_C4177_;
  assign new_C4154_ = new_C4176_ & ~new_C4177_;
  assign new_C4155_ = ~new_C4123_ & new_C4124_;
  assign new_C4156_ = new_C4123_ & ~new_C4124_;
  assign new_C4157_ = ~new_C4139_ | new_C4149_;
  assign new_C4158_ = new_C4139_ & new_C4149_;
  assign new_C4159_ = ~new_C4139_ & ~new_C4149_;
  assign new_C4160_ = new_C4181_ | new_C4180_;
  assign new_C4161_ = new_C4127_ | new_C4160_;
  assign new_C4162_ = new_C4185_ | new_C4184_;
  assign new_C4163_ = ~new_C4127_ & new_C4162_;
  assign new_C4164_ = new_C4183_ | new_C4182_;
  assign new_C4165_ = new_C4127_ & new_C4164_;
  assign new_C4166_ = new_C4125_ & ~new_C4135_;
  assign new_C4167_ = ~new_C4125_ & new_C4135_;
  assign new_C4168_ = ~new_C4124_ | ~new_C4149_;
  assign new_C4169_ = new_C4135_ & new_C4168_;
  assign new_C4170_ = ~new_C4135_ & ~new_C4169_;
  assign new_C4171_ = new_C4135_ | new_C4168_;
  assign new_C4172_ = ~new_C4125_ & new_C4126_;
  assign new_C4173_ = new_C4125_ & ~new_C4126_;
  assign new_C4174_ = new_C4142_ | new_C4179_;
  assign new_C4175_ = ~new_C4142_ & ~new_C4178_;
  assign new_C4176_ = new_C4125_ | new_C4142_;
  assign new_C4177_ = new_C4125_ | new_C4126_;
  assign new_C4178_ = new_C4142_ & new_C4179_;
  assign new_C4179_ = ~new_C4124_ | ~new_C4149_;
  assign new_C4180_ = new_C4157_ & new_C4177_;
  assign new_C4181_ = ~new_C4157_ & ~new_C4177_;
  assign new_C4182_ = new_C4186_ | new_C4187_;
  assign new_C4183_ = ~new_C4128_ & new_C4142_;
  assign new_C4184_ = new_C4188_ | new_C4189_;
  assign new_C4185_ = new_C4128_ & new_C4142_;
  assign new_C4186_ = ~new_C4128_ & ~new_C4142_;
  assign new_C4187_ = new_C4128_ & ~new_C4142_;
  assign new_C4188_ = new_C4128_ & ~new_C4142_;
  assign new_C4189_ = ~new_C4128_ & new_C4142_;
  assign new_C4190_ = new_E7045_;
  assign new_C4191_ = new_E7112_;
  assign new_C4192_ = new_E7179_;
  assign new_C4193_ = new_E7246_;
  assign new_C4194_ = new_E7313_;
  assign new_C4195_ = new_E7380_;
  assign new_C4196_ = new_C4203_ & new_C4202_;
  assign new_C4197_ = new_C4205_ | new_C4204_;
  assign new_C4198_ = new_C4207_ | new_C4206_;
  assign new_C4199_ = new_C4209_ & new_C4208_;
  assign new_C4200_ = new_C4209_ & new_C4210_;
  assign new_C4201_ = new_C4202_ | new_C4211_;
  assign new_C4202_ = new_C4191_ | new_C4214_;
  assign new_C4203_ = new_C4213_ | new_C4212_;
  assign new_C4204_ = new_C4218_ & new_C4217_;
  assign new_C4205_ = new_C4216_ & new_C4215_;
  assign new_C4206_ = new_C4221_ | new_C4220_;
  assign new_C4207_ = new_C4216_ & new_C4219_;
  assign new_C4208_ = new_C4191_ | new_C4224_;
  assign new_C4209_ = new_C4223_ | new_C4222_;
  assign new_C4210_ = new_C4226_ | new_C4225_;
  assign new_C4211_ = ~new_C4202_ & new_C4228_;
  assign new_C4212_ = ~new_C4204_ & new_C4216_;
  assign new_C4213_ = new_C4204_ & ~new_C4216_;
  assign new_C4214_ = new_C4190_ & ~new_C4191_;
  assign new_C4215_ = ~new_C4237_ | ~new_C4238_;
  assign new_C4216_ = new_C4230_ | new_C4232_;
  assign new_C4217_ = new_C4240_ | new_C4239_;
  assign new_C4218_ = new_C4234_ | new_C4233_;
  assign new_C4219_ = ~new_C4242_ | ~new_C4241_;
  assign new_C4220_ = ~new_C4243_ & new_C4244_;
  assign new_C4221_ = new_C4243_ & ~new_C4244_;
  assign new_C4222_ = ~new_C4190_ & new_C4191_;
  assign new_C4223_ = new_C4190_ & ~new_C4191_;
  assign new_C4224_ = ~new_C4206_ | new_C4216_;
  assign new_C4225_ = new_C4206_ & new_C4216_;
  assign new_C4226_ = ~new_C4206_ & ~new_C4216_;
  assign new_C4227_ = new_C4248_ | new_C4247_;
  assign new_C4228_ = new_C4194_ | new_C4227_;
  assign new_C4229_ = new_C4252_ | new_C4251_;
  assign new_C4230_ = ~new_C4194_ & new_C4229_;
  assign new_C4231_ = new_C4250_ | new_C4249_;
  assign new_C4232_ = new_C4194_ & new_C4231_;
  assign new_C4233_ = new_C4192_ & ~new_C4202_;
  assign new_C4234_ = ~new_C4192_ & new_C4202_;
  assign new_C4235_ = ~new_C4191_ | ~new_C4216_;
  assign new_C4236_ = new_C4202_ & new_C4235_;
  assign new_C4237_ = ~new_C4202_ & ~new_C4236_;
  assign new_C4238_ = new_C4202_ | new_C4235_;
  assign new_C4239_ = ~new_C4192_ & new_C4193_;
  assign new_C4240_ = new_C4192_ & ~new_C4193_;
  assign new_C4241_ = new_C4209_ | new_C4246_;
  assign new_C4242_ = ~new_C4209_ & ~new_C4245_;
  assign new_C4243_ = new_C4192_ | new_C4209_;
  assign new_C4244_ = new_C4192_ | new_C4193_;
  assign new_C4245_ = new_C4209_ & new_C4246_;
  assign new_C4246_ = ~new_C4191_ | ~new_C4216_;
  assign new_C4247_ = new_C4224_ & new_C4244_;
  assign new_C4248_ = ~new_C4224_ & ~new_C4244_;
  assign new_C4249_ = new_C4253_ | new_C4254_;
  assign new_C4250_ = ~new_C4195_ & new_C4209_;
  assign new_C4251_ = new_C4255_ | new_C4256_;
  assign new_C4252_ = new_C4195_ & new_C4209_;
  assign new_C4253_ = ~new_C4195_ & ~new_C4209_;
  assign new_C4254_ = new_C4195_ & ~new_C4209_;
  assign new_C4255_ = new_C4195_ & ~new_C4209_;
  assign new_C4256_ = ~new_C4195_ & new_C4209_;
  assign new_C4257_ = new_E7447_;
  assign new_C4258_ = new_E7514_;
  assign new_C4259_ = new_E7581_;
  assign new_C4260_ = new_E7648_;
  assign new_C4261_ = new_E7715_;
  assign new_C4262_ = new_E7782_;
  assign new_C4263_ = new_C4270_ & new_C4269_;
  assign new_C4264_ = new_C4272_ | new_C4271_;
  assign new_C4265_ = new_C4274_ | new_C4273_;
  assign new_C4266_ = new_C4276_ & new_C4275_;
  assign new_C4267_ = new_C4276_ & new_C4277_;
  assign new_C4268_ = new_C4269_ | new_C4278_;
  assign new_C4269_ = new_C4258_ | new_C4281_;
  assign new_C4270_ = new_C4280_ | new_C4279_;
  assign new_C4271_ = new_C4285_ & new_C4284_;
  assign new_C4272_ = new_C4283_ & new_C4282_;
  assign new_C4273_ = new_C4288_ | new_C4287_;
  assign new_C4274_ = new_C4283_ & new_C4286_;
  assign new_C4275_ = new_C4258_ | new_C4291_;
  assign new_C4276_ = new_C4290_ | new_C4289_;
  assign new_C4277_ = new_C4293_ | new_C4292_;
  assign new_C4278_ = ~new_C4269_ & new_C4295_;
  assign new_C4279_ = ~new_C4271_ & new_C4283_;
  assign new_C4280_ = new_C4271_ & ~new_C4283_;
  assign new_C4281_ = new_C4257_ & ~new_C4258_;
  assign new_C4282_ = ~new_C4304_ | ~new_C4305_;
  assign new_C4283_ = new_C4297_ | new_C4299_;
  assign new_C4284_ = new_C4307_ | new_C4306_;
  assign new_C4285_ = new_C4301_ | new_C4300_;
  assign new_C4286_ = ~new_C4309_ | ~new_C4308_;
  assign new_C4287_ = ~new_C4310_ & new_C4311_;
  assign new_C4288_ = new_C4310_ & ~new_C4311_;
  assign new_C4289_ = ~new_C4257_ & new_C4258_;
  assign new_C4290_ = new_C4257_ & ~new_C4258_;
  assign new_C4291_ = ~new_C4273_ | new_C4283_;
  assign new_C4292_ = new_C4273_ & new_C4283_;
  assign new_C4293_ = ~new_C4273_ & ~new_C4283_;
  assign new_C4294_ = new_C4315_ | new_C4314_;
  assign new_C4295_ = new_C4261_ | new_C4294_;
  assign new_C4296_ = new_C4319_ | new_C4318_;
  assign new_C4297_ = ~new_C4261_ & new_C4296_;
  assign new_C4298_ = new_C4317_ | new_C4316_;
  assign new_C4299_ = new_C4261_ & new_C4298_;
  assign new_C4300_ = new_C4259_ & ~new_C4269_;
  assign new_C4301_ = ~new_C4259_ & new_C4269_;
  assign new_C4302_ = ~new_C4258_ | ~new_C4283_;
  assign new_C4303_ = new_C4269_ & new_C4302_;
  assign new_C4304_ = ~new_C4269_ & ~new_C4303_;
  assign new_C4305_ = new_C4269_ | new_C4302_;
  assign new_C4306_ = ~new_C4259_ & new_C4260_;
  assign new_C4307_ = new_C4259_ & ~new_C4260_;
  assign new_C4308_ = new_C4276_ | new_C4313_;
  assign new_C4309_ = ~new_C4276_ & ~new_C4312_;
  assign new_C4310_ = new_C4259_ | new_C4276_;
  assign new_C4311_ = new_C4259_ | new_C4260_;
  assign new_C4312_ = new_C4276_ & new_C4313_;
  assign new_C4313_ = ~new_C4258_ | ~new_C4283_;
  assign new_C4314_ = new_C4291_ & new_C4311_;
  assign new_C4315_ = ~new_C4291_ & ~new_C4311_;
  assign new_C4316_ = new_C4320_ | new_C4321_;
  assign new_C4317_ = ~new_C4262_ & new_C4276_;
  assign new_C4318_ = new_C4322_ | new_C4323_;
  assign new_C4319_ = new_C4262_ & new_C4276_;
  assign new_C4320_ = ~new_C4262_ & ~new_C4276_;
  assign new_C4321_ = new_C4262_ & ~new_C4276_;
  assign new_C4322_ = new_C4262_ & ~new_C4276_;
  assign new_C4323_ = ~new_C4262_ & new_C4276_;
  assign new_C4324_ = new_E7849_;
  assign new_C4325_ = new_E7916_;
  assign new_C4326_ = new_E7983_;
  assign new_C4327_ = new_E8050_;
  assign new_C4328_ = new_E8117_;
  assign new_C4329_ = new_E8184_;
  assign new_C4330_ = new_C4337_ & new_C4336_;
  assign new_C4331_ = new_C4339_ | new_C4338_;
  assign new_C4332_ = new_C4341_ | new_C4340_;
  assign new_C4333_ = new_C4343_ & new_C4342_;
  assign new_C4334_ = new_C4343_ & new_C4344_;
  assign new_C4335_ = new_C4336_ | new_C4345_;
  assign new_C4336_ = new_C4325_ | new_C4348_;
  assign new_C4337_ = new_C4347_ | new_C4346_;
  assign new_C4338_ = new_C4352_ & new_C4351_;
  assign new_C4339_ = new_C4350_ & new_C4349_;
  assign new_C4340_ = new_C4355_ | new_C4354_;
  assign new_C4341_ = new_C4350_ & new_C4353_;
  assign new_C4342_ = new_C4325_ | new_C4358_;
  assign new_C4343_ = new_C4357_ | new_C4356_;
  assign new_C4344_ = new_C4360_ | new_C4359_;
  assign new_C4345_ = ~new_C4336_ & new_C4362_;
  assign new_C4346_ = ~new_C4338_ & new_C4350_;
  assign new_C4347_ = new_C4338_ & ~new_C4350_;
  assign new_C4348_ = new_C4324_ & ~new_C4325_;
  assign new_C4349_ = ~new_C4371_ | ~new_C4372_;
  assign new_C4350_ = new_C4364_ | new_C4366_;
  assign new_C4351_ = new_C4374_ | new_C4373_;
  assign new_C4352_ = new_C4368_ | new_C4367_;
  assign new_C4353_ = ~new_C4376_ | ~new_C4375_;
  assign new_C4354_ = ~new_C4377_ & new_C4378_;
  assign new_C4355_ = new_C4377_ & ~new_C4378_;
  assign new_C4356_ = ~new_C4324_ & new_C4325_;
  assign new_C4357_ = new_C4324_ & ~new_C4325_;
  assign new_C4358_ = ~new_C4340_ | new_C4350_;
  assign new_C4359_ = new_C4340_ & new_C4350_;
  assign new_C4360_ = ~new_C4340_ & ~new_C4350_;
  assign new_C4361_ = new_C4382_ | new_C4381_;
  assign new_C4362_ = new_C4328_ | new_C4361_;
  assign new_C4363_ = new_C4386_ | new_C4385_;
  assign new_C4364_ = ~new_C4328_ & new_C4363_;
  assign new_C4365_ = new_C4384_ | new_C4383_;
  assign new_C4366_ = new_C4328_ & new_C4365_;
  assign new_C4367_ = new_C4326_ & ~new_C4336_;
  assign new_C4368_ = ~new_C4326_ & new_C4336_;
  assign new_C4369_ = ~new_C4325_ | ~new_C4350_;
  assign new_C4370_ = new_C4336_ & new_C4369_;
  assign new_C4371_ = ~new_C4336_ & ~new_C4370_;
  assign new_C4372_ = new_C4336_ | new_C4369_;
  assign new_C4373_ = ~new_C4326_ & new_C4327_;
  assign new_C4374_ = new_C4326_ & ~new_C4327_;
  assign new_C4375_ = new_C4343_ | new_C4380_;
  assign new_C4376_ = ~new_C4343_ & ~new_C4379_;
  assign new_C4377_ = new_C4326_ | new_C4343_;
  assign new_C4378_ = new_C4326_ | new_C4327_;
  assign new_C4379_ = new_C4343_ & new_C4380_;
  assign new_C4380_ = ~new_C4325_ | ~new_C4350_;
  assign new_C4381_ = new_C4358_ & new_C4378_;
  assign new_C4382_ = ~new_C4358_ & ~new_C4378_;
  assign new_C4383_ = new_C4387_ | new_C4388_;
  assign new_C4384_ = ~new_C4329_ & new_C4343_;
  assign new_C4385_ = new_C4389_ | new_C4390_;
  assign new_C4386_ = new_C4329_ & new_C4343_;
  assign new_C4387_ = ~new_C4329_ & ~new_C4343_;
  assign new_C4388_ = new_C4329_ & ~new_C4343_;
  assign new_C4389_ = new_C4329_ & ~new_C4343_;
  assign new_C4390_ = ~new_C4329_ & new_C4343_;
  assign new_C4391_ = new_E8251_;
  assign new_C4392_ = new_E8318_;
  assign new_C4393_ = new_E8385_;
  assign new_C4394_ = new_E8452_;
  assign new_C4395_ = new_E8519_;
  assign new_C4396_ = new_E8586_;
  assign new_C4397_ = new_C4404_ & new_C4403_;
  assign new_C4398_ = new_C4406_ | new_C4405_;
  assign new_C4399_ = new_C4408_ | new_C4407_;
  assign new_C4400_ = new_C4410_ & new_C4409_;
  assign new_C4401_ = new_C4410_ & new_C4411_;
  assign new_C4402_ = new_C4403_ | new_C4412_;
  assign new_C4403_ = new_C4392_ | new_C4415_;
  assign new_C4404_ = new_C4414_ | new_C4413_;
  assign new_C4405_ = new_C4419_ & new_C4418_;
  assign new_C4406_ = new_C4417_ & new_C4416_;
  assign new_C4407_ = new_C4422_ | new_C4421_;
  assign new_C4408_ = new_C4417_ & new_C4420_;
  assign new_C4409_ = new_C4392_ | new_C4425_;
  assign new_C4410_ = new_C4424_ | new_C4423_;
  assign new_C4411_ = new_C4427_ | new_C4426_;
  assign new_C4412_ = ~new_C4403_ & new_C4429_;
  assign new_C4413_ = ~new_C4405_ & new_C4417_;
  assign new_C4414_ = new_C4405_ & ~new_C4417_;
  assign new_C4415_ = new_C4391_ & ~new_C4392_;
  assign new_C4416_ = ~new_C4438_ | ~new_C4439_;
  assign new_C4417_ = new_C4431_ | new_C4433_;
  assign new_C4418_ = new_C4441_ | new_C4440_;
  assign new_C4419_ = new_C4435_ | new_C4434_;
  assign new_C4420_ = ~new_C4443_ | ~new_C4442_;
  assign new_C4421_ = ~new_C4444_ & new_C4445_;
  assign new_C4422_ = new_C4444_ & ~new_C4445_;
  assign new_C4423_ = ~new_C4391_ & new_C4392_;
  assign new_C4424_ = new_C4391_ & ~new_C4392_;
  assign new_C4425_ = ~new_C4407_ | new_C4417_;
  assign new_C4426_ = new_C4407_ & new_C4417_;
  assign new_C4427_ = ~new_C4407_ & ~new_C4417_;
  assign new_C4428_ = new_C4449_ | new_C4448_;
  assign new_C4429_ = new_C4395_ | new_C4428_;
  assign new_C4430_ = new_C4453_ | new_C4452_;
  assign new_C4431_ = ~new_C4395_ & new_C4430_;
  assign new_C4432_ = new_C4451_ | new_C4450_;
  assign new_C4433_ = new_C4395_ & new_C4432_;
  assign new_C4434_ = new_C4393_ & ~new_C4403_;
  assign new_C4435_ = ~new_C4393_ & new_C4403_;
  assign new_C4436_ = ~new_C4392_ | ~new_C4417_;
  assign new_C4437_ = new_C4403_ & new_C4436_;
  assign new_C4438_ = ~new_C4403_ & ~new_C4437_;
  assign new_C4439_ = new_C4403_ | new_C4436_;
  assign new_C4440_ = ~new_C4393_ & new_C4394_;
  assign new_C4441_ = new_C4393_ & ~new_C4394_;
  assign new_C4442_ = new_C4410_ | new_C4447_;
  assign new_C4443_ = ~new_C4410_ & ~new_C4446_;
  assign new_C4444_ = new_C4393_ | new_C4410_;
  assign new_C4445_ = new_C4393_ | new_C4394_;
  assign new_C4446_ = new_C4410_ & new_C4447_;
  assign new_C4447_ = ~new_C4392_ | ~new_C4417_;
  assign new_C4448_ = new_C4425_ & new_C4445_;
  assign new_C4449_ = ~new_C4425_ & ~new_C4445_;
  assign new_C4450_ = new_C4454_ | new_C4455_;
  assign new_C4451_ = ~new_C4396_ & new_C4410_;
  assign new_C4452_ = new_C4456_ | new_C4457_;
  assign new_C4453_ = new_C4396_ & new_C4410_;
  assign new_C4454_ = ~new_C4396_ & ~new_C4410_;
  assign new_C4455_ = new_C4396_ & ~new_C4410_;
  assign new_C4456_ = new_C4396_ & ~new_C4410_;
  assign new_C4457_ = ~new_C4396_ & new_C4410_;
  assign new_C4458_ = new_E8653_;
  assign new_C4459_ = new_E8720_;
  assign new_C4460_ = new_E8787_;
  assign new_C4461_ = new_E8854_;
  assign new_C4462_ = new_E8921_;
  assign new_C4463_ = new_E8988_;
  assign new_C4464_ = new_C4471_ & new_C4470_;
  assign new_C4465_ = new_C4473_ | new_C4472_;
  assign new_C4466_ = new_C4475_ | new_C4474_;
  assign new_C4467_ = new_C4477_ & new_C4476_;
  assign new_C4468_ = new_C4477_ & new_C4478_;
  assign new_C4469_ = new_C4470_ | new_C4479_;
  assign new_C4470_ = new_C4459_ | new_C4482_;
  assign new_C4471_ = new_C4481_ | new_C4480_;
  assign new_C4472_ = new_C4486_ & new_C4485_;
  assign new_C4473_ = new_C4484_ & new_C4483_;
  assign new_C4474_ = new_C4489_ | new_C4488_;
  assign new_C4475_ = new_C4484_ & new_C4487_;
  assign new_C4476_ = new_C4459_ | new_C4492_;
  assign new_C4477_ = new_C4491_ | new_C4490_;
  assign new_C4478_ = new_C4494_ | new_C4493_;
  assign new_C4479_ = ~new_C4470_ & new_C4496_;
  assign new_C4480_ = ~new_C4472_ & new_C4484_;
  assign new_C4481_ = new_C4472_ & ~new_C4484_;
  assign new_C4482_ = new_C4458_ & ~new_C4459_;
  assign new_C4483_ = ~new_C4505_ | ~new_C4506_;
  assign new_C4484_ = new_C4498_ | new_C4500_;
  assign new_C4485_ = new_C4508_ | new_C4507_;
  assign new_C4486_ = new_C4502_ | new_C4501_;
  assign new_C4487_ = ~new_C4510_ | ~new_C4509_;
  assign new_C4488_ = ~new_C4511_ & new_C4512_;
  assign new_C4489_ = new_C4511_ & ~new_C4512_;
  assign new_C4490_ = ~new_C4458_ & new_C4459_;
  assign new_C4491_ = new_C4458_ & ~new_C4459_;
  assign new_C4492_ = ~new_C4474_ | new_C4484_;
  assign new_C4493_ = new_C4474_ & new_C4484_;
  assign new_C4494_ = ~new_C4474_ & ~new_C4484_;
  assign new_C4495_ = new_C4516_ | new_C4515_;
  assign new_C4496_ = new_C4462_ | new_C4495_;
  assign new_C4497_ = new_C4520_ | new_C4519_;
  assign new_C4498_ = ~new_C4462_ & new_C4497_;
  assign new_C4499_ = new_C4518_ | new_C4517_;
  assign new_C4500_ = new_C4462_ & new_C4499_;
  assign new_C4501_ = new_C4460_ & ~new_C4470_;
  assign new_C4502_ = ~new_C4460_ & new_C4470_;
  assign new_C4503_ = ~new_C4459_ | ~new_C4484_;
  assign new_C4504_ = new_C4470_ & new_C4503_;
  assign new_C4505_ = ~new_C4470_ & ~new_C4504_;
  assign new_C4506_ = new_C4470_ | new_C4503_;
  assign new_C4507_ = ~new_C4460_ & new_C4461_;
  assign new_C4508_ = new_C4460_ & ~new_C4461_;
  assign new_C4509_ = new_C4477_ | new_C4514_;
  assign new_C4510_ = ~new_C4477_ & ~new_C4513_;
  assign new_C4511_ = new_C4460_ | new_C4477_;
  assign new_C4512_ = new_C4460_ | new_C4461_;
  assign new_C4513_ = new_C4477_ & new_C4514_;
  assign new_C4514_ = ~new_C4459_ | ~new_C4484_;
  assign new_C4515_ = new_C4492_ & new_C4512_;
  assign new_C4516_ = ~new_C4492_ & ~new_C4512_;
  assign new_C4517_ = new_C4521_ | new_C4522_;
  assign new_C4518_ = ~new_C4463_ & new_C4477_;
  assign new_C4519_ = new_C4523_ | new_C4524_;
  assign new_C4520_ = new_C4463_ & new_C4477_;
  assign new_C4521_ = ~new_C4463_ & ~new_C4477_;
  assign new_C4522_ = new_C4463_ & ~new_C4477_;
  assign new_C4523_ = new_C4463_ & ~new_C4477_;
  assign new_C4524_ = ~new_C4463_ & new_C4477_;
  assign new_C4525_ = new_E9055_;
  assign new_C4526_ = new_E9122_;
  assign new_C4527_ = new_E9189_;
  assign new_C4528_ = new_E9256_;
  assign new_C4529_ = new_E9323_;
  assign new_C4530_ = new_E9390_;
  assign new_C4531_ = new_C4538_ & new_C4537_;
  assign new_C4532_ = new_C4540_ | new_C4539_;
  assign new_C4533_ = new_C4542_ | new_C4541_;
  assign new_C4534_ = new_C4544_ & new_C4543_;
  assign new_C4535_ = new_C4544_ & new_C4545_;
  assign new_C4536_ = new_C4537_ | new_C4546_;
  assign new_C4537_ = new_C4526_ | new_C4549_;
  assign new_C4538_ = new_C4548_ | new_C4547_;
  assign new_C4539_ = new_C4553_ & new_C4552_;
  assign new_C4540_ = new_C4551_ & new_C4550_;
  assign new_C4541_ = new_C4556_ | new_C4555_;
  assign new_C4542_ = new_C4551_ & new_C4554_;
  assign new_C4543_ = new_C4526_ | new_C4559_;
  assign new_C4544_ = new_C4558_ | new_C4557_;
  assign new_C4545_ = new_C4561_ | new_C4560_;
  assign new_C4546_ = ~new_C4537_ & new_C4563_;
  assign new_C4547_ = ~new_C4539_ & new_C4551_;
  assign new_C4548_ = new_C4539_ & ~new_C4551_;
  assign new_C4549_ = new_C4525_ & ~new_C4526_;
  assign new_C4550_ = ~new_C4572_ | ~new_C4573_;
  assign new_C4551_ = new_C4565_ | new_C4567_;
  assign new_C4552_ = new_C4575_ | new_C4574_;
  assign new_C4553_ = new_C4569_ | new_C4568_;
  assign new_C4554_ = ~new_C4577_ | ~new_C4576_;
  assign new_C4555_ = ~new_C4578_ & new_C4579_;
  assign new_C4556_ = new_C4578_ & ~new_C4579_;
  assign new_C4557_ = ~new_C4525_ & new_C4526_;
  assign new_C4558_ = new_C4525_ & ~new_C4526_;
  assign new_C4559_ = ~new_C4541_ | new_C4551_;
  assign new_C4560_ = new_C4541_ & new_C4551_;
  assign new_C4561_ = ~new_C4541_ & ~new_C4551_;
  assign new_C4562_ = new_C4583_ | new_C4582_;
  assign new_C4563_ = new_C4529_ | new_C4562_;
  assign new_C4564_ = new_C4587_ | new_C4586_;
  assign new_C4565_ = ~new_C4529_ & new_C4564_;
  assign new_C4566_ = new_C4585_ | new_C4584_;
  assign new_C4567_ = new_C4529_ & new_C4566_;
  assign new_C4568_ = new_C4527_ & ~new_C4537_;
  assign new_C4569_ = ~new_C4527_ & new_C4537_;
  assign new_C4570_ = ~new_C4526_ | ~new_C4551_;
  assign new_C4571_ = new_C4537_ & new_C4570_;
  assign new_C4572_ = ~new_C4537_ & ~new_C4571_;
  assign new_C4573_ = new_C4537_ | new_C4570_;
  assign new_C4574_ = ~new_C4527_ & new_C4528_;
  assign new_C4575_ = new_C4527_ & ~new_C4528_;
  assign new_C4576_ = new_C4544_ | new_C4581_;
  assign new_C4577_ = ~new_C4544_ & ~new_C4580_;
  assign new_C4578_ = new_C4527_ | new_C4544_;
  assign new_C4579_ = new_C4527_ | new_C4528_;
  assign new_C4580_ = new_C4544_ & new_C4581_;
  assign new_C4581_ = ~new_C4526_ | ~new_C4551_;
  assign new_C4582_ = new_C4559_ & new_C4579_;
  assign new_C4583_ = ~new_C4559_ & ~new_C4579_;
  assign new_C4584_ = new_C4588_ | new_C4589_;
  assign new_C4585_ = ~new_C4530_ & new_C4544_;
  assign new_C4586_ = new_C4590_ | new_C4591_;
  assign new_C4587_ = new_C4530_ & new_C4544_;
  assign new_C4588_ = ~new_C4530_ & ~new_C4544_;
  assign new_C4589_ = new_C4530_ & ~new_C4544_;
  assign new_C4590_ = new_C4530_ & ~new_C4544_;
  assign new_C4591_ = ~new_C4530_ & new_C4544_;
  assign new_C4592_ = new_E9457_;
  assign new_C4593_ = new_E9524_;
  assign new_C4594_ = new_E9591_;
  assign new_C4595_ = new_E9658_;
  assign new_C4596_ = new_E9725_;
  assign new_C4597_ = new_E9792_;
  assign new_C4598_ = new_C4605_ & new_C4604_;
  assign new_C4599_ = new_C4607_ | new_C4606_;
  assign new_C4600_ = new_C4609_ | new_C4608_;
  assign new_C4601_ = new_C4611_ & new_C4610_;
  assign new_C4602_ = new_C4611_ & new_C4612_;
  assign new_C4603_ = new_C4604_ | new_C4613_;
  assign new_C4604_ = new_C4593_ | new_C4616_;
  assign new_C4605_ = new_C4615_ | new_C4614_;
  assign new_C4606_ = new_C4620_ & new_C4619_;
  assign new_C4607_ = new_C4618_ & new_C4617_;
  assign new_C4608_ = new_C4623_ | new_C4622_;
  assign new_C4609_ = new_C4618_ & new_C4621_;
  assign new_C4610_ = new_C4593_ | new_C4626_;
  assign new_C4611_ = new_C4625_ | new_C4624_;
  assign new_C4612_ = new_C4628_ | new_C4627_;
  assign new_C4613_ = ~new_C4604_ & new_C4630_;
  assign new_C4614_ = ~new_C4606_ & new_C4618_;
  assign new_C4615_ = new_C4606_ & ~new_C4618_;
  assign new_C4616_ = new_C4592_ & ~new_C4593_;
  assign new_C4617_ = ~new_C4639_ | ~new_C4640_;
  assign new_C4618_ = new_C4632_ | new_C4634_;
  assign new_C4619_ = new_C4642_ | new_C4641_;
  assign new_C4620_ = new_C4636_ | new_C4635_;
  assign new_C4621_ = ~new_C4644_ | ~new_C4643_;
  assign new_C4622_ = ~new_C4645_ & new_C4646_;
  assign new_C4623_ = new_C4645_ & ~new_C4646_;
  assign new_C4624_ = ~new_C4592_ & new_C4593_;
  assign new_C4625_ = new_C4592_ & ~new_C4593_;
  assign new_C4626_ = ~new_C4608_ | new_C4618_;
  assign new_C4627_ = new_C4608_ & new_C4618_;
  assign new_C4628_ = ~new_C4608_ & ~new_C4618_;
  assign new_C4629_ = new_C4650_ | new_C4649_;
  assign new_C4630_ = new_C4596_ | new_C4629_;
  assign new_C4631_ = new_C4654_ | new_C4653_;
  assign new_C4632_ = ~new_C4596_ & new_C4631_;
  assign new_C4633_ = new_C4652_ | new_C4651_;
  assign new_C4634_ = new_C4596_ & new_C4633_;
  assign new_C4635_ = new_C4594_ & ~new_C4604_;
  assign new_C4636_ = ~new_C4594_ & new_C4604_;
  assign new_C4637_ = ~new_C4593_ | ~new_C4618_;
  assign new_C4638_ = new_C4604_ & new_C4637_;
  assign new_C4639_ = ~new_C4604_ & ~new_C4638_;
  assign new_C4640_ = new_C4604_ | new_C4637_;
  assign new_C4641_ = ~new_C4594_ & new_C4595_;
  assign new_C4642_ = new_C4594_ & ~new_C4595_;
  assign new_C4643_ = new_C4611_ | new_C4648_;
  assign new_C4644_ = ~new_C4611_ & ~new_C4647_;
  assign new_C4645_ = new_C4594_ | new_C4611_;
  assign new_C4646_ = new_C4594_ | new_C4595_;
  assign new_C4647_ = new_C4611_ & new_C4648_;
  assign new_C4648_ = ~new_C4593_ | ~new_C4618_;
  assign new_C4649_ = new_C4626_ & new_C4646_;
  assign new_C4650_ = ~new_C4626_ & ~new_C4646_;
  assign new_C4651_ = new_C4655_ | new_C4656_;
  assign new_C4652_ = ~new_C4597_ & new_C4611_;
  assign new_C4653_ = new_C4657_ | new_C4658_;
  assign new_C4654_ = new_C4597_ & new_C4611_;
  assign new_C4655_ = ~new_C4597_ & ~new_C4611_;
  assign new_C4656_ = new_C4597_ & ~new_C4611_;
  assign new_C4657_ = new_C4597_ & ~new_C4611_;
  assign new_C4658_ = ~new_C4597_ & new_C4611_;
  assign new_C4659_ = new_E9859_;
  assign new_C4660_ = new_E9926_;
  assign new_C4661_ = new_E9993_;
  assign new_C4662_ = new_F61_;
  assign new_C4663_ = new_F128_;
  assign new_C4664_ = new_F195_;
  assign new_C4665_ = new_C4672_ & new_C4671_;
  assign new_C4666_ = new_C4674_ | new_C4673_;
  assign new_C4667_ = new_C4676_ | new_C4675_;
  assign new_C4668_ = new_C4678_ & new_C4677_;
  assign new_C4669_ = new_C4678_ & new_C4679_;
  assign new_C4670_ = new_C4671_ | new_C4680_;
  assign new_C4671_ = new_C4660_ | new_C4683_;
  assign new_C4672_ = new_C4682_ | new_C4681_;
  assign new_C4673_ = new_C4687_ & new_C4686_;
  assign new_C4674_ = new_C4685_ & new_C4684_;
  assign new_C4675_ = new_C4690_ | new_C4689_;
  assign new_C4676_ = new_C4685_ & new_C4688_;
  assign new_C4677_ = new_C4660_ | new_C4693_;
  assign new_C4678_ = new_C4692_ | new_C4691_;
  assign new_C4679_ = new_C4695_ | new_C4694_;
  assign new_C4680_ = ~new_C4671_ & new_C4697_;
  assign new_C4681_ = ~new_C4673_ & new_C4685_;
  assign new_C4682_ = new_C4673_ & ~new_C4685_;
  assign new_C4683_ = new_C4659_ & ~new_C4660_;
  assign new_C4684_ = ~new_C4706_ | ~new_C4707_;
  assign new_C4685_ = new_C4699_ | new_C4701_;
  assign new_C4686_ = new_C4709_ | new_C4708_;
  assign new_C4687_ = new_C4703_ | new_C4702_;
  assign new_C4688_ = ~new_C4711_ | ~new_C4710_;
  assign new_C4689_ = ~new_C4712_ & new_C4713_;
  assign new_C4690_ = new_C4712_ & ~new_C4713_;
  assign new_C4691_ = ~new_C4659_ & new_C4660_;
  assign new_C4692_ = new_C4659_ & ~new_C4660_;
  assign new_C4693_ = ~new_C4675_ | new_C4685_;
  assign new_C4694_ = new_C4675_ & new_C4685_;
  assign new_C4695_ = ~new_C4675_ & ~new_C4685_;
  assign new_C4696_ = new_C4717_ | new_C4716_;
  assign new_C4697_ = new_C4663_ | new_C4696_;
  assign new_C4698_ = new_C4721_ | new_C4720_;
  assign new_C4699_ = ~new_C4663_ & new_C4698_;
  assign new_C4700_ = new_C4719_ | new_C4718_;
  assign new_C4701_ = new_C4663_ & new_C4700_;
  assign new_C4702_ = new_C4661_ & ~new_C4671_;
  assign new_C4703_ = ~new_C4661_ & new_C4671_;
  assign new_C4704_ = ~new_C4660_ | ~new_C4685_;
  assign new_C4705_ = new_C4671_ & new_C4704_;
  assign new_C4706_ = ~new_C4671_ & ~new_C4705_;
  assign new_C4707_ = new_C4671_ | new_C4704_;
  assign new_C4708_ = ~new_C4661_ & new_C4662_;
  assign new_C4709_ = new_C4661_ & ~new_C4662_;
  assign new_C4710_ = new_C4678_ | new_C4715_;
  assign new_C4711_ = ~new_C4678_ & ~new_C4714_;
  assign new_C4712_ = new_C4661_ | new_C4678_;
  assign new_C4713_ = new_C4661_ | new_C4662_;
  assign new_C4714_ = new_C4678_ & new_C4715_;
  assign new_C4715_ = ~new_C4660_ | ~new_C4685_;
  assign new_C4716_ = new_C4693_ & new_C4713_;
  assign new_C4717_ = ~new_C4693_ & ~new_C4713_;
  assign new_C4718_ = new_C4722_ | new_C4723_;
  assign new_C4719_ = ~new_C4664_ & new_C4678_;
  assign new_C4720_ = new_C4724_ | new_C4725_;
  assign new_C4721_ = new_C4664_ & new_C4678_;
  assign new_C4722_ = ~new_C4664_ & ~new_C4678_;
  assign new_C4723_ = new_C4664_ & ~new_C4678_;
  assign new_C4724_ = new_C4664_ & ~new_C4678_;
  assign new_C4725_ = ~new_C4664_ & new_C4678_;
  assign new_C4726_ = new_F262_;
  assign new_C4727_ = new_F329_;
  assign new_C4728_ = new_F396_;
  assign new_C4729_ = new_F463_;
  assign new_C4730_ = new_F530_;
  assign new_C4731_ = new_F597_;
  assign new_C4732_ = new_C4739_ & new_C4738_;
  assign new_C4733_ = new_C4741_ | new_C4740_;
  assign new_C4734_ = new_C4743_ | new_C4742_;
  assign new_C4735_ = new_C4745_ & new_C4744_;
  assign new_C4736_ = new_C4745_ & new_C4746_;
  assign new_C4737_ = new_C4738_ | new_C4747_;
  assign new_C4738_ = new_C4727_ | new_C4750_;
  assign new_C4739_ = new_C4749_ | new_C4748_;
  assign new_C4740_ = new_C4754_ & new_C4753_;
  assign new_C4741_ = new_C4752_ & new_C4751_;
  assign new_C4742_ = new_C4757_ | new_C4756_;
  assign new_C4743_ = new_C4752_ & new_C4755_;
  assign new_C4744_ = new_C4727_ | new_C4760_;
  assign new_C4745_ = new_C4759_ | new_C4758_;
  assign new_C4746_ = new_C4762_ | new_C4761_;
  assign new_C4747_ = ~new_C4738_ & new_C4764_;
  assign new_C4748_ = ~new_C4740_ & new_C4752_;
  assign new_C4749_ = new_C4740_ & ~new_C4752_;
  assign new_C4750_ = new_C4726_ & ~new_C4727_;
  assign new_C4751_ = ~new_C4773_ | ~new_C4774_;
  assign new_C4752_ = new_C4766_ | new_C4768_;
  assign new_C4753_ = new_C4776_ | new_C4775_;
  assign new_C4754_ = new_C4770_ | new_C4769_;
  assign new_C4755_ = ~new_C4778_ | ~new_C4777_;
  assign new_C4756_ = ~new_C4779_ & new_C4780_;
  assign new_C4757_ = new_C4779_ & ~new_C4780_;
  assign new_C4758_ = ~new_C4726_ & new_C4727_;
  assign new_C4759_ = new_C4726_ & ~new_C4727_;
  assign new_C4760_ = ~new_C4742_ | new_C4752_;
  assign new_C4761_ = new_C4742_ & new_C4752_;
  assign new_C4762_ = ~new_C4742_ & ~new_C4752_;
  assign new_C4763_ = new_C4784_ | new_C4783_;
  assign new_C4764_ = new_C4730_ | new_C4763_;
  assign new_C4765_ = new_C4788_ | new_C4787_;
  assign new_C4766_ = ~new_C4730_ & new_C4765_;
  assign new_C4767_ = new_C4786_ | new_C4785_;
  assign new_C4768_ = new_C4730_ & new_C4767_;
  assign new_C4769_ = new_C4728_ & ~new_C4738_;
  assign new_C4770_ = ~new_C4728_ & new_C4738_;
  assign new_C4771_ = ~new_C4727_ | ~new_C4752_;
  assign new_C4772_ = new_C4738_ & new_C4771_;
  assign new_C4773_ = ~new_C4738_ & ~new_C4772_;
  assign new_C4774_ = new_C4738_ | new_C4771_;
  assign new_C4775_ = ~new_C4728_ & new_C4729_;
  assign new_C4776_ = new_C4728_ & ~new_C4729_;
  assign new_C4777_ = new_C4745_ | new_C4782_;
  assign new_C4778_ = ~new_C4745_ & ~new_C4781_;
  assign new_C4779_ = new_C4728_ | new_C4745_;
  assign new_C4780_ = new_C4728_ | new_C4729_;
  assign new_C4781_ = new_C4745_ & new_C4782_;
  assign new_C4782_ = ~new_C4727_ | ~new_C4752_;
  assign new_C4783_ = new_C4760_ & new_C4780_;
  assign new_C4784_ = ~new_C4760_ & ~new_C4780_;
  assign new_C4785_ = new_C4789_ | new_C4790_;
  assign new_C4786_ = ~new_C4731_ & new_C4745_;
  assign new_C4787_ = new_C4791_ | new_C4792_;
  assign new_C4788_ = new_C4731_ & new_C4745_;
  assign new_C4789_ = ~new_C4731_ & ~new_C4745_;
  assign new_C4790_ = new_C4731_ & ~new_C4745_;
  assign new_C4791_ = new_C4731_ & ~new_C4745_;
  assign new_C4792_ = ~new_C4731_ & new_C4745_;
  assign new_C4793_ = new_F664_;
  assign new_C4794_ = new_F731_;
  assign new_C4795_ = new_F798_;
  assign new_C4796_ = new_F865_;
  assign new_C4797_ = new_F932_;
  assign new_C4798_ = new_F999_;
  assign new_C4799_ = new_C4806_ & new_C4805_;
  assign new_C4800_ = new_C4808_ | new_C4807_;
  assign new_C4801_ = new_C4810_ | new_C4809_;
  assign new_C4802_ = new_C4812_ & new_C4811_;
  assign new_C4803_ = new_C4812_ & new_C4813_;
  assign new_C4804_ = new_C4805_ | new_C4814_;
  assign new_C4805_ = new_C4794_ | new_C4817_;
  assign new_C4806_ = new_C4816_ | new_C4815_;
  assign new_C4807_ = new_C4821_ & new_C4820_;
  assign new_C4808_ = new_C4819_ & new_C4818_;
  assign new_C4809_ = new_C4824_ | new_C4823_;
  assign new_C4810_ = new_C4819_ & new_C4822_;
  assign new_C4811_ = new_C4794_ | new_C4827_;
  assign new_C4812_ = new_C4826_ | new_C4825_;
  assign new_C4813_ = new_C4829_ | new_C4828_;
  assign new_C4814_ = ~new_C4805_ & new_C4831_;
  assign new_C4815_ = ~new_C4807_ & new_C4819_;
  assign new_C4816_ = new_C4807_ & ~new_C4819_;
  assign new_C4817_ = new_C4793_ & ~new_C4794_;
  assign new_C4818_ = ~new_C4840_ | ~new_C4841_;
  assign new_C4819_ = new_C4833_ | new_C4835_;
  assign new_C4820_ = new_C4843_ | new_C4842_;
  assign new_C4821_ = new_C4837_ | new_C4836_;
  assign new_C4822_ = ~new_C4845_ | ~new_C4844_;
  assign new_C4823_ = ~new_C4846_ & new_C4847_;
  assign new_C4824_ = new_C4846_ & ~new_C4847_;
  assign new_C4825_ = ~new_C4793_ & new_C4794_;
  assign new_C4826_ = new_C4793_ & ~new_C4794_;
  assign new_C4827_ = ~new_C4809_ | new_C4819_;
  assign new_C4828_ = new_C4809_ & new_C4819_;
  assign new_C4829_ = ~new_C4809_ & ~new_C4819_;
  assign new_C4830_ = new_C4851_ | new_C4850_;
  assign new_C4831_ = new_C4797_ | new_C4830_;
  assign new_C4832_ = new_C4855_ | new_C4854_;
  assign new_C4833_ = ~new_C4797_ & new_C4832_;
  assign new_C4834_ = new_C4853_ | new_C4852_;
  assign new_C4835_ = new_C4797_ & new_C4834_;
  assign new_C4836_ = new_C4795_ & ~new_C4805_;
  assign new_C4837_ = ~new_C4795_ & new_C4805_;
  assign new_C4838_ = ~new_C4794_ | ~new_C4819_;
  assign new_C4839_ = new_C4805_ & new_C4838_;
  assign new_C4840_ = ~new_C4805_ & ~new_C4839_;
  assign new_C4841_ = new_C4805_ | new_C4838_;
  assign new_C4842_ = ~new_C4795_ & new_C4796_;
  assign new_C4843_ = new_C4795_ & ~new_C4796_;
  assign new_C4844_ = new_C4812_ | new_C4849_;
  assign new_C4845_ = ~new_C4812_ & ~new_C4848_;
  assign new_C4846_ = new_C4795_ | new_C4812_;
  assign new_C4847_ = new_C4795_ | new_C4796_;
  assign new_C4848_ = new_C4812_ & new_C4849_;
  assign new_C4849_ = ~new_C4794_ | ~new_C4819_;
  assign new_C4850_ = new_C4827_ & new_C4847_;
  assign new_C4851_ = ~new_C4827_ & ~new_C4847_;
  assign new_C4852_ = new_C4856_ | new_C4857_;
  assign new_C4853_ = ~new_C4798_ & new_C4812_;
  assign new_C4854_ = new_C4858_ | new_C4859_;
  assign new_C4855_ = new_C4798_ & new_C4812_;
  assign new_C4856_ = ~new_C4798_ & ~new_C4812_;
  assign new_C4857_ = new_C4798_ & ~new_C4812_;
  assign new_C4858_ = new_C4798_ & ~new_C4812_;
  assign new_C4859_ = ~new_C4798_ & new_C4812_;
  assign new_C4860_ = new_F1066_;
  assign new_C4861_ = new_F1133_;
  assign new_C4862_ = new_F1200_;
  assign new_C4863_ = new_F1267_;
  assign new_C4864_ = new_F1334_;
  assign new_C4865_ = new_F1401_;
  assign new_C4866_ = new_C4873_ & new_C4872_;
  assign new_C4867_ = new_C4875_ | new_C4874_;
  assign new_C4868_ = new_C4877_ | new_C4876_;
  assign new_C4869_ = new_C4879_ & new_C4878_;
  assign new_C4870_ = new_C4879_ & new_C4880_;
  assign new_C4871_ = new_C4872_ | new_C4881_;
  assign new_C4872_ = new_C4861_ | new_C4884_;
  assign new_C4873_ = new_C4883_ | new_C4882_;
  assign new_C4874_ = new_C4888_ & new_C4887_;
  assign new_C4875_ = new_C4886_ & new_C4885_;
  assign new_C4876_ = new_C4891_ | new_C4890_;
  assign new_C4877_ = new_C4886_ & new_C4889_;
  assign new_C4878_ = new_C4861_ | new_C4894_;
  assign new_C4879_ = new_C4893_ | new_C4892_;
  assign new_C4880_ = new_C4896_ | new_C4895_;
  assign new_C4881_ = ~new_C4872_ & new_C4898_;
  assign new_C4882_ = ~new_C4874_ & new_C4886_;
  assign new_C4883_ = new_C4874_ & ~new_C4886_;
  assign new_C4884_ = new_C4860_ & ~new_C4861_;
  assign new_C4885_ = ~new_C4907_ | ~new_C4908_;
  assign new_C4886_ = new_C4900_ | new_C4902_;
  assign new_C4887_ = new_C4910_ | new_C4909_;
  assign new_C4888_ = new_C4904_ | new_C4903_;
  assign new_C4889_ = ~new_C4912_ | ~new_C4911_;
  assign new_C4890_ = ~new_C4913_ & new_C4914_;
  assign new_C4891_ = new_C4913_ & ~new_C4914_;
  assign new_C4892_ = ~new_C4860_ & new_C4861_;
  assign new_C4893_ = new_C4860_ & ~new_C4861_;
  assign new_C4894_ = ~new_C4876_ | new_C4886_;
  assign new_C4895_ = new_C4876_ & new_C4886_;
  assign new_C4896_ = ~new_C4876_ & ~new_C4886_;
  assign new_C4897_ = new_C4918_ | new_C4917_;
  assign new_C4898_ = new_C4864_ | new_C4897_;
  assign new_C4899_ = new_C4922_ | new_C4921_;
  assign new_C4900_ = ~new_C4864_ & new_C4899_;
  assign new_C4901_ = new_C4920_ | new_C4919_;
  assign new_C4902_ = new_C4864_ & new_C4901_;
  assign new_C4903_ = new_C4862_ & ~new_C4872_;
  assign new_C4904_ = ~new_C4862_ & new_C4872_;
  assign new_C4905_ = ~new_C4861_ | ~new_C4886_;
  assign new_C4906_ = new_C4872_ & new_C4905_;
  assign new_C4907_ = ~new_C4872_ & ~new_C4906_;
  assign new_C4908_ = new_C4872_ | new_C4905_;
  assign new_C4909_ = ~new_C4862_ & new_C4863_;
  assign new_C4910_ = new_C4862_ & ~new_C4863_;
  assign new_C4911_ = new_C4879_ | new_C4916_;
  assign new_C4912_ = ~new_C4879_ & ~new_C4915_;
  assign new_C4913_ = new_C4862_ | new_C4879_;
  assign new_C4914_ = new_C4862_ | new_C4863_;
  assign new_C4915_ = new_C4879_ & new_C4916_;
  assign new_C4916_ = ~new_C4861_ | ~new_C4886_;
  assign new_C4917_ = new_C4894_ & new_C4914_;
  assign new_C4918_ = ~new_C4894_ & ~new_C4914_;
  assign new_C4919_ = new_C4923_ | new_C4924_;
  assign new_C4920_ = ~new_C4865_ & new_C4879_;
  assign new_C4921_ = new_C4925_ | new_C4926_;
  assign new_C4922_ = new_C4865_ & new_C4879_;
  assign new_C4923_ = ~new_C4865_ & ~new_C4879_;
  assign new_C4924_ = new_C4865_ & ~new_C4879_;
  assign new_C4925_ = new_C4865_ & ~new_C4879_;
  assign new_C4926_ = ~new_C4865_ & new_C4879_;
  assign new_C4927_ = new_D6998_;
  assign new_C4928_ = new_D7062_;
  assign new_C4929_ = new_D7129_;
  assign new_C4930_ = new_D7196_;
  assign new_C4931_ = new_D7263_;
  assign new_C4932_ = new_D7330_;
  assign new_C4933_ = new_C4940_ & new_C4939_;
  assign new_C4934_ = new_C4942_ | new_C4941_;
  assign new_C4935_ = new_C4944_ | new_C4943_;
  assign new_C4936_ = new_C4946_ & new_C4945_;
  assign new_C4937_ = new_C4946_ & new_C4947_;
  assign new_C4938_ = new_C4939_ | new_C4948_;
  assign new_C4939_ = new_C4928_ | new_C4951_;
  assign new_C4940_ = new_C4950_ | new_C4949_;
  assign new_C4941_ = new_C4955_ & new_C4954_;
  assign new_C4942_ = new_C4953_ & new_C4952_;
  assign new_C4943_ = new_C4958_ | new_C4957_;
  assign new_C4944_ = new_C4953_ & new_C4956_;
  assign new_C4945_ = new_C4928_ | new_C4961_;
  assign new_C4946_ = new_C4960_ | new_C4959_;
  assign new_C4947_ = new_C4963_ | new_C4962_;
  assign new_C4948_ = ~new_C4939_ & new_C4965_;
  assign new_C4949_ = ~new_C4941_ & new_C4953_;
  assign new_C4950_ = new_C4941_ & ~new_C4953_;
  assign new_C4951_ = new_C4927_ & ~new_C4928_;
  assign new_C4952_ = ~new_C4974_ | ~new_C4975_;
  assign new_C4953_ = new_C4967_ | new_C4969_;
  assign new_C4954_ = new_C4977_ | new_C4976_;
  assign new_C4955_ = new_C4971_ | new_C4970_;
  assign new_C4956_ = ~new_C4979_ | ~new_C4978_;
  assign new_C4957_ = ~new_C4980_ & new_C4981_;
  assign new_C4958_ = new_C4980_ & ~new_C4981_;
  assign new_C4959_ = ~new_C4927_ & new_C4928_;
  assign new_C4960_ = new_C4927_ & ~new_C4928_;
  assign new_C4961_ = ~new_C4943_ | new_C4953_;
  assign new_C4962_ = new_C4943_ & new_C4953_;
  assign new_C4963_ = ~new_C4943_ & ~new_C4953_;
  assign new_C4964_ = new_C4985_ | new_C4984_;
  assign new_C4965_ = new_C4931_ | new_C4964_;
  assign new_C4966_ = new_C4989_ | new_C4988_;
  assign new_C4967_ = ~new_C4931_ & new_C4966_;
  assign new_C4968_ = new_C4987_ | new_C4986_;
  assign new_C4969_ = new_C4931_ & new_C4968_;
  assign new_C4970_ = new_C4929_ & ~new_C4939_;
  assign new_C4971_ = ~new_C4929_ & new_C4939_;
  assign new_C4972_ = ~new_C4928_ | ~new_C4953_;
  assign new_C4973_ = new_C4939_ & new_C4972_;
  assign new_C4974_ = ~new_C4939_ & ~new_C4973_;
  assign new_C4975_ = new_C4939_ | new_C4972_;
  assign new_C4976_ = ~new_C4929_ & new_C4930_;
  assign new_C4977_ = new_C4929_ & ~new_C4930_;
  assign new_C4978_ = new_C4946_ | new_C4983_;
  assign new_C4979_ = ~new_C4946_ & ~new_C4982_;
  assign new_C4980_ = new_C4929_ | new_C4946_;
  assign new_C4981_ = new_C4929_ | new_C4930_;
  assign new_C4982_ = new_C4946_ & new_C4983_;
  assign new_C4983_ = ~new_C4928_ | ~new_C4953_;
  assign new_C4984_ = new_C4961_ & new_C4981_;
  assign new_C4985_ = ~new_C4961_ & ~new_C4981_;
  assign new_C4986_ = new_C4990_ | new_C4991_;
  assign new_C4987_ = ~new_C4932_ & new_C4946_;
  assign new_C4988_ = new_C4992_ | new_C4993_;
  assign new_C4989_ = new_C4932_ & new_C4946_;
  assign new_C4990_ = ~new_C4932_ & ~new_C4946_;
  assign new_C4991_ = new_C4932_ & ~new_C4946_;
  assign new_C4992_ = new_C4932_ & ~new_C4946_;
  assign new_C4993_ = ~new_C4932_ & new_C4946_;
  assign new_C4994_ = new_D7397_;
  assign new_C4995_ = new_D7464_;
  assign new_C4996_ = new_D7531_;
  assign new_C4997_ = new_D7598_;
  assign new_C4998_ = new_D7665_;
  assign new_C4999_ = new_D7732_;
  assign new_C5000_ = new_C5007_ & new_C5006_;
  assign new_C5001_ = new_C5009_ | new_C5008_;
  assign new_C5002_ = new_C5011_ | new_C5010_;
  assign new_C5003_ = new_C5013_ & new_C5012_;
  assign new_C5004_ = new_C5013_ & new_C5014_;
  assign new_C5005_ = new_C5006_ | new_C5015_;
  assign new_C5006_ = new_C4995_ | new_C5018_;
  assign new_C5007_ = new_C5017_ | new_C5016_;
  assign new_C5008_ = new_C5022_ & new_C5021_;
  assign new_C5009_ = new_C5020_ & new_C5019_;
  assign new_C5010_ = new_C5025_ | new_C5024_;
  assign new_C5011_ = new_C5020_ & new_C5023_;
  assign new_C5012_ = new_C4995_ | new_C5028_;
  assign new_C5013_ = new_C5027_ | new_C5026_;
  assign new_C5014_ = new_C5030_ | new_C5029_;
  assign new_C5015_ = ~new_C5006_ & new_C5032_;
  assign new_C5016_ = ~new_C5008_ & new_C5020_;
  assign new_C5017_ = new_C5008_ & ~new_C5020_;
  assign new_C5018_ = new_C4994_ & ~new_C4995_;
  assign new_C5019_ = ~new_C5041_ | ~new_C5042_;
  assign new_C5020_ = new_C5034_ | new_C5036_;
  assign new_C5021_ = new_C5044_ | new_C5043_;
  assign new_C5022_ = new_C5038_ | new_C5037_;
  assign new_C5023_ = ~new_C5046_ | ~new_C5045_;
  assign new_C5024_ = ~new_C5047_ & new_C5048_;
  assign new_C5025_ = new_C5047_ & ~new_C5048_;
  assign new_C5026_ = ~new_C4994_ & new_C4995_;
  assign new_C5027_ = new_C4994_ & ~new_C4995_;
  assign new_C5028_ = ~new_C5010_ | new_C5020_;
  assign new_C5029_ = new_C5010_ & new_C5020_;
  assign new_C5030_ = ~new_C5010_ & ~new_C5020_;
  assign new_C5031_ = new_C5052_ | new_C5051_;
  assign new_C5032_ = new_C4998_ | new_C5031_;
  assign new_C5033_ = new_C5056_ | new_C5055_;
  assign new_C5034_ = ~new_C4998_ & new_C5033_;
  assign new_C5035_ = new_C5054_ | new_C5053_;
  assign new_C5036_ = new_C4998_ & new_C5035_;
  assign new_C5037_ = new_C4996_ & ~new_C5006_;
  assign new_C5038_ = ~new_C4996_ & new_C5006_;
  assign new_C5039_ = ~new_C4995_ | ~new_C5020_;
  assign new_C5040_ = new_C5006_ & new_C5039_;
  assign new_C5041_ = ~new_C5006_ & ~new_C5040_;
  assign new_C5042_ = new_C5006_ | new_C5039_;
  assign new_C5043_ = ~new_C4996_ & new_C4997_;
  assign new_C5044_ = new_C4996_ & ~new_C4997_;
  assign new_C5045_ = new_C5013_ | new_C5050_;
  assign new_C5046_ = ~new_C5013_ & ~new_C5049_;
  assign new_C5047_ = new_C4996_ | new_C5013_;
  assign new_C5048_ = new_C4996_ | new_C4997_;
  assign new_C5049_ = new_C5013_ & new_C5050_;
  assign new_C5050_ = ~new_C4995_ | ~new_C5020_;
  assign new_C5051_ = new_C5028_ & new_C5048_;
  assign new_C5052_ = ~new_C5028_ & ~new_C5048_;
  assign new_C5053_ = new_C5057_ | new_C5058_;
  assign new_C5054_ = ~new_C4999_ & new_C5013_;
  assign new_C5055_ = new_C5059_ | new_C5060_;
  assign new_C5056_ = new_C4999_ & new_C5013_;
  assign new_C5057_ = ~new_C4999_ & ~new_C5013_;
  assign new_C5058_ = new_C4999_ & ~new_C5013_;
  assign new_C5059_ = new_C4999_ & ~new_C5013_;
  assign new_C5060_ = ~new_C4999_ & new_C5013_;
  assign new_C5061_ = new_D7799_;
  assign new_C5062_ = new_D7866_;
  assign new_C5063_ = new_D7933_;
  assign new_C5064_ = new_D8000_;
  assign new_C5065_ = new_D8067_;
  assign new_C5066_ = new_D8134_;
  assign new_C5067_ = new_C5074_ & new_C5073_;
  assign new_C5068_ = new_C5076_ | new_C5075_;
  assign new_C5069_ = new_C5078_ | new_C5077_;
  assign new_C5070_ = new_C5080_ & new_C5079_;
  assign new_C5071_ = new_C5080_ & new_C5081_;
  assign new_C5072_ = new_C5073_ | new_C5082_;
  assign new_C5073_ = new_C5062_ | new_C5085_;
  assign new_C5074_ = new_C5084_ | new_C5083_;
  assign new_C5075_ = new_C5089_ & new_C5088_;
  assign new_C5076_ = new_C5087_ & new_C5086_;
  assign new_C5077_ = new_C5092_ | new_C5091_;
  assign new_C5078_ = new_C5087_ & new_C5090_;
  assign new_C5079_ = new_C5062_ | new_C5095_;
  assign new_C5080_ = new_C5094_ | new_C5093_;
  assign new_C5081_ = new_C5097_ | new_C5096_;
  assign new_C5082_ = ~new_C5073_ & new_C5099_;
  assign new_C5083_ = ~new_C5075_ & new_C5087_;
  assign new_C5084_ = new_C5075_ & ~new_C5087_;
  assign new_C5085_ = new_C5061_ & ~new_C5062_;
  assign new_C5086_ = ~new_C5108_ | ~new_C5109_;
  assign new_C5087_ = new_C5101_ | new_C5103_;
  assign new_C5088_ = new_C5111_ | new_C5110_;
  assign new_C5089_ = new_C5105_ | new_C5104_;
  assign new_C5090_ = ~new_C5113_ | ~new_C5112_;
  assign new_C5091_ = ~new_C5114_ & new_C5115_;
  assign new_C5092_ = new_C5114_ & ~new_C5115_;
  assign new_C5093_ = ~new_C5061_ & new_C5062_;
  assign new_C5094_ = new_C5061_ & ~new_C5062_;
  assign new_C5095_ = ~new_C5077_ | new_C5087_;
  assign new_C5096_ = new_C5077_ & new_C5087_;
  assign new_C5097_ = ~new_C5077_ & ~new_C5087_;
  assign new_C5098_ = new_C5119_ | new_C5118_;
  assign new_C5099_ = new_C5065_ | new_C5098_;
  assign new_C5100_ = new_C5123_ | new_C5122_;
  assign new_C5101_ = ~new_C5065_ & new_C5100_;
  assign new_C5102_ = new_C5121_ | new_C5120_;
  assign new_C5103_ = new_C5065_ & new_C5102_;
  assign new_C5104_ = new_C5063_ & ~new_C5073_;
  assign new_C5105_ = ~new_C5063_ & new_C5073_;
  assign new_C5106_ = ~new_C5062_ | ~new_C5087_;
  assign new_C5107_ = new_C5073_ & new_C5106_;
  assign new_C5108_ = ~new_C5073_ & ~new_C5107_;
  assign new_C5109_ = new_C5073_ | new_C5106_;
  assign new_C5110_ = ~new_C5063_ & new_C5064_;
  assign new_C5111_ = new_C5063_ & ~new_C5064_;
  assign new_C5112_ = new_C5080_ | new_C5117_;
  assign new_C5113_ = ~new_C5080_ & ~new_C5116_;
  assign new_C5114_ = new_C5063_ | new_C5080_;
  assign new_C5115_ = new_C5063_ | new_C5064_;
  assign new_C5116_ = new_C5080_ & new_C5117_;
  assign new_C5117_ = ~new_C5062_ | ~new_C5087_;
  assign new_C5118_ = new_C5095_ & new_C5115_;
  assign new_C5119_ = ~new_C5095_ & ~new_C5115_;
  assign new_C5120_ = new_C5124_ | new_C5125_;
  assign new_C5121_ = ~new_C5066_ & new_C5080_;
  assign new_C5122_ = new_C5126_ | new_C5127_;
  assign new_C5123_ = new_C5066_ & new_C5080_;
  assign new_C5124_ = ~new_C5066_ & ~new_C5080_;
  assign new_C5125_ = new_C5066_ & ~new_C5080_;
  assign new_C5126_ = new_C5066_ & ~new_C5080_;
  assign new_C5127_ = ~new_C5066_ & new_C5080_;
  assign new_C5128_ = new_D8201_;
  assign new_C5129_ = new_D8268_;
  assign new_C5130_ = new_D8335_;
  assign new_C5131_ = new_D8402_;
  assign new_C5132_ = new_D8469_;
  assign new_C5133_ = new_D8536_;
  assign new_C5134_ = new_C5141_ & new_C5140_;
  assign new_C5135_ = new_C5143_ | new_C5142_;
  assign new_C5136_ = new_C5145_ | new_C5144_;
  assign new_C5137_ = new_C5147_ & new_C5146_;
  assign new_C5138_ = new_C5147_ & new_C5148_;
  assign new_C5139_ = new_C5140_ | new_C5149_;
  assign new_C5140_ = new_C5129_ | new_C5152_;
  assign new_C5141_ = new_C5151_ | new_C5150_;
  assign new_C5142_ = new_C5156_ & new_C5155_;
  assign new_C5143_ = new_C5154_ & new_C5153_;
  assign new_C5144_ = new_C5159_ | new_C5158_;
  assign new_C5145_ = new_C5154_ & new_C5157_;
  assign new_C5146_ = new_C5129_ | new_C5162_;
  assign new_C5147_ = new_C5161_ | new_C5160_;
  assign new_C5148_ = new_C5164_ | new_C5163_;
  assign new_C5149_ = ~new_C5140_ & new_C5166_;
  assign new_C5150_ = ~new_C5142_ & new_C5154_;
  assign new_C5151_ = new_C5142_ & ~new_C5154_;
  assign new_C5152_ = new_C5128_ & ~new_C5129_;
  assign new_C5153_ = ~new_C5175_ | ~new_C5176_;
  assign new_C5154_ = new_C5168_ | new_C5170_;
  assign new_C5155_ = new_C5178_ | new_C5177_;
  assign new_C5156_ = new_C5172_ | new_C5171_;
  assign new_C5157_ = ~new_C5180_ | ~new_C5179_;
  assign new_C5158_ = ~new_C5181_ & new_C5182_;
  assign new_C5159_ = new_C5181_ & ~new_C5182_;
  assign new_C5160_ = ~new_C5128_ & new_C5129_;
  assign new_C5161_ = new_C5128_ & ~new_C5129_;
  assign new_C5162_ = ~new_C5144_ | new_C5154_;
  assign new_C5163_ = new_C5144_ & new_C5154_;
  assign new_C5164_ = ~new_C5144_ & ~new_C5154_;
  assign new_C5165_ = new_C5186_ | new_C5185_;
  assign new_C5166_ = new_C5132_ | new_C5165_;
  assign new_C5167_ = new_C5190_ | new_C5189_;
  assign new_C5168_ = ~new_C5132_ & new_C5167_;
  assign new_C5169_ = new_C5188_ | new_C5187_;
  assign new_C5170_ = new_C5132_ & new_C5169_;
  assign new_C5171_ = new_C5130_ & ~new_C5140_;
  assign new_C5172_ = ~new_C5130_ & new_C5140_;
  assign new_C5173_ = ~new_C5129_ | ~new_C5154_;
  assign new_C5174_ = new_C5140_ & new_C5173_;
  assign new_C5175_ = ~new_C5140_ & ~new_C5174_;
  assign new_C5176_ = new_C5140_ | new_C5173_;
  assign new_C5177_ = ~new_C5130_ & new_C5131_;
  assign new_C5178_ = new_C5130_ & ~new_C5131_;
  assign new_C5179_ = new_C5147_ | new_C5184_;
  assign new_C5180_ = ~new_C5147_ & ~new_C5183_;
  assign new_C5181_ = new_C5130_ | new_C5147_;
  assign new_C5182_ = new_C5130_ | new_C5131_;
  assign new_C5183_ = new_C5147_ & new_C5184_;
  assign new_C5184_ = ~new_C5129_ | ~new_C5154_;
  assign new_C5185_ = new_C5162_ & new_C5182_;
  assign new_C5186_ = ~new_C5162_ & ~new_C5182_;
  assign new_C5187_ = new_C5191_ | new_C5192_;
  assign new_C5188_ = ~new_C5133_ & new_C5147_;
  assign new_C5189_ = new_C5193_ | new_C5194_;
  assign new_C5190_ = new_C5133_ & new_C5147_;
  assign new_C5191_ = ~new_C5133_ & ~new_C5147_;
  assign new_C5192_ = new_C5133_ & ~new_C5147_;
  assign new_C5193_ = new_C5133_ & ~new_C5147_;
  assign new_C5194_ = ~new_C5133_ & new_C5147_;
  assign new_C5195_ = new_D8603_;
  assign new_C5196_ = new_D8670_;
  assign new_C5197_ = new_D8737_;
  assign new_C5198_ = new_D8804_;
  assign new_C5199_ = new_D8871_;
  assign new_C5200_ = new_D8938_;
  assign new_C5201_ = new_C5208_ & new_C5207_;
  assign new_C5202_ = new_C5210_ | new_C5209_;
  assign new_C5203_ = new_C5212_ | new_C5211_;
  assign new_C5204_ = new_C5214_ & new_C5213_;
  assign new_C5205_ = new_C5214_ & new_C5215_;
  assign new_C5206_ = new_C5207_ | new_C5216_;
  assign new_C5207_ = new_C5196_ | new_C5219_;
  assign new_C5208_ = new_C5218_ | new_C5217_;
  assign new_C5209_ = new_C5223_ & new_C5222_;
  assign new_C5210_ = new_C5221_ & new_C5220_;
  assign new_C5211_ = new_C5226_ | new_C5225_;
  assign new_C5212_ = new_C5221_ & new_C5224_;
  assign new_C5213_ = new_C5196_ | new_C5229_;
  assign new_C5214_ = new_C5228_ | new_C5227_;
  assign new_C5215_ = new_C5231_ | new_C5230_;
  assign new_C5216_ = ~new_C5207_ & new_C5233_;
  assign new_C5217_ = ~new_C5209_ & new_C5221_;
  assign new_C5218_ = new_C5209_ & ~new_C5221_;
  assign new_C5219_ = new_C5195_ & ~new_C5196_;
  assign new_C5220_ = ~new_C5242_ | ~new_C5243_;
  assign new_C5221_ = new_C5235_ | new_C5237_;
  assign new_C5222_ = new_C5245_ | new_C5244_;
  assign new_C5223_ = new_C5239_ | new_C5238_;
  assign new_C5224_ = ~new_C5247_ | ~new_C5246_;
  assign new_C5225_ = ~new_C5248_ & new_C5249_;
  assign new_C5226_ = new_C5248_ & ~new_C5249_;
  assign new_C5227_ = ~new_C5195_ & new_C5196_;
  assign new_C5228_ = new_C5195_ & ~new_C5196_;
  assign new_C5229_ = ~new_C5211_ | new_C5221_;
  assign new_C5230_ = new_C5211_ & new_C5221_;
  assign new_C5231_ = ~new_C5211_ & ~new_C5221_;
  assign new_C5232_ = new_C5253_ | new_C5252_;
  assign new_C5233_ = new_C5199_ | new_C5232_;
  assign new_C5234_ = new_C5257_ | new_C5256_;
  assign new_C5235_ = ~new_C5199_ & new_C5234_;
  assign new_C5236_ = new_C5255_ | new_C5254_;
  assign new_C5237_ = new_C5199_ & new_C5236_;
  assign new_C5238_ = new_C5197_ & ~new_C5207_;
  assign new_C5239_ = ~new_C5197_ & new_C5207_;
  assign new_C5240_ = ~new_C5196_ | ~new_C5221_;
  assign new_C5241_ = new_C5207_ & new_C5240_;
  assign new_C5242_ = ~new_C5207_ & ~new_C5241_;
  assign new_C5243_ = new_C5207_ | new_C5240_;
  assign new_C5244_ = ~new_C5197_ & new_C5198_;
  assign new_C5245_ = new_C5197_ & ~new_C5198_;
  assign new_C5246_ = new_C5214_ | new_C5251_;
  assign new_C5247_ = ~new_C5214_ & ~new_C5250_;
  assign new_C5248_ = new_C5197_ | new_C5214_;
  assign new_C5249_ = new_C5197_ | new_C5198_;
  assign new_C5250_ = new_C5214_ & new_C5251_;
  assign new_C5251_ = ~new_C5196_ | ~new_C5221_;
  assign new_C5252_ = new_C5229_ & new_C5249_;
  assign new_C5253_ = ~new_C5229_ & ~new_C5249_;
  assign new_C5254_ = new_C5258_ | new_C5259_;
  assign new_C5255_ = ~new_C5200_ & new_C5214_;
  assign new_C5256_ = new_C5260_ | new_C5261_;
  assign new_C5257_ = new_C5200_ & new_C5214_;
  assign new_C5258_ = ~new_C5200_ & ~new_C5214_;
  assign new_C5259_ = new_C5200_ & ~new_C5214_;
  assign new_C5260_ = new_C5200_ & ~new_C5214_;
  assign new_C5261_ = ~new_C5200_ & new_C5214_;
  assign new_C5262_ = new_D9005_;
  assign new_C5263_ = new_D9072_;
  assign new_C5264_ = new_D9139_;
  assign new_C5265_ = new_D9206_;
  assign new_C5266_ = new_D9273_;
  assign new_C5267_ = new_D9340_;
  assign new_C5268_ = new_C5275_ & new_C5274_;
  assign new_C5269_ = new_C5277_ | new_C5276_;
  assign new_C5270_ = new_C5279_ | new_C5278_;
  assign new_C5271_ = new_C5281_ & new_C5280_;
  assign new_C5272_ = new_C5281_ & new_C5282_;
  assign new_C5273_ = new_C5274_ | new_C5283_;
  assign new_C5274_ = new_C5263_ | new_C5286_;
  assign new_C5275_ = new_C5285_ | new_C5284_;
  assign new_C5276_ = new_C5290_ & new_C5289_;
  assign new_C5277_ = new_C5288_ & new_C5287_;
  assign new_C5278_ = new_C5293_ | new_C5292_;
  assign new_C5279_ = new_C5288_ & new_C5291_;
  assign new_C5280_ = new_C5263_ | new_C5296_;
  assign new_C5281_ = new_C5295_ | new_C5294_;
  assign new_C5282_ = new_C5298_ | new_C5297_;
  assign new_C5283_ = ~new_C5274_ & new_C5300_;
  assign new_C5284_ = ~new_C5276_ & new_C5288_;
  assign new_C5285_ = new_C5276_ & ~new_C5288_;
  assign new_C5286_ = new_C5262_ & ~new_C5263_;
  assign new_C5287_ = ~new_C5309_ | ~new_C5310_;
  assign new_C5288_ = new_C5302_ | new_C5304_;
  assign new_C5289_ = new_C5312_ | new_C5311_;
  assign new_C5290_ = new_C5306_ | new_C5305_;
  assign new_C5291_ = ~new_C5314_ | ~new_C5313_;
  assign new_C5292_ = ~new_C5315_ & new_C5316_;
  assign new_C5293_ = new_C5315_ & ~new_C5316_;
  assign new_C5294_ = ~new_C5262_ & new_C5263_;
  assign new_C5295_ = new_C5262_ & ~new_C5263_;
  assign new_C5296_ = ~new_C5278_ | new_C5288_;
  assign new_C5297_ = new_C5278_ & new_C5288_;
  assign new_C5298_ = ~new_C5278_ & ~new_C5288_;
  assign new_C5299_ = new_C5320_ | new_C5319_;
  assign new_C5300_ = new_C5266_ | new_C5299_;
  assign new_C5301_ = new_C5324_ | new_C5323_;
  assign new_C5302_ = ~new_C5266_ & new_C5301_;
  assign new_C5303_ = new_C5322_ | new_C5321_;
  assign new_C5304_ = new_C5266_ & new_C5303_;
  assign new_C5305_ = new_C5264_ & ~new_C5274_;
  assign new_C5306_ = ~new_C5264_ & new_C5274_;
  assign new_C5307_ = ~new_C5263_ | ~new_C5288_;
  assign new_C5308_ = new_C5274_ & new_C5307_;
  assign new_C5309_ = ~new_C5274_ & ~new_C5308_;
  assign new_C5310_ = new_C5274_ | new_C5307_;
  assign new_C5311_ = ~new_C5264_ & new_C5265_;
  assign new_C5312_ = new_C5264_ & ~new_C5265_;
  assign new_C5313_ = new_C5281_ | new_C5318_;
  assign new_C5314_ = ~new_C5281_ & ~new_C5317_;
  assign new_C5315_ = new_C5264_ | new_C5281_;
  assign new_C5316_ = new_C5264_ | new_C5265_;
  assign new_C5317_ = new_C5281_ & new_C5318_;
  assign new_C5318_ = ~new_C5263_ | ~new_C5288_;
  assign new_C5319_ = new_C5296_ & new_C5316_;
  assign new_C5320_ = ~new_C5296_ & ~new_C5316_;
  assign new_C5321_ = new_C5325_ | new_C5326_;
  assign new_C5322_ = ~new_C5267_ & new_C5281_;
  assign new_C5323_ = new_C5327_ | new_C5328_;
  assign new_C5324_ = new_C5267_ & new_C5281_;
  assign new_C5325_ = ~new_C5267_ & ~new_C5281_;
  assign new_C5326_ = new_C5267_ & ~new_C5281_;
  assign new_C5327_ = new_C5267_ & ~new_C5281_;
  assign new_C5328_ = ~new_C5267_ & new_C5281_;
  assign new_C5329_ = new_D9407_;
  assign new_C5330_ = new_D9474_;
  assign new_C5331_ = new_D9541_;
  assign new_C5332_ = new_D9608_;
  assign new_C5333_ = new_D9675_;
  assign new_C5334_ = new_D9742_;
  assign new_C5335_ = new_C5342_ & new_C5341_;
  assign new_C5336_ = new_C5344_ | new_C5343_;
  assign new_C5337_ = new_C5346_ | new_C5345_;
  assign new_C5338_ = new_C5348_ & new_C5347_;
  assign new_C5339_ = new_C5348_ & new_C5349_;
  assign new_C5340_ = new_C5341_ | new_C5350_;
  assign new_C5341_ = new_C5330_ | new_C5353_;
  assign new_C5342_ = new_C5352_ | new_C5351_;
  assign new_C5343_ = new_C5357_ & new_C5356_;
  assign new_C5344_ = new_C5355_ & new_C5354_;
  assign new_C5345_ = new_C5360_ | new_C5359_;
  assign new_C5346_ = new_C5355_ & new_C5358_;
  assign new_C5347_ = new_C5330_ | new_C5363_;
  assign new_C5348_ = new_C5362_ | new_C5361_;
  assign new_C5349_ = new_C5365_ | new_C5364_;
  assign new_C5350_ = ~new_C5341_ & new_C5367_;
  assign new_C5351_ = ~new_C5343_ & new_C5355_;
  assign new_C5352_ = new_C5343_ & ~new_C5355_;
  assign new_C5353_ = new_C5329_ & ~new_C5330_;
  assign new_C5354_ = ~new_C5376_ | ~new_C5377_;
  assign new_C5355_ = new_C5369_ | new_C5371_;
  assign new_C5356_ = new_C5379_ | new_C5378_;
  assign new_C5357_ = new_C5373_ | new_C5372_;
  assign new_C5358_ = ~new_C5381_ | ~new_C5380_;
  assign new_C5359_ = ~new_C5382_ & new_C5383_;
  assign new_C5360_ = new_C5382_ & ~new_C5383_;
  assign new_C5361_ = ~new_C5329_ & new_C5330_;
  assign new_C5362_ = new_C5329_ & ~new_C5330_;
  assign new_C5363_ = ~new_C5345_ | new_C5355_;
  assign new_C5364_ = new_C5345_ & new_C5355_;
  assign new_C5365_ = ~new_C5345_ & ~new_C5355_;
  assign new_C5366_ = new_C5387_ | new_C5386_;
  assign new_C5367_ = new_C5333_ | new_C5366_;
  assign new_C5368_ = new_C5391_ | new_C5390_;
  assign new_C5369_ = ~new_C5333_ & new_C5368_;
  assign new_C5370_ = new_C5389_ | new_C5388_;
  assign new_C5371_ = new_C5333_ & new_C5370_;
  assign new_C5372_ = new_C5331_ & ~new_C5341_;
  assign new_C5373_ = ~new_C5331_ & new_C5341_;
  assign new_C5374_ = ~new_C5330_ | ~new_C5355_;
  assign new_C5375_ = new_C5341_ & new_C5374_;
  assign new_C5376_ = ~new_C5341_ & ~new_C5375_;
  assign new_C5377_ = new_C5341_ | new_C5374_;
  assign new_C5378_ = ~new_C5331_ & new_C5332_;
  assign new_C5379_ = new_C5331_ & ~new_C5332_;
  assign new_C5380_ = new_C5348_ | new_C5385_;
  assign new_C5381_ = ~new_C5348_ & ~new_C5384_;
  assign new_C5382_ = new_C5331_ | new_C5348_;
  assign new_C5383_ = new_C5331_ | new_C5332_;
  assign new_C5384_ = new_C5348_ & new_C5385_;
  assign new_C5385_ = ~new_C5330_ | ~new_C5355_;
  assign new_C5386_ = new_C5363_ & new_C5383_;
  assign new_C5387_ = ~new_C5363_ & ~new_C5383_;
  assign new_C5388_ = new_C5392_ | new_C5393_;
  assign new_C5389_ = ~new_C5334_ & new_C5348_;
  assign new_C5390_ = new_C5394_ | new_C5395_;
  assign new_C5391_ = new_C5334_ & new_C5348_;
  assign new_C5392_ = ~new_C5334_ & ~new_C5348_;
  assign new_C5393_ = new_C5334_ & ~new_C5348_;
  assign new_C5394_ = new_C5334_ & ~new_C5348_;
  assign new_C5395_ = ~new_C5334_ & new_C5348_;
  assign new_C5396_ = new_D9809_;
  assign new_C5397_ = new_D9876_;
  assign new_C5398_ = new_D9943_;
  assign new_C5399_ = new_E11_;
  assign new_C5400_ = new_E78_;
  assign new_C5401_ = new_E145_;
  assign new_C5402_ = new_C5409_ & new_C5408_;
  assign new_C5403_ = new_C5411_ | new_C5410_;
  assign new_C5404_ = new_C5413_ | new_C5412_;
  assign new_C5405_ = new_C5415_ & new_C5414_;
  assign new_C5406_ = new_C5415_ & new_C5416_;
  assign new_C5407_ = new_C5408_ | new_C5417_;
  assign new_C5408_ = new_C5397_ | new_C5420_;
  assign new_C5409_ = new_C5419_ | new_C5418_;
  assign new_C5410_ = new_C5424_ & new_C5423_;
  assign new_C5411_ = new_C5422_ & new_C5421_;
  assign new_C5412_ = new_C5427_ | new_C5426_;
  assign new_C5413_ = new_C5422_ & new_C5425_;
  assign new_C5414_ = new_C5397_ | new_C5430_;
  assign new_C5415_ = new_C5429_ | new_C5428_;
  assign new_C5416_ = new_C5432_ | new_C5431_;
  assign new_C5417_ = ~new_C5408_ & new_C5434_;
  assign new_C5418_ = ~new_C5410_ & new_C5422_;
  assign new_C5419_ = new_C5410_ & ~new_C5422_;
  assign new_C5420_ = new_C5396_ & ~new_C5397_;
  assign new_C5421_ = ~new_C5443_ | ~new_C5444_;
  assign new_C5422_ = new_C5436_ | new_C5438_;
  assign new_C5423_ = new_C5446_ | new_C5445_;
  assign new_C5424_ = new_C5440_ | new_C5439_;
  assign new_C5425_ = ~new_C5448_ | ~new_C5447_;
  assign new_C5426_ = ~new_C5449_ & new_C5450_;
  assign new_C5427_ = new_C5449_ & ~new_C5450_;
  assign new_C5428_ = ~new_C5396_ & new_C5397_;
  assign new_C5429_ = new_C5396_ & ~new_C5397_;
  assign new_C5430_ = ~new_C5412_ | new_C5422_;
  assign new_C5431_ = new_C5412_ & new_C5422_;
  assign new_C5432_ = ~new_C5412_ & ~new_C5422_;
  assign new_C5433_ = new_C5454_ | new_C5453_;
  assign new_C5434_ = new_C5400_ | new_C5433_;
  assign new_C5435_ = new_C5458_ | new_C5457_;
  assign new_C5436_ = ~new_C5400_ & new_C5435_;
  assign new_C5437_ = new_C5456_ | new_C5455_;
  assign new_C5438_ = new_C5400_ & new_C5437_;
  assign new_C5439_ = new_C5398_ & ~new_C5408_;
  assign new_C5440_ = ~new_C5398_ & new_C5408_;
  assign new_C5441_ = ~new_C5397_ | ~new_C5422_;
  assign new_C5442_ = new_C5408_ & new_C5441_;
  assign new_C5443_ = ~new_C5408_ & ~new_C5442_;
  assign new_C5444_ = new_C5408_ | new_C5441_;
  assign new_C5445_ = ~new_C5398_ & new_C5399_;
  assign new_C5446_ = new_C5398_ & ~new_C5399_;
  assign new_C5447_ = new_C5415_ | new_C5452_;
  assign new_C5448_ = ~new_C5415_ & ~new_C5451_;
  assign new_C5449_ = new_C5398_ | new_C5415_;
  assign new_C5450_ = new_C5398_ | new_C5399_;
  assign new_C5451_ = new_C5415_ & new_C5452_;
  assign new_C5452_ = ~new_C5397_ | ~new_C5422_;
  assign new_C5453_ = new_C5430_ & new_C5450_;
  assign new_C5454_ = ~new_C5430_ & ~new_C5450_;
  assign new_C5455_ = new_C5459_ | new_C5460_;
  assign new_C5456_ = ~new_C5401_ & new_C5415_;
  assign new_C5457_ = new_C5461_ | new_C5462_;
  assign new_C5458_ = new_C5401_ & new_C5415_;
  assign new_C5459_ = ~new_C5401_ & ~new_C5415_;
  assign new_C5460_ = new_C5401_ & ~new_C5415_;
  assign new_C5461_ = new_C5401_ & ~new_C5415_;
  assign new_C5462_ = ~new_C5401_ & new_C5415_;
  assign new_C5463_ = new_E212_;
  assign new_C5464_ = new_E279_;
  assign new_C5465_ = new_E346_;
  assign new_C5466_ = new_E413_;
  assign new_C5467_ = new_E480_;
  assign new_C5468_ = new_E547_;
  assign new_C5469_ = new_C5476_ & new_C5475_;
  assign new_C5470_ = new_C5478_ | new_C5477_;
  assign new_C5471_ = new_C5480_ | new_C5479_;
  assign new_C5472_ = new_C5482_ & new_C5481_;
  assign new_C5473_ = new_C5482_ & new_C5483_;
  assign new_C5474_ = new_C5475_ | new_C5484_;
  assign new_C5475_ = new_C5464_ | new_C5487_;
  assign new_C5476_ = new_C5486_ | new_C5485_;
  assign new_C5477_ = new_C5491_ & new_C5490_;
  assign new_C5478_ = new_C5489_ & new_C5488_;
  assign new_C5479_ = new_C5494_ | new_C5493_;
  assign new_C5480_ = new_C5489_ & new_C5492_;
  assign new_C5481_ = new_C5464_ | new_C5497_;
  assign new_C5482_ = new_C5496_ | new_C5495_;
  assign new_C5483_ = new_C5499_ | new_C5498_;
  assign new_C5484_ = ~new_C5475_ & new_C5501_;
  assign new_C5485_ = ~new_C5477_ & new_C5489_;
  assign new_C5486_ = new_C5477_ & ~new_C5489_;
  assign new_C5487_ = new_C5463_ & ~new_C5464_;
  assign new_C5488_ = ~new_C5510_ | ~new_C5511_;
  assign new_C5489_ = new_C5503_ | new_C5505_;
  assign new_C5490_ = new_C5513_ | new_C5512_;
  assign new_C5491_ = new_C5507_ | new_C5506_;
  assign new_C5492_ = ~new_C5515_ | ~new_C5514_;
  assign new_C5493_ = ~new_C5516_ & new_C5517_;
  assign new_C5494_ = new_C5516_ & ~new_C5517_;
  assign new_C5495_ = ~new_C5463_ & new_C5464_;
  assign new_C5496_ = new_C5463_ & ~new_C5464_;
  assign new_C5497_ = ~new_C5479_ | new_C5489_;
  assign new_C5498_ = new_C5479_ & new_C5489_;
  assign new_C5499_ = ~new_C5479_ & ~new_C5489_;
  assign new_C5500_ = new_C5521_ | new_C5520_;
  assign new_C5501_ = new_C5467_ | new_C5500_;
  assign new_C5502_ = new_C5525_ | new_C5524_;
  assign new_C5503_ = ~new_C5467_ & new_C5502_;
  assign new_C5504_ = new_C5523_ | new_C5522_;
  assign new_C5505_ = new_C5467_ & new_C5504_;
  assign new_C5506_ = new_C5465_ & ~new_C5475_;
  assign new_C5507_ = ~new_C5465_ & new_C5475_;
  assign new_C5508_ = ~new_C5464_ | ~new_C5489_;
  assign new_C5509_ = new_C5475_ & new_C5508_;
  assign new_C5510_ = ~new_C5475_ & ~new_C5509_;
  assign new_C5511_ = new_C5475_ | new_C5508_;
  assign new_C5512_ = ~new_C5465_ & new_C5466_;
  assign new_C5513_ = new_C5465_ & ~new_C5466_;
  assign new_C5514_ = new_C5482_ | new_C5519_;
  assign new_C5515_ = ~new_C5482_ & ~new_C5518_;
  assign new_C5516_ = new_C5465_ | new_C5482_;
  assign new_C5517_ = new_C5465_ | new_C5466_;
  assign new_C5518_ = new_C5482_ & new_C5519_;
  assign new_C5519_ = ~new_C5464_ | ~new_C5489_;
  assign new_C5520_ = new_C5497_ & new_C5517_;
  assign new_C5521_ = ~new_C5497_ & ~new_C5517_;
  assign new_C5522_ = new_C5526_ | new_C5527_;
  assign new_C5523_ = ~new_C5468_ & new_C5482_;
  assign new_C5524_ = new_C5528_ | new_C5529_;
  assign new_C5525_ = new_C5468_ & new_C5482_;
  assign new_C5526_ = ~new_C5468_ & ~new_C5482_;
  assign new_C5527_ = new_C5468_ & ~new_C5482_;
  assign new_C5528_ = new_C5468_ & ~new_C5482_;
  assign new_C5529_ = ~new_C5468_ & new_C5482_;
  assign new_C5530_ = new_E614_;
  assign new_C5531_ = new_E681_;
  assign new_C5532_ = new_E748_;
  assign new_C5533_ = new_E815_;
  assign new_C5534_ = new_E882_;
  assign new_C5535_ = new_E949_;
  assign new_C5536_ = new_C5543_ & new_C5542_;
  assign new_C5537_ = new_C5545_ | new_C5544_;
  assign new_C5538_ = new_C5547_ | new_C5546_;
  assign new_C5539_ = new_C5549_ & new_C5548_;
  assign new_C5540_ = new_C5549_ & new_C5550_;
  assign new_C5541_ = new_C5542_ | new_C5551_;
  assign new_C5542_ = new_C5531_ | new_C5554_;
  assign new_C5543_ = new_C5553_ | new_C5552_;
  assign new_C5544_ = new_C5558_ & new_C5557_;
  assign new_C5545_ = new_C5556_ & new_C5555_;
  assign new_C5546_ = new_C5561_ | new_C5560_;
  assign new_C5547_ = new_C5556_ & new_C5559_;
  assign new_C5548_ = new_C5531_ | new_C5564_;
  assign new_C5549_ = new_C5563_ | new_C5562_;
  assign new_C5550_ = new_C5566_ | new_C5565_;
  assign new_C5551_ = ~new_C5542_ & new_C5568_;
  assign new_C5552_ = ~new_C5544_ & new_C5556_;
  assign new_C5553_ = new_C5544_ & ~new_C5556_;
  assign new_C5554_ = new_C5530_ & ~new_C5531_;
  assign new_C5555_ = ~new_C5577_ | ~new_C5578_;
  assign new_C5556_ = new_C5570_ | new_C5572_;
  assign new_C5557_ = new_C5580_ | new_C5579_;
  assign new_C5558_ = new_C5574_ | new_C5573_;
  assign new_C5559_ = ~new_C5582_ | ~new_C5581_;
  assign new_C5560_ = ~new_C5583_ & new_C5584_;
  assign new_C5561_ = new_C5583_ & ~new_C5584_;
  assign new_C5562_ = ~new_C5530_ & new_C5531_;
  assign new_C5563_ = new_C5530_ & ~new_C5531_;
  assign new_C5564_ = ~new_C5546_ | new_C5556_;
  assign new_C5565_ = new_C5546_ & new_C5556_;
  assign new_C5566_ = ~new_C5546_ & ~new_C5556_;
  assign new_C5567_ = new_C5588_ | new_C5587_;
  assign new_C5568_ = new_C5534_ | new_C5567_;
  assign new_C5569_ = new_C5592_ | new_C5591_;
  assign new_C5570_ = ~new_C5534_ & new_C5569_;
  assign new_C5571_ = new_C5590_ | new_C5589_;
  assign new_C5572_ = new_C5534_ & new_C5571_;
  assign new_C5573_ = new_C5532_ & ~new_C5542_;
  assign new_C5574_ = ~new_C5532_ & new_C5542_;
  assign new_C5575_ = ~new_C5531_ | ~new_C5556_;
  assign new_C5576_ = new_C5542_ & new_C5575_;
  assign new_C5577_ = ~new_C5542_ & ~new_C5576_;
  assign new_C5578_ = new_C5542_ | new_C5575_;
  assign new_C5579_ = ~new_C5532_ & new_C5533_;
  assign new_C5580_ = new_C5532_ & ~new_C5533_;
  assign new_C5581_ = new_C5549_ | new_C5586_;
  assign new_C5582_ = ~new_C5549_ & ~new_C5585_;
  assign new_C5583_ = new_C5532_ | new_C5549_;
  assign new_C5584_ = new_C5532_ | new_C5533_;
  assign new_C5585_ = new_C5549_ & new_C5586_;
  assign new_C5586_ = ~new_C5531_ | ~new_C5556_;
  assign new_C5587_ = new_C5564_ & new_C5584_;
  assign new_C5588_ = ~new_C5564_ & ~new_C5584_;
  assign new_C5589_ = new_C5593_ | new_C5594_;
  assign new_C5590_ = ~new_C5535_ & new_C5549_;
  assign new_C5591_ = new_C5595_ | new_C5596_;
  assign new_C5592_ = new_C5535_ & new_C5549_;
  assign new_C5593_ = ~new_C5535_ & ~new_C5549_;
  assign new_C5594_ = new_C5535_ & ~new_C5549_;
  assign new_C5595_ = new_C5535_ & ~new_C5549_;
  assign new_C5596_ = ~new_C5535_ & new_C5549_;
  assign new_C5597_ = new_E1016_;
  assign new_C5598_ = new_E1083_;
  assign new_C5599_ = new_E1150_;
  assign new_C5600_ = new_E1217_;
  assign new_C5601_ = new_E1284_;
  assign new_C5602_ = new_E1351_;
  assign new_C5603_ = new_C5610_ & new_C5609_;
  assign new_C5604_ = new_C5612_ | new_C5611_;
  assign new_C5605_ = new_C5614_ | new_C5613_;
  assign new_C5606_ = new_C5616_ & new_C5615_;
  assign new_C5607_ = new_C5616_ & new_C5617_;
  assign new_C5608_ = new_C5609_ | new_C5618_;
  assign new_C5609_ = new_C5598_ | new_C5621_;
  assign new_C5610_ = new_C5620_ | new_C5619_;
  assign new_C5611_ = new_C5625_ & new_C5624_;
  assign new_C5612_ = new_C5623_ & new_C5622_;
  assign new_C5613_ = new_C5628_ | new_C5627_;
  assign new_C5614_ = new_C5623_ & new_C5626_;
  assign new_C5615_ = new_C5598_ | new_C5631_;
  assign new_C5616_ = new_C5630_ | new_C5629_;
  assign new_C5617_ = new_C5633_ | new_C5632_;
  assign new_C5618_ = ~new_C5609_ & new_C5635_;
  assign new_C5619_ = ~new_C5611_ & new_C5623_;
  assign new_C5620_ = new_C5611_ & ~new_C5623_;
  assign new_C5621_ = new_C5597_ & ~new_C5598_;
  assign new_C5622_ = ~new_C5644_ | ~new_C5645_;
  assign new_C5623_ = new_C5637_ | new_C5639_;
  assign new_C5624_ = new_C5647_ | new_C5646_;
  assign new_C5625_ = new_C5641_ | new_C5640_;
  assign new_C5626_ = ~new_C5649_ | ~new_C5648_;
  assign new_C5627_ = ~new_C5650_ & new_C5651_;
  assign new_C5628_ = new_C5650_ & ~new_C5651_;
  assign new_C5629_ = ~new_C5597_ & new_C5598_;
  assign new_C5630_ = new_C5597_ & ~new_C5598_;
  assign new_C5631_ = ~new_C5613_ | new_C5623_;
  assign new_C5632_ = new_C5613_ & new_C5623_;
  assign new_C5633_ = ~new_C5613_ & ~new_C5623_;
  assign new_C5634_ = new_C5655_ | new_C5654_;
  assign new_C5635_ = new_C5601_ | new_C5634_;
  assign new_C5636_ = new_C5659_ | new_C5658_;
  assign new_C5637_ = ~new_C5601_ & new_C5636_;
  assign new_C5638_ = new_C5657_ | new_C5656_;
  assign new_C5639_ = new_C5601_ & new_C5638_;
  assign new_C5640_ = new_C5599_ & ~new_C5609_;
  assign new_C5641_ = ~new_C5599_ & new_C5609_;
  assign new_C5642_ = ~new_C5598_ | ~new_C5623_;
  assign new_C5643_ = new_C5609_ & new_C5642_;
  assign new_C5644_ = ~new_C5609_ & ~new_C5643_;
  assign new_C5645_ = new_C5609_ | new_C5642_;
  assign new_C5646_ = ~new_C5599_ & new_C5600_;
  assign new_C5647_ = new_C5599_ & ~new_C5600_;
  assign new_C5648_ = new_C5616_ | new_C5653_;
  assign new_C5649_ = ~new_C5616_ & ~new_C5652_;
  assign new_C5650_ = new_C5599_ | new_C5616_;
  assign new_C5651_ = new_C5599_ | new_C5600_;
  assign new_C5652_ = new_C5616_ & new_C5653_;
  assign new_C5653_ = ~new_C5598_ | ~new_C5623_;
  assign new_C5654_ = new_C5631_ & new_C5651_;
  assign new_C5655_ = ~new_C5631_ & ~new_C5651_;
  assign new_C5656_ = new_C5660_ | new_C5661_;
  assign new_C5657_ = ~new_C5602_ & new_C5616_;
  assign new_C5658_ = new_C5662_ | new_C5663_;
  assign new_C5659_ = new_C5602_ & new_C5616_;
  assign new_C5660_ = ~new_C5602_ & ~new_C5616_;
  assign new_C5661_ = new_C5602_ & ~new_C5616_;
  assign new_C5662_ = new_C5602_ & ~new_C5616_;
  assign new_C5663_ = ~new_C5602_ & new_C5616_;
  assign new_C5664_ = new_E1418_;
  assign new_C5665_ = new_E1485_;
  assign new_C5666_ = new_E1552_;
  assign new_C5667_ = new_E1619_;
  assign new_C5668_ = new_E1686_;
  assign new_C5669_ = new_E1753_;
  assign new_C5670_ = new_C5677_ & new_C5676_;
  assign new_C5671_ = new_C5679_ | new_C5678_;
  assign new_C5672_ = new_C5681_ | new_C5680_;
  assign new_C5673_ = new_C5683_ & new_C5682_;
  assign new_C5674_ = new_C5683_ & new_C5684_;
  assign new_C5675_ = new_C5676_ | new_C5685_;
  assign new_C5676_ = new_C5665_ | new_C5688_;
  assign new_C5677_ = new_C5687_ | new_C5686_;
  assign new_C5678_ = new_C5692_ & new_C5691_;
  assign new_C5679_ = new_C5690_ & new_C5689_;
  assign new_C5680_ = new_C5695_ | new_C5694_;
  assign new_C5681_ = new_C5690_ & new_C5693_;
  assign new_C5682_ = new_C5665_ | new_C5698_;
  assign new_C5683_ = new_C5697_ | new_C5696_;
  assign new_C5684_ = new_C5700_ | new_C5699_;
  assign new_C5685_ = ~new_C5676_ & new_C5702_;
  assign new_C5686_ = ~new_C5678_ & new_C5690_;
  assign new_C5687_ = new_C5678_ & ~new_C5690_;
  assign new_C5688_ = new_C5664_ & ~new_C5665_;
  assign new_C5689_ = ~new_C5711_ | ~new_C5712_;
  assign new_C5690_ = new_C5704_ | new_C5706_;
  assign new_C5691_ = new_C5714_ | new_C5713_;
  assign new_C5692_ = new_C5708_ | new_C5707_;
  assign new_C5693_ = ~new_C5716_ | ~new_C5715_;
  assign new_C5694_ = ~new_C5717_ & new_C5718_;
  assign new_C5695_ = new_C5717_ & ~new_C5718_;
  assign new_C5696_ = ~new_C5664_ & new_C5665_;
  assign new_C5697_ = new_C5664_ & ~new_C5665_;
  assign new_C5698_ = ~new_C5680_ | new_C5690_;
  assign new_C5699_ = new_C5680_ & new_C5690_;
  assign new_C5700_ = ~new_C5680_ & ~new_C5690_;
  assign new_C5701_ = new_C5722_ | new_C5721_;
  assign new_C5702_ = new_C5668_ | new_C5701_;
  assign new_C5703_ = new_C5726_ | new_C5725_;
  assign new_C5704_ = ~new_C5668_ & new_C5703_;
  assign new_C5705_ = new_C5724_ | new_C5723_;
  assign new_C5706_ = new_C5668_ & new_C5705_;
  assign new_C5707_ = new_C5666_ & ~new_C5676_;
  assign new_C5708_ = ~new_C5666_ & new_C5676_;
  assign new_C5709_ = ~new_C5665_ | ~new_C5690_;
  assign new_C5710_ = new_C5676_ & new_C5709_;
  assign new_C5711_ = ~new_C5676_ & ~new_C5710_;
  assign new_C5712_ = new_C5676_ | new_C5709_;
  assign new_C5713_ = ~new_C5666_ & new_C5667_;
  assign new_C5714_ = new_C5666_ & ~new_C5667_;
  assign new_C5715_ = new_C5683_ | new_C5720_;
  assign new_C5716_ = ~new_C5683_ & ~new_C5719_;
  assign new_C5717_ = new_C5666_ | new_C5683_;
  assign new_C5718_ = new_C5666_ | new_C5667_;
  assign new_C5719_ = new_C5683_ & new_C5720_;
  assign new_C5720_ = ~new_C5665_ | ~new_C5690_;
  assign new_C5721_ = new_C5698_ & new_C5718_;
  assign new_C5722_ = ~new_C5698_ & ~new_C5718_;
  assign new_C5723_ = new_C5727_ | new_C5728_;
  assign new_C5724_ = ~new_C5669_ & new_C5683_;
  assign new_C5725_ = new_C5729_ | new_C5730_;
  assign new_C5726_ = new_C5669_ & new_C5683_;
  assign new_C5727_ = ~new_C5669_ & ~new_C5683_;
  assign new_C5728_ = new_C5669_ & ~new_C5683_;
  assign new_C5729_ = new_C5669_ & ~new_C5683_;
  assign new_C5730_ = ~new_C5669_ & new_C5683_;
  assign new_C5731_ = new_E1820_;
  assign new_C5732_ = new_E1887_;
  assign new_C5733_ = new_E1954_;
  assign new_C5734_ = new_E2021_;
  assign new_C5735_ = new_E2088_;
  assign new_C5736_ = new_E2155_;
  assign new_C5737_ = new_C5744_ & new_C5743_;
  assign new_C5738_ = new_C5746_ | new_C5745_;
  assign new_C5739_ = new_C5748_ | new_C5747_;
  assign new_C5740_ = new_C5750_ & new_C5749_;
  assign new_C5741_ = new_C5750_ & new_C5751_;
  assign new_C5742_ = new_C5743_ | new_C5752_;
  assign new_C5743_ = new_C5732_ | new_C5755_;
  assign new_C5744_ = new_C5754_ | new_C5753_;
  assign new_C5745_ = new_C5759_ & new_C5758_;
  assign new_C5746_ = new_C5757_ & new_C5756_;
  assign new_C5747_ = new_C5762_ | new_C5761_;
  assign new_C5748_ = new_C5757_ & new_C5760_;
  assign new_C5749_ = new_C5732_ | new_C5765_;
  assign new_C5750_ = new_C5764_ | new_C5763_;
  assign new_C5751_ = new_C5767_ | new_C5766_;
  assign new_C5752_ = ~new_C5743_ & new_C5769_;
  assign new_C5753_ = ~new_C5745_ & new_C5757_;
  assign new_C5754_ = new_C5745_ & ~new_C5757_;
  assign new_C5755_ = new_C5731_ & ~new_C5732_;
  assign new_C5756_ = ~new_C5778_ | ~new_C5779_;
  assign new_C5757_ = new_C5771_ | new_C5773_;
  assign new_C5758_ = new_C5781_ | new_C5780_;
  assign new_C5759_ = new_C5775_ | new_C5774_;
  assign new_C5760_ = ~new_C5783_ | ~new_C5782_;
  assign new_C5761_ = ~new_C5784_ & new_C5785_;
  assign new_C5762_ = new_C5784_ & ~new_C5785_;
  assign new_C5763_ = ~new_C5731_ & new_C5732_;
  assign new_C5764_ = new_C5731_ & ~new_C5732_;
  assign new_C5765_ = ~new_C5747_ | new_C5757_;
  assign new_C5766_ = new_C5747_ & new_C5757_;
  assign new_C5767_ = ~new_C5747_ & ~new_C5757_;
  assign new_C5768_ = new_C5789_ | new_C5788_;
  assign new_C5769_ = new_C5735_ | new_C5768_;
  assign new_C5770_ = new_C5793_ | new_C5792_;
  assign new_C5771_ = ~new_C5735_ & new_C5770_;
  assign new_C5772_ = new_C5791_ | new_C5790_;
  assign new_C5773_ = new_C5735_ & new_C5772_;
  assign new_C5774_ = new_C5733_ & ~new_C5743_;
  assign new_C5775_ = ~new_C5733_ & new_C5743_;
  assign new_C5776_ = ~new_C5732_ | ~new_C5757_;
  assign new_C5777_ = new_C5743_ & new_C5776_;
  assign new_C5778_ = ~new_C5743_ & ~new_C5777_;
  assign new_C5779_ = new_C5743_ | new_C5776_;
  assign new_C5780_ = ~new_C5733_ & new_C5734_;
  assign new_C5781_ = new_C5733_ & ~new_C5734_;
  assign new_C5782_ = new_C5750_ | new_C5787_;
  assign new_C5783_ = ~new_C5750_ & ~new_C5786_;
  assign new_C5784_ = new_C5733_ | new_C5750_;
  assign new_C5785_ = new_C5733_ | new_C5734_;
  assign new_C5786_ = new_C5750_ & new_C5787_;
  assign new_C5787_ = ~new_C5732_ | ~new_C5757_;
  assign new_C5788_ = new_C5765_ & new_C5785_;
  assign new_C5789_ = ~new_C5765_ & ~new_C5785_;
  assign new_C5790_ = new_C5794_ | new_C5795_;
  assign new_C5791_ = ~new_C5736_ & new_C5750_;
  assign new_C5792_ = new_C5796_ | new_C5797_;
  assign new_C5793_ = new_C5736_ & new_C5750_;
  assign new_C5794_ = ~new_C5736_ & ~new_C5750_;
  assign new_C5795_ = new_C5736_ & ~new_C5750_;
  assign new_C5796_ = new_C5736_ & ~new_C5750_;
  assign new_C5797_ = ~new_C5736_ & new_C5750_;
  assign new_C5798_ = new_E2222_;
  assign new_C5799_ = new_E2289_;
  assign new_C5800_ = new_E2356_;
  assign new_C5801_ = new_E2423_;
  assign new_C5802_ = new_E2490_;
  assign new_C5803_ = new_E2557_;
  assign new_C5804_ = new_C5811_ & new_C5810_;
  assign new_C5805_ = new_C5813_ | new_C5812_;
  assign new_C5806_ = new_C5815_ | new_C5814_;
  assign new_C5807_ = new_C5817_ & new_C5816_;
  assign new_C5808_ = new_C5817_ & new_C5818_;
  assign new_C5809_ = new_C5810_ | new_C5819_;
  assign new_C5810_ = new_C5799_ | new_C5822_;
  assign new_C5811_ = new_C5821_ | new_C5820_;
  assign new_C5812_ = new_C5826_ & new_C5825_;
  assign new_C5813_ = new_C5824_ & new_C5823_;
  assign new_C5814_ = new_C5829_ | new_C5828_;
  assign new_C5815_ = new_C5824_ & new_C5827_;
  assign new_C5816_ = new_C5799_ | new_C5832_;
  assign new_C5817_ = new_C5831_ | new_C5830_;
  assign new_C5818_ = new_C5834_ | new_C5833_;
  assign new_C5819_ = ~new_C5810_ & new_C5836_;
  assign new_C5820_ = ~new_C5812_ & new_C5824_;
  assign new_C5821_ = new_C5812_ & ~new_C5824_;
  assign new_C5822_ = new_C5798_ & ~new_C5799_;
  assign new_C5823_ = ~new_C5845_ | ~new_C5846_;
  assign new_C5824_ = new_C5838_ | new_C5840_;
  assign new_C5825_ = new_C5848_ | new_C5847_;
  assign new_C5826_ = new_C5842_ | new_C5841_;
  assign new_C5827_ = ~new_C5850_ | ~new_C5849_;
  assign new_C5828_ = ~new_C5851_ & new_C5852_;
  assign new_C5829_ = new_C5851_ & ~new_C5852_;
  assign new_C5830_ = ~new_C5798_ & new_C5799_;
  assign new_C5831_ = new_C5798_ & ~new_C5799_;
  assign new_C5832_ = ~new_C5814_ | new_C5824_;
  assign new_C5833_ = new_C5814_ & new_C5824_;
  assign new_C5834_ = ~new_C5814_ & ~new_C5824_;
  assign new_C5835_ = new_C5856_ | new_C5855_;
  assign new_C5836_ = new_C5802_ | new_C5835_;
  assign new_C5837_ = new_C5860_ | new_C5859_;
  assign new_C5838_ = ~new_C5802_ & new_C5837_;
  assign new_C5839_ = new_C5858_ | new_C5857_;
  assign new_C5840_ = new_C5802_ & new_C5839_;
  assign new_C5841_ = new_C5800_ & ~new_C5810_;
  assign new_C5842_ = ~new_C5800_ & new_C5810_;
  assign new_C5843_ = ~new_C5799_ | ~new_C5824_;
  assign new_C5844_ = new_C5810_ & new_C5843_;
  assign new_C5845_ = ~new_C5810_ & ~new_C5844_;
  assign new_C5846_ = new_C5810_ | new_C5843_;
  assign new_C5847_ = ~new_C5800_ & new_C5801_;
  assign new_C5848_ = new_C5800_ & ~new_C5801_;
  assign new_C5849_ = new_C5817_ | new_C5854_;
  assign new_C5850_ = ~new_C5817_ & ~new_C5853_;
  assign new_C5851_ = new_C5800_ | new_C5817_;
  assign new_C5852_ = new_C5800_ | new_C5801_;
  assign new_C5853_ = new_C5817_ & new_C5854_;
  assign new_C5854_ = ~new_C5799_ | ~new_C5824_;
  assign new_C5855_ = new_C5832_ & new_C5852_;
  assign new_C5856_ = ~new_C5832_ & ~new_C5852_;
  assign new_C5857_ = new_C5861_ | new_C5862_;
  assign new_C5858_ = ~new_C5803_ & new_C5817_;
  assign new_C5859_ = new_C5863_ | new_C5864_;
  assign new_C5860_ = new_C5803_ & new_C5817_;
  assign new_C5861_ = ~new_C5803_ & ~new_C5817_;
  assign new_C5862_ = new_C5803_ & ~new_C5817_;
  assign new_C5863_ = new_C5803_ & ~new_C5817_;
  assign new_C5864_ = ~new_C5803_ & new_C5817_;
  assign new_C5865_ = new_E2624_;
  assign new_C5866_ = new_E2691_;
  assign new_C5867_ = new_E2758_;
  assign new_C5868_ = new_E2825_;
  assign new_C5869_ = new_E2892_;
  assign new_C5870_ = new_E2959_;
  assign new_C5871_ = new_C5878_ & new_C5877_;
  assign new_C5872_ = new_C5880_ | new_C5879_;
  assign new_C5873_ = new_C5882_ | new_C5881_;
  assign new_C5874_ = new_C5884_ & new_C5883_;
  assign new_C5875_ = new_C5884_ & new_C5885_;
  assign new_C5876_ = new_C5877_ | new_C5886_;
  assign new_C5877_ = new_C5866_ | new_C5889_;
  assign new_C5878_ = new_C5888_ | new_C5887_;
  assign new_C5879_ = new_C5893_ & new_C5892_;
  assign new_C5880_ = new_C5891_ & new_C5890_;
  assign new_C5881_ = new_C5896_ | new_C5895_;
  assign new_C5882_ = new_C5891_ & new_C5894_;
  assign new_C5883_ = new_C5866_ | new_C5899_;
  assign new_C5884_ = new_C5898_ | new_C5897_;
  assign new_C5885_ = new_C5901_ | new_C5900_;
  assign new_C5886_ = ~new_C5877_ & new_C5903_;
  assign new_C5887_ = ~new_C5879_ & new_C5891_;
  assign new_C5888_ = new_C5879_ & ~new_C5891_;
  assign new_C5889_ = new_C5865_ & ~new_C5866_;
  assign new_C5890_ = ~new_C5912_ | ~new_C5913_;
  assign new_C5891_ = new_C5905_ | new_C5907_;
  assign new_C5892_ = new_C5915_ | new_C5914_;
  assign new_C5893_ = new_C5909_ | new_C5908_;
  assign new_C5894_ = ~new_C5917_ | ~new_C5916_;
  assign new_C5895_ = ~new_C5918_ & new_C5919_;
  assign new_C5896_ = new_C5918_ & ~new_C5919_;
  assign new_C5897_ = ~new_C5865_ & new_C5866_;
  assign new_C5898_ = new_C5865_ & ~new_C5866_;
  assign new_C5899_ = ~new_C5881_ | new_C5891_;
  assign new_C5900_ = new_C5881_ & new_C5891_;
  assign new_C5901_ = ~new_C5881_ & ~new_C5891_;
  assign new_C5902_ = new_C5923_ | new_C5922_;
  assign new_C5903_ = new_C5869_ | new_C5902_;
  assign new_C5904_ = new_C5927_ | new_C5926_;
  assign new_C5905_ = ~new_C5869_ & new_C5904_;
  assign new_C5906_ = new_C5925_ | new_C5924_;
  assign new_C5907_ = new_C5869_ & new_C5906_;
  assign new_C5908_ = new_C5867_ & ~new_C5877_;
  assign new_C5909_ = ~new_C5867_ & new_C5877_;
  assign new_C5910_ = ~new_C5866_ | ~new_C5891_;
  assign new_C5911_ = new_C5877_ & new_C5910_;
  assign new_C5912_ = ~new_C5877_ & ~new_C5911_;
  assign new_C5913_ = new_C5877_ | new_C5910_;
  assign new_C5914_ = ~new_C5867_ & new_C5868_;
  assign new_C5915_ = new_C5867_ & ~new_C5868_;
  assign new_C5916_ = new_C5884_ | new_C5921_;
  assign new_C5917_ = ~new_C5884_ & ~new_C5920_;
  assign new_C5918_ = new_C5867_ | new_C5884_;
  assign new_C5919_ = new_C5867_ | new_C5868_;
  assign new_C5920_ = new_C5884_ & new_C5921_;
  assign new_C5921_ = ~new_C5866_ | ~new_C5891_;
  assign new_C5922_ = new_C5899_ & new_C5919_;
  assign new_C5923_ = ~new_C5899_ & ~new_C5919_;
  assign new_C5924_ = new_C5928_ | new_C5929_;
  assign new_C5925_ = ~new_C5870_ & new_C5884_;
  assign new_C5926_ = new_C5930_ | new_C5931_;
  assign new_C5927_ = new_C5870_ & new_C5884_;
  assign new_C5928_ = ~new_C5870_ & ~new_C5884_;
  assign new_C5929_ = new_C5870_ & ~new_C5884_;
  assign new_C5930_ = new_C5870_ & ~new_C5884_;
  assign new_C5931_ = ~new_C5870_ & new_C5884_;
  assign new_C5932_ = new_E3026_;
  assign new_C5933_ = new_E3093_;
  assign new_C5934_ = new_E3160_;
  assign new_C5935_ = new_E3227_;
  assign new_C5936_ = new_E3294_;
  assign new_C5937_ = new_E3361_;
  assign new_C5938_ = new_C5945_ & new_C5944_;
  assign new_C5939_ = new_C5947_ | new_C5946_;
  assign new_C5940_ = new_C5949_ | new_C5948_;
  assign new_C5941_ = new_C5951_ & new_C5950_;
  assign new_C5942_ = new_C5951_ & new_C5952_;
  assign new_C5943_ = new_C5944_ | new_C5953_;
  assign new_C5944_ = new_C5933_ | new_C5956_;
  assign new_C5945_ = new_C5955_ | new_C5954_;
  assign new_C5946_ = new_C5960_ & new_C5959_;
  assign new_C5947_ = new_C5958_ & new_C5957_;
  assign new_C5948_ = new_C5963_ | new_C5962_;
  assign new_C5949_ = new_C5958_ & new_C5961_;
  assign new_C5950_ = new_C5933_ | new_C5966_;
  assign new_C5951_ = new_C5965_ | new_C5964_;
  assign new_C5952_ = new_C5968_ | new_C5967_;
  assign new_C5953_ = ~new_C5944_ & new_C5970_;
  assign new_C5954_ = ~new_C5946_ & new_C5958_;
  assign new_C5955_ = new_C5946_ & ~new_C5958_;
  assign new_C5956_ = new_C5932_ & ~new_C5933_;
  assign new_C5957_ = ~new_C5979_ | ~new_C5980_;
  assign new_C5958_ = new_C5972_ | new_C5974_;
  assign new_C5959_ = new_C5982_ | new_C5981_;
  assign new_C5960_ = new_C5976_ | new_C5975_;
  assign new_C5961_ = ~new_C5984_ | ~new_C5983_;
  assign new_C5962_ = ~new_C5985_ & new_C5986_;
  assign new_C5963_ = new_C5985_ & ~new_C5986_;
  assign new_C5964_ = ~new_C5932_ & new_C5933_;
  assign new_C5965_ = new_C5932_ & ~new_C5933_;
  assign new_C5966_ = ~new_C5948_ | new_C5958_;
  assign new_C5967_ = new_C5948_ & new_C5958_;
  assign new_C5968_ = ~new_C5948_ & ~new_C5958_;
  assign new_C5969_ = new_C5990_ | new_C5989_;
  assign new_C5970_ = new_C5936_ | new_C5969_;
  assign new_C5971_ = new_C5994_ | new_C5993_;
  assign new_C5972_ = ~new_C5936_ & new_C5971_;
  assign new_C5973_ = new_C5992_ | new_C5991_;
  assign new_C5974_ = new_C5936_ & new_C5973_;
  assign new_C5975_ = new_C5934_ & ~new_C5944_;
  assign new_C5976_ = ~new_C5934_ & new_C5944_;
  assign new_C5977_ = ~new_C5933_ | ~new_C5958_;
  assign new_C5978_ = new_C5944_ & new_C5977_;
  assign new_C5979_ = ~new_C5944_ & ~new_C5978_;
  assign new_C5980_ = new_C5944_ | new_C5977_;
  assign new_C5981_ = ~new_C5934_ & new_C5935_;
  assign new_C5982_ = new_C5934_ & ~new_C5935_;
  assign new_C5983_ = new_C5951_ | new_C5988_;
  assign new_C5984_ = ~new_C5951_ & ~new_C5987_;
  assign new_C5985_ = new_C5934_ | new_C5951_;
  assign new_C5986_ = new_C5934_ | new_C5935_;
  assign new_C5987_ = new_C5951_ & new_C5988_;
  assign new_C5988_ = ~new_C5933_ | ~new_C5958_;
  assign new_C5989_ = new_C5966_ & new_C5986_;
  assign new_C5990_ = ~new_C5966_ & ~new_C5986_;
  assign new_C5991_ = new_C5995_ | new_C5996_;
  assign new_C5992_ = ~new_C5937_ & new_C5951_;
  assign new_C5993_ = new_C5997_ | new_C5998_;
  assign new_C5994_ = new_C5937_ & new_C5951_;
  assign new_C5995_ = ~new_C5937_ & ~new_C5951_;
  assign new_C5996_ = new_C5937_ & ~new_C5951_;
  assign new_C5997_ = new_C5937_ & ~new_C5951_;
  assign new_C5998_ = ~new_C5937_ & new_C5951_;
  assign new_C5999_ = new_E3428_;
  assign new_C6000_ = new_E3495_;
  assign new_C6001_ = new_E3562_;
  assign new_C6002_ = new_E3629_;
  assign new_C6003_ = new_E3696_;
  assign new_C6004_ = new_E3763_;
  assign new_C6005_ = new_C6012_ & new_C6011_;
  assign new_C6006_ = new_C6014_ | new_C6013_;
  assign new_C6007_ = new_C6016_ | new_C6015_;
  assign new_C6008_ = new_C6018_ & new_C6017_;
  assign new_C6009_ = new_C6018_ & new_C6019_;
  assign new_C6010_ = new_C6011_ | new_C6020_;
  assign new_C6011_ = new_C6000_ | new_C6023_;
  assign new_C6012_ = new_C6022_ | new_C6021_;
  assign new_C6013_ = new_C6027_ & new_C6026_;
  assign new_C6014_ = new_C6025_ & new_C6024_;
  assign new_C6015_ = new_C6030_ | new_C6029_;
  assign new_C6016_ = new_C6025_ & new_C6028_;
  assign new_C6017_ = new_C6000_ | new_C6033_;
  assign new_C6018_ = new_C6032_ | new_C6031_;
  assign new_C6019_ = new_C6035_ | new_C6034_;
  assign new_C6020_ = ~new_C6011_ & new_C6037_;
  assign new_C6021_ = ~new_C6013_ & new_C6025_;
  assign new_C6022_ = new_C6013_ & ~new_C6025_;
  assign new_C6023_ = new_C5999_ & ~new_C6000_;
  assign new_C6024_ = ~new_C6046_ | ~new_C6047_;
  assign new_C6025_ = new_C6039_ | new_C6041_;
  assign new_C6026_ = new_C6049_ | new_C6048_;
  assign new_C6027_ = new_C6043_ | new_C6042_;
  assign new_C6028_ = ~new_C6051_ | ~new_C6050_;
  assign new_C6029_ = ~new_C6052_ & new_C6053_;
  assign new_C6030_ = new_C6052_ & ~new_C6053_;
  assign new_C6031_ = ~new_C5999_ & new_C6000_;
  assign new_C6032_ = new_C5999_ & ~new_C6000_;
  assign new_C6033_ = ~new_C6015_ | new_C6025_;
  assign new_C6034_ = new_C6015_ & new_C6025_;
  assign new_C6035_ = ~new_C6015_ & ~new_C6025_;
  assign new_C6036_ = new_C6057_ | new_C6056_;
  assign new_C6037_ = new_C6003_ | new_C6036_;
  assign new_C6038_ = new_C6061_ | new_C6060_;
  assign new_C6039_ = ~new_C6003_ & new_C6038_;
  assign new_C6040_ = new_C6059_ | new_C6058_;
  assign new_C6041_ = new_C6003_ & new_C6040_;
  assign new_C6042_ = new_C6001_ & ~new_C6011_;
  assign new_C6043_ = ~new_C6001_ & new_C6011_;
  assign new_C6044_ = ~new_C6000_ | ~new_C6025_;
  assign new_C6045_ = new_C6011_ & new_C6044_;
  assign new_C6046_ = ~new_C6011_ & ~new_C6045_;
  assign new_C6047_ = new_C6011_ | new_C6044_;
  assign new_C6048_ = ~new_C6001_ & new_C6002_;
  assign new_C6049_ = new_C6001_ & ~new_C6002_;
  assign new_C6050_ = new_C6018_ | new_C6055_;
  assign new_C6051_ = ~new_C6018_ & ~new_C6054_;
  assign new_C6052_ = new_C6001_ | new_C6018_;
  assign new_C6053_ = new_C6001_ | new_C6002_;
  assign new_C6054_ = new_C6018_ & new_C6055_;
  assign new_C6055_ = ~new_C6000_ | ~new_C6025_;
  assign new_C6056_ = new_C6033_ & new_C6053_;
  assign new_C6057_ = ~new_C6033_ & ~new_C6053_;
  assign new_C6058_ = new_C6062_ | new_C6063_;
  assign new_C6059_ = ~new_C6004_ & new_C6018_;
  assign new_C6060_ = new_C6064_ | new_C6065_;
  assign new_C6061_ = new_C6004_ & new_C6018_;
  assign new_C6062_ = ~new_C6004_ & ~new_C6018_;
  assign new_C6063_ = new_C6004_ & ~new_C6018_;
  assign new_C6064_ = new_C6004_ & ~new_C6018_;
  assign new_C6065_ = ~new_C6004_ & new_C6018_;
  assign new_C6066_ = new_E3830_;
  assign new_C6067_ = new_E3897_;
  assign new_C6068_ = new_E3964_;
  assign new_C6069_ = new_E4031_;
  assign new_C6070_ = new_E4098_;
  assign new_C6071_ = new_E4165_;
  assign new_C6072_ = new_C6079_ & new_C6078_;
  assign new_C6073_ = new_C6081_ | new_C6080_;
  assign new_C6074_ = new_C6083_ | new_C6082_;
  assign new_C6075_ = new_C6085_ & new_C6084_;
  assign new_C6076_ = new_C6085_ & new_C6086_;
  assign new_C6077_ = new_C6078_ | new_C6087_;
  assign new_C6078_ = new_C6067_ | new_C6090_;
  assign new_C6079_ = new_C6089_ | new_C6088_;
  assign new_C6080_ = new_C6094_ & new_C6093_;
  assign new_C6081_ = new_C6092_ & new_C6091_;
  assign new_C6082_ = new_C6097_ | new_C6096_;
  assign new_C6083_ = new_C6092_ & new_C6095_;
  assign new_C6084_ = new_C6067_ | new_C6100_;
  assign new_C6085_ = new_C6099_ | new_C6098_;
  assign new_C6086_ = new_C6102_ | new_C6101_;
  assign new_C6087_ = ~new_C6078_ & new_C6104_;
  assign new_C6088_ = ~new_C6080_ & new_C6092_;
  assign new_C6089_ = new_C6080_ & ~new_C6092_;
  assign new_C6090_ = new_C6066_ & ~new_C6067_;
  assign new_C6091_ = ~new_C6113_ | ~new_C6114_;
  assign new_C6092_ = new_C6106_ | new_C6108_;
  assign new_C6093_ = new_C6116_ | new_C6115_;
  assign new_C6094_ = new_C6110_ | new_C6109_;
  assign new_C6095_ = ~new_C6118_ | ~new_C6117_;
  assign new_C6096_ = ~new_C6119_ & new_C6120_;
  assign new_C6097_ = new_C6119_ & ~new_C6120_;
  assign new_C6098_ = ~new_C6066_ & new_C6067_;
  assign new_C6099_ = new_C6066_ & ~new_C6067_;
  assign new_C6100_ = ~new_C6082_ | new_C6092_;
  assign new_C6101_ = new_C6082_ & new_C6092_;
  assign new_C6102_ = ~new_C6082_ & ~new_C6092_;
  assign new_C6103_ = new_C6124_ | new_C6123_;
  assign new_C6104_ = new_C6070_ | new_C6103_;
  assign new_C6105_ = new_C6128_ | new_C6127_;
  assign new_C6106_ = ~new_C6070_ & new_C6105_;
  assign new_C6107_ = new_C6126_ | new_C6125_;
  assign new_C6108_ = new_C6070_ & new_C6107_;
  assign new_C6109_ = new_C6068_ & ~new_C6078_;
  assign new_C6110_ = ~new_C6068_ & new_C6078_;
  assign new_C6111_ = ~new_C6067_ | ~new_C6092_;
  assign new_C6112_ = new_C6078_ & new_C6111_;
  assign new_C6113_ = ~new_C6078_ & ~new_C6112_;
  assign new_C6114_ = new_C6078_ | new_C6111_;
  assign new_C6115_ = ~new_C6068_ & new_C6069_;
  assign new_C6116_ = new_C6068_ & ~new_C6069_;
  assign new_C6117_ = new_C6085_ | new_C6122_;
  assign new_C6118_ = ~new_C6085_ & ~new_C6121_;
  assign new_C6119_ = new_C6068_ | new_C6085_;
  assign new_C6120_ = new_C6068_ | new_C6069_;
  assign new_C6121_ = new_C6085_ & new_C6122_;
  assign new_C6122_ = ~new_C6067_ | ~new_C6092_;
  assign new_C6123_ = new_C6100_ & new_C6120_;
  assign new_C6124_ = ~new_C6100_ & ~new_C6120_;
  assign new_C6125_ = new_C6129_ | new_C6130_;
  assign new_C6126_ = ~new_C6071_ & new_C6085_;
  assign new_C6127_ = new_C6131_ | new_C6132_;
  assign new_C6128_ = new_C6071_ & new_C6085_;
  assign new_C6129_ = ~new_C6071_ & ~new_C6085_;
  assign new_C6130_ = new_C6071_ & ~new_C6085_;
  assign new_C6131_ = new_C6071_ & ~new_C6085_;
  assign new_C6132_ = ~new_C6071_ & new_C6085_;
  assign new_C6133_ = new_E4232_;
  assign new_C6134_ = new_E4299_;
  assign new_C6135_ = new_E4366_;
  assign new_C6136_ = new_E4433_;
  assign new_C6137_ = new_E4500_;
  assign new_C6138_ = new_E4567_;
  assign new_C6139_ = new_C6146_ & new_C6145_;
  assign new_C6140_ = new_C6148_ | new_C6147_;
  assign new_C6141_ = new_C6150_ | new_C6149_;
  assign new_C6142_ = new_C6152_ & new_C6151_;
  assign new_C6143_ = new_C6152_ & new_C6153_;
  assign new_C6144_ = new_C6145_ | new_C6154_;
  assign new_C6145_ = new_C6134_ | new_C6157_;
  assign new_C6146_ = new_C6156_ | new_C6155_;
  assign new_C6147_ = new_C6161_ & new_C6160_;
  assign new_C6148_ = new_C6159_ & new_C6158_;
  assign new_C6149_ = new_C6164_ | new_C6163_;
  assign new_C6150_ = new_C6159_ & new_C6162_;
  assign new_C6151_ = new_C6134_ | new_C6167_;
  assign new_C6152_ = new_C6166_ | new_C6165_;
  assign new_C6153_ = new_C6169_ | new_C6168_;
  assign new_C6154_ = ~new_C6145_ & new_C6171_;
  assign new_C6155_ = ~new_C6147_ & new_C6159_;
  assign new_C6156_ = new_C6147_ & ~new_C6159_;
  assign new_C6157_ = new_C6133_ & ~new_C6134_;
  assign new_C6158_ = ~new_C6180_ | ~new_C6181_;
  assign new_C6159_ = new_C6173_ | new_C6175_;
  assign new_C6160_ = new_C6183_ | new_C6182_;
  assign new_C6161_ = new_C6177_ | new_C6176_;
  assign new_C6162_ = ~new_C6185_ | ~new_C6184_;
  assign new_C6163_ = ~new_C6186_ & new_C6187_;
  assign new_C6164_ = new_C6186_ & ~new_C6187_;
  assign new_C6165_ = ~new_C6133_ & new_C6134_;
  assign new_C6166_ = new_C6133_ & ~new_C6134_;
  assign new_C6167_ = ~new_C6149_ | new_C6159_;
  assign new_C6168_ = new_C6149_ & new_C6159_;
  assign new_C6169_ = ~new_C6149_ & ~new_C6159_;
  assign new_C6170_ = new_C6191_ | new_C6190_;
  assign new_C6171_ = new_C6137_ | new_C6170_;
  assign new_C6172_ = new_C6195_ | new_C6194_;
  assign new_C6173_ = ~new_C6137_ & new_C6172_;
  assign new_C6174_ = new_C6193_ | new_C6192_;
  assign new_C6175_ = new_C6137_ & new_C6174_;
  assign new_C6176_ = new_C6135_ & ~new_C6145_;
  assign new_C6177_ = ~new_C6135_ & new_C6145_;
  assign new_C6178_ = ~new_C6134_ | ~new_C6159_;
  assign new_C6179_ = new_C6145_ & new_C6178_;
  assign new_C6180_ = ~new_C6145_ & ~new_C6179_;
  assign new_C6181_ = new_C6145_ | new_C6178_;
  assign new_C6182_ = ~new_C6135_ & new_C6136_;
  assign new_C6183_ = new_C6135_ & ~new_C6136_;
  assign new_C6184_ = new_C6152_ | new_C6189_;
  assign new_C6185_ = ~new_C6152_ & ~new_C6188_;
  assign new_C6186_ = new_C6135_ | new_C6152_;
  assign new_C6187_ = new_C6135_ | new_C6136_;
  assign new_C6188_ = new_C6152_ & new_C6189_;
  assign new_C6189_ = ~new_C6134_ | ~new_C6159_;
  assign new_C6190_ = new_C6167_ & new_C6187_;
  assign new_C6191_ = ~new_C6167_ & ~new_C6187_;
  assign new_C6192_ = new_C6196_ | new_C6197_;
  assign new_C6193_ = ~new_C6138_ & new_C6152_;
  assign new_C6194_ = new_C6198_ | new_C6199_;
  assign new_C6195_ = new_C6138_ & new_C6152_;
  assign new_C6196_ = ~new_C6138_ & ~new_C6152_;
  assign new_C6197_ = new_C6138_ & ~new_C6152_;
  assign new_C6198_ = new_C6138_ & ~new_C6152_;
  assign new_C6199_ = ~new_C6138_ & new_C6152_;
  assign new_C6200_ = new_E4634_;
  assign new_C6201_ = new_E4701_;
  assign new_C6202_ = new_E4768_;
  assign new_C6203_ = new_E4835_;
  assign new_C6204_ = new_E4902_;
  assign new_C6205_ = new_E4969_;
  assign new_C6206_ = new_C6213_ & new_C6212_;
  assign new_C6207_ = new_C6215_ | new_C6214_;
  assign new_C6208_ = new_C6217_ | new_C6216_;
  assign new_C6209_ = new_C6219_ & new_C6218_;
  assign new_C6210_ = new_C6219_ & new_C6220_;
  assign new_C6211_ = new_C6212_ | new_C6221_;
  assign new_C6212_ = new_C6201_ | new_C6224_;
  assign new_C6213_ = new_C6223_ | new_C6222_;
  assign new_C6214_ = new_C6228_ & new_C6227_;
  assign new_C6215_ = new_C6226_ & new_C6225_;
  assign new_C6216_ = new_C6231_ | new_C6230_;
  assign new_C6217_ = new_C6226_ & new_C6229_;
  assign new_C6218_ = new_C6201_ | new_C6234_;
  assign new_C6219_ = new_C6233_ | new_C6232_;
  assign new_C6220_ = new_C6236_ | new_C6235_;
  assign new_C6221_ = ~new_C6212_ & new_C6238_;
  assign new_C6222_ = ~new_C6214_ & new_C6226_;
  assign new_C6223_ = new_C6214_ & ~new_C6226_;
  assign new_C6224_ = new_C6200_ & ~new_C6201_;
  assign new_C6225_ = ~new_C6247_ | ~new_C6248_;
  assign new_C6226_ = new_C6240_ | new_C6242_;
  assign new_C6227_ = new_C6250_ | new_C6249_;
  assign new_C6228_ = new_C6244_ | new_C6243_;
  assign new_C6229_ = ~new_C6252_ | ~new_C6251_;
  assign new_C6230_ = ~new_C6253_ & new_C6254_;
  assign new_C6231_ = new_C6253_ & ~new_C6254_;
  assign new_C6232_ = ~new_C6200_ & new_C6201_;
  assign new_C6233_ = new_C6200_ & ~new_C6201_;
  assign new_C6234_ = ~new_C6216_ | new_C6226_;
  assign new_C6235_ = new_C6216_ & new_C6226_;
  assign new_C6236_ = ~new_C6216_ & ~new_C6226_;
  assign new_C6237_ = new_C6258_ | new_C6257_;
  assign new_C6238_ = new_C6204_ | new_C6237_;
  assign new_C6239_ = new_C6262_ | new_C6261_;
  assign new_C6240_ = ~new_C6204_ & new_C6239_;
  assign new_C6241_ = new_C6260_ | new_C6259_;
  assign new_C6242_ = new_C6204_ & new_C6241_;
  assign new_C6243_ = new_C6202_ & ~new_C6212_;
  assign new_C6244_ = ~new_C6202_ & new_C6212_;
  assign new_C6245_ = ~new_C6201_ | ~new_C6226_;
  assign new_C6246_ = new_C6212_ & new_C6245_;
  assign new_C6247_ = ~new_C6212_ & ~new_C6246_;
  assign new_C6248_ = new_C6212_ | new_C6245_;
  assign new_C6249_ = ~new_C6202_ & new_C6203_;
  assign new_C6250_ = new_C6202_ & ~new_C6203_;
  assign new_C6251_ = new_C6219_ | new_C6256_;
  assign new_C6252_ = ~new_C6219_ & ~new_C6255_;
  assign new_C6253_ = new_C6202_ | new_C6219_;
  assign new_C6254_ = new_C6202_ | new_C6203_;
  assign new_C6255_ = new_C6219_ & new_C6256_;
  assign new_C6256_ = ~new_C6201_ | ~new_C6226_;
  assign new_C6257_ = new_C6234_ & new_C6254_;
  assign new_C6258_ = ~new_C6234_ & ~new_C6254_;
  assign new_C6259_ = new_C6263_ | new_C6264_;
  assign new_C6260_ = ~new_C6205_ & new_C6219_;
  assign new_C6261_ = new_C6265_ | new_C6266_;
  assign new_C6262_ = new_C6205_ & new_C6219_;
  assign new_C6263_ = ~new_C6205_ & ~new_C6219_;
  assign new_C6264_ = new_C6205_ & ~new_C6219_;
  assign new_C6265_ = new_C6205_ & ~new_C6219_;
  assign new_C6266_ = ~new_C6205_ & new_C6219_;
  assign new_C6267_ = new_E5036_;
  assign new_C6268_ = new_E5103_;
  assign new_C6269_ = new_E5170_;
  assign new_C6270_ = new_E5237_;
  assign new_C6271_ = new_E5304_;
  assign new_C6272_ = new_E5371_;
  assign new_C6273_ = new_C6280_ & new_C6279_;
  assign new_C6274_ = new_C6282_ | new_C6281_;
  assign new_C6275_ = new_C6284_ | new_C6283_;
  assign new_C6276_ = new_C6286_ & new_C6285_;
  assign new_C6277_ = new_C6286_ & new_C6287_;
  assign new_C6278_ = new_C6279_ | new_C6288_;
  assign new_C6279_ = new_C6268_ | new_C6291_;
  assign new_C6280_ = new_C6290_ | new_C6289_;
  assign new_C6281_ = new_C6295_ & new_C6294_;
  assign new_C6282_ = new_C6293_ & new_C6292_;
  assign new_C6283_ = new_C6298_ | new_C6297_;
  assign new_C6284_ = new_C6293_ & new_C6296_;
  assign new_C6285_ = new_C6268_ | new_C6301_;
  assign new_C6286_ = new_C6300_ | new_C6299_;
  assign new_C6287_ = new_C6303_ | new_C6302_;
  assign new_C6288_ = ~new_C6279_ & new_C6305_;
  assign new_C6289_ = ~new_C6281_ & new_C6293_;
  assign new_C6290_ = new_C6281_ & ~new_C6293_;
  assign new_C6291_ = new_C6267_ & ~new_C6268_;
  assign new_C6292_ = ~new_C6314_ | ~new_C6315_;
  assign new_C6293_ = new_C6307_ | new_C6309_;
  assign new_C6294_ = new_C6317_ | new_C6316_;
  assign new_C6295_ = new_C6311_ | new_C6310_;
  assign new_C6296_ = ~new_C6319_ | ~new_C6318_;
  assign new_C6297_ = ~new_C6320_ & new_C6321_;
  assign new_C6298_ = new_C6320_ & ~new_C6321_;
  assign new_C6299_ = ~new_C6267_ & new_C6268_;
  assign new_C6300_ = new_C6267_ & ~new_C6268_;
  assign new_C6301_ = ~new_C6283_ | new_C6293_;
  assign new_C6302_ = new_C6283_ & new_C6293_;
  assign new_C6303_ = ~new_C6283_ & ~new_C6293_;
  assign new_C6304_ = new_C6325_ | new_C6324_;
  assign new_C6305_ = new_C6271_ | new_C6304_;
  assign new_C6306_ = new_C6329_ | new_C6328_;
  assign new_C6307_ = ~new_C6271_ & new_C6306_;
  assign new_C6308_ = new_C6327_ | new_C6326_;
  assign new_C6309_ = new_C6271_ & new_C6308_;
  assign new_C6310_ = new_C6269_ & ~new_C6279_;
  assign new_C6311_ = ~new_C6269_ & new_C6279_;
  assign new_C6312_ = ~new_C6268_ | ~new_C6293_;
  assign new_C6313_ = new_C6279_ & new_C6312_;
  assign new_C6314_ = ~new_C6279_ & ~new_C6313_;
  assign new_C6315_ = new_C6279_ | new_C6312_;
  assign new_C6316_ = ~new_C6269_ & new_C6270_;
  assign new_C6317_ = new_C6269_ & ~new_C6270_;
  assign new_C6318_ = new_C6286_ | new_C6323_;
  assign new_C6319_ = ~new_C6286_ & ~new_C6322_;
  assign new_C6320_ = new_C6269_ | new_C6286_;
  assign new_C6321_ = new_C6269_ | new_C6270_;
  assign new_C6322_ = new_C6286_ & new_C6323_;
  assign new_C6323_ = ~new_C6268_ | ~new_C6293_;
  assign new_C6324_ = new_C6301_ & new_C6321_;
  assign new_C6325_ = ~new_C6301_ & ~new_C6321_;
  assign new_C6326_ = new_C6330_ | new_C6331_;
  assign new_C6327_ = ~new_C6272_ & new_C6286_;
  assign new_C6328_ = new_C6332_ | new_C6333_;
  assign new_C6329_ = new_C6272_ & new_C6286_;
  assign new_C6330_ = ~new_C6272_ & ~new_C6286_;
  assign new_C6331_ = new_C6272_ & ~new_C6286_;
  assign new_C6332_ = new_C6272_ & ~new_C6286_;
  assign new_C6333_ = ~new_C6272_ & new_C6286_;
  assign new_C6334_ = new_E5438_;
  assign new_C6335_ = new_E5505_;
  assign new_C6336_ = new_E5572_;
  assign new_C6337_ = new_E5639_;
  assign new_C6338_ = new_E5706_;
  assign new_C6339_ = new_E5773_;
  assign new_C6340_ = new_C6347_ & new_C6346_;
  assign new_C6341_ = new_C6349_ | new_C6348_;
  assign new_C6342_ = new_C6351_ | new_C6350_;
  assign new_C6343_ = new_C6353_ & new_C6352_;
  assign new_C6344_ = new_C6353_ & new_C6354_;
  assign new_C6345_ = new_C6346_ | new_C6355_;
  assign new_C6346_ = new_C6335_ | new_C6358_;
  assign new_C6347_ = new_C6357_ | new_C6356_;
  assign new_C6348_ = new_C6362_ & new_C6361_;
  assign new_C6349_ = new_C6360_ & new_C6359_;
  assign new_C6350_ = new_C6365_ | new_C6364_;
  assign new_C6351_ = new_C6360_ & new_C6363_;
  assign new_C6352_ = new_C6335_ | new_C6368_;
  assign new_C6353_ = new_C6367_ | new_C6366_;
  assign new_C6354_ = new_C6370_ | new_C6369_;
  assign new_C6355_ = ~new_C6346_ & new_C6372_;
  assign new_C6356_ = ~new_C6348_ & new_C6360_;
  assign new_C6357_ = new_C6348_ & ~new_C6360_;
  assign new_C6358_ = new_C6334_ & ~new_C6335_;
  assign new_C6359_ = ~new_C6381_ | ~new_C6382_;
  assign new_C6360_ = new_C6374_ | new_C6376_;
  assign new_C6361_ = new_C6384_ | new_C6383_;
  assign new_C6362_ = new_C6378_ | new_C6377_;
  assign new_C6363_ = ~new_C6386_ | ~new_C6385_;
  assign new_C6364_ = ~new_C6387_ & new_C6388_;
  assign new_C6365_ = new_C6387_ & ~new_C6388_;
  assign new_C6366_ = ~new_C6334_ & new_C6335_;
  assign new_C6367_ = new_C6334_ & ~new_C6335_;
  assign new_C6368_ = ~new_C6350_ | new_C6360_;
  assign new_C6369_ = new_C6350_ & new_C6360_;
  assign new_C6370_ = ~new_C6350_ & ~new_C6360_;
  assign new_C6371_ = new_C6392_ | new_C6391_;
  assign new_C6372_ = new_C6338_ | new_C6371_;
  assign new_C6373_ = new_C6396_ | new_C6395_;
  assign new_C6374_ = ~new_C6338_ & new_C6373_;
  assign new_C6375_ = new_C6394_ | new_C6393_;
  assign new_C6376_ = new_C6338_ & new_C6375_;
  assign new_C6377_ = new_C6336_ & ~new_C6346_;
  assign new_C6378_ = ~new_C6336_ & new_C6346_;
  assign new_C6379_ = ~new_C6335_ | ~new_C6360_;
  assign new_C6380_ = new_C6346_ & new_C6379_;
  assign new_C6381_ = ~new_C6346_ & ~new_C6380_;
  assign new_C6382_ = new_C6346_ | new_C6379_;
  assign new_C6383_ = ~new_C6336_ & new_C6337_;
  assign new_C6384_ = new_C6336_ & ~new_C6337_;
  assign new_C6385_ = new_C6353_ | new_C6390_;
  assign new_C6386_ = ~new_C6353_ & ~new_C6389_;
  assign new_C6387_ = new_C6336_ | new_C6353_;
  assign new_C6388_ = new_C6336_ | new_C6337_;
  assign new_C6389_ = new_C6353_ & new_C6390_;
  assign new_C6390_ = ~new_C6335_ | ~new_C6360_;
  assign new_C6391_ = new_C6368_ & new_C6388_;
  assign new_C6392_ = ~new_C6368_ & ~new_C6388_;
  assign new_C6393_ = new_C6397_ | new_C6398_;
  assign new_C6394_ = ~new_C6339_ & new_C6353_;
  assign new_C6395_ = new_C6399_ | new_C6400_;
  assign new_C6396_ = new_C6339_ & new_C6353_;
  assign new_C6397_ = ~new_C6339_ & ~new_C6353_;
  assign new_C6398_ = new_C6339_ & ~new_C6353_;
  assign new_C6399_ = new_C6339_ & ~new_C6353_;
  assign new_C6400_ = ~new_C6339_ & new_C6353_;
  assign new_C6401_ = new_E5840_;
  assign new_C6402_ = new_E5907_;
  assign new_C6403_ = new_E5974_;
  assign new_C6404_ = new_E6041_;
  assign new_C6405_ = new_E6108_;
  assign new_C6406_ = new_E6175_;
  assign new_C6407_ = new_C6414_ & new_C6413_;
  assign new_C6408_ = new_C6416_ | new_C6415_;
  assign new_C6409_ = new_C6418_ | new_C6417_;
  assign new_C6410_ = new_C6420_ & new_C6419_;
  assign new_C6411_ = new_C6420_ & new_C6421_;
  assign new_C6412_ = new_C6413_ | new_C6422_;
  assign new_C6413_ = new_C6402_ | new_C6425_;
  assign new_C6414_ = new_C6424_ | new_C6423_;
  assign new_C6415_ = new_C6429_ & new_C6428_;
  assign new_C6416_ = new_C6427_ & new_C6426_;
  assign new_C6417_ = new_C6432_ | new_C6431_;
  assign new_C6418_ = new_C6427_ & new_C6430_;
  assign new_C6419_ = new_C6402_ | new_C6435_;
  assign new_C6420_ = new_C6434_ | new_C6433_;
  assign new_C6421_ = new_C6437_ | new_C6436_;
  assign new_C6422_ = ~new_C6413_ & new_C6439_;
  assign new_C6423_ = ~new_C6415_ & new_C6427_;
  assign new_C6424_ = new_C6415_ & ~new_C6427_;
  assign new_C6425_ = new_C6401_ & ~new_C6402_;
  assign new_C6426_ = ~new_C6448_ | ~new_C6449_;
  assign new_C6427_ = new_C6441_ | new_C6443_;
  assign new_C6428_ = new_C6451_ | new_C6450_;
  assign new_C6429_ = new_C6445_ | new_C6444_;
  assign new_C6430_ = ~new_C6453_ | ~new_C6452_;
  assign new_C6431_ = ~new_C6454_ & new_C6455_;
  assign new_C6432_ = new_C6454_ & ~new_C6455_;
  assign new_C6433_ = ~new_C6401_ & new_C6402_;
  assign new_C6434_ = new_C6401_ & ~new_C6402_;
  assign new_C6435_ = ~new_C6417_ | new_C6427_;
  assign new_C6436_ = new_C6417_ & new_C6427_;
  assign new_C6437_ = ~new_C6417_ & ~new_C6427_;
  assign new_C6438_ = new_C6459_ | new_C6458_;
  assign new_C6439_ = new_C6405_ | new_C6438_;
  assign new_C6440_ = new_C6463_ | new_C6462_;
  assign new_C6441_ = ~new_C6405_ & new_C6440_;
  assign new_C6442_ = new_C6461_ | new_C6460_;
  assign new_C6443_ = new_C6405_ & new_C6442_;
  assign new_C6444_ = new_C6403_ & ~new_C6413_;
  assign new_C6445_ = ~new_C6403_ & new_C6413_;
  assign new_C6446_ = ~new_C6402_ | ~new_C6427_;
  assign new_C6447_ = new_C6413_ & new_C6446_;
  assign new_C6448_ = ~new_C6413_ & ~new_C6447_;
  assign new_C6449_ = new_C6413_ | new_C6446_;
  assign new_C6450_ = ~new_C6403_ & new_C6404_;
  assign new_C6451_ = new_C6403_ & ~new_C6404_;
  assign new_C6452_ = new_C6420_ | new_C6457_;
  assign new_C6453_ = ~new_C6420_ & ~new_C6456_;
  assign new_C6454_ = new_C6403_ | new_C6420_;
  assign new_C6455_ = new_C6403_ | new_C6404_;
  assign new_C6456_ = new_C6420_ & new_C6457_;
  assign new_C6457_ = ~new_C6402_ | ~new_C6427_;
  assign new_C6458_ = new_C6435_ & new_C6455_;
  assign new_C6459_ = ~new_C6435_ & ~new_C6455_;
  assign new_C6460_ = new_C6464_ | new_C6465_;
  assign new_C6461_ = ~new_C6406_ & new_C6420_;
  assign new_C6462_ = new_C6466_ | new_C6467_;
  assign new_C6463_ = new_C6406_ & new_C6420_;
  assign new_C6464_ = ~new_C6406_ & ~new_C6420_;
  assign new_C6465_ = new_C6406_ & ~new_C6420_;
  assign new_C6466_ = new_C6406_ & ~new_C6420_;
  assign new_C6467_ = ~new_C6406_ & new_C6420_;
  assign new_C6468_ = new_E6242_;
  assign new_C6469_ = new_E6309_;
  assign new_C6470_ = new_E6376_;
  assign new_C6471_ = new_E6443_;
  assign new_C6472_ = new_E6510_;
  assign new_C6473_ = new_E6577_;
  assign new_C6474_ = new_C6481_ & new_C6480_;
  assign new_C6475_ = new_C6483_ | new_C6482_;
  assign new_C6476_ = new_C6485_ | new_C6484_;
  assign new_C6477_ = new_C6487_ & new_C6486_;
  assign new_C6478_ = new_C6487_ & new_C6488_;
  assign new_C6479_ = new_C6480_ | new_C6489_;
  assign new_C6480_ = new_C6469_ | new_C6492_;
  assign new_C6481_ = new_C6491_ | new_C6490_;
  assign new_C6482_ = new_C6496_ & new_C6495_;
  assign new_C6483_ = new_C6494_ & new_C6493_;
  assign new_C6484_ = new_C6499_ | new_C6498_;
  assign new_C6485_ = new_C6494_ & new_C6497_;
  assign new_C6486_ = new_C6469_ | new_C6502_;
  assign new_C6487_ = new_C6501_ | new_C6500_;
  assign new_C6488_ = new_C6504_ | new_C6503_;
  assign new_C6489_ = ~new_C6480_ & new_C6506_;
  assign new_C6490_ = ~new_C6482_ & new_C6494_;
  assign new_C6491_ = new_C6482_ & ~new_C6494_;
  assign new_C6492_ = new_C6468_ & ~new_C6469_;
  assign new_C6493_ = ~new_C6515_ | ~new_C6516_;
  assign new_C6494_ = new_C6508_ | new_C6510_;
  assign new_C6495_ = new_C6518_ | new_C6517_;
  assign new_C6496_ = new_C6512_ | new_C6511_;
  assign new_C6497_ = ~new_C6520_ | ~new_C6519_;
  assign new_C6498_ = ~new_C6521_ & new_C6522_;
  assign new_C6499_ = new_C6521_ & ~new_C6522_;
  assign new_C6500_ = ~new_C6468_ & new_C6469_;
  assign new_C6501_ = new_C6468_ & ~new_C6469_;
  assign new_C6502_ = ~new_C6484_ | new_C6494_;
  assign new_C6503_ = new_C6484_ & new_C6494_;
  assign new_C6504_ = ~new_C6484_ & ~new_C6494_;
  assign new_C6505_ = new_C6526_ | new_C6525_;
  assign new_C6506_ = new_C6472_ | new_C6505_;
  assign new_C6507_ = new_C6530_ | new_C6529_;
  assign new_C6508_ = ~new_C6472_ & new_C6507_;
  assign new_C6509_ = new_C6528_ | new_C6527_;
  assign new_C6510_ = new_C6472_ & new_C6509_;
  assign new_C6511_ = new_C6470_ & ~new_C6480_;
  assign new_C6512_ = ~new_C6470_ & new_C6480_;
  assign new_C6513_ = ~new_C6469_ | ~new_C6494_;
  assign new_C6514_ = new_C6480_ & new_C6513_;
  assign new_C6515_ = ~new_C6480_ & ~new_C6514_;
  assign new_C6516_ = new_C6480_ | new_C6513_;
  assign new_C6517_ = ~new_C6470_ & new_C6471_;
  assign new_C6518_ = new_C6470_ & ~new_C6471_;
  assign new_C6519_ = new_C6487_ | new_C6524_;
  assign new_C6520_ = ~new_C6487_ & ~new_C6523_;
  assign new_C6521_ = new_C6470_ | new_C6487_;
  assign new_C6522_ = new_C6470_ | new_C6471_;
  assign new_C6523_ = new_C6487_ & new_C6524_;
  assign new_C6524_ = ~new_C6469_ | ~new_C6494_;
  assign new_C6525_ = new_C6502_ & new_C6522_;
  assign new_C6526_ = ~new_C6502_ & ~new_C6522_;
  assign new_C6527_ = new_C6531_ | new_C6532_;
  assign new_C6528_ = ~new_C6473_ & new_C6487_;
  assign new_C6529_ = new_C6533_ | new_C6534_;
  assign new_C6530_ = new_C6473_ & new_C6487_;
  assign new_C6531_ = ~new_C6473_ & ~new_C6487_;
  assign new_C6532_ = new_C6473_ & ~new_C6487_;
  assign new_C6533_ = new_C6473_ & ~new_C6487_;
  assign new_C6534_ = ~new_C6473_ & new_C6487_;
  assign new_C6535_ = new_E6644_;
  assign new_C6536_ = new_E6711_;
  assign new_C6537_ = new_E6778_;
  assign new_C6538_ = new_E6845_;
  assign new_C6539_ = new_E6912_;
  assign new_C6540_ = new_E6979_;
  assign new_C6541_ = new_C6548_ & new_C6547_;
  assign new_C6542_ = new_C6550_ | new_C6549_;
  assign new_C6543_ = new_C6552_ | new_C6551_;
  assign new_C6544_ = new_C6554_ & new_C6553_;
  assign new_C6545_ = new_C6554_ & new_C6555_;
  assign new_C6546_ = new_C6547_ | new_C6556_;
  assign new_C6547_ = new_C6536_ | new_C6559_;
  assign new_C6548_ = new_C6558_ | new_C6557_;
  assign new_C6549_ = new_C6563_ & new_C6562_;
  assign new_C6550_ = new_C6561_ & new_C6560_;
  assign new_C6551_ = new_C6566_ | new_C6565_;
  assign new_C6552_ = new_C6561_ & new_C6564_;
  assign new_C6553_ = new_C6536_ | new_C6569_;
  assign new_C6554_ = new_C6568_ | new_C6567_;
  assign new_C6555_ = new_C6571_ | new_C6570_;
  assign new_C6556_ = ~new_C6547_ & new_C6573_;
  assign new_C6557_ = ~new_C6549_ & new_C6561_;
  assign new_C6558_ = new_C6549_ & ~new_C6561_;
  assign new_C6559_ = new_C6535_ & ~new_C6536_;
  assign new_C6560_ = ~new_C6582_ | ~new_C6583_;
  assign new_C6561_ = new_C6575_ | new_C6577_;
  assign new_C6562_ = new_C6585_ | new_C6584_;
  assign new_C6563_ = new_C6579_ | new_C6578_;
  assign new_C6564_ = ~new_C6587_ | ~new_C6586_;
  assign new_C6565_ = ~new_C6588_ & new_C6589_;
  assign new_C6566_ = new_C6588_ & ~new_C6589_;
  assign new_C6567_ = ~new_C6535_ & new_C6536_;
  assign new_C6568_ = new_C6535_ & ~new_C6536_;
  assign new_C6569_ = ~new_C6551_ | new_C6561_;
  assign new_C6570_ = new_C6551_ & new_C6561_;
  assign new_C6571_ = ~new_C6551_ & ~new_C6561_;
  assign new_C6572_ = new_C6593_ | new_C6592_;
  assign new_C6573_ = new_C6539_ | new_C6572_;
  assign new_C6574_ = new_C6597_ | new_C6596_;
  assign new_C6575_ = ~new_C6539_ & new_C6574_;
  assign new_C6576_ = new_C6595_ | new_C6594_;
  assign new_C6577_ = new_C6539_ & new_C6576_;
  assign new_C6578_ = new_C6537_ & ~new_C6547_;
  assign new_C6579_ = ~new_C6537_ & new_C6547_;
  assign new_C6580_ = ~new_C6536_ | ~new_C6561_;
  assign new_C6581_ = new_C6547_ & new_C6580_;
  assign new_C6582_ = ~new_C6547_ & ~new_C6581_;
  assign new_C6583_ = new_C6547_ | new_C6580_;
  assign new_C6584_ = ~new_C6537_ & new_C6538_;
  assign new_C6585_ = new_C6537_ & ~new_C6538_;
  assign new_C6586_ = new_C6554_ | new_C6591_;
  assign new_C6587_ = ~new_C6554_ & ~new_C6590_;
  assign new_C6588_ = new_C6537_ | new_C6554_;
  assign new_C6589_ = new_C6537_ | new_C6538_;
  assign new_C6590_ = new_C6554_ & new_C6591_;
  assign new_C6591_ = ~new_C6536_ | ~new_C6561_;
  assign new_C6592_ = new_C6569_ & new_C6589_;
  assign new_C6593_ = ~new_C6569_ & ~new_C6589_;
  assign new_C6594_ = new_C6598_ | new_C6599_;
  assign new_C6595_ = ~new_C6540_ & new_C6554_;
  assign new_C6596_ = new_C6600_ | new_C6601_;
  assign new_C6597_ = new_C6540_ & new_C6554_;
  assign new_C6598_ = ~new_C6540_ & ~new_C6554_;
  assign new_C6599_ = new_C6540_ & ~new_C6554_;
  assign new_C6600_ = new_C6540_ & ~new_C6554_;
  assign new_C6601_ = ~new_C6540_ & new_C6554_;
  assign new_C6602_ = new_E7046_;
  assign new_C6603_ = new_E7113_;
  assign new_C6604_ = new_E7180_;
  assign new_C6605_ = new_E7247_;
  assign new_C6606_ = new_E7314_;
  assign new_C6607_ = new_E7381_;
  assign new_C6608_ = new_C6615_ & new_C6614_;
  assign new_C6609_ = new_C6617_ | new_C6616_;
  assign new_C6610_ = new_C6619_ | new_C6618_;
  assign new_C6611_ = new_C6621_ & new_C6620_;
  assign new_C6612_ = new_C6621_ & new_C6622_;
  assign new_C6613_ = new_C6614_ | new_C6623_;
  assign new_C6614_ = new_C6603_ | new_C6626_;
  assign new_C6615_ = new_C6625_ | new_C6624_;
  assign new_C6616_ = new_C6630_ & new_C6629_;
  assign new_C6617_ = new_C6628_ & new_C6627_;
  assign new_C6618_ = new_C6633_ | new_C6632_;
  assign new_C6619_ = new_C6628_ & new_C6631_;
  assign new_C6620_ = new_C6603_ | new_C6636_;
  assign new_C6621_ = new_C6635_ | new_C6634_;
  assign new_C6622_ = new_C6638_ | new_C6637_;
  assign new_C6623_ = ~new_C6614_ & new_C6640_;
  assign new_C6624_ = ~new_C6616_ & new_C6628_;
  assign new_C6625_ = new_C6616_ & ~new_C6628_;
  assign new_C6626_ = new_C6602_ & ~new_C6603_;
  assign new_C6627_ = ~new_C6649_ | ~new_C6650_;
  assign new_C6628_ = new_C6642_ | new_C6644_;
  assign new_C6629_ = new_C6652_ | new_C6651_;
  assign new_C6630_ = new_C6646_ | new_C6645_;
  assign new_C6631_ = ~new_C6654_ | ~new_C6653_;
  assign new_C6632_ = ~new_C6655_ & new_C6656_;
  assign new_C6633_ = new_C6655_ & ~new_C6656_;
  assign new_C6634_ = ~new_C6602_ & new_C6603_;
  assign new_C6635_ = new_C6602_ & ~new_C6603_;
  assign new_C6636_ = ~new_C6618_ | new_C6628_;
  assign new_C6637_ = new_C6618_ & new_C6628_;
  assign new_C6638_ = ~new_C6618_ & ~new_C6628_;
  assign new_C6639_ = new_C6660_ | new_C6659_;
  assign new_C6640_ = new_C6606_ | new_C6639_;
  assign new_C6641_ = new_C6664_ | new_C6663_;
  assign new_C6642_ = ~new_C6606_ & new_C6641_;
  assign new_C6643_ = new_C6662_ | new_C6661_;
  assign new_C6644_ = new_C6606_ & new_C6643_;
  assign new_C6645_ = new_C6604_ & ~new_C6614_;
  assign new_C6646_ = ~new_C6604_ & new_C6614_;
  assign new_C6647_ = ~new_C6603_ | ~new_C6628_;
  assign new_C6648_ = new_C6614_ & new_C6647_;
  assign new_C6649_ = ~new_C6614_ & ~new_C6648_;
  assign new_C6650_ = new_C6614_ | new_C6647_;
  assign new_C6651_ = ~new_C6604_ & new_C6605_;
  assign new_C6652_ = new_C6604_ & ~new_C6605_;
  assign new_C6653_ = new_C6621_ | new_C6658_;
  assign new_C6654_ = ~new_C6621_ & ~new_C6657_;
  assign new_C6655_ = new_C6604_ | new_C6621_;
  assign new_C6656_ = new_C6604_ | new_C6605_;
  assign new_C6657_ = new_C6621_ & new_C6658_;
  assign new_C6658_ = ~new_C6603_ | ~new_C6628_;
  assign new_C6659_ = new_C6636_ & new_C6656_;
  assign new_C6660_ = ~new_C6636_ & ~new_C6656_;
  assign new_C6661_ = new_C6665_ | new_C6666_;
  assign new_C6662_ = ~new_C6607_ & new_C6621_;
  assign new_C6663_ = new_C6667_ | new_C6668_;
  assign new_C6664_ = new_C6607_ & new_C6621_;
  assign new_C6665_ = ~new_C6607_ & ~new_C6621_;
  assign new_C6666_ = new_C6607_ & ~new_C6621_;
  assign new_C6667_ = new_C6607_ & ~new_C6621_;
  assign new_C6668_ = ~new_C6607_ & new_C6621_;
  assign new_C6669_ = new_E7448_;
  assign new_C6670_ = new_E7515_;
  assign new_C6671_ = new_E7582_;
  assign new_C6672_ = new_E7649_;
  assign new_C6673_ = new_E7716_;
  assign new_C6674_ = new_E7783_;
  assign new_C6675_ = new_C6682_ & new_C6681_;
  assign new_C6676_ = new_C6684_ | new_C6683_;
  assign new_C6677_ = new_C6686_ | new_C6685_;
  assign new_C6678_ = new_C6688_ & new_C6687_;
  assign new_C6679_ = new_C6688_ & new_C6689_;
  assign new_C6680_ = new_C6681_ | new_C6690_;
  assign new_C6681_ = new_C6670_ | new_C6693_;
  assign new_C6682_ = new_C6692_ | new_C6691_;
  assign new_C6683_ = new_C6697_ & new_C6696_;
  assign new_C6684_ = new_C6695_ & new_C6694_;
  assign new_C6685_ = new_C6700_ | new_C6699_;
  assign new_C6686_ = new_C6695_ & new_C6698_;
  assign new_C6687_ = new_C6670_ | new_C6703_;
  assign new_C6688_ = new_C6702_ | new_C6701_;
  assign new_C6689_ = new_C6705_ | new_C6704_;
  assign new_C6690_ = ~new_C6681_ & new_C6707_;
  assign new_C6691_ = ~new_C6683_ & new_C6695_;
  assign new_C6692_ = new_C6683_ & ~new_C6695_;
  assign new_C6693_ = new_C6669_ & ~new_C6670_;
  assign new_C6694_ = ~new_C6716_ | ~new_C6717_;
  assign new_C6695_ = new_C6709_ | new_C6711_;
  assign new_C6696_ = new_C6719_ | new_C6718_;
  assign new_C6697_ = new_C6713_ | new_C6712_;
  assign new_C6698_ = ~new_C6721_ | ~new_C6720_;
  assign new_C6699_ = ~new_C6722_ & new_C6723_;
  assign new_C6700_ = new_C6722_ & ~new_C6723_;
  assign new_C6701_ = ~new_C6669_ & new_C6670_;
  assign new_C6702_ = new_C6669_ & ~new_C6670_;
  assign new_C6703_ = ~new_C6685_ | new_C6695_;
  assign new_C6704_ = new_C6685_ & new_C6695_;
  assign new_C6705_ = ~new_C6685_ & ~new_C6695_;
  assign new_C6706_ = new_C6727_ | new_C6726_;
  assign new_C6707_ = new_C6673_ | new_C6706_;
  assign new_C6708_ = new_C6731_ | new_C6730_;
  assign new_C6709_ = ~new_C6673_ & new_C6708_;
  assign new_C6710_ = new_C6729_ | new_C6728_;
  assign new_C6711_ = new_C6673_ & new_C6710_;
  assign new_C6712_ = new_C6671_ & ~new_C6681_;
  assign new_C6713_ = ~new_C6671_ & new_C6681_;
  assign new_C6714_ = ~new_C6670_ | ~new_C6695_;
  assign new_C6715_ = new_C6681_ & new_C6714_;
  assign new_C6716_ = ~new_C6681_ & ~new_C6715_;
  assign new_C6717_ = new_C6681_ | new_C6714_;
  assign new_C6718_ = ~new_C6671_ & new_C6672_;
  assign new_C6719_ = new_C6671_ & ~new_C6672_;
  assign new_C6720_ = new_C6688_ | new_C6725_;
  assign new_C6721_ = ~new_C6688_ & ~new_C6724_;
  assign new_C6722_ = new_C6671_ | new_C6688_;
  assign new_C6723_ = new_C6671_ | new_C6672_;
  assign new_C6724_ = new_C6688_ & new_C6725_;
  assign new_C6725_ = ~new_C6670_ | ~new_C6695_;
  assign new_C6726_ = new_C6703_ & new_C6723_;
  assign new_C6727_ = ~new_C6703_ & ~new_C6723_;
  assign new_C6728_ = new_C6732_ | new_C6733_;
  assign new_C6729_ = ~new_C6674_ & new_C6688_;
  assign new_C6730_ = new_C6734_ | new_C6735_;
  assign new_C6731_ = new_C6674_ & new_C6688_;
  assign new_C6732_ = ~new_C6674_ & ~new_C6688_;
  assign new_C6733_ = new_C6674_ & ~new_C6688_;
  assign new_C6734_ = new_C6674_ & ~new_C6688_;
  assign new_C6735_ = ~new_C6674_ & new_C6688_;
  assign new_C6736_ = new_E7850_;
  assign new_C6737_ = new_E7917_;
  assign new_C6738_ = new_E7984_;
  assign new_C6739_ = new_E8051_;
  assign new_C6740_ = new_E8118_;
  assign new_C6741_ = new_E8185_;
  assign new_C6742_ = new_C6749_ & new_C6748_;
  assign new_C6743_ = new_C6751_ | new_C6750_;
  assign new_C6744_ = new_C6753_ | new_C6752_;
  assign new_C6745_ = new_C6755_ & new_C6754_;
  assign new_C6746_ = new_C6755_ & new_C6756_;
  assign new_C6747_ = new_C6748_ | new_C6757_;
  assign new_C6748_ = new_C6737_ | new_C6760_;
  assign new_C6749_ = new_C6759_ | new_C6758_;
  assign new_C6750_ = new_C6764_ & new_C6763_;
  assign new_C6751_ = new_C6762_ & new_C6761_;
  assign new_C6752_ = new_C6767_ | new_C6766_;
  assign new_C6753_ = new_C6762_ & new_C6765_;
  assign new_C6754_ = new_C6737_ | new_C6770_;
  assign new_C6755_ = new_C6769_ | new_C6768_;
  assign new_C6756_ = new_C6772_ | new_C6771_;
  assign new_C6757_ = ~new_C6748_ & new_C6774_;
  assign new_C6758_ = ~new_C6750_ & new_C6762_;
  assign new_C6759_ = new_C6750_ & ~new_C6762_;
  assign new_C6760_ = new_C6736_ & ~new_C6737_;
  assign new_C6761_ = ~new_C6783_ | ~new_C6784_;
  assign new_C6762_ = new_C6776_ | new_C6778_;
  assign new_C6763_ = new_C6786_ | new_C6785_;
  assign new_C6764_ = new_C6780_ | new_C6779_;
  assign new_C6765_ = ~new_C6788_ | ~new_C6787_;
  assign new_C6766_ = ~new_C6789_ & new_C6790_;
  assign new_C6767_ = new_C6789_ & ~new_C6790_;
  assign new_C6768_ = ~new_C6736_ & new_C6737_;
  assign new_C6769_ = new_C6736_ & ~new_C6737_;
  assign new_C6770_ = ~new_C6752_ | new_C6762_;
  assign new_C6771_ = new_C6752_ & new_C6762_;
  assign new_C6772_ = ~new_C6752_ & ~new_C6762_;
  assign new_C6773_ = new_C6794_ | new_C6793_;
  assign new_C6774_ = new_C6740_ | new_C6773_;
  assign new_C6775_ = new_C6798_ | new_C6797_;
  assign new_C6776_ = ~new_C6740_ & new_C6775_;
  assign new_C6777_ = new_C6796_ | new_C6795_;
  assign new_C6778_ = new_C6740_ & new_C6777_;
  assign new_C6779_ = new_C6738_ & ~new_C6748_;
  assign new_C6780_ = ~new_C6738_ & new_C6748_;
  assign new_C6781_ = ~new_C6737_ | ~new_C6762_;
  assign new_C6782_ = new_C6748_ & new_C6781_;
  assign new_C6783_ = ~new_C6748_ & ~new_C6782_;
  assign new_C6784_ = new_C6748_ | new_C6781_;
  assign new_C6785_ = ~new_C6738_ & new_C6739_;
  assign new_C6786_ = new_C6738_ & ~new_C6739_;
  assign new_C6787_ = new_C6755_ | new_C6792_;
  assign new_C6788_ = ~new_C6755_ & ~new_C6791_;
  assign new_C6789_ = new_C6738_ | new_C6755_;
  assign new_C6790_ = new_C6738_ | new_C6739_;
  assign new_C6791_ = new_C6755_ & new_C6792_;
  assign new_C6792_ = ~new_C6737_ | ~new_C6762_;
  assign new_C6793_ = new_C6770_ & new_C6790_;
  assign new_C6794_ = ~new_C6770_ & ~new_C6790_;
  assign new_C6795_ = new_C6799_ | new_C6800_;
  assign new_C6796_ = ~new_C6741_ & new_C6755_;
  assign new_C6797_ = new_C6801_ | new_C6802_;
  assign new_C6798_ = new_C6741_ & new_C6755_;
  assign new_C6799_ = ~new_C6741_ & ~new_C6755_;
  assign new_C6800_ = new_C6741_ & ~new_C6755_;
  assign new_C6801_ = new_C6741_ & ~new_C6755_;
  assign new_C6802_ = ~new_C6741_ & new_C6755_;
  assign new_C6803_ = new_E8252_;
  assign new_C6804_ = new_E8319_;
  assign new_C6805_ = new_E8386_;
  assign new_C6806_ = new_E8453_;
  assign new_C6807_ = new_E8520_;
  assign new_C6808_ = new_E8587_;
  assign new_C6809_ = new_C6816_ & new_C6815_;
  assign new_C6810_ = new_C6818_ | new_C6817_;
  assign new_C6811_ = new_C6820_ | new_C6819_;
  assign new_C6812_ = new_C6822_ & new_C6821_;
  assign new_C6813_ = new_C6822_ & new_C6823_;
  assign new_C6814_ = new_C6815_ | new_C6824_;
  assign new_C6815_ = new_C6804_ | new_C6827_;
  assign new_C6816_ = new_C6826_ | new_C6825_;
  assign new_C6817_ = new_C6831_ & new_C6830_;
  assign new_C6818_ = new_C6829_ & new_C6828_;
  assign new_C6819_ = new_C6834_ | new_C6833_;
  assign new_C6820_ = new_C6829_ & new_C6832_;
  assign new_C6821_ = new_C6804_ | new_C6837_;
  assign new_C6822_ = new_C6836_ | new_C6835_;
  assign new_C6823_ = new_C6839_ | new_C6838_;
  assign new_C6824_ = ~new_C6815_ & new_C6841_;
  assign new_C6825_ = ~new_C6817_ & new_C6829_;
  assign new_C6826_ = new_C6817_ & ~new_C6829_;
  assign new_C6827_ = new_C6803_ & ~new_C6804_;
  assign new_C6828_ = ~new_C6850_ | ~new_C6851_;
  assign new_C6829_ = new_C6843_ | new_C6845_;
  assign new_C6830_ = new_C6853_ | new_C6852_;
  assign new_C6831_ = new_C6847_ | new_C6846_;
  assign new_C6832_ = ~new_C6855_ | ~new_C6854_;
  assign new_C6833_ = ~new_C6856_ & new_C6857_;
  assign new_C6834_ = new_C6856_ & ~new_C6857_;
  assign new_C6835_ = ~new_C6803_ & new_C6804_;
  assign new_C6836_ = new_C6803_ & ~new_C6804_;
  assign new_C6837_ = ~new_C6819_ | new_C6829_;
  assign new_C6838_ = new_C6819_ & new_C6829_;
  assign new_C6839_ = ~new_C6819_ & ~new_C6829_;
  assign new_C6840_ = new_C6861_ | new_C6860_;
  assign new_C6841_ = new_C6807_ | new_C6840_;
  assign new_C6842_ = new_C6865_ | new_C6864_;
  assign new_C6843_ = ~new_C6807_ & new_C6842_;
  assign new_C6844_ = new_C6863_ | new_C6862_;
  assign new_C6845_ = new_C6807_ & new_C6844_;
  assign new_C6846_ = new_C6805_ & ~new_C6815_;
  assign new_C6847_ = ~new_C6805_ & new_C6815_;
  assign new_C6848_ = ~new_C6804_ | ~new_C6829_;
  assign new_C6849_ = new_C6815_ & new_C6848_;
  assign new_C6850_ = ~new_C6815_ & ~new_C6849_;
  assign new_C6851_ = new_C6815_ | new_C6848_;
  assign new_C6852_ = ~new_C6805_ & new_C6806_;
  assign new_C6853_ = new_C6805_ & ~new_C6806_;
  assign new_C6854_ = new_C6822_ | new_C6859_;
  assign new_C6855_ = ~new_C6822_ & ~new_C6858_;
  assign new_C6856_ = new_C6805_ | new_C6822_;
  assign new_C6857_ = new_C6805_ | new_C6806_;
  assign new_C6858_ = new_C6822_ & new_C6859_;
  assign new_C6859_ = ~new_C6804_ | ~new_C6829_;
  assign new_C6860_ = new_C6837_ & new_C6857_;
  assign new_C6861_ = ~new_C6837_ & ~new_C6857_;
  assign new_C6862_ = new_C6866_ | new_C6867_;
  assign new_C6863_ = ~new_C6808_ & new_C6822_;
  assign new_C6864_ = new_C6868_ | new_C6869_;
  assign new_C6865_ = new_C6808_ & new_C6822_;
  assign new_C6866_ = ~new_C6808_ & ~new_C6822_;
  assign new_C6867_ = new_C6808_ & ~new_C6822_;
  assign new_C6868_ = new_C6808_ & ~new_C6822_;
  assign new_C6869_ = ~new_C6808_ & new_C6822_;
  assign new_C6870_ = new_E8654_;
  assign new_C6871_ = new_E8721_;
  assign new_C6872_ = new_E8788_;
  assign new_C6873_ = new_E8855_;
  assign new_C6874_ = new_E8922_;
  assign new_C6875_ = new_E8989_;
  assign new_C6876_ = new_C6883_ & new_C6882_;
  assign new_C6877_ = new_C6885_ | new_C6884_;
  assign new_C6878_ = new_C6887_ | new_C6886_;
  assign new_C6879_ = new_C6889_ & new_C6888_;
  assign new_C6880_ = new_C6889_ & new_C6890_;
  assign new_C6881_ = new_C6882_ | new_C6891_;
  assign new_C6882_ = new_C6871_ | new_C6894_;
  assign new_C6883_ = new_C6893_ | new_C6892_;
  assign new_C6884_ = new_C6898_ & new_C6897_;
  assign new_C6885_ = new_C6896_ & new_C6895_;
  assign new_C6886_ = new_C6901_ | new_C6900_;
  assign new_C6887_ = new_C6896_ & new_C6899_;
  assign new_C6888_ = new_C6871_ | new_C6904_;
  assign new_C6889_ = new_C6903_ | new_C6902_;
  assign new_C6890_ = new_C6906_ | new_C6905_;
  assign new_C6891_ = ~new_C6882_ & new_C6908_;
  assign new_C6892_ = ~new_C6884_ & new_C6896_;
  assign new_C6893_ = new_C6884_ & ~new_C6896_;
  assign new_C6894_ = new_C6870_ & ~new_C6871_;
  assign new_C6895_ = ~new_C6917_ | ~new_C6918_;
  assign new_C6896_ = new_C6910_ | new_C6912_;
  assign new_C6897_ = new_C6920_ | new_C6919_;
  assign new_C6898_ = new_C6914_ | new_C6913_;
  assign new_C6899_ = ~new_C6922_ | ~new_C6921_;
  assign new_C6900_ = ~new_C6923_ & new_C6924_;
  assign new_C6901_ = new_C6923_ & ~new_C6924_;
  assign new_C6902_ = ~new_C6870_ & new_C6871_;
  assign new_C6903_ = new_C6870_ & ~new_C6871_;
  assign new_C6904_ = ~new_C6886_ | new_C6896_;
  assign new_C6905_ = new_C6886_ & new_C6896_;
  assign new_C6906_ = ~new_C6886_ & ~new_C6896_;
  assign new_C6907_ = new_C6928_ | new_C6927_;
  assign new_C6908_ = new_C6874_ | new_C6907_;
  assign new_C6909_ = new_C6932_ | new_C6931_;
  assign new_C6910_ = ~new_C6874_ & new_C6909_;
  assign new_C6911_ = new_C6930_ | new_C6929_;
  assign new_C6912_ = new_C6874_ & new_C6911_;
  assign new_C6913_ = new_C6872_ & ~new_C6882_;
  assign new_C6914_ = ~new_C6872_ & new_C6882_;
  assign new_C6915_ = ~new_C6871_ | ~new_C6896_;
  assign new_C6916_ = new_C6882_ & new_C6915_;
  assign new_C6917_ = ~new_C6882_ & ~new_C6916_;
  assign new_C6918_ = new_C6882_ | new_C6915_;
  assign new_C6919_ = ~new_C6872_ & new_C6873_;
  assign new_C6920_ = new_C6872_ & ~new_C6873_;
  assign new_C6921_ = new_C6889_ | new_C6926_;
  assign new_C6922_ = ~new_C6889_ & ~new_C6925_;
  assign new_C6923_ = new_C6872_ | new_C6889_;
  assign new_C6924_ = new_C6872_ | new_C6873_;
  assign new_C6925_ = new_C6889_ & new_C6926_;
  assign new_C6926_ = ~new_C6871_ | ~new_C6896_;
  assign new_C6927_ = new_C6904_ & new_C6924_;
  assign new_C6928_ = ~new_C6904_ & ~new_C6924_;
  assign new_C6929_ = new_C6933_ | new_C6934_;
  assign new_C6930_ = ~new_C6875_ & new_C6889_;
  assign new_C6931_ = new_C6935_ | new_C6936_;
  assign new_C6932_ = new_C6875_ & new_C6889_;
  assign new_C6933_ = ~new_C6875_ & ~new_C6889_;
  assign new_C6934_ = new_C6875_ & ~new_C6889_;
  assign new_C6935_ = new_C6875_ & ~new_C6889_;
  assign new_C6936_ = ~new_C6875_ & new_C6889_;
  assign new_C6937_ = new_E9056_;
  assign new_C6938_ = new_E9123_;
  assign new_C6939_ = new_E9190_;
  assign new_C6940_ = new_E9257_;
  assign new_C6941_ = new_E9324_;
  assign new_C6942_ = new_E9391_;
  assign new_C6943_ = new_C6950_ & new_C6949_;
  assign new_C6944_ = new_C6952_ | new_C6951_;
  assign new_C6945_ = new_C6954_ | new_C6953_;
  assign new_C6946_ = new_C6956_ & new_C6955_;
  assign new_C6947_ = new_C6956_ & new_C6957_;
  assign new_C6948_ = new_C6949_ | new_C6958_;
  assign new_C6949_ = new_C6938_ | new_C6961_;
  assign new_C6950_ = new_C6960_ | new_C6959_;
  assign new_C6951_ = new_C6965_ & new_C6964_;
  assign new_C6952_ = new_C6963_ & new_C6962_;
  assign new_C6953_ = new_C6968_ | new_C6967_;
  assign new_C6954_ = new_C6963_ & new_C6966_;
  assign new_C6955_ = new_C6938_ | new_C6971_;
  assign new_C6956_ = new_C6970_ | new_C6969_;
  assign new_C6957_ = new_C6973_ | new_C6972_;
  assign new_C6958_ = ~new_C6949_ & new_C6975_;
  assign new_C6959_ = ~new_C6951_ & new_C6963_;
  assign new_C6960_ = new_C6951_ & ~new_C6963_;
  assign new_C6961_ = new_C6937_ & ~new_C6938_;
  assign new_C6962_ = ~new_C6984_ | ~new_C6985_;
  assign new_C6963_ = new_C6977_ | new_C6979_;
  assign new_C6964_ = new_C6987_ | new_C6986_;
  assign new_C6965_ = new_C6981_ | new_C6980_;
  assign new_C6966_ = ~new_C6989_ | ~new_C6988_;
  assign new_C6967_ = ~new_C6990_ & new_C6991_;
  assign new_C6968_ = new_C6990_ & ~new_C6991_;
  assign new_C6969_ = ~new_C6937_ & new_C6938_;
  assign new_C6970_ = new_C6937_ & ~new_C6938_;
  assign new_C6971_ = ~new_C6953_ | new_C6963_;
  assign new_C6972_ = new_C6953_ & new_C6963_;
  assign new_C6973_ = ~new_C6953_ & ~new_C6963_;
  assign new_C6974_ = new_C6995_ | new_C6994_;
  assign new_C6975_ = new_C6941_ | new_C6974_;
  assign new_C6976_ = new_C6999_ | new_C6998_;
  assign new_C6977_ = ~new_C6941_ & new_C6976_;
  assign new_C6978_ = new_C6997_ | new_C6996_;
  assign new_C6979_ = new_C6941_ & new_C6978_;
  assign new_C6980_ = new_C6939_ & ~new_C6949_;
  assign new_C6981_ = ~new_C6939_ & new_C6949_;
  assign new_C6982_ = ~new_C6938_ | ~new_C6963_;
  assign new_C6983_ = new_C6949_ & new_C6982_;
  assign new_C6984_ = ~new_C6949_ & ~new_C6983_;
  assign new_C6985_ = new_C6949_ | new_C6982_;
  assign new_C6986_ = ~new_C6939_ & new_C6940_;
  assign new_C6987_ = new_C6939_ & ~new_C6940_;
  assign new_C6988_ = new_C6956_ | new_C6993_;
  assign new_C6989_ = ~new_C6956_ & ~new_C6992_;
  assign new_C6990_ = new_C6939_ | new_C6956_;
  assign new_C6991_ = new_C6939_ | new_C6940_;
  assign new_C6992_ = new_C6956_ & new_C6993_;
  assign new_C6993_ = ~new_C6938_ | ~new_C6963_;
  assign new_C6994_ = new_C6971_ & new_C6991_;
  assign new_C6995_ = ~new_C6971_ & ~new_C6991_;
  assign new_C6996_ = new_C7000_ | new_C7001_;
  assign new_C6997_ = ~new_C6942_ & new_C6956_;
  assign new_C6998_ = new_C7002_ | new_C7003_;
  assign new_C6999_ = new_C6942_ & new_C6956_;
  assign new_C7000_ = ~new_C6942_ & ~new_C6956_;
  assign new_C7001_ = new_C6942_ & ~new_C6956_;
  assign new_C7002_ = new_C6942_ & ~new_C6956_;
  assign new_C7003_ = ~new_C6942_ & new_C6956_;
  assign new_C7004_ = new_E9458_;
  assign new_C7005_ = new_E9525_;
  assign new_C7006_ = new_E9592_;
  assign new_C7007_ = new_E9659_;
  assign new_C7008_ = new_E9726_;
  assign new_C7009_ = new_E9793_;
  assign new_C7010_ = new_C7017_ & new_C7016_;
  assign new_C7011_ = new_C7019_ | new_C7018_;
  assign new_C7012_ = new_C7021_ | new_C7020_;
  assign new_C7013_ = new_C7023_ & new_C7022_;
  assign new_C7014_ = new_C7023_ & new_C7024_;
  assign new_C7015_ = new_C7016_ | new_C7025_;
  assign new_C7016_ = new_C7005_ | new_C7028_;
  assign new_C7017_ = new_C7027_ | new_C7026_;
  assign new_C7018_ = new_C7032_ & new_C7031_;
  assign new_C7019_ = new_C7030_ & new_C7029_;
  assign new_C7020_ = new_C7035_ | new_C7034_;
  assign new_C7021_ = new_C7030_ & new_C7033_;
  assign new_C7022_ = new_C7005_ | new_C7038_;
  assign new_C7023_ = new_C7037_ | new_C7036_;
  assign new_C7024_ = new_C7040_ | new_C7039_;
  assign new_C7025_ = ~new_C7016_ & new_C7042_;
  assign new_C7026_ = ~new_C7018_ & new_C7030_;
  assign new_C7027_ = new_C7018_ & ~new_C7030_;
  assign new_C7028_ = new_C7004_ & ~new_C7005_;
  assign new_C7029_ = ~new_C7051_ | ~new_C7052_;
  assign new_C7030_ = new_C7044_ | new_C7046_;
  assign new_C7031_ = new_C7054_ | new_C7053_;
  assign new_C7032_ = new_C7048_ | new_C7047_;
  assign new_C7033_ = ~new_C7056_ | ~new_C7055_;
  assign new_C7034_ = ~new_C7057_ & new_C7058_;
  assign new_C7035_ = new_C7057_ & ~new_C7058_;
  assign new_C7036_ = ~new_C7004_ & new_C7005_;
  assign new_C7037_ = new_C7004_ & ~new_C7005_;
  assign new_C7038_ = ~new_C7020_ | new_C7030_;
  assign new_C7039_ = new_C7020_ & new_C7030_;
  assign new_C7040_ = ~new_C7020_ & ~new_C7030_;
  assign new_C7041_ = new_C7062_ | new_C7061_;
  assign new_C7042_ = new_C7008_ | new_C7041_;
  assign new_C7043_ = new_C7066_ | new_C7065_;
  assign new_C7044_ = ~new_C7008_ & new_C7043_;
  assign new_C7045_ = new_C7064_ | new_C7063_;
  assign new_C7046_ = new_C7008_ & new_C7045_;
  assign new_C7047_ = new_C7006_ & ~new_C7016_;
  assign new_C7048_ = ~new_C7006_ & new_C7016_;
  assign new_C7049_ = ~new_C7005_ | ~new_C7030_;
  assign new_C7050_ = new_C7016_ & new_C7049_;
  assign new_C7051_ = ~new_C7016_ & ~new_C7050_;
  assign new_C7052_ = new_C7016_ | new_C7049_;
  assign new_C7053_ = ~new_C7006_ & new_C7007_;
  assign new_C7054_ = new_C7006_ & ~new_C7007_;
  assign new_C7055_ = new_C7023_ | new_C7060_;
  assign new_C7056_ = ~new_C7023_ & ~new_C7059_;
  assign new_C7057_ = new_C7006_ | new_C7023_;
  assign new_C7058_ = new_C7006_ | new_C7007_;
  assign new_C7059_ = new_C7023_ & new_C7060_;
  assign new_C7060_ = ~new_C7005_ | ~new_C7030_;
  assign new_C7061_ = new_C7038_ & new_C7058_;
  assign new_C7062_ = ~new_C7038_ & ~new_C7058_;
  assign new_C7063_ = new_C7067_ | new_C7068_;
  assign new_C7064_ = ~new_C7009_ & new_C7023_;
  assign new_C7065_ = new_C7069_ | new_C7070_;
  assign new_C7066_ = new_C7009_ & new_C7023_;
  assign new_C7067_ = ~new_C7009_ & ~new_C7023_;
  assign new_C7068_ = new_C7009_ & ~new_C7023_;
  assign new_C7069_ = new_C7009_ & ~new_C7023_;
  assign new_C7070_ = ~new_C7009_ & new_C7023_;
  assign new_C7071_ = new_E9860_;
  assign new_C7072_ = new_E9927_;
  assign new_C7073_ = new_E9994_;
  assign new_C7074_ = new_F62_;
  assign new_C7075_ = new_F129_;
  assign new_C7076_ = new_F196_;
  assign new_C7077_ = new_C7084_ & new_C7083_;
  assign new_C7078_ = new_C7086_ | new_C7085_;
  assign new_C7079_ = new_C7088_ | new_C7087_;
  assign new_C7080_ = new_C7090_ & new_C7089_;
  assign new_C7081_ = new_C7090_ & new_C7091_;
  assign new_C7082_ = new_C7083_ | new_C7092_;
  assign new_C7083_ = new_C7072_ | new_C7095_;
  assign new_C7084_ = new_C7094_ | new_C7093_;
  assign new_C7085_ = new_C7099_ & new_C7098_;
  assign new_C7086_ = new_C7097_ & new_C7096_;
  assign new_C7087_ = new_C7102_ | new_C7101_;
  assign new_C7088_ = new_C7097_ & new_C7100_;
  assign new_C7089_ = new_C7072_ | new_C7105_;
  assign new_C7090_ = new_C7104_ | new_C7103_;
  assign new_C7091_ = new_C7107_ | new_C7106_;
  assign new_C7092_ = ~new_C7083_ & new_C7109_;
  assign new_C7093_ = ~new_C7085_ & new_C7097_;
  assign new_C7094_ = new_C7085_ & ~new_C7097_;
  assign new_C7095_ = new_C7071_ & ~new_C7072_;
  assign new_C7096_ = ~new_C7118_ | ~new_C7119_;
  assign new_C7097_ = new_C7111_ | new_C7113_;
  assign new_C7098_ = new_C7121_ | new_C7120_;
  assign new_C7099_ = new_C7115_ | new_C7114_;
  assign new_C7100_ = ~new_C7123_ | ~new_C7122_;
  assign new_C7101_ = ~new_C7124_ & new_C7125_;
  assign new_C7102_ = new_C7124_ & ~new_C7125_;
  assign new_C7103_ = ~new_C7071_ & new_C7072_;
  assign new_C7104_ = new_C7071_ & ~new_C7072_;
  assign new_C7105_ = ~new_C7087_ | new_C7097_;
  assign new_C7106_ = new_C7087_ & new_C7097_;
  assign new_C7107_ = ~new_C7087_ & ~new_C7097_;
  assign new_C7108_ = new_C7129_ | new_C7128_;
  assign new_C7109_ = new_C7075_ | new_C7108_;
  assign new_C7110_ = new_C7133_ | new_C7132_;
  assign new_C7111_ = ~new_C7075_ & new_C7110_;
  assign new_C7112_ = new_C7131_ | new_C7130_;
  assign new_C7113_ = new_C7075_ & new_C7112_;
  assign new_C7114_ = new_C7073_ & ~new_C7083_;
  assign new_C7115_ = ~new_C7073_ & new_C7083_;
  assign new_C7116_ = ~new_C7072_ | ~new_C7097_;
  assign new_C7117_ = new_C7083_ & new_C7116_;
  assign new_C7118_ = ~new_C7083_ & ~new_C7117_;
  assign new_C7119_ = new_C7083_ | new_C7116_;
  assign new_C7120_ = ~new_C7073_ & new_C7074_;
  assign new_C7121_ = new_C7073_ & ~new_C7074_;
  assign new_C7122_ = new_C7090_ | new_C7127_;
  assign new_C7123_ = ~new_C7090_ & ~new_C7126_;
  assign new_C7124_ = new_C7073_ | new_C7090_;
  assign new_C7125_ = new_C7073_ | new_C7074_;
  assign new_C7126_ = new_C7090_ & new_C7127_;
  assign new_C7127_ = ~new_C7072_ | ~new_C7097_;
  assign new_C7128_ = new_C7105_ & new_C7125_;
  assign new_C7129_ = ~new_C7105_ & ~new_C7125_;
  assign new_C7130_ = new_C7134_ | new_C7135_;
  assign new_C7131_ = ~new_C7076_ & new_C7090_;
  assign new_C7132_ = new_C7136_ | new_C7137_;
  assign new_C7133_ = new_C7076_ & new_C7090_;
  assign new_C7134_ = ~new_C7076_ & ~new_C7090_;
  assign new_C7135_ = new_C7076_ & ~new_C7090_;
  assign new_C7136_ = new_C7076_ & ~new_C7090_;
  assign new_C7137_ = ~new_C7076_ & new_C7090_;
  assign new_C7138_ = new_F263_;
  assign new_C7139_ = new_F330_;
  assign new_C7140_ = new_F397_;
  assign new_C7141_ = new_F464_;
  assign new_C7142_ = new_F531_;
  assign new_C7143_ = new_F598_;
  assign new_C7144_ = new_C7151_ & new_C7150_;
  assign new_C7145_ = new_C7153_ | new_C7152_;
  assign new_C7146_ = new_C7155_ | new_C7154_;
  assign new_C7147_ = new_C7157_ & new_C7156_;
  assign new_C7148_ = new_C7157_ & new_C7158_;
  assign new_C7149_ = new_C7150_ | new_C7159_;
  assign new_C7150_ = new_C7139_ | new_C7162_;
  assign new_C7151_ = new_C7161_ | new_C7160_;
  assign new_C7152_ = new_C7166_ & new_C7165_;
  assign new_C7153_ = new_C7164_ & new_C7163_;
  assign new_C7154_ = new_C7169_ | new_C7168_;
  assign new_C7155_ = new_C7164_ & new_C7167_;
  assign new_C7156_ = new_C7139_ | new_C7172_;
  assign new_C7157_ = new_C7171_ | new_C7170_;
  assign new_C7158_ = new_C7174_ | new_C7173_;
  assign new_C7159_ = ~new_C7150_ & new_C7176_;
  assign new_C7160_ = ~new_C7152_ & new_C7164_;
  assign new_C7161_ = new_C7152_ & ~new_C7164_;
  assign new_C7162_ = new_C7138_ & ~new_C7139_;
  assign new_C7163_ = ~new_C7185_ | ~new_C7186_;
  assign new_C7164_ = new_C7178_ | new_C7180_;
  assign new_C7165_ = new_C7188_ | new_C7187_;
  assign new_C7166_ = new_C7182_ | new_C7181_;
  assign new_C7167_ = ~new_C7190_ | ~new_C7189_;
  assign new_C7168_ = ~new_C7191_ & new_C7192_;
  assign new_C7169_ = new_C7191_ & ~new_C7192_;
  assign new_C7170_ = ~new_C7138_ & new_C7139_;
  assign new_C7171_ = new_C7138_ & ~new_C7139_;
  assign new_C7172_ = ~new_C7154_ | new_C7164_;
  assign new_C7173_ = new_C7154_ & new_C7164_;
  assign new_C7174_ = ~new_C7154_ & ~new_C7164_;
  assign new_C7175_ = new_C7196_ | new_C7195_;
  assign new_C7176_ = new_C7142_ | new_C7175_;
  assign new_C7177_ = new_C7200_ | new_C7199_;
  assign new_C7178_ = ~new_C7142_ & new_C7177_;
  assign new_C7179_ = new_C7198_ | new_C7197_;
  assign new_C7180_ = new_C7142_ & new_C7179_;
  assign new_C7181_ = new_C7140_ & ~new_C7150_;
  assign new_C7182_ = ~new_C7140_ & new_C7150_;
  assign new_C7183_ = ~new_C7139_ | ~new_C7164_;
  assign new_C7184_ = new_C7150_ & new_C7183_;
  assign new_C7185_ = ~new_C7150_ & ~new_C7184_;
  assign new_C7186_ = new_C7150_ | new_C7183_;
  assign new_C7187_ = ~new_C7140_ & new_C7141_;
  assign new_C7188_ = new_C7140_ & ~new_C7141_;
  assign new_C7189_ = new_C7157_ | new_C7194_;
  assign new_C7190_ = ~new_C7157_ & ~new_C7193_;
  assign new_C7191_ = new_C7140_ | new_C7157_;
  assign new_C7192_ = new_C7140_ | new_C7141_;
  assign new_C7193_ = new_C7157_ & new_C7194_;
  assign new_C7194_ = ~new_C7139_ | ~new_C7164_;
  assign new_C7195_ = new_C7172_ & new_C7192_;
  assign new_C7196_ = ~new_C7172_ & ~new_C7192_;
  assign new_C7197_ = new_C7201_ | new_C7202_;
  assign new_C7198_ = ~new_C7143_ & new_C7157_;
  assign new_C7199_ = new_C7203_ | new_C7204_;
  assign new_C7200_ = new_C7143_ & new_C7157_;
  assign new_C7201_ = ~new_C7143_ & ~new_C7157_;
  assign new_C7202_ = new_C7143_ & ~new_C7157_;
  assign new_C7203_ = new_C7143_ & ~new_C7157_;
  assign new_C7204_ = ~new_C7143_ & new_C7157_;
  assign new_C7205_ = new_F665_;
  assign new_C7206_ = new_F732_;
  assign new_C7207_ = new_F799_;
  assign new_C7208_ = new_F866_;
  assign new_C7209_ = new_F933_;
  assign new_C7210_ = new_F1000_;
  assign new_C7211_ = new_C7218_ & new_C7217_;
  assign new_C7212_ = new_C7220_ | new_C7219_;
  assign new_C7213_ = new_C7222_ | new_C7221_;
  assign new_C7214_ = new_C7224_ & new_C7223_;
  assign new_C7215_ = new_C7224_ & new_C7225_;
  assign new_C7216_ = new_C7217_ | new_C7226_;
  assign new_C7217_ = new_C7206_ | new_C7229_;
  assign new_C7218_ = new_C7228_ | new_C7227_;
  assign new_C7219_ = new_C7233_ & new_C7232_;
  assign new_C7220_ = new_C7231_ & new_C7230_;
  assign new_C7221_ = new_C7236_ | new_C7235_;
  assign new_C7222_ = new_C7231_ & new_C7234_;
  assign new_C7223_ = new_C7206_ | new_C7239_;
  assign new_C7224_ = new_C7238_ | new_C7237_;
  assign new_C7225_ = new_C7241_ | new_C7240_;
  assign new_C7226_ = ~new_C7217_ & new_C7243_;
  assign new_C7227_ = ~new_C7219_ & new_C7231_;
  assign new_C7228_ = new_C7219_ & ~new_C7231_;
  assign new_C7229_ = new_C7205_ & ~new_C7206_;
  assign new_C7230_ = ~new_C7252_ | ~new_C7253_;
  assign new_C7231_ = new_C7245_ | new_C7247_;
  assign new_C7232_ = new_C7255_ | new_C7254_;
  assign new_C7233_ = new_C7249_ | new_C7248_;
  assign new_C7234_ = ~new_C7257_ | ~new_C7256_;
  assign new_C7235_ = ~new_C7258_ & new_C7259_;
  assign new_C7236_ = new_C7258_ & ~new_C7259_;
  assign new_C7237_ = ~new_C7205_ & new_C7206_;
  assign new_C7238_ = new_C7205_ & ~new_C7206_;
  assign new_C7239_ = ~new_C7221_ | new_C7231_;
  assign new_C7240_ = new_C7221_ & new_C7231_;
  assign new_C7241_ = ~new_C7221_ & ~new_C7231_;
  assign new_C7242_ = new_C7263_ | new_C7262_;
  assign new_C7243_ = new_C7209_ | new_C7242_;
  assign new_C7244_ = new_C7267_ | new_C7266_;
  assign new_C7245_ = ~new_C7209_ & new_C7244_;
  assign new_C7246_ = new_C7265_ | new_C7264_;
  assign new_C7247_ = new_C7209_ & new_C7246_;
  assign new_C7248_ = new_C7207_ & ~new_C7217_;
  assign new_C7249_ = ~new_C7207_ & new_C7217_;
  assign new_C7250_ = ~new_C7206_ | ~new_C7231_;
  assign new_C7251_ = new_C7217_ & new_C7250_;
  assign new_C7252_ = ~new_C7217_ & ~new_C7251_;
  assign new_C7253_ = new_C7217_ | new_C7250_;
  assign new_C7254_ = ~new_C7207_ & new_C7208_;
  assign new_C7255_ = new_C7207_ & ~new_C7208_;
  assign new_C7256_ = new_C7224_ | new_C7261_;
  assign new_C7257_ = ~new_C7224_ & ~new_C7260_;
  assign new_C7258_ = new_C7207_ | new_C7224_;
  assign new_C7259_ = new_C7207_ | new_C7208_;
  assign new_C7260_ = new_C7224_ & new_C7261_;
  assign new_C7261_ = ~new_C7206_ | ~new_C7231_;
  assign new_C7262_ = new_C7239_ & new_C7259_;
  assign new_C7263_ = ~new_C7239_ & ~new_C7259_;
  assign new_C7264_ = new_C7268_ | new_C7269_;
  assign new_C7265_ = ~new_C7210_ & new_C7224_;
  assign new_C7266_ = new_C7270_ | new_C7271_;
  assign new_C7267_ = new_C7210_ & new_C7224_;
  assign new_C7268_ = ~new_C7210_ & ~new_C7224_;
  assign new_C7269_ = new_C7210_ & ~new_C7224_;
  assign new_C7270_ = new_C7210_ & ~new_C7224_;
  assign new_C7271_ = ~new_C7210_ & new_C7224_;
  assign new_C7272_ = new_F1067_;
  assign new_C7273_ = new_F1134_;
  assign new_C7274_ = new_F1201_;
  assign new_C7275_ = new_F1268_;
  assign new_C7276_ = new_F1335_;
  assign new_C7277_ = new_F1402_;
  assign new_C7278_ = new_C7285_ & new_C7284_;
  assign new_C7279_ = new_C7287_ | new_C7286_;
  assign new_C7280_ = new_C7289_ | new_C7288_;
  assign new_C7281_ = new_C7291_ & new_C7290_;
  assign new_C7282_ = new_C7291_ & new_C7292_;
  assign new_C7283_ = new_C7284_ | new_C7293_;
  assign new_C7284_ = new_C7273_ | new_C7296_;
  assign new_C7285_ = new_C7295_ | new_C7294_;
  assign new_C7286_ = new_C7300_ & new_C7299_;
  assign new_C7287_ = new_C7298_ & new_C7297_;
  assign new_C7288_ = new_C7303_ | new_C7302_;
  assign new_C7289_ = new_C7298_ & new_C7301_;
  assign new_C7290_ = new_C7273_ | new_C7306_;
  assign new_C7291_ = new_C7305_ | new_C7304_;
  assign new_C7292_ = new_C7308_ | new_C7307_;
  assign new_C7293_ = ~new_C7284_ & new_C7310_;
  assign new_C7294_ = ~new_C7286_ & new_C7298_;
  assign new_C7295_ = new_C7286_ & ~new_C7298_;
  assign new_C7296_ = new_C7272_ & ~new_C7273_;
  assign new_C7297_ = ~new_C7319_ | ~new_C7320_;
  assign new_C7298_ = new_C7312_ | new_C7314_;
  assign new_C7299_ = new_C7322_ | new_C7321_;
  assign new_C7300_ = new_C7316_ | new_C7315_;
  assign new_C7301_ = ~new_C7324_ | ~new_C7323_;
  assign new_C7302_ = ~new_C7325_ & new_C7326_;
  assign new_C7303_ = new_C7325_ & ~new_C7326_;
  assign new_C7304_ = ~new_C7272_ & new_C7273_;
  assign new_C7305_ = new_C7272_ & ~new_C7273_;
  assign new_C7306_ = ~new_C7288_ | new_C7298_;
  assign new_C7307_ = new_C7288_ & new_C7298_;
  assign new_C7308_ = ~new_C7288_ & ~new_C7298_;
  assign new_C7309_ = new_C7330_ | new_C7329_;
  assign new_C7310_ = new_C7276_ | new_C7309_;
  assign new_C7311_ = new_C7334_ | new_C7333_;
  assign new_C7312_ = ~new_C7276_ & new_C7311_;
  assign new_C7313_ = new_C7332_ | new_C7331_;
  assign new_C7314_ = new_C7276_ & new_C7313_;
  assign new_C7315_ = new_C7274_ & ~new_C7284_;
  assign new_C7316_ = ~new_C7274_ & new_C7284_;
  assign new_C7317_ = ~new_C7273_ | ~new_C7298_;
  assign new_C7318_ = new_C7284_ & new_C7317_;
  assign new_C7319_ = ~new_C7284_ & ~new_C7318_;
  assign new_C7320_ = new_C7284_ | new_C7317_;
  assign new_C7321_ = ~new_C7274_ & new_C7275_;
  assign new_C7322_ = new_C7274_ & ~new_C7275_;
  assign new_C7323_ = new_C7291_ | new_C7328_;
  assign new_C7324_ = ~new_C7291_ & ~new_C7327_;
  assign new_C7325_ = new_C7274_ | new_C7291_;
  assign new_C7326_ = new_C7274_ | new_C7275_;
  assign new_C7327_ = new_C7291_ & new_C7328_;
  assign new_C7328_ = ~new_C7273_ | ~new_C7298_;
  assign new_C7329_ = new_C7306_ & new_C7326_;
  assign new_C7330_ = ~new_C7306_ & ~new_C7326_;
  assign new_C7331_ = new_C7335_ | new_C7336_;
  assign new_C7332_ = ~new_C7277_ & new_C7291_;
  assign new_C7333_ = new_C7337_ | new_C7338_;
  assign new_C7334_ = new_C7277_ & new_C7291_;
  assign new_C7335_ = ~new_C7277_ & ~new_C7291_;
  assign new_C7336_ = new_C7277_ & ~new_C7291_;
  assign new_C7337_ = new_C7277_ & ~new_C7291_;
  assign new_C7338_ = ~new_C7277_ & new_C7291_;
  assign new_C7339_ = new_D6997_;
  assign new_C7340_ = new_D7063_;
  assign new_C7341_ = new_D7130_;
  assign new_C7342_ = new_D7197_;
  assign new_C7343_ = new_D7264_;
  assign new_C7344_ = new_D7331_;
  assign new_C7345_ = new_C7352_ & new_C7351_;
  assign new_C7346_ = new_C7354_ | new_C7353_;
  assign new_C7347_ = new_C7356_ | new_C7355_;
  assign new_C7348_ = new_C7358_ & new_C7357_;
  assign new_C7349_ = new_C7358_ & new_C7359_;
  assign new_C7350_ = new_C7351_ | new_C7360_;
  assign new_C7351_ = new_C7340_ | new_C7363_;
  assign new_C7352_ = new_C7362_ | new_C7361_;
  assign new_C7353_ = new_C7367_ & new_C7366_;
  assign new_C7354_ = new_C7365_ & new_C7364_;
  assign new_C7355_ = new_C7370_ | new_C7369_;
  assign new_C7356_ = new_C7365_ & new_C7368_;
  assign new_C7357_ = new_C7340_ | new_C7373_;
  assign new_C7358_ = new_C7372_ | new_C7371_;
  assign new_C7359_ = new_C7375_ | new_C7374_;
  assign new_C7360_ = ~new_C7351_ & new_C7377_;
  assign new_C7361_ = ~new_C7353_ & new_C7365_;
  assign new_C7362_ = new_C7353_ & ~new_C7365_;
  assign new_C7363_ = new_C7339_ & ~new_C7340_;
  assign new_C7364_ = ~new_C7386_ | ~new_C7387_;
  assign new_C7365_ = new_C7379_ | new_C7381_;
  assign new_C7366_ = new_C7389_ | new_C7388_;
  assign new_C7367_ = new_C7383_ | new_C7382_;
  assign new_C7368_ = ~new_C7391_ | ~new_C7390_;
  assign new_C7369_ = ~new_C7392_ & new_C7393_;
  assign new_C7370_ = new_C7392_ & ~new_C7393_;
  assign new_C7371_ = ~new_C7339_ & new_C7340_;
  assign new_C7372_ = new_C7339_ & ~new_C7340_;
  assign new_C7373_ = ~new_C7355_ | new_C7365_;
  assign new_C7374_ = new_C7355_ & new_C7365_;
  assign new_C7375_ = ~new_C7355_ & ~new_C7365_;
  assign new_C7376_ = new_C7397_ | new_C7396_;
  assign new_C7377_ = new_C7343_ | new_C7376_;
  assign new_C7378_ = new_C7401_ | new_C7400_;
  assign new_C7379_ = ~new_C7343_ & new_C7378_;
  assign new_C7380_ = new_C7399_ | new_C7398_;
  assign new_C7381_ = new_C7343_ & new_C7380_;
  assign new_C7382_ = new_C7341_ & ~new_C7351_;
  assign new_C7383_ = ~new_C7341_ & new_C7351_;
  assign new_C7384_ = ~new_C7340_ | ~new_C7365_;
  assign new_C7385_ = new_C7351_ & new_C7384_;
  assign new_C7386_ = ~new_C7351_ & ~new_C7385_;
  assign new_C7387_ = new_C7351_ | new_C7384_;
  assign new_C7388_ = ~new_C7341_ & new_C7342_;
  assign new_C7389_ = new_C7341_ & ~new_C7342_;
  assign new_C7390_ = new_C7358_ | new_C7395_;
  assign new_C7391_ = ~new_C7358_ & ~new_C7394_;
  assign new_C7392_ = new_C7341_ | new_C7358_;
  assign new_C7393_ = new_C7341_ | new_C7342_;
  assign new_C7394_ = new_C7358_ & new_C7395_;
  assign new_C7395_ = ~new_C7340_ | ~new_C7365_;
  assign new_C7396_ = new_C7373_ & new_C7393_;
  assign new_C7397_ = ~new_C7373_ & ~new_C7393_;
  assign new_C7398_ = new_C7402_ | new_C7403_;
  assign new_C7399_ = ~new_C7344_ & new_C7358_;
  assign new_C7400_ = new_C7404_ | new_C7405_;
  assign new_C7401_ = new_C7344_ & new_C7358_;
  assign new_C7402_ = ~new_C7344_ & ~new_C7358_;
  assign new_C7403_ = new_C7344_ & ~new_C7358_;
  assign new_C7404_ = new_C7344_ & ~new_C7358_;
  assign new_C7405_ = ~new_C7344_ & new_C7358_;
  assign new_C7406_ = new_D7398_;
  assign new_C7407_ = new_D7465_;
  assign new_C7408_ = new_D7532_;
  assign new_C7409_ = new_D7599_;
  assign new_C7410_ = new_D7666_;
  assign new_C7411_ = new_D7733_;
  assign new_C7412_ = new_C7419_ & new_C7418_;
  assign new_C7413_ = new_C7421_ | new_C7420_;
  assign new_C7414_ = new_C7423_ | new_C7422_;
  assign new_C7415_ = new_C7425_ & new_C7424_;
  assign new_C7416_ = new_C7425_ & new_C7426_;
  assign new_C7417_ = new_C7418_ | new_C7427_;
  assign new_C7418_ = new_C7407_ | new_C7430_;
  assign new_C7419_ = new_C7429_ | new_C7428_;
  assign new_C7420_ = new_C7434_ & new_C7433_;
  assign new_C7421_ = new_C7432_ & new_C7431_;
  assign new_C7422_ = new_C7437_ | new_C7436_;
  assign new_C7423_ = new_C7432_ & new_C7435_;
  assign new_C7424_ = new_C7407_ | new_C7440_;
  assign new_C7425_ = new_C7439_ | new_C7438_;
  assign new_C7426_ = new_C7442_ | new_C7441_;
  assign new_C7427_ = ~new_C7418_ & new_C7444_;
  assign new_C7428_ = ~new_C7420_ & new_C7432_;
  assign new_C7429_ = new_C7420_ & ~new_C7432_;
  assign new_C7430_ = new_C7406_ & ~new_C7407_;
  assign new_C7431_ = ~new_C7453_ | ~new_C7454_;
  assign new_C7432_ = new_C7446_ | new_C7448_;
  assign new_C7433_ = new_C7456_ | new_C7455_;
  assign new_C7434_ = new_C7450_ | new_C7449_;
  assign new_C7435_ = ~new_C7458_ | ~new_C7457_;
  assign new_C7436_ = ~new_C7459_ & new_C7460_;
  assign new_C7437_ = new_C7459_ & ~new_C7460_;
  assign new_C7438_ = ~new_C7406_ & new_C7407_;
  assign new_C7439_ = new_C7406_ & ~new_C7407_;
  assign new_C7440_ = ~new_C7422_ | new_C7432_;
  assign new_C7441_ = new_C7422_ & new_C7432_;
  assign new_C7442_ = ~new_C7422_ & ~new_C7432_;
  assign new_C7443_ = new_C7464_ | new_C7463_;
  assign new_C7444_ = new_C7410_ | new_C7443_;
  assign new_C7445_ = new_C7468_ | new_C7467_;
  assign new_C7446_ = ~new_C7410_ & new_C7445_;
  assign new_C7447_ = new_C7466_ | new_C7465_;
  assign new_C7448_ = new_C7410_ & new_C7447_;
  assign new_C7449_ = new_C7408_ & ~new_C7418_;
  assign new_C7450_ = ~new_C7408_ & new_C7418_;
  assign new_C7451_ = ~new_C7407_ | ~new_C7432_;
  assign new_C7452_ = new_C7418_ & new_C7451_;
  assign new_C7453_ = ~new_C7418_ & ~new_C7452_;
  assign new_C7454_ = new_C7418_ | new_C7451_;
  assign new_C7455_ = ~new_C7408_ & new_C7409_;
  assign new_C7456_ = new_C7408_ & ~new_C7409_;
  assign new_C7457_ = new_C7425_ | new_C7462_;
  assign new_C7458_ = ~new_C7425_ & ~new_C7461_;
  assign new_C7459_ = new_C7408_ | new_C7425_;
  assign new_C7460_ = new_C7408_ | new_C7409_;
  assign new_C7461_ = new_C7425_ & new_C7462_;
  assign new_C7462_ = ~new_C7407_ | ~new_C7432_;
  assign new_C7463_ = new_C7440_ & new_C7460_;
  assign new_C7464_ = ~new_C7440_ & ~new_C7460_;
  assign new_C7465_ = new_C7469_ | new_C7470_;
  assign new_C7466_ = ~new_C7411_ & new_C7425_;
  assign new_C7467_ = new_C7471_ | new_C7472_;
  assign new_C7468_ = new_C7411_ & new_C7425_;
  assign new_C7469_ = ~new_C7411_ & ~new_C7425_;
  assign new_C7470_ = new_C7411_ & ~new_C7425_;
  assign new_C7471_ = new_C7411_ & ~new_C7425_;
  assign new_C7472_ = ~new_C7411_ & new_C7425_;
  assign new_C7473_ = new_D7800_;
  assign new_C7474_ = new_D7867_;
  assign new_C7475_ = new_D7934_;
  assign new_C7476_ = new_D8001_;
  assign new_C7477_ = new_D8068_;
  assign new_C7478_ = new_D8135_;
  assign new_C7479_ = new_C7486_ & new_C7485_;
  assign new_C7480_ = new_C7488_ | new_C7487_;
  assign new_C7481_ = new_C7490_ | new_C7489_;
  assign new_C7482_ = new_C7492_ & new_C7491_;
  assign new_C7483_ = new_C7492_ & new_C7493_;
  assign new_C7484_ = new_C7485_ | new_C7494_;
  assign new_C7485_ = new_C7474_ | new_C7497_;
  assign new_C7486_ = new_C7496_ | new_C7495_;
  assign new_C7487_ = new_C7501_ & new_C7500_;
  assign new_C7488_ = new_C7499_ & new_C7498_;
  assign new_C7489_ = new_C7504_ | new_C7503_;
  assign new_C7490_ = new_C7499_ & new_C7502_;
  assign new_C7491_ = new_C7474_ | new_C7507_;
  assign new_C7492_ = new_C7506_ | new_C7505_;
  assign new_C7493_ = new_C7509_ | new_C7508_;
  assign new_C7494_ = ~new_C7485_ & new_C7511_;
  assign new_C7495_ = ~new_C7487_ & new_C7499_;
  assign new_C7496_ = new_C7487_ & ~new_C7499_;
  assign new_C7497_ = new_C7473_ & ~new_C7474_;
  assign new_C7498_ = ~new_C7520_ | ~new_C7521_;
  assign new_C7499_ = new_C7513_ | new_C7515_;
  assign new_C7500_ = new_C7523_ | new_C7522_;
  assign new_C7501_ = new_C7517_ | new_C7516_;
  assign new_C7502_ = ~new_C7525_ | ~new_C7524_;
  assign new_C7503_ = ~new_C7526_ & new_C7527_;
  assign new_C7504_ = new_C7526_ & ~new_C7527_;
  assign new_C7505_ = ~new_C7473_ & new_C7474_;
  assign new_C7506_ = new_C7473_ & ~new_C7474_;
  assign new_C7507_ = ~new_C7489_ | new_C7499_;
  assign new_C7508_ = new_C7489_ & new_C7499_;
  assign new_C7509_ = ~new_C7489_ & ~new_C7499_;
  assign new_C7510_ = new_C7531_ | new_C7530_;
  assign new_C7511_ = new_C7477_ | new_C7510_;
  assign new_C7512_ = new_C7535_ | new_C7534_;
  assign new_C7513_ = ~new_C7477_ & new_C7512_;
  assign new_C7514_ = new_C7533_ | new_C7532_;
  assign new_C7515_ = new_C7477_ & new_C7514_;
  assign new_C7516_ = new_C7475_ & ~new_C7485_;
  assign new_C7517_ = ~new_C7475_ & new_C7485_;
  assign new_C7518_ = ~new_C7474_ | ~new_C7499_;
  assign new_C7519_ = new_C7485_ & new_C7518_;
  assign new_C7520_ = ~new_C7485_ & ~new_C7519_;
  assign new_C7521_ = new_C7485_ | new_C7518_;
  assign new_C7522_ = ~new_C7475_ & new_C7476_;
  assign new_C7523_ = new_C7475_ & ~new_C7476_;
  assign new_C7524_ = new_C7492_ | new_C7529_;
  assign new_C7525_ = ~new_C7492_ & ~new_C7528_;
  assign new_C7526_ = new_C7475_ | new_C7492_;
  assign new_C7527_ = new_C7475_ | new_C7476_;
  assign new_C7528_ = new_C7492_ & new_C7529_;
  assign new_C7529_ = ~new_C7474_ | ~new_C7499_;
  assign new_C7530_ = new_C7507_ & new_C7527_;
  assign new_C7531_ = ~new_C7507_ & ~new_C7527_;
  assign new_C7532_ = new_C7536_ | new_C7537_;
  assign new_C7533_ = ~new_C7478_ & new_C7492_;
  assign new_C7534_ = new_C7538_ | new_C7539_;
  assign new_C7535_ = new_C7478_ & new_C7492_;
  assign new_C7536_ = ~new_C7478_ & ~new_C7492_;
  assign new_C7537_ = new_C7478_ & ~new_C7492_;
  assign new_C7538_ = new_C7478_ & ~new_C7492_;
  assign new_C7539_ = ~new_C7478_ & new_C7492_;
  assign new_C7540_ = new_D8202_;
  assign new_C7541_ = new_D8269_;
  assign new_C7542_ = new_D8336_;
  assign new_C7543_ = new_D8403_;
  assign new_C7544_ = new_D8470_;
  assign new_C7545_ = new_D8537_;
  assign new_C7546_ = new_C7553_ & new_C7552_;
  assign new_C7547_ = new_C7555_ | new_C7554_;
  assign new_C7548_ = new_C7557_ | new_C7556_;
  assign new_C7549_ = new_C7559_ & new_C7558_;
  assign new_C7550_ = new_C7559_ & new_C7560_;
  assign new_C7551_ = new_C7552_ | new_C7561_;
  assign new_C7552_ = new_C7541_ | new_C7564_;
  assign new_C7553_ = new_C7563_ | new_C7562_;
  assign new_C7554_ = new_C7568_ & new_C7567_;
  assign new_C7555_ = new_C7566_ & new_C7565_;
  assign new_C7556_ = new_C7571_ | new_C7570_;
  assign new_C7557_ = new_C7566_ & new_C7569_;
  assign new_C7558_ = new_C7541_ | new_C7574_;
  assign new_C7559_ = new_C7573_ | new_C7572_;
  assign new_C7560_ = new_C7576_ | new_C7575_;
  assign new_C7561_ = ~new_C7552_ & new_C7578_;
  assign new_C7562_ = ~new_C7554_ & new_C7566_;
  assign new_C7563_ = new_C7554_ & ~new_C7566_;
  assign new_C7564_ = new_C7540_ & ~new_C7541_;
  assign new_C7565_ = ~new_C7587_ | ~new_C7588_;
  assign new_C7566_ = new_C7580_ | new_C7582_;
  assign new_C7567_ = new_C7590_ | new_C7589_;
  assign new_C7568_ = new_C7584_ | new_C7583_;
  assign new_C7569_ = ~new_C7592_ | ~new_C7591_;
  assign new_C7570_ = ~new_C7593_ & new_C7594_;
  assign new_C7571_ = new_C7593_ & ~new_C7594_;
  assign new_C7572_ = ~new_C7540_ & new_C7541_;
  assign new_C7573_ = new_C7540_ & ~new_C7541_;
  assign new_C7574_ = ~new_C7556_ | new_C7566_;
  assign new_C7575_ = new_C7556_ & new_C7566_;
  assign new_C7576_ = ~new_C7556_ & ~new_C7566_;
  assign new_C7577_ = new_C7598_ | new_C7597_;
  assign new_C7578_ = new_C7544_ | new_C7577_;
  assign new_C7579_ = new_C7602_ | new_C7601_;
  assign new_C7580_ = ~new_C7544_ & new_C7579_;
  assign new_C7581_ = new_C7600_ | new_C7599_;
  assign new_C7582_ = new_C7544_ & new_C7581_;
  assign new_C7583_ = new_C7542_ & ~new_C7552_;
  assign new_C7584_ = ~new_C7542_ & new_C7552_;
  assign new_C7585_ = ~new_C7541_ | ~new_C7566_;
  assign new_C7586_ = new_C7552_ & new_C7585_;
  assign new_C7587_ = ~new_C7552_ & ~new_C7586_;
  assign new_C7588_ = new_C7552_ | new_C7585_;
  assign new_C7589_ = ~new_C7542_ & new_C7543_;
  assign new_C7590_ = new_C7542_ & ~new_C7543_;
  assign new_C7591_ = new_C7559_ | new_C7596_;
  assign new_C7592_ = ~new_C7559_ & ~new_C7595_;
  assign new_C7593_ = new_C7542_ | new_C7559_;
  assign new_C7594_ = new_C7542_ | new_C7543_;
  assign new_C7595_ = new_C7559_ & new_C7596_;
  assign new_C7596_ = ~new_C7541_ | ~new_C7566_;
  assign new_C7597_ = new_C7574_ & new_C7594_;
  assign new_C7598_ = ~new_C7574_ & ~new_C7594_;
  assign new_C7599_ = new_C7603_ | new_C7604_;
  assign new_C7600_ = ~new_C7545_ & new_C7559_;
  assign new_C7601_ = new_C7605_ | new_C7606_;
  assign new_C7602_ = new_C7545_ & new_C7559_;
  assign new_C7603_ = ~new_C7545_ & ~new_C7559_;
  assign new_C7604_ = new_C7545_ & ~new_C7559_;
  assign new_C7605_ = new_C7545_ & ~new_C7559_;
  assign new_C7606_ = ~new_C7545_ & new_C7559_;
  assign new_C7607_ = new_D8604_;
  assign new_C7608_ = new_D8671_;
  assign new_C7609_ = new_D8738_;
  assign new_C7610_ = new_D8805_;
  assign new_C7611_ = new_D8872_;
  assign new_C7612_ = new_D8939_;
  assign new_C7613_ = new_C7620_ & new_C7619_;
  assign new_C7614_ = new_C7622_ | new_C7621_;
  assign new_C7615_ = new_C7624_ | new_C7623_;
  assign new_C7616_ = new_C7626_ & new_C7625_;
  assign new_C7617_ = new_C7626_ & new_C7627_;
  assign new_C7618_ = new_C7619_ | new_C7628_;
  assign new_C7619_ = new_C7608_ | new_C7631_;
  assign new_C7620_ = new_C7630_ | new_C7629_;
  assign new_C7621_ = new_C7635_ & new_C7634_;
  assign new_C7622_ = new_C7633_ & new_C7632_;
  assign new_C7623_ = new_C7638_ | new_C7637_;
  assign new_C7624_ = new_C7633_ & new_C7636_;
  assign new_C7625_ = new_C7608_ | new_C7641_;
  assign new_C7626_ = new_C7640_ | new_C7639_;
  assign new_C7627_ = new_C7643_ | new_C7642_;
  assign new_C7628_ = ~new_C7619_ & new_C7645_;
  assign new_C7629_ = ~new_C7621_ & new_C7633_;
  assign new_C7630_ = new_C7621_ & ~new_C7633_;
  assign new_C7631_ = new_C7607_ & ~new_C7608_;
  assign new_C7632_ = ~new_C7654_ | ~new_C7655_;
  assign new_C7633_ = new_C7647_ | new_C7649_;
  assign new_C7634_ = new_C7657_ | new_C7656_;
  assign new_C7635_ = new_C7651_ | new_C7650_;
  assign new_C7636_ = ~new_C7659_ | ~new_C7658_;
  assign new_C7637_ = ~new_C7660_ & new_C7661_;
  assign new_C7638_ = new_C7660_ & ~new_C7661_;
  assign new_C7639_ = ~new_C7607_ & new_C7608_;
  assign new_C7640_ = new_C7607_ & ~new_C7608_;
  assign new_C7641_ = ~new_C7623_ | new_C7633_;
  assign new_C7642_ = new_C7623_ & new_C7633_;
  assign new_C7643_ = ~new_C7623_ & ~new_C7633_;
  assign new_C7644_ = new_C7665_ | new_C7664_;
  assign new_C7645_ = new_C7611_ | new_C7644_;
  assign new_C7646_ = new_C7669_ | new_C7668_;
  assign new_C7647_ = ~new_C7611_ & new_C7646_;
  assign new_C7648_ = new_C7667_ | new_C7666_;
  assign new_C7649_ = new_C7611_ & new_C7648_;
  assign new_C7650_ = new_C7609_ & ~new_C7619_;
  assign new_C7651_ = ~new_C7609_ & new_C7619_;
  assign new_C7652_ = ~new_C7608_ | ~new_C7633_;
  assign new_C7653_ = new_C7619_ & new_C7652_;
  assign new_C7654_ = ~new_C7619_ & ~new_C7653_;
  assign new_C7655_ = new_C7619_ | new_C7652_;
  assign new_C7656_ = ~new_C7609_ & new_C7610_;
  assign new_C7657_ = new_C7609_ & ~new_C7610_;
  assign new_C7658_ = new_C7626_ | new_C7663_;
  assign new_C7659_ = ~new_C7626_ & ~new_C7662_;
  assign new_C7660_ = new_C7609_ | new_C7626_;
  assign new_C7661_ = new_C7609_ | new_C7610_;
  assign new_C7662_ = new_C7626_ & new_C7663_;
  assign new_C7663_ = ~new_C7608_ | ~new_C7633_;
  assign new_C7664_ = new_C7641_ & new_C7661_;
  assign new_C7665_ = ~new_C7641_ & ~new_C7661_;
  assign new_C7666_ = new_C7670_ | new_C7671_;
  assign new_C7667_ = ~new_C7612_ & new_C7626_;
  assign new_C7668_ = new_C7672_ | new_C7673_;
  assign new_C7669_ = new_C7612_ & new_C7626_;
  assign new_C7670_ = ~new_C7612_ & ~new_C7626_;
  assign new_C7671_ = new_C7612_ & ~new_C7626_;
  assign new_C7672_ = new_C7612_ & ~new_C7626_;
  assign new_C7673_ = ~new_C7612_ & new_C7626_;
  assign new_C7674_ = new_D9006_;
  assign new_C7675_ = new_D9073_;
  assign new_C7676_ = new_D9140_;
  assign new_C7677_ = new_D9207_;
  assign new_C7678_ = new_D9274_;
  assign new_C7679_ = new_D9341_;
  assign new_C7680_ = new_C7687_ & new_C7686_;
  assign new_C7681_ = new_C7689_ | new_C7688_;
  assign new_C7682_ = new_C7691_ | new_C7690_;
  assign new_C7683_ = new_C7693_ & new_C7692_;
  assign new_C7684_ = new_C7693_ & new_C7694_;
  assign new_C7685_ = new_C7686_ | new_C7695_;
  assign new_C7686_ = new_C7675_ | new_C7698_;
  assign new_C7687_ = new_C7697_ | new_C7696_;
  assign new_C7688_ = new_C7702_ & new_C7701_;
  assign new_C7689_ = new_C7700_ & new_C7699_;
  assign new_C7690_ = new_C7705_ | new_C7704_;
  assign new_C7691_ = new_C7700_ & new_C7703_;
  assign new_C7692_ = new_C7675_ | new_C7708_;
  assign new_C7693_ = new_C7707_ | new_C7706_;
  assign new_C7694_ = new_C7710_ | new_C7709_;
  assign new_C7695_ = ~new_C7686_ & new_C7712_;
  assign new_C7696_ = ~new_C7688_ & new_C7700_;
  assign new_C7697_ = new_C7688_ & ~new_C7700_;
  assign new_C7698_ = new_C7674_ & ~new_C7675_;
  assign new_C7699_ = ~new_C7721_ | ~new_C7722_;
  assign new_C7700_ = new_C7714_ | new_C7716_;
  assign new_C7701_ = new_C7724_ | new_C7723_;
  assign new_C7702_ = new_C7718_ | new_C7717_;
  assign new_C7703_ = ~new_C7726_ | ~new_C7725_;
  assign new_C7704_ = ~new_C7727_ & new_C7728_;
  assign new_C7705_ = new_C7727_ & ~new_C7728_;
  assign new_C7706_ = ~new_C7674_ & new_C7675_;
  assign new_C7707_ = new_C7674_ & ~new_C7675_;
  assign new_C7708_ = ~new_C7690_ | new_C7700_;
  assign new_C7709_ = new_C7690_ & new_C7700_;
  assign new_C7710_ = ~new_C7690_ & ~new_C7700_;
  assign new_C7711_ = new_C7732_ | new_C7731_;
  assign new_C7712_ = new_C7678_ | new_C7711_;
  assign new_C7713_ = new_C7736_ | new_C7735_;
  assign new_C7714_ = ~new_C7678_ & new_C7713_;
  assign new_C7715_ = new_C7734_ | new_C7733_;
  assign new_C7716_ = new_C7678_ & new_C7715_;
  assign new_C7717_ = new_C7676_ & ~new_C7686_;
  assign new_C7718_ = ~new_C7676_ & new_C7686_;
  assign new_C7719_ = ~new_C7675_ | ~new_C7700_;
  assign new_C7720_ = new_C7686_ & new_C7719_;
  assign new_C7721_ = ~new_C7686_ & ~new_C7720_;
  assign new_C7722_ = new_C7686_ | new_C7719_;
  assign new_C7723_ = ~new_C7676_ & new_C7677_;
  assign new_C7724_ = new_C7676_ & ~new_C7677_;
  assign new_C7725_ = new_C7693_ | new_C7730_;
  assign new_C7726_ = ~new_C7693_ & ~new_C7729_;
  assign new_C7727_ = new_C7676_ | new_C7693_;
  assign new_C7728_ = new_C7676_ | new_C7677_;
  assign new_C7729_ = new_C7693_ & new_C7730_;
  assign new_C7730_ = ~new_C7675_ | ~new_C7700_;
  assign new_C7731_ = new_C7708_ & new_C7728_;
  assign new_C7732_ = ~new_C7708_ & ~new_C7728_;
  assign new_C7733_ = new_C7737_ | new_C7738_;
  assign new_C7734_ = ~new_C7679_ & new_C7693_;
  assign new_C7735_ = new_C7739_ | new_C7740_;
  assign new_C7736_ = new_C7679_ & new_C7693_;
  assign new_C7737_ = ~new_C7679_ & ~new_C7693_;
  assign new_C7738_ = new_C7679_ & ~new_C7693_;
  assign new_C7739_ = new_C7679_ & ~new_C7693_;
  assign new_C7740_ = ~new_C7679_ & new_C7693_;
  assign new_C7741_ = new_D9408_;
  assign new_C7742_ = new_D9475_;
  assign new_C7743_ = new_D9542_;
  assign new_C7744_ = new_D9609_;
  assign new_C7745_ = new_D9676_;
  assign new_C7746_ = new_D9743_;
  assign new_C7747_ = new_C7754_ & new_C7753_;
  assign new_C7748_ = new_C7756_ | new_C7755_;
  assign new_C7749_ = new_C7758_ | new_C7757_;
  assign new_C7750_ = new_C7760_ & new_C7759_;
  assign new_C7751_ = new_C7760_ & new_C7761_;
  assign new_C7752_ = new_C7753_ | new_C7762_;
  assign new_C7753_ = new_C7742_ | new_C7765_;
  assign new_C7754_ = new_C7764_ | new_C7763_;
  assign new_C7755_ = new_C7769_ & new_C7768_;
  assign new_C7756_ = new_C7767_ & new_C7766_;
  assign new_C7757_ = new_C7772_ | new_C7771_;
  assign new_C7758_ = new_C7767_ & new_C7770_;
  assign new_C7759_ = new_C7742_ | new_C7775_;
  assign new_C7760_ = new_C7774_ | new_C7773_;
  assign new_C7761_ = new_C7777_ | new_C7776_;
  assign new_C7762_ = ~new_C7753_ & new_C7779_;
  assign new_C7763_ = ~new_C7755_ & new_C7767_;
  assign new_C7764_ = new_C7755_ & ~new_C7767_;
  assign new_C7765_ = new_C7741_ & ~new_C7742_;
  assign new_C7766_ = ~new_C7788_ | ~new_C7789_;
  assign new_C7767_ = new_C7781_ | new_C7783_;
  assign new_C7768_ = new_C7791_ | new_C7790_;
  assign new_C7769_ = new_C7785_ | new_C7784_;
  assign new_C7770_ = ~new_C7793_ | ~new_C7792_;
  assign new_C7771_ = ~new_C7794_ & new_C7795_;
  assign new_C7772_ = new_C7794_ & ~new_C7795_;
  assign new_C7773_ = ~new_C7741_ & new_C7742_;
  assign new_C7774_ = new_C7741_ & ~new_C7742_;
  assign new_C7775_ = ~new_C7757_ | new_C7767_;
  assign new_C7776_ = new_C7757_ & new_C7767_;
  assign new_C7777_ = ~new_C7757_ & ~new_C7767_;
  assign new_C7778_ = new_C7799_ | new_C7798_;
  assign new_C7779_ = new_C7745_ | new_C7778_;
  assign new_C7780_ = new_C7803_ | new_C7802_;
  assign new_C7781_ = ~new_C7745_ & new_C7780_;
  assign new_C7782_ = new_C7801_ | new_C7800_;
  assign new_C7783_ = new_C7745_ & new_C7782_;
  assign new_C7784_ = new_C7743_ & ~new_C7753_;
  assign new_C7785_ = ~new_C7743_ & new_C7753_;
  assign new_C7786_ = ~new_C7742_ | ~new_C7767_;
  assign new_C7787_ = new_C7753_ & new_C7786_;
  assign new_C7788_ = ~new_C7753_ & ~new_C7787_;
  assign new_C7789_ = new_C7753_ | new_C7786_;
  assign new_C7790_ = ~new_C7743_ & new_C7744_;
  assign new_C7791_ = new_C7743_ & ~new_C7744_;
  assign new_C7792_ = new_C7760_ | new_C7797_;
  assign new_C7793_ = ~new_C7760_ & ~new_C7796_;
  assign new_C7794_ = new_C7743_ | new_C7760_;
  assign new_C7795_ = new_C7743_ | new_C7744_;
  assign new_C7796_ = new_C7760_ & new_C7797_;
  assign new_C7797_ = ~new_C7742_ | ~new_C7767_;
  assign new_C7798_ = new_C7775_ & new_C7795_;
  assign new_C7799_ = ~new_C7775_ & ~new_C7795_;
  assign new_C7800_ = new_C7804_ | new_C7805_;
  assign new_C7801_ = ~new_C7746_ & new_C7760_;
  assign new_C7802_ = new_C7806_ | new_C7807_;
  assign new_C7803_ = new_C7746_ & new_C7760_;
  assign new_C7804_ = ~new_C7746_ & ~new_C7760_;
  assign new_C7805_ = new_C7746_ & ~new_C7760_;
  assign new_C7806_ = new_C7746_ & ~new_C7760_;
  assign new_C7807_ = ~new_C7746_ & new_C7760_;
  assign new_C7808_ = new_D9810_;
  assign new_C7809_ = new_D9877_;
  assign new_C7810_ = new_D9944_;
  assign new_C7811_ = new_E12_;
  assign new_C7812_ = new_E79_;
  assign new_C7813_ = new_E146_;
  assign new_C7814_ = new_C7821_ & new_C7820_;
  assign new_C7815_ = new_C7823_ | new_C7822_;
  assign new_C7816_ = new_C7825_ | new_C7824_;
  assign new_C7817_ = new_C7827_ & new_C7826_;
  assign new_C7818_ = new_C7827_ & new_C7828_;
  assign new_C7819_ = new_C7820_ | new_C7829_;
  assign new_C7820_ = new_C7809_ | new_C7832_;
  assign new_C7821_ = new_C7831_ | new_C7830_;
  assign new_C7822_ = new_C7836_ & new_C7835_;
  assign new_C7823_ = new_C7834_ & new_C7833_;
  assign new_C7824_ = new_C7839_ | new_C7838_;
  assign new_C7825_ = new_C7834_ & new_C7837_;
  assign new_C7826_ = new_C7809_ | new_C7842_;
  assign new_C7827_ = new_C7841_ | new_C7840_;
  assign new_C7828_ = new_C7844_ | new_C7843_;
  assign new_C7829_ = ~new_C7820_ & new_C7846_;
  assign new_C7830_ = ~new_C7822_ & new_C7834_;
  assign new_C7831_ = new_C7822_ & ~new_C7834_;
  assign new_C7832_ = new_C7808_ & ~new_C7809_;
  assign new_C7833_ = ~new_C7855_ | ~new_C7856_;
  assign new_C7834_ = new_C7848_ | new_C7850_;
  assign new_C7835_ = new_C7858_ | new_C7857_;
  assign new_C7836_ = new_C7852_ | new_C7851_;
  assign new_C7837_ = ~new_C7860_ | ~new_C7859_;
  assign new_C7838_ = ~new_C7861_ & new_C7862_;
  assign new_C7839_ = new_C7861_ & ~new_C7862_;
  assign new_C7840_ = ~new_C7808_ & new_C7809_;
  assign new_C7841_ = new_C7808_ & ~new_C7809_;
  assign new_C7842_ = ~new_C7824_ | new_C7834_;
  assign new_C7843_ = new_C7824_ & new_C7834_;
  assign new_C7844_ = ~new_C7824_ & ~new_C7834_;
  assign new_C7845_ = new_C7866_ | new_C7865_;
  assign new_C7846_ = new_C7812_ | new_C7845_;
  assign new_C7847_ = new_C7870_ | new_C7869_;
  assign new_C7848_ = ~new_C7812_ & new_C7847_;
  assign new_C7849_ = new_C7868_ | new_C7867_;
  assign new_C7850_ = new_C7812_ & new_C7849_;
  assign new_C7851_ = new_C7810_ & ~new_C7820_;
  assign new_C7852_ = ~new_C7810_ & new_C7820_;
  assign new_C7853_ = ~new_C7809_ | ~new_C7834_;
  assign new_C7854_ = new_C7820_ & new_C7853_;
  assign new_C7855_ = ~new_C7820_ & ~new_C7854_;
  assign new_C7856_ = new_C7820_ | new_C7853_;
  assign new_C7857_ = ~new_C7810_ & new_C7811_;
  assign new_C7858_ = new_C7810_ & ~new_C7811_;
  assign new_C7859_ = new_C7827_ | new_C7864_;
  assign new_C7860_ = ~new_C7827_ & ~new_C7863_;
  assign new_C7861_ = new_C7810_ | new_C7827_;
  assign new_C7862_ = new_C7810_ | new_C7811_;
  assign new_C7863_ = new_C7827_ & new_C7864_;
  assign new_C7864_ = ~new_C7809_ | ~new_C7834_;
  assign new_C7865_ = new_C7842_ & new_C7862_;
  assign new_C7866_ = ~new_C7842_ & ~new_C7862_;
  assign new_C7867_ = new_C7871_ | new_C7872_;
  assign new_C7868_ = ~new_C7813_ & new_C7827_;
  assign new_C7869_ = new_C7873_ | new_C7874_;
  assign new_C7870_ = new_C7813_ & new_C7827_;
  assign new_C7871_ = ~new_C7813_ & ~new_C7827_;
  assign new_C7872_ = new_C7813_ & ~new_C7827_;
  assign new_C7873_ = new_C7813_ & ~new_C7827_;
  assign new_C7874_ = ~new_C7813_ & new_C7827_;
  assign new_C7875_ = new_E213_;
  assign new_C7876_ = new_E280_;
  assign new_C7877_ = new_E347_;
  assign new_C7878_ = new_E414_;
  assign new_C7879_ = new_E481_;
  assign new_C7880_ = new_E548_;
  assign new_C7881_ = new_C7888_ & new_C7887_;
  assign new_C7882_ = new_C7890_ | new_C7889_;
  assign new_C7883_ = new_C7892_ | new_C7891_;
  assign new_C7884_ = new_C7894_ & new_C7893_;
  assign new_C7885_ = new_C7894_ & new_C7895_;
  assign new_C7886_ = new_C7887_ | new_C7896_;
  assign new_C7887_ = new_C7876_ | new_C7899_;
  assign new_C7888_ = new_C7898_ | new_C7897_;
  assign new_C7889_ = new_C7903_ & new_C7902_;
  assign new_C7890_ = new_C7901_ & new_C7900_;
  assign new_C7891_ = new_C7906_ | new_C7905_;
  assign new_C7892_ = new_C7901_ & new_C7904_;
  assign new_C7893_ = new_C7876_ | new_C7909_;
  assign new_C7894_ = new_C7908_ | new_C7907_;
  assign new_C7895_ = new_C7911_ | new_C7910_;
  assign new_C7896_ = ~new_C7887_ & new_C7913_;
  assign new_C7897_ = ~new_C7889_ & new_C7901_;
  assign new_C7898_ = new_C7889_ & ~new_C7901_;
  assign new_C7899_ = new_C7875_ & ~new_C7876_;
  assign new_C7900_ = ~new_C7922_ | ~new_C7923_;
  assign new_C7901_ = new_C7915_ | new_C7917_;
  assign new_C7902_ = new_C7925_ | new_C7924_;
  assign new_C7903_ = new_C7919_ | new_C7918_;
  assign new_C7904_ = ~new_C7927_ | ~new_C7926_;
  assign new_C7905_ = ~new_C7928_ & new_C7929_;
  assign new_C7906_ = new_C7928_ & ~new_C7929_;
  assign new_C7907_ = ~new_C7875_ & new_C7876_;
  assign new_C7908_ = new_C7875_ & ~new_C7876_;
  assign new_C7909_ = ~new_C7891_ | new_C7901_;
  assign new_C7910_ = new_C7891_ & new_C7901_;
  assign new_C7911_ = ~new_C7891_ & ~new_C7901_;
  assign new_C7912_ = new_C7933_ | new_C7932_;
  assign new_C7913_ = new_C7879_ | new_C7912_;
  assign new_C7914_ = new_C7937_ | new_C7936_;
  assign new_C7915_ = ~new_C7879_ & new_C7914_;
  assign new_C7916_ = new_C7935_ | new_C7934_;
  assign new_C7917_ = new_C7879_ & new_C7916_;
  assign new_C7918_ = new_C7877_ & ~new_C7887_;
  assign new_C7919_ = ~new_C7877_ & new_C7887_;
  assign new_C7920_ = ~new_C7876_ | ~new_C7901_;
  assign new_C7921_ = new_C7887_ & new_C7920_;
  assign new_C7922_ = ~new_C7887_ & ~new_C7921_;
  assign new_C7923_ = new_C7887_ | new_C7920_;
  assign new_C7924_ = ~new_C7877_ & new_C7878_;
  assign new_C7925_ = new_C7877_ & ~new_C7878_;
  assign new_C7926_ = new_C7894_ | new_C7931_;
  assign new_C7927_ = ~new_C7894_ & ~new_C7930_;
  assign new_C7928_ = new_C7877_ | new_C7894_;
  assign new_C7929_ = new_C7877_ | new_C7878_;
  assign new_C7930_ = new_C7894_ & new_C7931_;
  assign new_C7931_ = ~new_C7876_ | ~new_C7901_;
  assign new_C7932_ = new_C7909_ & new_C7929_;
  assign new_C7933_ = ~new_C7909_ & ~new_C7929_;
  assign new_C7934_ = new_C7938_ | new_C7939_;
  assign new_C7935_ = ~new_C7880_ & new_C7894_;
  assign new_C7936_ = new_C7940_ | new_C7941_;
  assign new_C7937_ = new_C7880_ & new_C7894_;
  assign new_C7938_ = ~new_C7880_ & ~new_C7894_;
  assign new_C7939_ = new_C7880_ & ~new_C7894_;
  assign new_C7940_ = new_C7880_ & ~new_C7894_;
  assign new_C7941_ = ~new_C7880_ & new_C7894_;
  assign new_C7942_ = new_E615_;
  assign new_C7943_ = new_E682_;
  assign new_C7944_ = new_E749_;
  assign new_C7945_ = new_E816_;
  assign new_C7946_ = new_E883_;
  assign new_C7947_ = new_E950_;
  assign new_C7948_ = new_C7955_ & new_C7954_;
  assign new_C7949_ = new_C7957_ | new_C7956_;
  assign new_C7950_ = new_C7959_ | new_C7958_;
  assign new_C7951_ = new_C7961_ & new_C7960_;
  assign new_C7952_ = new_C7961_ & new_C7962_;
  assign new_C7953_ = new_C7954_ | new_C7963_;
  assign new_C7954_ = new_C7943_ | new_C7966_;
  assign new_C7955_ = new_C7965_ | new_C7964_;
  assign new_C7956_ = new_C7970_ & new_C7969_;
  assign new_C7957_ = new_C7968_ & new_C7967_;
  assign new_C7958_ = new_C7973_ | new_C7972_;
  assign new_C7959_ = new_C7968_ & new_C7971_;
  assign new_C7960_ = new_C7943_ | new_C7976_;
  assign new_C7961_ = new_C7975_ | new_C7974_;
  assign new_C7962_ = new_C7978_ | new_C7977_;
  assign new_C7963_ = ~new_C7954_ & new_C7980_;
  assign new_C7964_ = ~new_C7956_ & new_C7968_;
  assign new_C7965_ = new_C7956_ & ~new_C7968_;
  assign new_C7966_ = new_C7942_ & ~new_C7943_;
  assign new_C7967_ = ~new_C7989_ | ~new_C7990_;
  assign new_C7968_ = new_C7982_ | new_C7984_;
  assign new_C7969_ = new_C7992_ | new_C7991_;
  assign new_C7970_ = new_C7986_ | new_C7985_;
  assign new_C7971_ = ~new_C7994_ | ~new_C7993_;
  assign new_C7972_ = ~new_C7995_ & new_C7996_;
  assign new_C7973_ = new_C7995_ & ~new_C7996_;
  assign new_C7974_ = ~new_C7942_ & new_C7943_;
  assign new_C7975_ = new_C7942_ & ~new_C7943_;
  assign new_C7976_ = ~new_C7958_ | new_C7968_;
  assign new_C7977_ = new_C7958_ & new_C7968_;
  assign new_C7978_ = ~new_C7958_ & ~new_C7968_;
  assign new_C7979_ = new_C8000_ | new_C7999_;
  assign new_C7980_ = new_C7946_ | new_C7979_;
  assign new_C7981_ = new_C8004_ | new_C8003_;
  assign new_C7982_ = ~new_C7946_ & new_C7981_;
  assign new_C7983_ = new_C8002_ | new_C8001_;
  assign new_C7984_ = new_C7946_ & new_C7983_;
  assign new_C7985_ = new_C7944_ & ~new_C7954_;
  assign new_C7986_ = ~new_C7944_ & new_C7954_;
  assign new_C7987_ = ~new_C7943_ | ~new_C7968_;
  assign new_C7988_ = new_C7954_ & new_C7987_;
  assign new_C7989_ = ~new_C7954_ & ~new_C7988_;
  assign new_C7990_ = new_C7954_ | new_C7987_;
  assign new_C7991_ = ~new_C7944_ & new_C7945_;
  assign new_C7992_ = new_C7944_ & ~new_C7945_;
  assign new_C7993_ = new_C7961_ | new_C7998_;
  assign new_C7994_ = ~new_C7961_ & ~new_C7997_;
  assign new_C7995_ = new_C7944_ | new_C7961_;
  assign new_C7996_ = new_C7944_ | new_C7945_;
  assign new_C7997_ = new_C7961_ & new_C7998_;
  assign new_C7998_ = ~new_C7943_ | ~new_C7968_;
  assign new_C7999_ = new_C7976_ & new_C7996_;
  assign new_C8000_ = ~new_C7976_ & ~new_C7996_;
  assign new_C8001_ = new_C8005_ | new_C8006_;
  assign new_C8002_ = ~new_C7947_ & new_C7961_;
  assign new_C8003_ = new_C8007_ | new_C8008_;
  assign new_C8004_ = new_C7947_ & new_C7961_;
  assign new_C8005_ = ~new_C7947_ & ~new_C7961_;
  assign new_C8006_ = new_C7947_ & ~new_C7961_;
  assign new_C8007_ = new_C7947_ & ~new_C7961_;
  assign new_C8008_ = ~new_C7947_ & new_C7961_;
  assign new_C8009_ = new_E1017_;
  assign new_C8010_ = new_E1084_;
  assign new_C8011_ = new_E1151_;
  assign new_C8012_ = new_E1218_;
  assign new_C8013_ = new_E1285_;
  assign new_C8014_ = new_E1352_;
  assign new_C8015_ = new_C8022_ & new_C8021_;
  assign new_C8016_ = new_C8024_ | new_C8023_;
  assign new_C8017_ = new_C8026_ | new_C8025_;
  assign new_C8018_ = new_C8028_ & new_C8027_;
  assign new_C8019_ = new_C8028_ & new_C8029_;
  assign new_C8020_ = new_C8021_ | new_C8030_;
  assign new_C8021_ = new_C8010_ | new_C8033_;
  assign new_C8022_ = new_C8032_ | new_C8031_;
  assign new_C8023_ = new_C8037_ & new_C8036_;
  assign new_C8024_ = new_C8035_ & new_C8034_;
  assign new_C8025_ = new_C8040_ | new_C8039_;
  assign new_C8026_ = new_C8035_ & new_C8038_;
  assign new_C8027_ = new_C8010_ | new_C8043_;
  assign new_C8028_ = new_C8042_ | new_C8041_;
  assign new_C8029_ = new_C8045_ | new_C8044_;
  assign new_C8030_ = ~new_C8021_ & new_C8047_;
  assign new_C8031_ = ~new_C8023_ & new_C8035_;
  assign new_C8032_ = new_C8023_ & ~new_C8035_;
  assign new_C8033_ = new_C8009_ & ~new_C8010_;
  assign new_C8034_ = ~new_C8056_ | ~new_C8057_;
  assign new_C8035_ = new_C8049_ | new_C8051_;
  assign new_C8036_ = new_C8059_ | new_C8058_;
  assign new_C8037_ = new_C8053_ | new_C8052_;
  assign new_C8038_ = ~new_C8061_ | ~new_C8060_;
  assign new_C8039_ = ~new_C8062_ & new_C8063_;
  assign new_C8040_ = new_C8062_ & ~new_C8063_;
  assign new_C8041_ = ~new_C8009_ & new_C8010_;
  assign new_C8042_ = new_C8009_ & ~new_C8010_;
  assign new_C8043_ = ~new_C8025_ | new_C8035_;
  assign new_C8044_ = new_C8025_ & new_C8035_;
  assign new_C8045_ = ~new_C8025_ & ~new_C8035_;
  assign new_C8046_ = new_C8067_ | new_C8066_;
  assign new_C8047_ = new_C8013_ | new_C8046_;
  assign new_C8048_ = new_C8071_ | new_C8070_;
  assign new_C8049_ = ~new_C8013_ & new_C8048_;
  assign new_C8050_ = new_C8069_ | new_C8068_;
  assign new_C8051_ = new_C8013_ & new_C8050_;
  assign new_C8052_ = new_C8011_ & ~new_C8021_;
  assign new_C8053_ = ~new_C8011_ & new_C8021_;
  assign new_C8054_ = ~new_C8010_ | ~new_C8035_;
  assign new_C8055_ = new_C8021_ & new_C8054_;
  assign new_C8056_ = ~new_C8021_ & ~new_C8055_;
  assign new_C8057_ = new_C8021_ | new_C8054_;
  assign new_C8058_ = ~new_C8011_ & new_C8012_;
  assign new_C8059_ = new_C8011_ & ~new_C8012_;
  assign new_C8060_ = new_C8028_ | new_C8065_;
  assign new_C8061_ = ~new_C8028_ & ~new_C8064_;
  assign new_C8062_ = new_C8011_ | new_C8028_;
  assign new_C8063_ = new_C8011_ | new_C8012_;
  assign new_C8064_ = new_C8028_ & new_C8065_;
  assign new_C8065_ = ~new_C8010_ | ~new_C8035_;
  assign new_C8066_ = new_C8043_ & new_C8063_;
  assign new_C8067_ = ~new_C8043_ & ~new_C8063_;
  assign new_C8068_ = new_C8072_ | new_C8073_;
  assign new_C8069_ = ~new_C8014_ & new_C8028_;
  assign new_C8070_ = new_C8074_ | new_C8075_;
  assign new_C8071_ = new_C8014_ & new_C8028_;
  assign new_C8072_ = ~new_C8014_ & ~new_C8028_;
  assign new_C8073_ = new_C8014_ & ~new_C8028_;
  assign new_C8074_ = new_C8014_ & ~new_C8028_;
  assign new_C8075_ = ~new_C8014_ & new_C8028_;
  assign new_C8076_ = new_E1419_;
  assign new_C8077_ = new_E1486_;
  assign new_C8078_ = new_E1553_;
  assign new_C8079_ = new_E1620_;
  assign new_C8080_ = new_E1687_;
  assign new_C8081_ = new_E1754_;
  assign new_C8082_ = new_C8089_ & new_C8088_;
  assign new_C8083_ = new_C8091_ | new_C8090_;
  assign new_C8084_ = new_C8093_ | new_C8092_;
  assign new_C8085_ = new_C8095_ & new_C8094_;
  assign new_C8086_ = new_C8095_ & new_C8096_;
  assign new_C8087_ = new_C8088_ | new_C8097_;
  assign new_C8088_ = new_C8077_ | new_C8100_;
  assign new_C8089_ = new_C8099_ | new_C8098_;
  assign new_C8090_ = new_C8104_ & new_C8103_;
  assign new_C8091_ = new_C8102_ & new_C8101_;
  assign new_C8092_ = new_C8107_ | new_C8106_;
  assign new_C8093_ = new_C8102_ & new_C8105_;
  assign new_C8094_ = new_C8077_ | new_C8110_;
  assign new_C8095_ = new_C8109_ | new_C8108_;
  assign new_C8096_ = new_C8112_ | new_C8111_;
  assign new_C8097_ = ~new_C8088_ & new_C8114_;
  assign new_C8098_ = ~new_C8090_ & new_C8102_;
  assign new_C8099_ = new_C8090_ & ~new_C8102_;
  assign new_C8100_ = new_C8076_ & ~new_C8077_;
  assign new_C8101_ = ~new_C8123_ | ~new_C8124_;
  assign new_C8102_ = new_C8116_ | new_C8118_;
  assign new_C8103_ = new_C8126_ | new_C8125_;
  assign new_C8104_ = new_C8120_ | new_C8119_;
  assign new_C8105_ = ~new_C8128_ | ~new_C8127_;
  assign new_C8106_ = ~new_C8129_ & new_C8130_;
  assign new_C8107_ = new_C8129_ & ~new_C8130_;
  assign new_C8108_ = ~new_C8076_ & new_C8077_;
  assign new_C8109_ = new_C8076_ & ~new_C8077_;
  assign new_C8110_ = ~new_C8092_ | new_C8102_;
  assign new_C8111_ = new_C8092_ & new_C8102_;
  assign new_C8112_ = ~new_C8092_ & ~new_C8102_;
  assign new_C8113_ = new_C8134_ | new_C8133_;
  assign new_C8114_ = new_C8080_ | new_C8113_;
  assign new_C8115_ = new_C8138_ | new_C8137_;
  assign new_C8116_ = ~new_C8080_ & new_C8115_;
  assign new_C8117_ = new_C8136_ | new_C8135_;
  assign new_C8118_ = new_C8080_ & new_C8117_;
  assign new_C8119_ = new_C8078_ & ~new_C8088_;
  assign new_C8120_ = ~new_C8078_ & new_C8088_;
  assign new_C8121_ = ~new_C8077_ | ~new_C8102_;
  assign new_C8122_ = new_C8088_ & new_C8121_;
  assign new_C8123_ = ~new_C8088_ & ~new_C8122_;
  assign new_C8124_ = new_C8088_ | new_C8121_;
  assign new_C8125_ = ~new_C8078_ & new_C8079_;
  assign new_C8126_ = new_C8078_ & ~new_C8079_;
  assign new_C8127_ = new_C8095_ | new_C8132_;
  assign new_C8128_ = ~new_C8095_ & ~new_C8131_;
  assign new_C8129_ = new_C8078_ | new_C8095_;
  assign new_C8130_ = new_C8078_ | new_C8079_;
  assign new_C8131_ = new_C8095_ & new_C8132_;
  assign new_C8132_ = ~new_C8077_ | ~new_C8102_;
  assign new_C8133_ = new_C8110_ & new_C8130_;
  assign new_C8134_ = ~new_C8110_ & ~new_C8130_;
  assign new_C8135_ = new_C8139_ | new_C8140_;
  assign new_C8136_ = ~new_C8081_ & new_C8095_;
  assign new_C8137_ = new_C8141_ | new_C8142_;
  assign new_C8138_ = new_C8081_ & new_C8095_;
  assign new_C8139_ = ~new_C8081_ & ~new_C8095_;
  assign new_C8140_ = new_C8081_ & ~new_C8095_;
  assign new_C8141_ = new_C8081_ & ~new_C8095_;
  assign new_C8142_ = ~new_C8081_ & new_C8095_;
  assign new_C8143_ = new_E1821_;
  assign new_C8144_ = new_E1888_;
  assign new_C8145_ = new_E1955_;
  assign new_C8146_ = new_E2022_;
  assign new_C8147_ = new_E2089_;
  assign new_C8148_ = new_E2156_;
  assign new_C8149_ = new_C8156_ & new_C8155_;
  assign new_C8150_ = new_C8158_ | new_C8157_;
  assign new_C8151_ = new_C8160_ | new_C8159_;
  assign new_C8152_ = new_C8162_ & new_C8161_;
  assign new_C8153_ = new_C8162_ & new_C8163_;
  assign new_C8154_ = new_C8155_ | new_C8164_;
  assign new_C8155_ = new_C8144_ | new_C8167_;
  assign new_C8156_ = new_C8166_ | new_C8165_;
  assign new_C8157_ = new_C8171_ & new_C8170_;
  assign new_C8158_ = new_C8169_ & new_C8168_;
  assign new_C8159_ = new_C8174_ | new_C8173_;
  assign new_C8160_ = new_C8169_ & new_C8172_;
  assign new_C8161_ = new_C8144_ | new_C8177_;
  assign new_C8162_ = new_C8176_ | new_C8175_;
  assign new_C8163_ = new_C8179_ | new_C8178_;
  assign new_C8164_ = ~new_C8155_ & new_C8181_;
  assign new_C8165_ = ~new_C8157_ & new_C8169_;
  assign new_C8166_ = new_C8157_ & ~new_C8169_;
  assign new_C8167_ = new_C8143_ & ~new_C8144_;
  assign new_C8168_ = ~new_C8190_ | ~new_C8191_;
  assign new_C8169_ = new_C8183_ | new_C8185_;
  assign new_C8170_ = new_C8193_ | new_C8192_;
  assign new_C8171_ = new_C8187_ | new_C8186_;
  assign new_C8172_ = ~new_C8195_ | ~new_C8194_;
  assign new_C8173_ = ~new_C8196_ & new_C8197_;
  assign new_C8174_ = new_C8196_ & ~new_C8197_;
  assign new_C8175_ = ~new_C8143_ & new_C8144_;
  assign new_C8176_ = new_C8143_ & ~new_C8144_;
  assign new_C8177_ = ~new_C8159_ | new_C8169_;
  assign new_C8178_ = new_C8159_ & new_C8169_;
  assign new_C8179_ = ~new_C8159_ & ~new_C8169_;
  assign new_C8180_ = new_C8201_ | new_C8200_;
  assign new_C8181_ = new_C8147_ | new_C8180_;
  assign new_C8182_ = new_C8205_ | new_C8204_;
  assign new_C8183_ = ~new_C8147_ & new_C8182_;
  assign new_C8184_ = new_C8203_ | new_C8202_;
  assign new_C8185_ = new_C8147_ & new_C8184_;
  assign new_C8186_ = new_C8145_ & ~new_C8155_;
  assign new_C8187_ = ~new_C8145_ & new_C8155_;
  assign new_C8188_ = ~new_C8144_ | ~new_C8169_;
  assign new_C8189_ = new_C8155_ & new_C8188_;
  assign new_C8190_ = ~new_C8155_ & ~new_C8189_;
  assign new_C8191_ = new_C8155_ | new_C8188_;
  assign new_C8192_ = ~new_C8145_ & new_C8146_;
  assign new_C8193_ = new_C8145_ & ~new_C8146_;
  assign new_C8194_ = new_C8162_ | new_C8199_;
  assign new_C8195_ = ~new_C8162_ & ~new_C8198_;
  assign new_C8196_ = new_C8145_ | new_C8162_;
  assign new_C8197_ = new_C8145_ | new_C8146_;
  assign new_C8198_ = new_C8162_ & new_C8199_;
  assign new_C8199_ = ~new_C8144_ | ~new_C8169_;
  assign new_C8200_ = new_C8177_ & new_C8197_;
  assign new_C8201_ = ~new_C8177_ & ~new_C8197_;
  assign new_C8202_ = new_C8206_ | new_C8207_;
  assign new_C8203_ = ~new_C8148_ & new_C8162_;
  assign new_C8204_ = new_C8208_ | new_C8209_;
  assign new_C8205_ = new_C8148_ & new_C8162_;
  assign new_C8206_ = ~new_C8148_ & ~new_C8162_;
  assign new_C8207_ = new_C8148_ & ~new_C8162_;
  assign new_C8208_ = new_C8148_ & ~new_C8162_;
  assign new_C8209_ = ~new_C8148_ & new_C8162_;
  assign new_C8210_ = new_E2223_;
  assign new_C8211_ = new_E2290_;
  assign new_C8212_ = new_E2357_;
  assign new_C8213_ = new_E2424_;
  assign new_C8214_ = new_E2491_;
  assign new_C8215_ = new_E2558_;
  assign new_C8216_ = new_C8223_ & new_C8222_;
  assign new_C8217_ = new_C8225_ | new_C8224_;
  assign new_C8218_ = new_C8227_ | new_C8226_;
  assign new_C8219_ = new_C8229_ & new_C8228_;
  assign new_C8220_ = new_C8229_ & new_C8230_;
  assign new_C8221_ = new_C8222_ | new_C8231_;
  assign new_C8222_ = new_C8211_ | new_C8234_;
  assign new_C8223_ = new_C8233_ | new_C8232_;
  assign new_C8224_ = new_C8238_ & new_C8237_;
  assign new_C8225_ = new_C8236_ & new_C8235_;
  assign new_C8226_ = new_C8241_ | new_C8240_;
  assign new_C8227_ = new_C8236_ & new_C8239_;
  assign new_C8228_ = new_C8211_ | new_C8244_;
  assign new_C8229_ = new_C8243_ | new_C8242_;
  assign new_C8230_ = new_C8246_ | new_C8245_;
  assign new_C8231_ = ~new_C8222_ & new_C8248_;
  assign new_C8232_ = ~new_C8224_ & new_C8236_;
  assign new_C8233_ = new_C8224_ & ~new_C8236_;
  assign new_C8234_ = new_C8210_ & ~new_C8211_;
  assign new_C8235_ = ~new_C8257_ | ~new_C8258_;
  assign new_C8236_ = new_C8250_ | new_C8252_;
  assign new_C8237_ = new_C8260_ | new_C8259_;
  assign new_C8238_ = new_C8254_ | new_C8253_;
  assign new_C8239_ = ~new_C8262_ | ~new_C8261_;
  assign new_C8240_ = ~new_C8263_ & new_C8264_;
  assign new_C8241_ = new_C8263_ & ~new_C8264_;
  assign new_C8242_ = ~new_C8210_ & new_C8211_;
  assign new_C8243_ = new_C8210_ & ~new_C8211_;
  assign new_C8244_ = ~new_C8226_ | new_C8236_;
  assign new_C8245_ = new_C8226_ & new_C8236_;
  assign new_C8246_ = ~new_C8226_ & ~new_C8236_;
  assign new_C8247_ = new_C8268_ | new_C8267_;
  assign new_C8248_ = new_C8214_ | new_C8247_;
  assign new_C8249_ = new_C8272_ | new_C8271_;
  assign new_C8250_ = ~new_C8214_ & new_C8249_;
  assign new_C8251_ = new_C8270_ | new_C8269_;
  assign new_C8252_ = new_C8214_ & new_C8251_;
  assign new_C8253_ = new_C8212_ & ~new_C8222_;
  assign new_C8254_ = ~new_C8212_ & new_C8222_;
  assign new_C8255_ = ~new_C8211_ | ~new_C8236_;
  assign new_C8256_ = new_C8222_ & new_C8255_;
  assign new_C8257_ = ~new_C8222_ & ~new_C8256_;
  assign new_C8258_ = new_C8222_ | new_C8255_;
  assign new_C8259_ = ~new_C8212_ & new_C8213_;
  assign new_C8260_ = new_C8212_ & ~new_C8213_;
  assign new_C8261_ = new_C8229_ | new_C8266_;
  assign new_C8262_ = ~new_C8229_ & ~new_C8265_;
  assign new_C8263_ = new_C8212_ | new_C8229_;
  assign new_C8264_ = new_C8212_ | new_C8213_;
  assign new_C8265_ = new_C8229_ & new_C8266_;
  assign new_C8266_ = ~new_C8211_ | ~new_C8236_;
  assign new_C8267_ = new_C8244_ & new_C8264_;
  assign new_C8268_ = ~new_C8244_ & ~new_C8264_;
  assign new_C8269_ = new_C8273_ | new_C8274_;
  assign new_C8270_ = ~new_C8215_ & new_C8229_;
  assign new_C8271_ = new_C8275_ | new_C8276_;
  assign new_C8272_ = new_C8215_ & new_C8229_;
  assign new_C8273_ = ~new_C8215_ & ~new_C8229_;
  assign new_C8274_ = new_C8215_ & ~new_C8229_;
  assign new_C8275_ = new_C8215_ & ~new_C8229_;
  assign new_C8276_ = ~new_C8215_ & new_C8229_;
  assign new_C8277_ = new_E2625_;
  assign new_C8278_ = new_E2692_;
  assign new_C8279_ = new_E2759_;
  assign new_C8280_ = new_E2826_;
  assign new_C8281_ = new_E2893_;
  assign new_C8282_ = new_E2960_;
  assign new_C8283_ = new_C8290_ & new_C8289_;
  assign new_C8284_ = new_C8292_ | new_C8291_;
  assign new_C8285_ = new_C8294_ | new_C8293_;
  assign new_C8286_ = new_C8296_ & new_C8295_;
  assign new_C8287_ = new_C8296_ & new_C8297_;
  assign new_C8288_ = new_C8289_ | new_C8298_;
  assign new_C8289_ = new_C8278_ | new_C8301_;
  assign new_C8290_ = new_C8300_ | new_C8299_;
  assign new_C8291_ = new_C8305_ & new_C8304_;
  assign new_C8292_ = new_C8303_ & new_C8302_;
  assign new_C8293_ = new_C8308_ | new_C8307_;
  assign new_C8294_ = new_C8303_ & new_C8306_;
  assign new_C8295_ = new_C8278_ | new_C8311_;
  assign new_C8296_ = new_C8310_ | new_C8309_;
  assign new_C8297_ = new_C8313_ | new_C8312_;
  assign new_C8298_ = ~new_C8289_ & new_C8315_;
  assign new_C8299_ = ~new_C8291_ & new_C8303_;
  assign new_C8300_ = new_C8291_ & ~new_C8303_;
  assign new_C8301_ = new_C8277_ & ~new_C8278_;
  assign new_C8302_ = ~new_C8324_ | ~new_C8325_;
  assign new_C8303_ = new_C8317_ | new_C8319_;
  assign new_C8304_ = new_C8327_ | new_C8326_;
  assign new_C8305_ = new_C8321_ | new_C8320_;
  assign new_C8306_ = ~new_C8329_ | ~new_C8328_;
  assign new_C8307_ = ~new_C8330_ & new_C8331_;
  assign new_C8308_ = new_C8330_ & ~new_C8331_;
  assign new_C8309_ = ~new_C8277_ & new_C8278_;
  assign new_C8310_ = new_C8277_ & ~new_C8278_;
  assign new_C8311_ = ~new_C8293_ | new_C8303_;
  assign new_C8312_ = new_C8293_ & new_C8303_;
  assign new_C8313_ = ~new_C8293_ & ~new_C8303_;
  assign new_C8314_ = new_C8335_ | new_C8334_;
  assign new_C8315_ = new_C8281_ | new_C8314_;
  assign new_C8316_ = new_C8339_ | new_C8338_;
  assign new_C8317_ = ~new_C8281_ & new_C8316_;
  assign new_C8318_ = new_C8337_ | new_C8336_;
  assign new_C8319_ = new_C8281_ & new_C8318_;
  assign new_C8320_ = new_C8279_ & ~new_C8289_;
  assign new_C8321_ = ~new_C8279_ & new_C8289_;
  assign new_C8322_ = ~new_C8278_ | ~new_C8303_;
  assign new_C8323_ = new_C8289_ & new_C8322_;
  assign new_C8324_ = ~new_C8289_ & ~new_C8323_;
  assign new_C8325_ = new_C8289_ | new_C8322_;
  assign new_C8326_ = ~new_C8279_ & new_C8280_;
  assign new_C8327_ = new_C8279_ & ~new_C8280_;
  assign new_C8328_ = new_C8296_ | new_C8333_;
  assign new_C8329_ = ~new_C8296_ & ~new_C8332_;
  assign new_C8330_ = new_C8279_ | new_C8296_;
  assign new_C8331_ = new_C8279_ | new_C8280_;
  assign new_C8332_ = new_C8296_ & new_C8333_;
  assign new_C8333_ = ~new_C8278_ | ~new_C8303_;
  assign new_C8334_ = new_C8311_ & new_C8331_;
  assign new_C8335_ = ~new_C8311_ & ~new_C8331_;
  assign new_C8336_ = new_C8340_ | new_C8341_;
  assign new_C8337_ = ~new_C8282_ & new_C8296_;
  assign new_C8338_ = new_C8342_ | new_C8343_;
  assign new_C8339_ = new_C8282_ & new_C8296_;
  assign new_C8340_ = ~new_C8282_ & ~new_C8296_;
  assign new_C8341_ = new_C8282_ & ~new_C8296_;
  assign new_C8342_ = new_C8282_ & ~new_C8296_;
  assign new_C8343_ = ~new_C8282_ & new_C8296_;
  assign new_C8344_ = new_E3027_;
  assign new_C8345_ = new_E3094_;
  assign new_C8346_ = new_E3161_;
  assign new_C8347_ = new_E3228_;
  assign new_C8348_ = new_E3295_;
  assign new_C8349_ = new_E3362_;
  assign new_C8350_ = new_C8357_ & new_C8356_;
  assign new_C8351_ = new_C8359_ | new_C8358_;
  assign new_C8352_ = new_C8361_ | new_C8360_;
  assign new_C8353_ = new_C8363_ & new_C8362_;
  assign new_C8354_ = new_C8363_ & new_C8364_;
  assign new_C8355_ = new_C8356_ | new_C8365_;
  assign new_C8356_ = new_C8345_ | new_C8368_;
  assign new_C8357_ = new_C8367_ | new_C8366_;
  assign new_C8358_ = new_C8372_ & new_C8371_;
  assign new_C8359_ = new_C8370_ & new_C8369_;
  assign new_C8360_ = new_C8375_ | new_C8374_;
  assign new_C8361_ = new_C8370_ & new_C8373_;
  assign new_C8362_ = new_C8345_ | new_C8378_;
  assign new_C8363_ = new_C8377_ | new_C8376_;
  assign new_C8364_ = new_C8380_ | new_C8379_;
  assign new_C8365_ = ~new_C8356_ & new_C8382_;
  assign new_C8366_ = ~new_C8358_ & new_C8370_;
  assign new_C8367_ = new_C8358_ & ~new_C8370_;
  assign new_C8368_ = new_C8344_ & ~new_C8345_;
  assign new_C8369_ = ~new_C8391_ | ~new_C8392_;
  assign new_C8370_ = new_C8384_ | new_C8386_;
  assign new_C8371_ = new_C8394_ | new_C8393_;
  assign new_C8372_ = new_C8388_ | new_C8387_;
  assign new_C8373_ = ~new_C8396_ | ~new_C8395_;
  assign new_C8374_ = ~new_C8397_ & new_C8398_;
  assign new_C8375_ = new_C8397_ & ~new_C8398_;
  assign new_C8376_ = ~new_C8344_ & new_C8345_;
  assign new_C8377_ = new_C8344_ & ~new_C8345_;
  assign new_C8378_ = ~new_C8360_ | new_C8370_;
  assign new_C8379_ = new_C8360_ & new_C8370_;
  assign new_C8380_ = ~new_C8360_ & ~new_C8370_;
  assign new_C8381_ = new_C8402_ | new_C8401_;
  assign new_C8382_ = new_C8348_ | new_C8381_;
  assign new_C8383_ = new_C8406_ | new_C8405_;
  assign new_C8384_ = ~new_C8348_ & new_C8383_;
  assign new_C8385_ = new_C8404_ | new_C8403_;
  assign new_C8386_ = new_C8348_ & new_C8385_;
  assign new_C8387_ = new_C8346_ & ~new_C8356_;
  assign new_C8388_ = ~new_C8346_ & new_C8356_;
  assign new_C8389_ = ~new_C8345_ | ~new_C8370_;
  assign new_C8390_ = new_C8356_ & new_C8389_;
  assign new_C8391_ = ~new_C8356_ & ~new_C8390_;
  assign new_C8392_ = new_C8356_ | new_C8389_;
  assign new_C8393_ = ~new_C8346_ & new_C8347_;
  assign new_C8394_ = new_C8346_ & ~new_C8347_;
  assign new_C8395_ = new_C8363_ | new_C8400_;
  assign new_C8396_ = ~new_C8363_ & ~new_C8399_;
  assign new_C8397_ = new_C8346_ | new_C8363_;
  assign new_C8398_ = new_C8346_ | new_C8347_;
  assign new_C8399_ = new_C8363_ & new_C8400_;
  assign new_C8400_ = ~new_C8345_ | ~new_C8370_;
  assign new_C8401_ = new_C8378_ & new_C8398_;
  assign new_C8402_ = ~new_C8378_ & ~new_C8398_;
  assign new_C8403_ = new_C8407_ | new_C8408_;
  assign new_C8404_ = ~new_C8349_ & new_C8363_;
  assign new_C8405_ = new_C8409_ | new_C8410_;
  assign new_C8406_ = new_C8349_ & new_C8363_;
  assign new_C8407_ = ~new_C8349_ & ~new_C8363_;
  assign new_C8408_ = new_C8349_ & ~new_C8363_;
  assign new_C8409_ = new_C8349_ & ~new_C8363_;
  assign new_C8410_ = ~new_C8349_ & new_C8363_;
  assign new_C8411_ = new_E3429_;
  assign new_C8412_ = new_E3496_;
  assign new_C8413_ = new_E3563_;
  assign new_C8414_ = new_E3630_;
  assign new_C8415_ = new_E3697_;
  assign new_C8416_ = new_E3764_;
  assign new_C8417_ = new_C8424_ & new_C8423_;
  assign new_C8418_ = new_C8426_ | new_C8425_;
  assign new_C8419_ = new_C8428_ | new_C8427_;
  assign new_C8420_ = new_C8430_ & new_C8429_;
  assign new_C8421_ = new_C8430_ & new_C8431_;
  assign new_C8422_ = new_C8423_ | new_C8432_;
  assign new_C8423_ = new_C8412_ | new_C8435_;
  assign new_C8424_ = new_C8434_ | new_C8433_;
  assign new_C8425_ = new_C8439_ & new_C8438_;
  assign new_C8426_ = new_C8437_ & new_C8436_;
  assign new_C8427_ = new_C8442_ | new_C8441_;
  assign new_C8428_ = new_C8437_ & new_C8440_;
  assign new_C8429_ = new_C8412_ | new_C8445_;
  assign new_C8430_ = new_C8444_ | new_C8443_;
  assign new_C8431_ = new_C8447_ | new_C8446_;
  assign new_C8432_ = ~new_C8423_ & new_C8449_;
  assign new_C8433_ = ~new_C8425_ & new_C8437_;
  assign new_C8434_ = new_C8425_ & ~new_C8437_;
  assign new_C8435_ = new_C8411_ & ~new_C8412_;
  assign new_C8436_ = ~new_C8458_ | ~new_C8459_;
  assign new_C8437_ = new_C8451_ | new_C8453_;
  assign new_C8438_ = new_C8461_ | new_C8460_;
  assign new_C8439_ = new_C8455_ | new_C8454_;
  assign new_C8440_ = ~new_C8463_ | ~new_C8462_;
  assign new_C8441_ = ~new_C8464_ & new_C8465_;
  assign new_C8442_ = new_C8464_ & ~new_C8465_;
  assign new_C8443_ = ~new_C8411_ & new_C8412_;
  assign new_C8444_ = new_C8411_ & ~new_C8412_;
  assign new_C8445_ = ~new_C8427_ | new_C8437_;
  assign new_C8446_ = new_C8427_ & new_C8437_;
  assign new_C8447_ = ~new_C8427_ & ~new_C8437_;
  assign new_C8448_ = new_C8469_ | new_C8468_;
  assign new_C8449_ = new_C8415_ | new_C8448_;
  assign new_C8450_ = new_C8473_ | new_C8472_;
  assign new_C8451_ = ~new_C8415_ & new_C8450_;
  assign new_C8452_ = new_C8471_ | new_C8470_;
  assign new_C8453_ = new_C8415_ & new_C8452_;
  assign new_C8454_ = new_C8413_ & ~new_C8423_;
  assign new_C8455_ = ~new_C8413_ & new_C8423_;
  assign new_C8456_ = ~new_C8412_ | ~new_C8437_;
  assign new_C8457_ = new_C8423_ & new_C8456_;
  assign new_C8458_ = ~new_C8423_ & ~new_C8457_;
  assign new_C8459_ = new_C8423_ | new_C8456_;
  assign new_C8460_ = ~new_C8413_ & new_C8414_;
  assign new_C8461_ = new_C8413_ & ~new_C8414_;
  assign new_C8462_ = new_C8430_ | new_C8467_;
  assign new_C8463_ = ~new_C8430_ & ~new_C8466_;
  assign new_C8464_ = new_C8413_ | new_C8430_;
  assign new_C8465_ = new_C8413_ | new_C8414_;
  assign new_C8466_ = new_C8430_ & new_C8467_;
  assign new_C8467_ = ~new_C8412_ | ~new_C8437_;
  assign new_C8468_ = new_C8445_ & new_C8465_;
  assign new_C8469_ = ~new_C8445_ & ~new_C8465_;
  assign new_C8470_ = new_C8474_ | new_C8475_;
  assign new_C8471_ = ~new_C8416_ & new_C8430_;
  assign new_C8472_ = new_C8476_ | new_C8477_;
  assign new_C8473_ = new_C8416_ & new_C8430_;
  assign new_C8474_ = ~new_C8416_ & ~new_C8430_;
  assign new_C8475_ = new_C8416_ & ~new_C8430_;
  assign new_C8476_ = new_C8416_ & ~new_C8430_;
  assign new_C8477_ = ~new_C8416_ & new_C8430_;
  assign new_C8478_ = new_E3831_;
  assign new_C8479_ = new_E3898_;
  assign new_C8480_ = new_E3965_;
  assign new_C8481_ = new_E4032_;
  assign new_C8482_ = new_E4099_;
  assign new_C8483_ = new_E4166_;
  assign new_C8484_ = new_C8491_ & new_C8490_;
  assign new_C8485_ = new_C8493_ | new_C8492_;
  assign new_C8486_ = new_C8495_ | new_C8494_;
  assign new_C8487_ = new_C8497_ & new_C8496_;
  assign new_C8488_ = new_C8497_ & new_C8498_;
  assign new_C8489_ = new_C8490_ | new_C8499_;
  assign new_C8490_ = new_C8479_ | new_C8502_;
  assign new_C8491_ = new_C8501_ | new_C8500_;
  assign new_C8492_ = new_C8506_ & new_C8505_;
  assign new_C8493_ = new_C8504_ & new_C8503_;
  assign new_C8494_ = new_C8509_ | new_C8508_;
  assign new_C8495_ = new_C8504_ & new_C8507_;
  assign new_C8496_ = new_C8479_ | new_C8512_;
  assign new_C8497_ = new_C8511_ | new_C8510_;
  assign new_C8498_ = new_C8514_ | new_C8513_;
  assign new_C8499_ = ~new_C8490_ & new_C8516_;
  assign new_C8500_ = ~new_C8492_ & new_C8504_;
  assign new_C8501_ = new_C8492_ & ~new_C8504_;
  assign new_C8502_ = new_C8478_ & ~new_C8479_;
  assign new_C8503_ = ~new_C8525_ | ~new_C8526_;
  assign new_C8504_ = new_C8518_ | new_C8520_;
  assign new_C8505_ = new_C8528_ | new_C8527_;
  assign new_C8506_ = new_C8522_ | new_C8521_;
  assign new_C8507_ = ~new_C8530_ | ~new_C8529_;
  assign new_C8508_ = ~new_C8531_ & new_C8532_;
  assign new_C8509_ = new_C8531_ & ~new_C8532_;
  assign new_C8510_ = ~new_C8478_ & new_C8479_;
  assign new_C8511_ = new_C8478_ & ~new_C8479_;
  assign new_C8512_ = ~new_C8494_ | new_C8504_;
  assign new_C8513_ = new_C8494_ & new_C8504_;
  assign new_C8514_ = ~new_C8494_ & ~new_C8504_;
  assign new_C8515_ = new_C8536_ | new_C8535_;
  assign new_C8516_ = new_C8482_ | new_C8515_;
  assign new_C8517_ = new_C8540_ | new_C8539_;
  assign new_C8518_ = ~new_C8482_ & new_C8517_;
  assign new_C8519_ = new_C8538_ | new_C8537_;
  assign new_C8520_ = new_C8482_ & new_C8519_;
  assign new_C8521_ = new_C8480_ & ~new_C8490_;
  assign new_C8522_ = ~new_C8480_ & new_C8490_;
  assign new_C8523_ = ~new_C8479_ | ~new_C8504_;
  assign new_C8524_ = new_C8490_ & new_C8523_;
  assign new_C8525_ = ~new_C8490_ & ~new_C8524_;
  assign new_C8526_ = new_C8490_ | new_C8523_;
  assign new_C8527_ = ~new_C8480_ & new_C8481_;
  assign new_C8528_ = new_C8480_ & ~new_C8481_;
  assign new_C8529_ = new_C8497_ | new_C8534_;
  assign new_C8530_ = ~new_C8497_ & ~new_C8533_;
  assign new_C8531_ = new_C8480_ | new_C8497_;
  assign new_C8532_ = new_C8480_ | new_C8481_;
  assign new_C8533_ = new_C8497_ & new_C8534_;
  assign new_C8534_ = ~new_C8479_ | ~new_C8504_;
  assign new_C8535_ = new_C8512_ & new_C8532_;
  assign new_C8536_ = ~new_C8512_ & ~new_C8532_;
  assign new_C8537_ = new_C8541_ | new_C8542_;
  assign new_C8538_ = ~new_C8483_ & new_C8497_;
  assign new_C8539_ = new_C8543_ | new_C8544_;
  assign new_C8540_ = new_C8483_ & new_C8497_;
  assign new_C8541_ = ~new_C8483_ & ~new_C8497_;
  assign new_C8542_ = new_C8483_ & ~new_C8497_;
  assign new_C8543_ = new_C8483_ & ~new_C8497_;
  assign new_C8544_ = ~new_C8483_ & new_C8497_;
  assign new_C8545_ = new_E4233_;
  assign new_C8546_ = new_E4300_;
  assign new_C8547_ = new_E4367_;
  assign new_C8548_ = new_E4434_;
  assign new_C8549_ = new_E4501_;
  assign new_C8550_ = new_E4568_;
  assign new_C8551_ = new_C8558_ & new_C8557_;
  assign new_C8552_ = new_C8560_ | new_C8559_;
  assign new_C8553_ = new_C8562_ | new_C8561_;
  assign new_C8554_ = new_C8564_ & new_C8563_;
  assign new_C8555_ = new_C8564_ & new_C8565_;
  assign new_C8556_ = new_C8557_ | new_C8566_;
  assign new_C8557_ = new_C8546_ | new_C8569_;
  assign new_C8558_ = new_C8568_ | new_C8567_;
  assign new_C8559_ = new_C8573_ & new_C8572_;
  assign new_C8560_ = new_C8571_ & new_C8570_;
  assign new_C8561_ = new_C8576_ | new_C8575_;
  assign new_C8562_ = new_C8571_ & new_C8574_;
  assign new_C8563_ = new_C8546_ | new_C8579_;
  assign new_C8564_ = new_C8578_ | new_C8577_;
  assign new_C8565_ = new_C8581_ | new_C8580_;
  assign new_C8566_ = ~new_C8557_ & new_C8583_;
  assign new_C8567_ = ~new_C8559_ & new_C8571_;
  assign new_C8568_ = new_C8559_ & ~new_C8571_;
  assign new_C8569_ = new_C8545_ & ~new_C8546_;
  assign new_C8570_ = ~new_C8592_ | ~new_C8593_;
  assign new_C8571_ = new_C8585_ | new_C8587_;
  assign new_C8572_ = new_C8595_ | new_C8594_;
  assign new_C8573_ = new_C8589_ | new_C8588_;
  assign new_C8574_ = ~new_C8597_ | ~new_C8596_;
  assign new_C8575_ = ~new_C8598_ & new_C8599_;
  assign new_C8576_ = new_C8598_ & ~new_C8599_;
  assign new_C8577_ = ~new_C8545_ & new_C8546_;
  assign new_C8578_ = new_C8545_ & ~new_C8546_;
  assign new_C8579_ = ~new_C8561_ | new_C8571_;
  assign new_C8580_ = new_C8561_ & new_C8571_;
  assign new_C8581_ = ~new_C8561_ & ~new_C8571_;
  assign new_C8582_ = new_C8603_ | new_C8602_;
  assign new_C8583_ = new_C8549_ | new_C8582_;
  assign new_C8584_ = new_C8607_ | new_C8606_;
  assign new_C8585_ = ~new_C8549_ & new_C8584_;
  assign new_C8586_ = new_C8605_ | new_C8604_;
  assign new_C8587_ = new_C8549_ & new_C8586_;
  assign new_C8588_ = new_C8547_ & ~new_C8557_;
  assign new_C8589_ = ~new_C8547_ & new_C8557_;
  assign new_C8590_ = ~new_C8546_ | ~new_C8571_;
  assign new_C8591_ = new_C8557_ & new_C8590_;
  assign new_C8592_ = ~new_C8557_ & ~new_C8591_;
  assign new_C8593_ = new_C8557_ | new_C8590_;
  assign new_C8594_ = ~new_C8547_ & new_C8548_;
  assign new_C8595_ = new_C8547_ & ~new_C8548_;
  assign new_C8596_ = new_C8564_ | new_C8601_;
  assign new_C8597_ = ~new_C8564_ & ~new_C8600_;
  assign new_C8598_ = new_C8547_ | new_C8564_;
  assign new_C8599_ = new_C8547_ | new_C8548_;
  assign new_C8600_ = new_C8564_ & new_C8601_;
  assign new_C8601_ = ~new_C8546_ | ~new_C8571_;
  assign new_C8602_ = new_C8579_ & new_C8599_;
  assign new_C8603_ = ~new_C8579_ & ~new_C8599_;
  assign new_C8604_ = new_C8608_ | new_C8609_;
  assign new_C8605_ = ~new_C8550_ & new_C8564_;
  assign new_C8606_ = new_C8610_ | new_C8611_;
  assign new_C8607_ = new_C8550_ & new_C8564_;
  assign new_C8608_ = ~new_C8550_ & ~new_C8564_;
  assign new_C8609_ = new_C8550_ & ~new_C8564_;
  assign new_C8610_ = new_C8550_ & ~new_C8564_;
  assign new_C8611_ = ~new_C8550_ & new_C8564_;
  assign new_C8612_ = new_E4635_;
  assign new_C8613_ = new_E4702_;
  assign new_C8614_ = new_E4769_;
  assign new_C8615_ = new_E4836_;
  assign new_C8616_ = new_E4903_;
  assign new_C8617_ = new_E4970_;
  assign new_C8618_ = new_C8625_ & new_C8624_;
  assign new_C8619_ = new_C8627_ | new_C8626_;
  assign new_C8620_ = new_C8629_ | new_C8628_;
  assign new_C8621_ = new_C8631_ & new_C8630_;
  assign new_C8622_ = new_C8631_ & new_C8632_;
  assign new_C8623_ = new_C8624_ | new_C8633_;
  assign new_C8624_ = new_C8613_ | new_C8636_;
  assign new_C8625_ = new_C8635_ | new_C8634_;
  assign new_C8626_ = new_C8640_ & new_C8639_;
  assign new_C8627_ = new_C8638_ & new_C8637_;
  assign new_C8628_ = new_C8643_ | new_C8642_;
  assign new_C8629_ = new_C8638_ & new_C8641_;
  assign new_C8630_ = new_C8613_ | new_C8646_;
  assign new_C8631_ = new_C8645_ | new_C8644_;
  assign new_C8632_ = new_C8648_ | new_C8647_;
  assign new_C8633_ = ~new_C8624_ & new_C8650_;
  assign new_C8634_ = ~new_C8626_ & new_C8638_;
  assign new_C8635_ = new_C8626_ & ~new_C8638_;
  assign new_C8636_ = new_C8612_ & ~new_C8613_;
  assign new_C8637_ = ~new_C8659_ | ~new_C8660_;
  assign new_C8638_ = new_C8652_ | new_C8654_;
  assign new_C8639_ = new_C8662_ | new_C8661_;
  assign new_C8640_ = new_C8656_ | new_C8655_;
  assign new_C8641_ = ~new_C8664_ | ~new_C8663_;
  assign new_C8642_ = ~new_C8665_ & new_C8666_;
  assign new_C8643_ = new_C8665_ & ~new_C8666_;
  assign new_C8644_ = ~new_C8612_ & new_C8613_;
  assign new_C8645_ = new_C8612_ & ~new_C8613_;
  assign new_C8646_ = ~new_C8628_ | new_C8638_;
  assign new_C8647_ = new_C8628_ & new_C8638_;
  assign new_C8648_ = ~new_C8628_ & ~new_C8638_;
  assign new_C8649_ = new_C8670_ | new_C8669_;
  assign new_C8650_ = new_C8616_ | new_C8649_;
  assign new_C8651_ = new_C8674_ | new_C8673_;
  assign new_C8652_ = ~new_C8616_ & new_C8651_;
  assign new_C8653_ = new_C8672_ | new_C8671_;
  assign new_C8654_ = new_C8616_ & new_C8653_;
  assign new_C8655_ = new_C8614_ & ~new_C8624_;
  assign new_C8656_ = ~new_C8614_ & new_C8624_;
  assign new_C8657_ = ~new_C8613_ | ~new_C8638_;
  assign new_C8658_ = new_C8624_ & new_C8657_;
  assign new_C8659_ = ~new_C8624_ & ~new_C8658_;
  assign new_C8660_ = new_C8624_ | new_C8657_;
  assign new_C8661_ = ~new_C8614_ & new_C8615_;
  assign new_C8662_ = new_C8614_ & ~new_C8615_;
  assign new_C8663_ = new_C8631_ | new_C8668_;
  assign new_C8664_ = ~new_C8631_ & ~new_C8667_;
  assign new_C8665_ = new_C8614_ | new_C8631_;
  assign new_C8666_ = new_C8614_ | new_C8615_;
  assign new_C8667_ = new_C8631_ & new_C8668_;
  assign new_C8668_ = ~new_C8613_ | ~new_C8638_;
  assign new_C8669_ = new_C8646_ & new_C8666_;
  assign new_C8670_ = ~new_C8646_ & ~new_C8666_;
  assign new_C8671_ = new_C8675_ | new_C8676_;
  assign new_C8672_ = ~new_C8617_ & new_C8631_;
  assign new_C8673_ = new_C8677_ | new_C8678_;
  assign new_C8674_ = new_C8617_ & new_C8631_;
  assign new_C8675_ = ~new_C8617_ & ~new_C8631_;
  assign new_C8676_ = new_C8617_ & ~new_C8631_;
  assign new_C8677_ = new_C8617_ & ~new_C8631_;
  assign new_C8678_ = ~new_C8617_ & new_C8631_;
  assign new_C8679_ = new_E5037_;
  assign new_C8680_ = new_E5104_;
  assign new_C8681_ = new_E5171_;
  assign new_C8682_ = new_E5238_;
  assign new_C8683_ = new_E5305_;
  assign new_C8684_ = new_E5372_;
  assign new_C8685_ = new_C8692_ & new_C8691_;
  assign new_C8686_ = new_C8694_ | new_C8693_;
  assign new_C8687_ = new_C8696_ | new_C8695_;
  assign new_C8688_ = new_C8698_ & new_C8697_;
  assign new_C8689_ = new_C8698_ & new_C8699_;
  assign new_C8690_ = new_C8691_ | new_C8700_;
  assign new_C8691_ = new_C8680_ | new_C8703_;
  assign new_C8692_ = new_C8702_ | new_C8701_;
  assign new_C8693_ = new_C8707_ & new_C8706_;
  assign new_C8694_ = new_C8705_ & new_C8704_;
  assign new_C8695_ = new_C8710_ | new_C8709_;
  assign new_C8696_ = new_C8705_ & new_C8708_;
  assign new_C8697_ = new_C8680_ | new_C8713_;
  assign new_C8698_ = new_C8712_ | new_C8711_;
  assign new_C8699_ = new_C8715_ | new_C8714_;
  assign new_C8700_ = ~new_C8691_ & new_C8717_;
  assign new_C8701_ = ~new_C8693_ & new_C8705_;
  assign new_C8702_ = new_C8693_ & ~new_C8705_;
  assign new_C8703_ = new_C8679_ & ~new_C8680_;
  assign new_C8704_ = ~new_C8726_ | ~new_C8727_;
  assign new_C8705_ = new_C8719_ | new_C8721_;
  assign new_C8706_ = new_C8729_ | new_C8728_;
  assign new_C8707_ = new_C8723_ | new_C8722_;
  assign new_C8708_ = ~new_C8731_ | ~new_C8730_;
  assign new_C8709_ = ~new_C8732_ & new_C8733_;
  assign new_C8710_ = new_C8732_ & ~new_C8733_;
  assign new_C8711_ = ~new_C8679_ & new_C8680_;
  assign new_C8712_ = new_C8679_ & ~new_C8680_;
  assign new_C8713_ = ~new_C8695_ | new_C8705_;
  assign new_C8714_ = new_C8695_ & new_C8705_;
  assign new_C8715_ = ~new_C8695_ & ~new_C8705_;
  assign new_C8716_ = new_C8737_ | new_C8736_;
  assign new_C8717_ = new_C8683_ | new_C8716_;
  assign new_C8718_ = new_C8741_ | new_C8740_;
  assign new_C8719_ = ~new_C8683_ & new_C8718_;
  assign new_C8720_ = new_C8739_ | new_C8738_;
  assign new_C8721_ = new_C8683_ & new_C8720_;
  assign new_C8722_ = new_C8681_ & ~new_C8691_;
  assign new_C8723_ = ~new_C8681_ & new_C8691_;
  assign new_C8724_ = ~new_C8680_ | ~new_C8705_;
  assign new_C8725_ = new_C8691_ & new_C8724_;
  assign new_C8726_ = ~new_C8691_ & ~new_C8725_;
  assign new_C8727_ = new_C8691_ | new_C8724_;
  assign new_C8728_ = ~new_C8681_ & new_C8682_;
  assign new_C8729_ = new_C8681_ & ~new_C8682_;
  assign new_C8730_ = new_C8698_ | new_C8735_;
  assign new_C8731_ = ~new_C8698_ & ~new_C8734_;
  assign new_C8732_ = new_C8681_ | new_C8698_;
  assign new_C8733_ = new_C8681_ | new_C8682_;
  assign new_C8734_ = new_C8698_ & new_C8735_;
  assign new_C8735_ = ~new_C8680_ | ~new_C8705_;
  assign new_C8736_ = new_C8713_ & new_C8733_;
  assign new_C8737_ = ~new_C8713_ & ~new_C8733_;
  assign new_C8738_ = new_C8742_ | new_C8743_;
  assign new_C8739_ = ~new_C8684_ & new_C8698_;
  assign new_C8740_ = new_C8744_ | new_C8745_;
  assign new_C8741_ = new_C8684_ & new_C8698_;
  assign new_C8742_ = ~new_C8684_ & ~new_C8698_;
  assign new_C8743_ = new_C8684_ & ~new_C8698_;
  assign new_C8744_ = new_C8684_ & ~new_C8698_;
  assign new_C8745_ = ~new_C8684_ & new_C8698_;
  assign new_C8746_ = new_E5439_;
  assign new_C8747_ = new_E5506_;
  assign new_C8748_ = new_E5573_;
  assign new_C8749_ = new_E5640_;
  assign new_C8750_ = new_E5707_;
  assign new_C8751_ = new_E5774_;
  assign new_C8752_ = new_C8759_ & new_C8758_;
  assign new_C8753_ = new_C8761_ | new_C8760_;
  assign new_C8754_ = new_C8763_ | new_C8762_;
  assign new_C8755_ = new_C8765_ & new_C8764_;
  assign new_C8756_ = new_C8765_ & new_C8766_;
  assign new_C8757_ = new_C8758_ | new_C8767_;
  assign new_C8758_ = new_C8747_ | new_C8770_;
  assign new_C8759_ = new_C8769_ | new_C8768_;
  assign new_C8760_ = new_C8774_ & new_C8773_;
  assign new_C8761_ = new_C8772_ & new_C8771_;
  assign new_C8762_ = new_C8777_ | new_C8776_;
  assign new_C8763_ = new_C8772_ & new_C8775_;
  assign new_C8764_ = new_C8747_ | new_C8780_;
  assign new_C8765_ = new_C8779_ | new_C8778_;
  assign new_C8766_ = new_C8782_ | new_C8781_;
  assign new_C8767_ = ~new_C8758_ & new_C8784_;
  assign new_C8768_ = ~new_C8760_ & new_C8772_;
  assign new_C8769_ = new_C8760_ & ~new_C8772_;
  assign new_C8770_ = new_C8746_ & ~new_C8747_;
  assign new_C8771_ = ~new_C8793_ | ~new_C8794_;
  assign new_C8772_ = new_C8786_ | new_C8788_;
  assign new_C8773_ = new_C8796_ | new_C8795_;
  assign new_C8774_ = new_C8790_ | new_C8789_;
  assign new_C8775_ = ~new_C8798_ | ~new_C8797_;
  assign new_C8776_ = ~new_C8799_ & new_C8800_;
  assign new_C8777_ = new_C8799_ & ~new_C8800_;
  assign new_C8778_ = ~new_C8746_ & new_C8747_;
  assign new_C8779_ = new_C8746_ & ~new_C8747_;
  assign new_C8780_ = ~new_C8762_ | new_C8772_;
  assign new_C8781_ = new_C8762_ & new_C8772_;
  assign new_C8782_ = ~new_C8762_ & ~new_C8772_;
  assign new_C8783_ = new_C8804_ | new_C8803_;
  assign new_C8784_ = new_C8750_ | new_C8783_;
  assign new_C8785_ = new_C8808_ | new_C8807_;
  assign new_C8786_ = ~new_C8750_ & new_C8785_;
  assign new_C8787_ = new_C8806_ | new_C8805_;
  assign new_C8788_ = new_C8750_ & new_C8787_;
  assign new_C8789_ = new_C8748_ & ~new_C8758_;
  assign new_C8790_ = ~new_C8748_ & new_C8758_;
  assign new_C8791_ = ~new_C8747_ | ~new_C8772_;
  assign new_C8792_ = new_C8758_ & new_C8791_;
  assign new_C8793_ = ~new_C8758_ & ~new_C8792_;
  assign new_C8794_ = new_C8758_ | new_C8791_;
  assign new_C8795_ = ~new_C8748_ & new_C8749_;
  assign new_C8796_ = new_C8748_ & ~new_C8749_;
  assign new_C8797_ = new_C8765_ | new_C8802_;
  assign new_C8798_ = ~new_C8765_ & ~new_C8801_;
  assign new_C8799_ = new_C8748_ | new_C8765_;
  assign new_C8800_ = new_C8748_ | new_C8749_;
  assign new_C8801_ = new_C8765_ & new_C8802_;
  assign new_C8802_ = ~new_C8747_ | ~new_C8772_;
  assign new_C8803_ = new_C8780_ & new_C8800_;
  assign new_C8804_ = ~new_C8780_ & ~new_C8800_;
  assign new_C8805_ = new_C8809_ | new_C8810_;
  assign new_C8806_ = ~new_C8751_ & new_C8765_;
  assign new_C8807_ = new_C8811_ | new_C8812_;
  assign new_C8808_ = new_C8751_ & new_C8765_;
  assign new_C8809_ = ~new_C8751_ & ~new_C8765_;
  assign new_C8810_ = new_C8751_ & ~new_C8765_;
  assign new_C8811_ = new_C8751_ & ~new_C8765_;
  assign new_C8812_ = ~new_C8751_ & new_C8765_;
  assign new_C8813_ = new_E5841_;
  assign new_C8814_ = new_E5908_;
  assign new_C8815_ = new_E5975_;
  assign new_C8816_ = new_E6042_;
  assign new_C8817_ = new_E6109_;
  assign new_C8818_ = new_E6176_;
  assign new_C8819_ = new_C8826_ & new_C8825_;
  assign new_C8820_ = new_C8828_ | new_C8827_;
  assign new_C8821_ = new_C8830_ | new_C8829_;
  assign new_C8822_ = new_C8832_ & new_C8831_;
  assign new_C8823_ = new_C8832_ & new_C8833_;
  assign new_C8824_ = new_C8825_ | new_C8834_;
  assign new_C8825_ = new_C8814_ | new_C8837_;
  assign new_C8826_ = new_C8836_ | new_C8835_;
  assign new_C8827_ = new_C8841_ & new_C8840_;
  assign new_C8828_ = new_C8839_ & new_C8838_;
  assign new_C8829_ = new_C8844_ | new_C8843_;
  assign new_C8830_ = new_C8839_ & new_C8842_;
  assign new_C8831_ = new_C8814_ | new_C8847_;
  assign new_C8832_ = new_C8846_ | new_C8845_;
  assign new_C8833_ = new_C8849_ | new_C8848_;
  assign new_C8834_ = ~new_C8825_ & new_C8851_;
  assign new_C8835_ = ~new_C8827_ & new_C8839_;
  assign new_C8836_ = new_C8827_ & ~new_C8839_;
  assign new_C8837_ = new_C8813_ & ~new_C8814_;
  assign new_C8838_ = ~new_C8860_ | ~new_C8861_;
  assign new_C8839_ = new_C8853_ | new_C8855_;
  assign new_C8840_ = new_C8863_ | new_C8862_;
  assign new_C8841_ = new_C8857_ | new_C8856_;
  assign new_C8842_ = ~new_C8865_ | ~new_C8864_;
  assign new_C8843_ = ~new_C8866_ & new_C8867_;
  assign new_C8844_ = new_C8866_ & ~new_C8867_;
  assign new_C8845_ = ~new_C8813_ & new_C8814_;
  assign new_C8846_ = new_C8813_ & ~new_C8814_;
  assign new_C8847_ = ~new_C8829_ | new_C8839_;
  assign new_C8848_ = new_C8829_ & new_C8839_;
  assign new_C8849_ = ~new_C8829_ & ~new_C8839_;
  assign new_C8850_ = new_C8871_ | new_C8870_;
  assign new_C8851_ = new_C8817_ | new_C8850_;
  assign new_C8852_ = new_C8875_ | new_C8874_;
  assign new_C8853_ = ~new_C8817_ & new_C8852_;
  assign new_C8854_ = new_C8873_ | new_C8872_;
  assign new_C8855_ = new_C8817_ & new_C8854_;
  assign new_C8856_ = new_C8815_ & ~new_C8825_;
  assign new_C8857_ = ~new_C8815_ & new_C8825_;
  assign new_C8858_ = ~new_C8814_ | ~new_C8839_;
  assign new_C8859_ = new_C8825_ & new_C8858_;
  assign new_C8860_ = ~new_C8825_ & ~new_C8859_;
  assign new_C8861_ = new_C8825_ | new_C8858_;
  assign new_C8862_ = ~new_C8815_ & new_C8816_;
  assign new_C8863_ = new_C8815_ & ~new_C8816_;
  assign new_C8864_ = new_C8832_ | new_C8869_;
  assign new_C8865_ = ~new_C8832_ & ~new_C8868_;
  assign new_C8866_ = new_C8815_ | new_C8832_;
  assign new_C8867_ = new_C8815_ | new_C8816_;
  assign new_C8868_ = new_C8832_ & new_C8869_;
  assign new_C8869_ = ~new_C8814_ | ~new_C8839_;
  assign new_C8870_ = new_C8847_ & new_C8867_;
  assign new_C8871_ = ~new_C8847_ & ~new_C8867_;
  assign new_C8872_ = new_C8876_ | new_C8877_;
  assign new_C8873_ = ~new_C8818_ & new_C8832_;
  assign new_C8874_ = new_C8878_ | new_C8879_;
  assign new_C8875_ = new_C8818_ & new_C8832_;
  assign new_C8876_ = ~new_C8818_ & ~new_C8832_;
  assign new_C8877_ = new_C8818_ & ~new_C8832_;
  assign new_C8878_ = new_C8818_ & ~new_C8832_;
  assign new_C8879_ = ~new_C8818_ & new_C8832_;
  assign new_C8880_ = new_E6243_;
  assign new_C8881_ = new_E6310_;
  assign new_C8882_ = new_E6377_;
  assign new_C8883_ = new_E6444_;
  assign new_C8884_ = new_E6511_;
  assign new_C8885_ = new_E6578_;
  assign new_C8886_ = new_C8893_ & new_C8892_;
  assign new_C8887_ = new_C8895_ | new_C8894_;
  assign new_C8888_ = new_C8897_ | new_C8896_;
  assign new_C8889_ = new_C8899_ & new_C8898_;
  assign new_C8890_ = new_C8899_ & new_C8900_;
  assign new_C8891_ = new_C8892_ | new_C8901_;
  assign new_C8892_ = new_C8881_ | new_C8904_;
  assign new_C8893_ = new_C8903_ | new_C8902_;
  assign new_C8894_ = new_C8908_ & new_C8907_;
  assign new_C8895_ = new_C8906_ & new_C8905_;
  assign new_C8896_ = new_C8911_ | new_C8910_;
  assign new_C8897_ = new_C8906_ & new_C8909_;
  assign new_C8898_ = new_C8881_ | new_C8914_;
  assign new_C8899_ = new_C8913_ | new_C8912_;
  assign new_C8900_ = new_C8916_ | new_C8915_;
  assign new_C8901_ = ~new_C8892_ & new_C8918_;
  assign new_C8902_ = ~new_C8894_ & new_C8906_;
  assign new_C8903_ = new_C8894_ & ~new_C8906_;
  assign new_C8904_ = new_C8880_ & ~new_C8881_;
  assign new_C8905_ = ~new_C8927_ | ~new_C8928_;
  assign new_C8906_ = new_C8920_ | new_C8922_;
  assign new_C8907_ = new_C8930_ | new_C8929_;
  assign new_C8908_ = new_C8924_ | new_C8923_;
  assign new_C8909_ = ~new_C8932_ | ~new_C8931_;
  assign new_C8910_ = ~new_C8933_ & new_C8934_;
  assign new_C8911_ = new_C8933_ & ~new_C8934_;
  assign new_C8912_ = ~new_C8880_ & new_C8881_;
  assign new_C8913_ = new_C8880_ & ~new_C8881_;
  assign new_C8914_ = ~new_C8896_ | new_C8906_;
  assign new_C8915_ = new_C8896_ & new_C8906_;
  assign new_C8916_ = ~new_C8896_ & ~new_C8906_;
  assign new_C8917_ = new_C8938_ | new_C8937_;
  assign new_C8918_ = new_C8884_ | new_C8917_;
  assign new_C8919_ = new_C8942_ | new_C8941_;
  assign new_C8920_ = ~new_C8884_ & new_C8919_;
  assign new_C8921_ = new_C8940_ | new_C8939_;
  assign new_C8922_ = new_C8884_ & new_C8921_;
  assign new_C8923_ = new_C8882_ & ~new_C8892_;
  assign new_C8924_ = ~new_C8882_ & new_C8892_;
  assign new_C8925_ = ~new_C8881_ | ~new_C8906_;
  assign new_C8926_ = new_C8892_ & new_C8925_;
  assign new_C8927_ = ~new_C8892_ & ~new_C8926_;
  assign new_C8928_ = new_C8892_ | new_C8925_;
  assign new_C8929_ = ~new_C8882_ & new_C8883_;
  assign new_C8930_ = new_C8882_ & ~new_C8883_;
  assign new_C8931_ = new_C8899_ | new_C8936_;
  assign new_C8932_ = ~new_C8899_ & ~new_C8935_;
  assign new_C8933_ = new_C8882_ | new_C8899_;
  assign new_C8934_ = new_C8882_ | new_C8883_;
  assign new_C8935_ = new_C8899_ & new_C8936_;
  assign new_C8936_ = ~new_C8881_ | ~new_C8906_;
  assign new_C8937_ = new_C8914_ & new_C8934_;
  assign new_C8938_ = ~new_C8914_ & ~new_C8934_;
  assign new_C8939_ = new_C8943_ | new_C8944_;
  assign new_C8940_ = ~new_C8885_ & new_C8899_;
  assign new_C8941_ = new_C8945_ | new_C8946_;
  assign new_C8942_ = new_C8885_ & new_C8899_;
  assign new_C8943_ = ~new_C8885_ & ~new_C8899_;
  assign new_C8944_ = new_C8885_ & ~new_C8899_;
  assign new_C8945_ = new_C8885_ & ~new_C8899_;
  assign new_C8946_ = ~new_C8885_ & new_C8899_;
  assign new_C8947_ = new_E6645_;
  assign new_C8948_ = new_E6712_;
  assign new_C8949_ = new_E6779_;
  assign new_C8950_ = new_E6846_;
  assign new_C8951_ = new_E6913_;
  assign new_C8952_ = new_E6980_;
  assign new_C8953_ = new_C8960_ & new_C8959_;
  assign new_C8954_ = new_C8962_ | new_C8961_;
  assign new_C8955_ = new_C8964_ | new_C8963_;
  assign new_C8956_ = new_C8966_ & new_C8965_;
  assign new_C8957_ = new_C8966_ & new_C8967_;
  assign new_C8958_ = new_C8959_ | new_C8968_;
  assign new_C8959_ = new_C8948_ | new_C8971_;
  assign new_C8960_ = new_C8970_ | new_C8969_;
  assign new_C8961_ = new_C8975_ & new_C8974_;
  assign new_C8962_ = new_C8973_ & new_C8972_;
  assign new_C8963_ = new_C8978_ | new_C8977_;
  assign new_C8964_ = new_C8973_ & new_C8976_;
  assign new_C8965_ = new_C8948_ | new_C8981_;
  assign new_C8966_ = new_C8980_ | new_C8979_;
  assign new_C8967_ = new_C8983_ | new_C8982_;
  assign new_C8968_ = ~new_C8959_ & new_C8985_;
  assign new_C8969_ = ~new_C8961_ & new_C8973_;
  assign new_C8970_ = new_C8961_ & ~new_C8973_;
  assign new_C8971_ = new_C8947_ & ~new_C8948_;
  assign new_C8972_ = ~new_C8994_ | ~new_C8995_;
  assign new_C8973_ = new_C8987_ | new_C8989_;
  assign new_C8974_ = new_C8997_ | new_C8996_;
  assign new_C8975_ = new_C8991_ | new_C8990_;
  assign new_C8976_ = ~new_C8999_ | ~new_C8998_;
  assign new_C8977_ = ~new_C9000_ & new_C9001_;
  assign new_C8978_ = new_C9000_ & ~new_C9001_;
  assign new_C8979_ = ~new_C8947_ & new_C8948_;
  assign new_C8980_ = new_C8947_ & ~new_C8948_;
  assign new_C8981_ = ~new_C8963_ | new_C8973_;
  assign new_C8982_ = new_C8963_ & new_C8973_;
  assign new_C8983_ = ~new_C8963_ & ~new_C8973_;
  assign new_C8984_ = new_C9005_ | new_C9004_;
  assign new_C8985_ = new_C8951_ | new_C8984_;
  assign new_C8986_ = new_C9009_ | new_C9008_;
  assign new_C8987_ = ~new_C8951_ & new_C8986_;
  assign new_C8988_ = new_C9007_ | new_C9006_;
  assign new_C8989_ = new_C8951_ & new_C8988_;
  assign new_C8990_ = new_C8949_ & ~new_C8959_;
  assign new_C8991_ = ~new_C8949_ & new_C8959_;
  assign new_C8992_ = ~new_C8948_ | ~new_C8973_;
  assign new_C8993_ = new_C8959_ & new_C8992_;
  assign new_C8994_ = ~new_C8959_ & ~new_C8993_;
  assign new_C8995_ = new_C8959_ | new_C8992_;
  assign new_C8996_ = ~new_C8949_ & new_C8950_;
  assign new_C8997_ = new_C8949_ & ~new_C8950_;
  assign new_C8998_ = new_C8966_ | new_C9003_;
  assign new_C8999_ = ~new_C8966_ & ~new_C9002_;
  assign new_C9000_ = new_C8949_ | new_C8966_;
  assign new_C9001_ = new_C8949_ | new_C8950_;
  assign new_C9002_ = new_C8966_ & new_C9003_;
  assign new_C9003_ = ~new_C8948_ | ~new_C8973_;
  assign new_C9004_ = new_C8981_ & new_C9001_;
  assign new_C9005_ = ~new_C8981_ & ~new_C9001_;
  assign new_C9006_ = new_C9010_ | new_C9011_;
  assign new_C9007_ = ~new_C8952_ & new_C8966_;
  assign new_C9008_ = new_C9012_ | new_C9013_;
  assign new_C9009_ = new_C8952_ & new_C8966_;
  assign new_C9010_ = ~new_C8952_ & ~new_C8966_;
  assign new_C9011_ = new_C8952_ & ~new_C8966_;
  assign new_C9012_ = new_C8952_ & ~new_C8966_;
  assign new_C9013_ = ~new_C8952_ & new_C8966_;
  assign new_C9014_ = new_E7047_;
  assign new_C9015_ = new_E7114_;
  assign new_C9016_ = new_E7181_;
  assign new_C9017_ = new_E7248_;
  assign new_C9018_ = new_E7315_;
  assign new_C9019_ = new_E7382_;
  assign new_C9020_ = new_C9027_ & new_C9026_;
  assign new_C9021_ = new_C9029_ | new_C9028_;
  assign new_C9022_ = new_C9031_ | new_C9030_;
  assign new_C9023_ = new_C9033_ & new_C9032_;
  assign new_C9024_ = new_C9033_ & new_C9034_;
  assign new_C9025_ = new_C9026_ | new_C9035_;
  assign new_C9026_ = new_C9015_ | new_C9038_;
  assign new_C9027_ = new_C9037_ | new_C9036_;
  assign new_C9028_ = new_C9042_ & new_C9041_;
  assign new_C9029_ = new_C9040_ & new_C9039_;
  assign new_C9030_ = new_C9045_ | new_C9044_;
  assign new_C9031_ = new_C9040_ & new_C9043_;
  assign new_C9032_ = new_C9015_ | new_C9048_;
  assign new_C9033_ = new_C9047_ | new_C9046_;
  assign new_C9034_ = new_C9050_ | new_C9049_;
  assign new_C9035_ = ~new_C9026_ & new_C9052_;
  assign new_C9036_ = ~new_C9028_ & new_C9040_;
  assign new_C9037_ = new_C9028_ & ~new_C9040_;
  assign new_C9038_ = new_C9014_ & ~new_C9015_;
  assign new_C9039_ = ~new_C9061_ | ~new_C9062_;
  assign new_C9040_ = new_C9054_ | new_C9056_;
  assign new_C9041_ = new_C9064_ | new_C9063_;
  assign new_C9042_ = new_C9058_ | new_C9057_;
  assign new_C9043_ = ~new_C9066_ | ~new_C9065_;
  assign new_C9044_ = ~new_C9067_ & new_C9068_;
  assign new_C9045_ = new_C9067_ & ~new_C9068_;
  assign new_C9046_ = ~new_C9014_ & new_C9015_;
  assign new_C9047_ = new_C9014_ & ~new_C9015_;
  assign new_C9048_ = ~new_C9030_ | new_C9040_;
  assign new_C9049_ = new_C9030_ & new_C9040_;
  assign new_C9050_ = ~new_C9030_ & ~new_C9040_;
  assign new_C9051_ = new_C9072_ | new_C9071_;
  assign new_C9052_ = new_C9018_ | new_C9051_;
  assign new_C9053_ = new_C9076_ | new_C9075_;
  assign new_C9054_ = ~new_C9018_ & new_C9053_;
  assign new_C9055_ = new_C9074_ | new_C9073_;
  assign new_C9056_ = new_C9018_ & new_C9055_;
  assign new_C9057_ = new_C9016_ & ~new_C9026_;
  assign new_C9058_ = ~new_C9016_ & new_C9026_;
  assign new_C9059_ = ~new_C9015_ | ~new_C9040_;
  assign new_C9060_ = new_C9026_ & new_C9059_;
  assign new_C9061_ = ~new_C9026_ & ~new_C9060_;
  assign new_C9062_ = new_C9026_ | new_C9059_;
  assign new_C9063_ = ~new_C9016_ & new_C9017_;
  assign new_C9064_ = new_C9016_ & ~new_C9017_;
  assign new_C9065_ = new_C9033_ | new_C9070_;
  assign new_C9066_ = ~new_C9033_ & ~new_C9069_;
  assign new_C9067_ = new_C9016_ | new_C9033_;
  assign new_C9068_ = new_C9016_ | new_C9017_;
  assign new_C9069_ = new_C9033_ & new_C9070_;
  assign new_C9070_ = ~new_C9015_ | ~new_C9040_;
  assign new_C9071_ = new_C9048_ & new_C9068_;
  assign new_C9072_ = ~new_C9048_ & ~new_C9068_;
  assign new_C9073_ = new_C9077_ | new_C9078_;
  assign new_C9074_ = ~new_C9019_ & new_C9033_;
  assign new_C9075_ = new_C9079_ | new_C9080_;
  assign new_C9076_ = new_C9019_ & new_C9033_;
  assign new_C9077_ = ~new_C9019_ & ~new_C9033_;
  assign new_C9078_ = new_C9019_ & ~new_C9033_;
  assign new_C9079_ = new_C9019_ & ~new_C9033_;
  assign new_C9080_ = ~new_C9019_ & new_C9033_;
  assign new_C9081_ = new_E7449_;
  assign new_C9082_ = new_E7516_;
  assign new_C9083_ = new_E7583_;
  assign new_C9084_ = new_E7650_;
  assign new_C9085_ = new_E7717_;
  assign new_C9086_ = new_E7784_;
  assign new_C9087_ = new_C9094_ & new_C9093_;
  assign new_C9088_ = new_C9096_ | new_C9095_;
  assign new_C9089_ = new_C9098_ | new_C9097_;
  assign new_C9090_ = new_C9100_ & new_C9099_;
  assign new_C9091_ = new_C9100_ & new_C9101_;
  assign new_C9092_ = new_C9093_ | new_C9102_;
  assign new_C9093_ = new_C9082_ | new_C9105_;
  assign new_C9094_ = new_C9104_ | new_C9103_;
  assign new_C9095_ = new_C9109_ & new_C9108_;
  assign new_C9096_ = new_C9107_ & new_C9106_;
  assign new_C9097_ = new_C9112_ | new_C9111_;
  assign new_C9098_ = new_C9107_ & new_C9110_;
  assign new_C9099_ = new_C9082_ | new_C9115_;
  assign new_C9100_ = new_C9114_ | new_C9113_;
  assign new_C9101_ = new_C9117_ | new_C9116_;
  assign new_C9102_ = ~new_C9093_ & new_C9119_;
  assign new_C9103_ = ~new_C9095_ & new_C9107_;
  assign new_C9104_ = new_C9095_ & ~new_C9107_;
  assign new_C9105_ = new_C9081_ & ~new_C9082_;
  assign new_C9106_ = ~new_C9128_ | ~new_C9129_;
  assign new_C9107_ = new_C9121_ | new_C9123_;
  assign new_C9108_ = new_C9131_ | new_C9130_;
  assign new_C9109_ = new_C9125_ | new_C9124_;
  assign new_C9110_ = ~new_C9133_ | ~new_C9132_;
  assign new_C9111_ = ~new_C9134_ & new_C9135_;
  assign new_C9112_ = new_C9134_ & ~new_C9135_;
  assign new_C9113_ = ~new_C9081_ & new_C9082_;
  assign new_C9114_ = new_C9081_ & ~new_C9082_;
  assign new_C9115_ = ~new_C9097_ | new_C9107_;
  assign new_C9116_ = new_C9097_ & new_C9107_;
  assign new_C9117_ = ~new_C9097_ & ~new_C9107_;
  assign new_C9118_ = new_C9139_ | new_C9138_;
  assign new_C9119_ = new_C9085_ | new_C9118_;
  assign new_C9120_ = new_C9143_ | new_C9142_;
  assign new_C9121_ = ~new_C9085_ & new_C9120_;
  assign new_C9122_ = new_C9141_ | new_C9140_;
  assign new_C9123_ = new_C9085_ & new_C9122_;
  assign new_C9124_ = new_C9083_ & ~new_C9093_;
  assign new_C9125_ = ~new_C9083_ & new_C9093_;
  assign new_C9126_ = ~new_C9082_ | ~new_C9107_;
  assign new_C9127_ = new_C9093_ & new_C9126_;
  assign new_C9128_ = ~new_C9093_ & ~new_C9127_;
  assign new_C9129_ = new_C9093_ | new_C9126_;
  assign new_C9130_ = ~new_C9083_ & new_C9084_;
  assign new_C9131_ = new_C9083_ & ~new_C9084_;
  assign new_C9132_ = new_C9100_ | new_C9137_;
  assign new_C9133_ = ~new_C9100_ & ~new_C9136_;
  assign new_C9134_ = new_C9083_ | new_C9100_;
  assign new_C9135_ = new_C9083_ | new_C9084_;
  assign new_C9136_ = new_C9100_ & new_C9137_;
  assign new_C9137_ = ~new_C9082_ | ~new_C9107_;
  assign new_C9138_ = new_C9115_ & new_C9135_;
  assign new_C9139_ = ~new_C9115_ & ~new_C9135_;
  assign new_C9140_ = new_C9144_ | new_C9145_;
  assign new_C9141_ = ~new_C9086_ & new_C9100_;
  assign new_C9142_ = new_C9146_ | new_C9147_;
  assign new_C9143_ = new_C9086_ & new_C9100_;
  assign new_C9144_ = ~new_C9086_ & ~new_C9100_;
  assign new_C9145_ = new_C9086_ & ~new_C9100_;
  assign new_C9146_ = new_C9086_ & ~new_C9100_;
  assign new_C9147_ = ~new_C9086_ & new_C9100_;
  assign new_C9148_ = new_E7851_;
  assign new_C9149_ = new_E7918_;
  assign new_C9150_ = new_E7985_;
  assign new_C9151_ = new_E8052_;
  assign new_C9152_ = new_E8119_;
  assign new_C9153_ = new_E8186_;
  assign new_C9154_ = new_C9161_ & new_C9160_;
  assign new_C9155_ = new_C9163_ | new_C9162_;
  assign new_C9156_ = new_C9165_ | new_C9164_;
  assign new_C9157_ = new_C9167_ & new_C9166_;
  assign new_C9158_ = new_C9167_ & new_C9168_;
  assign new_C9159_ = new_C9160_ | new_C9169_;
  assign new_C9160_ = new_C9149_ | new_C9172_;
  assign new_C9161_ = new_C9171_ | new_C9170_;
  assign new_C9162_ = new_C9176_ & new_C9175_;
  assign new_C9163_ = new_C9174_ & new_C9173_;
  assign new_C9164_ = new_C9179_ | new_C9178_;
  assign new_C9165_ = new_C9174_ & new_C9177_;
  assign new_C9166_ = new_C9149_ | new_C9182_;
  assign new_C9167_ = new_C9181_ | new_C9180_;
  assign new_C9168_ = new_C9184_ | new_C9183_;
  assign new_C9169_ = ~new_C9160_ & new_C9186_;
  assign new_C9170_ = ~new_C9162_ & new_C9174_;
  assign new_C9171_ = new_C9162_ & ~new_C9174_;
  assign new_C9172_ = new_C9148_ & ~new_C9149_;
  assign new_C9173_ = ~new_C9195_ | ~new_C9196_;
  assign new_C9174_ = new_C9188_ | new_C9190_;
  assign new_C9175_ = new_C9198_ | new_C9197_;
  assign new_C9176_ = new_C9192_ | new_C9191_;
  assign new_C9177_ = ~new_C9200_ | ~new_C9199_;
  assign new_C9178_ = ~new_C9201_ & new_C9202_;
  assign new_C9179_ = new_C9201_ & ~new_C9202_;
  assign new_C9180_ = ~new_C9148_ & new_C9149_;
  assign new_C9181_ = new_C9148_ & ~new_C9149_;
  assign new_C9182_ = ~new_C9164_ | new_C9174_;
  assign new_C9183_ = new_C9164_ & new_C9174_;
  assign new_C9184_ = ~new_C9164_ & ~new_C9174_;
  assign new_C9185_ = new_C9206_ | new_C9205_;
  assign new_C9186_ = new_C9152_ | new_C9185_;
  assign new_C9187_ = new_C9210_ | new_C9209_;
  assign new_C9188_ = ~new_C9152_ & new_C9187_;
  assign new_C9189_ = new_C9208_ | new_C9207_;
  assign new_C9190_ = new_C9152_ & new_C9189_;
  assign new_C9191_ = new_C9150_ & ~new_C9160_;
  assign new_C9192_ = ~new_C9150_ & new_C9160_;
  assign new_C9193_ = ~new_C9149_ | ~new_C9174_;
  assign new_C9194_ = new_C9160_ & new_C9193_;
  assign new_C9195_ = ~new_C9160_ & ~new_C9194_;
  assign new_C9196_ = new_C9160_ | new_C9193_;
  assign new_C9197_ = ~new_C9150_ & new_C9151_;
  assign new_C9198_ = new_C9150_ & ~new_C9151_;
  assign new_C9199_ = new_C9167_ | new_C9204_;
  assign new_C9200_ = ~new_C9167_ & ~new_C9203_;
  assign new_C9201_ = new_C9150_ | new_C9167_;
  assign new_C9202_ = new_C9150_ | new_C9151_;
  assign new_C9203_ = new_C9167_ & new_C9204_;
  assign new_C9204_ = ~new_C9149_ | ~new_C9174_;
  assign new_C9205_ = new_C9182_ & new_C9202_;
  assign new_C9206_ = ~new_C9182_ & ~new_C9202_;
  assign new_C9207_ = new_C9211_ | new_C9212_;
  assign new_C9208_ = ~new_C9153_ & new_C9167_;
  assign new_C9209_ = new_C9213_ | new_C9214_;
  assign new_C9210_ = new_C9153_ & new_C9167_;
  assign new_C9211_ = ~new_C9153_ & ~new_C9167_;
  assign new_C9212_ = new_C9153_ & ~new_C9167_;
  assign new_C9213_ = new_C9153_ & ~new_C9167_;
  assign new_C9214_ = ~new_C9153_ & new_C9167_;
  assign new_C9215_ = new_E8253_;
  assign new_C9216_ = new_E8320_;
  assign new_C9217_ = new_E8387_;
  assign new_C9218_ = new_E8454_;
  assign new_C9219_ = new_E8521_;
  assign new_C9220_ = new_E8588_;
  assign new_C9221_ = new_C9228_ & new_C9227_;
  assign new_C9222_ = new_C9230_ | new_C9229_;
  assign new_C9223_ = new_C9232_ | new_C9231_;
  assign new_C9224_ = new_C9234_ & new_C9233_;
  assign new_C9225_ = new_C9234_ & new_C9235_;
  assign new_C9226_ = new_C9227_ | new_C9236_;
  assign new_C9227_ = new_C9216_ | new_C9239_;
  assign new_C9228_ = new_C9238_ | new_C9237_;
  assign new_C9229_ = new_C9243_ & new_C9242_;
  assign new_C9230_ = new_C9241_ & new_C9240_;
  assign new_C9231_ = new_C9246_ | new_C9245_;
  assign new_C9232_ = new_C9241_ & new_C9244_;
  assign new_C9233_ = new_C9216_ | new_C9249_;
  assign new_C9234_ = new_C9248_ | new_C9247_;
  assign new_C9235_ = new_C9251_ | new_C9250_;
  assign new_C9236_ = ~new_C9227_ & new_C9253_;
  assign new_C9237_ = ~new_C9229_ & new_C9241_;
  assign new_C9238_ = new_C9229_ & ~new_C9241_;
  assign new_C9239_ = new_C9215_ & ~new_C9216_;
  assign new_C9240_ = ~new_C9262_ | ~new_C9263_;
  assign new_C9241_ = new_C9255_ | new_C9257_;
  assign new_C9242_ = new_C9265_ | new_C9264_;
  assign new_C9243_ = new_C9259_ | new_C9258_;
  assign new_C9244_ = ~new_C9267_ | ~new_C9266_;
  assign new_C9245_ = ~new_C9268_ & new_C9269_;
  assign new_C9246_ = new_C9268_ & ~new_C9269_;
  assign new_C9247_ = ~new_C9215_ & new_C9216_;
  assign new_C9248_ = new_C9215_ & ~new_C9216_;
  assign new_C9249_ = ~new_C9231_ | new_C9241_;
  assign new_C9250_ = new_C9231_ & new_C9241_;
  assign new_C9251_ = ~new_C9231_ & ~new_C9241_;
  assign new_C9252_ = new_C9273_ | new_C9272_;
  assign new_C9253_ = new_C9219_ | new_C9252_;
  assign new_C9254_ = new_C9277_ | new_C9276_;
  assign new_C9255_ = ~new_C9219_ & new_C9254_;
  assign new_C9256_ = new_C9275_ | new_C9274_;
  assign new_C9257_ = new_C9219_ & new_C9256_;
  assign new_C9258_ = new_C9217_ & ~new_C9227_;
  assign new_C9259_ = ~new_C9217_ & new_C9227_;
  assign new_C9260_ = ~new_C9216_ | ~new_C9241_;
  assign new_C9261_ = new_C9227_ & new_C9260_;
  assign new_C9262_ = ~new_C9227_ & ~new_C9261_;
  assign new_C9263_ = new_C9227_ | new_C9260_;
  assign new_C9264_ = ~new_C9217_ & new_C9218_;
  assign new_C9265_ = new_C9217_ & ~new_C9218_;
  assign new_C9266_ = new_C9234_ | new_C9271_;
  assign new_C9267_ = ~new_C9234_ & ~new_C9270_;
  assign new_C9268_ = new_C9217_ | new_C9234_;
  assign new_C9269_ = new_C9217_ | new_C9218_;
  assign new_C9270_ = new_C9234_ & new_C9271_;
  assign new_C9271_ = ~new_C9216_ | ~new_C9241_;
  assign new_C9272_ = new_C9249_ & new_C9269_;
  assign new_C9273_ = ~new_C9249_ & ~new_C9269_;
  assign new_C9274_ = new_C9278_ | new_C9279_;
  assign new_C9275_ = ~new_C9220_ & new_C9234_;
  assign new_C9276_ = new_C9280_ | new_C9281_;
  assign new_C9277_ = new_C9220_ & new_C9234_;
  assign new_C9278_ = ~new_C9220_ & ~new_C9234_;
  assign new_C9279_ = new_C9220_ & ~new_C9234_;
  assign new_C9280_ = new_C9220_ & ~new_C9234_;
  assign new_C9281_ = ~new_C9220_ & new_C9234_;
  assign new_C9282_ = new_E8655_;
  assign new_C9283_ = new_E8722_;
  assign new_C9284_ = new_E8789_;
  assign new_C9285_ = new_E8856_;
  assign new_C9286_ = new_E8923_;
  assign new_C9287_ = new_E8990_;
  assign new_C9288_ = new_C9295_ & new_C9294_;
  assign new_C9289_ = new_C9297_ | new_C9296_;
  assign new_C9290_ = new_C9299_ | new_C9298_;
  assign new_C9291_ = new_C9301_ & new_C9300_;
  assign new_C9292_ = new_C9301_ & new_C9302_;
  assign new_C9293_ = new_C9294_ | new_C9303_;
  assign new_C9294_ = new_C9283_ | new_C9306_;
  assign new_C9295_ = new_C9305_ | new_C9304_;
  assign new_C9296_ = new_C9310_ & new_C9309_;
  assign new_C9297_ = new_C9308_ & new_C9307_;
  assign new_C9298_ = new_C9313_ | new_C9312_;
  assign new_C9299_ = new_C9308_ & new_C9311_;
  assign new_C9300_ = new_C9283_ | new_C9316_;
  assign new_C9301_ = new_C9315_ | new_C9314_;
  assign new_C9302_ = new_C9318_ | new_C9317_;
  assign new_C9303_ = ~new_C9294_ & new_C9320_;
  assign new_C9304_ = ~new_C9296_ & new_C9308_;
  assign new_C9305_ = new_C9296_ & ~new_C9308_;
  assign new_C9306_ = new_C9282_ & ~new_C9283_;
  assign new_C9307_ = ~new_C9329_ | ~new_C9330_;
  assign new_C9308_ = new_C9322_ | new_C9324_;
  assign new_C9309_ = new_C9332_ | new_C9331_;
  assign new_C9310_ = new_C9326_ | new_C9325_;
  assign new_C9311_ = ~new_C9334_ | ~new_C9333_;
  assign new_C9312_ = ~new_C9335_ & new_C9336_;
  assign new_C9313_ = new_C9335_ & ~new_C9336_;
  assign new_C9314_ = ~new_C9282_ & new_C9283_;
  assign new_C9315_ = new_C9282_ & ~new_C9283_;
  assign new_C9316_ = ~new_C9298_ | new_C9308_;
  assign new_C9317_ = new_C9298_ & new_C9308_;
  assign new_C9318_ = ~new_C9298_ & ~new_C9308_;
  assign new_C9319_ = new_C9340_ | new_C9339_;
  assign new_C9320_ = new_C9286_ | new_C9319_;
  assign new_C9321_ = new_C9344_ | new_C9343_;
  assign new_C9322_ = ~new_C9286_ & new_C9321_;
  assign new_C9323_ = new_C9342_ | new_C9341_;
  assign new_C9324_ = new_C9286_ & new_C9323_;
  assign new_C9325_ = new_C9284_ & ~new_C9294_;
  assign new_C9326_ = ~new_C9284_ & new_C9294_;
  assign new_C9327_ = ~new_C9283_ | ~new_C9308_;
  assign new_C9328_ = new_C9294_ & new_C9327_;
  assign new_C9329_ = ~new_C9294_ & ~new_C9328_;
  assign new_C9330_ = new_C9294_ | new_C9327_;
  assign new_C9331_ = ~new_C9284_ & new_C9285_;
  assign new_C9332_ = new_C9284_ & ~new_C9285_;
  assign new_C9333_ = new_C9301_ | new_C9338_;
  assign new_C9334_ = ~new_C9301_ & ~new_C9337_;
  assign new_C9335_ = new_C9284_ | new_C9301_;
  assign new_C9336_ = new_C9284_ | new_C9285_;
  assign new_C9337_ = new_C9301_ & new_C9338_;
  assign new_C9338_ = ~new_C9283_ | ~new_C9308_;
  assign new_C9339_ = new_C9316_ & new_C9336_;
  assign new_C9340_ = ~new_C9316_ & ~new_C9336_;
  assign new_C9341_ = new_C9345_ | new_C9346_;
  assign new_C9342_ = ~new_C9287_ & new_C9301_;
  assign new_C9343_ = new_C9347_ | new_C9348_;
  assign new_C9344_ = new_C9287_ & new_C9301_;
  assign new_C9345_ = ~new_C9287_ & ~new_C9301_;
  assign new_C9346_ = new_C9287_ & ~new_C9301_;
  assign new_C9347_ = new_C9287_ & ~new_C9301_;
  assign new_C9348_ = ~new_C9287_ & new_C9301_;
  assign new_C9349_ = new_E9057_;
  assign new_C9350_ = new_E9124_;
  assign new_C9351_ = new_E9191_;
  assign new_C9352_ = new_E9258_;
  assign new_C9353_ = new_E9325_;
  assign new_C9354_ = new_E9392_;
  assign new_C9355_ = new_C9362_ & new_C9361_;
  assign new_C9356_ = new_C9364_ | new_C9363_;
  assign new_C9357_ = new_C9366_ | new_C9365_;
  assign new_C9358_ = new_C9368_ & new_C9367_;
  assign new_C9359_ = new_C9368_ & new_C9369_;
  assign new_C9360_ = new_C9361_ | new_C9370_;
  assign new_C9361_ = new_C9350_ | new_C9373_;
  assign new_C9362_ = new_C9372_ | new_C9371_;
  assign new_C9363_ = new_C9377_ & new_C9376_;
  assign new_C9364_ = new_C9375_ & new_C9374_;
  assign new_C9365_ = new_C9380_ | new_C9379_;
  assign new_C9366_ = new_C9375_ & new_C9378_;
  assign new_C9367_ = new_C9350_ | new_C9383_;
  assign new_C9368_ = new_C9382_ | new_C9381_;
  assign new_C9369_ = new_C9385_ | new_C9384_;
  assign new_C9370_ = ~new_C9361_ & new_C9387_;
  assign new_C9371_ = ~new_C9363_ & new_C9375_;
  assign new_C9372_ = new_C9363_ & ~new_C9375_;
  assign new_C9373_ = new_C9349_ & ~new_C9350_;
  assign new_C9374_ = ~new_C9396_ | ~new_C9397_;
  assign new_C9375_ = new_C9389_ | new_C9391_;
  assign new_C9376_ = new_C9399_ | new_C9398_;
  assign new_C9377_ = new_C9393_ | new_C9392_;
  assign new_C9378_ = ~new_C9401_ | ~new_C9400_;
  assign new_C9379_ = ~new_C9402_ & new_C9403_;
  assign new_C9380_ = new_C9402_ & ~new_C9403_;
  assign new_C9381_ = ~new_C9349_ & new_C9350_;
  assign new_C9382_ = new_C9349_ & ~new_C9350_;
  assign new_C9383_ = ~new_C9365_ | new_C9375_;
  assign new_C9384_ = new_C9365_ & new_C9375_;
  assign new_C9385_ = ~new_C9365_ & ~new_C9375_;
  assign new_C9386_ = new_C9407_ | new_C9406_;
  assign new_C9387_ = new_C9353_ | new_C9386_;
  assign new_C9388_ = new_C9411_ | new_C9410_;
  assign new_C9389_ = ~new_C9353_ & new_C9388_;
  assign new_C9390_ = new_C9409_ | new_C9408_;
  assign new_C9391_ = new_C9353_ & new_C9390_;
  assign new_C9392_ = new_C9351_ & ~new_C9361_;
  assign new_C9393_ = ~new_C9351_ & new_C9361_;
  assign new_C9394_ = ~new_C9350_ | ~new_C9375_;
  assign new_C9395_ = new_C9361_ & new_C9394_;
  assign new_C9396_ = ~new_C9361_ & ~new_C9395_;
  assign new_C9397_ = new_C9361_ | new_C9394_;
  assign new_C9398_ = ~new_C9351_ & new_C9352_;
  assign new_C9399_ = new_C9351_ & ~new_C9352_;
  assign new_C9400_ = new_C9368_ | new_C9405_;
  assign new_C9401_ = ~new_C9368_ & ~new_C9404_;
  assign new_C9402_ = new_C9351_ | new_C9368_;
  assign new_C9403_ = new_C9351_ | new_C9352_;
  assign new_C9404_ = new_C9368_ & new_C9405_;
  assign new_C9405_ = ~new_C9350_ | ~new_C9375_;
  assign new_C9406_ = new_C9383_ & new_C9403_;
  assign new_C9407_ = ~new_C9383_ & ~new_C9403_;
  assign new_C9408_ = new_C9412_ | new_C9413_;
  assign new_C9409_ = ~new_C9354_ & new_C9368_;
  assign new_C9410_ = new_C9414_ | new_C9415_;
  assign new_C9411_ = new_C9354_ & new_C9368_;
  assign new_C9412_ = ~new_C9354_ & ~new_C9368_;
  assign new_C9413_ = new_C9354_ & ~new_C9368_;
  assign new_C9414_ = new_C9354_ & ~new_C9368_;
  assign new_C9415_ = ~new_C9354_ & new_C9368_;
  assign new_C9416_ = new_E9459_;
  assign new_C9417_ = new_E9526_;
  assign new_C9418_ = new_E9593_;
  assign new_C9419_ = new_E9660_;
  assign new_C9420_ = new_E9727_;
  assign new_C9421_ = new_E9794_;
  assign new_C9422_ = new_C9429_ & new_C9428_;
  assign new_C9423_ = new_C9431_ | new_C9430_;
  assign new_C9424_ = new_C9433_ | new_C9432_;
  assign new_C9425_ = new_C9435_ & new_C9434_;
  assign new_C9426_ = new_C9435_ & new_C9436_;
  assign new_C9427_ = new_C9428_ | new_C9437_;
  assign new_C9428_ = new_C9417_ | new_C9440_;
  assign new_C9429_ = new_C9439_ | new_C9438_;
  assign new_C9430_ = new_C9444_ & new_C9443_;
  assign new_C9431_ = new_C9442_ & new_C9441_;
  assign new_C9432_ = new_C9447_ | new_C9446_;
  assign new_C9433_ = new_C9442_ & new_C9445_;
  assign new_C9434_ = new_C9417_ | new_C9450_;
  assign new_C9435_ = new_C9449_ | new_C9448_;
  assign new_C9436_ = new_C9452_ | new_C9451_;
  assign new_C9437_ = ~new_C9428_ & new_C9454_;
  assign new_C9438_ = ~new_C9430_ & new_C9442_;
  assign new_C9439_ = new_C9430_ & ~new_C9442_;
  assign new_C9440_ = new_C9416_ & ~new_C9417_;
  assign new_C9441_ = ~new_C9463_ | ~new_C9464_;
  assign new_C9442_ = new_C9456_ | new_C9458_;
  assign new_C9443_ = new_C9466_ | new_C9465_;
  assign new_C9444_ = new_C9460_ | new_C9459_;
  assign new_C9445_ = ~new_C9468_ | ~new_C9467_;
  assign new_C9446_ = ~new_C9469_ & new_C9470_;
  assign new_C9447_ = new_C9469_ & ~new_C9470_;
  assign new_C9448_ = ~new_C9416_ & new_C9417_;
  assign new_C9449_ = new_C9416_ & ~new_C9417_;
  assign new_C9450_ = ~new_C9432_ | new_C9442_;
  assign new_C9451_ = new_C9432_ & new_C9442_;
  assign new_C9452_ = ~new_C9432_ & ~new_C9442_;
  assign new_C9453_ = new_C9474_ | new_C9473_;
  assign new_C9454_ = new_C9420_ | new_C9453_;
  assign new_C9455_ = new_C9478_ | new_C9477_;
  assign new_C9456_ = ~new_C9420_ & new_C9455_;
  assign new_C9457_ = new_C9476_ | new_C9475_;
  assign new_C9458_ = new_C9420_ & new_C9457_;
  assign new_C9459_ = new_C9418_ & ~new_C9428_;
  assign new_C9460_ = ~new_C9418_ & new_C9428_;
  assign new_C9461_ = ~new_C9417_ | ~new_C9442_;
  assign new_C9462_ = new_C9428_ & new_C9461_;
  assign new_C9463_ = ~new_C9428_ & ~new_C9462_;
  assign new_C9464_ = new_C9428_ | new_C9461_;
  assign new_C9465_ = ~new_C9418_ & new_C9419_;
  assign new_C9466_ = new_C9418_ & ~new_C9419_;
  assign new_C9467_ = new_C9435_ | new_C9472_;
  assign new_C9468_ = ~new_C9435_ & ~new_C9471_;
  assign new_C9469_ = new_C9418_ | new_C9435_;
  assign new_C9470_ = new_C9418_ | new_C9419_;
  assign new_C9471_ = new_C9435_ & new_C9472_;
  assign new_C9472_ = ~new_C9417_ | ~new_C9442_;
  assign new_C9473_ = new_C9450_ & new_C9470_;
  assign new_C9474_ = ~new_C9450_ & ~new_C9470_;
  assign new_C9475_ = new_C9479_ | new_C9480_;
  assign new_C9476_ = ~new_C9421_ & new_C9435_;
  assign new_C9477_ = new_C9481_ | new_C9482_;
  assign new_C9478_ = new_C9421_ & new_C9435_;
  assign new_C9479_ = ~new_C9421_ & ~new_C9435_;
  assign new_C9480_ = new_C9421_ & ~new_C9435_;
  assign new_C9481_ = new_C9421_ & ~new_C9435_;
  assign new_C9482_ = ~new_C9421_ & new_C9435_;
  assign new_C9483_ = new_E9861_;
  assign new_C9484_ = new_E9928_;
  assign new_C9485_ = new_E9995_;
  assign new_C9486_ = new_F63_;
  assign new_C9487_ = new_F130_;
  assign new_C9488_ = new_F197_;
  assign new_C9489_ = new_C9496_ & new_C9495_;
  assign new_C9490_ = new_C9498_ | new_C9497_;
  assign new_C9491_ = new_C9500_ | new_C9499_;
  assign new_C9492_ = new_C9502_ & new_C9501_;
  assign new_C9493_ = new_C9502_ & new_C9503_;
  assign new_C9494_ = new_C9495_ | new_C9504_;
  assign new_C9495_ = new_C9484_ | new_C9507_;
  assign new_C9496_ = new_C9506_ | new_C9505_;
  assign new_C9497_ = new_C9511_ & new_C9510_;
  assign new_C9498_ = new_C9509_ & new_C9508_;
  assign new_C9499_ = new_C9514_ | new_C9513_;
  assign new_C9500_ = new_C9509_ & new_C9512_;
  assign new_C9501_ = new_C9484_ | new_C9517_;
  assign new_C9502_ = new_C9516_ | new_C9515_;
  assign new_C9503_ = new_C9519_ | new_C9518_;
  assign new_C9504_ = ~new_C9495_ & new_C9521_;
  assign new_C9505_ = ~new_C9497_ & new_C9509_;
  assign new_C9506_ = new_C9497_ & ~new_C9509_;
  assign new_C9507_ = new_C9483_ & ~new_C9484_;
  assign new_C9508_ = ~new_C9530_ | ~new_C9531_;
  assign new_C9509_ = new_C9523_ | new_C9525_;
  assign new_C9510_ = new_C9533_ | new_C9532_;
  assign new_C9511_ = new_C9527_ | new_C9526_;
  assign new_C9512_ = ~new_C9535_ | ~new_C9534_;
  assign new_C9513_ = ~new_C9536_ & new_C9537_;
  assign new_C9514_ = new_C9536_ & ~new_C9537_;
  assign new_C9515_ = ~new_C9483_ & new_C9484_;
  assign new_C9516_ = new_C9483_ & ~new_C9484_;
  assign new_C9517_ = ~new_C9499_ | new_C9509_;
  assign new_C9518_ = new_C9499_ & new_C9509_;
  assign new_C9519_ = ~new_C9499_ & ~new_C9509_;
  assign new_C9520_ = new_C9541_ | new_C9540_;
  assign new_C9521_ = new_C9487_ | new_C9520_;
  assign new_C9522_ = new_C9545_ | new_C9544_;
  assign new_C9523_ = ~new_C9487_ & new_C9522_;
  assign new_C9524_ = new_C9543_ | new_C9542_;
  assign new_C9525_ = new_C9487_ & new_C9524_;
  assign new_C9526_ = new_C9485_ & ~new_C9495_;
  assign new_C9527_ = ~new_C9485_ & new_C9495_;
  assign new_C9528_ = ~new_C9484_ | ~new_C9509_;
  assign new_C9529_ = new_C9495_ & new_C9528_;
  assign new_C9530_ = ~new_C9495_ & ~new_C9529_;
  assign new_C9531_ = new_C9495_ | new_C9528_;
  assign new_C9532_ = ~new_C9485_ & new_C9486_;
  assign new_C9533_ = new_C9485_ & ~new_C9486_;
  assign new_C9534_ = new_C9502_ | new_C9539_;
  assign new_C9535_ = ~new_C9502_ & ~new_C9538_;
  assign new_C9536_ = new_C9485_ | new_C9502_;
  assign new_C9537_ = new_C9485_ | new_C9486_;
  assign new_C9538_ = new_C9502_ & new_C9539_;
  assign new_C9539_ = ~new_C9484_ | ~new_C9509_;
  assign new_C9540_ = new_C9517_ & new_C9537_;
  assign new_C9541_ = ~new_C9517_ & ~new_C9537_;
  assign new_C9542_ = new_C9546_ | new_C9547_;
  assign new_C9543_ = ~new_C9488_ & new_C9502_;
  assign new_C9544_ = new_C9548_ | new_C9549_;
  assign new_C9545_ = new_C9488_ & new_C9502_;
  assign new_C9546_ = ~new_C9488_ & ~new_C9502_;
  assign new_C9547_ = new_C9488_ & ~new_C9502_;
  assign new_C9548_ = new_C9488_ & ~new_C9502_;
  assign new_C9549_ = ~new_C9488_ & new_C9502_;
  assign new_C9550_ = new_F264_;
  assign new_C9551_ = new_F331_;
  assign new_C9552_ = new_F398_;
  assign new_C9553_ = new_F465_;
  assign new_C9554_ = new_F532_;
  assign new_C9555_ = new_F599_;
  assign new_C9556_ = new_C9563_ & new_C9562_;
  assign new_C9557_ = new_C9565_ | new_C9564_;
  assign new_C9558_ = new_C9567_ | new_C9566_;
  assign new_C9559_ = new_C9569_ & new_C9568_;
  assign new_C9560_ = new_C9569_ & new_C9570_;
  assign new_C9561_ = new_C9562_ | new_C9571_;
  assign new_C9562_ = new_C9551_ | new_C9574_;
  assign new_C9563_ = new_C9573_ | new_C9572_;
  assign new_C9564_ = new_C9578_ & new_C9577_;
  assign new_C9565_ = new_C9576_ & new_C9575_;
  assign new_C9566_ = new_C9581_ | new_C9580_;
  assign new_C9567_ = new_C9576_ & new_C9579_;
  assign new_C9568_ = new_C9551_ | new_C9584_;
  assign new_C9569_ = new_C9583_ | new_C9582_;
  assign new_C9570_ = new_C9586_ | new_C9585_;
  assign new_C9571_ = ~new_C9562_ & new_C9588_;
  assign new_C9572_ = ~new_C9564_ & new_C9576_;
  assign new_C9573_ = new_C9564_ & ~new_C9576_;
  assign new_C9574_ = new_C9550_ & ~new_C9551_;
  assign new_C9575_ = ~new_C9597_ | ~new_C9598_;
  assign new_C9576_ = new_C9590_ | new_C9592_;
  assign new_C9577_ = new_C9600_ | new_C9599_;
  assign new_C9578_ = new_C9594_ | new_C9593_;
  assign new_C9579_ = ~new_C9602_ | ~new_C9601_;
  assign new_C9580_ = ~new_C9603_ & new_C9604_;
  assign new_C9581_ = new_C9603_ & ~new_C9604_;
  assign new_C9582_ = ~new_C9550_ & new_C9551_;
  assign new_C9583_ = new_C9550_ & ~new_C9551_;
  assign new_C9584_ = ~new_C9566_ | new_C9576_;
  assign new_C9585_ = new_C9566_ & new_C9576_;
  assign new_C9586_ = ~new_C9566_ & ~new_C9576_;
  assign new_C9587_ = new_C9608_ | new_C9607_;
  assign new_C9588_ = new_C9554_ | new_C9587_;
  assign new_C9589_ = new_C9612_ | new_C9611_;
  assign new_C9590_ = ~new_C9554_ & new_C9589_;
  assign new_C9591_ = new_C9610_ | new_C9609_;
  assign new_C9592_ = new_C9554_ & new_C9591_;
  assign new_C9593_ = new_C9552_ & ~new_C9562_;
  assign new_C9594_ = ~new_C9552_ & new_C9562_;
  assign new_C9595_ = ~new_C9551_ | ~new_C9576_;
  assign new_C9596_ = new_C9562_ & new_C9595_;
  assign new_C9597_ = ~new_C9562_ & ~new_C9596_;
  assign new_C9598_ = new_C9562_ | new_C9595_;
  assign new_C9599_ = ~new_C9552_ & new_C9553_;
  assign new_C9600_ = new_C9552_ & ~new_C9553_;
  assign new_C9601_ = new_C9569_ | new_C9606_;
  assign new_C9602_ = ~new_C9569_ & ~new_C9605_;
  assign new_C9603_ = new_C9552_ | new_C9569_;
  assign new_C9604_ = new_C9552_ | new_C9553_;
  assign new_C9605_ = new_C9569_ & new_C9606_;
  assign new_C9606_ = ~new_C9551_ | ~new_C9576_;
  assign new_C9607_ = new_C9584_ & new_C9604_;
  assign new_C9608_ = ~new_C9584_ & ~new_C9604_;
  assign new_C9609_ = new_C9613_ | new_C9614_;
  assign new_C9610_ = ~new_C9555_ & new_C9569_;
  assign new_C9611_ = new_C9615_ | new_C9616_;
  assign new_C9612_ = new_C9555_ & new_C9569_;
  assign new_C9613_ = ~new_C9555_ & ~new_C9569_;
  assign new_C9614_ = new_C9555_ & ~new_C9569_;
  assign new_C9615_ = new_C9555_ & ~new_C9569_;
  assign new_C9616_ = ~new_C9555_ & new_C9569_;
  assign new_C9617_ = new_F666_;
  assign new_C9618_ = new_F733_;
  assign new_C9619_ = new_F800_;
  assign new_C9620_ = new_F867_;
  assign new_C9621_ = new_F934_;
  assign new_C9622_ = new_F1001_;
  assign new_C9623_ = new_C9630_ & new_C9629_;
  assign new_C9624_ = new_C9632_ | new_C9631_;
  assign new_C9625_ = new_C9634_ | new_C9633_;
  assign new_C9626_ = new_C9636_ & new_C9635_;
  assign new_C9627_ = new_C9636_ & new_C9637_;
  assign new_C9628_ = new_C9629_ | new_C9638_;
  assign new_C9629_ = new_C9618_ | new_C9641_;
  assign new_C9630_ = new_C9640_ | new_C9639_;
  assign new_C9631_ = new_C9645_ & new_C9644_;
  assign new_C9632_ = new_C9643_ & new_C9642_;
  assign new_C9633_ = new_C9648_ | new_C9647_;
  assign new_C9634_ = new_C9643_ & new_C9646_;
  assign new_C9635_ = new_C9618_ | new_C9651_;
  assign new_C9636_ = new_C9650_ | new_C9649_;
  assign new_C9637_ = new_C9653_ | new_C9652_;
  assign new_C9638_ = ~new_C9629_ & new_C9655_;
  assign new_C9639_ = ~new_C9631_ & new_C9643_;
  assign new_C9640_ = new_C9631_ & ~new_C9643_;
  assign new_C9641_ = new_C9617_ & ~new_C9618_;
  assign new_C9642_ = ~new_C9664_ | ~new_C9665_;
  assign new_C9643_ = new_C9657_ | new_C9659_;
  assign new_C9644_ = new_C9667_ | new_C9666_;
  assign new_C9645_ = new_C9661_ | new_C9660_;
  assign new_C9646_ = ~new_C9669_ | ~new_C9668_;
  assign new_C9647_ = ~new_C9670_ & new_C9671_;
  assign new_C9648_ = new_C9670_ & ~new_C9671_;
  assign new_C9649_ = ~new_C9617_ & new_C9618_;
  assign new_C9650_ = new_C9617_ & ~new_C9618_;
  assign new_C9651_ = ~new_C9633_ | new_C9643_;
  assign new_C9652_ = new_C9633_ & new_C9643_;
  assign new_C9653_ = ~new_C9633_ & ~new_C9643_;
  assign new_C9654_ = new_C9675_ | new_C9674_;
  assign new_C9655_ = new_C9621_ | new_C9654_;
  assign new_C9656_ = new_C9679_ | new_C9678_;
  assign new_C9657_ = ~new_C9621_ & new_C9656_;
  assign new_C9658_ = new_C9677_ | new_C9676_;
  assign new_C9659_ = new_C9621_ & new_C9658_;
  assign new_C9660_ = new_C9619_ & ~new_C9629_;
  assign new_C9661_ = ~new_C9619_ & new_C9629_;
  assign new_C9662_ = ~new_C9618_ | ~new_C9643_;
  assign new_C9663_ = new_C9629_ & new_C9662_;
  assign new_C9664_ = ~new_C9629_ & ~new_C9663_;
  assign new_C9665_ = new_C9629_ | new_C9662_;
  assign new_C9666_ = ~new_C9619_ & new_C9620_;
  assign new_C9667_ = new_C9619_ & ~new_C9620_;
  assign new_C9668_ = new_C9636_ | new_C9673_;
  assign new_C9669_ = ~new_C9636_ & ~new_C9672_;
  assign new_C9670_ = new_C9619_ | new_C9636_;
  assign new_C9671_ = new_C9619_ | new_C9620_;
  assign new_C9672_ = new_C9636_ & new_C9673_;
  assign new_C9673_ = ~new_C9618_ | ~new_C9643_;
  assign new_C9674_ = new_C9651_ & new_C9671_;
  assign new_C9675_ = ~new_C9651_ & ~new_C9671_;
  assign new_C9676_ = new_C9680_ | new_C9681_;
  assign new_C9677_ = ~new_C9622_ & new_C9636_;
  assign new_C9678_ = new_C9682_ | new_C9683_;
  assign new_C9679_ = new_C9622_ & new_C9636_;
  assign new_C9680_ = ~new_C9622_ & ~new_C9636_;
  assign new_C9681_ = new_C9622_ & ~new_C9636_;
  assign new_C9682_ = new_C9622_ & ~new_C9636_;
  assign new_C9683_ = ~new_C9622_ & new_C9636_;
  assign new_C9684_ = new_F1068_;
  assign new_C9685_ = new_F1135_;
  assign new_C9686_ = new_F1202_;
  assign new_C9687_ = new_F1269_;
  assign new_C9688_ = new_F1336_;
  assign new_C9689_ = new_F1403_;
  assign new_C9690_ = new_C9697_ & new_C9696_;
  assign new_C9691_ = new_C9699_ | new_C9698_;
  assign new_C9692_ = new_C9701_ | new_C9700_;
  assign new_C9693_ = new_C9703_ & new_C9702_;
  assign new_C9694_ = new_C9703_ & new_C9704_;
  assign new_C9695_ = new_C9696_ | new_C9705_;
  assign new_C9696_ = new_C9685_ | new_C9708_;
  assign new_C9697_ = new_C9707_ | new_C9706_;
  assign new_C9698_ = new_C9712_ & new_C9711_;
  assign new_C9699_ = new_C9710_ & new_C9709_;
  assign new_C9700_ = new_C9715_ | new_C9714_;
  assign new_C9701_ = new_C9710_ & new_C9713_;
  assign new_C9702_ = new_C9685_ | new_C9718_;
  assign new_C9703_ = new_C9717_ | new_C9716_;
  assign new_C9704_ = new_C9720_ | new_C9719_;
  assign new_C9705_ = ~new_C9696_ & new_C9722_;
  assign new_C9706_ = ~new_C9698_ & new_C9710_;
  assign new_C9707_ = new_C9698_ & ~new_C9710_;
  assign new_C9708_ = new_C9684_ & ~new_C9685_;
  assign new_C9709_ = ~new_C9731_ | ~new_C9732_;
  assign new_C9710_ = new_C9724_ | new_C9726_;
  assign new_C9711_ = new_C9734_ | new_C9733_;
  assign new_C9712_ = new_C9728_ | new_C9727_;
  assign new_C9713_ = ~new_C9736_ | ~new_C9735_;
  assign new_C9714_ = ~new_C9737_ & new_C9738_;
  assign new_C9715_ = new_C9737_ & ~new_C9738_;
  assign new_C9716_ = ~new_C9684_ & new_C9685_;
  assign new_C9717_ = new_C9684_ & ~new_C9685_;
  assign new_C9718_ = ~new_C9700_ | new_C9710_;
  assign new_C9719_ = new_C9700_ & new_C9710_;
  assign new_C9720_ = ~new_C9700_ & ~new_C9710_;
  assign new_C9721_ = new_C9742_ | new_C9741_;
  assign new_C9722_ = new_C9688_ | new_C9721_;
  assign new_C9723_ = new_C9746_ | new_C9745_;
  assign new_C9724_ = ~new_C9688_ & new_C9723_;
  assign new_C9725_ = new_C9744_ | new_C9743_;
  assign new_C9726_ = new_C9688_ & new_C9725_;
  assign new_C9727_ = new_C9686_ & ~new_C9696_;
  assign new_C9728_ = ~new_C9686_ & new_C9696_;
  assign new_C9729_ = ~new_C9685_ | ~new_C9710_;
  assign new_C9730_ = new_C9696_ & new_C9729_;
  assign new_C9731_ = ~new_C9696_ & ~new_C9730_;
  assign new_C9732_ = new_C9696_ | new_C9729_;
  assign new_C9733_ = ~new_C9686_ & new_C9687_;
  assign new_C9734_ = new_C9686_ & ~new_C9687_;
  assign new_C9735_ = new_C9703_ | new_C9740_;
  assign new_C9736_ = ~new_C9703_ & ~new_C9739_;
  assign new_C9737_ = new_C9686_ | new_C9703_;
  assign new_C9738_ = new_C9686_ | new_C9687_;
  assign new_C9739_ = new_C9703_ & new_C9740_;
  assign new_C9740_ = ~new_C9685_ | ~new_C9710_;
  assign new_C9741_ = new_C9718_ & new_C9738_;
  assign new_C9742_ = ~new_C9718_ & ~new_C9738_;
  assign new_C9743_ = new_C9747_ | new_C9748_;
  assign new_C9744_ = ~new_C9689_ & new_C9703_;
  assign new_C9745_ = new_C9749_ | new_C9750_;
  assign new_C9746_ = new_C9689_ & new_C9703_;
  assign new_C9747_ = ~new_C9689_ & ~new_C9703_;
  assign new_C9748_ = new_C9689_ & ~new_C9703_;
  assign new_C9749_ = new_C9689_ & ~new_C9703_;
  assign new_C9750_ = ~new_C9689_ & new_C9703_;
  assign new_C9751_ = new_D6996_;
  assign new_C9752_ = new_D7064_;
  assign new_C9753_ = new_D7131_;
  assign new_C9754_ = new_D7198_;
  assign new_C9755_ = new_D7265_;
  assign new_C9756_ = new_D7332_;
  assign new_C9757_ = new_C9764_ & new_C9763_;
  assign new_C9758_ = new_C9766_ | new_C9765_;
  assign new_C9759_ = new_C9768_ | new_C9767_;
  assign new_C9760_ = new_C9770_ & new_C9769_;
  assign new_C9761_ = new_C9770_ & new_C9771_;
  assign new_C9762_ = new_C9763_ | new_C9772_;
  assign new_C9763_ = new_C9752_ | new_C9775_;
  assign new_C9764_ = new_C9774_ | new_C9773_;
  assign new_C9765_ = new_C9779_ & new_C9778_;
  assign new_C9766_ = new_C9777_ & new_C9776_;
  assign new_C9767_ = new_C9782_ | new_C9781_;
  assign new_C9768_ = new_C9777_ & new_C9780_;
  assign new_C9769_ = new_C9752_ | new_C9785_;
  assign new_C9770_ = new_C9784_ | new_C9783_;
  assign new_C9771_ = new_C9787_ | new_C9786_;
  assign new_C9772_ = ~new_C9763_ & new_C9789_;
  assign new_C9773_ = ~new_C9765_ & new_C9777_;
  assign new_C9774_ = new_C9765_ & ~new_C9777_;
  assign new_C9775_ = new_C9751_ & ~new_C9752_;
  assign new_C9776_ = ~new_C9798_ | ~new_C9799_;
  assign new_C9777_ = new_C9791_ | new_C9793_;
  assign new_C9778_ = new_C9801_ | new_C9800_;
  assign new_C9779_ = new_C9795_ | new_C9794_;
  assign new_C9780_ = ~new_C9803_ | ~new_C9802_;
  assign new_C9781_ = ~new_C9804_ & new_C9805_;
  assign new_C9782_ = new_C9804_ & ~new_C9805_;
  assign new_C9783_ = ~new_C9751_ & new_C9752_;
  assign new_C9784_ = new_C9751_ & ~new_C9752_;
  assign new_C9785_ = ~new_C9767_ | new_C9777_;
  assign new_C9786_ = new_C9767_ & new_C9777_;
  assign new_C9787_ = ~new_C9767_ & ~new_C9777_;
  assign new_C9788_ = new_C9809_ | new_C9808_;
  assign new_C9789_ = new_C9755_ | new_C9788_;
  assign new_C9790_ = new_C9813_ | new_C9812_;
  assign new_C9791_ = ~new_C9755_ & new_C9790_;
  assign new_C9792_ = new_C9811_ | new_C9810_;
  assign new_C9793_ = new_C9755_ & new_C9792_;
  assign new_C9794_ = new_C9753_ & ~new_C9763_;
  assign new_C9795_ = ~new_C9753_ & new_C9763_;
  assign new_C9796_ = ~new_C9752_ | ~new_C9777_;
  assign new_C9797_ = new_C9763_ & new_C9796_;
  assign new_C9798_ = ~new_C9763_ & ~new_C9797_;
  assign new_C9799_ = new_C9763_ | new_C9796_;
  assign new_C9800_ = ~new_C9753_ & new_C9754_;
  assign new_C9801_ = new_C9753_ & ~new_C9754_;
  assign new_C9802_ = new_C9770_ | new_C9807_;
  assign new_C9803_ = ~new_C9770_ & ~new_C9806_;
  assign new_C9804_ = new_C9753_ | new_C9770_;
  assign new_C9805_ = new_C9753_ | new_C9754_;
  assign new_C9806_ = new_C9770_ & new_C9807_;
  assign new_C9807_ = ~new_C9752_ | ~new_C9777_;
  assign new_C9808_ = new_C9785_ & new_C9805_;
  assign new_C9809_ = ~new_C9785_ & ~new_C9805_;
  assign new_C9810_ = new_C9814_ | new_C9815_;
  assign new_C9811_ = ~new_C9756_ & new_C9770_;
  assign new_C9812_ = new_C9816_ | new_C9817_;
  assign new_C9813_ = new_C9756_ & new_C9770_;
  assign new_C9814_ = ~new_C9756_ & ~new_C9770_;
  assign new_C9815_ = new_C9756_ & ~new_C9770_;
  assign new_C9816_ = new_C9756_ & ~new_C9770_;
  assign new_C9817_ = ~new_C9756_ & new_C9770_;
  assign new_C9818_ = new_D7399_;
  assign new_C9819_ = new_D7466_;
  assign new_C9820_ = new_D7533_;
  assign new_C9821_ = new_D7600_;
  assign new_C9822_ = new_D7667_;
  assign new_C9823_ = new_D7734_;
  assign new_C9824_ = new_C9831_ & new_C9830_;
  assign new_C9825_ = new_C9833_ | new_C9832_;
  assign new_C9826_ = new_C9835_ | new_C9834_;
  assign new_C9827_ = new_C9837_ & new_C9836_;
  assign new_C9828_ = new_C9837_ & new_C9838_;
  assign new_C9829_ = new_C9830_ | new_C9839_;
  assign new_C9830_ = new_C9819_ | new_C9842_;
  assign new_C9831_ = new_C9841_ | new_C9840_;
  assign new_C9832_ = new_C9846_ & new_C9845_;
  assign new_C9833_ = new_C9844_ & new_C9843_;
  assign new_C9834_ = new_C9849_ | new_C9848_;
  assign new_C9835_ = new_C9844_ & new_C9847_;
  assign new_C9836_ = new_C9819_ | new_C9852_;
  assign new_C9837_ = new_C9851_ | new_C9850_;
  assign new_C9838_ = new_C9854_ | new_C9853_;
  assign new_C9839_ = ~new_C9830_ & new_C9856_;
  assign new_C9840_ = ~new_C9832_ & new_C9844_;
  assign new_C9841_ = new_C9832_ & ~new_C9844_;
  assign new_C9842_ = new_C9818_ & ~new_C9819_;
  assign new_C9843_ = ~new_C9865_ | ~new_C9866_;
  assign new_C9844_ = new_C9858_ | new_C9860_;
  assign new_C9845_ = new_C9868_ | new_C9867_;
  assign new_C9846_ = new_C9862_ | new_C9861_;
  assign new_C9847_ = ~new_C9870_ | ~new_C9869_;
  assign new_C9848_ = ~new_C9871_ & new_C9872_;
  assign new_C9849_ = new_C9871_ & ~new_C9872_;
  assign new_C9850_ = ~new_C9818_ & new_C9819_;
  assign new_C9851_ = new_C9818_ & ~new_C9819_;
  assign new_C9852_ = ~new_C9834_ | new_C9844_;
  assign new_C9853_ = new_C9834_ & new_C9844_;
  assign new_C9854_ = ~new_C9834_ & ~new_C9844_;
  assign new_C9855_ = new_C9876_ | new_C9875_;
  assign new_C9856_ = new_C9822_ | new_C9855_;
  assign new_C9857_ = new_C9880_ | new_C9879_;
  assign new_C9858_ = ~new_C9822_ & new_C9857_;
  assign new_C9859_ = new_C9878_ | new_C9877_;
  assign new_C9860_ = new_C9822_ & new_C9859_;
  assign new_C9861_ = new_C9820_ & ~new_C9830_;
  assign new_C9862_ = ~new_C9820_ & new_C9830_;
  assign new_C9863_ = ~new_C9819_ | ~new_C9844_;
  assign new_C9864_ = new_C9830_ & new_C9863_;
  assign new_C9865_ = ~new_C9830_ & ~new_C9864_;
  assign new_C9866_ = new_C9830_ | new_C9863_;
  assign new_C9867_ = ~new_C9820_ & new_C9821_;
  assign new_C9868_ = new_C9820_ & ~new_C9821_;
  assign new_C9869_ = new_C9837_ | new_C9874_;
  assign new_C9870_ = ~new_C9837_ & ~new_C9873_;
  assign new_C9871_ = new_C9820_ | new_C9837_;
  assign new_C9872_ = new_C9820_ | new_C9821_;
  assign new_C9873_ = new_C9837_ & new_C9874_;
  assign new_C9874_ = ~new_C9819_ | ~new_C9844_;
  assign new_C9875_ = new_C9852_ & new_C9872_;
  assign new_C9876_ = ~new_C9852_ & ~new_C9872_;
  assign new_C9877_ = new_C9881_ | new_C9882_;
  assign new_C9878_ = ~new_C9823_ & new_C9837_;
  assign new_C9879_ = new_C9883_ | new_C9884_;
  assign new_C9880_ = new_C9823_ & new_C9837_;
  assign new_C9881_ = ~new_C9823_ & ~new_C9837_;
  assign new_C9882_ = new_C9823_ & ~new_C9837_;
  assign new_C9883_ = new_C9823_ & ~new_C9837_;
  assign new_C9884_ = ~new_C9823_ & new_C9837_;
  assign new_C9885_ = new_D7801_;
  assign new_C9886_ = new_D7868_;
  assign new_C9887_ = new_D7935_;
  assign new_C9888_ = new_D8002_;
  assign new_C9889_ = new_D8069_;
  assign new_C9890_ = new_D8136_;
  assign new_C9891_ = new_C9898_ & new_C9897_;
  assign new_C9892_ = new_C9900_ | new_C9899_;
  assign new_C9893_ = new_C9902_ | new_C9901_;
  assign new_C9894_ = new_C9904_ & new_C9903_;
  assign new_C9895_ = new_C9904_ & new_C9905_;
  assign new_C9896_ = new_C9897_ | new_C9906_;
  assign new_C9897_ = new_C9886_ | new_C9909_;
  assign new_C9898_ = new_C9908_ | new_C9907_;
  assign new_C9899_ = new_C9913_ & new_C9912_;
  assign new_C9900_ = new_C9911_ & new_C9910_;
  assign new_C9901_ = new_C9916_ | new_C9915_;
  assign new_C9902_ = new_C9911_ & new_C9914_;
  assign new_C9903_ = new_C9886_ | new_C9919_;
  assign new_C9904_ = new_C9918_ | new_C9917_;
  assign new_C9905_ = new_C9921_ | new_C9920_;
  assign new_C9906_ = ~new_C9897_ & new_C9923_;
  assign new_C9907_ = ~new_C9899_ & new_C9911_;
  assign new_C9908_ = new_C9899_ & ~new_C9911_;
  assign new_C9909_ = new_C9885_ & ~new_C9886_;
  assign new_C9910_ = ~new_C9932_ | ~new_C9933_;
  assign new_C9911_ = new_C9925_ | new_C9927_;
  assign new_C9912_ = new_C9935_ | new_C9934_;
  assign new_C9913_ = new_C9929_ | new_C9928_;
  assign new_C9914_ = ~new_C9937_ | ~new_C9936_;
  assign new_C9915_ = ~new_C9938_ & new_C9939_;
  assign new_C9916_ = new_C9938_ & ~new_C9939_;
  assign new_C9917_ = ~new_C9885_ & new_C9886_;
  assign new_C9918_ = new_C9885_ & ~new_C9886_;
  assign new_C9919_ = ~new_C9901_ | new_C9911_;
  assign new_C9920_ = new_C9901_ & new_C9911_;
  assign new_C9921_ = ~new_C9901_ & ~new_C9911_;
  assign new_C9922_ = new_C9943_ | new_C9942_;
  assign new_C9923_ = new_C9889_ | new_C9922_;
  assign new_C9924_ = new_C9947_ | new_C9946_;
  assign new_C9925_ = ~new_C9889_ & new_C9924_;
  assign new_C9926_ = new_C9945_ | new_C9944_;
  assign new_C9927_ = new_C9889_ & new_C9926_;
  assign new_C9928_ = new_C9887_ & ~new_C9897_;
  assign new_C9929_ = ~new_C9887_ & new_C9897_;
  assign new_C9930_ = ~new_C9886_ | ~new_C9911_;
  assign new_C9931_ = new_C9897_ & new_C9930_;
  assign new_C9932_ = ~new_C9897_ & ~new_C9931_;
  assign new_C9933_ = new_C9897_ | new_C9930_;
  assign new_C9934_ = ~new_C9887_ & new_C9888_;
  assign new_C9935_ = new_C9887_ & ~new_C9888_;
  assign new_C9936_ = new_C9904_ | new_C9941_;
  assign new_C9937_ = ~new_C9904_ & ~new_C9940_;
  assign new_C9938_ = new_C9887_ | new_C9904_;
  assign new_C9939_ = new_C9887_ | new_C9888_;
  assign new_C9940_ = new_C9904_ & new_C9941_;
  assign new_C9941_ = ~new_C9886_ | ~new_C9911_;
  assign new_C9942_ = new_C9919_ & new_C9939_;
  assign new_C9943_ = ~new_C9919_ & ~new_C9939_;
  assign new_C9944_ = new_C9948_ | new_C9949_;
  assign new_C9945_ = ~new_C9890_ & new_C9904_;
  assign new_C9946_ = new_C9950_ | new_C9951_;
  assign new_C9947_ = new_C9890_ & new_C9904_;
  assign new_C9948_ = ~new_C9890_ & ~new_C9904_;
  assign new_C9949_ = new_C9890_ & ~new_C9904_;
  assign new_C9950_ = new_C9890_ & ~new_C9904_;
  assign new_C9951_ = ~new_C9890_ & new_C9904_;
  assign new_C9952_ = new_D8203_;
  assign new_C9953_ = new_D8270_;
  assign new_C9954_ = new_D8337_;
  assign new_C9955_ = new_D8404_;
  assign new_C9956_ = new_D8471_;
  assign new_C9957_ = new_D8538_;
  assign new_C9958_ = new_C9965_ & new_C9964_;
  assign new_C9959_ = new_C9967_ | new_C9966_;
  assign new_C9960_ = new_C9969_ | new_C9968_;
  assign new_C9961_ = new_C9971_ & new_C9970_;
  assign new_C9962_ = new_C9971_ & new_C9972_;
  assign new_C9963_ = new_C9964_ | new_C9973_;
  assign new_C9964_ = new_C9953_ | new_C9976_;
  assign new_C9965_ = new_C9975_ | new_C9974_;
  assign new_C9966_ = new_C9980_ & new_C9979_;
  assign new_C9967_ = new_C9978_ & new_C9977_;
  assign new_C9968_ = new_C9983_ | new_C9982_;
  assign new_C9969_ = new_C9978_ & new_C9981_;
  assign new_C9970_ = new_C9953_ | new_C9986_;
  assign new_C9971_ = new_C9985_ | new_C9984_;
  assign new_C9972_ = new_C9988_ | new_C9987_;
  assign new_C9973_ = ~new_C9964_ & new_C9990_;
  assign new_C9974_ = ~new_C9966_ & new_C9978_;
  assign new_C9975_ = new_C9966_ & ~new_C9978_;
  assign new_C9976_ = new_C9952_ & ~new_C9953_;
  assign new_C9977_ = ~new_C9999_ | ~new_D1_;
  assign new_C9978_ = new_C9992_ | new_C9994_;
  assign new_C9979_ = new_D3_ | new_D2_;
  assign new_C9980_ = new_C9996_ | new_C9995_;
  assign new_C9981_ = ~new_D5_ | ~new_D4_;
  assign new_C9982_ = ~new_D6_ & new_D7_;
  assign new_C9983_ = new_D6_ & ~new_D7_;
  assign new_C9984_ = ~new_C9952_ & new_C9953_;
  assign new_C9985_ = new_C9952_ & ~new_C9953_;
  assign new_C9986_ = ~new_C9968_ | new_C9978_;
  assign new_C9987_ = new_C9968_ & new_C9978_;
  assign new_C9988_ = ~new_C9968_ & ~new_C9978_;
  assign new_C9989_ = new_D11_ | new_D10_;
  assign new_C9990_ = new_C9956_ | new_C9989_;
  assign new_C9991_ = new_D15_ | new_D14_;
  assign new_C9992_ = ~new_C9956_ & new_C9991_;
  assign new_C9993_ = new_D13_ | new_D12_;
  assign new_C9994_ = new_C9956_ & new_C9993_;
  assign new_C9995_ = new_C9954_ & ~new_C9964_;
  assign new_C9996_ = ~new_C9954_ & new_C9964_;
  assign new_C9997_ = ~new_C9953_ | ~new_C9978_;
  assign new_C9998_ = new_C9964_ & new_C9997_;
  assign new_C9999_ = ~new_C9964_ & ~new_C9998_;
  assign new_D1_ = new_C9964_ | new_C9997_;
  assign new_D2_ = ~new_C9954_ & new_C9955_;
  assign new_D3_ = new_C9954_ & ~new_C9955_;
  assign new_D4_ = new_C9971_ | new_D9_;
  assign new_D5_ = ~new_C9971_ & ~new_D8_;
  assign new_D6_ = new_C9954_ | new_C9971_;
  assign new_D7_ = new_C9954_ | new_C9955_;
  assign new_D8_ = new_C9971_ & new_D9_;
  assign new_D9_ = ~new_C9953_ | ~new_C9978_;
  assign new_D10_ = new_C9986_ & new_D7_;
  assign new_D11_ = ~new_C9986_ & ~new_D7_;
  assign new_D12_ = new_D16_ | new_D17_;
  assign new_D13_ = ~new_C9957_ & new_C9971_;
  assign new_D14_ = new_D18_ | new_D19_;
  assign new_D15_ = new_C9957_ & new_C9971_;
  assign new_D16_ = ~new_C9957_ & ~new_C9971_;
  assign new_D17_ = new_C9957_ & ~new_C9971_;
  assign new_D18_ = new_C9957_ & ~new_C9971_;
  assign new_D19_ = ~new_C9957_ & new_C9971_;
  assign new_D20_ = new_D8605_;
  assign new_D21_ = new_D8672_;
  assign new_D22_ = new_D8739_;
  assign new_D23_ = new_D8806_;
  assign new_D24_ = new_D8873_;
  assign new_D25_ = new_D8940_;
  assign new_D26_ = new_D33_ & new_D32_;
  assign new_D27_ = new_D35_ | new_D34_;
  assign new_D28_ = new_D37_ | new_D36_;
  assign new_D29_ = new_D39_ & new_D38_;
  assign new_D30_ = new_D39_ & new_D40_;
  assign new_D31_ = new_D32_ | new_D41_;
  assign new_D32_ = new_D21_ | new_D44_;
  assign new_D33_ = new_D43_ | new_D42_;
  assign new_D34_ = new_D48_ & new_D47_;
  assign new_D35_ = new_D46_ & new_D45_;
  assign new_D36_ = new_D51_ | new_D50_;
  assign new_D37_ = new_D46_ & new_D49_;
  assign new_D38_ = new_D21_ | new_D54_;
  assign new_D39_ = new_D53_ | new_D52_;
  assign new_D40_ = new_D56_ | new_D55_;
  assign new_D41_ = ~new_D32_ & new_D58_;
  assign new_D42_ = ~new_D34_ & new_D46_;
  assign new_D43_ = new_D34_ & ~new_D46_;
  assign new_D44_ = new_D20_ & ~new_D21_;
  assign new_D45_ = ~new_D67_ | ~new_D68_;
  assign new_D46_ = new_D60_ | new_D62_;
  assign new_D47_ = new_D70_ | new_D69_;
  assign new_D48_ = new_D64_ | new_D63_;
  assign new_D49_ = ~new_D72_ | ~new_D71_;
  assign new_D50_ = ~new_D73_ & new_D74_;
  assign new_D51_ = new_D73_ & ~new_D74_;
  assign new_D52_ = ~new_D20_ & new_D21_;
  assign new_D53_ = new_D20_ & ~new_D21_;
  assign new_D54_ = ~new_D36_ | new_D46_;
  assign new_D55_ = new_D36_ & new_D46_;
  assign new_D56_ = ~new_D36_ & ~new_D46_;
  assign new_D57_ = new_D78_ | new_D77_;
  assign new_D58_ = new_D24_ | new_D57_;
  assign new_D59_ = new_D82_ | new_D81_;
  assign new_D60_ = ~new_D24_ & new_D59_;
  assign new_D61_ = new_D80_ | new_D79_;
  assign new_D62_ = new_D24_ & new_D61_;
  assign new_D63_ = new_D22_ & ~new_D32_;
  assign new_D64_ = ~new_D22_ & new_D32_;
  assign new_D65_ = ~new_D21_ | ~new_D46_;
  assign new_D66_ = new_D32_ & new_D65_;
  assign new_D67_ = ~new_D32_ & ~new_D66_;
  assign new_D68_ = new_D32_ | new_D65_;
  assign new_D69_ = ~new_D22_ & new_D23_;
  assign new_D70_ = new_D22_ & ~new_D23_;
  assign new_D71_ = new_D39_ | new_D76_;
  assign new_D72_ = ~new_D39_ & ~new_D75_;
  assign new_D73_ = new_D22_ | new_D39_;
  assign new_D74_ = new_D22_ | new_D23_;
  assign new_D75_ = new_D39_ & new_D76_;
  assign new_D76_ = ~new_D21_ | ~new_D46_;
  assign new_D77_ = new_D54_ & new_D74_;
  assign new_D78_ = ~new_D54_ & ~new_D74_;
  assign new_D79_ = new_D83_ | new_D84_;
  assign new_D80_ = ~new_D25_ & new_D39_;
  assign new_D81_ = new_D85_ | new_D86_;
  assign new_D82_ = new_D25_ & new_D39_;
  assign new_D83_ = ~new_D25_ & ~new_D39_;
  assign new_D84_ = new_D25_ & ~new_D39_;
  assign new_D85_ = new_D25_ & ~new_D39_;
  assign new_D86_ = ~new_D25_ & new_D39_;
  assign new_D87_ = new_D9007_;
  assign new_D88_ = new_D9074_;
  assign new_D89_ = new_D9141_;
  assign new_D90_ = new_D9208_;
  assign new_D91_ = new_D9275_;
  assign new_D92_ = new_D9342_;
  assign new_D93_ = new_D100_ & new_D99_;
  assign new_D94_ = new_D102_ | new_D101_;
  assign new_D95_ = new_D104_ | new_D103_;
  assign new_D96_ = new_D106_ & new_D105_;
  assign new_D97_ = new_D106_ & new_D107_;
  assign new_D98_ = new_D99_ | new_D108_;
  assign new_D99_ = new_D88_ | new_D111_;
  assign new_D100_ = new_D110_ | new_D109_;
  assign new_D101_ = new_D115_ & new_D114_;
  assign new_D102_ = new_D113_ & new_D112_;
  assign new_D103_ = new_D118_ | new_D117_;
  assign new_D104_ = new_D113_ & new_D116_;
  assign new_D105_ = new_D88_ | new_D121_;
  assign new_D106_ = new_D120_ | new_D119_;
  assign new_D107_ = new_D123_ | new_D122_;
  assign new_D108_ = ~new_D99_ & new_D125_;
  assign new_D109_ = ~new_D101_ & new_D113_;
  assign new_D110_ = new_D101_ & ~new_D113_;
  assign new_D111_ = new_D87_ & ~new_D88_;
  assign new_D112_ = ~new_D134_ | ~new_D135_;
  assign new_D113_ = new_D127_ | new_D129_;
  assign new_D114_ = new_D137_ | new_D136_;
  assign new_D115_ = new_D131_ | new_D130_;
  assign new_D116_ = ~new_D139_ | ~new_D138_;
  assign new_D117_ = ~new_D140_ & new_D141_;
  assign new_D118_ = new_D140_ & ~new_D141_;
  assign new_D119_ = ~new_D87_ & new_D88_;
  assign new_D120_ = new_D87_ & ~new_D88_;
  assign new_D121_ = ~new_D103_ | new_D113_;
  assign new_D122_ = new_D103_ & new_D113_;
  assign new_D123_ = ~new_D103_ & ~new_D113_;
  assign new_D124_ = new_D145_ | new_D144_;
  assign new_D125_ = new_D91_ | new_D124_;
  assign new_D126_ = new_D149_ | new_D148_;
  assign new_D127_ = ~new_D91_ & new_D126_;
  assign new_D128_ = new_D147_ | new_D146_;
  assign new_D129_ = new_D91_ & new_D128_;
  assign new_D130_ = new_D89_ & ~new_D99_;
  assign new_D131_ = ~new_D89_ & new_D99_;
  assign new_D132_ = ~new_D88_ | ~new_D113_;
  assign new_D133_ = new_D99_ & new_D132_;
  assign new_D134_ = ~new_D99_ & ~new_D133_;
  assign new_D135_ = new_D99_ | new_D132_;
  assign new_D136_ = ~new_D89_ & new_D90_;
  assign new_D137_ = new_D89_ & ~new_D90_;
  assign new_D138_ = new_D106_ | new_D143_;
  assign new_D139_ = ~new_D106_ & ~new_D142_;
  assign new_D140_ = new_D89_ | new_D106_;
  assign new_D141_ = new_D89_ | new_D90_;
  assign new_D142_ = new_D106_ & new_D143_;
  assign new_D143_ = ~new_D88_ | ~new_D113_;
  assign new_D144_ = new_D121_ & new_D141_;
  assign new_D145_ = ~new_D121_ & ~new_D141_;
  assign new_D146_ = new_D150_ | new_D151_;
  assign new_D147_ = ~new_D92_ & new_D106_;
  assign new_D148_ = new_D152_ | new_D153_;
  assign new_D149_ = new_D92_ & new_D106_;
  assign new_D150_ = ~new_D92_ & ~new_D106_;
  assign new_D151_ = new_D92_ & ~new_D106_;
  assign new_D152_ = new_D92_ & ~new_D106_;
  assign new_D153_ = ~new_D92_ & new_D106_;
  assign new_D154_ = new_D9409_;
  assign new_D155_ = new_D9476_;
  assign new_D156_ = new_D9543_;
  assign new_D157_ = new_D9610_;
  assign new_D158_ = new_D9677_;
  assign new_D159_ = new_D9744_;
  assign new_D160_ = new_D167_ & new_D166_;
  assign new_D161_ = new_D169_ | new_D168_;
  assign new_D162_ = new_D171_ | new_D170_;
  assign new_D163_ = new_D173_ & new_D172_;
  assign new_D164_ = new_D173_ & new_D174_;
  assign new_D165_ = new_D166_ | new_D175_;
  assign new_D166_ = new_D155_ | new_D178_;
  assign new_D167_ = new_D177_ | new_D176_;
  assign new_D168_ = new_D182_ & new_D181_;
  assign new_D169_ = new_D180_ & new_D179_;
  assign new_D170_ = new_D185_ | new_D184_;
  assign new_D171_ = new_D180_ & new_D183_;
  assign new_D172_ = new_D155_ | new_D188_;
  assign new_D173_ = new_D187_ | new_D186_;
  assign new_D174_ = new_D190_ | new_D189_;
  assign new_D175_ = ~new_D166_ & new_D192_;
  assign new_D176_ = ~new_D168_ & new_D180_;
  assign new_D177_ = new_D168_ & ~new_D180_;
  assign new_D178_ = new_D154_ & ~new_D155_;
  assign new_D179_ = ~new_D201_ | ~new_D202_;
  assign new_D180_ = new_D194_ | new_D196_;
  assign new_D181_ = new_D204_ | new_D203_;
  assign new_D182_ = new_D198_ | new_D197_;
  assign new_D183_ = ~new_D206_ | ~new_D205_;
  assign new_D184_ = ~new_D207_ & new_D208_;
  assign new_D185_ = new_D207_ & ~new_D208_;
  assign new_D186_ = ~new_D154_ & new_D155_;
  assign new_D187_ = new_D154_ & ~new_D155_;
  assign new_D188_ = ~new_D170_ | new_D180_;
  assign new_D189_ = new_D170_ & new_D180_;
  assign new_D190_ = ~new_D170_ & ~new_D180_;
  assign new_D191_ = new_D212_ | new_D211_;
  assign new_D192_ = new_D158_ | new_D191_;
  assign new_D193_ = new_D216_ | new_D215_;
  assign new_D194_ = ~new_D158_ & new_D193_;
  assign new_D195_ = new_D214_ | new_D213_;
  assign new_D196_ = new_D158_ & new_D195_;
  assign new_D197_ = new_D156_ & ~new_D166_;
  assign new_D198_ = ~new_D156_ & new_D166_;
  assign new_D199_ = ~new_D155_ | ~new_D180_;
  assign new_D200_ = new_D166_ & new_D199_;
  assign new_D201_ = ~new_D166_ & ~new_D200_;
  assign new_D202_ = new_D166_ | new_D199_;
  assign new_D203_ = ~new_D156_ & new_D157_;
  assign new_D204_ = new_D156_ & ~new_D157_;
  assign new_D205_ = new_D173_ | new_D210_;
  assign new_D206_ = ~new_D173_ & ~new_D209_;
  assign new_D207_ = new_D156_ | new_D173_;
  assign new_D208_ = new_D156_ | new_D157_;
  assign new_D209_ = new_D173_ & new_D210_;
  assign new_D210_ = ~new_D155_ | ~new_D180_;
  assign new_D211_ = new_D188_ & new_D208_;
  assign new_D212_ = ~new_D188_ & ~new_D208_;
  assign new_D213_ = new_D217_ | new_D218_;
  assign new_D214_ = ~new_D159_ & new_D173_;
  assign new_D215_ = new_D219_ | new_D220_;
  assign new_D216_ = new_D159_ & new_D173_;
  assign new_D217_ = ~new_D159_ & ~new_D173_;
  assign new_D218_ = new_D159_ & ~new_D173_;
  assign new_D219_ = new_D159_ & ~new_D173_;
  assign new_D220_ = ~new_D159_ & new_D173_;
  assign new_D221_ = new_D9811_;
  assign new_D222_ = new_D9878_;
  assign new_D223_ = new_D9945_;
  assign new_D224_ = new_E13_;
  assign new_D225_ = new_E80_;
  assign new_D226_ = new_E147_;
  assign new_D227_ = new_D234_ & new_D233_;
  assign new_D228_ = new_D236_ | new_D235_;
  assign new_D229_ = new_D238_ | new_D237_;
  assign new_D230_ = new_D240_ & new_D239_;
  assign new_D231_ = new_D240_ & new_D241_;
  assign new_D232_ = new_D233_ | new_D242_;
  assign new_D233_ = new_D222_ | new_D245_;
  assign new_D234_ = new_D244_ | new_D243_;
  assign new_D235_ = new_D249_ & new_D248_;
  assign new_D236_ = new_D247_ & new_D246_;
  assign new_D237_ = new_D252_ | new_D251_;
  assign new_D238_ = new_D247_ & new_D250_;
  assign new_D239_ = new_D222_ | new_D255_;
  assign new_D240_ = new_D254_ | new_D253_;
  assign new_D241_ = new_D257_ | new_D256_;
  assign new_D242_ = ~new_D233_ & new_D259_;
  assign new_D243_ = ~new_D235_ & new_D247_;
  assign new_D244_ = new_D235_ & ~new_D247_;
  assign new_D245_ = new_D221_ & ~new_D222_;
  assign new_D246_ = ~new_D268_ | ~new_D269_;
  assign new_D247_ = new_D261_ | new_D263_;
  assign new_D248_ = new_D271_ | new_D270_;
  assign new_D249_ = new_D265_ | new_D264_;
  assign new_D250_ = ~new_D273_ | ~new_D272_;
  assign new_D251_ = ~new_D274_ & new_D275_;
  assign new_D252_ = new_D274_ & ~new_D275_;
  assign new_D253_ = ~new_D221_ & new_D222_;
  assign new_D254_ = new_D221_ & ~new_D222_;
  assign new_D255_ = ~new_D237_ | new_D247_;
  assign new_D256_ = new_D237_ & new_D247_;
  assign new_D257_ = ~new_D237_ & ~new_D247_;
  assign new_D258_ = new_D279_ | new_D278_;
  assign new_D259_ = new_D225_ | new_D258_;
  assign new_D260_ = new_D283_ | new_D282_;
  assign new_D261_ = ~new_D225_ & new_D260_;
  assign new_D262_ = new_D281_ | new_D280_;
  assign new_D263_ = new_D225_ & new_D262_;
  assign new_D264_ = new_D223_ & ~new_D233_;
  assign new_D265_ = ~new_D223_ & new_D233_;
  assign new_D266_ = ~new_D222_ | ~new_D247_;
  assign new_D267_ = new_D233_ & new_D266_;
  assign new_D268_ = ~new_D233_ & ~new_D267_;
  assign new_D269_ = new_D233_ | new_D266_;
  assign new_D270_ = ~new_D223_ & new_D224_;
  assign new_D271_ = new_D223_ & ~new_D224_;
  assign new_D272_ = new_D240_ | new_D277_;
  assign new_D273_ = ~new_D240_ & ~new_D276_;
  assign new_D274_ = new_D223_ | new_D240_;
  assign new_D275_ = new_D223_ | new_D224_;
  assign new_D276_ = new_D240_ & new_D277_;
  assign new_D277_ = ~new_D222_ | ~new_D247_;
  assign new_D278_ = new_D255_ & new_D275_;
  assign new_D279_ = ~new_D255_ & ~new_D275_;
  assign new_D280_ = new_D284_ | new_D285_;
  assign new_D281_ = ~new_D226_ & new_D240_;
  assign new_D282_ = new_D286_ | new_D287_;
  assign new_D283_ = new_D226_ & new_D240_;
  assign new_D284_ = ~new_D226_ & ~new_D240_;
  assign new_D285_ = new_D226_ & ~new_D240_;
  assign new_D286_ = new_D226_ & ~new_D240_;
  assign new_D287_ = ~new_D226_ & new_D240_;
  assign new_D288_ = new_E214_;
  assign new_D289_ = new_E281_;
  assign new_D290_ = new_E348_;
  assign new_D291_ = new_E415_;
  assign new_D292_ = new_E482_;
  assign new_D293_ = new_E549_;
  assign new_D294_ = new_D301_ & new_D300_;
  assign new_D295_ = new_D303_ | new_D302_;
  assign new_D296_ = new_D305_ | new_D304_;
  assign new_D297_ = new_D307_ & new_D306_;
  assign new_D298_ = new_D307_ & new_D308_;
  assign new_D299_ = new_D300_ | new_D309_;
  assign new_D300_ = new_D289_ | new_D312_;
  assign new_D301_ = new_D311_ | new_D310_;
  assign new_D302_ = new_D316_ & new_D315_;
  assign new_D303_ = new_D314_ & new_D313_;
  assign new_D304_ = new_D319_ | new_D318_;
  assign new_D305_ = new_D314_ & new_D317_;
  assign new_D306_ = new_D289_ | new_D322_;
  assign new_D307_ = new_D321_ | new_D320_;
  assign new_D308_ = new_D324_ | new_D323_;
  assign new_D309_ = ~new_D300_ & new_D326_;
  assign new_D310_ = ~new_D302_ & new_D314_;
  assign new_D311_ = new_D302_ & ~new_D314_;
  assign new_D312_ = new_D288_ & ~new_D289_;
  assign new_D313_ = ~new_D335_ | ~new_D336_;
  assign new_D314_ = new_D328_ | new_D330_;
  assign new_D315_ = new_D338_ | new_D337_;
  assign new_D316_ = new_D332_ | new_D331_;
  assign new_D317_ = ~new_D340_ | ~new_D339_;
  assign new_D318_ = ~new_D341_ & new_D342_;
  assign new_D319_ = new_D341_ & ~new_D342_;
  assign new_D320_ = ~new_D288_ & new_D289_;
  assign new_D321_ = new_D288_ & ~new_D289_;
  assign new_D322_ = ~new_D304_ | new_D314_;
  assign new_D323_ = new_D304_ & new_D314_;
  assign new_D324_ = ~new_D304_ & ~new_D314_;
  assign new_D325_ = new_D346_ | new_D345_;
  assign new_D326_ = new_D292_ | new_D325_;
  assign new_D327_ = new_D350_ | new_D349_;
  assign new_D328_ = ~new_D292_ & new_D327_;
  assign new_D329_ = new_D348_ | new_D347_;
  assign new_D330_ = new_D292_ & new_D329_;
  assign new_D331_ = new_D290_ & ~new_D300_;
  assign new_D332_ = ~new_D290_ & new_D300_;
  assign new_D333_ = ~new_D289_ | ~new_D314_;
  assign new_D334_ = new_D300_ & new_D333_;
  assign new_D335_ = ~new_D300_ & ~new_D334_;
  assign new_D336_ = new_D300_ | new_D333_;
  assign new_D337_ = ~new_D290_ & new_D291_;
  assign new_D338_ = new_D290_ & ~new_D291_;
  assign new_D339_ = new_D307_ | new_D344_;
  assign new_D340_ = ~new_D307_ & ~new_D343_;
  assign new_D341_ = new_D290_ | new_D307_;
  assign new_D342_ = new_D290_ | new_D291_;
  assign new_D343_ = new_D307_ & new_D344_;
  assign new_D344_ = ~new_D289_ | ~new_D314_;
  assign new_D345_ = new_D322_ & new_D342_;
  assign new_D346_ = ~new_D322_ & ~new_D342_;
  assign new_D347_ = new_D351_ | new_D352_;
  assign new_D348_ = ~new_D293_ & new_D307_;
  assign new_D349_ = new_D353_ | new_D354_;
  assign new_D350_ = new_D293_ & new_D307_;
  assign new_D351_ = ~new_D293_ & ~new_D307_;
  assign new_D352_ = new_D293_ & ~new_D307_;
  assign new_D353_ = new_D293_ & ~new_D307_;
  assign new_D354_ = ~new_D293_ & new_D307_;
  assign new_D355_ = new_E616_;
  assign new_D356_ = new_E683_;
  assign new_D357_ = new_E750_;
  assign new_D358_ = new_E817_;
  assign new_D359_ = new_E884_;
  assign new_D360_ = new_E951_;
  assign new_D361_ = new_D368_ & new_D367_;
  assign new_D362_ = new_D370_ | new_D369_;
  assign new_D363_ = new_D372_ | new_D371_;
  assign new_D364_ = new_D374_ & new_D373_;
  assign new_D365_ = new_D374_ & new_D375_;
  assign new_D366_ = new_D367_ | new_D376_;
  assign new_D367_ = new_D356_ | new_D379_;
  assign new_D368_ = new_D378_ | new_D377_;
  assign new_D369_ = new_D383_ & new_D382_;
  assign new_D370_ = new_D381_ & new_D380_;
  assign new_D371_ = new_D386_ | new_D385_;
  assign new_D372_ = new_D381_ & new_D384_;
  assign new_D373_ = new_D356_ | new_D389_;
  assign new_D374_ = new_D388_ | new_D387_;
  assign new_D375_ = new_D391_ | new_D390_;
  assign new_D376_ = ~new_D367_ & new_D393_;
  assign new_D377_ = ~new_D369_ & new_D381_;
  assign new_D378_ = new_D369_ & ~new_D381_;
  assign new_D379_ = new_D355_ & ~new_D356_;
  assign new_D380_ = ~new_D402_ | ~new_D403_;
  assign new_D381_ = new_D395_ | new_D397_;
  assign new_D382_ = new_D405_ | new_D404_;
  assign new_D383_ = new_D399_ | new_D398_;
  assign new_D384_ = ~new_D407_ | ~new_D406_;
  assign new_D385_ = ~new_D408_ & new_D409_;
  assign new_D386_ = new_D408_ & ~new_D409_;
  assign new_D387_ = ~new_D355_ & new_D356_;
  assign new_D388_ = new_D355_ & ~new_D356_;
  assign new_D389_ = ~new_D371_ | new_D381_;
  assign new_D390_ = new_D371_ & new_D381_;
  assign new_D391_ = ~new_D371_ & ~new_D381_;
  assign new_D392_ = new_D413_ | new_D412_;
  assign new_D393_ = new_D359_ | new_D392_;
  assign new_D394_ = new_D417_ | new_D416_;
  assign new_D395_ = ~new_D359_ & new_D394_;
  assign new_D396_ = new_D415_ | new_D414_;
  assign new_D397_ = new_D359_ & new_D396_;
  assign new_D398_ = new_D357_ & ~new_D367_;
  assign new_D399_ = ~new_D357_ & new_D367_;
  assign new_D400_ = ~new_D356_ | ~new_D381_;
  assign new_D401_ = new_D367_ & new_D400_;
  assign new_D402_ = ~new_D367_ & ~new_D401_;
  assign new_D403_ = new_D367_ | new_D400_;
  assign new_D404_ = ~new_D357_ & new_D358_;
  assign new_D405_ = new_D357_ & ~new_D358_;
  assign new_D406_ = new_D374_ | new_D411_;
  assign new_D407_ = ~new_D374_ & ~new_D410_;
  assign new_D408_ = new_D357_ | new_D374_;
  assign new_D409_ = new_D357_ | new_D358_;
  assign new_D410_ = new_D374_ & new_D411_;
  assign new_D411_ = ~new_D356_ | ~new_D381_;
  assign new_D412_ = new_D389_ & new_D409_;
  assign new_D413_ = ~new_D389_ & ~new_D409_;
  assign new_D414_ = new_D418_ | new_D419_;
  assign new_D415_ = ~new_D360_ & new_D374_;
  assign new_D416_ = new_D420_ | new_D421_;
  assign new_D417_ = new_D360_ & new_D374_;
  assign new_D418_ = ~new_D360_ & ~new_D374_;
  assign new_D419_ = new_D360_ & ~new_D374_;
  assign new_D420_ = new_D360_ & ~new_D374_;
  assign new_D421_ = ~new_D360_ & new_D374_;
  assign new_D422_ = new_E1018_;
  assign new_D423_ = new_E1085_;
  assign new_D424_ = new_E1152_;
  assign new_D425_ = new_E1219_;
  assign new_D426_ = new_E1286_;
  assign new_D427_ = new_E1353_;
  assign new_D428_ = new_D435_ & new_D434_;
  assign new_D429_ = new_D437_ | new_D436_;
  assign new_D430_ = new_D439_ | new_D438_;
  assign new_D431_ = new_D441_ & new_D440_;
  assign new_D432_ = new_D441_ & new_D442_;
  assign new_D433_ = new_D434_ | new_D443_;
  assign new_D434_ = new_D423_ | new_D446_;
  assign new_D435_ = new_D445_ | new_D444_;
  assign new_D436_ = new_D450_ & new_D449_;
  assign new_D437_ = new_D448_ & new_D447_;
  assign new_D438_ = new_D453_ | new_D452_;
  assign new_D439_ = new_D448_ & new_D451_;
  assign new_D440_ = new_D423_ | new_D456_;
  assign new_D441_ = new_D455_ | new_D454_;
  assign new_D442_ = new_D458_ | new_D457_;
  assign new_D443_ = ~new_D434_ & new_D460_;
  assign new_D444_ = ~new_D436_ & new_D448_;
  assign new_D445_ = new_D436_ & ~new_D448_;
  assign new_D446_ = new_D422_ & ~new_D423_;
  assign new_D447_ = ~new_D469_ | ~new_D470_;
  assign new_D448_ = new_D462_ | new_D464_;
  assign new_D449_ = new_D472_ | new_D471_;
  assign new_D450_ = new_D466_ | new_D465_;
  assign new_D451_ = ~new_D474_ | ~new_D473_;
  assign new_D452_ = ~new_D475_ & new_D476_;
  assign new_D453_ = new_D475_ & ~new_D476_;
  assign new_D454_ = ~new_D422_ & new_D423_;
  assign new_D455_ = new_D422_ & ~new_D423_;
  assign new_D456_ = ~new_D438_ | new_D448_;
  assign new_D457_ = new_D438_ & new_D448_;
  assign new_D458_ = ~new_D438_ & ~new_D448_;
  assign new_D459_ = new_D480_ | new_D479_;
  assign new_D460_ = new_D426_ | new_D459_;
  assign new_D461_ = new_D484_ | new_D483_;
  assign new_D462_ = ~new_D426_ & new_D461_;
  assign new_D463_ = new_D482_ | new_D481_;
  assign new_D464_ = new_D426_ & new_D463_;
  assign new_D465_ = new_D424_ & ~new_D434_;
  assign new_D466_ = ~new_D424_ & new_D434_;
  assign new_D467_ = ~new_D423_ | ~new_D448_;
  assign new_D468_ = new_D434_ & new_D467_;
  assign new_D469_ = ~new_D434_ & ~new_D468_;
  assign new_D470_ = new_D434_ | new_D467_;
  assign new_D471_ = ~new_D424_ & new_D425_;
  assign new_D472_ = new_D424_ & ~new_D425_;
  assign new_D473_ = new_D441_ | new_D478_;
  assign new_D474_ = ~new_D441_ & ~new_D477_;
  assign new_D475_ = new_D424_ | new_D441_;
  assign new_D476_ = new_D424_ | new_D425_;
  assign new_D477_ = new_D441_ & new_D478_;
  assign new_D478_ = ~new_D423_ | ~new_D448_;
  assign new_D479_ = new_D456_ & new_D476_;
  assign new_D480_ = ~new_D456_ & ~new_D476_;
  assign new_D481_ = new_D485_ | new_D486_;
  assign new_D482_ = ~new_D427_ & new_D441_;
  assign new_D483_ = new_D487_ | new_D488_;
  assign new_D484_ = new_D427_ & new_D441_;
  assign new_D485_ = ~new_D427_ & ~new_D441_;
  assign new_D486_ = new_D427_ & ~new_D441_;
  assign new_D487_ = new_D427_ & ~new_D441_;
  assign new_D488_ = ~new_D427_ & new_D441_;
  assign new_D489_ = new_E1420_;
  assign new_D490_ = new_E1487_;
  assign new_D491_ = new_E1554_;
  assign new_D492_ = new_E1621_;
  assign new_D493_ = new_E1688_;
  assign new_D494_ = new_E1755_;
  assign new_D495_ = new_D502_ & new_D501_;
  assign new_D496_ = new_D504_ | new_D503_;
  assign new_D497_ = new_D506_ | new_D505_;
  assign new_D498_ = new_D508_ & new_D507_;
  assign new_D499_ = new_D508_ & new_D509_;
  assign new_D500_ = new_D501_ | new_D510_;
  assign new_D501_ = new_D490_ | new_D513_;
  assign new_D502_ = new_D512_ | new_D511_;
  assign new_D503_ = new_D517_ & new_D516_;
  assign new_D504_ = new_D515_ & new_D514_;
  assign new_D505_ = new_D520_ | new_D519_;
  assign new_D506_ = new_D515_ & new_D518_;
  assign new_D507_ = new_D490_ | new_D523_;
  assign new_D508_ = new_D522_ | new_D521_;
  assign new_D509_ = new_D525_ | new_D524_;
  assign new_D510_ = ~new_D501_ & new_D527_;
  assign new_D511_ = ~new_D503_ & new_D515_;
  assign new_D512_ = new_D503_ & ~new_D515_;
  assign new_D513_ = new_D489_ & ~new_D490_;
  assign new_D514_ = ~new_D536_ | ~new_D537_;
  assign new_D515_ = new_D529_ | new_D531_;
  assign new_D516_ = new_D539_ | new_D538_;
  assign new_D517_ = new_D533_ | new_D532_;
  assign new_D518_ = ~new_D541_ | ~new_D540_;
  assign new_D519_ = ~new_D542_ & new_D543_;
  assign new_D520_ = new_D542_ & ~new_D543_;
  assign new_D521_ = ~new_D489_ & new_D490_;
  assign new_D522_ = new_D489_ & ~new_D490_;
  assign new_D523_ = ~new_D505_ | new_D515_;
  assign new_D524_ = new_D505_ & new_D515_;
  assign new_D525_ = ~new_D505_ & ~new_D515_;
  assign new_D526_ = new_D547_ | new_D546_;
  assign new_D527_ = new_D493_ | new_D526_;
  assign new_D528_ = new_D551_ | new_D550_;
  assign new_D529_ = ~new_D493_ & new_D528_;
  assign new_D530_ = new_D549_ | new_D548_;
  assign new_D531_ = new_D493_ & new_D530_;
  assign new_D532_ = new_D491_ & ~new_D501_;
  assign new_D533_ = ~new_D491_ & new_D501_;
  assign new_D534_ = ~new_D490_ | ~new_D515_;
  assign new_D535_ = new_D501_ & new_D534_;
  assign new_D536_ = ~new_D501_ & ~new_D535_;
  assign new_D537_ = new_D501_ | new_D534_;
  assign new_D538_ = ~new_D491_ & new_D492_;
  assign new_D539_ = new_D491_ & ~new_D492_;
  assign new_D540_ = new_D508_ | new_D545_;
  assign new_D541_ = ~new_D508_ & ~new_D544_;
  assign new_D542_ = new_D491_ | new_D508_;
  assign new_D543_ = new_D491_ | new_D492_;
  assign new_D544_ = new_D508_ & new_D545_;
  assign new_D545_ = ~new_D490_ | ~new_D515_;
  assign new_D546_ = new_D523_ & new_D543_;
  assign new_D547_ = ~new_D523_ & ~new_D543_;
  assign new_D548_ = new_D552_ | new_D553_;
  assign new_D549_ = ~new_D494_ & new_D508_;
  assign new_D550_ = new_D554_ | new_D555_;
  assign new_D551_ = new_D494_ & new_D508_;
  assign new_D552_ = ~new_D494_ & ~new_D508_;
  assign new_D553_ = new_D494_ & ~new_D508_;
  assign new_D554_ = new_D494_ & ~new_D508_;
  assign new_D555_ = ~new_D494_ & new_D508_;
  assign new_D556_ = new_E1822_;
  assign new_D557_ = new_E1889_;
  assign new_D558_ = new_E1956_;
  assign new_D559_ = new_E2023_;
  assign new_D560_ = new_E2090_;
  assign new_D561_ = new_E2157_;
  assign new_D562_ = new_D569_ & new_D568_;
  assign new_D563_ = new_D571_ | new_D570_;
  assign new_D564_ = new_D573_ | new_D572_;
  assign new_D565_ = new_D575_ & new_D574_;
  assign new_D566_ = new_D575_ & new_D576_;
  assign new_D567_ = new_D568_ | new_D577_;
  assign new_D568_ = new_D557_ | new_D580_;
  assign new_D569_ = new_D579_ | new_D578_;
  assign new_D570_ = new_D584_ & new_D583_;
  assign new_D571_ = new_D582_ & new_D581_;
  assign new_D572_ = new_D587_ | new_D586_;
  assign new_D573_ = new_D582_ & new_D585_;
  assign new_D574_ = new_D557_ | new_D590_;
  assign new_D575_ = new_D589_ | new_D588_;
  assign new_D576_ = new_D592_ | new_D591_;
  assign new_D577_ = ~new_D568_ & new_D594_;
  assign new_D578_ = ~new_D570_ & new_D582_;
  assign new_D579_ = new_D570_ & ~new_D582_;
  assign new_D580_ = new_D556_ & ~new_D557_;
  assign new_D581_ = ~new_D603_ | ~new_D604_;
  assign new_D582_ = new_D596_ | new_D598_;
  assign new_D583_ = new_D606_ | new_D605_;
  assign new_D584_ = new_D600_ | new_D599_;
  assign new_D585_ = ~new_D608_ | ~new_D607_;
  assign new_D586_ = ~new_D609_ & new_D610_;
  assign new_D587_ = new_D609_ & ~new_D610_;
  assign new_D588_ = ~new_D556_ & new_D557_;
  assign new_D589_ = new_D556_ & ~new_D557_;
  assign new_D590_ = ~new_D572_ | new_D582_;
  assign new_D591_ = new_D572_ & new_D582_;
  assign new_D592_ = ~new_D572_ & ~new_D582_;
  assign new_D593_ = new_D614_ | new_D613_;
  assign new_D594_ = new_D560_ | new_D593_;
  assign new_D595_ = new_D618_ | new_D617_;
  assign new_D596_ = ~new_D560_ & new_D595_;
  assign new_D597_ = new_D616_ | new_D615_;
  assign new_D598_ = new_D560_ & new_D597_;
  assign new_D599_ = new_D558_ & ~new_D568_;
  assign new_D600_ = ~new_D558_ & new_D568_;
  assign new_D601_ = ~new_D557_ | ~new_D582_;
  assign new_D602_ = new_D568_ & new_D601_;
  assign new_D603_ = ~new_D568_ & ~new_D602_;
  assign new_D604_ = new_D568_ | new_D601_;
  assign new_D605_ = ~new_D558_ & new_D559_;
  assign new_D606_ = new_D558_ & ~new_D559_;
  assign new_D607_ = new_D575_ | new_D612_;
  assign new_D608_ = ~new_D575_ & ~new_D611_;
  assign new_D609_ = new_D558_ | new_D575_;
  assign new_D610_ = new_D558_ | new_D559_;
  assign new_D611_ = new_D575_ & new_D612_;
  assign new_D612_ = ~new_D557_ | ~new_D582_;
  assign new_D613_ = new_D590_ & new_D610_;
  assign new_D614_ = ~new_D590_ & ~new_D610_;
  assign new_D615_ = new_D619_ | new_D620_;
  assign new_D616_ = ~new_D561_ & new_D575_;
  assign new_D617_ = new_D621_ | new_D622_;
  assign new_D618_ = new_D561_ & new_D575_;
  assign new_D619_ = ~new_D561_ & ~new_D575_;
  assign new_D620_ = new_D561_ & ~new_D575_;
  assign new_D621_ = new_D561_ & ~new_D575_;
  assign new_D622_ = ~new_D561_ & new_D575_;
  assign new_D623_ = new_E2224_;
  assign new_D624_ = new_E2291_;
  assign new_D625_ = new_E2358_;
  assign new_D626_ = new_E2425_;
  assign new_D627_ = new_E2492_;
  assign new_D628_ = new_E2559_;
  assign new_D629_ = new_D636_ & new_D635_;
  assign new_D630_ = new_D638_ | new_D637_;
  assign new_D631_ = new_D640_ | new_D639_;
  assign new_D632_ = new_D642_ & new_D641_;
  assign new_D633_ = new_D642_ & new_D643_;
  assign new_D634_ = new_D635_ | new_D644_;
  assign new_D635_ = new_D624_ | new_D647_;
  assign new_D636_ = new_D646_ | new_D645_;
  assign new_D637_ = new_D651_ & new_D650_;
  assign new_D638_ = new_D649_ & new_D648_;
  assign new_D639_ = new_D654_ | new_D653_;
  assign new_D640_ = new_D649_ & new_D652_;
  assign new_D641_ = new_D624_ | new_D657_;
  assign new_D642_ = new_D656_ | new_D655_;
  assign new_D643_ = new_D659_ | new_D658_;
  assign new_D644_ = ~new_D635_ & new_D661_;
  assign new_D645_ = ~new_D637_ & new_D649_;
  assign new_D646_ = new_D637_ & ~new_D649_;
  assign new_D647_ = new_D623_ & ~new_D624_;
  assign new_D648_ = ~new_D670_ | ~new_D671_;
  assign new_D649_ = new_D663_ | new_D665_;
  assign new_D650_ = new_D673_ | new_D672_;
  assign new_D651_ = new_D667_ | new_D666_;
  assign new_D652_ = ~new_D675_ | ~new_D674_;
  assign new_D653_ = ~new_D676_ & new_D677_;
  assign new_D654_ = new_D676_ & ~new_D677_;
  assign new_D655_ = ~new_D623_ & new_D624_;
  assign new_D656_ = new_D623_ & ~new_D624_;
  assign new_D657_ = ~new_D639_ | new_D649_;
  assign new_D658_ = new_D639_ & new_D649_;
  assign new_D659_ = ~new_D639_ & ~new_D649_;
  assign new_D660_ = new_D681_ | new_D680_;
  assign new_D661_ = new_D627_ | new_D660_;
  assign new_D662_ = new_D685_ | new_D684_;
  assign new_D663_ = ~new_D627_ & new_D662_;
  assign new_D664_ = new_D683_ | new_D682_;
  assign new_D665_ = new_D627_ & new_D664_;
  assign new_D666_ = new_D625_ & ~new_D635_;
  assign new_D667_ = ~new_D625_ & new_D635_;
  assign new_D668_ = ~new_D624_ | ~new_D649_;
  assign new_D669_ = new_D635_ & new_D668_;
  assign new_D670_ = ~new_D635_ & ~new_D669_;
  assign new_D671_ = new_D635_ | new_D668_;
  assign new_D672_ = ~new_D625_ & new_D626_;
  assign new_D673_ = new_D625_ & ~new_D626_;
  assign new_D674_ = new_D642_ | new_D679_;
  assign new_D675_ = ~new_D642_ & ~new_D678_;
  assign new_D676_ = new_D625_ | new_D642_;
  assign new_D677_ = new_D625_ | new_D626_;
  assign new_D678_ = new_D642_ & new_D679_;
  assign new_D679_ = ~new_D624_ | ~new_D649_;
  assign new_D680_ = new_D657_ & new_D677_;
  assign new_D681_ = ~new_D657_ & ~new_D677_;
  assign new_D682_ = new_D686_ | new_D687_;
  assign new_D683_ = ~new_D628_ & new_D642_;
  assign new_D684_ = new_D688_ | new_D689_;
  assign new_D685_ = new_D628_ & new_D642_;
  assign new_D686_ = ~new_D628_ & ~new_D642_;
  assign new_D687_ = new_D628_ & ~new_D642_;
  assign new_D688_ = new_D628_ & ~new_D642_;
  assign new_D689_ = ~new_D628_ & new_D642_;
  assign new_D690_ = new_E2626_;
  assign new_D691_ = new_E2693_;
  assign new_D692_ = new_E2760_;
  assign new_D693_ = new_E2827_;
  assign new_D694_ = new_E2894_;
  assign new_D695_ = new_E2961_;
  assign new_D696_ = new_D703_ & new_D702_;
  assign new_D697_ = new_D705_ | new_D704_;
  assign new_D698_ = new_D707_ | new_D706_;
  assign new_D699_ = new_D709_ & new_D708_;
  assign new_D700_ = new_D709_ & new_D710_;
  assign new_D701_ = new_D702_ | new_D711_;
  assign new_D702_ = new_D691_ | new_D714_;
  assign new_D703_ = new_D713_ | new_D712_;
  assign new_D704_ = new_D718_ & new_D717_;
  assign new_D705_ = new_D716_ & new_D715_;
  assign new_D706_ = new_D721_ | new_D720_;
  assign new_D707_ = new_D716_ & new_D719_;
  assign new_D708_ = new_D691_ | new_D724_;
  assign new_D709_ = new_D723_ | new_D722_;
  assign new_D710_ = new_D726_ | new_D725_;
  assign new_D711_ = ~new_D702_ & new_D728_;
  assign new_D712_ = ~new_D704_ & new_D716_;
  assign new_D713_ = new_D704_ & ~new_D716_;
  assign new_D714_ = new_D690_ & ~new_D691_;
  assign new_D715_ = ~new_D737_ | ~new_D738_;
  assign new_D716_ = new_D730_ | new_D732_;
  assign new_D717_ = new_D740_ | new_D739_;
  assign new_D718_ = new_D734_ | new_D733_;
  assign new_D719_ = ~new_D742_ | ~new_D741_;
  assign new_D720_ = ~new_D743_ & new_D744_;
  assign new_D721_ = new_D743_ & ~new_D744_;
  assign new_D722_ = ~new_D690_ & new_D691_;
  assign new_D723_ = new_D690_ & ~new_D691_;
  assign new_D724_ = ~new_D706_ | new_D716_;
  assign new_D725_ = new_D706_ & new_D716_;
  assign new_D726_ = ~new_D706_ & ~new_D716_;
  assign new_D727_ = new_D748_ | new_D747_;
  assign new_D728_ = new_D694_ | new_D727_;
  assign new_D729_ = new_D752_ | new_D751_;
  assign new_D730_ = ~new_D694_ & new_D729_;
  assign new_D731_ = new_D750_ | new_D749_;
  assign new_D732_ = new_D694_ & new_D731_;
  assign new_D733_ = new_D692_ & ~new_D702_;
  assign new_D734_ = ~new_D692_ & new_D702_;
  assign new_D735_ = ~new_D691_ | ~new_D716_;
  assign new_D736_ = new_D702_ & new_D735_;
  assign new_D737_ = ~new_D702_ & ~new_D736_;
  assign new_D738_ = new_D702_ | new_D735_;
  assign new_D739_ = ~new_D692_ & new_D693_;
  assign new_D740_ = new_D692_ & ~new_D693_;
  assign new_D741_ = new_D709_ | new_D746_;
  assign new_D742_ = ~new_D709_ & ~new_D745_;
  assign new_D743_ = new_D692_ | new_D709_;
  assign new_D744_ = new_D692_ | new_D693_;
  assign new_D745_ = new_D709_ & new_D746_;
  assign new_D746_ = ~new_D691_ | ~new_D716_;
  assign new_D747_ = new_D724_ & new_D744_;
  assign new_D748_ = ~new_D724_ & ~new_D744_;
  assign new_D749_ = new_D753_ | new_D754_;
  assign new_D750_ = ~new_D695_ & new_D709_;
  assign new_D751_ = new_D755_ | new_D756_;
  assign new_D752_ = new_D695_ & new_D709_;
  assign new_D753_ = ~new_D695_ & ~new_D709_;
  assign new_D754_ = new_D695_ & ~new_D709_;
  assign new_D755_ = new_D695_ & ~new_D709_;
  assign new_D756_ = ~new_D695_ & new_D709_;
  assign new_D757_ = new_E3028_;
  assign new_D758_ = new_E3095_;
  assign new_D759_ = new_E3162_;
  assign new_D760_ = new_E3229_;
  assign new_D761_ = new_E3296_;
  assign new_D762_ = new_E3363_;
  assign new_D763_ = new_D770_ & new_D769_;
  assign new_D764_ = new_D772_ | new_D771_;
  assign new_D765_ = new_D774_ | new_D773_;
  assign new_D766_ = new_D776_ & new_D775_;
  assign new_D767_ = new_D776_ & new_D777_;
  assign new_D768_ = new_D769_ | new_D778_;
  assign new_D769_ = new_D758_ | new_D781_;
  assign new_D770_ = new_D780_ | new_D779_;
  assign new_D771_ = new_D785_ & new_D784_;
  assign new_D772_ = new_D783_ & new_D782_;
  assign new_D773_ = new_D788_ | new_D787_;
  assign new_D774_ = new_D783_ & new_D786_;
  assign new_D775_ = new_D758_ | new_D791_;
  assign new_D776_ = new_D790_ | new_D789_;
  assign new_D777_ = new_D793_ | new_D792_;
  assign new_D778_ = ~new_D769_ & new_D795_;
  assign new_D779_ = ~new_D771_ & new_D783_;
  assign new_D780_ = new_D771_ & ~new_D783_;
  assign new_D781_ = new_D757_ & ~new_D758_;
  assign new_D782_ = ~new_D804_ | ~new_D805_;
  assign new_D783_ = new_D797_ | new_D799_;
  assign new_D784_ = new_D807_ | new_D806_;
  assign new_D785_ = new_D801_ | new_D800_;
  assign new_D786_ = ~new_D809_ | ~new_D808_;
  assign new_D787_ = ~new_D810_ & new_D811_;
  assign new_D788_ = new_D810_ & ~new_D811_;
  assign new_D789_ = ~new_D757_ & new_D758_;
  assign new_D790_ = new_D757_ & ~new_D758_;
  assign new_D791_ = ~new_D773_ | new_D783_;
  assign new_D792_ = new_D773_ & new_D783_;
  assign new_D793_ = ~new_D773_ & ~new_D783_;
  assign new_D794_ = new_D815_ | new_D814_;
  assign new_D795_ = new_D761_ | new_D794_;
  assign new_D796_ = new_D819_ | new_D818_;
  assign new_D797_ = ~new_D761_ & new_D796_;
  assign new_D798_ = new_D817_ | new_D816_;
  assign new_D799_ = new_D761_ & new_D798_;
  assign new_D800_ = new_D759_ & ~new_D769_;
  assign new_D801_ = ~new_D759_ & new_D769_;
  assign new_D802_ = ~new_D758_ | ~new_D783_;
  assign new_D803_ = new_D769_ & new_D802_;
  assign new_D804_ = ~new_D769_ & ~new_D803_;
  assign new_D805_ = new_D769_ | new_D802_;
  assign new_D806_ = ~new_D759_ & new_D760_;
  assign new_D807_ = new_D759_ & ~new_D760_;
  assign new_D808_ = new_D776_ | new_D813_;
  assign new_D809_ = ~new_D776_ & ~new_D812_;
  assign new_D810_ = new_D759_ | new_D776_;
  assign new_D811_ = new_D759_ | new_D760_;
  assign new_D812_ = new_D776_ & new_D813_;
  assign new_D813_ = ~new_D758_ | ~new_D783_;
  assign new_D814_ = new_D791_ & new_D811_;
  assign new_D815_ = ~new_D791_ & ~new_D811_;
  assign new_D816_ = new_D820_ | new_D821_;
  assign new_D817_ = ~new_D762_ & new_D776_;
  assign new_D818_ = new_D822_ | new_D823_;
  assign new_D819_ = new_D762_ & new_D776_;
  assign new_D820_ = ~new_D762_ & ~new_D776_;
  assign new_D821_ = new_D762_ & ~new_D776_;
  assign new_D822_ = new_D762_ & ~new_D776_;
  assign new_D823_ = ~new_D762_ & new_D776_;
  assign new_D824_ = new_E3430_;
  assign new_D825_ = new_E3497_;
  assign new_D826_ = new_E3564_;
  assign new_D827_ = new_E3631_;
  assign new_D828_ = new_E3698_;
  assign new_D829_ = new_E3765_;
  assign new_D830_ = new_D837_ & new_D836_;
  assign new_D831_ = new_D839_ | new_D838_;
  assign new_D832_ = new_D841_ | new_D840_;
  assign new_D833_ = new_D843_ & new_D842_;
  assign new_D834_ = new_D843_ & new_D844_;
  assign new_D835_ = new_D836_ | new_D845_;
  assign new_D836_ = new_D825_ | new_D848_;
  assign new_D837_ = new_D847_ | new_D846_;
  assign new_D838_ = new_D852_ & new_D851_;
  assign new_D839_ = new_D850_ & new_D849_;
  assign new_D840_ = new_D855_ | new_D854_;
  assign new_D841_ = new_D850_ & new_D853_;
  assign new_D842_ = new_D825_ | new_D858_;
  assign new_D843_ = new_D857_ | new_D856_;
  assign new_D844_ = new_D860_ | new_D859_;
  assign new_D845_ = ~new_D836_ & new_D862_;
  assign new_D846_ = ~new_D838_ & new_D850_;
  assign new_D847_ = new_D838_ & ~new_D850_;
  assign new_D848_ = new_D824_ & ~new_D825_;
  assign new_D849_ = ~new_D871_ | ~new_D872_;
  assign new_D850_ = new_D864_ | new_D866_;
  assign new_D851_ = new_D874_ | new_D873_;
  assign new_D852_ = new_D868_ | new_D867_;
  assign new_D853_ = ~new_D876_ | ~new_D875_;
  assign new_D854_ = ~new_D877_ & new_D878_;
  assign new_D855_ = new_D877_ & ~new_D878_;
  assign new_D856_ = ~new_D824_ & new_D825_;
  assign new_D857_ = new_D824_ & ~new_D825_;
  assign new_D858_ = ~new_D840_ | new_D850_;
  assign new_D859_ = new_D840_ & new_D850_;
  assign new_D860_ = ~new_D840_ & ~new_D850_;
  assign new_D861_ = new_D882_ | new_D881_;
  assign new_D862_ = new_D828_ | new_D861_;
  assign new_D863_ = new_D886_ | new_D885_;
  assign new_D864_ = ~new_D828_ & new_D863_;
  assign new_D865_ = new_D884_ | new_D883_;
  assign new_D866_ = new_D828_ & new_D865_;
  assign new_D867_ = new_D826_ & ~new_D836_;
  assign new_D868_ = ~new_D826_ & new_D836_;
  assign new_D869_ = ~new_D825_ | ~new_D850_;
  assign new_D870_ = new_D836_ & new_D869_;
  assign new_D871_ = ~new_D836_ & ~new_D870_;
  assign new_D872_ = new_D836_ | new_D869_;
  assign new_D873_ = ~new_D826_ & new_D827_;
  assign new_D874_ = new_D826_ & ~new_D827_;
  assign new_D875_ = new_D843_ | new_D880_;
  assign new_D876_ = ~new_D843_ & ~new_D879_;
  assign new_D877_ = new_D826_ | new_D843_;
  assign new_D878_ = new_D826_ | new_D827_;
  assign new_D879_ = new_D843_ & new_D880_;
  assign new_D880_ = ~new_D825_ | ~new_D850_;
  assign new_D881_ = new_D858_ & new_D878_;
  assign new_D882_ = ~new_D858_ & ~new_D878_;
  assign new_D883_ = new_D887_ | new_D888_;
  assign new_D884_ = ~new_D829_ & new_D843_;
  assign new_D885_ = new_D889_ | new_D890_;
  assign new_D886_ = new_D829_ & new_D843_;
  assign new_D887_ = ~new_D829_ & ~new_D843_;
  assign new_D888_ = new_D829_ & ~new_D843_;
  assign new_D889_ = new_D829_ & ~new_D843_;
  assign new_D890_ = ~new_D829_ & new_D843_;
  assign new_D891_ = new_E3832_;
  assign new_D892_ = new_E3899_;
  assign new_D893_ = new_E3966_;
  assign new_D894_ = new_E4033_;
  assign new_D895_ = new_E4100_;
  assign new_D896_ = new_E4167_;
  assign new_D897_ = new_D904_ & new_D903_;
  assign new_D898_ = new_D906_ | new_D905_;
  assign new_D899_ = new_D908_ | new_D907_;
  assign new_D900_ = new_D910_ & new_D909_;
  assign new_D901_ = new_D910_ & new_D911_;
  assign new_D902_ = new_D903_ | new_D912_;
  assign new_D903_ = new_D892_ | new_D915_;
  assign new_D904_ = new_D914_ | new_D913_;
  assign new_D905_ = new_D919_ & new_D918_;
  assign new_D906_ = new_D917_ & new_D916_;
  assign new_D907_ = new_D922_ | new_D921_;
  assign new_D908_ = new_D917_ & new_D920_;
  assign new_D909_ = new_D892_ | new_D925_;
  assign new_D910_ = new_D924_ | new_D923_;
  assign new_D911_ = new_D927_ | new_D926_;
  assign new_D912_ = ~new_D903_ & new_D929_;
  assign new_D913_ = ~new_D905_ & new_D917_;
  assign new_D914_ = new_D905_ & ~new_D917_;
  assign new_D915_ = new_D891_ & ~new_D892_;
  assign new_D916_ = ~new_D938_ | ~new_D939_;
  assign new_D917_ = new_D931_ | new_D933_;
  assign new_D918_ = new_D941_ | new_D940_;
  assign new_D919_ = new_D935_ | new_D934_;
  assign new_D920_ = ~new_D943_ | ~new_D942_;
  assign new_D921_ = ~new_D944_ & new_D945_;
  assign new_D922_ = new_D944_ & ~new_D945_;
  assign new_D923_ = ~new_D891_ & new_D892_;
  assign new_D924_ = new_D891_ & ~new_D892_;
  assign new_D925_ = ~new_D907_ | new_D917_;
  assign new_D926_ = new_D907_ & new_D917_;
  assign new_D927_ = ~new_D907_ & ~new_D917_;
  assign new_D928_ = new_D949_ | new_D948_;
  assign new_D929_ = new_D895_ | new_D928_;
  assign new_D930_ = new_D953_ | new_D952_;
  assign new_D931_ = ~new_D895_ & new_D930_;
  assign new_D932_ = new_D951_ | new_D950_;
  assign new_D933_ = new_D895_ & new_D932_;
  assign new_D934_ = new_D893_ & ~new_D903_;
  assign new_D935_ = ~new_D893_ & new_D903_;
  assign new_D936_ = ~new_D892_ | ~new_D917_;
  assign new_D937_ = new_D903_ & new_D936_;
  assign new_D938_ = ~new_D903_ & ~new_D937_;
  assign new_D939_ = new_D903_ | new_D936_;
  assign new_D940_ = ~new_D893_ & new_D894_;
  assign new_D941_ = new_D893_ & ~new_D894_;
  assign new_D942_ = new_D910_ | new_D947_;
  assign new_D943_ = ~new_D910_ & ~new_D946_;
  assign new_D944_ = new_D893_ | new_D910_;
  assign new_D945_ = new_D893_ | new_D894_;
  assign new_D946_ = new_D910_ & new_D947_;
  assign new_D947_ = ~new_D892_ | ~new_D917_;
  assign new_D948_ = new_D925_ & new_D945_;
  assign new_D949_ = ~new_D925_ & ~new_D945_;
  assign new_D950_ = new_D954_ | new_D955_;
  assign new_D951_ = ~new_D896_ & new_D910_;
  assign new_D952_ = new_D956_ | new_D957_;
  assign new_D953_ = new_D896_ & new_D910_;
  assign new_D954_ = ~new_D896_ & ~new_D910_;
  assign new_D955_ = new_D896_ & ~new_D910_;
  assign new_D956_ = new_D896_ & ~new_D910_;
  assign new_D957_ = ~new_D896_ & new_D910_;
  assign new_D958_ = new_E4234_;
  assign new_D959_ = new_E4301_;
  assign new_D960_ = new_E4368_;
  assign new_D961_ = new_E4435_;
  assign new_D962_ = new_E4502_;
  assign new_D963_ = new_E4569_;
  assign new_D964_ = new_D971_ & new_D970_;
  assign new_D965_ = new_D973_ | new_D972_;
  assign new_D966_ = new_D975_ | new_D974_;
  assign new_D967_ = new_D977_ & new_D976_;
  assign new_D968_ = new_D977_ & new_D978_;
  assign new_D969_ = new_D970_ | new_D979_;
  assign new_D970_ = new_D959_ | new_D982_;
  assign new_D971_ = new_D981_ | new_D980_;
  assign new_D972_ = new_D986_ & new_D985_;
  assign new_D973_ = new_D984_ & new_D983_;
  assign new_D974_ = new_D989_ | new_D988_;
  assign new_D975_ = new_D984_ & new_D987_;
  assign new_D976_ = new_D959_ | new_D992_;
  assign new_D977_ = new_D991_ | new_D990_;
  assign new_D978_ = new_D994_ | new_D993_;
  assign new_D979_ = ~new_D970_ & new_D996_;
  assign new_D980_ = ~new_D972_ & new_D984_;
  assign new_D981_ = new_D972_ & ~new_D984_;
  assign new_D982_ = new_D958_ & ~new_D959_;
  assign new_D983_ = ~new_D1005_ | ~new_D1006_;
  assign new_D984_ = new_D998_ | new_D1000_;
  assign new_D985_ = new_D1008_ | new_D1007_;
  assign new_D986_ = new_D1002_ | new_D1001_;
  assign new_D987_ = ~new_D1010_ | ~new_D1009_;
  assign new_D988_ = ~new_D1011_ & new_D1012_;
  assign new_D989_ = new_D1011_ & ~new_D1012_;
  assign new_D990_ = ~new_D958_ & new_D959_;
  assign new_D991_ = new_D958_ & ~new_D959_;
  assign new_D992_ = ~new_D974_ | new_D984_;
  assign new_D993_ = new_D974_ & new_D984_;
  assign new_D994_ = ~new_D974_ & ~new_D984_;
  assign new_D995_ = new_D1016_ | new_D1015_;
  assign new_D996_ = new_D962_ | new_D995_;
  assign new_D997_ = new_D1020_ | new_D1019_;
  assign new_D998_ = ~new_D962_ & new_D997_;
  assign new_D999_ = new_D1018_ | new_D1017_;
  assign new_D1000_ = new_D962_ & new_D999_;
  assign new_D1001_ = new_D960_ & ~new_D970_;
  assign new_D1002_ = ~new_D960_ & new_D970_;
  assign new_D1003_ = ~new_D959_ | ~new_D984_;
  assign new_D1004_ = new_D970_ & new_D1003_;
  assign new_D1005_ = ~new_D970_ & ~new_D1004_;
  assign new_D1006_ = new_D970_ | new_D1003_;
  assign new_D1007_ = ~new_D960_ & new_D961_;
  assign new_D1008_ = new_D960_ & ~new_D961_;
  assign new_D1009_ = new_D977_ | new_D1014_;
  assign new_D1010_ = ~new_D977_ & ~new_D1013_;
  assign new_D1011_ = new_D960_ | new_D977_;
  assign new_D1012_ = new_D960_ | new_D961_;
  assign new_D1013_ = new_D977_ & new_D1014_;
  assign new_D1014_ = ~new_D959_ | ~new_D984_;
  assign new_D1015_ = new_D992_ & new_D1012_;
  assign new_D1016_ = ~new_D992_ & ~new_D1012_;
  assign new_D1017_ = new_D1021_ | new_D1022_;
  assign new_D1018_ = ~new_D963_ & new_D977_;
  assign new_D1019_ = new_D1023_ | new_D1024_;
  assign new_D1020_ = new_D963_ & new_D977_;
  assign new_D1021_ = ~new_D963_ & ~new_D977_;
  assign new_D1022_ = new_D963_ & ~new_D977_;
  assign new_D1023_ = new_D963_ & ~new_D977_;
  assign new_D1024_ = ~new_D963_ & new_D977_;
  assign new_D1025_ = new_E4636_;
  assign new_D1026_ = new_E4703_;
  assign new_D1027_ = new_E4770_;
  assign new_D1028_ = new_E4837_;
  assign new_D1029_ = new_E4904_;
  assign new_D1030_ = new_E4971_;
  assign new_D1031_ = new_D1038_ & new_D1037_;
  assign new_D1032_ = new_D1040_ | new_D1039_;
  assign new_D1033_ = new_D1042_ | new_D1041_;
  assign new_D1034_ = new_D1044_ & new_D1043_;
  assign new_D1035_ = new_D1044_ & new_D1045_;
  assign new_D1036_ = new_D1037_ | new_D1046_;
  assign new_D1037_ = new_D1026_ | new_D1049_;
  assign new_D1038_ = new_D1048_ | new_D1047_;
  assign new_D1039_ = new_D1053_ & new_D1052_;
  assign new_D1040_ = new_D1051_ & new_D1050_;
  assign new_D1041_ = new_D1056_ | new_D1055_;
  assign new_D1042_ = new_D1051_ & new_D1054_;
  assign new_D1043_ = new_D1026_ | new_D1059_;
  assign new_D1044_ = new_D1058_ | new_D1057_;
  assign new_D1045_ = new_D1061_ | new_D1060_;
  assign new_D1046_ = ~new_D1037_ & new_D1063_;
  assign new_D1047_ = ~new_D1039_ & new_D1051_;
  assign new_D1048_ = new_D1039_ & ~new_D1051_;
  assign new_D1049_ = new_D1025_ & ~new_D1026_;
  assign new_D1050_ = ~new_D1072_ | ~new_D1073_;
  assign new_D1051_ = new_D1065_ | new_D1067_;
  assign new_D1052_ = new_D1075_ | new_D1074_;
  assign new_D1053_ = new_D1069_ | new_D1068_;
  assign new_D1054_ = ~new_D1077_ | ~new_D1076_;
  assign new_D1055_ = ~new_D1078_ & new_D1079_;
  assign new_D1056_ = new_D1078_ & ~new_D1079_;
  assign new_D1057_ = ~new_D1025_ & new_D1026_;
  assign new_D1058_ = new_D1025_ & ~new_D1026_;
  assign new_D1059_ = ~new_D1041_ | new_D1051_;
  assign new_D1060_ = new_D1041_ & new_D1051_;
  assign new_D1061_ = ~new_D1041_ & ~new_D1051_;
  assign new_D1062_ = new_D1083_ | new_D1082_;
  assign new_D1063_ = new_D1029_ | new_D1062_;
  assign new_D1064_ = new_D1087_ | new_D1086_;
  assign new_D1065_ = ~new_D1029_ & new_D1064_;
  assign new_D1066_ = new_D1085_ | new_D1084_;
  assign new_D1067_ = new_D1029_ & new_D1066_;
  assign new_D1068_ = new_D1027_ & ~new_D1037_;
  assign new_D1069_ = ~new_D1027_ & new_D1037_;
  assign new_D1070_ = ~new_D1026_ | ~new_D1051_;
  assign new_D1071_ = new_D1037_ & new_D1070_;
  assign new_D1072_ = ~new_D1037_ & ~new_D1071_;
  assign new_D1073_ = new_D1037_ | new_D1070_;
  assign new_D1074_ = ~new_D1027_ & new_D1028_;
  assign new_D1075_ = new_D1027_ & ~new_D1028_;
  assign new_D1076_ = new_D1044_ | new_D1081_;
  assign new_D1077_ = ~new_D1044_ & ~new_D1080_;
  assign new_D1078_ = new_D1027_ | new_D1044_;
  assign new_D1079_ = new_D1027_ | new_D1028_;
  assign new_D1080_ = new_D1044_ & new_D1081_;
  assign new_D1081_ = ~new_D1026_ | ~new_D1051_;
  assign new_D1082_ = new_D1059_ & new_D1079_;
  assign new_D1083_ = ~new_D1059_ & ~new_D1079_;
  assign new_D1084_ = new_D1088_ | new_D1089_;
  assign new_D1085_ = ~new_D1030_ & new_D1044_;
  assign new_D1086_ = new_D1090_ | new_D1091_;
  assign new_D1087_ = new_D1030_ & new_D1044_;
  assign new_D1088_ = ~new_D1030_ & ~new_D1044_;
  assign new_D1089_ = new_D1030_ & ~new_D1044_;
  assign new_D1090_ = new_D1030_ & ~new_D1044_;
  assign new_D1091_ = ~new_D1030_ & new_D1044_;
  assign new_D1092_ = new_E5038_;
  assign new_D1093_ = new_E5105_;
  assign new_D1094_ = new_E5172_;
  assign new_D1095_ = new_E5239_;
  assign new_D1096_ = new_E5306_;
  assign new_D1097_ = new_E5373_;
  assign new_D1098_ = new_D1105_ & new_D1104_;
  assign new_D1099_ = new_D1107_ | new_D1106_;
  assign new_D1100_ = new_D1109_ | new_D1108_;
  assign new_D1101_ = new_D1111_ & new_D1110_;
  assign new_D1102_ = new_D1111_ & new_D1112_;
  assign new_D1103_ = new_D1104_ | new_D1113_;
  assign new_D1104_ = new_D1093_ | new_D1116_;
  assign new_D1105_ = new_D1115_ | new_D1114_;
  assign new_D1106_ = new_D1120_ & new_D1119_;
  assign new_D1107_ = new_D1118_ & new_D1117_;
  assign new_D1108_ = new_D1123_ | new_D1122_;
  assign new_D1109_ = new_D1118_ & new_D1121_;
  assign new_D1110_ = new_D1093_ | new_D1126_;
  assign new_D1111_ = new_D1125_ | new_D1124_;
  assign new_D1112_ = new_D1128_ | new_D1127_;
  assign new_D1113_ = ~new_D1104_ & new_D1130_;
  assign new_D1114_ = ~new_D1106_ & new_D1118_;
  assign new_D1115_ = new_D1106_ & ~new_D1118_;
  assign new_D1116_ = new_D1092_ & ~new_D1093_;
  assign new_D1117_ = ~new_D1139_ | ~new_D1140_;
  assign new_D1118_ = new_D1132_ | new_D1134_;
  assign new_D1119_ = new_D1142_ | new_D1141_;
  assign new_D1120_ = new_D1136_ | new_D1135_;
  assign new_D1121_ = ~new_D1144_ | ~new_D1143_;
  assign new_D1122_ = ~new_D1145_ & new_D1146_;
  assign new_D1123_ = new_D1145_ & ~new_D1146_;
  assign new_D1124_ = ~new_D1092_ & new_D1093_;
  assign new_D1125_ = new_D1092_ & ~new_D1093_;
  assign new_D1126_ = ~new_D1108_ | new_D1118_;
  assign new_D1127_ = new_D1108_ & new_D1118_;
  assign new_D1128_ = ~new_D1108_ & ~new_D1118_;
  assign new_D1129_ = new_D1150_ | new_D1149_;
  assign new_D1130_ = new_D1096_ | new_D1129_;
  assign new_D1131_ = new_D1154_ | new_D1153_;
  assign new_D1132_ = ~new_D1096_ & new_D1131_;
  assign new_D1133_ = new_D1152_ | new_D1151_;
  assign new_D1134_ = new_D1096_ & new_D1133_;
  assign new_D1135_ = new_D1094_ & ~new_D1104_;
  assign new_D1136_ = ~new_D1094_ & new_D1104_;
  assign new_D1137_ = ~new_D1093_ | ~new_D1118_;
  assign new_D1138_ = new_D1104_ & new_D1137_;
  assign new_D1139_ = ~new_D1104_ & ~new_D1138_;
  assign new_D1140_ = new_D1104_ | new_D1137_;
  assign new_D1141_ = ~new_D1094_ & new_D1095_;
  assign new_D1142_ = new_D1094_ & ~new_D1095_;
  assign new_D1143_ = new_D1111_ | new_D1148_;
  assign new_D1144_ = ~new_D1111_ & ~new_D1147_;
  assign new_D1145_ = new_D1094_ | new_D1111_;
  assign new_D1146_ = new_D1094_ | new_D1095_;
  assign new_D1147_ = new_D1111_ & new_D1148_;
  assign new_D1148_ = ~new_D1093_ | ~new_D1118_;
  assign new_D1149_ = new_D1126_ & new_D1146_;
  assign new_D1150_ = ~new_D1126_ & ~new_D1146_;
  assign new_D1151_ = new_D1155_ | new_D1156_;
  assign new_D1152_ = ~new_D1097_ & new_D1111_;
  assign new_D1153_ = new_D1157_ | new_D1158_;
  assign new_D1154_ = new_D1097_ & new_D1111_;
  assign new_D1155_ = ~new_D1097_ & ~new_D1111_;
  assign new_D1156_ = new_D1097_ & ~new_D1111_;
  assign new_D1157_ = new_D1097_ & ~new_D1111_;
  assign new_D1158_ = ~new_D1097_ & new_D1111_;
  assign new_D1159_ = new_E5440_;
  assign new_D1160_ = new_E5507_;
  assign new_D1161_ = new_E5574_;
  assign new_D1162_ = new_E5641_;
  assign new_D1163_ = new_E5708_;
  assign new_D1164_ = new_E5775_;
  assign new_D1165_ = new_D1172_ & new_D1171_;
  assign new_D1166_ = new_D1174_ | new_D1173_;
  assign new_D1167_ = new_D1176_ | new_D1175_;
  assign new_D1168_ = new_D1178_ & new_D1177_;
  assign new_D1169_ = new_D1178_ & new_D1179_;
  assign new_D1170_ = new_D1171_ | new_D1180_;
  assign new_D1171_ = new_D1160_ | new_D1183_;
  assign new_D1172_ = new_D1182_ | new_D1181_;
  assign new_D1173_ = new_D1187_ & new_D1186_;
  assign new_D1174_ = new_D1185_ & new_D1184_;
  assign new_D1175_ = new_D1190_ | new_D1189_;
  assign new_D1176_ = new_D1185_ & new_D1188_;
  assign new_D1177_ = new_D1160_ | new_D1193_;
  assign new_D1178_ = new_D1192_ | new_D1191_;
  assign new_D1179_ = new_D1195_ | new_D1194_;
  assign new_D1180_ = ~new_D1171_ & new_D1197_;
  assign new_D1181_ = ~new_D1173_ & new_D1185_;
  assign new_D1182_ = new_D1173_ & ~new_D1185_;
  assign new_D1183_ = new_D1159_ & ~new_D1160_;
  assign new_D1184_ = ~new_D1206_ | ~new_D1207_;
  assign new_D1185_ = new_D1199_ | new_D1201_;
  assign new_D1186_ = new_D1209_ | new_D1208_;
  assign new_D1187_ = new_D1203_ | new_D1202_;
  assign new_D1188_ = ~new_D1211_ | ~new_D1210_;
  assign new_D1189_ = ~new_D1212_ & new_D1213_;
  assign new_D1190_ = new_D1212_ & ~new_D1213_;
  assign new_D1191_ = ~new_D1159_ & new_D1160_;
  assign new_D1192_ = new_D1159_ & ~new_D1160_;
  assign new_D1193_ = ~new_D1175_ | new_D1185_;
  assign new_D1194_ = new_D1175_ & new_D1185_;
  assign new_D1195_ = ~new_D1175_ & ~new_D1185_;
  assign new_D1196_ = new_D1217_ | new_D1216_;
  assign new_D1197_ = new_D1163_ | new_D1196_;
  assign new_D1198_ = new_D1221_ | new_D1220_;
  assign new_D1199_ = ~new_D1163_ & new_D1198_;
  assign new_D1200_ = new_D1219_ | new_D1218_;
  assign new_D1201_ = new_D1163_ & new_D1200_;
  assign new_D1202_ = new_D1161_ & ~new_D1171_;
  assign new_D1203_ = ~new_D1161_ & new_D1171_;
  assign new_D1204_ = ~new_D1160_ | ~new_D1185_;
  assign new_D1205_ = new_D1171_ & new_D1204_;
  assign new_D1206_ = ~new_D1171_ & ~new_D1205_;
  assign new_D1207_ = new_D1171_ | new_D1204_;
  assign new_D1208_ = ~new_D1161_ & new_D1162_;
  assign new_D1209_ = new_D1161_ & ~new_D1162_;
  assign new_D1210_ = new_D1178_ | new_D1215_;
  assign new_D1211_ = ~new_D1178_ & ~new_D1214_;
  assign new_D1212_ = new_D1161_ | new_D1178_;
  assign new_D1213_ = new_D1161_ | new_D1162_;
  assign new_D1214_ = new_D1178_ & new_D1215_;
  assign new_D1215_ = ~new_D1160_ | ~new_D1185_;
  assign new_D1216_ = new_D1193_ & new_D1213_;
  assign new_D1217_ = ~new_D1193_ & ~new_D1213_;
  assign new_D1218_ = new_D1222_ | new_D1223_;
  assign new_D1219_ = ~new_D1164_ & new_D1178_;
  assign new_D1220_ = new_D1224_ | new_D1225_;
  assign new_D1221_ = new_D1164_ & new_D1178_;
  assign new_D1222_ = ~new_D1164_ & ~new_D1178_;
  assign new_D1223_ = new_D1164_ & ~new_D1178_;
  assign new_D1224_ = new_D1164_ & ~new_D1178_;
  assign new_D1225_ = ~new_D1164_ & new_D1178_;
  assign new_D1226_ = new_E5842_;
  assign new_D1227_ = new_E5909_;
  assign new_D1228_ = new_E5976_;
  assign new_D1229_ = new_E6043_;
  assign new_D1230_ = new_E6110_;
  assign new_D1231_ = new_E6177_;
  assign new_D1232_ = new_D1239_ & new_D1238_;
  assign new_D1233_ = new_D1241_ | new_D1240_;
  assign new_D1234_ = new_D1243_ | new_D1242_;
  assign new_D1235_ = new_D1245_ & new_D1244_;
  assign new_D1236_ = new_D1245_ & new_D1246_;
  assign new_D1237_ = new_D1238_ | new_D1247_;
  assign new_D1238_ = new_D1227_ | new_D1250_;
  assign new_D1239_ = new_D1249_ | new_D1248_;
  assign new_D1240_ = new_D1254_ & new_D1253_;
  assign new_D1241_ = new_D1252_ & new_D1251_;
  assign new_D1242_ = new_D1257_ | new_D1256_;
  assign new_D1243_ = new_D1252_ & new_D1255_;
  assign new_D1244_ = new_D1227_ | new_D1260_;
  assign new_D1245_ = new_D1259_ | new_D1258_;
  assign new_D1246_ = new_D1262_ | new_D1261_;
  assign new_D1247_ = ~new_D1238_ & new_D1264_;
  assign new_D1248_ = ~new_D1240_ & new_D1252_;
  assign new_D1249_ = new_D1240_ & ~new_D1252_;
  assign new_D1250_ = new_D1226_ & ~new_D1227_;
  assign new_D1251_ = ~new_D1273_ | ~new_D1274_;
  assign new_D1252_ = new_D1266_ | new_D1268_;
  assign new_D1253_ = new_D1276_ | new_D1275_;
  assign new_D1254_ = new_D1270_ | new_D1269_;
  assign new_D1255_ = ~new_D1278_ | ~new_D1277_;
  assign new_D1256_ = ~new_D1279_ & new_D1280_;
  assign new_D1257_ = new_D1279_ & ~new_D1280_;
  assign new_D1258_ = ~new_D1226_ & new_D1227_;
  assign new_D1259_ = new_D1226_ & ~new_D1227_;
  assign new_D1260_ = ~new_D1242_ | new_D1252_;
  assign new_D1261_ = new_D1242_ & new_D1252_;
  assign new_D1262_ = ~new_D1242_ & ~new_D1252_;
  assign new_D1263_ = new_D1284_ | new_D1283_;
  assign new_D1264_ = new_D1230_ | new_D1263_;
  assign new_D1265_ = new_D1288_ | new_D1287_;
  assign new_D1266_ = ~new_D1230_ & new_D1265_;
  assign new_D1267_ = new_D1286_ | new_D1285_;
  assign new_D1268_ = new_D1230_ & new_D1267_;
  assign new_D1269_ = new_D1228_ & ~new_D1238_;
  assign new_D1270_ = ~new_D1228_ & new_D1238_;
  assign new_D1271_ = ~new_D1227_ | ~new_D1252_;
  assign new_D1272_ = new_D1238_ & new_D1271_;
  assign new_D1273_ = ~new_D1238_ & ~new_D1272_;
  assign new_D1274_ = new_D1238_ | new_D1271_;
  assign new_D1275_ = ~new_D1228_ & new_D1229_;
  assign new_D1276_ = new_D1228_ & ~new_D1229_;
  assign new_D1277_ = new_D1245_ | new_D1282_;
  assign new_D1278_ = ~new_D1245_ & ~new_D1281_;
  assign new_D1279_ = new_D1228_ | new_D1245_;
  assign new_D1280_ = new_D1228_ | new_D1229_;
  assign new_D1281_ = new_D1245_ & new_D1282_;
  assign new_D1282_ = ~new_D1227_ | ~new_D1252_;
  assign new_D1283_ = new_D1260_ & new_D1280_;
  assign new_D1284_ = ~new_D1260_ & ~new_D1280_;
  assign new_D1285_ = new_D1289_ | new_D1290_;
  assign new_D1286_ = ~new_D1231_ & new_D1245_;
  assign new_D1287_ = new_D1291_ | new_D1292_;
  assign new_D1288_ = new_D1231_ & new_D1245_;
  assign new_D1289_ = ~new_D1231_ & ~new_D1245_;
  assign new_D1290_ = new_D1231_ & ~new_D1245_;
  assign new_D1291_ = new_D1231_ & ~new_D1245_;
  assign new_D1292_ = ~new_D1231_ & new_D1245_;
  assign new_D1293_ = new_E6244_;
  assign new_D1294_ = new_E6311_;
  assign new_D1295_ = new_E6378_;
  assign new_D1296_ = new_E6445_;
  assign new_D1297_ = new_E6512_;
  assign new_D1298_ = new_E6579_;
  assign new_D1299_ = new_D1306_ & new_D1305_;
  assign new_D1300_ = new_D1308_ | new_D1307_;
  assign new_D1301_ = new_D1310_ | new_D1309_;
  assign new_D1302_ = new_D1312_ & new_D1311_;
  assign new_D1303_ = new_D1312_ & new_D1313_;
  assign new_D1304_ = new_D1305_ | new_D1314_;
  assign new_D1305_ = new_D1294_ | new_D1317_;
  assign new_D1306_ = new_D1316_ | new_D1315_;
  assign new_D1307_ = new_D1321_ & new_D1320_;
  assign new_D1308_ = new_D1319_ & new_D1318_;
  assign new_D1309_ = new_D1324_ | new_D1323_;
  assign new_D1310_ = new_D1319_ & new_D1322_;
  assign new_D1311_ = new_D1294_ | new_D1327_;
  assign new_D1312_ = new_D1326_ | new_D1325_;
  assign new_D1313_ = new_D1329_ | new_D1328_;
  assign new_D1314_ = ~new_D1305_ & new_D1331_;
  assign new_D1315_ = ~new_D1307_ & new_D1319_;
  assign new_D1316_ = new_D1307_ & ~new_D1319_;
  assign new_D1317_ = new_D1293_ & ~new_D1294_;
  assign new_D1318_ = ~new_D1340_ | ~new_D1341_;
  assign new_D1319_ = new_D1333_ | new_D1335_;
  assign new_D1320_ = new_D1343_ | new_D1342_;
  assign new_D1321_ = new_D1337_ | new_D1336_;
  assign new_D1322_ = ~new_D1345_ | ~new_D1344_;
  assign new_D1323_ = ~new_D1346_ & new_D1347_;
  assign new_D1324_ = new_D1346_ & ~new_D1347_;
  assign new_D1325_ = ~new_D1293_ & new_D1294_;
  assign new_D1326_ = new_D1293_ & ~new_D1294_;
  assign new_D1327_ = ~new_D1309_ | new_D1319_;
  assign new_D1328_ = new_D1309_ & new_D1319_;
  assign new_D1329_ = ~new_D1309_ & ~new_D1319_;
  assign new_D1330_ = new_D1351_ | new_D1350_;
  assign new_D1331_ = new_D1297_ | new_D1330_;
  assign new_D1332_ = new_D1355_ | new_D1354_;
  assign new_D1333_ = ~new_D1297_ & new_D1332_;
  assign new_D1334_ = new_D1353_ | new_D1352_;
  assign new_D1335_ = new_D1297_ & new_D1334_;
  assign new_D1336_ = new_D1295_ & ~new_D1305_;
  assign new_D1337_ = ~new_D1295_ & new_D1305_;
  assign new_D1338_ = ~new_D1294_ | ~new_D1319_;
  assign new_D1339_ = new_D1305_ & new_D1338_;
  assign new_D1340_ = ~new_D1305_ & ~new_D1339_;
  assign new_D1341_ = new_D1305_ | new_D1338_;
  assign new_D1342_ = ~new_D1295_ & new_D1296_;
  assign new_D1343_ = new_D1295_ & ~new_D1296_;
  assign new_D1344_ = new_D1312_ | new_D1349_;
  assign new_D1345_ = ~new_D1312_ & ~new_D1348_;
  assign new_D1346_ = new_D1295_ | new_D1312_;
  assign new_D1347_ = new_D1295_ | new_D1296_;
  assign new_D1348_ = new_D1312_ & new_D1349_;
  assign new_D1349_ = ~new_D1294_ | ~new_D1319_;
  assign new_D1350_ = new_D1327_ & new_D1347_;
  assign new_D1351_ = ~new_D1327_ & ~new_D1347_;
  assign new_D1352_ = new_D1356_ | new_D1357_;
  assign new_D1353_ = ~new_D1298_ & new_D1312_;
  assign new_D1354_ = new_D1358_ | new_D1359_;
  assign new_D1355_ = new_D1298_ & new_D1312_;
  assign new_D1356_ = ~new_D1298_ & ~new_D1312_;
  assign new_D1357_ = new_D1298_ & ~new_D1312_;
  assign new_D1358_ = new_D1298_ & ~new_D1312_;
  assign new_D1359_ = ~new_D1298_ & new_D1312_;
  assign new_D1360_ = new_E6646_;
  assign new_D1361_ = new_E6713_;
  assign new_D1362_ = new_E6780_;
  assign new_D1363_ = new_E6847_;
  assign new_D1364_ = new_E6914_;
  assign new_D1365_ = new_E6981_;
  assign new_D1366_ = new_D1373_ & new_D1372_;
  assign new_D1367_ = new_D1375_ | new_D1374_;
  assign new_D1368_ = new_D1377_ | new_D1376_;
  assign new_D1369_ = new_D1379_ & new_D1378_;
  assign new_D1370_ = new_D1379_ & new_D1380_;
  assign new_D1371_ = new_D1372_ | new_D1381_;
  assign new_D1372_ = new_D1361_ | new_D1384_;
  assign new_D1373_ = new_D1383_ | new_D1382_;
  assign new_D1374_ = new_D1388_ & new_D1387_;
  assign new_D1375_ = new_D1386_ & new_D1385_;
  assign new_D1376_ = new_D1391_ | new_D1390_;
  assign new_D1377_ = new_D1386_ & new_D1389_;
  assign new_D1378_ = new_D1361_ | new_D1394_;
  assign new_D1379_ = new_D1393_ | new_D1392_;
  assign new_D1380_ = new_D1396_ | new_D1395_;
  assign new_D1381_ = ~new_D1372_ & new_D1398_;
  assign new_D1382_ = ~new_D1374_ & new_D1386_;
  assign new_D1383_ = new_D1374_ & ~new_D1386_;
  assign new_D1384_ = new_D1360_ & ~new_D1361_;
  assign new_D1385_ = ~new_D1407_ | ~new_D1408_;
  assign new_D1386_ = new_D1400_ | new_D1402_;
  assign new_D1387_ = new_D1410_ | new_D1409_;
  assign new_D1388_ = new_D1404_ | new_D1403_;
  assign new_D1389_ = ~new_D1412_ | ~new_D1411_;
  assign new_D1390_ = ~new_D1413_ & new_D1414_;
  assign new_D1391_ = new_D1413_ & ~new_D1414_;
  assign new_D1392_ = ~new_D1360_ & new_D1361_;
  assign new_D1393_ = new_D1360_ & ~new_D1361_;
  assign new_D1394_ = ~new_D1376_ | new_D1386_;
  assign new_D1395_ = new_D1376_ & new_D1386_;
  assign new_D1396_ = ~new_D1376_ & ~new_D1386_;
  assign new_D1397_ = new_D1418_ | new_D1417_;
  assign new_D1398_ = new_D1364_ | new_D1397_;
  assign new_D1399_ = new_D1422_ | new_D1421_;
  assign new_D1400_ = ~new_D1364_ & new_D1399_;
  assign new_D1401_ = new_D1420_ | new_D1419_;
  assign new_D1402_ = new_D1364_ & new_D1401_;
  assign new_D1403_ = new_D1362_ & ~new_D1372_;
  assign new_D1404_ = ~new_D1362_ & new_D1372_;
  assign new_D1405_ = ~new_D1361_ | ~new_D1386_;
  assign new_D1406_ = new_D1372_ & new_D1405_;
  assign new_D1407_ = ~new_D1372_ & ~new_D1406_;
  assign new_D1408_ = new_D1372_ | new_D1405_;
  assign new_D1409_ = ~new_D1362_ & new_D1363_;
  assign new_D1410_ = new_D1362_ & ~new_D1363_;
  assign new_D1411_ = new_D1379_ | new_D1416_;
  assign new_D1412_ = ~new_D1379_ & ~new_D1415_;
  assign new_D1413_ = new_D1362_ | new_D1379_;
  assign new_D1414_ = new_D1362_ | new_D1363_;
  assign new_D1415_ = new_D1379_ & new_D1416_;
  assign new_D1416_ = ~new_D1361_ | ~new_D1386_;
  assign new_D1417_ = new_D1394_ & new_D1414_;
  assign new_D1418_ = ~new_D1394_ & ~new_D1414_;
  assign new_D1419_ = new_D1423_ | new_D1424_;
  assign new_D1420_ = ~new_D1365_ & new_D1379_;
  assign new_D1421_ = new_D1425_ | new_D1426_;
  assign new_D1422_ = new_D1365_ & new_D1379_;
  assign new_D1423_ = ~new_D1365_ & ~new_D1379_;
  assign new_D1424_ = new_D1365_ & ~new_D1379_;
  assign new_D1425_ = new_D1365_ & ~new_D1379_;
  assign new_D1426_ = ~new_D1365_ & new_D1379_;
  assign new_D1427_ = new_E7048_;
  assign new_D1428_ = new_E7115_;
  assign new_D1429_ = new_E7182_;
  assign new_D1430_ = new_E7249_;
  assign new_D1431_ = new_E7316_;
  assign new_D1432_ = new_E7383_;
  assign new_D1433_ = new_D1440_ & new_D1439_;
  assign new_D1434_ = new_D1442_ | new_D1441_;
  assign new_D1435_ = new_D1444_ | new_D1443_;
  assign new_D1436_ = new_D1446_ & new_D1445_;
  assign new_D1437_ = new_D1446_ & new_D1447_;
  assign new_D1438_ = new_D1439_ | new_D1448_;
  assign new_D1439_ = new_D1428_ | new_D1451_;
  assign new_D1440_ = new_D1450_ | new_D1449_;
  assign new_D1441_ = new_D1455_ & new_D1454_;
  assign new_D1442_ = new_D1453_ & new_D1452_;
  assign new_D1443_ = new_D1458_ | new_D1457_;
  assign new_D1444_ = new_D1453_ & new_D1456_;
  assign new_D1445_ = new_D1428_ | new_D1461_;
  assign new_D1446_ = new_D1460_ | new_D1459_;
  assign new_D1447_ = new_D1463_ | new_D1462_;
  assign new_D1448_ = ~new_D1439_ & new_D1465_;
  assign new_D1449_ = ~new_D1441_ & new_D1453_;
  assign new_D1450_ = new_D1441_ & ~new_D1453_;
  assign new_D1451_ = new_D1427_ & ~new_D1428_;
  assign new_D1452_ = ~new_D1474_ | ~new_D1475_;
  assign new_D1453_ = new_D1467_ | new_D1469_;
  assign new_D1454_ = new_D1477_ | new_D1476_;
  assign new_D1455_ = new_D1471_ | new_D1470_;
  assign new_D1456_ = ~new_D1479_ | ~new_D1478_;
  assign new_D1457_ = ~new_D1480_ & new_D1481_;
  assign new_D1458_ = new_D1480_ & ~new_D1481_;
  assign new_D1459_ = ~new_D1427_ & new_D1428_;
  assign new_D1460_ = new_D1427_ & ~new_D1428_;
  assign new_D1461_ = ~new_D1443_ | new_D1453_;
  assign new_D1462_ = new_D1443_ & new_D1453_;
  assign new_D1463_ = ~new_D1443_ & ~new_D1453_;
  assign new_D1464_ = new_D1485_ | new_D1484_;
  assign new_D1465_ = new_D1431_ | new_D1464_;
  assign new_D1466_ = new_D1489_ | new_D1488_;
  assign new_D1467_ = ~new_D1431_ & new_D1466_;
  assign new_D1468_ = new_D1487_ | new_D1486_;
  assign new_D1469_ = new_D1431_ & new_D1468_;
  assign new_D1470_ = new_D1429_ & ~new_D1439_;
  assign new_D1471_ = ~new_D1429_ & new_D1439_;
  assign new_D1472_ = ~new_D1428_ | ~new_D1453_;
  assign new_D1473_ = new_D1439_ & new_D1472_;
  assign new_D1474_ = ~new_D1439_ & ~new_D1473_;
  assign new_D1475_ = new_D1439_ | new_D1472_;
  assign new_D1476_ = ~new_D1429_ & new_D1430_;
  assign new_D1477_ = new_D1429_ & ~new_D1430_;
  assign new_D1478_ = new_D1446_ | new_D1483_;
  assign new_D1479_ = ~new_D1446_ & ~new_D1482_;
  assign new_D1480_ = new_D1429_ | new_D1446_;
  assign new_D1481_ = new_D1429_ | new_D1430_;
  assign new_D1482_ = new_D1446_ & new_D1483_;
  assign new_D1483_ = ~new_D1428_ | ~new_D1453_;
  assign new_D1484_ = new_D1461_ & new_D1481_;
  assign new_D1485_ = ~new_D1461_ & ~new_D1481_;
  assign new_D1486_ = new_D1490_ | new_D1491_;
  assign new_D1487_ = ~new_D1432_ & new_D1446_;
  assign new_D1488_ = new_D1492_ | new_D1493_;
  assign new_D1489_ = new_D1432_ & new_D1446_;
  assign new_D1490_ = ~new_D1432_ & ~new_D1446_;
  assign new_D1491_ = new_D1432_ & ~new_D1446_;
  assign new_D1492_ = new_D1432_ & ~new_D1446_;
  assign new_D1493_ = ~new_D1432_ & new_D1446_;
  assign new_D1494_ = new_E7450_;
  assign new_D1495_ = new_E7517_;
  assign new_D1496_ = new_E7584_;
  assign new_D1497_ = new_E7651_;
  assign new_D1498_ = new_E7718_;
  assign new_D1499_ = new_E7785_;
  assign new_D1500_ = new_D1507_ & new_D1506_;
  assign new_D1501_ = new_D1509_ | new_D1508_;
  assign new_D1502_ = new_D1511_ | new_D1510_;
  assign new_D1503_ = new_D1513_ & new_D1512_;
  assign new_D1504_ = new_D1513_ & new_D1514_;
  assign new_D1505_ = new_D1506_ | new_D1515_;
  assign new_D1506_ = new_D1495_ | new_D1518_;
  assign new_D1507_ = new_D1517_ | new_D1516_;
  assign new_D1508_ = new_D1522_ & new_D1521_;
  assign new_D1509_ = new_D1520_ & new_D1519_;
  assign new_D1510_ = new_D1525_ | new_D1524_;
  assign new_D1511_ = new_D1520_ & new_D1523_;
  assign new_D1512_ = new_D1495_ | new_D1528_;
  assign new_D1513_ = new_D1527_ | new_D1526_;
  assign new_D1514_ = new_D1530_ | new_D1529_;
  assign new_D1515_ = ~new_D1506_ & new_D1532_;
  assign new_D1516_ = ~new_D1508_ & new_D1520_;
  assign new_D1517_ = new_D1508_ & ~new_D1520_;
  assign new_D1518_ = new_D1494_ & ~new_D1495_;
  assign new_D1519_ = ~new_D1541_ | ~new_D1542_;
  assign new_D1520_ = new_D1534_ | new_D1536_;
  assign new_D1521_ = new_D1544_ | new_D1543_;
  assign new_D1522_ = new_D1538_ | new_D1537_;
  assign new_D1523_ = ~new_D1546_ | ~new_D1545_;
  assign new_D1524_ = ~new_D1547_ & new_D1548_;
  assign new_D1525_ = new_D1547_ & ~new_D1548_;
  assign new_D1526_ = ~new_D1494_ & new_D1495_;
  assign new_D1527_ = new_D1494_ & ~new_D1495_;
  assign new_D1528_ = ~new_D1510_ | new_D1520_;
  assign new_D1529_ = new_D1510_ & new_D1520_;
  assign new_D1530_ = ~new_D1510_ & ~new_D1520_;
  assign new_D1531_ = new_D1552_ | new_D1551_;
  assign new_D1532_ = new_D1498_ | new_D1531_;
  assign new_D1533_ = new_D1556_ | new_D1555_;
  assign new_D1534_ = ~new_D1498_ & new_D1533_;
  assign new_D1535_ = new_D1554_ | new_D1553_;
  assign new_D1536_ = new_D1498_ & new_D1535_;
  assign new_D1537_ = new_D1496_ & ~new_D1506_;
  assign new_D1538_ = ~new_D1496_ & new_D1506_;
  assign new_D1539_ = ~new_D1495_ | ~new_D1520_;
  assign new_D1540_ = new_D1506_ & new_D1539_;
  assign new_D1541_ = ~new_D1506_ & ~new_D1540_;
  assign new_D1542_ = new_D1506_ | new_D1539_;
  assign new_D1543_ = ~new_D1496_ & new_D1497_;
  assign new_D1544_ = new_D1496_ & ~new_D1497_;
  assign new_D1545_ = new_D1513_ | new_D1550_;
  assign new_D1546_ = ~new_D1513_ & ~new_D1549_;
  assign new_D1547_ = new_D1496_ | new_D1513_;
  assign new_D1548_ = new_D1496_ | new_D1497_;
  assign new_D1549_ = new_D1513_ & new_D1550_;
  assign new_D1550_ = ~new_D1495_ | ~new_D1520_;
  assign new_D1551_ = new_D1528_ & new_D1548_;
  assign new_D1552_ = ~new_D1528_ & ~new_D1548_;
  assign new_D1553_ = new_D1557_ | new_D1558_;
  assign new_D1554_ = ~new_D1499_ & new_D1513_;
  assign new_D1555_ = new_D1559_ | new_D1560_;
  assign new_D1556_ = new_D1499_ & new_D1513_;
  assign new_D1557_ = ~new_D1499_ & ~new_D1513_;
  assign new_D1558_ = new_D1499_ & ~new_D1513_;
  assign new_D1559_ = new_D1499_ & ~new_D1513_;
  assign new_D1560_ = ~new_D1499_ & new_D1513_;
  assign new_D1561_ = new_E7852_;
  assign new_D1562_ = new_E7919_;
  assign new_D1563_ = new_E7986_;
  assign new_D1564_ = new_E8053_;
  assign new_D1565_ = new_E8120_;
  assign new_D1566_ = new_E8187_;
  assign new_D1567_ = new_D1574_ & new_D1573_;
  assign new_D1568_ = new_D1576_ | new_D1575_;
  assign new_D1569_ = new_D1578_ | new_D1577_;
  assign new_D1570_ = new_D1580_ & new_D1579_;
  assign new_D1571_ = new_D1580_ & new_D1581_;
  assign new_D1572_ = new_D1573_ | new_D1582_;
  assign new_D1573_ = new_D1562_ | new_D1585_;
  assign new_D1574_ = new_D1584_ | new_D1583_;
  assign new_D1575_ = new_D1589_ & new_D1588_;
  assign new_D1576_ = new_D1587_ & new_D1586_;
  assign new_D1577_ = new_D1592_ | new_D1591_;
  assign new_D1578_ = new_D1587_ & new_D1590_;
  assign new_D1579_ = new_D1562_ | new_D1595_;
  assign new_D1580_ = new_D1594_ | new_D1593_;
  assign new_D1581_ = new_D1597_ | new_D1596_;
  assign new_D1582_ = ~new_D1573_ & new_D1599_;
  assign new_D1583_ = ~new_D1575_ & new_D1587_;
  assign new_D1584_ = new_D1575_ & ~new_D1587_;
  assign new_D1585_ = new_D1561_ & ~new_D1562_;
  assign new_D1586_ = ~new_D1608_ | ~new_D1609_;
  assign new_D1587_ = new_D1601_ | new_D1603_;
  assign new_D1588_ = new_D1611_ | new_D1610_;
  assign new_D1589_ = new_D1605_ | new_D1604_;
  assign new_D1590_ = ~new_D1613_ | ~new_D1612_;
  assign new_D1591_ = ~new_D1614_ & new_D1615_;
  assign new_D1592_ = new_D1614_ & ~new_D1615_;
  assign new_D1593_ = ~new_D1561_ & new_D1562_;
  assign new_D1594_ = new_D1561_ & ~new_D1562_;
  assign new_D1595_ = ~new_D1577_ | new_D1587_;
  assign new_D1596_ = new_D1577_ & new_D1587_;
  assign new_D1597_ = ~new_D1577_ & ~new_D1587_;
  assign new_D1598_ = new_D1619_ | new_D1618_;
  assign new_D1599_ = new_D1565_ | new_D1598_;
  assign new_D1600_ = new_D1623_ | new_D1622_;
  assign new_D1601_ = ~new_D1565_ & new_D1600_;
  assign new_D1602_ = new_D1621_ | new_D1620_;
  assign new_D1603_ = new_D1565_ & new_D1602_;
  assign new_D1604_ = new_D1563_ & ~new_D1573_;
  assign new_D1605_ = ~new_D1563_ & new_D1573_;
  assign new_D1606_ = ~new_D1562_ | ~new_D1587_;
  assign new_D1607_ = new_D1573_ & new_D1606_;
  assign new_D1608_ = ~new_D1573_ & ~new_D1607_;
  assign new_D1609_ = new_D1573_ | new_D1606_;
  assign new_D1610_ = ~new_D1563_ & new_D1564_;
  assign new_D1611_ = new_D1563_ & ~new_D1564_;
  assign new_D1612_ = new_D1580_ | new_D1617_;
  assign new_D1613_ = ~new_D1580_ & ~new_D1616_;
  assign new_D1614_ = new_D1563_ | new_D1580_;
  assign new_D1615_ = new_D1563_ | new_D1564_;
  assign new_D1616_ = new_D1580_ & new_D1617_;
  assign new_D1617_ = ~new_D1562_ | ~new_D1587_;
  assign new_D1618_ = new_D1595_ & new_D1615_;
  assign new_D1619_ = ~new_D1595_ & ~new_D1615_;
  assign new_D1620_ = new_D1624_ | new_D1625_;
  assign new_D1621_ = ~new_D1566_ & new_D1580_;
  assign new_D1622_ = new_D1626_ | new_D1627_;
  assign new_D1623_ = new_D1566_ & new_D1580_;
  assign new_D1624_ = ~new_D1566_ & ~new_D1580_;
  assign new_D1625_ = new_D1566_ & ~new_D1580_;
  assign new_D1626_ = new_D1566_ & ~new_D1580_;
  assign new_D1627_ = ~new_D1566_ & new_D1580_;
  assign new_D1628_ = new_E8254_;
  assign new_D1629_ = new_E8321_;
  assign new_D1630_ = new_E8388_;
  assign new_D1631_ = new_E8455_;
  assign new_D1632_ = new_E8522_;
  assign new_D1633_ = new_E8589_;
  assign new_D1634_ = new_D1641_ & new_D1640_;
  assign new_D1635_ = new_D1643_ | new_D1642_;
  assign new_D1636_ = new_D1645_ | new_D1644_;
  assign new_D1637_ = new_D1647_ & new_D1646_;
  assign new_D1638_ = new_D1647_ & new_D1648_;
  assign new_D1639_ = new_D1640_ | new_D1649_;
  assign new_D1640_ = new_D1629_ | new_D1652_;
  assign new_D1641_ = new_D1651_ | new_D1650_;
  assign new_D1642_ = new_D1656_ & new_D1655_;
  assign new_D1643_ = new_D1654_ & new_D1653_;
  assign new_D1644_ = new_D1659_ | new_D1658_;
  assign new_D1645_ = new_D1654_ & new_D1657_;
  assign new_D1646_ = new_D1629_ | new_D1662_;
  assign new_D1647_ = new_D1661_ | new_D1660_;
  assign new_D1648_ = new_D1664_ | new_D1663_;
  assign new_D1649_ = ~new_D1640_ & new_D1666_;
  assign new_D1650_ = ~new_D1642_ & new_D1654_;
  assign new_D1651_ = new_D1642_ & ~new_D1654_;
  assign new_D1652_ = new_D1628_ & ~new_D1629_;
  assign new_D1653_ = ~new_D1675_ | ~new_D1676_;
  assign new_D1654_ = new_D1668_ | new_D1670_;
  assign new_D1655_ = new_D1678_ | new_D1677_;
  assign new_D1656_ = new_D1672_ | new_D1671_;
  assign new_D1657_ = ~new_D1680_ | ~new_D1679_;
  assign new_D1658_ = ~new_D1681_ & new_D1682_;
  assign new_D1659_ = new_D1681_ & ~new_D1682_;
  assign new_D1660_ = ~new_D1628_ & new_D1629_;
  assign new_D1661_ = new_D1628_ & ~new_D1629_;
  assign new_D1662_ = ~new_D1644_ | new_D1654_;
  assign new_D1663_ = new_D1644_ & new_D1654_;
  assign new_D1664_ = ~new_D1644_ & ~new_D1654_;
  assign new_D1665_ = new_D1686_ | new_D1685_;
  assign new_D1666_ = new_D1632_ | new_D1665_;
  assign new_D1667_ = new_D1690_ | new_D1689_;
  assign new_D1668_ = ~new_D1632_ & new_D1667_;
  assign new_D1669_ = new_D1688_ | new_D1687_;
  assign new_D1670_ = new_D1632_ & new_D1669_;
  assign new_D1671_ = new_D1630_ & ~new_D1640_;
  assign new_D1672_ = ~new_D1630_ & new_D1640_;
  assign new_D1673_ = ~new_D1629_ | ~new_D1654_;
  assign new_D1674_ = new_D1640_ & new_D1673_;
  assign new_D1675_ = ~new_D1640_ & ~new_D1674_;
  assign new_D1676_ = new_D1640_ | new_D1673_;
  assign new_D1677_ = ~new_D1630_ & new_D1631_;
  assign new_D1678_ = new_D1630_ & ~new_D1631_;
  assign new_D1679_ = new_D1647_ | new_D1684_;
  assign new_D1680_ = ~new_D1647_ & ~new_D1683_;
  assign new_D1681_ = new_D1630_ | new_D1647_;
  assign new_D1682_ = new_D1630_ | new_D1631_;
  assign new_D1683_ = new_D1647_ & new_D1684_;
  assign new_D1684_ = ~new_D1629_ | ~new_D1654_;
  assign new_D1685_ = new_D1662_ & new_D1682_;
  assign new_D1686_ = ~new_D1662_ & ~new_D1682_;
  assign new_D1687_ = new_D1691_ | new_D1692_;
  assign new_D1688_ = ~new_D1633_ & new_D1647_;
  assign new_D1689_ = new_D1693_ | new_D1694_;
  assign new_D1690_ = new_D1633_ & new_D1647_;
  assign new_D1691_ = ~new_D1633_ & ~new_D1647_;
  assign new_D1692_ = new_D1633_ & ~new_D1647_;
  assign new_D1693_ = new_D1633_ & ~new_D1647_;
  assign new_D1694_ = ~new_D1633_ & new_D1647_;
  assign new_D1695_ = new_E8656_;
  assign new_D1696_ = new_E8723_;
  assign new_D1697_ = new_E8790_;
  assign new_D1698_ = new_E8857_;
  assign new_D1699_ = new_E8924_;
  assign new_D1700_ = new_E8991_;
  assign new_D1701_ = new_D1708_ & new_D1707_;
  assign new_D1702_ = new_D1710_ | new_D1709_;
  assign new_D1703_ = new_D1712_ | new_D1711_;
  assign new_D1704_ = new_D1714_ & new_D1713_;
  assign new_D1705_ = new_D1714_ & new_D1715_;
  assign new_D1706_ = new_D1707_ | new_D1716_;
  assign new_D1707_ = new_D1696_ | new_D1719_;
  assign new_D1708_ = new_D1718_ | new_D1717_;
  assign new_D1709_ = new_D1723_ & new_D1722_;
  assign new_D1710_ = new_D1721_ & new_D1720_;
  assign new_D1711_ = new_D1726_ | new_D1725_;
  assign new_D1712_ = new_D1721_ & new_D1724_;
  assign new_D1713_ = new_D1696_ | new_D1729_;
  assign new_D1714_ = new_D1728_ | new_D1727_;
  assign new_D1715_ = new_D1731_ | new_D1730_;
  assign new_D1716_ = ~new_D1707_ & new_D1733_;
  assign new_D1717_ = ~new_D1709_ & new_D1721_;
  assign new_D1718_ = new_D1709_ & ~new_D1721_;
  assign new_D1719_ = new_D1695_ & ~new_D1696_;
  assign new_D1720_ = ~new_D1742_ | ~new_D1743_;
  assign new_D1721_ = new_D1735_ | new_D1737_;
  assign new_D1722_ = new_D1745_ | new_D1744_;
  assign new_D1723_ = new_D1739_ | new_D1738_;
  assign new_D1724_ = ~new_D1747_ | ~new_D1746_;
  assign new_D1725_ = ~new_D1748_ & new_D1749_;
  assign new_D1726_ = new_D1748_ & ~new_D1749_;
  assign new_D1727_ = ~new_D1695_ & new_D1696_;
  assign new_D1728_ = new_D1695_ & ~new_D1696_;
  assign new_D1729_ = ~new_D1711_ | new_D1721_;
  assign new_D1730_ = new_D1711_ & new_D1721_;
  assign new_D1731_ = ~new_D1711_ & ~new_D1721_;
  assign new_D1732_ = new_D1753_ | new_D1752_;
  assign new_D1733_ = new_D1699_ | new_D1732_;
  assign new_D1734_ = new_D1757_ | new_D1756_;
  assign new_D1735_ = ~new_D1699_ & new_D1734_;
  assign new_D1736_ = new_D1755_ | new_D1754_;
  assign new_D1737_ = new_D1699_ & new_D1736_;
  assign new_D1738_ = new_D1697_ & ~new_D1707_;
  assign new_D1739_ = ~new_D1697_ & new_D1707_;
  assign new_D1740_ = ~new_D1696_ | ~new_D1721_;
  assign new_D1741_ = new_D1707_ & new_D1740_;
  assign new_D1742_ = ~new_D1707_ & ~new_D1741_;
  assign new_D1743_ = new_D1707_ | new_D1740_;
  assign new_D1744_ = ~new_D1697_ & new_D1698_;
  assign new_D1745_ = new_D1697_ & ~new_D1698_;
  assign new_D1746_ = new_D1714_ | new_D1751_;
  assign new_D1747_ = ~new_D1714_ & ~new_D1750_;
  assign new_D1748_ = new_D1697_ | new_D1714_;
  assign new_D1749_ = new_D1697_ | new_D1698_;
  assign new_D1750_ = new_D1714_ & new_D1751_;
  assign new_D1751_ = ~new_D1696_ | ~new_D1721_;
  assign new_D1752_ = new_D1729_ & new_D1749_;
  assign new_D1753_ = ~new_D1729_ & ~new_D1749_;
  assign new_D1754_ = new_D1758_ | new_D1759_;
  assign new_D1755_ = ~new_D1700_ & new_D1714_;
  assign new_D1756_ = new_D1760_ | new_D1761_;
  assign new_D1757_ = new_D1700_ & new_D1714_;
  assign new_D1758_ = ~new_D1700_ & ~new_D1714_;
  assign new_D1759_ = new_D1700_ & ~new_D1714_;
  assign new_D1760_ = new_D1700_ & ~new_D1714_;
  assign new_D1761_ = ~new_D1700_ & new_D1714_;
  assign new_D1762_ = new_E9058_;
  assign new_D1763_ = new_E9125_;
  assign new_D1764_ = new_E9192_;
  assign new_D1765_ = new_E9259_;
  assign new_D1766_ = new_E9326_;
  assign new_D1767_ = new_E9393_;
  assign new_D1768_ = new_D1775_ & new_D1774_;
  assign new_D1769_ = new_D1777_ | new_D1776_;
  assign new_D1770_ = new_D1779_ | new_D1778_;
  assign new_D1771_ = new_D1781_ & new_D1780_;
  assign new_D1772_ = new_D1781_ & new_D1782_;
  assign new_D1773_ = new_D1774_ | new_D1783_;
  assign new_D1774_ = new_D1763_ | new_D1786_;
  assign new_D1775_ = new_D1785_ | new_D1784_;
  assign new_D1776_ = new_D1790_ & new_D1789_;
  assign new_D1777_ = new_D1788_ & new_D1787_;
  assign new_D1778_ = new_D1793_ | new_D1792_;
  assign new_D1779_ = new_D1788_ & new_D1791_;
  assign new_D1780_ = new_D1763_ | new_D1796_;
  assign new_D1781_ = new_D1795_ | new_D1794_;
  assign new_D1782_ = new_D1798_ | new_D1797_;
  assign new_D1783_ = ~new_D1774_ & new_D1800_;
  assign new_D1784_ = ~new_D1776_ & new_D1788_;
  assign new_D1785_ = new_D1776_ & ~new_D1788_;
  assign new_D1786_ = new_D1762_ & ~new_D1763_;
  assign new_D1787_ = ~new_D1809_ | ~new_D1810_;
  assign new_D1788_ = new_D1802_ | new_D1804_;
  assign new_D1789_ = new_D1812_ | new_D1811_;
  assign new_D1790_ = new_D1806_ | new_D1805_;
  assign new_D1791_ = ~new_D1814_ | ~new_D1813_;
  assign new_D1792_ = ~new_D1815_ & new_D1816_;
  assign new_D1793_ = new_D1815_ & ~new_D1816_;
  assign new_D1794_ = ~new_D1762_ & new_D1763_;
  assign new_D1795_ = new_D1762_ & ~new_D1763_;
  assign new_D1796_ = ~new_D1778_ | new_D1788_;
  assign new_D1797_ = new_D1778_ & new_D1788_;
  assign new_D1798_ = ~new_D1778_ & ~new_D1788_;
  assign new_D1799_ = new_D1820_ | new_D1819_;
  assign new_D1800_ = new_D1766_ | new_D1799_;
  assign new_D1801_ = new_D1824_ | new_D1823_;
  assign new_D1802_ = ~new_D1766_ & new_D1801_;
  assign new_D1803_ = new_D1822_ | new_D1821_;
  assign new_D1804_ = new_D1766_ & new_D1803_;
  assign new_D1805_ = new_D1764_ & ~new_D1774_;
  assign new_D1806_ = ~new_D1764_ & new_D1774_;
  assign new_D1807_ = ~new_D1763_ | ~new_D1788_;
  assign new_D1808_ = new_D1774_ & new_D1807_;
  assign new_D1809_ = ~new_D1774_ & ~new_D1808_;
  assign new_D1810_ = new_D1774_ | new_D1807_;
  assign new_D1811_ = ~new_D1764_ & new_D1765_;
  assign new_D1812_ = new_D1764_ & ~new_D1765_;
  assign new_D1813_ = new_D1781_ | new_D1818_;
  assign new_D1814_ = ~new_D1781_ & ~new_D1817_;
  assign new_D1815_ = new_D1764_ | new_D1781_;
  assign new_D1816_ = new_D1764_ | new_D1765_;
  assign new_D1817_ = new_D1781_ & new_D1818_;
  assign new_D1818_ = ~new_D1763_ | ~new_D1788_;
  assign new_D1819_ = new_D1796_ & new_D1816_;
  assign new_D1820_ = ~new_D1796_ & ~new_D1816_;
  assign new_D1821_ = new_D1825_ | new_D1826_;
  assign new_D1822_ = ~new_D1767_ & new_D1781_;
  assign new_D1823_ = new_D1827_ | new_D1828_;
  assign new_D1824_ = new_D1767_ & new_D1781_;
  assign new_D1825_ = ~new_D1767_ & ~new_D1781_;
  assign new_D1826_ = new_D1767_ & ~new_D1781_;
  assign new_D1827_ = new_D1767_ & ~new_D1781_;
  assign new_D1828_ = ~new_D1767_ & new_D1781_;
  assign new_D1829_ = new_E9460_;
  assign new_D1830_ = new_E9527_;
  assign new_D1831_ = new_E9594_;
  assign new_D1832_ = new_E9661_;
  assign new_D1833_ = new_E9728_;
  assign new_D1834_ = new_E9795_;
  assign new_D1835_ = new_D1842_ & new_D1841_;
  assign new_D1836_ = new_D1844_ | new_D1843_;
  assign new_D1837_ = new_D1846_ | new_D1845_;
  assign new_D1838_ = new_D1848_ & new_D1847_;
  assign new_D1839_ = new_D1848_ & new_D1849_;
  assign new_D1840_ = new_D1841_ | new_D1850_;
  assign new_D1841_ = new_D1830_ | new_D1853_;
  assign new_D1842_ = new_D1852_ | new_D1851_;
  assign new_D1843_ = new_D1857_ & new_D1856_;
  assign new_D1844_ = new_D1855_ & new_D1854_;
  assign new_D1845_ = new_D1860_ | new_D1859_;
  assign new_D1846_ = new_D1855_ & new_D1858_;
  assign new_D1847_ = new_D1830_ | new_D1863_;
  assign new_D1848_ = new_D1862_ | new_D1861_;
  assign new_D1849_ = new_D1865_ | new_D1864_;
  assign new_D1850_ = ~new_D1841_ & new_D1867_;
  assign new_D1851_ = ~new_D1843_ & new_D1855_;
  assign new_D1852_ = new_D1843_ & ~new_D1855_;
  assign new_D1853_ = new_D1829_ & ~new_D1830_;
  assign new_D1854_ = ~new_D1876_ | ~new_D1877_;
  assign new_D1855_ = new_D1869_ | new_D1871_;
  assign new_D1856_ = new_D1879_ | new_D1878_;
  assign new_D1857_ = new_D1873_ | new_D1872_;
  assign new_D1858_ = ~new_D1881_ | ~new_D1880_;
  assign new_D1859_ = ~new_D1882_ & new_D1883_;
  assign new_D1860_ = new_D1882_ & ~new_D1883_;
  assign new_D1861_ = ~new_D1829_ & new_D1830_;
  assign new_D1862_ = new_D1829_ & ~new_D1830_;
  assign new_D1863_ = ~new_D1845_ | new_D1855_;
  assign new_D1864_ = new_D1845_ & new_D1855_;
  assign new_D1865_ = ~new_D1845_ & ~new_D1855_;
  assign new_D1866_ = new_D1887_ | new_D1886_;
  assign new_D1867_ = new_D1833_ | new_D1866_;
  assign new_D1868_ = new_D1891_ | new_D1890_;
  assign new_D1869_ = ~new_D1833_ & new_D1868_;
  assign new_D1870_ = new_D1889_ | new_D1888_;
  assign new_D1871_ = new_D1833_ & new_D1870_;
  assign new_D1872_ = new_D1831_ & ~new_D1841_;
  assign new_D1873_ = ~new_D1831_ & new_D1841_;
  assign new_D1874_ = ~new_D1830_ | ~new_D1855_;
  assign new_D1875_ = new_D1841_ & new_D1874_;
  assign new_D1876_ = ~new_D1841_ & ~new_D1875_;
  assign new_D1877_ = new_D1841_ | new_D1874_;
  assign new_D1878_ = ~new_D1831_ & new_D1832_;
  assign new_D1879_ = new_D1831_ & ~new_D1832_;
  assign new_D1880_ = new_D1848_ | new_D1885_;
  assign new_D1881_ = ~new_D1848_ & ~new_D1884_;
  assign new_D1882_ = new_D1831_ | new_D1848_;
  assign new_D1883_ = new_D1831_ | new_D1832_;
  assign new_D1884_ = new_D1848_ & new_D1885_;
  assign new_D1885_ = ~new_D1830_ | ~new_D1855_;
  assign new_D1886_ = new_D1863_ & new_D1883_;
  assign new_D1887_ = ~new_D1863_ & ~new_D1883_;
  assign new_D1888_ = new_D1892_ | new_D1893_;
  assign new_D1889_ = ~new_D1834_ & new_D1848_;
  assign new_D1890_ = new_D1894_ | new_D1895_;
  assign new_D1891_ = new_D1834_ & new_D1848_;
  assign new_D1892_ = ~new_D1834_ & ~new_D1848_;
  assign new_D1893_ = new_D1834_ & ~new_D1848_;
  assign new_D1894_ = new_D1834_ & ~new_D1848_;
  assign new_D1895_ = ~new_D1834_ & new_D1848_;
  assign new_D1896_ = new_E9862_;
  assign new_D1897_ = new_E9929_;
  assign new_D1898_ = new_E9996_;
  assign new_D1899_ = new_F64_;
  assign new_D1900_ = new_F131_;
  assign new_D1901_ = new_F198_;
  assign new_D1902_ = new_D1909_ & new_D1908_;
  assign new_D1903_ = new_D1911_ | new_D1910_;
  assign new_D1904_ = new_D1913_ | new_D1912_;
  assign new_D1905_ = new_D1915_ & new_D1914_;
  assign new_D1906_ = new_D1915_ & new_D1916_;
  assign new_D1907_ = new_D1908_ | new_D1917_;
  assign new_D1908_ = new_D1897_ | new_D1920_;
  assign new_D1909_ = new_D1919_ | new_D1918_;
  assign new_D1910_ = new_D1924_ & new_D1923_;
  assign new_D1911_ = new_D1922_ & new_D1921_;
  assign new_D1912_ = new_D1927_ | new_D1926_;
  assign new_D1913_ = new_D1922_ & new_D1925_;
  assign new_D1914_ = new_D1897_ | new_D1930_;
  assign new_D1915_ = new_D1929_ | new_D1928_;
  assign new_D1916_ = new_D1932_ | new_D1931_;
  assign new_D1917_ = ~new_D1908_ & new_D1934_;
  assign new_D1918_ = ~new_D1910_ & new_D1922_;
  assign new_D1919_ = new_D1910_ & ~new_D1922_;
  assign new_D1920_ = new_D1896_ & ~new_D1897_;
  assign new_D1921_ = ~new_D1943_ | ~new_D1944_;
  assign new_D1922_ = new_D1936_ | new_D1938_;
  assign new_D1923_ = new_D1946_ | new_D1945_;
  assign new_D1924_ = new_D1940_ | new_D1939_;
  assign new_D1925_ = ~new_D1948_ | ~new_D1947_;
  assign new_D1926_ = ~new_D1949_ & new_D1950_;
  assign new_D1927_ = new_D1949_ & ~new_D1950_;
  assign new_D1928_ = ~new_D1896_ & new_D1897_;
  assign new_D1929_ = new_D1896_ & ~new_D1897_;
  assign new_D1930_ = ~new_D1912_ | new_D1922_;
  assign new_D1931_ = new_D1912_ & new_D1922_;
  assign new_D1932_ = ~new_D1912_ & ~new_D1922_;
  assign new_D1933_ = new_D1954_ | new_D1953_;
  assign new_D1934_ = new_D1900_ | new_D1933_;
  assign new_D1935_ = new_D1958_ | new_D1957_;
  assign new_D1936_ = ~new_D1900_ & new_D1935_;
  assign new_D1937_ = new_D1956_ | new_D1955_;
  assign new_D1938_ = new_D1900_ & new_D1937_;
  assign new_D1939_ = new_D1898_ & ~new_D1908_;
  assign new_D1940_ = ~new_D1898_ & new_D1908_;
  assign new_D1941_ = ~new_D1897_ | ~new_D1922_;
  assign new_D1942_ = new_D1908_ & new_D1941_;
  assign new_D1943_ = ~new_D1908_ & ~new_D1942_;
  assign new_D1944_ = new_D1908_ | new_D1941_;
  assign new_D1945_ = ~new_D1898_ & new_D1899_;
  assign new_D1946_ = new_D1898_ & ~new_D1899_;
  assign new_D1947_ = new_D1915_ | new_D1952_;
  assign new_D1948_ = ~new_D1915_ & ~new_D1951_;
  assign new_D1949_ = new_D1898_ | new_D1915_;
  assign new_D1950_ = new_D1898_ | new_D1899_;
  assign new_D1951_ = new_D1915_ & new_D1952_;
  assign new_D1952_ = ~new_D1897_ | ~new_D1922_;
  assign new_D1953_ = new_D1930_ & new_D1950_;
  assign new_D1954_ = ~new_D1930_ & ~new_D1950_;
  assign new_D1955_ = new_D1959_ | new_D1960_;
  assign new_D1956_ = ~new_D1901_ & new_D1915_;
  assign new_D1957_ = new_D1961_ | new_D1962_;
  assign new_D1958_ = new_D1901_ & new_D1915_;
  assign new_D1959_ = ~new_D1901_ & ~new_D1915_;
  assign new_D1960_ = new_D1901_ & ~new_D1915_;
  assign new_D1961_ = new_D1901_ & ~new_D1915_;
  assign new_D1962_ = ~new_D1901_ & new_D1915_;
  assign new_D1963_ = new_F265_;
  assign new_D1964_ = new_F332_;
  assign new_D1965_ = new_F399_;
  assign new_D1966_ = new_F466_;
  assign new_D1967_ = new_F533_;
  assign new_D1968_ = new_F600_;
  assign new_D1969_ = new_D1976_ & new_D1975_;
  assign new_D1970_ = new_D1978_ | new_D1977_;
  assign new_D1971_ = new_D1980_ | new_D1979_;
  assign new_D1972_ = new_D1982_ & new_D1981_;
  assign new_D1973_ = new_D1982_ & new_D1983_;
  assign new_D1974_ = new_D1975_ | new_D1984_;
  assign new_D1975_ = new_D1964_ | new_D1987_;
  assign new_D1976_ = new_D1986_ | new_D1985_;
  assign new_D1977_ = new_D1991_ & new_D1990_;
  assign new_D1978_ = new_D1989_ & new_D1988_;
  assign new_D1979_ = new_D1994_ | new_D1993_;
  assign new_D1980_ = new_D1989_ & new_D1992_;
  assign new_D1981_ = new_D1964_ | new_D1997_;
  assign new_D1982_ = new_D1996_ | new_D1995_;
  assign new_D1983_ = new_D1999_ | new_D1998_;
  assign new_D1984_ = ~new_D1975_ & new_D2001_;
  assign new_D1985_ = ~new_D1977_ & new_D1989_;
  assign new_D1986_ = new_D1977_ & ~new_D1989_;
  assign new_D1987_ = new_D1963_ & ~new_D1964_;
  assign new_D1988_ = ~new_D2010_ | ~new_D2011_;
  assign new_D1989_ = new_D2003_ | new_D2005_;
  assign new_D1990_ = new_D2013_ | new_D2012_;
  assign new_D1991_ = new_D2007_ | new_D2006_;
  assign new_D1992_ = ~new_D2015_ | ~new_D2014_;
  assign new_D1993_ = ~new_D2016_ & new_D2017_;
  assign new_D1994_ = new_D2016_ & ~new_D2017_;
  assign new_D1995_ = ~new_D1963_ & new_D1964_;
  assign new_D1996_ = new_D1963_ & ~new_D1964_;
  assign new_D1997_ = ~new_D1979_ | new_D1989_;
  assign new_D1998_ = new_D1979_ & new_D1989_;
  assign new_D1999_ = ~new_D1979_ & ~new_D1989_;
  assign new_D2000_ = new_D2021_ | new_D2020_;
  assign new_D2001_ = new_D1967_ | new_D2000_;
  assign new_D2002_ = new_D2025_ | new_D2024_;
  assign new_D2003_ = ~new_D1967_ & new_D2002_;
  assign new_D2004_ = new_D2023_ | new_D2022_;
  assign new_D2005_ = new_D1967_ & new_D2004_;
  assign new_D2006_ = new_D1965_ & ~new_D1975_;
  assign new_D2007_ = ~new_D1965_ & new_D1975_;
  assign new_D2008_ = ~new_D1964_ | ~new_D1989_;
  assign new_D2009_ = new_D1975_ & new_D2008_;
  assign new_D2010_ = ~new_D1975_ & ~new_D2009_;
  assign new_D2011_ = new_D1975_ | new_D2008_;
  assign new_D2012_ = ~new_D1965_ & new_D1966_;
  assign new_D2013_ = new_D1965_ & ~new_D1966_;
  assign new_D2014_ = new_D1982_ | new_D2019_;
  assign new_D2015_ = ~new_D1982_ & ~new_D2018_;
  assign new_D2016_ = new_D1965_ | new_D1982_;
  assign new_D2017_ = new_D1965_ | new_D1966_;
  assign new_D2018_ = new_D1982_ & new_D2019_;
  assign new_D2019_ = ~new_D1964_ | ~new_D1989_;
  assign new_D2020_ = new_D1997_ & new_D2017_;
  assign new_D2021_ = ~new_D1997_ & ~new_D2017_;
  assign new_D2022_ = new_D2026_ | new_D2027_;
  assign new_D2023_ = ~new_D1968_ & new_D1982_;
  assign new_D2024_ = new_D2028_ | new_D2029_;
  assign new_D2025_ = new_D1968_ & new_D1982_;
  assign new_D2026_ = ~new_D1968_ & ~new_D1982_;
  assign new_D2027_ = new_D1968_ & ~new_D1982_;
  assign new_D2028_ = new_D1968_ & ~new_D1982_;
  assign new_D2029_ = ~new_D1968_ & new_D1982_;
  assign new_D2030_ = new_F667_;
  assign new_D2031_ = new_F734_;
  assign new_D2032_ = new_F801_;
  assign new_D2033_ = new_F868_;
  assign new_D2034_ = new_F935_;
  assign new_D2035_ = new_F1002_;
  assign new_D2036_ = new_D2043_ & new_D2042_;
  assign new_D2037_ = new_D2045_ | new_D2044_;
  assign new_D2038_ = new_D2047_ | new_D2046_;
  assign new_D2039_ = new_D2049_ & new_D2048_;
  assign new_D2040_ = new_D2049_ & new_D2050_;
  assign new_D2041_ = new_D2042_ | new_D2051_;
  assign new_D2042_ = new_D2031_ | new_D2054_;
  assign new_D2043_ = new_D2053_ | new_D2052_;
  assign new_D2044_ = new_D2058_ & new_D2057_;
  assign new_D2045_ = new_D2056_ & new_D2055_;
  assign new_D2046_ = new_D2061_ | new_D2060_;
  assign new_D2047_ = new_D2056_ & new_D2059_;
  assign new_D2048_ = new_D2031_ | new_D2064_;
  assign new_D2049_ = new_D2063_ | new_D2062_;
  assign new_D2050_ = new_D2066_ | new_D2065_;
  assign new_D2051_ = ~new_D2042_ & new_D2068_;
  assign new_D2052_ = ~new_D2044_ & new_D2056_;
  assign new_D2053_ = new_D2044_ & ~new_D2056_;
  assign new_D2054_ = new_D2030_ & ~new_D2031_;
  assign new_D2055_ = ~new_D2077_ | ~new_D2078_;
  assign new_D2056_ = new_D2070_ | new_D2072_;
  assign new_D2057_ = new_D2080_ | new_D2079_;
  assign new_D2058_ = new_D2074_ | new_D2073_;
  assign new_D2059_ = ~new_D2082_ | ~new_D2081_;
  assign new_D2060_ = ~new_D2083_ & new_D2084_;
  assign new_D2061_ = new_D2083_ & ~new_D2084_;
  assign new_D2062_ = ~new_D2030_ & new_D2031_;
  assign new_D2063_ = new_D2030_ & ~new_D2031_;
  assign new_D2064_ = ~new_D2046_ | new_D2056_;
  assign new_D2065_ = new_D2046_ & new_D2056_;
  assign new_D2066_ = ~new_D2046_ & ~new_D2056_;
  assign new_D2067_ = new_D2088_ | new_D2087_;
  assign new_D2068_ = new_D2034_ | new_D2067_;
  assign new_D2069_ = new_D2092_ | new_D2091_;
  assign new_D2070_ = ~new_D2034_ & new_D2069_;
  assign new_D2071_ = new_D2090_ | new_D2089_;
  assign new_D2072_ = new_D2034_ & new_D2071_;
  assign new_D2073_ = new_D2032_ & ~new_D2042_;
  assign new_D2074_ = ~new_D2032_ & new_D2042_;
  assign new_D2075_ = ~new_D2031_ | ~new_D2056_;
  assign new_D2076_ = new_D2042_ & new_D2075_;
  assign new_D2077_ = ~new_D2042_ & ~new_D2076_;
  assign new_D2078_ = new_D2042_ | new_D2075_;
  assign new_D2079_ = ~new_D2032_ & new_D2033_;
  assign new_D2080_ = new_D2032_ & ~new_D2033_;
  assign new_D2081_ = new_D2049_ | new_D2086_;
  assign new_D2082_ = ~new_D2049_ & ~new_D2085_;
  assign new_D2083_ = new_D2032_ | new_D2049_;
  assign new_D2084_ = new_D2032_ | new_D2033_;
  assign new_D2085_ = new_D2049_ & new_D2086_;
  assign new_D2086_ = ~new_D2031_ | ~new_D2056_;
  assign new_D2087_ = new_D2064_ & new_D2084_;
  assign new_D2088_ = ~new_D2064_ & ~new_D2084_;
  assign new_D2089_ = new_D2093_ | new_D2094_;
  assign new_D2090_ = ~new_D2035_ & new_D2049_;
  assign new_D2091_ = new_D2095_ | new_D2096_;
  assign new_D2092_ = new_D2035_ & new_D2049_;
  assign new_D2093_ = ~new_D2035_ & ~new_D2049_;
  assign new_D2094_ = new_D2035_ & ~new_D2049_;
  assign new_D2095_ = new_D2035_ & ~new_D2049_;
  assign new_D2096_ = ~new_D2035_ & new_D2049_;
  assign new_D2097_ = new_F1069_;
  assign new_D2098_ = new_F1136_;
  assign new_D2099_ = new_F1203_;
  assign new_D2100_ = new_F1270_;
  assign new_D2101_ = new_F1337_;
  assign new_D2102_ = new_F1404_;
  assign new_D2103_ = new_D2110_ & new_D2109_;
  assign new_D2104_ = new_D2112_ | new_D2111_;
  assign new_D2105_ = new_D2114_ | new_D2113_;
  assign new_D2106_ = new_D2116_ & new_D2115_;
  assign new_D2107_ = new_D2116_ & new_D2117_;
  assign new_D2108_ = new_D2109_ | new_D2118_;
  assign new_D2109_ = new_D2098_ | new_D2121_;
  assign new_D2110_ = new_D2120_ | new_D2119_;
  assign new_D2111_ = new_D2125_ & new_D2124_;
  assign new_D2112_ = new_D2123_ & new_D2122_;
  assign new_D2113_ = new_D2128_ | new_D2127_;
  assign new_D2114_ = new_D2123_ & new_D2126_;
  assign new_D2115_ = new_D2098_ | new_D2131_;
  assign new_D2116_ = new_D2130_ | new_D2129_;
  assign new_D2117_ = new_D2133_ | new_D2132_;
  assign new_D2118_ = ~new_D2109_ & new_D2135_;
  assign new_D2119_ = ~new_D2111_ & new_D2123_;
  assign new_D2120_ = new_D2111_ & ~new_D2123_;
  assign new_D2121_ = new_D2097_ & ~new_D2098_;
  assign new_D2122_ = ~new_D2144_ | ~new_D2145_;
  assign new_D2123_ = new_D2137_ | new_D2139_;
  assign new_D2124_ = new_D2147_ | new_D2146_;
  assign new_D2125_ = new_D2141_ | new_D2140_;
  assign new_D2126_ = ~new_D2149_ | ~new_D2148_;
  assign new_D2127_ = ~new_D2150_ & new_D2151_;
  assign new_D2128_ = new_D2150_ & ~new_D2151_;
  assign new_D2129_ = ~new_D2097_ & new_D2098_;
  assign new_D2130_ = new_D2097_ & ~new_D2098_;
  assign new_D2131_ = ~new_D2113_ | new_D2123_;
  assign new_D2132_ = new_D2113_ & new_D2123_;
  assign new_D2133_ = ~new_D2113_ & ~new_D2123_;
  assign new_D2134_ = new_D2155_ | new_D2154_;
  assign new_D2135_ = new_D2101_ | new_D2134_;
  assign new_D2136_ = new_D2159_ | new_D2158_;
  assign new_D2137_ = ~new_D2101_ & new_D2136_;
  assign new_D2138_ = new_D2157_ | new_D2156_;
  assign new_D2139_ = new_D2101_ & new_D2138_;
  assign new_D2140_ = new_D2099_ & ~new_D2109_;
  assign new_D2141_ = ~new_D2099_ & new_D2109_;
  assign new_D2142_ = ~new_D2098_ | ~new_D2123_;
  assign new_D2143_ = new_D2109_ & new_D2142_;
  assign new_D2144_ = ~new_D2109_ & ~new_D2143_;
  assign new_D2145_ = new_D2109_ | new_D2142_;
  assign new_D2146_ = ~new_D2099_ & new_D2100_;
  assign new_D2147_ = new_D2099_ & ~new_D2100_;
  assign new_D2148_ = new_D2116_ | new_D2153_;
  assign new_D2149_ = ~new_D2116_ & ~new_D2152_;
  assign new_D2150_ = new_D2099_ | new_D2116_;
  assign new_D2151_ = new_D2099_ | new_D2100_;
  assign new_D2152_ = new_D2116_ & new_D2153_;
  assign new_D2153_ = ~new_D2098_ | ~new_D2123_;
  assign new_D2154_ = new_D2131_ & new_D2151_;
  assign new_D2155_ = ~new_D2131_ & ~new_D2151_;
  assign new_D2156_ = new_D2160_ | new_D2161_;
  assign new_D2157_ = ~new_D2102_ & new_D2116_;
  assign new_D2158_ = new_D2162_ | new_D2163_;
  assign new_D2159_ = new_D2102_ & new_D2116_;
  assign new_D2160_ = ~new_D2102_ & ~new_D2116_;
  assign new_D2161_ = new_D2102_ & ~new_D2116_;
  assign new_D2162_ = new_D2102_ & ~new_D2116_;
  assign new_D2163_ = ~new_D2102_ & new_D2116_;
  assign new_D2164_ = new_D6995_;
  assign new_D2165_ = new_D7065_;
  assign new_D2166_ = new_D7132_;
  assign new_D2167_ = new_D7199_;
  assign new_D2168_ = new_D7266_;
  assign new_D2169_ = new_D7333_;
  assign new_D2170_ = new_D2177_ & new_D2176_;
  assign new_D2171_ = new_D2179_ | new_D2178_;
  assign new_D2172_ = new_D2181_ | new_D2180_;
  assign new_D2173_ = new_D2183_ & new_D2182_;
  assign new_D2174_ = new_D2183_ & new_D2184_;
  assign new_D2175_ = new_D2176_ | new_D2185_;
  assign new_D2176_ = new_D2165_ | new_D2188_;
  assign new_D2177_ = new_D2187_ | new_D2186_;
  assign new_D2178_ = new_D2192_ & new_D2191_;
  assign new_D2179_ = new_D2190_ & new_D2189_;
  assign new_D2180_ = new_D2195_ | new_D2194_;
  assign new_D2181_ = new_D2190_ & new_D2193_;
  assign new_D2182_ = new_D2165_ | new_D2198_;
  assign new_D2183_ = new_D2197_ | new_D2196_;
  assign new_D2184_ = new_D2200_ | new_D2199_;
  assign new_D2185_ = ~new_D2176_ & new_D2202_;
  assign new_D2186_ = ~new_D2178_ & new_D2190_;
  assign new_D2187_ = new_D2178_ & ~new_D2190_;
  assign new_D2188_ = new_D2164_ & ~new_D2165_;
  assign new_D2189_ = ~new_D2211_ | ~new_D2212_;
  assign new_D2190_ = new_D2204_ | new_D2206_;
  assign new_D2191_ = new_D2214_ | new_D2213_;
  assign new_D2192_ = new_D2208_ | new_D2207_;
  assign new_D2193_ = ~new_D2216_ | ~new_D2215_;
  assign new_D2194_ = ~new_D2217_ & new_D2218_;
  assign new_D2195_ = new_D2217_ & ~new_D2218_;
  assign new_D2196_ = ~new_D2164_ & new_D2165_;
  assign new_D2197_ = new_D2164_ & ~new_D2165_;
  assign new_D2198_ = ~new_D2180_ | new_D2190_;
  assign new_D2199_ = new_D2180_ & new_D2190_;
  assign new_D2200_ = ~new_D2180_ & ~new_D2190_;
  assign new_D2201_ = new_D2222_ | new_D2221_;
  assign new_D2202_ = new_D2168_ | new_D2201_;
  assign new_D2203_ = new_D2226_ | new_D2225_;
  assign new_D2204_ = ~new_D2168_ & new_D2203_;
  assign new_D2205_ = new_D2224_ | new_D2223_;
  assign new_D2206_ = new_D2168_ & new_D2205_;
  assign new_D2207_ = new_D2166_ & ~new_D2176_;
  assign new_D2208_ = ~new_D2166_ & new_D2176_;
  assign new_D2209_ = ~new_D2165_ | ~new_D2190_;
  assign new_D2210_ = new_D2176_ & new_D2209_;
  assign new_D2211_ = ~new_D2176_ & ~new_D2210_;
  assign new_D2212_ = new_D2176_ | new_D2209_;
  assign new_D2213_ = ~new_D2166_ & new_D2167_;
  assign new_D2214_ = new_D2166_ & ~new_D2167_;
  assign new_D2215_ = new_D2183_ | new_D2220_;
  assign new_D2216_ = ~new_D2183_ & ~new_D2219_;
  assign new_D2217_ = new_D2166_ | new_D2183_;
  assign new_D2218_ = new_D2166_ | new_D2167_;
  assign new_D2219_ = new_D2183_ & new_D2220_;
  assign new_D2220_ = ~new_D2165_ | ~new_D2190_;
  assign new_D2221_ = new_D2198_ & new_D2218_;
  assign new_D2222_ = ~new_D2198_ & ~new_D2218_;
  assign new_D2223_ = new_D2227_ | new_D2228_;
  assign new_D2224_ = ~new_D2169_ & new_D2183_;
  assign new_D2225_ = new_D2229_ | new_D2230_;
  assign new_D2226_ = new_D2169_ & new_D2183_;
  assign new_D2227_ = ~new_D2169_ & ~new_D2183_;
  assign new_D2228_ = new_D2169_ & ~new_D2183_;
  assign new_D2229_ = new_D2169_ & ~new_D2183_;
  assign new_D2230_ = ~new_D2169_ & new_D2183_;
  assign new_D2231_ = new_D7400_;
  assign new_D2232_ = new_D7467_;
  assign new_D2233_ = new_D7534_;
  assign new_D2234_ = new_D7601_;
  assign new_D2235_ = new_D7668_;
  assign new_D2236_ = new_D7735_;
  assign new_D2237_ = new_D2244_ & new_D2243_;
  assign new_D2238_ = new_D2246_ | new_D2245_;
  assign new_D2239_ = new_D2248_ | new_D2247_;
  assign new_D2240_ = new_D2250_ & new_D2249_;
  assign new_D2241_ = new_D2250_ & new_D2251_;
  assign new_D2242_ = new_D2243_ | new_D2252_;
  assign new_D2243_ = new_D2232_ | new_D2255_;
  assign new_D2244_ = new_D2254_ | new_D2253_;
  assign new_D2245_ = new_D2259_ & new_D2258_;
  assign new_D2246_ = new_D2257_ & new_D2256_;
  assign new_D2247_ = new_D2262_ | new_D2261_;
  assign new_D2248_ = new_D2257_ & new_D2260_;
  assign new_D2249_ = new_D2232_ | new_D2265_;
  assign new_D2250_ = new_D2264_ | new_D2263_;
  assign new_D2251_ = new_D2267_ | new_D2266_;
  assign new_D2252_ = ~new_D2243_ & new_D2269_;
  assign new_D2253_ = ~new_D2245_ & new_D2257_;
  assign new_D2254_ = new_D2245_ & ~new_D2257_;
  assign new_D2255_ = new_D2231_ & ~new_D2232_;
  assign new_D2256_ = ~new_D2278_ | ~new_D2279_;
  assign new_D2257_ = new_D2271_ | new_D2273_;
  assign new_D2258_ = new_D2281_ | new_D2280_;
  assign new_D2259_ = new_D2275_ | new_D2274_;
  assign new_D2260_ = ~new_D2283_ | ~new_D2282_;
  assign new_D2261_ = ~new_D2284_ & new_D2285_;
  assign new_D2262_ = new_D2284_ & ~new_D2285_;
  assign new_D2263_ = ~new_D2231_ & new_D2232_;
  assign new_D2264_ = new_D2231_ & ~new_D2232_;
  assign new_D2265_ = ~new_D2247_ | new_D2257_;
  assign new_D2266_ = new_D2247_ & new_D2257_;
  assign new_D2267_ = ~new_D2247_ & ~new_D2257_;
  assign new_D2268_ = new_D2289_ | new_D2288_;
  assign new_D2269_ = new_D2235_ | new_D2268_;
  assign new_D2270_ = new_D2293_ | new_D2292_;
  assign new_D2271_ = ~new_D2235_ & new_D2270_;
  assign new_D2272_ = new_D2291_ | new_D2290_;
  assign new_D2273_ = new_D2235_ & new_D2272_;
  assign new_D2274_ = new_D2233_ & ~new_D2243_;
  assign new_D2275_ = ~new_D2233_ & new_D2243_;
  assign new_D2276_ = ~new_D2232_ | ~new_D2257_;
  assign new_D2277_ = new_D2243_ & new_D2276_;
  assign new_D2278_ = ~new_D2243_ & ~new_D2277_;
  assign new_D2279_ = new_D2243_ | new_D2276_;
  assign new_D2280_ = ~new_D2233_ & new_D2234_;
  assign new_D2281_ = new_D2233_ & ~new_D2234_;
  assign new_D2282_ = new_D2250_ | new_D2287_;
  assign new_D2283_ = ~new_D2250_ & ~new_D2286_;
  assign new_D2284_ = new_D2233_ | new_D2250_;
  assign new_D2285_ = new_D2233_ | new_D2234_;
  assign new_D2286_ = new_D2250_ & new_D2287_;
  assign new_D2287_ = ~new_D2232_ | ~new_D2257_;
  assign new_D2288_ = new_D2265_ & new_D2285_;
  assign new_D2289_ = ~new_D2265_ & ~new_D2285_;
  assign new_D2290_ = new_D2294_ | new_D2295_;
  assign new_D2291_ = ~new_D2236_ & new_D2250_;
  assign new_D2292_ = new_D2296_ | new_D2297_;
  assign new_D2293_ = new_D2236_ & new_D2250_;
  assign new_D2294_ = ~new_D2236_ & ~new_D2250_;
  assign new_D2295_ = new_D2236_ & ~new_D2250_;
  assign new_D2296_ = new_D2236_ & ~new_D2250_;
  assign new_D2297_ = ~new_D2236_ & new_D2250_;
  assign new_D2298_ = new_D7802_;
  assign new_D2299_ = new_D7869_;
  assign new_D2300_ = new_D7936_;
  assign new_D2301_ = new_D8003_;
  assign new_D2302_ = new_D8070_;
  assign new_D2303_ = new_D8137_;
  assign new_D2304_ = new_D2311_ & new_D2310_;
  assign new_D2305_ = new_D2313_ | new_D2312_;
  assign new_D2306_ = new_D2315_ | new_D2314_;
  assign new_D2307_ = new_D2317_ & new_D2316_;
  assign new_D2308_ = new_D2317_ & new_D2318_;
  assign new_D2309_ = new_D2310_ | new_D2319_;
  assign new_D2310_ = new_D2299_ | new_D2322_;
  assign new_D2311_ = new_D2321_ | new_D2320_;
  assign new_D2312_ = new_D2326_ & new_D2325_;
  assign new_D2313_ = new_D2324_ & new_D2323_;
  assign new_D2314_ = new_D2329_ | new_D2328_;
  assign new_D2315_ = new_D2324_ & new_D2327_;
  assign new_D2316_ = new_D2299_ | new_D2332_;
  assign new_D2317_ = new_D2331_ | new_D2330_;
  assign new_D2318_ = new_D2334_ | new_D2333_;
  assign new_D2319_ = ~new_D2310_ & new_D2336_;
  assign new_D2320_ = ~new_D2312_ & new_D2324_;
  assign new_D2321_ = new_D2312_ & ~new_D2324_;
  assign new_D2322_ = new_D2298_ & ~new_D2299_;
  assign new_D2323_ = ~new_D2345_ | ~new_D2346_;
  assign new_D2324_ = new_D2338_ | new_D2340_;
  assign new_D2325_ = new_D2348_ | new_D2347_;
  assign new_D2326_ = new_D2342_ | new_D2341_;
  assign new_D2327_ = ~new_D2350_ | ~new_D2349_;
  assign new_D2328_ = ~new_D2351_ & new_D2352_;
  assign new_D2329_ = new_D2351_ & ~new_D2352_;
  assign new_D2330_ = ~new_D2298_ & new_D2299_;
  assign new_D2331_ = new_D2298_ & ~new_D2299_;
  assign new_D2332_ = ~new_D2314_ | new_D2324_;
  assign new_D2333_ = new_D2314_ & new_D2324_;
  assign new_D2334_ = ~new_D2314_ & ~new_D2324_;
  assign new_D2335_ = new_D2356_ | new_D2355_;
  assign new_D2336_ = new_D2302_ | new_D2335_;
  assign new_D2337_ = new_D2360_ | new_D2359_;
  assign new_D2338_ = ~new_D2302_ & new_D2337_;
  assign new_D2339_ = new_D2358_ | new_D2357_;
  assign new_D2340_ = new_D2302_ & new_D2339_;
  assign new_D2341_ = new_D2300_ & ~new_D2310_;
  assign new_D2342_ = ~new_D2300_ & new_D2310_;
  assign new_D2343_ = ~new_D2299_ | ~new_D2324_;
  assign new_D2344_ = new_D2310_ & new_D2343_;
  assign new_D2345_ = ~new_D2310_ & ~new_D2344_;
  assign new_D2346_ = new_D2310_ | new_D2343_;
  assign new_D2347_ = ~new_D2300_ & new_D2301_;
  assign new_D2348_ = new_D2300_ & ~new_D2301_;
  assign new_D2349_ = new_D2317_ | new_D2354_;
  assign new_D2350_ = ~new_D2317_ & ~new_D2353_;
  assign new_D2351_ = new_D2300_ | new_D2317_;
  assign new_D2352_ = new_D2300_ | new_D2301_;
  assign new_D2353_ = new_D2317_ & new_D2354_;
  assign new_D2354_ = ~new_D2299_ | ~new_D2324_;
  assign new_D2355_ = new_D2332_ & new_D2352_;
  assign new_D2356_ = ~new_D2332_ & ~new_D2352_;
  assign new_D2357_ = new_D2361_ | new_D2362_;
  assign new_D2358_ = ~new_D2303_ & new_D2317_;
  assign new_D2359_ = new_D2363_ | new_D2364_;
  assign new_D2360_ = new_D2303_ & new_D2317_;
  assign new_D2361_ = ~new_D2303_ & ~new_D2317_;
  assign new_D2362_ = new_D2303_ & ~new_D2317_;
  assign new_D2363_ = new_D2303_ & ~new_D2317_;
  assign new_D2364_ = ~new_D2303_ & new_D2317_;
  assign new_D2365_ = new_D8204_;
  assign new_D2366_ = new_D8271_;
  assign new_D2367_ = new_D8338_;
  assign new_D2368_ = new_D8405_;
  assign new_D2369_ = new_D8472_;
  assign new_D2370_ = new_D8539_;
  assign new_D2371_ = new_D2378_ & new_D2377_;
  assign new_D2372_ = new_D2380_ | new_D2379_;
  assign new_D2373_ = new_D2382_ | new_D2381_;
  assign new_D2374_ = new_D2384_ & new_D2383_;
  assign new_D2375_ = new_D2384_ & new_D2385_;
  assign new_D2376_ = new_D2377_ | new_D2386_;
  assign new_D2377_ = new_D2366_ | new_D2389_;
  assign new_D2378_ = new_D2388_ | new_D2387_;
  assign new_D2379_ = new_D2393_ & new_D2392_;
  assign new_D2380_ = new_D2391_ & new_D2390_;
  assign new_D2381_ = new_D2396_ | new_D2395_;
  assign new_D2382_ = new_D2391_ & new_D2394_;
  assign new_D2383_ = new_D2366_ | new_D2399_;
  assign new_D2384_ = new_D2398_ | new_D2397_;
  assign new_D2385_ = new_D2401_ | new_D2400_;
  assign new_D2386_ = ~new_D2377_ & new_D2403_;
  assign new_D2387_ = ~new_D2379_ & new_D2391_;
  assign new_D2388_ = new_D2379_ & ~new_D2391_;
  assign new_D2389_ = new_D2365_ & ~new_D2366_;
  assign new_D2390_ = ~new_D2412_ | ~new_D2413_;
  assign new_D2391_ = new_D2405_ | new_D2407_;
  assign new_D2392_ = new_D2415_ | new_D2414_;
  assign new_D2393_ = new_D2409_ | new_D2408_;
  assign new_D2394_ = ~new_D2417_ | ~new_D2416_;
  assign new_D2395_ = ~new_D2418_ & new_D2419_;
  assign new_D2396_ = new_D2418_ & ~new_D2419_;
  assign new_D2397_ = ~new_D2365_ & new_D2366_;
  assign new_D2398_ = new_D2365_ & ~new_D2366_;
  assign new_D2399_ = ~new_D2381_ | new_D2391_;
  assign new_D2400_ = new_D2381_ & new_D2391_;
  assign new_D2401_ = ~new_D2381_ & ~new_D2391_;
  assign new_D2402_ = new_D2423_ | new_D2422_;
  assign new_D2403_ = new_D2369_ | new_D2402_;
  assign new_D2404_ = new_D2427_ | new_D2426_;
  assign new_D2405_ = ~new_D2369_ & new_D2404_;
  assign new_D2406_ = new_D2425_ | new_D2424_;
  assign new_D2407_ = new_D2369_ & new_D2406_;
  assign new_D2408_ = new_D2367_ & ~new_D2377_;
  assign new_D2409_ = ~new_D2367_ & new_D2377_;
  assign new_D2410_ = ~new_D2366_ | ~new_D2391_;
  assign new_D2411_ = new_D2377_ & new_D2410_;
  assign new_D2412_ = ~new_D2377_ & ~new_D2411_;
  assign new_D2413_ = new_D2377_ | new_D2410_;
  assign new_D2414_ = ~new_D2367_ & new_D2368_;
  assign new_D2415_ = new_D2367_ & ~new_D2368_;
  assign new_D2416_ = new_D2384_ | new_D2421_;
  assign new_D2417_ = ~new_D2384_ & ~new_D2420_;
  assign new_D2418_ = new_D2367_ | new_D2384_;
  assign new_D2419_ = new_D2367_ | new_D2368_;
  assign new_D2420_ = new_D2384_ & new_D2421_;
  assign new_D2421_ = ~new_D2366_ | ~new_D2391_;
  assign new_D2422_ = new_D2399_ & new_D2419_;
  assign new_D2423_ = ~new_D2399_ & ~new_D2419_;
  assign new_D2424_ = new_D2428_ | new_D2429_;
  assign new_D2425_ = ~new_D2370_ & new_D2384_;
  assign new_D2426_ = new_D2430_ | new_D2431_;
  assign new_D2427_ = new_D2370_ & new_D2384_;
  assign new_D2428_ = ~new_D2370_ & ~new_D2384_;
  assign new_D2429_ = new_D2370_ & ~new_D2384_;
  assign new_D2430_ = new_D2370_ & ~new_D2384_;
  assign new_D2431_ = ~new_D2370_ & new_D2384_;
  assign new_D2432_ = new_D8606_;
  assign new_D2433_ = new_D8673_;
  assign new_D2434_ = new_D8740_;
  assign new_D2435_ = new_D8807_;
  assign new_D2436_ = new_D8874_;
  assign new_D2437_ = new_D8941_;
  assign new_D2438_ = new_D2445_ & new_D2444_;
  assign new_D2439_ = new_D2447_ | new_D2446_;
  assign new_D2440_ = new_D2449_ | new_D2448_;
  assign new_D2441_ = new_D2451_ & new_D2450_;
  assign new_D2442_ = new_D2451_ & new_D2452_;
  assign new_D2443_ = new_D2444_ | new_D2453_;
  assign new_D2444_ = new_D2433_ | new_D2456_;
  assign new_D2445_ = new_D2455_ | new_D2454_;
  assign new_D2446_ = new_D2460_ & new_D2459_;
  assign new_D2447_ = new_D2458_ & new_D2457_;
  assign new_D2448_ = new_D2463_ | new_D2462_;
  assign new_D2449_ = new_D2458_ & new_D2461_;
  assign new_D2450_ = new_D2433_ | new_D2466_;
  assign new_D2451_ = new_D2465_ | new_D2464_;
  assign new_D2452_ = new_D2468_ | new_D2467_;
  assign new_D2453_ = ~new_D2444_ & new_D2470_;
  assign new_D2454_ = ~new_D2446_ & new_D2458_;
  assign new_D2455_ = new_D2446_ & ~new_D2458_;
  assign new_D2456_ = new_D2432_ & ~new_D2433_;
  assign new_D2457_ = ~new_D2479_ | ~new_D2480_;
  assign new_D2458_ = new_D2472_ | new_D2474_;
  assign new_D2459_ = new_D2482_ | new_D2481_;
  assign new_D2460_ = new_D2476_ | new_D2475_;
  assign new_D2461_ = ~new_D2484_ | ~new_D2483_;
  assign new_D2462_ = ~new_D2485_ & new_D2486_;
  assign new_D2463_ = new_D2485_ & ~new_D2486_;
  assign new_D2464_ = ~new_D2432_ & new_D2433_;
  assign new_D2465_ = new_D2432_ & ~new_D2433_;
  assign new_D2466_ = ~new_D2448_ | new_D2458_;
  assign new_D2467_ = new_D2448_ & new_D2458_;
  assign new_D2468_ = ~new_D2448_ & ~new_D2458_;
  assign new_D2469_ = new_D2490_ | new_D2489_;
  assign new_D2470_ = new_D2436_ | new_D2469_;
  assign new_D2471_ = new_D2494_ | new_D2493_;
  assign new_D2472_ = ~new_D2436_ & new_D2471_;
  assign new_D2473_ = new_D2492_ | new_D2491_;
  assign new_D2474_ = new_D2436_ & new_D2473_;
  assign new_D2475_ = new_D2434_ & ~new_D2444_;
  assign new_D2476_ = ~new_D2434_ & new_D2444_;
  assign new_D2477_ = ~new_D2433_ | ~new_D2458_;
  assign new_D2478_ = new_D2444_ & new_D2477_;
  assign new_D2479_ = ~new_D2444_ & ~new_D2478_;
  assign new_D2480_ = new_D2444_ | new_D2477_;
  assign new_D2481_ = ~new_D2434_ & new_D2435_;
  assign new_D2482_ = new_D2434_ & ~new_D2435_;
  assign new_D2483_ = new_D2451_ | new_D2488_;
  assign new_D2484_ = ~new_D2451_ & ~new_D2487_;
  assign new_D2485_ = new_D2434_ | new_D2451_;
  assign new_D2486_ = new_D2434_ | new_D2435_;
  assign new_D2487_ = new_D2451_ & new_D2488_;
  assign new_D2488_ = ~new_D2433_ | ~new_D2458_;
  assign new_D2489_ = new_D2466_ & new_D2486_;
  assign new_D2490_ = ~new_D2466_ & ~new_D2486_;
  assign new_D2491_ = new_D2495_ | new_D2496_;
  assign new_D2492_ = ~new_D2437_ & new_D2451_;
  assign new_D2493_ = new_D2497_ | new_D2498_;
  assign new_D2494_ = new_D2437_ & new_D2451_;
  assign new_D2495_ = ~new_D2437_ & ~new_D2451_;
  assign new_D2496_ = new_D2437_ & ~new_D2451_;
  assign new_D2497_ = new_D2437_ & ~new_D2451_;
  assign new_D2498_ = ~new_D2437_ & new_D2451_;
  assign new_D2499_ = new_D9008_;
  assign new_D2500_ = new_D9075_;
  assign new_D2501_ = new_D9142_;
  assign new_D2502_ = new_D9209_;
  assign new_D2503_ = new_D9276_;
  assign new_D2504_ = new_D9343_;
  assign new_D2505_ = new_D2512_ & new_D2511_;
  assign new_D2506_ = new_D2514_ | new_D2513_;
  assign new_D2507_ = new_D2516_ | new_D2515_;
  assign new_D2508_ = new_D2518_ & new_D2517_;
  assign new_D2509_ = new_D2518_ & new_D2519_;
  assign new_D2510_ = new_D2511_ | new_D2520_;
  assign new_D2511_ = new_D2500_ | new_D2523_;
  assign new_D2512_ = new_D2522_ | new_D2521_;
  assign new_D2513_ = new_D2527_ & new_D2526_;
  assign new_D2514_ = new_D2525_ & new_D2524_;
  assign new_D2515_ = new_D2530_ | new_D2529_;
  assign new_D2516_ = new_D2525_ & new_D2528_;
  assign new_D2517_ = new_D2500_ | new_D2533_;
  assign new_D2518_ = new_D2532_ | new_D2531_;
  assign new_D2519_ = new_D2535_ | new_D2534_;
  assign new_D2520_ = ~new_D2511_ & new_D2537_;
  assign new_D2521_ = ~new_D2513_ & new_D2525_;
  assign new_D2522_ = new_D2513_ & ~new_D2525_;
  assign new_D2523_ = new_D2499_ & ~new_D2500_;
  assign new_D2524_ = ~new_D2546_ | ~new_D2547_;
  assign new_D2525_ = new_D2539_ | new_D2541_;
  assign new_D2526_ = new_D2549_ | new_D2548_;
  assign new_D2527_ = new_D2543_ | new_D2542_;
  assign new_D2528_ = ~new_D2551_ | ~new_D2550_;
  assign new_D2529_ = ~new_D2552_ & new_D2553_;
  assign new_D2530_ = new_D2552_ & ~new_D2553_;
  assign new_D2531_ = ~new_D2499_ & new_D2500_;
  assign new_D2532_ = new_D2499_ & ~new_D2500_;
  assign new_D2533_ = ~new_D2515_ | new_D2525_;
  assign new_D2534_ = new_D2515_ & new_D2525_;
  assign new_D2535_ = ~new_D2515_ & ~new_D2525_;
  assign new_D2536_ = new_D2557_ | new_D2556_;
  assign new_D2537_ = new_D2503_ | new_D2536_;
  assign new_D2538_ = new_D2561_ | new_D2560_;
  assign new_D2539_ = ~new_D2503_ & new_D2538_;
  assign new_D2540_ = new_D2559_ | new_D2558_;
  assign new_D2541_ = new_D2503_ & new_D2540_;
  assign new_D2542_ = new_D2501_ & ~new_D2511_;
  assign new_D2543_ = ~new_D2501_ & new_D2511_;
  assign new_D2544_ = ~new_D2500_ | ~new_D2525_;
  assign new_D2545_ = new_D2511_ & new_D2544_;
  assign new_D2546_ = ~new_D2511_ & ~new_D2545_;
  assign new_D2547_ = new_D2511_ | new_D2544_;
  assign new_D2548_ = ~new_D2501_ & new_D2502_;
  assign new_D2549_ = new_D2501_ & ~new_D2502_;
  assign new_D2550_ = new_D2518_ | new_D2555_;
  assign new_D2551_ = ~new_D2518_ & ~new_D2554_;
  assign new_D2552_ = new_D2501_ | new_D2518_;
  assign new_D2553_ = new_D2501_ | new_D2502_;
  assign new_D2554_ = new_D2518_ & new_D2555_;
  assign new_D2555_ = ~new_D2500_ | ~new_D2525_;
  assign new_D2556_ = new_D2533_ & new_D2553_;
  assign new_D2557_ = ~new_D2533_ & ~new_D2553_;
  assign new_D2558_ = new_D2562_ | new_D2563_;
  assign new_D2559_ = ~new_D2504_ & new_D2518_;
  assign new_D2560_ = new_D2564_ | new_D2565_;
  assign new_D2561_ = new_D2504_ & new_D2518_;
  assign new_D2562_ = ~new_D2504_ & ~new_D2518_;
  assign new_D2563_ = new_D2504_ & ~new_D2518_;
  assign new_D2564_ = new_D2504_ & ~new_D2518_;
  assign new_D2565_ = ~new_D2504_ & new_D2518_;
  assign new_D2566_ = new_D9410_;
  assign new_D2567_ = new_D9477_;
  assign new_D2568_ = new_D9544_;
  assign new_D2569_ = new_D9611_;
  assign new_D2570_ = new_D9678_;
  assign new_D2571_ = new_D9745_;
  assign new_D2572_ = new_D2579_ & new_D2578_;
  assign new_D2573_ = new_D2581_ | new_D2580_;
  assign new_D2574_ = new_D2583_ | new_D2582_;
  assign new_D2575_ = new_D2585_ & new_D2584_;
  assign new_D2576_ = new_D2585_ & new_D2586_;
  assign new_D2577_ = new_D2578_ | new_D2587_;
  assign new_D2578_ = new_D2567_ | new_D2590_;
  assign new_D2579_ = new_D2589_ | new_D2588_;
  assign new_D2580_ = new_D2594_ & new_D2593_;
  assign new_D2581_ = new_D2592_ & new_D2591_;
  assign new_D2582_ = new_D2597_ | new_D2596_;
  assign new_D2583_ = new_D2592_ & new_D2595_;
  assign new_D2584_ = new_D2567_ | new_D2600_;
  assign new_D2585_ = new_D2599_ | new_D2598_;
  assign new_D2586_ = new_D2602_ | new_D2601_;
  assign new_D2587_ = ~new_D2578_ & new_D2604_;
  assign new_D2588_ = ~new_D2580_ & new_D2592_;
  assign new_D2589_ = new_D2580_ & ~new_D2592_;
  assign new_D2590_ = new_D2566_ & ~new_D2567_;
  assign new_D2591_ = ~new_D2613_ | ~new_D2614_;
  assign new_D2592_ = new_D2606_ | new_D2608_;
  assign new_D2593_ = new_D2616_ | new_D2615_;
  assign new_D2594_ = new_D2610_ | new_D2609_;
  assign new_D2595_ = ~new_D2618_ | ~new_D2617_;
  assign new_D2596_ = ~new_D2619_ & new_D2620_;
  assign new_D2597_ = new_D2619_ & ~new_D2620_;
  assign new_D2598_ = ~new_D2566_ & new_D2567_;
  assign new_D2599_ = new_D2566_ & ~new_D2567_;
  assign new_D2600_ = ~new_D2582_ | new_D2592_;
  assign new_D2601_ = new_D2582_ & new_D2592_;
  assign new_D2602_ = ~new_D2582_ & ~new_D2592_;
  assign new_D2603_ = new_D2624_ | new_D2623_;
  assign new_D2604_ = new_D2570_ | new_D2603_;
  assign new_D2605_ = new_D2628_ | new_D2627_;
  assign new_D2606_ = ~new_D2570_ & new_D2605_;
  assign new_D2607_ = new_D2626_ | new_D2625_;
  assign new_D2608_ = new_D2570_ & new_D2607_;
  assign new_D2609_ = new_D2568_ & ~new_D2578_;
  assign new_D2610_ = ~new_D2568_ & new_D2578_;
  assign new_D2611_ = ~new_D2567_ | ~new_D2592_;
  assign new_D2612_ = new_D2578_ & new_D2611_;
  assign new_D2613_ = ~new_D2578_ & ~new_D2612_;
  assign new_D2614_ = new_D2578_ | new_D2611_;
  assign new_D2615_ = ~new_D2568_ & new_D2569_;
  assign new_D2616_ = new_D2568_ & ~new_D2569_;
  assign new_D2617_ = new_D2585_ | new_D2622_;
  assign new_D2618_ = ~new_D2585_ & ~new_D2621_;
  assign new_D2619_ = new_D2568_ | new_D2585_;
  assign new_D2620_ = new_D2568_ | new_D2569_;
  assign new_D2621_ = new_D2585_ & new_D2622_;
  assign new_D2622_ = ~new_D2567_ | ~new_D2592_;
  assign new_D2623_ = new_D2600_ & new_D2620_;
  assign new_D2624_ = ~new_D2600_ & ~new_D2620_;
  assign new_D2625_ = new_D2629_ | new_D2630_;
  assign new_D2626_ = ~new_D2571_ & new_D2585_;
  assign new_D2627_ = new_D2631_ | new_D2632_;
  assign new_D2628_ = new_D2571_ & new_D2585_;
  assign new_D2629_ = ~new_D2571_ & ~new_D2585_;
  assign new_D2630_ = new_D2571_ & ~new_D2585_;
  assign new_D2631_ = new_D2571_ & ~new_D2585_;
  assign new_D2632_ = ~new_D2571_ & new_D2585_;
  assign new_D2633_ = new_D9812_;
  assign new_D2634_ = new_D9879_;
  assign new_D2635_ = new_D9946_;
  assign new_D2636_ = new_E14_;
  assign new_D2637_ = new_E81_;
  assign new_D2638_ = new_E148_;
  assign new_D2639_ = new_D2646_ & new_D2645_;
  assign new_D2640_ = new_D2648_ | new_D2647_;
  assign new_D2641_ = new_D2650_ | new_D2649_;
  assign new_D2642_ = new_D2652_ & new_D2651_;
  assign new_D2643_ = new_D2652_ & new_D2653_;
  assign new_D2644_ = new_D2645_ | new_D2654_;
  assign new_D2645_ = new_D2634_ | new_D2657_;
  assign new_D2646_ = new_D2656_ | new_D2655_;
  assign new_D2647_ = new_D2661_ & new_D2660_;
  assign new_D2648_ = new_D2659_ & new_D2658_;
  assign new_D2649_ = new_D2664_ | new_D2663_;
  assign new_D2650_ = new_D2659_ & new_D2662_;
  assign new_D2651_ = new_D2634_ | new_D2667_;
  assign new_D2652_ = new_D2666_ | new_D2665_;
  assign new_D2653_ = new_D2669_ | new_D2668_;
  assign new_D2654_ = ~new_D2645_ & new_D2671_;
  assign new_D2655_ = ~new_D2647_ & new_D2659_;
  assign new_D2656_ = new_D2647_ & ~new_D2659_;
  assign new_D2657_ = new_D2633_ & ~new_D2634_;
  assign new_D2658_ = ~new_D2680_ | ~new_D2681_;
  assign new_D2659_ = new_D2673_ | new_D2675_;
  assign new_D2660_ = new_D2683_ | new_D2682_;
  assign new_D2661_ = new_D2677_ | new_D2676_;
  assign new_D2662_ = ~new_D2685_ | ~new_D2684_;
  assign new_D2663_ = ~new_D2686_ & new_D2687_;
  assign new_D2664_ = new_D2686_ & ~new_D2687_;
  assign new_D2665_ = ~new_D2633_ & new_D2634_;
  assign new_D2666_ = new_D2633_ & ~new_D2634_;
  assign new_D2667_ = ~new_D2649_ | new_D2659_;
  assign new_D2668_ = new_D2649_ & new_D2659_;
  assign new_D2669_ = ~new_D2649_ & ~new_D2659_;
  assign new_D2670_ = new_D2691_ | new_D2690_;
  assign new_D2671_ = new_D2637_ | new_D2670_;
  assign new_D2672_ = new_D2695_ | new_D2694_;
  assign new_D2673_ = ~new_D2637_ & new_D2672_;
  assign new_D2674_ = new_D2693_ | new_D2692_;
  assign new_D2675_ = new_D2637_ & new_D2674_;
  assign new_D2676_ = new_D2635_ & ~new_D2645_;
  assign new_D2677_ = ~new_D2635_ & new_D2645_;
  assign new_D2678_ = ~new_D2634_ | ~new_D2659_;
  assign new_D2679_ = new_D2645_ & new_D2678_;
  assign new_D2680_ = ~new_D2645_ & ~new_D2679_;
  assign new_D2681_ = new_D2645_ | new_D2678_;
  assign new_D2682_ = ~new_D2635_ & new_D2636_;
  assign new_D2683_ = new_D2635_ & ~new_D2636_;
  assign new_D2684_ = new_D2652_ | new_D2689_;
  assign new_D2685_ = ~new_D2652_ & ~new_D2688_;
  assign new_D2686_ = new_D2635_ | new_D2652_;
  assign new_D2687_ = new_D2635_ | new_D2636_;
  assign new_D2688_ = new_D2652_ & new_D2689_;
  assign new_D2689_ = ~new_D2634_ | ~new_D2659_;
  assign new_D2690_ = new_D2667_ & new_D2687_;
  assign new_D2691_ = ~new_D2667_ & ~new_D2687_;
  assign new_D2692_ = new_D2696_ | new_D2697_;
  assign new_D2693_ = ~new_D2638_ & new_D2652_;
  assign new_D2694_ = new_D2698_ | new_D2699_;
  assign new_D2695_ = new_D2638_ & new_D2652_;
  assign new_D2696_ = ~new_D2638_ & ~new_D2652_;
  assign new_D2697_ = new_D2638_ & ~new_D2652_;
  assign new_D2698_ = new_D2638_ & ~new_D2652_;
  assign new_D2699_ = ~new_D2638_ & new_D2652_;
  assign new_D2700_ = new_E215_;
  assign new_D2701_ = new_E282_;
  assign new_D2702_ = new_E349_;
  assign new_D2703_ = new_E416_;
  assign new_D2704_ = new_E483_;
  assign new_D2705_ = new_E550_;
  assign new_D2706_ = new_D2713_ & new_D2712_;
  assign new_D2707_ = new_D2715_ | new_D2714_;
  assign new_D2708_ = new_D2717_ | new_D2716_;
  assign new_D2709_ = new_D2719_ & new_D2718_;
  assign new_D2710_ = new_D2719_ & new_D2720_;
  assign new_D2711_ = new_D2712_ | new_D2721_;
  assign new_D2712_ = new_D2701_ | new_D2724_;
  assign new_D2713_ = new_D2723_ | new_D2722_;
  assign new_D2714_ = new_D2728_ & new_D2727_;
  assign new_D2715_ = new_D2726_ & new_D2725_;
  assign new_D2716_ = new_D2731_ | new_D2730_;
  assign new_D2717_ = new_D2726_ & new_D2729_;
  assign new_D2718_ = new_D2701_ | new_D2734_;
  assign new_D2719_ = new_D2733_ | new_D2732_;
  assign new_D2720_ = new_D2736_ | new_D2735_;
  assign new_D2721_ = ~new_D2712_ & new_D2738_;
  assign new_D2722_ = ~new_D2714_ & new_D2726_;
  assign new_D2723_ = new_D2714_ & ~new_D2726_;
  assign new_D2724_ = new_D2700_ & ~new_D2701_;
  assign new_D2725_ = ~new_D2747_ | ~new_D2748_;
  assign new_D2726_ = new_D2740_ | new_D2742_;
  assign new_D2727_ = new_D2750_ | new_D2749_;
  assign new_D2728_ = new_D2744_ | new_D2743_;
  assign new_D2729_ = ~new_D2752_ | ~new_D2751_;
  assign new_D2730_ = ~new_D2753_ & new_D2754_;
  assign new_D2731_ = new_D2753_ & ~new_D2754_;
  assign new_D2732_ = ~new_D2700_ & new_D2701_;
  assign new_D2733_ = new_D2700_ & ~new_D2701_;
  assign new_D2734_ = ~new_D2716_ | new_D2726_;
  assign new_D2735_ = new_D2716_ & new_D2726_;
  assign new_D2736_ = ~new_D2716_ & ~new_D2726_;
  assign new_D2737_ = new_D2758_ | new_D2757_;
  assign new_D2738_ = new_D2704_ | new_D2737_;
  assign new_D2739_ = new_D2762_ | new_D2761_;
  assign new_D2740_ = ~new_D2704_ & new_D2739_;
  assign new_D2741_ = new_D2760_ | new_D2759_;
  assign new_D2742_ = new_D2704_ & new_D2741_;
  assign new_D2743_ = new_D2702_ & ~new_D2712_;
  assign new_D2744_ = ~new_D2702_ & new_D2712_;
  assign new_D2745_ = ~new_D2701_ | ~new_D2726_;
  assign new_D2746_ = new_D2712_ & new_D2745_;
  assign new_D2747_ = ~new_D2712_ & ~new_D2746_;
  assign new_D2748_ = new_D2712_ | new_D2745_;
  assign new_D2749_ = ~new_D2702_ & new_D2703_;
  assign new_D2750_ = new_D2702_ & ~new_D2703_;
  assign new_D2751_ = new_D2719_ | new_D2756_;
  assign new_D2752_ = ~new_D2719_ & ~new_D2755_;
  assign new_D2753_ = new_D2702_ | new_D2719_;
  assign new_D2754_ = new_D2702_ | new_D2703_;
  assign new_D2755_ = new_D2719_ & new_D2756_;
  assign new_D2756_ = ~new_D2701_ | ~new_D2726_;
  assign new_D2757_ = new_D2734_ & new_D2754_;
  assign new_D2758_ = ~new_D2734_ & ~new_D2754_;
  assign new_D2759_ = new_D2763_ | new_D2764_;
  assign new_D2760_ = ~new_D2705_ & new_D2719_;
  assign new_D2761_ = new_D2765_ | new_D2766_;
  assign new_D2762_ = new_D2705_ & new_D2719_;
  assign new_D2763_ = ~new_D2705_ & ~new_D2719_;
  assign new_D2764_ = new_D2705_ & ~new_D2719_;
  assign new_D2765_ = new_D2705_ & ~new_D2719_;
  assign new_D2766_ = ~new_D2705_ & new_D2719_;
  assign new_D2767_ = new_E617_;
  assign new_D2768_ = new_E684_;
  assign new_D2769_ = new_E751_;
  assign new_D2770_ = new_E818_;
  assign new_D2771_ = new_E885_;
  assign new_D2772_ = new_E952_;
  assign new_D2773_ = new_D2780_ & new_D2779_;
  assign new_D2774_ = new_D2782_ | new_D2781_;
  assign new_D2775_ = new_D2784_ | new_D2783_;
  assign new_D2776_ = new_D2786_ & new_D2785_;
  assign new_D2777_ = new_D2786_ & new_D2787_;
  assign new_D2778_ = new_D2779_ | new_D2788_;
  assign new_D2779_ = new_D2768_ | new_D2791_;
  assign new_D2780_ = new_D2790_ | new_D2789_;
  assign new_D2781_ = new_D2795_ & new_D2794_;
  assign new_D2782_ = new_D2793_ & new_D2792_;
  assign new_D2783_ = new_D2798_ | new_D2797_;
  assign new_D2784_ = new_D2793_ & new_D2796_;
  assign new_D2785_ = new_D2768_ | new_D2801_;
  assign new_D2786_ = new_D2800_ | new_D2799_;
  assign new_D2787_ = new_D2803_ | new_D2802_;
  assign new_D2788_ = ~new_D2779_ & new_D2805_;
  assign new_D2789_ = ~new_D2781_ & new_D2793_;
  assign new_D2790_ = new_D2781_ & ~new_D2793_;
  assign new_D2791_ = new_D2767_ & ~new_D2768_;
  assign new_D2792_ = ~new_D2814_ | ~new_D2815_;
  assign new_D2793_ = new_D2807_ | new_D2809_;
  assign new_D2794_ = new_D2817_ | new_D2816_;
  assign new_D2795_ = new_D2811_ | new_D2810_;
  assign new_D2796_ = ~new_D2819_ | ~new_D2818_;
  assign new_D2797_ = ~new_D2820_ & new_D2821_;
  assign new_D2798_ = new_D2820_ & ~new_D2821_;
  assign new_D2799_ = ~new_D2767_ & new_D2768_;
  assign new_D2800_ = new_D2767_ & ~new_D2768_;
  assign new_D2801_ = ~new_D2783_ | new_D2793_;
  assign new_D2802_ = new_D2783_ & new_D2793_;
  assign new_D2803_ = ~new_D2783_ & ~new_D2793_;
  assign new_D2804_ = new_D2825_ | new_D2824_;
  assign new_D2805_ = new_D2771_ | new_D2804_;
  assign new_D2806_ = new_D2829_ | new_D2828_;
  assign new_D2807_ = ~new_D2771_ & new_D2806_;
  assign new_D2808_ = new_D2827_ | new_D2826_;
  assign new_D2809_ = new_D2771_ & new_D2808_;
  assign new_D2810_ = new_D2769_ & ~new_D2779_;
  assign new_D2811_ = ~new_D2769_ & new_D2779_;
  assign new_D2812_ = ~new_D2768_ | ~new_D2793_;
  assign new_D2813_ = new_D2779_ & new_D2812_;
  assign new_D2814_ = ~new_D2779_ & ~new_D2813_;
  assign new_D2815_ = new_D2779_ | new_D2812_;
  assign new_D2816_ = ~new_D2769_ & new_D2770_;
  assign new_D2817_ = new_D2769_ & ~new_D2770_;
  assign new_D2818_ = new_D2786_ | new_D2823_;
  assign new_D2819_ = ~new_D2786_ & ~new_D2822_;
  assign new_D2820_ = new_D2769_ | new_D2786_;
  assign new_D2821_ = new_D2769_ | new_D2770_;
  assign new_D2822_ = new_D2786_ & new_D2823_;
  assign new_D2823_ = ~new_D2768_ | ~new_D2793_;
  assign new_D2824_ = new_D2801_ & new_D2821_;
  assign new_D2825_ = ~new_D2801_ & ~new_D2821_;
  assign new_D2826_ = new_D2830_ | new_D2831_;
  assign new_D2827_ = ~new_D2772_ & new_D2786_;
  assign new_D2828_ = new_D2832_ | new_D2833_;
  assign new_D2829_ = new_D2772_ & new_D2786_;
  assign new_D2830_ = ~new_D2772_ & ~new_D2786_;
  assign new_D2831_ = new_D2772_ & ~new_D2786_;
  assign new_D2832_ = new_D2772_ & ~new_D2786_;
  assign new_D2833_ = ~new_D2772_ & new_D2786_;
  assign new_D2834_ = new_E1019_;
  assign new_D2835_ = new_E1086_;
  assign new_D2836_ = new_E1153_;
  assign new_D2837_ = new_E1220_;
  assign new_D2838_ = new_E1287_;
  assign new_D2839_ = new_E1354_;
  assign new_D2840_ = new_D2847_ & new_D2846_;
  assign new_D2841_ = new_D2849_ | new_D2848_;
  assign new_D2842_ = new_D2851_ | new_D2850_;
  assign new_D2843_ = new_D2853_ & new_D2852_;
  assign new_D2844_ = new_D2853_ & new_D2854_;
  assign new_D2845_ = new_D2846_ | new_D2855_;
  assign new_D2846_ = new_D2835_ | new_D2858_;
  assign new_D2847_ = new_D2857_ | new_D2856_;
  assign new_D2848_ = new_D2862_ & new_D2861_;
  assign new_D2849_ = new_D2860_ & new_D2859_;
  assign new_D2850_ = new_D2865_ | new_D2864_;
  assign new_D2851_ = new_D2860_ & new_D2863_;
  assign new_D2852_ = new_D2835_ | new_D2868_;
  assign new_D2853_ = new_D2867_ | new_D2866_;
  assign new_D2854_ = new_D2870_ | new_D2869_;
  assign new_D2855_ = ~new_D2846_ & new_D2872_;
  assign new_D2856_ = ~new_D2848_ & new_D2860_;
  assign new_D2857_ = new_D2848_ & ~new_D2860_;
  assign new_D2858_ = new_D2834_ & ~new_D2835_;
  assign new_D2859_ = ~new_D2881_ | ~new_D2882_;
  assign new_D2860_ = new_D2874_ | new_D2876_;
  assign new_D2861_ = new_D2884_ | new_D2883_;
  assign new_D2862_ = new_D2878_ | new_D2877_;
  assign new_D2863_ = ~new_D2886_ | ~new_D2885_;
  assign new_D2864_ = ~new_D2887_ & new_D2888_;
  assign new_D2865_ = new_D2887_ & ~new_D2888_;
  assign new_D2866_ = ~new_D2834_ & new_D2835_;
  assign new_D2867_ = new_D2834_ & ~new_D2835_;
  assign new_D2868_ = ~new_D2850_ | new_D2860_;
  assign new_D2869_ = new_D2850_ & new_D2860_;
  assign new_D2870_ = ~new_D2850_ & ~new_D2860_;
  assign new_D2871_ = new_D2892_ | new_D2891_;
  assign new_D2872_ = new_D2838_ | new_D2871_;
  assign new_D2873_ = new_D2896_ | new_D2895_;
  assign new_D2874_ = ~new_D2838_ & new_D2873_;
  assign new_D2875_ = new_D2894_ | new_D2893_;
  assign new_D2876_ = new_D2838_ & new_D2875_;
  assign new_D2877_ = new_D2836_ & ~new_D2846_;
  assign new_D2878_ = ~new_D2836_ & new_D2846_;
  assign new_D2879_ = ~new_D2835_ | ~new_D2860_;
  assign new_D2880_ = new_D2846_ & new_D2879_;
  assign new_D2881_ = ~new_D2846_ & ~new_D2880_;
  assign new_D2882_ = new_D2846_ | new_D2879_;
  assign new_D2883_ = ~new_D2836_ & new_D2837_;
  assign new_D2884_ = new_D2836_ & ~new_D2837_;
  assign new_D2885_ = new_D2853_ | new_D2890_;
  assign new_D2886_ = ~new_D2853_ & ~new_D2889_;
  assign new_D2887_ = new_D2836_ | new_D2853_;
  assign new_D2888_ = new_D2836_ | new_D2837_;
  assign new_D2889_ = new_D2853_ & new_D2890_;
  assign new_D2890_ = ~new_D2835_ | ~new_D2860_;
  assign new_D2891_ = new_D2868_ & new_D2888_;
  assign new_D2892_ = ~new_D2868_ & ~new_D2888_;
  assign new_D2893_ = new_D2897_ | new_D2898_;
  assign new_D2894_ = ~new_D2839_ & new_D2853_;
  assign new_D2895_ = new_D2899_ | new_D2900_;
  assign new_D2896_ = new_D2839_ & new_D2853_;
  assign new_D2897_ = ~new_D2839_ & ~new_D2853_;
  assign new_D2898_ = new_D2839_ & ~new_D2853_;
  assign new_D2899_ = new_D2839_ & ~new_D2853_;
  assign new_D2900_ = ~new_D2839_ & new_D2853_;
  assign new_D2901_ = new_E1421_;
  assign new_D2902_ = new_E1488_;
  assign new_D2903_ = new_E1555_;
  assign new_D2904_ = new_E1622_;
  assign new_D2905_ = new_E1689_;
  assign new_D2906_ = new_E1756_;
  assign new_D2907_ = new_D2914_ & new_D2913_;
  assign new_D2908_ = new_D2916_ | new_D2915_;
  assign new_D2909_ = new_D2918_ | new_D2917_;
  assign new_D2910_ = new_D2920_ & new_D2919_;
  assign new_D2911_ = new_D2920_ & new_D2921_;
  assign new_D2912_ = new_D2913_ | new_D2922_;
  assign new_D2913_ = new_D2902_ | new_D2925_;
  assign new_D2914_ = new_D2924_ | new_D2923_;
  assign new_D2915_ = new_D2929_ & new_D2928_;
  assign new_D2916_ = new_D2927_ & new_D2926_;
  assign new_D2917_ = new_D2932_ | new_D2931_;
  assign new_D2918_ = new_D2927_ & new_D2930_;
  assign new_D2919_ = new_D2902_ | new_D2935_;
  assign new_D2920_ = new_D2934_ | new_D2933_;
  assign new_D2921_ = new_D2937_ | new_D2936_;
  assign new_D2922_ = ~new_D2913_ & new_D2939_;
  assign new_D2923_ = ~new_D2915_ & new_D2927_;
  assign new_D2924_ = new_D2915_ & ~new_D2927_;
  assign new_D2925_ = new_D2901_ & ~new_D2902_;
  assign new_D2926_ = ~new_D2948_ | ~new_D2949_;
  assign new_D2927_ = new_D2941_ | new_D2943_;
  assign new_D2928_ = new_D2951_ | new_D2950_;
  assign new_D2929_ = new_D2945_ | new_D2944_;
  assign new_D2930_ = ~new_D2953_ | ~new_D2952_;
  assign new_D2931_ = ~new_D2954_ & new_D2955_;
  assign new_D2932_ = new_D2954_ & ~new_D2955_;
  assign new_D2933_ = ~new_D2901_ & new_D2902_;
  assign new_D2934_ = new_D2901_ & ~new_D2902_;
  assign new_D2935_ = ~new_D2917_ | new_D2927_;
  assign new_D2936_ = new_D2917_ & new_D2927_;
  assign new_D2937_ = ~new_D2917_ & ~new_D2927_;
  assign new_D2938_ = new_D2959_ | new_D2958_;
  assign new_D2939_ = new_D2905_ | new_D2938_;
  assign new_D2940_ = new_D2963_ | new_D2962_;
  assign new_D2941_ = ~new_D2905_ & new_D2940_;
  assign new_D2942_ = new_D2961_ | new_D2960_;
  assign new_D2943_ = new_D2905_ & new_D2942_;
  assign new_D2944_ = new_D2903_ & ~new_D2913_;
  assign new_D2945_ = ~new_D2903_ & new_D2913_;
  assign new_D2946_ = ~new_D2902_ | ~new_D2927_;
  assign new_D2947_ = new_D2913_ & new_D2946_;
  assign new_D2948_ = ~new_D2913_ & ~new_D2947_;
  assign new_D2949_ = new_D2913_ | new_D2946_;
  assign new_D2950_ = ~new_D2903_ & new_D2904_;
  assign new_D2951_ = new_D2903_ & ~new_D2904_;
  assign new_D2952_ = new_D2920_ | new_D2957_;
  assign new_D2953_ = ~new_D2920_ & ~new_D2956_;
  assign new_D2954_ = new_D2903_ | new_D2920_;
  assign new_D2955_ = new_D2903_ | new_D2904_;
  assign new_D2956_ = new_D2920_ & new_D2957_;
  assign new_D2957_ = ~new_D2902_ | ~new_D2927_;
  assign new_D2958_ = new_D2935_ & new_D2955_;
  assign new_D2959_ = ~new_D2935_ & ~new_D2955_;
  assign new_D2960_ = new_D2964_ | new_D2965_;
  assign new_D2961_ = ~new_D2906_ & new_D2920_;
  assign new_D2962_ = new_D2966_ | new_D2967_;
  assign new_D2963_ = new_D2906_ & new_D2920_;
  assign new_D2964_ = ~new_D2906_ & ~new_D2920_;
  assign new_D2965_ = new_D2906_ & ~new_D2920_;
  assign new_D2966_ = new_D2906_ & ~new_D2920_;
  assign new_D2967_ = ~new_D2906_ & new_D2920_;
  assign new_D2968_ = new_E1823_;
  assign new_D2969_ = new_E1890_;
  assign new_D2970_ = new_E1957_;
  assign new_D2971_ = new_E2024_;
  assign new_D2972_ = new_E2091_;
  assign new_D2973_ = new_E2158_;
  assign new_D2974_ = new_D2981_ & new_D2980_;
  assign new_D2975_ = new_D2983_ | new_D2982_;
  assign new_D2976_ = new_D2985_ | new_D2984_;
  assign new_D2977_ = new_D2987_ & new_D2986_;
  assign new_D2978_ = new_D2987_ & new_D2988_;
  assign new_D2979_ = new_D2980_ | new_D2989_;
  assign new_D2980_ = new_D2969_ | new_D2992_;
  assign new_D2981_ = new_D2991_ | new_D2990_;
  assign new_D2982_ = new_D2996_ & new_D2995_;
  assign new_D2983_ = new_D2994_ & new_D2993_;
  assign new_D2984_ = new_D2999_ | new_D2998_;
  assign new_D2985_ = new_D2994_ & new_D2997_;
  assign new_D2986_ = new_D2969_ | new_D3002_;
  assign new_D2987_ = new_D3001_ | new_D3000_;
  assign new_D2988_ = new_D3004_ | new_D3003_;
  assign new_D2989_ = ~new_D2980_ & new_D3006_;
  assign new_D2990_ = ~new_D2982_ & new_D2994_;
  assign new_D2991_ = new_D2982_ & ~new_D2994_;
  assign new_D2992_ = new_D2968_ & ~new_D2969_;
  assign new_D2993_ = ~new_D3015_ | ~new_D3016_;
  assign new_D2994_ = new_D3008_ | new_D3010_;
  assign new_D2995_ = new_D3018_ | new_D3017_;
  assign new_D2996_ = new_D3012_ | new_D3011_;
  assign new_D2997_ = ~new_D3020_ | ~new_D3019_;
  assign new_D2998_ = ~new_D3021_ & new_D3022_;
  assign new_D2999_ = new_D3021_ & ~new_D3022_;
  assign new_D3000_ = ~new_D2968_ & new_D2969_;
  assign new_D3001_ = new_D2968_ & ~new_D2969_;
  assign new_D3002_ = ~new_D2984_ | new_D2994_;
  assign new_D3003_ = new_D2984_ & new_D2994_;
  assign new_D3004_ = ~new_D2984_ & ~new_D2994_;
  assign new_D3005_ = new_D3026_ | new_D3025_;
  assign new_D3006_ = new_D2972_ | new_D3005_;
  assign new_D3007_ = new_D3030_ | new_D3029_;
  assign new_D3008_ = ~new_D2972_ & new_D3007_;
  assign new_D3009_ = new_D3028_ | new_D3027_;
  assign new_D3010_ = new_D2972_ & new_D3009_;
  assign new_D3011_ = new_D2970_ & ~new_D2980_;
  assign new_D3012_ = ~new_D2970_ & new_D2980_;
  assign new_D3013_ = ~new_D2969_ | ~new_D2994_;
  assign new_D3014_ = new_D2980_ & new_D3013_;
  assign new_D3015_ = ~new_D2980_ & ~new_D3014_;
  assign new_D3016_ = new_D2980_ | new_D3013_;
  assign new_D3017_ = ~new_D2970_ & new_D2971_;
  assign new_D3018_ = new_D2970_ & ~new_D2971_;
  assign new_D3019_ = new_D2987_ | new_D3024_;
  assign new_D3020_ = ~new_D2987_ & ~new_D3023_;
  assign new_D3021_ = new_D2970_ | new_D2987_;
  assign new_D3022_ = new_D2970_ | new_D2971_;
  assign new_D3023_ = new_D2987_ & new_D3024_;
  assign new_D3024_ = ~new_D2969_ | ~new_D2994_;
  assign new_D3025_ = new_D3002_ & new_D3022_;
  assign new_D3026_ = ~new_D3002_ & ~new_D3022_;
  assign new_D3027_ = new_D3031_ | new_D3032_;
  assign new_D3028_ = ~new_D2973_ & new_D2987_;
  assign new_D3029_ = new_D3033_ | new_D3034_;
  assign new_D3030_ = new_D2973_ & new_D2987_;
  assign new_D3031_ = ~new_D2973_ & ~new_D2987_;
  assign new_D3032_ = new_D2973_ & ~new_D2987_;
  assign new_D3033_ = new_D2973_ & ~new_D2987_;
  assign new_D3034_ = ~new_D2973_ & new_D2987_;
  assign new_D3035_ = new_E2225_;
  assign new_D3036_ = new_E2292_;
  assign new_D3037_ = new_E2359_;
  assign new_D3038_ = new_E2426_;
  assign new_D3039_ = new_E2493_;
  assign new_D3040_ = new_E2560_;
  assign new_D3041_ = new_D3048_ & new_D3047_;
  assign new_D3042_ = new_D3050_ | new_D3049_;
  assign new_D3043_ = new_D3052_ | new_D3051_;
  assign new_D3044_ = new_D3054_ & new_D3053_;
  assign new_D3045_ = new_D3054_ & new_D3055_;
  assign new_D3046_ = new_D3047_ | new_D3056_;
  assign new_D3047_ = new_D3036_ | new_D3059_;
  assign new_D3048_ = new_D3058_ | new_D3057_;
  assign new_D3049_ = new_D3063_ & new_D3062_;
  assign new_D3050_ = new_D3061_ & new_D3060_;
  assign new_D3051_ = new_D3066_ | new_D3065_;
  assign new_D3052_ = new_D3061_ & new_D3064_;
  assign new_D3053_ = new_D3036_ | new_D3069_;
  assign new_D3054_ = new_D3068_ | new_D3067_;
  assign new_D3055_ = new_D3071_ | new_D3070_;
  assign new_D3056_ = ~new_D3047_ & new_D3073_;
  assign new_D3057_ = ~new_D3049_ & new_D3061_;
  assign new_D3058_ = new_D3049_ & ~new_D3061_;
  assign new_D3059_ = new_D3035_ & ~new_D3036_;
  assign new_D3060_ = ~new_D3082_ | ~new_D3083_;
  assign new_D3061_ = new_D3075_ | new_D3077_;
  assign new_D3062_ = new_D3085_ | new_D3084_;
  assign new_D3063_ = new_D3079_ | new_D3078_;
  assign new_D3064_ = ~new_D3087_ | ~new_D3086_;
  assign new_D3065_ = ~new_D3088_ & new_D3089_;
  assign new_D3066_ = new_D3088_ & ~new_D3089_;
  assign new_D3067_ = ~new_D3035_ & new_D3036_;
  assign new_D3068_ = new_D3035_ & ~new_D3036_;
  assign new_D3069_ = ~new_D3051_ | new_D3061_;
  assign new_D3070_ = new_D3051_ & new_D3061_;
  assign new_D3071_ = ~new_D3051_ & ~new_D3061_;
  assign new_D3072_ = new_D3093_ | new_D3092_;
  assign new_D3073_ = new_D3039_ | new_D3072_;
  assign new_D3074_ = new_D3097_ | new_D3096_;
  assign new_D3075_ = ~new_D3039_ & new_D3074_;
  assign new_D3076_ = new_D3095_ | new_D3094_;
  assign new_D3077_ = new_D3039_ & new_D3076_;
  assign new_D3078_ = new_D3037_ & ~new_D3047_;
  assign new_D3079_ = ~new_D3037_ & new_D3047_;
  assign new_D3080_ = ~new_D3036_ | ~new_D3061_;
  assign new_D3081_ = new_D3047_ & new_D3080_;
  assign new_D3082_ = ~new_D3047_ & ~new_D3081_;
  assign new_D3083_ = new_D3047_ | new_D3080_;
  assign new_D3084_ = ~new_D3037_ & new_D3038_;
  assign new_D3085_ = new_D3037_ & ~new_D3038_;
  assign new_D3086_ = new_D3054_ | new_D3091_;
  assign new_D3087_ = ~new_D3054_ & ~new_D3090_;
  assign new_D3088_ = new_D3037_ | new_D3054_;
  assign new_D3089_ = new_D3037_ | new_D3038_;
  assign new_D3090_ = new_D3054_ & new_D3091_;
  assign new_D3091_ = ~new_D3036_ | ~new_D3061_;
  assign new_D3092_ = new_D3069_ & new_D3089_;
  assign new_D3093_ = ~new_D3069_ & ~new_D3089_;
  assign new_D3094_ = new_D3098_ | new_D3099_;
  assign new_D3095_ = ~new_D3040_ & new_D3054_;
  assign new_D3096_ = new_D3100_ | new_D3101_;
  assign new_D3097_ = new_D3040_ & new_D3054_;
  assign new_D3098_ = ~new_D3040_ & ~new_D3054_;
  assign new_D3099_ = new_D3040_ & ~new_D3054_;
  assign new_D3100_ = new_D3040_ & ~new_D3054_;
  assign new_D3101_ = ~new_D3040_ & new_D3054_;
  assign new_D3102_ = new_E2627_;
  assign new_D3103_ = new_E2694_;
  assign new_D3104_ = new_E2761_;
  assign new_D3105_ = new_E2828_;
  assign new_D3106_ = new_E2895_;
  assign new_D3107_ = new_E2962_;
  assign new_D3108_ = new_D3115_ & new_D3114_;
  assign new_D3109_ = new_D3117_ | new_D3116_;
  assign new_D3110_ = new_D3119_ | new_D3118_;
  assign new_D3111_ = new_D3121_ & new_D3120_;
  assign new_D3112_ = new_D3121_ & new_D3122_;
  assign new_D3113_ = new_D3114_ | new_D3123_;
  assign new_D3114_ = new_D3103_ | new_D3126_;
  assign new_D3115_ = new_D3125_ | new_D3124_;
  assign new_D3116_ = new_D3130_ & new_D3129_;
  assign new_D3117_ = new_D3128_ & new_D3127_;
  assign new_D3118_ = new_D3133_ | new_D3132_;
  assign new_D3119_ = new_D3128_ & new_D3131_;
  assign new_D3120_ = new_D3103_ | new_D3136_;
  assign new_D3121_ = new_D3135_ | new_D3134_;
  assign new_D3122_ = new_D3138_ | new_D3137_;
  assign new_D3123_ = ~new_D3114_ & new_D3140_;
  assign new_D3124_ = ~new_D3116_ & new_D3128_;
  assign new_D3125_ = new_D3116_ & ~new_D3128_;
  assign new_D3126_ = new_D3102_ & ~new_D3103_;
  assign new_D3127_ = ~new_D3149_ | ~new_D3150_;
  assign new_D3128_ = new_D3142_ | new_D3144_;
  assign new_D3129_ = new_D3152_ | new_D3151_;
  assign new_D3130_ = new_D3146_ | new_D3145_;
  assign new_D3131_ = ~new_D3154_ | ~new_D3153_;
  assign new_D3132_ = ~new_D3155_ & new_D3156_;
  assign new_D3133_ = new_D3155_ & ~new_D3156_;
  assign new_D3134_ = ~new_D3102_ & new_D3103_;
  assign new_D3135_ = new_D3102_ & ~new_D3103_;
  assign new_D3136_ = ~new_D3118_ | new_D3128_;
  assign new_D3137_ = new_D3118_ & new_D3128_;
  assign new_D3138_ = ~new_D3118_ & ~new_D3128_;
  assign new_D3139_ = new_D3160_ | new_D3159_;
  assign new_D3140_ = new_D3106_ | new_D3139_;
  assign new_D3141_ = new_D3164_ | new_D3163_;
  assign new_D3142_ = ~new_D3106_ & new_D3141_;
  assign new_D3143_ = new_D3162_ | new_D3161_;
  assign new_D3144_ = new_D3106_ & new_D3143_;
  assign new_D3145_ = new_D3104_ & ~new_D3114_;
  assign new_D3146_ = ~new_D3104_ & new_D3114_;
  assign new_D3147_ = ~new_D3103_ | ~new_D3128_;
  assign new_D3148_ = new_D3114_ & new_D3147_;
  assign new_D3149_ = ~new_D3114_ & ~new_D3148_;
  assign new_D3150_ = new_D3114_ | new_D3147_;
  assign new_D3151_ = ~new_D3104_ & new_D3105_;
  assign new_D3152_ = new_D3104_ & ~new_D3105_;
  assign new_D3153_ = new_D3121_ | new_D3158_;
  assign new_D3154_ = ~new_D3121_ & ~new_D3157_;
  assign new_D3155_ = new_D3104_ | new_D3121_;
  assign new_D3156_ = new_D3104_ | new_D3105_;
  assign new_D3157_ = new_D3121_ & new_D3158_;
  assign new_D3158_ = ~new_D3103_ | ~new_D3128_;
  assign new_D3159_ = new_D3136_ & new_D3156_;
  assign new_D3160_ = ~new_D3136_ & ~new_D3156_;
  assign new_D3161_ = new_D3165_ | new_D3166_;
  assign new_D3162_ = ~new_D3107_ & new_D3121_;
  assign new_D3163_ = new_D3167_ | new_D3168_;
  assign new_D3164_ = new_D3107_ & new_D3121_;
  assign new_D3165_ = ~new_D3107_ & ~new_D3121_;
  assign new_D3166_ = new_D3107_ & ~new_D3121_;
  assign new_D3167_ = new_D3107_ & ~new_D3121_;
  assign new_D3168_ = ~new_D3107_ & new_D3121_;
  assign new_D3169_ = new_E3029_;
  assign new_D3170_ = new_E3096_;
  assign new_D3171_ = new_E3163_;
  assign new_D3172_ = new_E3230_;
  assign new_D3173_ = new_E3297_;
  assign new_D3174_ = new_E3364_;
  assign new_D3175_ = new_D3182_ & new_D3181_;
  assign new_D3176_ = new_D3184_ | new_D3183_;
  assign new_D3177_ = new_D3186_ | new_D3185_;
  assign new_D3178_ = new_D3188_ & new_D3187_;
  assign new_D3179_ = new_D3188_ & new_D3189_;
  assign new_D3180_ = new_D3181_ | new_D3190_;
  assign new_D3181_ = new_D3170_ | new_D3193_;
  assign new_D3182_ = new_D3192_ | new_D3191_;
  assign new_D3183_ = new_D3197_ & new_D3196_;
  assign new_D3184_ = new_D3195_ & new_D3194_;
  assign new_D3185_ = new_D3200_ | new_D3199_;
  assign new_D3186_ = new_D3195_ & new_D3198_;
  assign new_D3187_ = new_D3170_ | new_D3203_;
  assign new_D3188_ = new_D3202_ | new_D3201_;
  assign new_D3189_ = new_D3205_ | new_D3204_;
  assign new_D3190_ = ~new_D3181_ & new_D3207_;
  assign new_D3191_ = ~new_D3183_ & new_D3195_;
  assign new_D3192_ = new_D3183_ & ~new_D3195_;
  assign new_D3193_ = new_D3169_ & ~new_D3170_;
  assign new_D3194_ = ~new_D3216_ | ~new_D3217_;
  assign new_D3195_ = new_D3209_ | new_D3211_;
  assign new_D3196_ = new_D3219_ | new_D3218_;
  assign new_D3197_ = new_D3213_ | new_D3212_;
  assign new_D3198_ = ~new_D3221_ | ~new_D3220_;
  assign new_D3199_ = ~new_D3222_ & new_D3223_;
  assign new_D3200_ = new_D3222_ & ~new_D3223_;
  assign new_D3201_ = ~new_D3169_ & new_D3170_;
  assign new_D3202_ = new_D3169_ & ~new_D3170_;
  assign new_D3203_ = ~new_D3185_ | new_D3195_;
  assign new_D3204_ = new_D3185_ & new_D3195_;
  assign new_D3205_ = ~new_D3185_ & ~new_D3195_;
  assign new_D3206_ = new_D3227_ | new_D3226_;
  assign new_D3207_ = new_D3173_ | new_D3206_;
  assign new_D3208_ = new_D3231_ | new_D3230_;
  assign new_D3209_ = ~new_D3173_ & new_D3208_;
  assign new_D3210_ = new_D3229_ | new_D3228_;
  assign new_D3211_ = new_D3173_ & new_D3210_;
  assign new_D3212_ = new_D3171_ & ~new_D3181_;
  assign new_D3213_ = ~new_D3171_ & new_D3181_;
  assign new_D3214_ = ~new_D3170_ | ~new_D3195_;
  assign new_D3215_ = new_D3181_ & new_D3214_;
  assign new_D3216_ = ~new_D3181_ & ~new_D3215_;
  assign new_D3217_ = new_D3181_ | new_D3214_;
  assign new_D3218_ = ~new_D3171_ & new_D3172_;
  assign new_D3219_ = new_D3171_ & ~new_D3172_;
  assign new_D3220_ = new_D3188_ | new_D3225_;
  assign new_D3221_ = ~new_D3188_ & ~new_D3224_;
  assign new_D3222_ = new_D3171_ | new_D3188_;
  assign new_D3223_ = new_D3171_ | new_D3172_;
  assign new_D3224_ = new_D3188_ & new_D3225_;
  assign new_D3225_ = ~new_D3170_ | ~new_D3195_;
  assign new_D3226_ = new_D3203_ & new_D3223_;
  assign new_D3227_ = ~new_D3203_ & ~new_D3223_;
  assign new_D3228_ = new_D3232_ | new_D3233_;
  assign new_D3229_ = ~new_D3174_ & new_D3188_;
  assign new_D3230_ = new_D3234_ | new_D3235_;
  assign new_D3231_ = new_D3174_ & new_D3188_;
  assign new_D3232_ = ~new_D3174_ & ~new_D3188_;
  assign new_D3233_ = new_D3174_ & ~new_D3188_;
  assign new_D3234_ = new_D3174_ & ~new_D3188_;
  assign new_D3235_ = ~new_D3174_ & new_D3188_;
  assign new_D3236_ = new_E3431_;
  assign new_D3237_ = new_E3498_;
  assign new_D3238_ = new_E3565_;
  assign new_D3239_ = new_E3632_;
  assign new_D3240_ = new_E3699_;
  assign new_D3241_ = new_E3766_;
  assign new_D3242_ = new_D3249_ & new_D3248_;
  assign new_D3243_ = new_D3251_ | new_D3250_;
  assign new_D3244_ = new_D3253_ | new_D3252_;
  assign new_D3245_ = new_D3255_ & new_D3254_;
  assign new_D3246_ = new_D3255_ & new_D3256_;
  assign new_D3247_ = new_D3248_ | new_D3257_;
  assign new_D3248_ = new_D3237_ | new_D3260_;
  assign new_D3249_ = new_D3259_ | new_D3258_;
  assign new_D3250_ = new_D3264_ & new_D3263_;
  assign new_D3251_ = new_D3262_ & new_D3261_;
  assign new_D3252_ = new_D3267_ | new_D3266_;
  assign new_D3253_ = new_D3262_ & new_D3265_;
  assign new_D3254_ = new_D3237_ | new_D3270_;
  assign new_D3255_ = new_D3269_ | new_D3268_;
  assign new_D3256_ = new_D3272_ | new_D3271_;
  assign new_D3257_ = ~new_D3248_ & new_D3274_;
  assign new_D3258_ = ~new_D3250_ & new_D3262_;
  assign new_D3259_ = new_D3250_ & ~new_D3262_;
  assign new_D3260_ = new_D3236_ & ~new_D3237_;
  assign new_D3261_ = ~new_D3283_ | ~new_D3284_;
  assign new_D3262_ = new_D3276_ | new_D3278_;
  assign new_D3263_ = new_D3286_ | new_D3285_;
  assign new_D3264_ = new_D3280_ | new_D3279_;
  assign new_D3265_ = ~new_D3288_ | ~new_D3287_;
  assign new_D3266_ = ~new_D3289_ & new_D3290_;
  assign new_D3267_ = new_D3289_ & ~new_D3290_;
  assign new_D3268_ = ~new_D3236_ & new_D3237_;
  assign new_D3269_ = new_D3236_ & ~new_D3237_;
  assign new_D3270_ = ~new_D3252_ | new_D3262_;
  assign new_D3271_ = new_D3252_ & new_D3262_;
  assign new_D3272_ = ~new_D3252_ & ~new_D3262_;
  assign new_D3273_ = new_D3294_ | new_D3293_;
  assign new_D3274_ = new_D3240_ | new_D3273_;
  assign new_D3275_ = new_D3298_ | new_D3297_;
  assign new_D3276_ = ~new_D3240_ & new_D3275_;
  assign new_D3277_ = new_D3296_ | new_D3295_;
  assign new_D3278_ = new_D3240_ & new_D3277_;
  assign new_D3279_ = new_D3238_ & ~new_D3248_;
  assign new_D3280_ = ~new_D3238_ & new_D3248_;
  assign new_D3281_ = ~new_D3237_ | ~new_D3262_;
  assign new_D3282_ = new_D3248_ & new_D3281_;
  assign new_D3283_ = ~new_D3248_ & ~new_D3282_;
  assign new_D3284_ = new_D3248_ | new_D3281_;
  assign new_D3285_ = ~new_D3238_ & new_D3239_;
  assign new_D3286_ = new_D3238_ & ~new_D3239_;
  assign new_D3287_ = new_D3255_ | new_D3292_;
  assign new_D3288_ = ~new_D3255_ & ~new_D3291_;
  assign new_D3289_ = new_D3238_ | new_D3255_;
  assign new_D3290_ = new_D3238_ | new_D3239_;
  assign new_D3291_ = new_D3255_ & new_D3292_;
  assign new_D3292_ = ~new_D3237_ | ~new_D3262_;
  assign new_D3293_ = new_D3270_ & new_D3290_;
  assign new_D3294_ = ~new_D3270_ & ~new_D3290_;
  assign new_D3295_ = new_D3299_ | new_D3300_;
  assign new_D3296_ = ~new_D3241_ & new_D3255_;
  assign new_D3297_ = new_D3301_ | new_D3302_;
  assign new_D3298_ = new_D3241_ & new_D3255_;
  assign new_D3299_ = ~new_D3241_ & ~new_D3255_;
  assign new_D3300_ = new_D3241_ & ~new_D3255_;
  assign new_D3301_ = new_D3241_ & ~new_D3255_;
  assign new_D3302_ = ~new_D3241_ & new_D3255_;
  assign new_D3303_ = new_E3833_;
  assign new_D3304_ = new_E3900_;
  assign new_D3305_ = new_E3967_;
  assign new_D3306_ = new_E4034_;
  assign new_D3307_ = new_E4101_;
  assign new_D3308_ = new_E4168_;
  assign new_D3309_ = new_D3316_ & new_D3315_;
  assign new_D3310_ = new_D3318_ | new_D3317_;
  assign new_D3311_ = new_D3320_ | new_D3319_;
  assign new_D3312_ = new_D3322_ & new_D3321_;
  assign new_D3313_ = new_D3322_ & new_D3323_;
  assign new_D3314_ = new_D3315_ | new_D3324_;
  assign new_D3315_ = new_D3304_ | new_D3327_;
  assign new_D3316_ = new_D3326_ | new_D3325_;
  assign new_D3317_ = new_D3331_ & new_D3330_;
  assign new_D3318_ = new_D3329_ & new_D3328_;
  assign new_D3319_ = new_D3334_ | new_D3333_;
  assign new_D3320_ = new_D3329_ & new_D3332_;
  assign new_D3321_ = new_D3304_ | new_D3337_;
  assign new_D3322_ = new_D3336_ | new_D3335_;
  assign new_D3323_ = new_D3339_ | new_D3338_;
  assign new_D3324_ = ~new_D3315_ & new_D3341_;
  assign new_D3325_ = ~new_D3317_ & new_D3329_;
  assign new_D3326_ = new_D3317_ & ~new_D3329_;
  assign new_D3327_ = new_D3303_ & ~new_D3304_;
  assign new_D3328_ = ~new_D3350_ | ~new_D3351_;
  assign new_D3329_ = new_D3343_ | new_D3345_;
  assign new_D3330_ = new_D3353_ | new_D3352_;
  assign new_D3331_ = new_D3347_ | new_D3346_;
  assign new_D3332_ = ~new_D3355_ | ~new_D3354_;
  assign new_D3333_ = ~new_D3356_ & new_D3357_;
  assign new_D3334_ = new_D3356_ & ~new_D3357_;
  assign new_D3335_ = ~new_D3303_ & new_D3304_;
  assign new_D3336_ = new_D3303_ & ~new_D3304_;
  assign new_D3337_ = ~new_D3319_ | new_D3329_;
  assign new_D3338_ = new_D3319_ & new_D3329_;
  assign new_D3339_ = ~new_D3319_ & ~new_D3329_;
  assign new_D3340_ = new_D3361_ | new_D3360_;
  assign new_D3341_ = new_D3307_ | new_D3340_;
  assign new_D3342_ = new_D3365_ | new_D3364_;
  assign new_D3343_ = ~new_D3307_ & new_D3342_;
  assign new_D3344_ = new_D3363_ | new_D3362_;
  assign new_D3345_ = new_D3307_ & new_D3344_;
  assign new_D3346_ = new_D3305_ & ~new_D3315_;
  assign new_D3347_ = ~new_D3305_ & new_D3315_;
  assign new_D3348_ = ~new_D3304_ | ~new_D3329_;
  assign new_D3349_ = new_D3315_ & new_D3348_;
  assign new_D3350_ = ~new_D3315_ & ~new_D3349_;
  assign new_D3351_ = new_D3315_ | new_D3348_;
  assign new_D3352_ = ~new_D3305_ & new_D3306_;
  assign new_D3353_ = new_D3305_ & ~new_D3306_;
  assign new_D3354_ = new_D3322_ | new_D3359_;
  assign new_D3355_ = ~new_D3322_ & ~new_D3358_;
  assign new_D3356_ = new_D3305_ | new_D3322_;
  assign new_D3357_ = new_D3305_ | new_D3306_;
  assign new_D3358_ = new_D3322_ & new_D3359_;
  assign new_D3359_ = ~new_D3304_ | ~new_D3329_;
  assign new_D3360_ = new_D3337_ & new_D3357_;
  assign new_D3361_ = ~new_D3337_ & ~new_D3357_;
  assign new_D3362_ = new_D3366_ | new_D3367_;
  assign new_D3363_ = ~new_D3308_ & new_D3322_;
  assign new_D3364_ = new_D3368_ | new_D3369_;
  assign new_D3365_ = new_D3308_ & new_D3322_;
  assign new_D3366_ = ~new_D3308_ & ~new_D3322_;
  assign new_D3367_ = new_D3308_ & ~new_D3322_;
  assign new_D3368_ = new_D3308_ & ~new_D3322_;
  assign new_D3369_ = ~new_D3308_ & new_D3322_;
  assign new_D3370_ = new_E4235_;
  assign new_D3371_ = new_E4302_;
  assign new_D3372_ = new_E4369_;
  assign new_D3373_ = new_E4436_;
  assign new_D3374_ = new_E4503_;
  assign new_D3375_ = new_E4570_;
  assign new_D3376_ = new_D3383_ & new_D3382_;
  assign new_D3377_ = new_D3385_ | new_D3384_;
  assign new_D3378_ = new_D3387_ | new_D3386_;
  assign new_D3379_ = new_D3389_ & new_D3388_;
  assign new_D3380_ = new_D3389_ & new_D3390_;
  assign new_D3381_ = new_D3382_ | new_D3391_;
  assign new_D3382_ = new_D3371_ | new_D3394_;
  assign new_D3383_ = new_D3393_ | new_D3392_;
  assign new_D3384_ = new_D3398_ & new_D3397_;
  assign new_D3385_ = new_D3396_ & new_D3395_;
  assign new_D3386_ = new_D3401_ | new_D3400_;
  assign new_D3387_ = new_D3396_ & new_D3399_;
  assign new_D3388_ = new_D3371_ | new_D3404_;
  assign new_D3389_ = new_D3403_ | new_D3402_;
  assign new_D3390_ = new_D3406_ | new_D3405_;
  assign new_D3391_ = ~new_D3382_ & new_D3408_;
  assign new_D3392_ = ~new_D3384_ & new_D3396_;
  assign new_D3393_ = new_D3384_ & ~new_D3396_;
  assign new_D3394_ = new_D3370_ & ~new_D3371_;
  assign new_D3395_ = ~new_D3417_ | ~new_D3418_;
  assign new_D3396_ = new_D3410_ | new_D3412_;
  assign new_D3397_ = new_D3420_ | new_D3419_;
  assign new_D3398_ = new_D3414_ | new_D3413_;
  assign new_D3399_ = ~new_D3422_ | ~new_D3421_;
  assign new_D3400_ = ~new_D3423_ & new_D3424_;
  assign new_D3401_ = new_D3423_ & ~new_D3424_;
  assign new_D3402_ = ~new_D3370_ & new_D3371_;
  assign new_D3403_ = new_D3370_ & ~new_D3371_;
  assign new_D3404_ = ~new_D3386_ | new_D3396_;
  assign new_D3405_ = new_D3386_ & new_D3396_;
  assign new_D3406_ = ~new_D3386_ & ~new_D3396_;
  assign new_D3407_ = new_D3428_ | new_D3427_;
  assign new_D3408_ = new_D3374_ | new_D3407_;
  assign new_D3409_ = new_D3432_ | new_D3431_;
  assign new_D3410_ = ~new_D3374_ & new_D3409_;
  assign new_D3411_ = new_D3430_ | new_D3429_;
  assign new_D3412_ = new_D3374_ & new_D3411_;
  assign new_D3413_ = new_D3372_ & ~new_D3382_;
  assign new_D3414_ = ~new_D3372_ & new_D3382_;
  assign new_D3415_ = ~new_D3371_ | ~new_D3396_;
  assign new_D3416_ = new_D3382_ & new_D3415_;
  assign new_D3417_ = ~new_D3382_ & ~new_D3416_;
  assign new_D3418_ = new_D3382_ | new_D3415_;
  assign new_D3419_ = ~new_D3372_ & new_D3373_;
  assign new_D3420_ = new_D3372_ & ~new_D3373_;
  assign new_D3421_ = new_D3389_ | new_D3426_;
  assign new_D3422_ = ~new_D3389_ & ~new_D3425_;
  assign new_D3423_ = new_D3372_ | new_D3389_;
  assign new_D3424_ = new_D3372_ | new_D3373_;
  assign new_D3425_ = new_D3389_ & new_D3426_;
  assign new_D3426_ = ~new_D3371_ | ~new_D3396_;
  assign new_D3427_ = new_D3404_ & new_D3424_;
  assign new_D3428_ = ~new_D3404_ & ~new_D3424_;
  assign new_D3429_ = new_D3433_ | new_D3434_;
  assign new_D3430_ = ~new_D3375_ & new_D3389_;
  assign new_D3431_ = new_D3435_ | new_D3436_;
  assign new_D3432_ = new_D3375_ & new_D3389_;
  assign new_D3433_ = ~new_D3375_ & ~new_D3389_;
  assign new_D3434_ = new_D3375_ & ~new_D3389_;
  assign new_D3435_ = new_D3375_ & ~new_D3389_;
  assign new_D3436_ = ~new_D3375_ & new_D3389_;
  assign new_D3437_ = new_E4637_;
  assign new_D3438_ = new_E4704_;
  assign new_D3439_ = new_E4771_;
  assign new_D3440_ = new_E4838_;
  assign new_D3441_ = new_E4905_;
  assign new_D3442_ = new_E4972_;
  assign new_D3443_ = new_D3450_ & new_D3449_;
  assign new_D3444_ = new_D3452_ | new_D3451_;
  assign new_D3445_ = new_D3454_ | new_D3453_;
  assign new_D3446_ = new_D3456_ & new_D3455_;
  assign new_D3447_ = new_D3456_ & new_D3457_;
  assign new_D3448_ = new_D3449_ | new_D3458_;
  assign new_D3449_ = new_D3438_ | new_D3461_;
  assign new_D3450_ = new_D3460_ | new_D3459_;
  assign new_D3451_ = new_D3465_ & new_D3464_;
  assign new_D3452_ = new_D3463_ & new_D3462_;
  assign new_D3453_ = new_D3468_ | new_D3467_;
  assign new_D3454_ = new_D3463_ & new_D3466_;
  assign new_D3455_ = new_D3438_ | new_D3471_;
  assign new_D3456_ = new_D3470_ | new_D3469_;
  assign new_D3457_ = new_D3473_ | new_D3472_;
  assign new_D3458_ = ~new_D3449_ & new_D3475_;
  assign new_D3459_ = ~new_D3451_ & new_D3463_;
  assign new_D3460_ = new_D3451_ & ~new_D3463_;
  assign new_D3461_ = new_D3437_ & ~new_D3438_;
  assign new_D3462_ = ~new_D3484_ | ~new_D3485_;
  assign new_D3463_ = new_D3477_ | new_D3479_;
  assign new_D3464_ = new_D3487_ | new_D3486_;
  assign new_D3465_ = new_D3481_ | new_D3480_;
  assign new_D3466_ = ~new_D3489_ | ~new_D3488_;
  assign new_D3467_ = ~new_D3490_ & new_D3491_;
  assign new_D3468_ = new_D3490_ & ~new_D3491_;
  assign new_D3469_ = ~new_D3437_ & new_D3438_;
  assign new_D3470_ = new_D3437_ & ~new_D3438_;
  assign new_D3471_ = ~new_D3453_ | new_D3463_;
  assign new_D3472_ = new_D3453_ & new_D3463_;
  assign new_D3473_ = ~new_D3453_ & ~new_D3463_;
  assign new_D3474_ = new_D3495_ | new_D3494_;
  assign new_D3475_ = new_D3441_ | new_D3474_;
  assign new_D3476_ = new_D3499_ | new_D3498_;
  assign new_D3477_ = ~new_D3441_ & new_D3476_;
  assign new_D3478_ = new_D3497_ | new_D3496_;
  assign new_D3479_ = new_D3441_ & new_D3478_;
  assign new_D3480_ = new_D3439_ & ~new_D3449_;
  assign new_D3481_ = ~new_D3439_ & new_D3449_;
  assign new_D3482_ = ~new_D3438_ | ~new_D3463_;
  assign new_D3483_ = new_D3449_ & new_D3482_;
  assign new_D3484_ = ~new_D3449_ & ~new_D3483_;
  assign new_D3485_ = new_D3449_ | new_D3482_;
  assign new_D3486_ = ~new_D3439_ & new_D3440_;
  assign new_D3487_ = new_D3439_ & ~new_D3440_;
  assign new_D3488_ = new_D3456_ | new_D3493_;
  assign new_D3489_ = ~new_D3456_ & ~new_D3492_;
  assign new_D3490_ = new_D3439_ | new_D3456_;
  assign new_D3491_ = new_D3439_ | new_D3440_;
  assign new_D3492_ = new_D3456_ & new_D3493_;
  assign new_D3493_ = ~new_D3438_ | ~new_D3463_;
  assign new_D3494_ = new_D3471_ & new_D3491_;
  assign new_D3495_ = ~new_D3471_ & ~new_D3491_;
  assign new_D3496_ = new_D3500_ | new_D3501_;
  assign new_D3497_ = ~new_D3442_ & new_D3456_;
  assign new_D3498_ = new_D3502_ | new_D3503_;
  assign new_D3499_ = new_D3442_ & new_D3456_;
  assign new_D3500_ = ~new_D3442_ & ~new_D3456_;
  assign new_D3501_ = new_D3442_ & ~new_D3456_;
  assign new_D3502_ = new_D3442_ & ~new_D3456_;
  assign new_D3503_ = ~new_D3442_ & new_D3456_;
  assign new_D3504_ = new_E5039_;
  assign new_D3505_ = new_E5106_;
  assign new_D3506_ = new_E5173_;
  assign new_D3507_ = new_E5240_;
  assign new_D3508_ = new_E5307_;
  assign new_D3509_ = new_E5374_;
  assign new_D3510_ = new_D3517_ & new_D3516_;
  assign new_D3511_ = new_D3519_ | new_D3518_;
  assign new_D3512_ = new_D3521_ | new_D3520_;
  assign new_D3513_ = new_D3523_ & new_D3522_;
  assign new_D3514_ = new_D3523_ & new_D3524_;
  assign new_D3515_ = new_D3516_ | new_D3525_;
  assign new_D3516_ = new_D3505_ | new_D3528_;
  assign new_D3517_ = new_D3527_ | new_D3526_;
  assign new_D3518_ = new_D3532_ & new_D3531_;
  assign new_D3519_ = new_D3530_ & new_D3529_;
  assign new_D3520_ = new_D3535_ | new_D3534_;
  assign new_D3521_ = new_D3530_ & new_D3533_;
  assign new_D3522_ = new_D3505_ | new_D3538_;
  assign new_D3523_ = new_D3537_ | new_D3536_;
  assign new_D3524_ = new_D3540_ | new_D3539_;
  assign new_D3525_ = ~new_D3516_ & new_D3542_;
  assign new_D3526_ = ~new_D3518_ & new_D3530_;
  assign new_D3527_ = new_D3518_ & ~new_D3530_;
  assign new_D3528_ = new_D3504_ & ~new_D3505_;
  assign new_D3529_ = ~new_D3551_ | ~new_D3552_;
  assign new_D3530_ = new_D3544_ | new_D3546_;
  assign new_D3531_ = new_D3554_ | new_D3553_;
  assign new_D3532_ = new_D3548_ | new_D3547_;
  assign new_D3533_ = ~new_D3556_ | ~new_D3555_;
  assign new_D3534_ = ~new_D3557_ & new_D3558_;
  assign new_D3535_ = new_D3557_ & ~new_D3558_;
  assign new_D3536_ = ~new_D3504_ & new_D3505_;
  assign new_D3537_ = new_D3504_ & ~new_D3505_;
  assign new_D3538_ = ~new_D3520_ | new_D3530_;
  assign new_D3539_ = new_D3520_ & new_D3530_;
  assign new_D3540_ = ~new_D3520_ & ~new_D3530_;
  assign new_D3541_ = new_D3562_ | new_D3561_;
  assign new_D3542_ = new_D3508_ | new_D3541_;
  assign new_D3543_ = new_D3566_ | new_D3565_;
  assign new_D3544_ = ~new_D3508_ & new_D3543_;
  assign new_D3545_ = new_D3564_ | new_D3563_;
  assign new_D3546_ = new_D3508_ & new_D3545_;
  assign new_D3547_ = new_D3506_ & ~new_D3516_;
  assign new_D3548_ = ~new_D3506_ & new_D3516_;
  assign new_D3549_ = ~new_D3505_ | ~new_D3530_;
  assign new_D3550_ = new_D3516_ & new_D3549_;
  assign new_D3551_ = ~new_D3516_ & ~new_D3550_;
  assign new_D3552_ = new_D3516_ | new_D3549_;
  assign new_D3553_ = ~new_D3506_ & new_D3507_;
  assign new_D3554_ = new_D3506_ & ~new_D3507_;
  assign new_D3555_ = new_D3523_ | new_D3560_;
  assign new_D3556_ = ~new_D3523_ & ~new_D3559_;
  assign new_D3557_ = new_D3506_ | new_D3523_;
  assign new_D3558_ = new_D3506_ | new_D3507_;
  assign new_D3559_ = new_D3523_ & new_D3560_;
  assign new_D3560_ = ~new_D3505_ | ~new_D3530_;
  assign new_D3561_ = new_D3538_ & new_D3558_;
  assign new_D3562_ = ~new_D3538_ & ~new_D3558_;
  assign new_D3563_ = new_D3567_ | new_D3568_;
  assign new_D3564_ = ~new_D3509_ & new_D3523_;
  assign new_D3565_ = new_D3569_ | new_D3570_;
  assign new_D3566_ = new_D3509_ & new_D3523_;
  assign new_D3567_ = ~new_D3509_ & ~new_D3523_;
  assign new_D3568_ = new_D3509_ & ~new_D3523_;
  assign new_D3569_ = new_D3509_ & ~new_D3523_;
  assign new_D3570_ = ~new_D3509_ & new_D3523_;
  assign new_D3571_ = new_E5441_;
  assign new_D3572_ = new_E5508_;
  assign new_D3573_ = new_E5575_;
  assign new_D3574_ = new_E5642_;
  assign new_D3575_ = new_E5709_;
  assign new_D3576_ = new_E5776_;
  assign new_D3577_ = new_D3584_ & new_D3583_;
  assign new_D3578_ = new_D3586_ | new_D3585_;
  assign new_D3579_ = new_D3588_ | new_D3587_;
  assign new_D3580_ = new_D3590_ & new_D3589_;
  assign new_D3581_ = new_D3590_ & new_D3591_;
  assign new_D3582_ = new_D3583_ | new_D3592_;
  assign new_D3583_ = new_D3572_ | new_D3595_;
  assign new_D3584_ = new_D3594_ | new_D3593_;
  assign new_D3585_ = new_D3599_ & new_D3598_;
  assign new_D3586_ = new_D3597_ & new_D3596_;
  assign new_D3587_ = new_D3602_ | new_D3601_;
  assign new_D3588_ = new_D3597_ & new_D3600_;
  assign new_D3589_ = new_D3572_ | new_D3605_;
  assign new_D3590_ = new_D3604_ | new_D3603_;
  assign new_D3591_ = new_D3607_ | new_D3606_;
  assign new_D3592_ = ~new_D3583_ & new_D3609_;
  assign new_D3593_ = ~new_D3585_ & new_D3597_;
  assign new_D3594_ = new_D3585_ & ~new_D3597_;
  assign new_D3595_ = new_D3571_ & ~new_D3572_;
  assign new_D3596_ = ~new_D3618_ | ~new_D3619_;
  assign new_D3597_ = new_D3611_ | new_D3613_;
  assign new_D3598_ = new_D3621_ | new_D3620_;
  assign new_D3599_ = new_D3615_ | new_D3614_;
  assign new_D3600_ = ~new_D3623_ | ~new_D3622_;
  assign new_D3601_ = ~new_D3624_ & new_D3625_;
  assign new_D3602_ = new_D3624_ & ~new_D3625_;
  assign new_D3603_ = ~new_D3571_ & new_D3572_;
  assign new_D3604_ = new_D3571_ & ~new_D3572_;
  assign new_D3605_ = ~new_D3587_ | new_D3597_;
  assign new_D3606_ = new_D3587_ & new_D3597_;
  assign new_D3607_ = ~new_D3587_ & ~new_D3597_;
  assign new_D3608_ = new_D3629_ | new_D3628_;
  assign new_D3609_ = new_D3575_ | new_D3608_;
  assign new_D3610_ = new_D3633_ | new_D3632_;
  assign new_D3611_ = ~new_D3575_ & new_D3610_;
  assign new_D3612_ = new_D3631_ | new_D3630_;
  assign new_D3613_ = new_D3575_ & new_D3612_;
  assign new_D3614_ = new_D3573_ & ~new_D3583_;
  assign new_D3615_ = ~new_D3573_ & new_D3583_;
  assign new_D3616_ = ~new_D3572_ | ~new_D3597_;
  assign new_D3617_ = new_D3583_ & new_D3616_;
  assign new_D3618_ = ~new_D3583_ & ~new_D3617_;
  assign new_D3619_ = new_D3583_ | new_D3616_;
  assign new_D3620_ = ~new_D3573_ & new_D3574_;
  assign new_D3621_ = new_D3573_ & ~new_D3574_;
  assign new_D3622_ = new_D3590_ | new_D3627_;
  assign new_D3623_ = ~new_D3590_ & ~new_D3626_;
  assign new_D3624_ = new_D3573_ | new_D3590_;
  assign new_D3625_ = new_D3573_ | new_D3574_;
  assign new_D3626_ = new_D3590_ & new_D3627_;
  assign new_D3627_ = ~new_D3572_ | ~new_D3597_;
  assign new_D3628_ = new_D3605_ & new_D3625_;
  assign new_D3629_ = ~new_D3605_ & ~new_D3625_;
  assign new_D3630_ = new_D3634_ | new_D3635_;
  assign new_D3631_ = ~new_D3576_ & new_D3590_;
  assign new_D3632_ = new_D3636_ | new_D3637_;
  assign new_D3633_ = new_D3576_ & new_D3590_;
  assign new_D3634_ = ~new_D3576_ & ~new_D3590_;
  assign new_D3635_ = new_D3576_ & ~new_D3590_;
  assign new_D3636_ = new_D3576_ & ~new_D3590_;
  assign new_D3637_ = ~new_D3576_ & new_D3590_;
  assign new_D3638_ = new_E5843_;
  assign new_D3639_ = new_E5910_;
  assign new_D3640_ = new_E5977_;
  assign new_D3641_ = new_E6044_;
  assign new_D3642_ = new_E6111_;
  assign new_D3643_ = new_E6178_;
  assign new_D3644_ = new_D3651_ & new_D3650_;
  assign new_D3645_ = new_D3653_ | new_D3652_;
  assign new_D3646_ = new_D3655_ | new_D3654_;
  assign new_D3647_ = new_D3657_ & new_D3656_;
  assign new_D3648_ = new_D3657_ & new_D3658_;
  assign new_D3649_ = new_D3650_ | new_D3659_;
  assign new_D3650_ = new_D3639_ | new_D3662_;
  assign new_D3651_ = new_D3661_ | new_D3660_;
  assign new_D3652_ = new_D3666_ & new_D3665_;
  assign new_D3653_ = new_D3664_ & new_D3663_;
  assign new_D3654_ = new_D3669_ | new_D3668_;
  assign new_D3655_ = new_D3664_ & new_D3667_;
  assign new_D3656_ = new_D3639_ | new_D3672_;
  assign new_D3657_ = new_D3671_ | new_D3670_;
  assign new_D3658_ = new_D3674_ | new_D3673_;
  assign new_D3659_ = ~new_D3650_ & new_D3676_;
  assign new_D3660_ = ~new_D3652_ & new_D3664_;
  assign new_D3661_ = new_D3652_ & ~new_D3664_;
  assign new_D3662_ = new_D3638_ & ~new_D3639_;
  assign new_D3663_ = ~new_D3685_ | ~new_D3686_;
  assign new_D3664_ = new_D3678_ | new_D3680_;
  assign new_D3665_ = new_D3688_ | new_D3687_;
  assign new_D3666_ = new_D3682_ | new_D3681_;
  assign new_D3667_ = ~new_D3690_ | ~new_D3689_;
  assign new_D3668_ = ~new_D3691_ & new_D3692_;
  assign new_D3669_ = new_D3691_ & ~new_D3692_;
  assign new_D3670_ = ~new_D3638_ & new_D3639_;
  assign new_D3671_ = new_D3638_ & ~new_D3639_;
  assign new_D3672_ = ~new_D3654_ | new_D3664_;
  assign new_D3673_ = new_D3654_ & new_D3664_;
  assign new_D3674_ = ~new_D3654_ & ~new_D3664_;
  assign new_D3675_ = new_D3696_ | new_D3695_;
  assign new_D3676_ = new_D3642_ | new_D3675_;
  assign new_D3677_ = new_D3700_ | new_D3699_;
  assign new_D3678_ = ~new_D3642_ & new_D3677_;
  assign new_D3679_ = new_D3698_ | new_D3697_;
  assign new_D3680_ = new_D3642_ & new_D3679_;
  assign new_D3681_ = new_D3640_ & ~new_D3650_;
  assign new_D3682_ = ~new_D3640_ & new_D3650_;
  assign new_D3683_ = ~new_D3639_ | ~new_D3664_;
  assign new_D3684_ = new_D3650_ & new_D3683_;
  assign new_D3685_ = ~new_D3650_ & ~new_D3684_;
  assign new_D3686_ = new_D3650_ | new_D3683_;
  assign new_D3687_ = ~new_D3640_ & new_D3641_;
  assign new_D3688_ = new_D3640_ & ~new_D3641_;
  assign new_D3689_ = new_D3657_ | new_D3694_;
  assign new_D3690_ = ~new_D3657_ & ~new_D3693_;
  assign new_D3691_ = new_D3640_ | new_D3657_;
  assign new_D3692_ = new_D3640_ | new_D3641_;
  assign new_D3693_ = new_D3657_ & new_D3694_;
  assign new_D3694_ = ~new_D3639_ | ~new_D3664_;
  assign new_D3695_ = new_D3672_ & new_D3692_;
  assign new_D3696_ = ~new_D3672_ & ~new_D3692_;
  assign new_D3697_ = new_D3701_ | new_D3702_;
  assign new_D3698_ = ~new_D3643_ & new_D3657_;
  assign new_D3699_ = new_D3703_ | new_D3704_;
  assign new_D3700_ = new_D3643_ & new_D3657_;
  assign new_D3701_ = ~new_D3643_ & ~new_D3657_;
  assign new_D3702_ = new_D3643_ & ~new_D3657_;
  assign new_D3703_ = new_D3643_ & ~new_D3657_;
  assign new_D3704_ = ~new_D3643_ & new_D3657_;
  assign new_D3705_ = new_E6245_;
  assign new_D3706_ = new_E6312_;
  assign new_D3707_ = new_E6379_;
  assign new_D3708_ = new_E6446_;
  assign new_D3709_ = new_E6513_;
  assign new_D3710_ = new_E6580_;
  assign new_D3711_ = new_D3718_ & new_D3717_;
  assign new_D3712_ = new_D3720_ | new_D3719_;
  assign new_D3713_ = new_D3722_ | new_D3721_;
  assign new_D3714_ = new_D3724_ & new_D3723_;
  assign new_D3715_ = new_D3724_ & new_D3725_;
  assign new_D3716_ = new_D3717_ | new_D3726_;
  assign new_D3717_ = new_D3706_ | new_D3729_;
  assign new_D3718_ = new_D3728_ | new_D3727_;
  assign new_D3719_ = new_D3733_ & new_D3732_;
  assign new_D3720_ = new_D3731_ & new_D3730_;
  assign new_D3721_ = new_D3736_ | new_D3735_;
  assign new_D3722_ = new_D3731_ & new_D3734_;
  assign new_D3723_ = new_D3706_ | new_D3739_;
  assign new_D3724_ = new_D3738_ | new_D3737_;
  assign new_D3725_ = new_D3741_ | new_D3740_;
  assign new_D3726_ = ~new_D3717_ & new_D3743_;
  assign new_D3727_ = ~new_D3719_ & new_D3731_;
  assign new_D3728_ = new_D3719_ & ~new_D3731_;
  assign new_D3729_ = new_D3705_ & ~new_D3706_;
  assign new_D3730_ = ~new_D3752_ | ~new_D3753_;
  assign new_D3731_ = new_D3745_ | new_D3747_;
  assign new_D3732_ = new_D3755_ | new_D3754_;
  assign new_D3733_ = new_D3749_ | new_D3748_;
  assign new_D3734_ = ~new_D3757_ | ~new_D3756_;
  assign new_D3735_ = ~new_D3758_ & new_D3759_;
  assign new_D3736_ = new_D3758_ & ~new_D3759_;
  assign new_D3737_ = ~new_D3705_ & new_D3706_;
  assign new_D3738_ = new_D3705_ & ~new_D3706_;
  assign new_D3739_ = ~new_D3721_ | new_D3731_;
  assign new_D3740_ = new_D3721_ & new_D3731_;
  assign new_D3741_ = ~new_D3721_ & ~new_D3731_;
  assign new_D3742_ = new_D3763_ | new_D3762_;
  assign new_D3743_ = new_D3709_ | new_D3742_;
  assign new_D3744_ = new_D3767_ | new_D3766_;
  assign new_D3745_ = ~new_D3709_ & new_D3744_;
  assign new_D3746_ = new_D3765_ | new_D3764_;
  assign new_D3747_ = new_D3709_ & new_D3746_;
  assign new_D3748_ = new_D3707_ & ~new_D3717_;
  assign new_D3749_ = ~new_D3707_ & new_D3717_;
  assign new_D3750_ = ~new_D3706_ | ~new_D3731_;
  assign new_D3751_ = new_D3717_ & new_D3750_;
  assign new_D3752_ = ~new_D3717_ & ~new_D3751_;
  assign new_D3753_ = new_D3717_ | new_D3750_;
  assign new_D3754_ = ~new_D3707_ & new_D3708_;
  assign new_D3755_ = new_D3707_ & ~new_D3708_;
  assign new_D3756_ = new_D3724_ | new_D3761_;
  assign new_D3757_ = ~new_D3724_ & ~new_D3760_;
  assign new_D3758_ = new_D3707_ | new_D3724_;
  assign new_D3759_ = new_D3707_ | new_D3708_;
  assign new_D3760_ = new_D3724_ & new_D3761_;
  assign new_D3761_ = ~new_D3706_ | ~new_D3731_;
  assign new_D3762_ = new_D3739_ & new_D3759_;
  assign new_D3763_ = ~new_D3739_ & ~new_D3759_;
  assign new_D3764_ = new_D3768_ | new_D3769_;
  assign new_D3765_ = ~new_D3710_ & new_D3724_;
  assign new_D3766_ = new_D3770_ | new_D3771_;
  assign new_D3767_ = new_D3710_ & new_D3724_;
  assign new_D3768_ = ~new_D3710_ & ~new_D3724_;
  assign new_D3769_ = new_D3710_ & ~new_D3724_;
  assign new_D3770_ = new_D3710_ & ~new_D3724_;
  assign new_D3771_ = ~new_D3710_ & new_D3724_;
  assign new_D3772_ = new_E6647_;
  assign new_D3773_ = new_E6714_;
  assign new_D3774_ = new_E6781_;
  assign new_D3775_ = new_E6848_;
  assign new_D3776_ = new_E6915_;
  assign new_D3777_ = new_E6982_;
  assign new_D3778_ = new_D3785_ & new_D3784_;
  assign new_D3779_ = new_D3787_ | new_D3786_;
  assign new_D3780_ = new_D3789_ | new_D3788_;
  assign new_D3781_ = new_D3791_ & new_D3790_;
  assign new_D3782_ = new_D3791_ & new_D3792_;
  assign new_D3783_ = new_D3784_ | new_D3793_;
  assign new_D3784_ = new_D3773_ | new_D3796_;
  assign new_D3785_ = new_D3795_ | new_D3794_;
  assign new_D3786_ = new_D3800_ & new_D3799_;
  assign new_D3787_ = new_D3798_ & new_D3797_;
  assign new_D3788_ = new_D3803_ | new_D3802_;
  assign new_D3789_ = new_D3798_ & new_D3801_;
  assign new_D3790_ = new_D3773_ | new_D3806_;
  assign new_D3791_ = new_D3805_ | new_D3804_;
  assign new_D3792_ = new_D3808_ | new_D3807_;
  assign new_D3793_ = ~new_D3784_ & new_D3810_;
  assign new_D3794_ = ~new_D3786_ & new_D3798_;
  assign new_D3795_ = new_D3786_ & ~new_D3798_;
  assign new_D3796_ = new_D3772_ & ~new_D3773_;
  assign new_D3797_ = ~new_D3819_ | ~new_D3820_;
  assign new_D3798_ = new_D3812_ | new_D3814_;
  assign new_D3799_ = new_D3822_ | new_D3821_;
  assign new_D3800_ = new_D3816_ | new_D3815_;
  assign new_D3801_ = ~new_D3824_ | ~new_D3823_;
  assign new_D3802_ = ~new_D3825_ & new_D3826_;
  assign new_D3803_ = new_D3825_ & ~new_D3826_;
  assign new_D3804_ = ~new_D3772_ & new_D3773_;
  assign new_D3805_ = new_D3772_ & ~new_D3773_;
  assign new_D3806_ = ~new_D3788_ | new_D3798_;
  assign new_D3807_ = new_D3788_ & new_D3798_;
  assign new_D3808_ = ~new_D3788_ & ~new_D3798_;
  assign new_D3809_ = new_D3830_ | new_D3829_;
  assign new_D3810_ = new_D3776_ | new_D3809_;
  assign new_D3811_ = new_D3834_ | new_D3833_;
  assign new_D3812_ = ~new_D3776_ & new_D3811_;
  assign new_D3813_ = new_D3832_ | new_D3831_;
  assign new_D3814_ = new_D3776_ & new_D3813_;
  assign new_D3815_ = new_D3774_ & ~new_D3784_;
  assign new_D3816_ = ~new_D3774_ & new_D3784_;
  assign new_D3817_ = ~new_D3773_ | ~new_D3798_;
  assign new_D3818_ = new_D3784_ & new_D3817_;
  assign new_D3819_ = ~new_D3784_ & ~new_D3818_;
  assign new_D3820_ = new_D3784_ | new_D3817_;
  assign new_D3821_ = ~new_D3774_ & new_D3775_;
  assign new_D3822_ = new_D3774_ & ~new_D3775_;
  assign new_D3823_ = new_D3791_ | new_D3828_;
  assign new_D3824_ = ~new_D3791_ & ~new_D3827_;
  assign new_D3825_ = new_D3774_ | new_D3791_;
  assign new_D3826_ = new_D3774_ | new_D3775_;
  assign new_D3827_ = new_D3791_ & new_D3828_;
  assign new_D3828_ = ~new_D3773_ | ~new_D3798_;
  assign new_D3829_ = new_D3806_ & new_D3826_;
  assign new_D3830_ = ~new_D3806_ & ~new_D3826_;
  assign new_D3831_ = new_D3835_ | new_D3836_;
  assign new_D3832_ = ~new_D3777_ & new_D3791_;
  assign new_D3833_ = new_D3837_ | new_D3838_;
  assign new_D3834_ = new_D3777_ & new_D3791_;
  assign new_D3835_ = ~new_D3777_ & ~new_D3791_;
  assign new_D3836_ = new_D3777_ & ~new_D3791_;
  assign new_D3837_ = new_D3777_ & ~new_D3791_;
  assign new_D3838_ = ~new_D3777_ & new_D3791_;
  assign new_D3839_ = new_E7049_;
  assign new_D3840_ = new_E7116_;
  assign new_D3841_ = new_E7183_;
  assign new_D3842_ = new_E7250_;
  assign new_D3843_ = new_E7317_;
  assign new_D3844_ = new_E7384_;
  assign new_D3845_ = new_D3852_ & new_D3851_;
  assign new_D3846_ = new_D3854_ | new_D3853_;
  assign new_D3847_ = new_D3856_ | new_D3855_;
  assign new_D3848_ = new_D3858_ & new_D3857_;
  assign new_D3849_ = new_D3858_ & new_D3859_;
  assign new_D3850_ = new_D3851_ | new_D3860_;
  assign new_D3851_ = new_D3840_ | new_D3863_;
  assign new_D3852_ = new_D3862_ | new_D3861_;
  assign new_D3853_ = new_D3867_ & new_D3866_;
  assign new_D3854_ = new_D3865_ & new_D3864_;
  assign new_D3855_ = new_D3870_ | new_D3869_;
  assign new_D3856_ = new_D3865_ & new_D3868_;
  assign new_D3857_ = new_D3840_ | new_D3873_;
  assign new_D3858_ = new_D3872_ | new_D3871_;
  assign new_D3859_ = new_D3875_ | new_D3874_;
  assign new_D3860_ = ~new_D3851_ & new_D3877_;
  assign new_D3861_ = ~new_D3853_ & new_D3865_;
  assign new_D3862_ = new_D3853_ & ~new_D3865_;
  assign new_D3863_ = new_D3839_ & ~new_D3840_;
  assign new_D3864_ = ~new_D3886_ | ~new_D3887_;
  assign new_D3865_ = new_D3879_ | new_D3881_;
  assign new_D3866_ = new_D3889_ | new_D3888_;
  assign new_D3867_ = new_D3883_ | new_D3882_;
  assign new_D3868_ = ~new_D3891_ | ~new_D3890_;
  assign new_D3869_ = ~new_D3892_ & new_D3893_;
  assign new_D3870_ = new_D3892_ & ~new_D3893_;
  assign new_D3871_ = ~new_D3839_ & new_D3840_;
  assign new_D3872_ = new_D3839_ & ~new_D3840_;
  assign new_D3873_ = ~new_D3855_ | new_D3865_;
  assign new_D3874_ = new_D3855_ & new_D3865_;
  assign new_D3875_ = ~new_D3855_ & ~new_D3865_;
  assign new_D3876_ = new_D3897_ | new_D3896_;
  assign new_D3877_ = new_D3843_ | new_D3876_;
  assign new_D3878_ = new_D3901_ | new_D3900_;
  assign new_D3879_ = ~new_D3843_ & new_D3878_;
  assign new_D3880_ = new_D3899_ | new_D3898_;
  assign new_D3881_ = new_D3843_ & new_D3880_;
  assign new_D3882_ = new_D3841_ & ~new_D3851_;
  assign new_D3883_ = ~new_D3841_ & new_D3851_;
  assign new_D3884_ = ~new_D3840_ | ~new_D3865_;
  assign new_D3885_ = new_D3851_ & new_D3884_;
  assign new_D3886_ = ~new_D3851_ & ~new_D3885_;
  assign new_D3887_ = new_D3851_ | new_D3884_;
  assign new_D3888_ = ~new_D3841_ & new_D3842_;
  assign new_D3889_ = new_D3841_ & ~new_D3842_;
  assign new_D3890_ = new_D3858_ | new_D3895_;
  assign new_D3891_ = ~new_D3858_ & ~new_D3894_;
  assign new_D3892_ = new_D3841_ | new_D3858_;
  assign new_D3893_ = new_D3841_ | new_D3842_;
  assign new_D3894_ = new_D3858_ & new_D3895_;
  assign new_D3895_ = ~new_D3840_ | ~new_D3865_;
  assign new_D3896_ = new_D3873_ & new_D3893_;
  assign new_D3897_ = ~new_D3873_ & ~new_D3893_;
  assign new_D3898_ = new_D3902_ | new_D3903_;
  assign new_D3899_ = ~new_D3844_ & new_D3858_;
  assign new_D3900_ = new_D3904_ | new_D3905_;
  assign new_D3901_ = new_D3844_ & new_D3858_;
  assign new_D3902_ = ~new_D3844_ & ~new_D3858_;
  assign new_D3903_ = new_D3844_ & ~new_D3858_;
  assign new_D3904_ = new_D3844_ & ~new_D3858_;
  assign new_D3905_ = ~new_D3844_ & new_D3858_;
  assign new_D3906_ = new_E7451_;
  assign new_D3907_ = new_E7518_;
  assign new_D3908_ = new_E7585_;
  assign new_D3909_ = new_E7652_;
  assign new_D3910_ = new_E7719_;
  assign new_D3911_ = new_E7786_;
  assign new_D3912_ = new_D3919_ & new_D3918_;
  assign new_D3913_ = new_D3921_ | new_D3920_;
  assign new_D3914_ = new_D3923_ | new_D3922_;
  assign new_D3915_ = new_D3925_ & new_D3924_;
  assign new_D3916_ = new_D3925_ & new_D3926_;
  assign new_D3917_ = new_D3918_ | new_D3927_;
  assign new_D3918_ = new_D3907_ | new_D3930_;
  assign new_D3919_ = new_D3929_ | new_D3928_;
  assign new_D3920_ = new_D3934_ & new_D3933_;
  assign new_D3921_ = new_D3932_ & new_D3931_;
  assign new_D3922_ = new_D3937_ | new_D3936_;
  assign new_D3923_ = new_D3932_ & new_D3935_;
  assign new_D3924_ = new_D3907_ | new_D3940_;
  assign new_D3925_ = new_D3939_ | new_D3938_;
  assign new_D3926_ = new_D3942_ | new_D3941_;
  assign new_D3927_ = ~new_D3918_ & new_D3944_;
  assign new_D3928_ = ~new_D3920_ & new_D3932_;
  assign new_D3929_ = new_D3920_ & ~new_D3932_;
  assign new_D3930_ = new_D3906_ & ~new_D3907_;
  assign new_D3931_ = ~new_D3953_ | ~new_D3954_;
  assign new_D3932_ = new_D3946_ | new_D3948_;
  assign new_D3933_ = new_D3956_ | new_D3955_;
  assign new_D3934_ = new_D3950_ | new_D3949_;
  assign new_D3935_ = ~new_D3958_ | ~new_D3957_;
  assign new_D3936_ = ~new_D3959_ & new_D3960_;
  assign new_D3937_ = new_D3959_ & ~new_D3960_;
  assign new_D3938_ = ~new_D3906_ & new_D3907_;
  assign new_D3939_ = new_D3906_ & ~new_D3907_;
  assign new_D3940_ = ~new_D3922_ | new_D3932_;
  assign new_D3941_ = new_D3922_ & new_D3932_;
  assign new_D3942_ = ~new_D3922_ & ~new_D3932_;
  assign new_D3943_ = new_D3964_ | new_D3963_;
  assign new_D3944_ = new_D3910_ | new_D3943_;
  assign new_D3945_ = new_D3968_ | new_D3967_;
  assign new_D3946_ = ~new_D3910_ & new_D3945_;
  assign new_D3947_ = new_D3966_ | new_D3965_;
  assign new_D3948_ = new_D3910_ & new_D3947_;
  assign new_D3949_ = new_D3908_ & ~new_D3918_;
  assign new_D3950_ = ~new_D3908_ & new_D3918_;
  assign new_D3951_ = ~new_D3907_ | ~new_D3932_;
  assign new_D3952_ = new_D3918_ & new_D3951_;
  assign new_D3953_ = ~new_D3918_ & ~new_D3952_;
  assign new_D3954_ = new_D3918_ | new_D3951_;
  assign new_D3955_ = ~new_D3908_ & new_D3909_;
  assign new_D3956_ = new_D3908_ & ~new_D3909_;
  assign new_D3957_ = new_D3925_ | new_D3962_;
  assign new_D3958_ = ~new_D3925_ & ~new_D3961_;
  assign new_D3959_ = new_D3908_ | new_D3925_;
  assign new_D3960_ = new_D3908_ | new_D3909_;
  assign new_D3961_ = new_D3925_ & new_D3962_;
  assign new_D3962_ = ~new_D3907_ | ~new_D3932_;
  assign new_D3963_ = new_D3940_ & new_D3960_;
  assign new_D3964_ = ~new_D3940_ & ~new_D3960_;
  assign new_D3965_ = new_D3969_ | new_D3970_;
  assign new_D3966_ = ~new_D3911_ & new_D3925_;
  assign new_D3967_ = new_D3971_ | new_D3972_;
  assign new_D3968_ = new_D3911_ & new_D3925_;
  assign new_D3969_ = ~new_D3911_ & ~new_D3925_;
  assign new_D3970_ = new_D3911_ & ~new_D3925_;
  assign new_D3971_ = new_D3911_ & ~new_D3925_;
  assign new_D3972_ = ~new_D3911_ & new_D3925_;
  assign new_D3973_ = new_E7853_;
  assign new_D3974_ = new_E7920_;
  assign new_D3975_ = new_E7987_;
  assign new_D3976_ = new_E8054_;
  assign new_D3977_ = new_E8121_;
  assign new_D3978_ = new_E8188_;
  assign new_D3979_ = new_D3986_ & new_D3985_;
  assign new_D3980_ = new_D3988_ | new_D3987_;
  assign new_D3981_ = new_D3990_ | new_D3989_;
  assign new_D3982_ = new_D3992_ & new_D3991_;
  assign new_D3983_ = new_D3992_ & new_D3993_;
  assign new_D3984_ = new_D3985_ | new_D3994_;
  assign new_D3985_ = new_D3974_ | new_D3997_;
  assign new_D3986_ = new_D3996_ | new_D3995_;
  assign new_D3987_ = new_D4001_ & new_D4000_;
  assign new_D3988_ = new_D3999_ & new_D3998_;
  assign new_D3989_ = new_D4004_ | new_D4003_;
  assign new_D3990_ = new_D3999_ & new_D4002_;
  assign new_D3991_ = new_D3974_ | new_D4007_;
  assign new_D3992_ = new_D4006_ | new_D4005_;
  assign new_D3993_ = new_D4009_ | new_D4008_;
  assign new_D3994_ = ~new_D3985_ & new_D4011_;
  assign new_D3995_ = ~new_D3987_ & new_D3999_;
  assign new_D3996_ = new_D3987_ & ~new_D3999_;
  assign new_D3997_ = new_D3973_ & ~new_D3974_;
  assign new_D3998_ = ~new_D4020_ | ~new_D4021_;
  assign new_D3999_ = new_D4013_ | new_D4015_;
  assign new_D4000_ = new_D4023_ | new_D4022_;
  assign new_D4001_ = new_D4017_ | new_D4016_;
  assign new_D4002_ = ~new_D4025_ | ~new_D4024_;
  assign new_D4003_ = ~new_D4026_ & new_D4027_;
  assign new_D4004_ = new_D4026_ & ~new_D4027_;
  assign new_D4005_ = ~new_D3973_ & new_D3974_;
  assign new_D4006_ = new_D3973_ & ~new_D3974_;
  assign new_D4007_ = ~new_D3989_ | new_D3999_;
  assign new_D4008_ = new_D3989_ & new_D3999_;
  assign new_D4009_ = ~new_D3989_ & ~new_D3999_;
  assign new_D4010_ = new_D4031_ | new_D4030_;
  assign new_D4011_ = new_D3977_ | new_D4010_;
  assign new_D4012_ = new_D4035_ | new_D4034_;
  assign new_D4013_ = ~new_D3977_ & new_D4012_;
  assign new_D4014_ = new_D4033_ | new_D4032_;
  assign new_D4015_ = new_D3977_ & new_D4014_;
  assign new_D4016_ = new_D3975_ & ~new_D3985_;
  assign new_D4017_ = ~new_D3975_ & new_D3985_;
  assign new_D4018_ = ~new_D3974_ | ~new_D3999_;
  assign new_D4019_ = new_D3985_ & new_D4018_;
  assign new_D4020_ = ~new_D3985_ & ~new_D4019_;
  assign new_D4021_ = new_D3985_ | new_D4018_;
  assign new_D4022_ = ~new_D3975_ & new_D3976_;
  assign new_D4023_ = new_D3975_ & ~new_D3976_;
  assign new_D4024_ = new_D3992_ | new_D4029_;
  assign new_D4025_ = ~new_D3992_ & ~new_D4028_;
  assign new_D4026_ = new_D3975_ | new_D3992_;
  assign new_D4027_ = new_D3975_ | new_D3976_;
  assign new_D4028_ = new_D3992_ & new_D4029_;
  assign new_D4029_ = ~new_D3974_ | ~new_D3999_;
  assign new_D4030_ = new_D4007_ & new_D4027_;
  assign new_D4031_ = ~new_D4007_ & ~new_D4027_;
  assign new_D4032_ = new_D4036_ | new_D4037_;
  assign new_D4033_ = ~new_D3978_ & new_D3992_;
  assign new_D4034_ = new_D4038_ | new_D4039_;
  assign new_D4035_ = new_D3978_ & new_D3992_;
  assign new_D4036_ = ~new_D3978_ & ~new_D3992_;
  assign new_D4037_ = new_D3978_ & ~new_D3992_;
  assign new_D4038_ = new_D3978_ & ~new_D3992_;
  assign new_D4039_ = ~new_D3978_ & new_D3992_;
  assign new_D4040_ = new_E8255_;
  assign new_D4041_ = new_E8322_;
  assign new_D4042_ = new_E8389_;
  assign new_D4043_ = new_E8456_;
  assign new_D4044_ = new_E8523_;
  assign new_D4045_ = new_E8590_;
  assign new_D4046_ = new_D4053_ & new_D4052_;
  assign new_D4047_ = new_D4055_ | new_D4054_;
  assign new_D4048_ = new_D4057_ | new_D4056_;
  assign new_D4049_ = new_D4059_ & new_D4058_;
  assign new_D4050_ = new_D4059_ & new_D4060_;
  assign new_D4051_ = new_D4052_ | new_D4061_;
  assign new_D4052_ = new_D4041_ | new_D4064_;
  assign new_D4053_ = new_D4063_ | new_D4062_;
  assign new_D4054_ = new_D4068_ & new_D4067_;
  assign new_D4055_ = new_D4066_ & new_D4065_;
  assign new_D4056_ = new_D4071_ | new_D4070_;
  assign new_D4057_ = new_D4066_ & new_D4069_;
  assign new_D4058_ = new_D4041_ | new_D4074_;
  assign new_D4059_ = new_D4073_ | new_D4072_;
  assign new_D4060_ = new_D4076_ | new_D4075_;
  assign new_D4061_ = ~new_D4052_ & new_D4078_;
  assign new_D4062_ = ~new_D4054_ & new_D4066_;
  assign new_D4063_ = new_D4054_ & ~new_D4066_;
  assign new_D4064_ = new_D4040_ & ~new_D4041_;
  assign new_D4065_ = ~new_D4087_ | ~new_D4088_;
  assign new_D4066_ = new_D4080_ | new_D4082_;
  assign new_D4067_ = new_D4090_ | new_D4089_;
  assign new_D4068_ = new_D4084_ | new_D4083_;
  assign new_D4069_ = ~new_D4092_ | ~new_D4091_;
  assign new_D4070_ = ~new_D4093_ & new_D4094_;
  assign new_D4071_ = new_D4093_ & ~new_D4094_;
  assign new_D4072_ = ~new_D4040_ & new_D4041_;
  assign new_D4073_ = new_D4040_ & ~new_D4041_;
  assign new_D4074_ = ~new_D4056_ | new_D4066_;
  assign new_D4075_ = new_D4056_ & new_D4066_;
  assign new_D4076_ = ~new_D4056_ & ~new_D4066_;
  assign new_D4077_ = new_D4098_ | new_D4097_;
  assign new_D4078_ = new_D4044_ | new_D4077_;
  assign new_D4079_ = new_D4102_ | new_D4101_;
  assign new_D4080_ = ~new_D4044_ & new_D4079_;
  assign new_D4081_ = new_D4100_ | new_D4099_;
  assign new_D4082_ = new_D4044_ & new_D4081_;
  assign new_D4083_ = new_D4042_ & ~new_D4052_;
  assign new_D4084_ = ~new_D4042_ & new_D4052_;
  assign new_D4085_ = ~new_D4041_ | ~new_D4066_;
  assign new_D4086_ = new_D4052_ & new_D4085_;
  assign new_D4087_ = ~new_D4052_ & ~new_D4086_;
  assign new_D4088_ = new_D4052_ | new_D4085_;
  assign new_D4089_ = ~new_D4042_ & new_D4043_;
  assign new_D4090_ = new_D4042_ & ~new_D4043_;
  assign new_D4091_ = new_D4059_ | new_D4096_;
  assign new_D4092_ = ~new_D4059_ & ~new_D4095_;
  assign new_D4093_ = new_D4042_ | new_D4059_;
  assign new_D4094_ = new_D4042_ | new_D4043_;
  assign new_D4095_ = new_D4059_ & new_D4096_;
  assign new_D4096_ = ~new_D4041_ | ~new_D4066_;
  assign new_D4097_ = new_D4074_ & new_D4094_;
  assign new_D4098_ = ~new_D4074_ & ~new_D4094_;
  assign new_D4099_ = new_D4103_ | new_D4104_;
  assign new_D4100_ = ~new_D4045_ & new_D4059_;
  assign new_D4101_ = new_D4105_ | new_D4106_;
  assign new_D4102_ = new_D4045_ & new_D4059_;
  assign new_D4103_ = ~new_D4045_ & ~new_D4059_;
  assign new_D4104_ = new_D4045_ & ~new_D4059_;
  assign new_D4105_ = new_D4045_ & ~new_D4059_;
  assign new_D4106_ = ~new_D4045_ & new_D4059_;
  assign new_D4107_ = new_E8657_;
  assign new_D4108_ = new_E8724_;
  assign new_D4109_ = new_E8791_;
  assign new_D4110_ = new_E8858_;
  assign new_D4111_ = new_E8925_;
  assign new_D4112_ = new_E8992_;
  assign new_D4113_ = new_D4120_ & new_D4119_;
  assign new_D4114_ = new_D4122_ | new_D4121_;
  assign new_D4115_ = new_D4124_ | new_D4123_;
  assign new_D4116_ = new_D4126_ & new_D4125_;
  assign new_D4117_ = new_D4126_ & new_D4127_;
  assign new_D4118_ = new_D4119_ | new_D4128_;
  assign new_D4119_ = new_D4108_ | new_D4131_;
  assign new_D4120_ = new_D4130_ | new_D4129_;
  assign new_D4121_ = new_D4135_ & new_D4134_;
  assign new_D4122_ = new_D4133_ & new_D4132_;
  assign new_D4123_ = new_D4138_ | new_D4137_;
  assign new_D4124_ = new_D4133_ & new_D4136_;
  assign new_D4125_ = new_D4108_ | new_D4141_;
  assign new_D4126_ = new_D4140_ | new_D4139_;
  assign new_D4127_ = new_D4143_ | new_D4142_;
  assign new_D4128_ = ~new_D4119_ & new_D4145_;
  assign new_D4129_ = ~new_D4121_ & new_D4133_;
  assign new_D4130_ = new_D4121_ & ~new_D4133_;
  assign new_D4131_ = new_D4107_ & ~new_D4108_;
  assign new_D4132_ = ~new_D4154_ | ~new_D4155_;
  assign new_D4133_ = new_D4147_ | new_D4149_;
  assign new_D4134_ = new_D4157_ | new_D4156_;
  assign new_D4135_ = new_D4151_ | new_D4150_;
  assign new_D4136_ = ~new_D4159_ | ~new_D4158_;
  assign new_D4137_ = ~new_D4160_ & new_D4161_;
  assign new_D4138_ = new_D4160_ & ~new_D4161_;
  assign new_D4139_ = ~new_D4107_ & new_D4108_;
  assign new_D4140_ = new_D4107_ & ~new_D4108_;
  assign new_D4141_ = ~new_D4123_ | new_D4133_;
  assign new_D4142_ = new_D4123_ & new_D4133_;
  assign new_D4143_ = ~new_D4123_ & ~new_D4133_;
  assign new_D4144_ = new_D4165_ | new_D4164_;
  assign new_D4145_ = new_D4111_ | new_D4144_;
  assign new_D4146_ = new_D4169_ | new_D4168_;
  assign new_D4147_ = ~new_D4111_ & new_D4146_;
  assign new_D4148_ = new_D4167_ | new_D4166_;
  assign new_D4149_ = new_D4111_ & new_D4148_;
  assign new_D4150_ = new_D4109_ & ~new_D4119_;
  assign new_D4151_ = ~new_D4109_ & new_D4119_;
  assign new_D4152_ = ~new_D4108_ | ~new_D4133_;
  assign new_D4153_ = new_D4119_ & new_D4152_;
  assign new_D4154_ = ~new_D4119_ & ~new_D4153_;
  assign new_D4155_ = new_D4119_ | new_D4152_;
  assign new_D4156_ = ~new_D4109_ & new_D4110_;
  assign new_D4157_ = new_D4109_ & ~new_D4110_;
  assign new_D4158_ = new_D4126_ | new_D4163_;
  assign new_D4159_ = ~new_D4126_ & ~new_D4162_;
  assign new_D4160_ = new_D4109_ | new_D4126_;
  assign new_D4161_ = new_D4109_ | new_D4110_;
  assign new_D4162_ = new_D4126_ & new_D4163_;
  assign new_D4163_ = ~new_D4108_ | ~new_D4133_;
  assign new_D4164_ = new_D4141_ & new_D4161_;
  assign new_D4165_ = ~new_D4141_ & ~new_D4161_;
  assign new_D4166_ = new_D4170_ | new_D4171_;
  assign new_D4167_ = ~new_D4112_ & new_D4126_;
  assign new_D4168_ = new_D4172_ | new_D4173_;
  assign new_D4169_ = new_D4112_ & new_D4126_;
  assign new_D4170_ = ~new_D4112_ & ~new_D4126_;
  assign new_D4171_ = new_D4112_ & ~new_D4126_;
  assign new_D4172_ = new_D4112_ & ~new_D4126_;
  assign new_D4173_ = ~new_D4112_ & new_D4126_;
  assign new_D4174_ = new_E9059_;
  assign new_D4175_ = new_E9126_;
  assign new_D4176_ = new_E9193_;
  assign new_D4177_ = new_E9260_;
  assign new_D4178_ = new_E9327_;
  assign new_D4179_ = new_E9394_;
  assign new_D4180_ = new_D4187_ & new_D4186_;
  assign new_D4181_ = new_D4189_ | new_D4188_;
  assign new_D4182_ = new_D4191_ | new_D4190_;
  assign new_D4183_ = new_D4193_ & new_D4192_;
  assign new_D4184_ = new_D4193_ & new_D4194_;
  assign new_D4185_ = new_D4186_ | new_D4195_;
  assign new_D4186_ = new_D4175_ | new_D4198_;
  assign new_D4187_ = new_D4197_ | new_D4196_;
  assign new_D4188_ = new_D4202_ & new_D4201_;
  assign new_D4189_ = new_D4200_ & new_D4199_;
  assign new_D4190_ = new_D4205_ | new_D4204_;
  assign new_D4191_ = new_D4200_ & new_D4203_;
  assign new_D4192_ = new_D4175_ | new_D4208_;
  assign new_D4193_ = new_D4207_ | new_D4206_;
  assign new_D4194_ = new_D4210_ | new_D4209_;
  assign new_D4195_ = ~new_D4186_ & new_D4212_;
  assign new_D4196_ = ~new_D4188_ & new_D4200_;
  assign new_D4197_ = new_D4188_ & ~new_D4200_;
  assign new_D4198_ = new_D4174_ & ~new_D4175_;
  assign new_D4199_ = ~new_D4221_ | ~new_D4222_;
  assign new_D4200_ = new_D4214_ | new_D4216_;
  assign new_D4201_ = new_D4224_ | new_D4223_;
  assign new_D4202_ = new_D4218_ | new_D4217_;
  assign new_D4203_ = ~new_D4226_ | ~new_D4225_;
  assign new_D4204_ = ~new_D4227_ & new_D4228_;
  assign new_D4205_ = new_D4227_ & ~new_D4228_;
  assign new_D4206_ = ~new_D4174_ & new_D4175_;
  assign new_D4207_ = new_D4174_ & ~new_D4175_;
  assign new_D4208_ = ~new_D4190_ | new_D4200_;
  assign new_D4209_ = new_D4190_ & new_D4200_;
  assign new_D4210_ = ~new_D4190_ & ~new_D4200_;
  assign new_D4211_ = new_D4232_ | new_D4231_;
  assign new_D4212_ = new_D4178_ | new_D4211_;
  assign new_D4213_ = new_D4236_ | new_D4235_;
  assign new_D4214_ = ~new_D4178_ & new_D4213_;
  assign new_D4215_ = new_D4234_ | new_D4233_;
  assign new_D4216_ = new_D4178_ & new_D4215_;
  assign new_D4217_ = new_D4176_ & ~new_D4186_;
  assign new_D4218_ = ~new_D4176_ & new_D4186_;
  assign new_D4219_ = ~new_D4175_ | ~new_D4200_;
  assign new_D4220_ = new_D4186_ & new_D4219_;
  assign new_D4221_ = ~new_D4186_ & ~new_D4220_;
  assign new_D4222_ = new_D4186_ | new_D4219_;
  assign new_D4223_ = ~new_D4176_ & new_D4177_;
  assign new_D4224_ = new_D4176_ & ~new_D4177_;
  assign new_D4225_ = new_D4193_ | new_D4230_;
  assign new_D4226_ = ~new_D4193_ & ~new_D4229_;
  assign new_D4227_ = new_D4176_ | new_D4193_;
  assign new_D4228_ = new_D4176_ | new_D4177_;
  assign new_D4229_ = new_D4193_ & new_D4230_;
  assign new_D4230_ = ~new_D4175_ | ~new_D4200_;
  assign new_D4231_ = new_D4208_ & new_D4228_;
  assign new_D4232_ = ~new_D4208_ & ~new_D4228_;
  assign new_D4233_ = new_D4237_ | new_D4238_;
  assign new_D4234_ = ~new_D4179_ & new_D4193_;
  assign new_D4235_ = new_D4239_ | new_D4240_;
  assign new_D4236_ = new_D4179_ & new_D4193_;
  assign new_D4237_ = ~new_D4179_ & ~new_D4193_;
  assign new_D4238_ = new_D4179_ & ~new_D4193_;
  assign new_D4239_ = new_D4179_ & ~new_D4193_;
  assign new_D4240_ = ~new_D4179_ & new_D4193_;
  assign new_D4241_ = new_E9461_;
  assign new_D4242_ = new_E9528_;
  assign new_D4243_ = new_E9595_;
  assign new_D4244_ = new_E9662_;
  assign new_D4245_ = new_E9729_;
  assign new_D4246_ = new_E9796_;
  assign new_D4247_ = new_D4254_ & new_D4253_;
  assign new_D4248_ = new_D4256_ | new_D4255_;
  assign new_D4249_ = new_D4258_ | new_D4257_;
  assign new_D4250_ = new_D4260_ & new_D4259_;
  assign new_D4251_ = new_D4260_ & new_D4261_;
  assign new_D4252_ = new_D4253_ | new_D4262_;
  assign new_D4253_ = new_D4242_ | new_D4265_;
  assign new_D4254_ = new_D4264_ | new_D4263_;
  assign new_D4255_ = new_D4269_ & new_D4268_;
  assign new_D4256_ = new_D4267_ & new_D4266_;
  assign new_D4257_ = new_D4272_ | new_D4271_;
  assign new_D4258_ = new_D4267_ & new_D4270_;
  assign new_D4259_ = new_D4242_ | new_D4275_;
  assign new_D4260_ = new_D4274_ | new_D4273_;
  assign new_D4261_ = new_D4277_ | new_D4276_;
  assign new_D4262_ = ~new_D4253_ & new_D4279_;
  assign new_D4263_ = ~new_D4255_ & new_D4267_;
  assign new_D4264_ = new_D4255_ & ~new_D4267_;
  assign new_D4265_ = new_D4241_ & ~new_D4242_;
  assign new_D4266_ = ~new_D4288_ | ~new_D4289_;
  assign new_D4267_ = new_D4281_ | new_D4283_;
  assign new_D4268_ = new_D4291_ | new_D4290_;
  assign new_D4269_ = new_D4285_ | new_D4284_;
  assign new_D4270_ = ~new_D4293_ | ~new_D4292_;
  assign new_D4271_ = ~new_D4294_ & new_D4295_;
  assign new_D4272_ = new_D4294_ & ~new_D4295_;
  assign new_D4273_ = ~new_D4241_ & new_D4242_;
  assign new_D4274_ = new_D4241_ & ~new_D4242_;
  assign new_D4275_ = ~new_D4257_ | new_D4267_;
  assign new_D4276_ = new_D4257_ & new_D4267_;
  assign new_D4277_ = ~new_D4257_ & ~new_D4267_;
  assign new_D4278_ = new_D4299_ | new_D4298_;
  assign new_D4279_ = new_D4245_ | new_D4278_;
  assign new_D4280_ = new_D4303_ | new_D4302_;
  assign new_D4281_ = ~new_D4245_ & new_D4280_;
  assign new_D4282_ = new_D4301_ | new_D4300_;
  assign new_D4283_ = new_D4245_ & new_D4282_;
  assign new_D4284_ = new_D4243_ & ~new_D4253_;
  assign new_D4285_ = ~new_D4243_ & new_D4253_;
  assign new_D4286_ = ~new_D4242_ | ~new_D4267_;
  assign new_D4287_ = new_D4253_ & new_D4286_;
  assign new_D4288_ = ~new_D4253_ & ~new_D4287_;
  assign new_D4289_ = new_D4253_ | new_D4286_;
  assign new_D4290_ = ~new_D4243_ & new_D4244_;
  assign new_D4291_ = new_D4243_ & ~new_D4244_;
  assign new_D4292_ = new_D4260_ | new_D4297_;
  assign new_D4293_ = ~new_D4260_ & ~new_D4296_;
  assign new_D4294_ = new_D4243_ | new_D4260_;
  assign new_D4295_ = new_D4243_ | new_D4244_;
  assign new_D4296_ = new_D4260_ & new_D4297_;
  assign new_D4297_ = ~new_D4242_ | ~new_D4267_;
  assign new_D4298_ = new_D4275_ & new_D4295_;
  assign new_D4299_ = ~new_D4275_ & ~new_D4295_;
  assign new_D4300_ = new_D4304_ | new_D4305_;
  assign new_D4301_ = ~new_D4246_ & new_D4260_;
  assign new_D4302_ = new_D4306_ | new_D4307_;
  assign new_D4303_ = new_D4246_ & new_D4260_;
  assign new_D4304_ = ~new_D4246_ & ~new_D4260_;
  assign new_D4305_ = new_D4246_ & ~new_D4260_;
  assign new_D4306_ = new_D4246_ & ~new_D4260_;
  assign new_D4307_ = ~new_D4246_ & new_D4260_;
  assign new_D4308_ = new_E9863_;
  assign new_D4309_ = new_E9930_;
  assign new_D4310_ = new_E9997_;
  assign new_D4311_ = new_F65_;
  assign new_D4312_ = new_F132_;
  assign new_D4313_ = new_F199_;
  assign new_D4314_ = new_D4321_ & new_D4320_;
  assign new_D4315_ = new_D4323_ | new_D4322_;
  assign new_D4316_ = new_D4325_ | new_D4324_;
  assign new_D4317_ = new_D4327_ & new_D4326_;
  assign new_D4318_ = new_D4327_ & new_D4328_;
  assign new_D4319_ = new_D4320_ | new_D4329_;
  assign new_D4320_ = new_D4309_ | new_D4332_;
  assign new_D4321_ = new_D4331_ | new_D4330_;
  assign new_D4322_ = new_D4336_ & new_D4335_;
  assign new_D4323_ = new_D4334_ & new_D4333_;
  assign new_D4324_ = new_D4339_ | new_D4338_;
  assign new_D4325_ = new_D4334_ & new_D4337_;
  assign new_D4326_ = new_D4309_ | new_D4342_;
  assign new_D4327_ = new_D4341_ | new_D4340_;
  assign new_D4328_ = new_D4344_ | new_D4343_;
  assign new_D4329_ = ~new_D4320_ & new_D4346_;
  assign new_D4330_ = ~new_D4322_ & new_D4334_;
  assign new_D4331_ = new_D4322_ & ~new_D4334_;
  assign new_D4332_ = new_D4308_ & ~new_D4309_;
  assign new_D4333_ = ~new_D4355_ | ~new_D4356_;
  assign new_D4334_ = new_D4348_ | new_D4350_;
  assign new_D4335_ = new_D4358_ | new_D4357_;
  assign new_D4336_ = new_D4352_ | new_D4351_;
  assign new_D4337_ = ~new_D4360_ | ~new_D4359_;
  assign new_D4338_ = ~new_D4361_ & new_D4362_;
  assign new_D4339_ = new_D4361_ & ~new_D4362_;
  assign new_D4340_ = ~new_D4308_ & new_D4309_;
  assign new_D4341_ = new_D4308_ & ~new_D4309_;
  assign new_D4342_ = ~new_D4324_ | new_D4334_;
  assign new_D4343_ = new_D4324_ & new_D4334_;
  assign new_D4344_ = ~new_D4324_ & ~new_D4334_;
  assign new_D4345_ = new_D4366_ | new_D4365_;
  assign new_D4346_ = new_D4312_ | new_D4345_;
  assign new_D4347_ = new_D4370_ | new_D4369_;
  assign new_D4348_ = ~new_D4312_ & new_D4347_;
  assign new_D4349_ = new_D4368_ | new_D4367_;
  assign new_D4350_ = new_D4312_ & new_D4349_;
  assign new_D4351_ = new_D4310_ & ~new_D4320_;
  assign new_D4352_ = ~new_D4310_ & new_D4320_;
  assign new_D4353_ = ~new_D4309_ | ~new_D4334_;
  assign new_D4354_ = new_D4320_ & new_D4353_;
  assign new_D4355_ = ~new_D4320_ & ~new_D4354_;
  assign new_D4356_ = new_D4320_ | new_D4353_;
  assign new_D4357_ = ~new_D4310_ & new_D4311_;
  assign new_D4358_ = new_D4310_ & ~new_D4311_;
  assign new_D4359_ = new_D4327_ | new_D4364_;
  assign new_D4360_ = ~new_D4327_ & ~new_D4363_;
  assign new_D4361_ = new_D4310_ | new_D4327_;
  assign new_D4362_ = new_D4310_ | new_D4311_;
  assign new_D4363_ = new_D4327_ & new_D4364_;
  assign new_D4364_ = ~new_D4309_ | ~new_D4334_;
  assign new_D4365_ = new_D4342_ & new_D4362_;
  assign new_D4366_ = ~new_D4342_ & ~new_D4362_;
  assign new_D4367_ = new_D4371_ | new_D4372_;
  assign new_D4368_ = ~new_D4313_ & new_D4327_;
  assign new_D4369_ = new_D4373_ | new_D4374_;
  assign new_D4370_ = new_D4313_ & new_D4327_;
  assign new_D4371_ = ~new_D4313_ & ~new_D4327_;
  assign new_D4372_ = new_D4313_ & ~new_D4327_;
  assign new_D4373_ = new_D4313_ & ~new_D4327_;
  assign new_D4374_ = ~new_D4313_ & new_D4327_;
  assign new_D4375_ = new_F266_;
  assign new_D4376_ = new_F333_;
  assign new_D4377_ = new_F400_;
  assign new_D4378_ = new_F467_;
  assign new_D4379_ = new_F534_;
  assign new_D4380_ = new_F601_;
  assign new_D4381_ = new_D4388_ & new_D4387_;
  assign new_D4382_ = new_D4390_ | new_D4389_;
  assign new_D4383_ = new_D4392_ | new_D4391_;
  assign new_D4384_ = new_D4394_ & new_D4393_;
  assign new_D4385_ = new_D4394_ & new_D4395_;
  assign new_D4386_ = new_D4387_ | new_D4396_;
  assign new_D4387_ = new_D4376_ | new_D4399_;
  assign new_D4388_ = new_D4398_ | new_D4397_;
  assign new_D4389_ = new_D4403_ & new_D4402_;
  assign new_D4390_ = new_D4401_ & new_D4400_;
  assign new_D4391_ = new_D4406_ | new_D4405_;
  assign new_D4392_ = new_D4401_ & new_D4404_;
  assign new_D4393_ = new_D4376_ | new_D4409_;
  assign new_D4394_ = new_D4408_ | new_D4407_;
  assign new_D4395_ = new_D4411_ | new_D4410_;
  assign new_D4396_ = ~new_D4387_ & new_D4413_;
  assign new_D4397_ = ~new_D4389_ & new_D4401_;
  assign new_D4398_ = new_D4389_ & ~new_D4401_;
  assign new_D4399_ = new_D4375_ & ~new_D4376_;
  assign new_D4400_ = ~new_D4422_ | ~new_D4423_;
  assign new_D4401_ = new_D4415_ | new_D4417_;
  assign new_D4402_ = new_D4425_ | new_D4424_;
  assign new_D4403_ = new_D4419_ | new_D4418_;
  assign new_D4404_ = ~new_D4427_ | ~new_D4426_;
  assign new_D4405_ = ~new_D4428_ & new_D4429_;
  assign new_D4406_ = new_D4428_ & ~new_D4429_;
  assign new_D4407_ = ~new_D4375_ & new_D4376_;
  assign new_D4408_ = new_D4375_ & ~new_D4376_;
  assign new_D4409_ = ~new_D4391_ | new_D4401_;
  assign new_D4410_ = new_D4391_ & new_D4401_;
  assign new_D4411_ = ~new_D4391_ & ~new_D4401_;
  assign new_D4412_ = new_D4433_ | new_D4432_;
  assign new_D4413_ = new_D4379_ | new_D4412_;
  assign new_D4414_ = new_D4437_ | new_D4436_;
  assign new_D4415_ = ~new_D4379_ & new_D4414_;
  assign new_D4416_ = new_D4435_ | new_D4434_;
  assign new_D4417_ = new_D4379_ & new_D4416_;
  assign new_D4418_ = new_D4377_ & ~new_D4387_;
  assign new_D4419_ = ~new_D4377_ & new_D4387_;
  assign new_D4420_ = ~new_D4376_ | ~new_D4401_;
  assign new_D4421_ = new_D4387_ & new_D4420_;
  assign new_D4422_ = ~new_D4387_ & ~new_D4421_;
  assign new_D4423_ = new_D4387_ | new_D4420_;
  assign new_D4424_ = ~new_D4377_ & new_D4378_;
  assign new_D4425_ = new_D4377_ & ~new_D4378_;
  assign new_D4426_ = new_D4394_ | new_D4431_;
  assign new_D4427_ = ~new_D4394_ & ~new_D4430_;
  assign new_D4428_ = new_D4377_ | new_D4394_;
  assign new_D4429_ = new_D4377_ | new_D4378_;
  assign new_D4430_ = new_D4394_ & new_D4431_;
  assign new_D4431_ = ~new_D4376_ | ~new_D4401_;
  assign new_D4432_ = new_D4409_ & new_D4429_;
  assign new_D4433_ = ~new_D4409_ & ~new_D4429_;
  assign new_D4434_ = new_D4438_ | new_D4439_;
  assign new_D4435_ = ~new_D4380_ & new_D4394_;
  assign new_D4436_ = new_D4440_ | new_D4441_;
  assign new_D4437_ = new_D4380_ & new_D4394_;
  assign new_D4438_ = ~new_D4380_ & ~new_D4394_;
  assign new_D4439_ = new_D4380_ & ~new_D4394_;
  assign new_D4440_ = new_D4380_ & ~new_D4394_;
  assign new_D4441_ = ~new_D4380_ & new_D4394_;
  assign new_D4442_ = new_F668_;
  assign new_D4443_ = new_F735_;
  assign new_D4444_ = new_F802_;
  assign new_D4445_ = new_F869_;
  assign new_D4446_ = new_F936_;
  assign new_D4447_ = new_F1003_;
  assign new_D4448_ = new_D4455_ & new_D4454_;
  assign new_D4449_ = new_D4457_ | new_D4456_;
  assign new_D4450_ = new_D4459_ | new_D4458_;
  assign new_D4451_ = new_D4461_ & new_D4460_;
  assign new_D4452_ = new_D4461_ & new_D4462_;
  assign new_D4453_ = new_D4454_ | new_D4463_;
  assign new_D4454_ = new_D4443_ | new_D4466_;
  assign new_D4455_ = new_D4465_ | new_D4464_;
  assign new_D4456_ = new_D4470_ & new_D4469_;
  assign new_D4457_ = new_D4468_ & new_D4467_;
  assign new_D4458_ = new_D4473_ | new_D4472_;
  assign new_D4459_ = new_D4468_ & new_D4471_;
  assign new_D4460_ = new_D4443_ | new_D4476_;
  assign new_D4461_ = new_D4475_ | new_D4474_;
  assign new_D4462_ = new_D4478_ | new_D4477_;
  assign new_D4463_ = ~new_D4454_ & new_D4480_;
  assign new_D4464_ = ~new_D4456_ & new_D4468_;
  assign new_D4465_ = new_D4456_ & ~new_D4468_;
  assign new_D4466_ = new_D4442_ & ~new_D4443_;
  assign new_D4467_ = ~new_D4489_ | ~new_D4490_;
  assign new_D4468_ = new_D4482_ | new_D4484_;
  assign new_D4469_ = new_D4492_ | new_D4491_;
  assign new_D4470_ = new_D4486_ | new_D4485_;
  assign new_D4471_ = ~new_D4494_ | ~new_D4493_;
  assign new_D4472_ = ~new_D4495_ & new_D4496_;
  assign new_D4473_ = new_D4495_ & ~new_D4496_;
  assign new_D4474_ = ~new_D4442_ & new_D4443_;
  assign new_D4475_ = new_D4442_ & ~new_D4443_;
  assign new_D4476_ = ~new_D4458_ | new_D4468_;
  assign new_D4477_ = new_D4458_ & new_D4468_;
  assign new_D4478_ = ~new_D4458_ & ~new_D4468_;
  assign new_D4479_ = new_D4500_ | new_D4499_;
  assign new_D4480_ = new_D4446_ | new_D4479_;
  assign new_D4481_ = new_D4504_ | new_D4503_;
  assign new_D4482_ = ~new_D4446_ & new_D4481_;
  assign new_D4483_ = new_D4502_ | new_D4501_;
  assign new_D4484_ = new_D4446_ & new_D4483_;
  assign new_D4485_ = new_D4444_ & ~new_D4454_;
  assign new_D4486_ = ~new_D4444_ & new_D4454_;
  assign new_D4487_ = ~new_D4443_ | ~new_D4468_;
  assign new_D4488_ = new_D4454_ & new_D4487_;
  assign new_D4489_ = ~new_D4454_ & ~new_D4488_;
  assign new_D4490_ = new_D4454_ | new_D4487_;
  assign new_D4491_ = ~new_D4444_ & new_D4445_;
  assign new_D4492_ = new_D4444_ & ~new_D4445_;
  assign new_D4493_ = new_D4461_ | new_D4498_;
  assign new_D4494_ = ~new_D4461_ & ~new_D4497_;
  assign new_D4495_ = new_D4444_ | new_D4461_;
  assign new_D4496_ = new_D4444_ | new_D4445_;
  assign new_D4497_ = new_D4461_ & new_D4498_;
  assign new_D4498_ = ~new_D4443_ | ~new_D4468_;
  assign new_D4499_ = new_D4476_ & new_D4496_;
  assign new_D4500_ = ~new_D4476_ & ~new_D4496_;
  assign new_D4501_ = new_D4505_ | new_D4506_;
  assign new_D4502_ = ~new_D4447_ & new_D4461_;
  assign new_D4503_ = new_D4507_ | new_D4508_;
  assign new_D4504_ = new_D4447_ & new_D4461_;
  assign new_D4505_ = ~new_D4447_ & ~new_D4461_;
  assign new_D4506_ = new_D4447_ & ~new_D4461_;
  assign new_D4507_ = new_D4447_ & ~new_D4461_;
  assign new_D4508_ = ~new_D4447_ & new_D4461_;
  assign new_D4509_ = new_F1070_;
  assign new_D4510_ = new_F1137_;
  assign new_D4511_ = new_F1204_;
  assign new_D4512_ = new_F1271_;
  assign new_D4513_ = new_F1338_;
  assign new_D4514_ = new_F1405_;
  assign new_D4515_ = new_D4522_ & new_D4521_;
  assign new_D4516_ = new_D4524_ | new_D4523_;
  assign new_D4517_ = new_D4526_ | new_D4525_;
  assign new_D4518_ = new_D4528_ & new_D4527_;
  assign new_D4519_ = new_D4528_ & new_D4529_;
  assign new_D4520_ = new_D4521_ | new_D4530_;
  assign new_D4521_ = new_D4510_ | new_D4533_;
  assign new_D4522_ = new_D4532_ | new_D4531_;
  assign new_D4523_ = new_D4537_ & new_D4536_;
  assign new_D4524_ = new_D4535_ & new_D4534_;
  assign new_D4525_ = new_D4540_ | new_D4539_;
  assign new_D4526_ = new_D4535_ & new_D4538_;
  assign new_D4527_ = new_D4510_ | new_D4543_;
  assign new_D4528_ = new_D4542_ | new_D4541_;
  assign new_D4529_ = new_D4545_ | new_D4544_;
  assign new_D4530_ = ~new_D4521_ & new_D4547_;
  assign new_D4531_ = ~new_D4523_ & new_D4535_;
  assign new_D4532_ = new_D4523_ & ~new_D4535_;
  assign new_D4533_ = new_D4509_ & ~new_D4510_;
  assign new_D4534_ = ~new_D4556_ | ~new_D4557_;
  assign new_D4535_ = new_D4549_ | new_D4551_;
  assign new_D4536_ = new_D4559_ | new_D4558_;
  assign new_D4537_ = new_D4553_ | new_D4552_;
  assign new_D4538_ = ~new_D4561_ | ~new_D4560_;
  assign new_D4539_ = ~new_D4562_ & new_D4563_;
  assign new_D4540_ = new_D4562_ & ~new_D4563_;
  assign new_D4541_ = ~new_D4509_ & new_D4510_;
  assign new_D4542_ = new_D4509_ & ~new_D4510_;
  assign new_D4543_ = ~new_D4525_ | new_D4535_;
  assign new_D4544_ = new_D4525_ & new_D4535_;
  assign new_D4545_ = ~new_D4525_ & ~new_D4535_;
  assign new_D4546_ = new_D4567_ | new_D4566_;
  assign new_D4547_ = new_D4513_ | new_D4546_;
  assign new_D4548_ = new_D4571_ | new_D4570_;
  assign new_D4549_ = ~new_D4513_ & new_D4548_;
  assign new_D4550_ = new_D4569_ | new_D4568_;
  assign new_D4551_ = new_D4513_ & new_D4550_;
  assign new_D4552_ = new_D4511_ & ~new_D4521_;
  assign new_D4553_ = ~new_D4511_ & new_D4521_;
  assign new_D4554_ = ~new_D4510_ | ~new_D4535_;
  assign new_D4555_ = new_D4521_ & new_D4554_;
  assign new_D4556_ = ~new_D4521_ & ~new_D4555_;
  assign new_D4557_ = new_D4521_ | new_D4554_;
  assign new_D4558_ = ~new_D4511_ & new_D4512_;
  assign new_D4559_ = new_D4511_ & ~new_D4512_;
  assign new_D4560_ = new_D4528_ | new_D4565_;
  assign new_D4561_ = ~new_D4528_ & ~new_D4564_;
  assign new_D4562_ = new_D4511_ | new_D4528_;
  assign new_D4563_ = new_D4511_ | new_D4512_;
  assign new_D4564_ = new_D4528_ & new_D4565_;
  assign new_D4565_ = ~new_D4510_ | ~new_D4535_;
  assign new_D4566_ = new_D4543_ & new_D4563_;
  assign new_D4567_ = ~new_D4543_ & ~new_D4563_;
  assign new_D4568_ = new_D4572_ | new_D4573_;
  assign new_D4569_ = ~new_D4514_ & new_D4528_;
  assign new_D4570_ = new_D4574_ | new_D4575_;
  assign new_D4571_ = new_D4514_ & new_D4528_;
  assign new_D4572_ = ~new_D4514_ & ~new_D4528_;
  assign new_D4573_ = new_D4514_ & ~new_D4528_;
  assign new_D4574_ = new_D4514_ & ~new_D4528_;
  assign new_D4575_ = ~new_D4514_ & new_D4528_;
  assign new_D4576_ = new_D6994_;
  assign new_D4577_ = new_D7066_;
  assign new_D4578_ = new_D7133_;
  assign new_D4579_ = new_D7200_;
  assign new_D4580_ = new_D7267_;
  assign new_D4581_ = new_D7334_;
  assign new_D4582_ = new_D4589_ & new_D4588_;
  assign new_D4583_ = new_D4591_ | new_D4590_;
  assign new_D4584_ = new_D4593_ | new_D4592_;
  assign new_D4585_ = new_D4595_ & new_D4594_;
  assign new_D4586_ = new_D4595_ & new_D4596_;
  assign new_D4587_ = new_D4588_ | new_D4597_;
  assign new_D4588_ = new_D4577_ | new_D4600_;
  assign new_D4589_ = new_D4599_ | new_D4598_;
  assign new_D4590_ = new_D4604_ & new_D4603_;
  assign new_D4591_ = new_D4602_ & new_D4601_;
  assign new_D4592_ = new_D4607_ | new_D4606_;
  assign new_D4593_ = new_D4602_ & new_D4605_;
  assign new_D4594_ = new_D4577_ | new_D4610_;
  assign new_D4595_ = new_D4609_ | new_D4608_;
  assign new_D4596_ = new_D4612_ | new_D4611_;
  assign new_D4597_ = ~new_D4588_ & new_D4614_;
  assign new_D4598_ = ~new_D4590_ & new_D4602_;
  assign new_D4599_ = new_D4590_ & ~new_D4602_;
  assign new_D4600_ = new_D4576_ & ~new_D4577_;
  assign new_D4601_ = ~new_D4623_ | ~new_D4624_;
  assign new_D4602_ = new_D4616_ | new_D4618_;
  assign new_D4603_ = new_D4626_ | new_D4625_;
  assign new_D4604_ = new_D4620_ | new_D4619_;
  assign new_D4605_ = ~new_D4628_ | ~new_D4627_;
  assign new_D4606_ = ~new_D4629_ & new_D4630_;
  assign new_D4607_ = new_D4629_ & ~new_D4630_;
  assign new_D4608_ = ~new_D4576_ & new_D4577_;
  assign new_D4609_ = new_D4576_ & ~new_D4577_;
  assign new_D4610_ = ~new_D4592_ | new_D4602_;
  assign new_D4611_ = new_D4592_ & new_D4602_;
  assign new_D4612_ = ~new_D4592_ & ~new_D4602_;
  assign new_D4613_ = new_D4634_ | new_D4633_;
  assign new_D4614_ = new_D4580_ | new_D4613_;
  assign new_D4615_ = new_D4638_ | new_D4637_;
  assign new_D4616_ = ~new_D4580_ & new_D4615_;
  assign new_D4617_ = new_D4636_ | new_D4635_;
  assign new_D4618_ = new_D4580_ & new_D4617_;
  assign new_D4619_ = new_D4578_ & ~new_D4588_;
  assign new_D4620_ = ~new_D4578_ & new_D4588_;
  assign new_D4621_ = ~new_D4577_ | ~new_D4602_;
  assign new_D4622_ = new_D4588_ & new_D4621_;
  assign new_D4623_ = ~new_D4588_ & ~new_D4622_;
  assign new_D4624_ = new_D4588_ | new_D4621_;
  assign new_D4625_ = ~new_D4578_ & new_D4579_;
  assign new_D4626_ = new_D4578_ & ~new_D4579_;
  assign new_D4627_ = new_D4595_ | new_D4632_;
  assign new_D4628_ = ~new_D4595_ & ~new_D4631_;
  assign new_D4629_ = new_D4578_ | new_D4595_;
  assign new_D4630_ = new_D4578_ | new_D4579_;
  assign new_D4631_ = new_D4595_ & new_D4632_;
  assign new_D4632_ = ~new_D4577_ | ~new_D4602_;
  assign new_D4633_ = new_D4610_ & new_D4630_;
  assign new_D4634_ = ~new_D4610_ & ~new_D4630_;
  assign new_D4635_ = new_D4639_ | new_D4640_;
  assign new_D4636_ = ~new_D4581_ & new_D4595_;
  assign new_D4637_ = new_D4641_ | new_D4642_;
  assign new_D4638_ = new_D4581_ & new_D4595_;
  assign new_D4639_ = ~new_D4581_ & ~new_D4595_;
  assign new_D4640_ = new_D4581_ & ~new_D4595_;
  assign new_D4641_ = new_D4581_ & ~new_D4595_;
  assign new_D4642_ = ~new_D4581_ & new_D4595_;
  assign new_D4643_ = new_D7401_;
  assign new_D4644_ = new_D7468_;
  assign new_D4645_ = new_D7535_;
  assign new_D4646_ = new_D7602_;
  assign new_D4647_ = new_D7669_;
  assign new_D4648_ = new_D7736_;
  assign new_D4649_ = new_D4656_ & new_D4655_;
  assign new_D4650_ = new_D4658_ | new_D4657_;
  assign new_D4651_ = new_D4660_ | new_D4659_;
  assign new_D4652_ = new_D4662_ & new_D4661_;
  assign new_D4653_ = new_D4662_ & new_D4663_;
  assign new_D4654_ = new_D4655_ | new_D4664_;
  assign new_D4655_ = new_D4644_ | new_D4667_;
  assign new_D4656_ = new_D4666_ | new_D4665_;
  assign new_D4657_ = new_D4671_ & new_D4670_;
  assign new_D4658_ = new_D4669_ & new_D4668_;
  assign new_D4659_ = new_D4674_ | new_D4673_;
  assign new_D4660_ = new_D4669_ & new_D4672_;
  assign new_D4661_ = new_D4644_ | new_D4677_;
  assign new_D4662_ = new_D4676_ | new_D4675_;
  assign new_D4663_ = new_D4679_ | new_D4678_;
  assign new_D4664_ = ~new_D4655_ & new_D4681_;
  assign new_D4665_ = ~new_D4657_ & new_D4669_;
  assign new_D4666_ = new_D4657_ & ~new_D4669_;
  assign new_D4667_ = new_D4643_ & ~new_D4644_;
  assign new_D4668_ = ~new_D4690_ | ~new_D4691_;
  assign new_D4669_ = new_D4683_ | new_D4685_;
  assign new_D4670_ = new_D4693_ | new_D4692_;
  assign new_D4671_ = new_D4687_ | new_D4686_;
  assign new_D4672_ = ~new_D4695_ | ~new_D4694_;
  assign new_D4673_ = ~new_D4696_ & new_D4697_;
  assign new_D4674_ = new_D4696_ & ~new_D4697_;
  assign new_D4675_ = ~new_D4643_ & new_D4644_;
  assign new_D4676_ = new_D4643_ & ~new_D4644_;
  assign new_D4677_ = ~new_D4659_ | new_D4669_;
  assign new_D4678_ = new_D4659_ & new_D4669_;
  assign new_D4679_ = ~new_D4659_ & ~new_D4669_;
  assign new_D4680_ = new_D4701_ | new_D4700_;
  assign new_D4681_ = new_D4647_ | new_D4680_;
  assign new_D4682_ = new_D4705_ | new_D4704_;
  assign new_D4683_ = ~new_D4647_ & new_D4682_;
  assign new_D4684_ = new_D4703_ | new_D4702_;
  assign new_D4685_ = new_D4647_ & new_D4684_;
  assign new_D4686_ = new_D4645_ & ~new_D4655_;
  assign new_D4687_ = ~new_D4645_ & new_D4655_;
  assign new_D4688_ = ~new_D4644_ | ~new_D4669_;
  assign new_D4689_ = new_D4655_ & new_D4688_;
  assign new_D4690_ = ~new_D4655_ & ~new_D4689_;
  assign new_D4691_ = new_D4655_ | new_D4688_;
  assign new_D4692_ = ~new_D4645_ & new_D4646_;
  assign new_D4693_ = new_D4645_ & ~new_D4646_;
  assign new_D4694_ = new_D4662_ | new_D4699_;
  assign new_D4695_ = ~new_D4662_ & ~new_D4698_;
  assign new_D4696_ = new_D4645_ | new_D4662_;
  assign new_D4697_ = new_D4645_ | new_D4646_;
  assign new_D4698_ = new_D4662_ & new_D4699_;
  assign new_D4699_ = ~new_D4644_ | ~new_D4669_;
  assign new_D4700_ = new_D4677_ & new_D4697_;
  assign new_D4701_ = ~new_D4677_ & ~new_D4697_;
  assign new_D4702_ = new_D4706_ | new_D4707_;
  assign new_D4703_ = ~new_D4648_ & new_D4662_;
  assign new_D4704_ = new_D4708_ | new_D4709_;
  assign new_D4705_ = new_D4648_ & new_D4662_;
  assign new_D4706_ = ~new_D4648_ & ~new_D4662_;
  assign new_D4707_ = new_D4648_ & ~new_D4662_;
  assign new_D4708_ = new_D4648_ & ~new_D4662_;
  assign new_D4709_ = ~new_D4648_ & new_D4662_;
  assign new_D4710_ = new_D7803_;
  assign new_D4711_ = new_D7870_;
  assign new_D4712_ = new_D7937_;
  assign new_D4713_ = new_D8004_;
  assign new_D4714_ = new_D8071_;
  assign new_D4715_ = new_D8138_;
  assign new_D4716_ = new_D4723_ & new_D4722_;
  assign new_D4717_ = new_D4725_ | new_D4724_;
  assign new_D4718_ = new_D4727_ | new_D4726_;
  assign new_D4719_ = new_D4729_ & new_D4728_;
  assign new_D4720_ = new_D4729_ & new_D4730_;
  assign new_D4721_ = new_D4722_ | new_D4731_;
  assign new_D4722_ = new_D4711_ | new_D4734_;
  assign new_D4723_ = new_D4733_ | new_D4732_;
  assign new_D4724_ = new_D4738_ & new_D4737_;
  assign new_D4725_ = new_D4736_ & new_D4735_;
  assign new_D4726_ = new_D4741_ | new_D4740_;
  assign new_D4727_ = new_D4736_ & new_D4739_;
  assign new_D4728_ = new_D4711_ | new_D4744_;
  assign new_D4729_ = new_D4743_ | new_D4742_;
  assign new_D4730_ = new_D4746_ | new_D4745_;
  assign new_D4731_ = ~new_D4722_ & new_D4748_;
  assign new_D4732_ = ~new_D4724_ & new_D4736_;
  assign new_D4733_ = new_D4724_ & ~new_D4736_;
  assign new_D4734_ = new_D4710_ & ~new_D4711_;
  assign new_D4735_ = ~new_D4757_ | ~new_D4758_;
  assign new_D4736_ = new_D4750_ | new_D4752_;
  assign new_D4737_ = new_D4760_ | new_D4759_;
  assign new_D4738_ = new_D4754_ | new_D4753_;
  assign new_D4739_ = ~new_D4762_ | ~new_D4761_;
  assign new_D4740_ = ~new_D4763_ & new_D4764_;
  assign new_D4741_ = new_D4763_ & ~new_D4764_;
  assign new_D4742_ = ~new_D4710_ & new_D4711_;
  assign new_D4743_ = new_D4710_ & ~new_D4711_;
  assign new_D4744_ = ~new_D4726_ | new_D4736_;
  assign new_D4745_ = new_D4726_ & new_D4736_;
  assign new_D4746_ = ~new_D4726_ & ~new_D4736_;
  assign new_D4747_ = new_D4768_ | new_D4767_;
  assign new_D4748_ = new_D4714_ | new_D4747_;
  assign new_D4749_ = new_D4772_ | new_D4771_;
  assign new_D4750_ = ~new_D4714_ & new_D4749_;
  assign new_D4751_ = new_D4770_ | new_D4769_;
  assign new_D4752_ = new_D4714_ & new_D4751_;
  assign new_D4753_ = new_D4712_ & ~new_D4722_;
  assign new_D4754_ = ~new_D4712_ & new_D4722_;
  assign new_D4755_ = ~new_D4711_ | ~new_D4736_;
  assign new_D4756_ = new_D4722_ & new_D4755_;
  assign new_D4757_ = ~new_D4722_ & ~new_D4756_;
  assign new_D4758_ = new_D4722_ | new_D4755_;
  assign new_D4759_ = ~new_D4712_ & new_D4713_;
  assign new_D4760_ = new_D4712_ & ~new_D4713_;
  assign new_D4761_ = new_D4729_ | new_D4766_;
  assign new_D4762_ = ~new_D4729_ & ~new_D4765_;
  assign new_D4763_ = new_D4712_ | new_D4729_;
  assign new_D4764_ = new_D4712_ | new_D4713_;
  assign new_D4765_ = new_D4729_ & new_D4766_;
  assign new_D4766_ = ~new_D4711_ | ~new_D4736_;
  assign new_D4767_ = new_D4744_ & new_D4764_;
  assign new_D4768_ = ~new_D4744_ & ~new_D4764_;
  assign new_D4769_ = new_D4773_ | new_D4774_;
  assign new_D4770_ = ~new_D4715_ & new_D4729_;
  assign new_D4771_ = new_D4775_ | new_D4776_;
  assign new_D4772_ = new_D4715_ & new_D4729_;
  assign new_D4773_ = ~new_D4715_ & ~new_D4729_;
  assign new_D4774_ = new_D4715_ & ~new_D4729_;
  assign new_D4775_ = new_D4715_ & ~new_D4729_;
  assign new_D4776_ = ~new_D4715_ & new_D4729_;
  assign new_D4777_ = new_D8205_;
  assign new_D4778_ = new_D8272_;
  assign new_D4779_ = new_D8339_;
  assign new_D4780_ = new_D8406_;
  assign new_D4781_ = new_D8473_;
  assign new_D4782_ = new_D8540_;
  assign new_D4783_ = new_D4790_ & new_D4789_;
  assign new_D4784_ = new_D4792_ | new_D4791_;
  assign new_D4785_ = new_D4794_ | new_D4793_;
  assign new_D4786_ = new_D4796_ & new_D4795_;
  assign new_D4787_ = new_D4796_ & new_D4797_;
  assign new_D4788_ = new_D4789_ | new_D4798_;
  assign new_D4789_ = new_D4778_ | new_D4801_;
  assign new_D4790_ = new_D4800_ | new_D4799_;
  assign new_D4791_ = new_D4805_ & new_D4804_;
  assign new_D4792_ = new_D4803_ & new_D4802_;
  assign new_D4793_ = new_D4808_ | new_D4807_;
  assign new_D4794_ = new_D4803_ & new_D4806_;
  assign new_D4795_ = new_D4778_ | new_D4811_;
  assign new_D4796_ = new_D4810_ | new_D4809_;
  assign new_D4797_ = new_D4813_ | new_D4812_;
  assign new_D4798_ = ~new_D4789_ & new_D4815_;
  assign new_D4799_ = ~new_D4791_ & new_D4803_;
  assign new_D4800_ = new_D4791_ & ~new_D4803_;
  assign new_D4801_ = new_D4777_ & ~new_D4778_;
  assign new_D4802_ = ~new_D4824_ | ~new_D4825_;
  assign new_D4803_ = new_D4817_ | new_D4819_;
  assign new_D4804_ = new_D4827_ | new_D4826_;
  assign new_D4805_ = new_D4821_ | new_D4820_;
  assign new_D4806_ = ~new_D4829_ | ~new_D4828_;
  assign new_D4807_ = ~new_D4830_ & new_D4831_;
  assign new_D4808_ = new_D4830_ & ~new_D4831_;
  assign new_D4809_ = ~new_D4777_ & new_D4778_;
  assign new_D4810_ = new_D4777_ & ~new_D4778_;
  assign new_D4811_ = ~new_D4793_ | new_D4803_;
  assign new_D4812_ = new_D4793_ & new_D4803_;
  assign new_D4813_ = ~new_D4793_ & ~new_D4803_;
  assign new_D4814_ = new_D4835_ | new_D4834_;
  assign new_D4815_ = new_D4781_ | new_D4814_;
  assign new_D4816_ = new_D4839_ | new_D4838_;
  assign new_D4817_ = ~new_D4781_ & new_D4816_;
  assign new_D4818_ = new_D4837_ | new_D4836_;
  assign new_D4819_ = new_D4781_ & new_D4818_;
  assign new_D4820_ = new_D4779_ & ~new_D4789_;
  assign new_D4821_ = ~new_D4779_ & new_D4789_;
  assign new_D4822_ = ~new_D4778_ | ~new_D4803_;
  assign new_D4823_ = new_D4789_ & new_D4822_;
  assign new_D4824_ = ~new_D4789_ & ~new_D4823_;
  assign new_D4825_ = new_D4789_ | new_D4822_;
  assign new_D4826_ = ~new_D4779_ & new_D4780_;
  assign new_D4827_ = new_D4779_ & ~new_D4780_;
  assign new_D4828_ = new_D4796_ | new_D4833_;
  assign new_D4829_ = ~new_D4796_ & ~new_D4832_;
  assign new_D4830_ = new_D4779_ | new_D4796_;
  assign new_D4831_ = new_D4779_ | new_D4780_;
  assign new_D4832_ = new_D4796_ & new_D4833_;
  assign new_D4833_ = ~new_D4778_ | ~new_D4803_;
  assign new_D4834_ = new_D4811_ & new_D4831_;
  assign new_D4835_ = ~new_D4811_ & ~new_D4831_;
  assign new_D4836_ = new_D4840_ | new_D4841_;
  assign new_D4837_ = ~new_D4782_ & new_D4796_;
  assign new_D4838_ = new_D4842_ | new_D4843_;
  assign new_D4839_ = new_D4782_ & new_D4796_;
  assign new_D4840_ = ~new_D4782_ & ~new_D4796_;
  assign new_D4841_ = new_D4782_ & ~new_D4796_;
  assign new_D4842_ = new_D4782_ & ~new_D4796_;
  assign new_D4843_ = ~new_D4782_ & new_D4796_;
  assign new_D4844_ = new_D8607_;
  assign new_D4845_ = new_D8674_;
  assign new_D4846_ = new_D8741_;
  assign new_D4847_ = new_D8808_;
  assign new_D4848_ = new_D8875_;
  assign new_D4849_ = new_D8942_;
  assign new_D4850_ = new_D4857_ & new_D4856_;
  assign new_D4851_ = new_D4859_ | new_D4858_;
  assign new_D4852_ = new_D4861_ | new_D4860_;
  assign new_D4853_ = new_D4863_ & new_D4862_;
  assign new_D4854_ = new_D4863_ & new_D4864_;
  assign new_D4855_ = new_D4856_ | new_D4865_;
  assign new_D4856_ = new_D4845_ | new_D4868_;
  assign new_D4857_ = new_D4867_ | new_D4866_;
  assign new_D4858_ = new_D4872_ & new_D4871_;
  assign new_D4859_ = new_D4870_ & new_D4869_;
  assign new_D4860_ = new_D4875_ | new_D4874_;
  assign new_D4861_ = new_D4870_ & new_D4873_;
  assign new_D4862_ = new_D4845_ | new_D4878_;
  assign new_D4863_ = new_D4877_ | new_D4876_;
  assign new_D4864_ = new_D4880_ | new_D4879_;
  assign new_D4865_ = ~new_D4856_ & new_D4882_;
  assign new_D4866_ = ~new_D4858_ & new_D4870_;
  assign new_D4867_ = new_D4858_ & ~new_D4870_;
  assign new_D4868_ = new_D4844_ & ~new_D4845_;
  assign new_D4869_ = ~new_D4891_ | ~new_D4892_;
  assign new_D4870_ = new_D4884_ | new_D4886_;
  assign new_D4871_ = new_D4894_ | new_D4893_;
  assign new_D4872_ = new_D4888_ | new_D4887_;
  assign new_D4873_ = ~new_D4896_ | ~new_D4895_;
  assign new_D4874_ = ~new_D4897_ & new_D4898_;
  assign new_D4875_ = new_D4897_ & ~new_D4898_;
  assign new_D4876_ = ~new_D4844_ & new_D4845_;
  assign new_D4877_ = new_D4844_ & ~new_D4845_;
  assign new_D4878_ = ~new_D4860_ | new_D4870_;
  assign new_D4879_ = new_D4860_ & new_D4870_;
  assign new_D4880_ = ~new_D4860_ & ~new_D4870_;
  assign new_D4881_ = new_D4902_ | new_D4901_;
  assign new_D4882_ = new_D4848_ | new_D4881_;
  assign new_D4883_ = new_D4906_ | new_D4905_;
  assign new_D4884_ = ~new_D4848_ & new_D4883_;
  assign new_D4885_ = new_D4904_ | new_D4903_;
  assign new_D4886_ = new_D4848_ & new_D4885_;
  assign new_D4887_ = new_D4846_ & ~new_D4856_;
  assign new_D4888_ = ~new_D4846_ & new_D4856_;
  assign new_D4889_ = ~new_D4845_ | ~new_D4870_;
  assign new_D4890_ = new_D4856_ & new_D4889_;
  assign new_D4891_ = ~new_D4856_ & ~new_D4890_;
  assign new_D4892_ = new_D4856_ | new_D4889_;
  assign new_D4893_ = ~new_D4846_ & new_D4847_;
  assign new_D4894_ = new_D4846_ & ~new_D4847_;
  assign new_D4895_ = new_D4863_ | new_D4900_;
  assign new_D4896_ = ~new_D4863_ & ~new_D4899_;
  assign new_D4897_ = new_D4846_ | new_D4863_;
  assign new_D4898_ = new_D4846_ | new_D4847_;
  assign new_D4899_ = new_D4863_ & new_D4900_;
  assign new_D4900_ = ~new_D4845_ | ~new_D4870_;
  assign new_D4901_ = new_D4878_ & new_D4898_;
  assign new_D4902_ = ~new_D4878_ & ~new_D4898_;
  assign new_D4903_ = new_D4907_ | new_D4908_;
  assign new_D4904_ = ~new_D4849_ & new_D4863_;
  assign new_D4905_ = new_D4909_ | new_D4910_;
  assign new_D4906_ = new_D4849_ & new_D4863_;
  assign new_D4907_ = ~new_D4849_ & ~new_D4863_;
  assign new_D4908_ = new_D4849_ & ~new_D4863_;
  assign new_D4909_ = new_D4849_ & ~new_D4863_;
  assign new_D4910_ = ~new_D4849_ & new_D4863_;
  assign new_D4911_ = new_D9009_;
  assign new_D4912_ = new_D9076_;
  assign new_D4913_ = new_D9143_;
  assign new_D4914_ = new_D9210_;
  assign new_D4915_ = new_D9277_;
  assign new_D4916_ = new_D9344_;
  assign new_D4917_ = new_D4924_ & new_D4923_;
  assign new_D4918_ = new_D4926_ | new_D4925_;
  assign new_D4919_ = new_D4928_ | new_D4927_;
  assign new_D4920_ = new_D4930_ & new_D4929_;
  assign new_D4921_ = new_D4930_ & new_D4931_;
  assign new_D4922_ = new_D4923_ | new_D4932_;
  assign new_D4923_ = new_D4912_ | new_D4935_;
  assign new_D4924_ = new_D4934_ | new_D4933_;
  assign new_D4925_ = new_D4939_ & new_D4938_;
  assign new_D4926_ = new_D4937_ & new_D4936_;
  assign new_D4927_ = new_D4942_ | new_D4941_;
  assign new_D4928_ = new_D4937_ & new_D4940_;
  assign new_D4929_ = new_D4912_ | new_D4945_;
  assign new_D4930_ = new_D4944_ | new_D4943_;
  assign new_D4931_ = new_D4947_ | new_D4946_;
  assign new_D4932_ = ~new_D4923_ & new_D4949_;
  assign new_D4933_ = ~new_D4925_ & new_D4937_;
  assign new_D4934_ = new_D4925_ & ~new_D4937_;
  assign new_D4935_ = new_D4911_ & ~new_D4912_;
  assign new_D4936_ = ~new_D4958_ | ~new_D4959_;
  assign new_D4937_ = new_D4951_ | new_D4953_;
  assign new_D4938_ = new_D4961_ | new_D4960_;
  assign new_D4939_ = new_D4955_ | new_D4954_;
  assign new_D4940_ = ~new_D4963_ | ~new_D4962_;
  assign new_D4941_ = ~new_D4964_ & new_D4965_;
  assign new_D4942_ = new_D4964_ & ~new_D4965_;
  assign new_D4943_ = ~new_D4911_ & new_D4912_;
  assign new_D4944_ = new_D4911_ & ~new_D4912_;
  assign new_D4945_ = ~new_D4927_ | new_D4937_;
  assign new_D4946_ = new_D4927_ & new_D4937_;
  assign new_D4947_ = ~new_D4927_ & ~new_D4937_;
  assign new_D4948_ = new_D4969_ | new_D4968_;
  assign new_D4949_ = new_D4915_ | new_D4948_;
  assign new_D4950_ = new_D4973_ | new_D4972_;
  assign new_D4951_ = ~new_D4915_ & new_D4950_;
  assign new_D4952_ = new_D4971_ | new_D4970_;
  assign new_D4953_ = new_D4915_ & new_D4952_;
  assign new_D4954_ = new_D4913_ & ~new_D4923_;
  assign new_D4955_ = ~new_D4913_ & new_D4923_;
  assign new_D4956_ = ~new_D4912_ | ~new_D4937_;
  assign new_D4957_ = new_D4923_ & new_D4956_;
  assign new_D4958_ = ~new_D4923_ & ~new_D4957_;
  assign new_D4959_ = new_D4923_ | new_D4956_;
  assign new_D4960_ = ~new_D4913_ & new_D4914_;
  assign new_D4961_ = new_D4913_ & ~new_D4914_;
  assign new_D4962_ = new_D4930_ | new_D4967_;
  assign new_D4963_ = ~new_D4930_ & ~new_D4966_;
  assign new_D4964_ = new_D4913_ | new_D4930_;
  assign new_D4965_ = new_D4913_ | new_D4914_;
  assign new_D4966_ = new_D4930_ & new_D4967_;
  assign new_D4967_ = ~new_D4912_ | ~new_D4937_;
  assign new_D4968_ = new_D4945_ & new_D4965_;
  assign new_D4969_ = ~new_D4945_ & ~new_D4965_;
  assign new_D4970_ = new_D4974_ | new_D4975_;
  assign new_D4971_ = ~new_D4916_ & new_D4930_;
  assign new_D4972_ = new_D4976_ | new_D4977_;
  assign new_D4973_ = new_D4916_ & new_D4930_;
  assign new_D4974_ = ~new_D4916_ & ~new_D4930_;
  assign new_D4975_ = new_D4916_ & ~new_D4930_;
  assign new_D4976_ = new_D4916_ & ~new_D4930_;
  assign new_D4977_ = ~new_D4916_ & new_D4930_;
  assign new_D4978_ = new_D9411_;
  assign new_D4979_ = new_D9478_;
  assign new_D4980_ = new_D9545_;
  assign new_D4981_ = new_D9612_;
  assign new_D4982_ = new_D9679_;
  assign new_D4983_ = new_D9746_;
  assign new_D4984_ = new_D4991_ & new_D4990_;
  assign new_D4985_ = new_D4993_ | new_D4992_;
  assign new_D4986_ = new_D4995_ | new_D4994_;
  assign new_D4987_ = new_D4997_ & new_D4996_;
  assign new_D4988_ = new_D4997_ & new_D4998_;
  assign new_D4989_ = new_D4990_ | new_D4999_;
  assign new_D4990_ = new_D4979_ | new_D5002_;
  assign new_D4991_ = new_D5001_ | new_D5000_;
  assign new_D4992_ = new_D5006_ & new_D5005_;
  assign new_D4993_ = new_D5004_ & new_D5003_;
  assign new_D4994_ = new_D5009_ | new_D5008_;
  assign new_D4995_ = new_D5004_ & new_D5007_;
  assign new_D4996_ = new_D4979_ | new_D5012_;
  assign new_D4997_ = new_D5011_ | new_D5010_;
  assign new_D4998_ = new_D5014_ | new_D5013_;
  assign new_D4999_ = ~new_D4990_ & new_D5016_;
  assign new_D5000_ = ~new_D4992_ & new_D5004_;
  assign new_D5001_ = new_D4992_ & ~new_D5004_;
  assign new_D5002_ = new_D4978_ & ~new_D4979_;
  assign new_D5003_ = ~new_D5025_ | ~new_D5026_;
  assign new_D5004_ = new_D5018_ | new_D5020_;
  assign new_D5005_ = new_D5028_ | new_D5027_;
  assign new_D5006_ = new_D5022_ | new_D5021_;
  assign new_D5007_ = ~new_D5030_ | ~new_D5029_;
  assign new_D5008_ = ~new_D5031_ & new_D5032_;
  assign new_D5009_ = new_D5031_ & ~new_D5032_;
  assign new_D5010_ = ~new_D4978_ & new_D4979_;
  assign new_D5011_ = new_D4978_ & ~new_D4979_;
  assign new_D5012_ = ~new_D4994_ | new_D5004_;
  assign new_D5013_ = new_D4994_ & new_D5004_;
  assign new_D5014_ = ~new_D4994_ & ~new_D5004_;
  assign new_D5015_ = new_D5036_ | new_D5035_;
  assign new_D5016_ = new_D4982_ | new_D5015_;
  assign new_D5017_ = new_D5040_ | new_D5039_;
  assign new_D5018_ = ~new_D4982_ & new_D5017_;
  assign new_D5019_ = new_D5038_ | new_D5037_;
  assign new_D5020_ = new_D4982_ & new_D5019_;
  assign new_D5021_ = new_D4980_ & ~new_D4990_;
  assign new_D5022_ = ~new_D4980_ & new_D4990_;
  assign new_D5023_ = ~new_D4979_ | ~new_D5004_;
  assign new_D5024_ = new_D4990_ & new_D5023_;
  assign new_D5025_ = ~new_D4990_ & ~new_D5024_;
  assign new_D5026_ = new_D4990_ | new_D5023_;
  assign new_D5027_ = ~new_D4980_ & new_D4981_;
  assign new_D5028_ = new_D4980_ & ~new_D4981_;
  assign new_D5029_ = new_D4997_ | new_D5034_;
  assign new_D5030_ = ~new_D4997_ & ~new_D5033_;
  assign new_D5031_ = new_D4980_ | new_D4997_;
  assign new_D5032_ = new_D4980_ | new_D4981_;
  assign new_D5033_ = new_D4997_ & new_D5034_;
  assign new_D5034_ = ~new_D4979_ | ~new_D5004_;
  assign new_D5035_ = new_D5012_ & new_D5032_;
  assign new_D5036_ = ~new_D5012_ & ~new_D5032_;
  assign new_D5037_ = new_D5041_ | new_D5042_;
  assign new_D5038_ = ~new_D4983_ & new_D4997_;
  assign new_D5039_ = new_D5043_ | new_D5044_;
  assign new_D5040_ = new_D4983_ & new_D4997_;
  assign new_D5041_ = ~new_D4983_ & ~new_D4997_;
  assign new_D5042_ = new_D4983_ & ~new_D4997_;
  assign new_D5043_ = new_D4983_ & ~new_D4997_;
  assign new_D5044_ = ~new_D4983_ & new_D4997_;
  assign new_D5045_ = new_D9813_;
  assign new_D5046_ = new_D9880_;
  assign new_D5047_ = new_D9947_;
  assign new_D5048_ = new_E15_;
  assign new_D5049_ = new_E82_;
  assign new_D5050_ = new_E149_;
  assign new_D5051_ = new_D5058_ & new_D5057_;
  assign new_D5052_ = new_D5060_ | new_D5059_;
  assign new_D5053_ = new_D5062_ | new_D5061_;
  assign new_D5054_ = new_D5064_ & new_D5063_;
  assign new_D5055_ = new_D5064_ & new_D5065_;
  assign new_D5056_ = new_D5057_ | new_D5066_;
  assign new_D5057_ = new_D5046_ | new_D5069_;
  assign new_D5058_ = new_D5068_ | new_D5067_;
  assign new_D5059_ = new_D5073_ & new_D5072_;
  assign new_D5060_ = new_D5071_ & new_D5070_;
  assign new_D5061_ = new_D5076_ | new_D5075_;
  assign new_D5062_ = new_D5071_ & new_D5074_;
  assign new_D5063_ = new_D5046_ | new_D5079_;
  assign new_D5064_ = new_D5078_ | new_D5077_;
  assign new_D5065_ = new_D5081_ | new_D5080_;
  assign new_D5066_ = ~new_D5057_ & new_D5083_;
  assign new_D5067_ = ~new_D5059_ & new_D5071_;
  assign new_D5068_ = new_D5059_ & ~new_D5071_;
  assign new_D5069_ = new_D5045_ & ~new_D5046_;
  assign new_D5070_ = ~new_D5092_ | ~new_D5093_;
  assign new_D5071_ = new_D5085_ | new_D5087_;
  assign new_D5072_ = new_D5095_ | new_D5094_;
  assign new_D5073_ = new_D5089_ | new_D5088_;
  assign new_D5074_ = ~new_D5097_ | ~new_D5096_;
  assign new_D5075_ = ~new_D5098_ & new_D5099_;
  assign new_D5076_ = new_D5098_ & ~new_D5099_;
  assign new_D5077_ = ~new_D5045_ & new_D5046_;
  assign new_D5078_ = new_D5045_ & ~new_D5046_;
  assign new_D5079_ = ~new_D5061_ | new_D5071_;
  assign new_D5080_ = new_D5061_ & new_D5071_;
  assign new_D5081_ = ~new_D5061_ & ~new_D5071_;
  assign new_D5082_ = new_D5103_ | new_D5102_;
  assign new_D5083_ = new_D5049_ | new_D5082_;
  assign new_D5084_ = new_D5107_ | new_D5106_;
  assign new_D5085_ = ~new_D5049_ & new_D5084_;
  assign new_D5086_ = new_D5105_ | new_D5104_;
  assign new_D5087_ = new_D5049_ & new_D5086_;
  assign new_D5088_ = new_D5047_ & ~new_D5057_;
  assign new_D5089_ = ~new_D5047_ & new_D5057_;
  assign new_D5090_ = ~new_D5046_ | ~new_D5071_;
  assign new_D5091_ = new_D5057_ & new_D5090_;
  assign new_D5092_ = ~new_D5057_ & ~new_D5091_;
  assign new_D5093_ = new_D5057_ | new_D5090_;
  assign new_D5094_ = ~new_D5047_ & new_D5048_;
  assign new_D5095_ = new_D5047_ & ~new_D5048_;
  assign new_D5096_ = new_D5064_ | new_D5101_;
  assign new_D5097_ = ~new_D5064_ & ~new_D5100_;
  assign new_D5098_ = new_D5047_ | new_D5064_;
  assign new_D5099_ = new_D5047_ | new_D5048_;
  assign new_D5100_ = new_D5064_ & new_D5101_;
  assign new_D5101_ = ~new_D5046_ | ~new_D5071_;
  assign new_D5102_ = new_D5079_ & new_D5099_;
  assign new_D5103_ = ~new_D5079_ & ~new_D5099_;
  assign new_D5104_ = new_D5108_ | new_D5109_;
  assign new_D5105_ = ~new_D5050_ & new_D5064_;
  assign new_D5106_ = new_D5110_ | new_D5111_;
  assign new_D5107_ = new_D5050_ & new_D5064_;
  assign new_D5108_ = ~new_D5050_ & ~new_D5064_;
  assign new_D5109_ = new_D5050_ & ~new_D5064_;
  assign new_D5110_ = new_D5050_ & ~new_D5064_;
  assign new_D5111_ = ~new_D5050_ & new_D5064_;
  assign new_D5112_ = new_E216_;
  assign new_D5113_ = new_E283_;
  assign new_D5114_ = new_E350_;
  assign new_D5115_ = new_E417_;
  assign new_D5116_ = new_E484_;
  assign new_D5117_ = new_E551_;
  assign new_D5118_ = new_D5125_ & new_D5124_;
  assign new_D5119_ = new_D5127_ | new_D5126_;
  assign new_D5120_ = new_D5129_ | new_D5128_;
  assign new_D5121_ = new_D5131_ & new_D5130_;
  assign new_D5122_ = new_D5131_ & new_D5132_;
  assign new_D5123_ = new_D5124_ | new_D5133_;
  assign new_D5124_ = new_D5113_ | new_D5136_;
  assign new_D5125_ = new_D5135_ | new_D5134_;
  assign new_D5126_ = new_D5140_ & new_D5139_;
  assign new_D5127_ = new_D5138_ & new_D5137_;
  assign new_D5128_ = new_D5143_ | new_D5142_;
  assign new_D5129_ = new_D5138_ & new_D5141_;
  assign new_D5130_ = new_D5113_ | new_D5146_;
  assign new_D5131_ = new_D5145_ | new_D5144_;
  assign new_D5132_ = new_D5148_ | new_D5147_;
  assign new_D5133_ = ~new_D5124_ & new_D5150_;
  assign new_D5134_ = ~new_D5126_ & new_D5138_;
  assign new_D5135_ = new_D5126_ & ~new_D5138_;
  assign new_D5136_ = new_D5112_ & ~new_D5113_;
  assign new_D5137_ = ~new_D5159_ | ~new_D5160_;
  assign new_D5138_ = new_D5152_ | new_D5154_;
  assign new_D5139_ = new_D5162_ | new_D5161_;
  assign new_D5140_ = new_D5156_ | new_D5155_;
  assign new_D5141_ = ~new_D5164_ | ~new_D5163_;
  assign new_D5142_ = ~new_D5165_ & new_D5166_;
  assign new_D5143_ = new_D5165_ & ~new_D5166_;
  assign new_D5144_ = ~new_D5112_ & new_D5113_;
  assign new_D5145_ = new_D5112_ & ~new_D5113_;
  assign new_D5146_ = ~new_D5128_ | new_D5138_;
  assign new_D5147_ = new_D5128_ & new_D5138_;
  assign new_D5148_ = ~new_D5128_ & ~new_D5138_;
  assign new_D5149_ = new_D5170_ | new_D5169_;
  assign new_D5150_ = new_D5116_ | new_D5149_;
  assign new_D5151_ = new_D5174_ | new_D5173_;
  assign new_D5152_ = ~new_D5116_ & new_D5151_;
  assign new_D5153_ = new_D5172_ | new_D5171_;
  assign new_D5154_ = new_D5116_ & new_D5153_;
  assign new_D5155_ = new_D5114_ & ~new_D5124_;
  assign new_D5156_ = ~new_D5114_ & new_D5124_;
  assign new_D5157_ = ~new_D5113_ | ~new_D5138_;
  assign new_D5158_ = new_D5124_ & new_D5157_;
  assign new_D5159_ = ~new_D5124_ & ~new_D5158_;
  assign new_D5160_ = new_D5124_ | new_D5157_;
  assign new_D5161_ = ~new_D5114_ & new_D5115_;
  assign new_D5162_ = new_D5114_ & ~new_D5115_;
  assign new_D5163_ = new_D5131_ | new_D5168_;
  assign new_D5164_ = ~new_D5131_ & ~new_D5167_;
  assign new_D5165_ = new_D5114_ | new_D5131_;
  assign new_D5166_ = new_D5114_ | new_D5115_;
  assign new_D5167_ = new_D5131_ & new_D5168_;
  assign new_D5168_ = ~new_D5113_ | ~new_D5138_;
  assign new_D5169_ = new_D5146_ & new_D5166_;
  assign new_D5170_ = ~new_D5146_ & ~new_D5166_;
  assign new_D5171_ = new_D5175_ | new_D5176_;
  assign new_D5172_ = ~new_D5117_ & new_D5131_;
  assign new_D5173_ = new_D5177_ | new_D5178_;
  assign new_D5174_ = new_D5117_ & new_D5131_;
  assign new_D5175_ = ~new_D5117_ & ~new_D5131_;
  assign new_D5176_ = new_D5117_ & ~new_D5131_;
  assign new_D5177_ = new_D5117_ & ~new_D5131_;
  assign new_D5178_ = ~new_D5117_ & new_D5131_;
  assign new_D5179_ = new_E618_;
  assign new_D5180_ = new_E685_;
  assign new_D5181_ = new_E752_;
  assign new_D5182_ = new_E819_;
  assign new_D5183_ = new_E886_;
  assign new_D5184_ = new_E953_;
  assign new_D5185_ = new_D5192_ & new_D5191_;
  assign new_D5186_ = new_D5194_ | new_D5193_;
  assign new_D5187_ = new_D5196_ | new_D5195_;
  assign new_D5188_ = new_D5198_ & new_D5197_;
  assign new_D5189_ = new_D5198_ & new_D5199_;
  assign new_D5190_ = new_D5191_ | new_D5200_;
  assign new_D5191_ = new_D5180_ | new_D5203_;
  assign new_D5192_ = new_D5202_ | new_D5201_;
  assign new_D5193_ = new_D5207_ & new_D5206_;
  assign new_D5194_ = new_D5205_ & new_D5204_;
  assign new_D5195_ = new_D5210_ | new_D5209_;
  assign new_D5196_ = new_D5205_ & new_D5208_;
  assign new_D5197_ = new_D5180_ | new_D5213_;
  assign new_D5198_ = new_D5212_ | new_D5211_;
  assign new_D5199_ = new_D5215_ | new_D5214_;
  assign new_D5200_ = ~new_D5191_ & new_D5217_;
  assign new_D5201_ = ~new_D5193_ & new_D5205_;
  assign new_D5202_ = new_D5193_ & ~new_D5205_;
  assign new_D5203_ = new_D5179_ & ~new_D5180_;
  assign new_D5204_ = ~new_D5226_ | ~new_D5227_;
  assign new_D5205_ = new_D5219_ | new_D5221_;
  assign new_D5206_ = new_D5229_ | new_D5228_;
  assign new_D5207_ = new_D5223_ | new_D5222_;
  assign new_D5208_ = ~new_D5231_ | ~new_D5230_;
  assign new_D5209_ = ~new_D5232_ & new_D5233_;
  assign new_D5210_ = new_D5232_ & ~new_D5233_;
  assign new_D5211_ = ~new_D5179_ & new_D5180_;
  assign new_D5212_ = new_D5179_ & ~new_D5180_;
  assign new_D5213_ = ~new_D5195_ | new_D5205_;
  assign new_D5214_ = new_D5195_ & new_D5205_;
  assign new_D5215_ = ~new_D5195_ & ~new_D5205_;
  assign new_D5216_ = new_D5237_ | new_D5236_;
  assign new_D5217_ = new_D5183_ | new_D5216_;
  assign new_D5218_ = new_D5241_ | new_D5240_;
  assign new_D5219_ = ~new_D5183_ & new_D5218_;
  assign new_D5220_ = new_D5239_ | new_D5238_;
  assign new_D5221_ = new_D5183_ & new_D5220_;
  assign new_D5222_ = new_D5181_ & ~new_D5191_;
  assign new_D5223_ = ~new_D5181_ & new_D5191_;
  assign new_D5224_ = ~new_D5180_ | ~new_D5205_;
  assign new_D5225_ = new_D5191_ & new_D5224_;
  assign new_D5226_ = ~new_D5191_ & ~new_D5225_;
  assign new_D5227_ = new_D5191_ | new_D5224_;
  assign new_D5228_ = ~new_D5181_ & new_D5182_;
  assign new_D5229_ = new_D5181_ & ~new_D5182_;
  assign new_D5230_ = new_D5198_ | new_D5235_;
  assign new_D5231_ = ~new_D5198_ & ~new_D5234_;
  assign new_D5232_ = new_D5181_ | new_D5198_;
  assign new_D5233_ = new_D5181_ | new_D5182_;
  assign new_D5234_ = new_D5198_ & new_D5235_;
  assign new_D5235_ = ~new_D5180_ | ~new_D5205_;
  assign new_D5236_ = new_D5213_ & new_D5233_;
  assign new_D5237_ = ~new_D5213_ & ~new_D5233_;
  assign new_D5238_ = new_D5242_ | new_D5243_;
  assign new_D5239_ = ~new_D5184_ & new_D5198_;
  assign new_D5240_ = new_D5244_ | new_D5245_;
  assign new_D5241_ = new_D5184_ & new_D5198_;
  assign new_D5242_ = ~new_D5184_ & ~new_D5198_;
  assign new_D5243_ = new_D5184_ & ~new_D5198_;
  assign new_D5244_ = new_D5184_ & ~new_D5198_;
  assign new_D5245_ = ~new_D5184_ & new_D5198_;
  assign new_D5246_ = new_E1020_;
  assign new_D5247_ = new_E1087_;
  assign new_D5248_ = new_E1154_;
  assign new_D5249_ = new_E1221_;
  assign new_D5250_ = new_E1288_;
  assign new_D5251_ = new_E1355_;
  assign new_D5252_ = new_D5259_ & new_D5258_;
  assign new_D5253_ = new_D5261_ | new_D5260_;
  assign new_D5254_ = new_D5263_ | new_D5262_;
  assign new_D5255_ = new_D5265_ & new_D5264_;
  assign new_D5256_ = new_D5265_ & new_D5266_;
  assign new_D5257_ = new_D5258_ | new_D5267_;
  assign new_D5258_ = new_D5247_ | new_D5270_;
  assign new_D5259_ = new_D5269_ | new_D5268_;
  assign new_D5260_ = new_D5274_ & new_D5273_;
  assign new_D5261_ = new_D5272_ & new_D5271_;
  assign new_D5262_ = new_D5277_ | new_D5276_;
  assign new_D5263_ = new_D5272_ & new_D5275_;
  assign new_D5264_ = new_D5247_ | new_D5280_;
  assign new_D5265_ = new_D5279_ | new_D5278_;
  assign new_D5266_ = new_D5282_ | new_D5281_;
  assign new_D5267_ = ~new_D5258_ & new_D5284_;
  assign new_D5268_ = ~new_D5260_ & new_D5272_;
  assign new_D5269_ = new_D5260_ & ~new_D5272_;
  assign new_D5270_ = new_D5246_ & ~new_D5247_;
  assign new_D5271_ = ~new_D5293_ | ~new_D5294_;
  assign new_D5272_ = new_D5286_ | new_D5288_;
  assign new_D5273_ = new_D5296_ | new_D5295_;
  assign new_D5274_ = new_D5290_ | new_D5289_;
  assign new_D5275_ = ~new_D5298_ | ~new_D5297_;
  assign new_D5276_ = ~new_D5299_ & new_D5300_;
  assign new_D5277_ = new_D5299_ & ~new_D5300_;
  assign new_D5278_ = ~new_D5246_ & new_D5247_;
  assign new_D5279_ = new_D5246_ & ~new_D5247_;
  assign new_D5280_ = ~new_D5262_ | new_D5272_;
  assign new_D5281_ = new_D5262_ & new_D5272_;
  assign new_D5282_ = ~new_D5262_ & ~new_D5272_;
  assign new_D5283_ = new_D5304_ | new_D5303_;
  assign new_D5284_ = new_D5250_ | new_D5283_;
  assign new_D5285_ = new_D5308_ | new_D5307_;
  assign new_D5286_ = ~new_D5250_ & new_D5285_;
  assign new_D5287_ = new_D5306_ | new_D5305_;
  assign new_D5288_ = new_D5250_ & new_D5287_;
  assign new_D5289_ = new_D5248_ & ~new_D5258_;
  assign new_D5290_ = ~new_D5248_ & new_D5258_;
  assign new_D5291_ = ~new_D5247_ | ~new_D5272_;
  assign new_D5292_ = new_D5258_ & new_D5291_;
  assign new_D5293_ = ~new_D5258_ & ~new_D5292_;
  assign new_D5294_ = new_D5258_ | new_D5291_;
  assign new_D5295_ = ~new_D5248_ & new_D5249_;
  assign new_D5296_ = new_D5248_ & ~new_D5249_;
  assign new_D5297_ = new_D5265_ | new_D5302_;
  assign new_D5298_ = ~new_D5265_ & ~new_D5301_;
  assign new_D5299_ = new_D5248_ | new_D5265_;
  assign new_D5300_ = new_D5248_ | new_D5249_;
  assign new_D5301_ = new_D5265_ & new_D5302_;
  assign new_D5302_ = ~new_D5247_ | ~new_D5272_;
  assign new_D5303_ = new_D5280_ & new_D5300_;
  assign new_D5304_ = ~new_D5280_ & ~new_D5300_;
  assign new_D5305_ = new_D5309_ | new_D5310_;
  assign new_D5306_ = ~new_D5251_ & new_D5265_;
  assign new_D5307_ = new_D5311_ | new_D5312_;
  assign new_D5308_ = new_D5251_ & new_D5265_;
  assign new_D5309_ = ~new_D5251_ & ~new_D5265_;
  assign new_D5310_ = new_D5251_ & ~new_D5265_;
  assign new_D5311_ = new_D5251_ & ~new_D5265_;
  assign new_D5312_ = ~new_D5251_ & new_D5265_;
  assign new_D5313_ = new_E1422_;
  assign new_D5314_ = new_E1489_;
  assign new_D5315_ = new_E1556_;
  assign new_D5316_ = new_E1623_;
  assign new_D5317_ = new_E1690_;
  assign new_D5318_ = new_E1757_;
  assign new_D5319_ = new_D5326_ & new_D5325_;
  assign new_D5320_ = new_D5328_ | new_D5327_;
  assign new_D5321_ = new_D5330_ | new_D5329_;
  assign new_D5322_ = new_D5332_ & new_D5331_;
  assign new_D5323_ = new_D5332_ & new_D5333_;
  assign new_D5324_ = new_D5325_ | new_D5334_;
  assign new_D5325_ = new_D5314_ | new_D5337_;
  assign new_D5326_ = new_D5336_ | new_D5335_;
  assign new_D5327_ = new_D5341_ & new_D5340_;
  assign new_D5328_ = new_D5339_ & new_D5338_;
  assign new_D5329_ = new_D5344_ | new_D5343_;
  assign new_D5330_ = new_D5339_ & new_D5342_;
  assign new_D5331_ = new_D5314_ | new_D5347_;
  assign new_D5332_ = new_D5346_ | new_D5345_;
  assign new_D5333_ = new_D5349_ | new_D5348_;
  assign new_D5334_ = ~new_D5325_ & new_D5351_;
  assign new_D5335_ = ~new_D5327_ & new_D5339_;
  assign new_D5336_ = new_D5327_ & ~new_D5339_;
  assign new_D5337_ = new_D5313_ & ~new_D5314_;
  assign new_D5338_ = ~new_D5360_ | ~new_D5361_;
  assign new_D5339_ = new_D5353_ | new_D5355_;
  assign new_D5340_ = new_D5363_ | new_D5362_;
  assign new_D5341_ = new_D5357_ | new_D5356_;
  assign new_D5342_ = ~new_D5365_ | ~new_D5364_;
  assign new_D5343_ = ~new_D5366_ & new_D5367_;
  assign new_D5344_ = new_D5366_ & ~new_D5367_;
  assign new_D5345_ = ~new_D5313_ & new_D5314_;
  assign new_D5346_ = new_D5313_ & ~new_D5314_;
  assign new_D5347_ = ~new_D5329_ | new_D5339_;
  assign new_D5348_ = new_D5329_ & new_D5339_;
  assign new_D5349_ = ~new_D5329_ & ~new_D5339_;
  assign new_D5350_ = new_D5371_ | new_D5370_;
  assign new_D5351_ = new_D5317_ | new_D5350_;
  assign new_D5352_ = new_D5375_ | new_D5374_;
  assign new_D5353_ = ~new_D5317_ & new_D5352_;
  assign new_D5354_ = new_D5373_ | new_D5372_;
  assign new_D5355_ = new_D5317_ & new_D5354_;
  assign new_D5356_ = new_D5315_ & ~new_D5325_;
  assign new_D5357_ = ~new_D5315_ & new_D5325_;
  assign new_D5358_ = ~new_D5314_ | ~new_D5339_;
  assign new_D5359_ = new_D5325_ & new_D5358_;
  assign new_D5360_ = ~new_D5325_ & ~new_D5359_;
  assign new_D5361_ = new_D5325_ | new_D5358_;
  assign new_D5362_ = ~new_D5315_ & new_D5316_;
  assign new_D5363_ = new_D5315_ & ~new_D5316_;
  assign new_D5364_ = new_D5332_ | new_D5369_;
  assign new_D5365_ = ~new_D5332_ & ~new_D5368_;
  assign new_D5366_ = new_D5315_ | new_D5332_;
  assign new_D5367_ = new_D5315_ | new_D5316_;
  assign new_D5368_ = new_D5332_ & new_D5369_;
  assign new_D5369_ = ~new_D5314_ | ~new_D5339_;
  assign new_D5370_ = new_D5347_ & new_D5367_;
  assign new_D5371_ = ~new_D5347_ & ~new_D5367_;
  assign new_D5372_ = new_D5376_ | new_D5377_;
  assign new_D5373_ = ~new_D5318_ & new_D5332_;
  assign new_D5374_ = new_D5378_ | new_D5379_;
  assign new_D5375_ = new_D5318_ & new_D5332_;
  assign new_D5376_ = ~new_D5318_ & ~new_D5332_;
  assign new_D5377_ = new_D5318_ & ~new_D5332_;
  assign new_D5378_ = new_D5318_ & ~new_D5332_;
  assign new_D5379_ = ~new_D5318_ & new_D5332_;
  assign new_D5380_ = new_E1824_;
  assign new_D5381_ = new_E1891_;
  assign new_D5382_ = new_E1958_;
  assign new_D5383_ = new_E2025_;
  assign new_D5384_ = new_E2092_;
  assign new_D5385_ = new_E2159_;
  assign new_D5386_ = new_D5393_ & new_D5392_;
  assign new_D5387_ = new_D5395_ | new_D5394_;
  assign new_D5388_ = new_D5397_ | new_D5396_;
  assign new_D5389_ = new_D5399_ & new_D5398_;
  assign new_D5390_ = new_D5399_ & new_D5400_;
  assign new_D5391_ = new_D5392_ | new_D5401_;
  assign new_D5392_ = new_D5381_ | new_D5404_;
  assign new_D5393_ = new_D5403_ | new_D5402_;
  assign new_D5394_ = new_D5408_ & new_D5407_;
  assign new_D5395_ = new_D5406_ & new_D5405_;
  assign new_D5396_ = new_D5411_ | new_D5410_;
  assign new_D5397_ = new_D5406_ & new_D5409_;
  assign new_D5398_ = new_D5381_ | new_D5414_;
  assign new_D5399_ = new_D5413_ | new_D5412_;
  assign new_D5400_ = new_D5416_ | new_D5415_;
  assign new_D5401_ = ~new_D5392_ & new_D5418_;
  assign new_D5402_ = ~new_D5394_ & new_D5406_;
  assign new_D5403_ = new_D5394_ & ~new_D5406_;
  assign new_D5404_ = new_D5380_ & ~new_D5381_;
  assign new_D5405_ = ~new_D5427_ | ~new_D5428_;
  assign new_D5406_ = new_D5420_ | new_D5422_;
  assign new_D5407_ = new_D5430_ | new_D5429_;
  assign new_D5408_ = new_D5424_ | new_D5423_;
  assign new_D5409_ = ~new_D5432_ | ~new_D5431_;
  assign new_D5410_ = ~new_D5433_ & new_D5434_;
  assign new_D5411_ = new_D5433_ & ~new_D5434_;
  assign new_D5412_ = ~new_D5380_ & new_D5381_;
  assign new_D5413_ = new_D5380_ & ~new_D5381_;
  assign new_D5414_ = ~new_D5396_ | new_D5406_;
  assign new_D5415_ = new_D5396_ & new_D5406_;
  assign new_D5416_ = ~new_D5396_ & ~new_D5406_;
  assign new_D5417_ = new_D5438_ | new_D5437_;
  assign new_D5418_ = new_D5384_ | new_D5417_;
  assign new_D5419_ = new_D5442_ | new_D5441_;
  assign new_D5420_ = ~new_D5384_ & new_D5419_;
  assign new_D5421_ = new_D5440_ | new_D5439_;
  assign new_D5422_ = new_D5384_ & new_D5421_;
  assign new_D5423_ = new_D5382_ & ~new_D5392_;
  assign new_D5424_ = ~new_D5382_ & new_D5392_;
  assign new_D5425_ = ~new_D5381_ | ~new_D5406_;
  assign new_D5426_ = new_D5392_ & new_D5425_;
  assign new_D5427_ = ~new_D5392_ & ~new_D5426_;
  assign new_D5428_ = new_D5392_ | new_D5425_;
  assign new_D5429_ = ~new_D5382_ & new_D5383_;
  assign new_D5430_ = new_D5382_ & ~new_D5383_;
  assign new_D5431_ = new_D5399_ | new_D5436_;
  assign new_D5432_ = ~new_D5399_ & ~new_D5435_;
  assign new_D5433_ = new_D5382_ | new_D5399_;
  assign new_D5434_ = new_D5382_ | new_D5383_;
  assign new_D5435_ = new_D5399_ & new_D5436_;
  assign new_D5436_ = ~new_D5381_ | ~new_D5406_;
  assign new_D5437_ = new_D5414_ & new_D5434_;
  assign new_D5438_ = ~new_D5414_ & ~new_D5434_;
  assign new_D5439_ = new_D5443_ | new_D5444_;
  assign new_D5440_ = ~new_D5385_ & new_D5399_;
  assign new_D5441_ = new_D5445_ | new_D5446_;
  assign new_D5442_ = new_D5385_ & new_D5399_;
  assign new_D5443_ = ~new_D5385_ & ~new_D5399_;
  assign new_D5444_ = new_D5385_ & ~new_D5399_;
  assign new_D5445_ = new_D5385_ & ~new_D5399_;
  assign new_D5446_ = ~new_D5385_ & new_D5399_;
  assign new_D5447_ = new_E2226_;
  assign new_D5448_ = new_E2293_;
  assign new_D5449_ = new_E2360_;
  assign new_D5450_ = new_E2427_;
  assign new_D5451_ = new_E2494_;
  assign new_D5452_ = new_E2561_;
  assign new_D5453_ = new_D5460_ & new_D5459_;
  assign new_D5454_ = new_D5462_ | new_D5461_;
  assign new_D5455_ = new_D5464_ | new_D5463_;
  assign new_D5456_ = new_D5466_ & new_D5465_;
  assign new_D5457_ = new_D5466_ & new_D5467_;
  assign new_D5458_ = new_D5459_ | new_D5468_;
  assign new_D5459_ = new_D5448_ | new_D5471_;
  assign new_D5460_ = new_D5470_ | new_D5469_;
  assign new_D5461_ = new_D5475_ & new_D5474_;
  assign new_D5462_ = new_D5473_ & new_D5472_;
  assign new_D5463_ = new_D5478_ | new_D5477_;
  assign new_D5464_ = new_D5473_ & new_D5476_;
  assign new_D5465_ = new_D5448_ | new_D5481_;
  assign new_D5466_ = new_D5480_ | new_D5479_;
  assign new_D5467_ = new_D5483_ | new_D5482_;
  assign new_D5468_ = ~new_D5459_ & new_D5485_;
  assign new_D5469_ = ~new_D5461_ & new_D5473_;
  assign new_D5470_ = new_D5461_ & ~new_D5473_;
  assign new_D5471_ = new_D5447_ & ~new_D5448_;
  assign new_D5472_ = ~new_D5494_ | ~new_D5495_;
  assign new_D5473_ = new_D5487_ | new_D5489_;
  assign new_D5474_ = new_D5497_ | new_D5496_;
  assign new_D5475_ = new_D5491_ | new_D5490_;
  assign new_D5476_ = ~new_D5499_ | ~new_D5498_;
  assign new_D5477_ = ~new_D5500_ & new_D5501_;
  assign new_D5478_ = new_D5500_ & ~new_D5501_;
  assign new_D5479_ = ~new_D5447_ & new_D5448_;
  assign new_D5480_ = new_D5447_ & ~new_D5448_;
  assign new_D5481_ = ~new_D5463_ | new_D5473_;
  assign new_D5482_ = new_D5463_ & new_D5473_;
  assign new_D5483_ = ~new_D5463_ & ~new_D5473_;
  assign new_D5484_ = new_D5505_ | new_D5504_;
  assign new_D5485_ = new_D5451_ | new_D5484_;
  assign new_D5486_ = new_D5509_ | new_D5508_;
  assign new_D5487_ = ~new_D5451_ & new_D5486_;
  assign new_D5488_ = new_D5507_ | new_D5506_;
  assign new_D5489_ = new_D5451_ & new_D5488_;
  assign new_D5490_ = new_D5449_ & ~new_D5459_;
  assign new_D5491_ = ~new_D5449_ & new_D5459_;
  assign new_D5492_ = ~new_D5448_ | ~new_D5473_;
  assign new_D5493_ = new_D5459_ & new_D5492_;
  assign new_D5494_ = ~new_D5459_ & ~new_D5493_;
  assign new_D5495_ = new_D5459_ | new_D5492_;
  assign new_D5496_ = ~new_D5449_ & new_D5450_;
  assign new_D5497_ = new_D5449_ & ~new_D5450_;
  assign new_D5498_ = new_D5466_ | new_D5503_;
  assign new_D5499_ = ~new_D5466_ & ~new_D5502_;
  assign new_D5500_ = new_D5449_ | new_D5466_;
  assign new_D5501_ = new_D5449_ | new_D5450_;
  assign new_D5502_ = new_D5466_ & new_D5503_;
  assign new_D5503_ = ~new_D5448_ | ~new_D5473_;
  assign new_D5504_ = new_D5481_ & new_D5501_;
  assign new_D5505_ = ~new_D5481_ & ~new_D5501_;
  assign new_D5506_ = new_D5510_ | new_D5511_;
  assign new_D5507_ = ~new_D5452_ & new_D5466_;
  assign new_D5508_ = new_D5512_ | new_D5513_;
  assign new_D5509_ = new_D5452_ & new_D5466_;
  assign new_D5510_ = ~new_D5452_ & ~new_D5466_;
  assign new_D5511_ = new_D5452_ & ~new_D5466_;
  assign new_D5512_ = new_D5452_ & ~new_D5466_;
  assign new_D5513_ = ~new_D5452_ & new_D5466_;
  assign new_D5514_ = new_E2628_;
  assign new_D5515_ = new_E2695_;
  assign new_D5516_ = new_E2762_;
  assign new_D5517_ = new_E2829_;
  assign new_D5518_ = new_E2896_;
  assign new_D5519_ = new_E2963_;
  assign new_D5520_ = new_D5527_ & new_D5526_;
  assign new_D5521_ = new_D5529_ | new_D5528_;
  assign new_D5522_ = new_D5531_ | new_D5530_;
  assign new_D5523_ = new_D5533_ & new_D5532_;
  assign new_D5524_ = new_D5533_ & new_D5534_;
  assign new_D5525_ = new_D5526_ | new_D5535_;
  assign new_D5526_ = new_D5515_ | new_D5538_;
  assign new_D5527_ = new_D5537_ | new_D5536_;
  assign new_D5528_ = new_D5542_ & new_D5541_;
  assign new_D5529_ = new_D5540_ & new_D5539_;
  assign new_D5530_ = new_D5545_ | new_D5544_;
  assign new_D5531_ = new_D5540_ & new_D5543_;
  assign new_D5532_ = new_D5515_ | new_D5548_;
  assign new_D5533_ = new_D5547_ | new_D5546_;
  assign new_D5534_ = new_D5550_ | new_D5549_;
  assign new_D5535_ = ~new_D5526_ & new_D5552_;
  assign new_D5536_ = ~new_D5528_ & new_D5540_;
  assign new_D5537_ = new_D5528_ & ~new_D5540_;
  assign new_D5538_ = new_D5514_ & ~new_D5515_;
  assign new_D5539_ = ~new_D5561_ | ~new_D5562_;
  assign new_D5540_ = new_D5554_ | new_D5556_;
  assign new_D5541_ = new_D5564_ | new_D5563_;
  assign new_D5542_ = new_D5558_ | new_D5557_;
  assign new_D5543_ = ~new_D5566_ | ~new_D5565_;
  assign new_D5544_ = ~new_D5567_ & new_D5568_;
  assign new_D5545_ = new_D5567_ & ~new_D5568_;
  assign new_D5546_ = ~new_D5514_ & new_D5515_;
  assign new_D5547_ = new_D5514_ & ~new_D5515_;
  assign new_D5548_ = ~new_D5530_ | new_D5540_;
  assign new_D5549_ = new_D5530_ & new_D5540_;
  assign new_D5550_ = ~new_D5530_ & ~new_D5540_;
  assign new_D5551_ = new_D5572_ | new_D5571_;
  assign new_D5552_ = new_D5518_ | new_D5551_;
  assign new_D5553_ = new_D5576_ | new_D5575_;
  assign new_D5554_ = ~new_D5518_ & new_D5553_;
  assign new_D5555_ = new_D5574_ | new_D5573_;
  assign new_D5556_ = new_D5518_ & new_D5555_;
  assign new_D5557_ = new_D5516_ & ~new_D5526_;
  assign new_D5558_ = ~new_D5516_ & new_D5526_;
  assign new_D5559_ = ~new_D5515_ | ~new_D5540_;
  assign new_D5560_ = new_D5526_ & new_D5559_;
  assign new_D5561_ = ~new_D5526_ & ~new_D5560_;
  assign new_D5562_ = new_D5526_ | new_D5559_;
  assign new_D5563_ = ~new_D5516_ & new_D5517_;
  assign new_D5564_ = new_D5516_ & ~new_D5517_;
  assign new_D5565_ = new_D5533_ | new_D5570_;
  assign new_D5566_ = ~new_D5533_ & ~new_D5569_;
  assign new_D5567_ = new_D5516_ | new_D5533_;
  assign new_D5568_ = new_D5516_ | new_D5517_;
  assign new_D5569_ = new_D5533_ & new_D5570_;
  assign new_D5570_ = ~new_D5515_ | ~new_D5540_;
  assign new_D5571_ = new_D5548_ & new_D5568_;
  assign new_D5572_ = ~new_D5548_ & ~new_D5568_;
  assign new_D5573_ = new_D5577_ | new_D5578_;
  assign new_D5574_ = ~new_D5519_ & new_D5533_;
  assign new_D5575_ = new_D5579_ | new_D5580_;
  assign new_D5576_ = new_D5519_ & new_D5533_;
  assign new_D5577_ = ~new_D5519_ & ~new_D5533_;
  assign new_D5578_ = new_D5519_ & ~new_D5533_;
  assign new_D5579_ = new_D5519_ & ~new_D5533_;
  assign new_D5580_ = ~new_D5519_ & new_D5533_;
  assign new_D5581_ = new_E3030_;
  assign new_D5582_ = new_E3097_;
  assign new_D5583_ = new_E3164_;
  assign new_D5584_ = new_E3231_;
  assign new_D5585_ = new_E3298_;
  assign new_D5586_ = new_E3365_;
  assign new_D5587_ = new_D5594_ & new_D5593_;
  assign new_D5588_ = new_D5596_ | new_D5595_;
  assign new_D5589_ = new_D5598_ | new_D5597_;
  assign new_D5590_ = new_D5600_ & new_D5599_;
  assign new_D5591_ = new_D5600_ & new_D5601_;
  assign new_D5592_ = new_D5593_ | new_D5602_;
  assign new_D5593_ = new_D5582_ | new_D5605_;
  assign new_D5594_ = new_D5604_ | new_D5603_;
  assign new_D5595_ = new_D5609_ & new_D5608_;
  assign new_D5596_ = new_D5607_ & new_D5606_;
  assign new_D5597_ = new_D5612_ | new_D5611_;
  assign new_D5598_ = new_D5607_ & new_D5610_;
  assign new_D5599_ = new_D5582_ | new_D5615_;
  assign new_D5600_ = new_D5614_ | new_D5613_;
  assign new_D5601_ = new_D5617_ | new_D5616_;
  assign new_D5602_ = ~new_D5593_ & new_D5619_;
  assign new_D5603_ = ~new_D5595_ & new_D5607_;
  assign new_D5604_ = new_D5595_ & ~new_D5607_;
  assign new_D5605_ = new_D5581_ & ~new_D5582_;
  assign new_D5606_ = ~new_D5628_ | ~new_D5629_;
  assign new_D5607_ = new_D5621_ | new_D5623_;
  assign new_D5608_ = new_D5631_ | new_D5630_;
  assign new_D5609_ = new_D5625_ | new_D5624_;
  assign new_D5610_ = ~new_D5633_ | ~new_D5632_;
  assign new_D5611_ = ~new_D5634_ & new_D5635_;
  assign new_D5612_ = new_D5634_ & ~new_D5635_;
  assign new_D5613_ = ~new_D5581_ & new_D5582_;
  assign new_D5614_ = new_D5581_ & ~new_D5582_;
  assign new_D5615_ = ~new_D5597_ | new_D5607_;
  assign new_D5616_ = new_D5597_ & new_D5607_;
  assign new_D5617_ = ~new_D5597_ & ~new_D5607_;
  assign new_D5618_ = new_D5639_ | new_D5638_;
  assign new_D5619_ = new_D5585_ | new_D5618_;
  assign new_D5620_ = new_D5643_ | new_D5642_;
  assign new_D5621_ = ~new_D5585_ & new_D5620_;
  assign new_D5622_ = new_D5641_ | new_D5640_;
  assign new_D5623_ = new_D5585_ & new_D5622_;
  assign new_D5624_ = new_D5583_ & ~new_D5593_;
  assign new_D5625_ = ~new_D5583_ & new_D5593_;
  assign new_D5626_ = ~new_D5582_ | ~new_D5607_;
  assign new_D5627_ = new_D5593_ & new_D5626_;
  assign new_D5628_ = ~new_D5593_ & ~new_D5627_;
  assign new_D5629_ = new_D5593_ | new_D5626_;
  assign new_D5630_ = ~new_D5583_ & new_D5584_;
  assign new_D5631_ = new_D5583_ & ~new_D5584_;
  assign new_D5632_ = new_D5600_ | new_D5637_;
  assign new_D5633_ = ~new_D5600_ & ~new_D5636_;
  assign new_D5634_ = new_D5583_ | new_D5600_;
  assign new_D5635_ = new_D5583_ | new_D5584_;
  assign new_D5636_ = new_D5600_ & new_D5637_;
  assign new_D5637_ = ~new_D5582_ | ~new_D5607_;
  assign new_D5638_ = new_D5615_ & new_D5635_;
  assign new_D5639_ = ~new_D5615_ & ~new_D5635_;
  assign new_D5640_ = new_D5644_ | new_D5645_;
  assign new_D5641_ = ~new_D5586_ & new_D5600_;
  assign new_D5642_ = new_D5646_ | new_D5647_;
  assign new_D5643_ = new_D5586_ & new_D5600_;
  assign new_D5644_ = ~new_D5586_ & ~new_D5600_;
  assign new_D5645_ = new_D5586_ & ~new_D5600_;
  assign new_D5646_ = new_D5586_ & ~new_D5600_;
  assign new_D5647_ = ~new_D5586_ & new_D5600_;
  assign new_D5648_ = new_E3432_;
  assign new_D5649_ = new_E3499_;
  assign new_D5650_ = new_E3566_;
  assign new_D5651_ = new_E3633_;
  assign new_D5652_ = new_E3700_;
  assign new_D5653_ = new_E3767_;
  assign new_D5654_ = new_D5661_ & new_D5660_;
  assign new_D5655_ = new_D5663_ | new_D5662_;
  assign new_D5656_ = new_D5665_ | new_D5664_;
  assign new_D5657_ = new_D5667_ & new_D5666_;
  assign new_D5658_ = new_D5667_ & new_D5668_;
  assign new_D5659_ = new_D5660_ | new_D5669_;
  assign new_D5660_ = new_D5649_ | new_D5672_;
  assign new_D5661_ = new_D5671_ | new_D5670_;
  assign new_D5662_ = new_D5676_ & new_D5675_;
  assign new_D5663_ = new_D5674_ & new_D5673_;
  assign new_D5664_ = new_D5679_ | new_D5678_;
  assign new_D5665_ = new_D5674_ & new_D5677_;
  assign new_D5666_ = new_D5649_ | new_D5682_;
  assign new_D5667_ = new_D5681_ | new_D5680_;
  assign new_D5668_ = new_D5684_ | new_D5683_;
  assign new_D5669_ = ~new_D5660_ & new_D5686_;
  assign new_D5670_ = ~new_D5662_ & new_D5674_;
  assign new_D5671_ = new_D5662_ & ~new_D5674_;
  assign new_D5672_ = new_D5648_ & ~new_D5649_;
  assign new_D5673_ = ~new_D5695_ | ~new_D5696_;
  assign new_D5674_ = new_D5688_ | new_D5690_;
  assign new_D5675_ = new_D5698_ | new_D5697_;
  assign new_D5676_ = new_D5692_ | new_D5691_;
  assign new_D5677_ = ~new_D5700_ | ~new_D5699_;
  assign new_D5678_ = ~new_D5701_ & new_D5702_;
  assign new_D5679_ = new_D5701_ & ~new_D5702_;
  assign new_D5680_ = ~new_D5648_ & new_D5649_;
  assign new_D5681_ = new_D5648_ & ~new_D5649_;
  assign new_D5682_ = ~new_D5664_ | new_D5674_;
  assign new_D5683_ = new_D5664_ & new_D5674_;
  assign new_D5684_ = ~new_D5664_ & ~new_D5674_;
  assign new_D5685_ = new_D5706_ | new_D5705_;
  assign new_D5686_ = new_D5652_ | new_D5685_;
  assign new_D5687_ = new_D5710_ | new_D5709_;
  assign new_D5688_ = ~new_D5652_ & new_D5687_;
  assign new_D5689_ = new_D5708_ | new_D5707_;
  assign new_D5690_ = new_D5652_ & new_D5689_;
  assign new_D5691_ = new_D5650_ & ~new_D5660_;
  assign new_D5692_ = ~new_D5650_ & new_D5660_;
  assign new_D5693_ = ~new_D5649_ | ~new_D5674_;
  assign new_D5694_ = new_D5660_ & new_D5693_;
  assign new_D5695_ = ~new_D5660_ & ~new_D5694_;
  assign new_D5696_ = new_D5660_ | new_D5693_;
  assign new_D5697_ = ~new_D5650_ & new_D5651_;
  assign new_D5698_ = new_D5650_ & ~new_D5651_;
  assign new_D5699_ = new_D5667_ | new_D5704_;
  assign new_D5700_ = ~new_D5667_ & ~new_D5703_;
  assign new_D5701_ = new_D5650_ | new_D5667_;
  assign new_D5702_ = new_D5650_ | new_D5651_;
  assign new_D5703_ = new_D5667_ & new_D5704_;
  assign new_D5704_ = ~new_D5649_ | ~new_D5674_;
  assign new_D5705_ = new_D5682_ & new_D5702_;
  assign new_D5706_ = ~new_D5682_ & ~new_D5702_;
  assign new_D5707_ = new_D5711_ | new_D5712_;
  assign new_D5708_ = ~new_D5653_ & new_D5667_;
  assign new_D5709_ = new_D5713_ | new_D5714_;
  assign new_D5710_ = new_D5653_ & new_D5667_;
  assign new_D5711_ = ~new_D5653_ & ~new_D5667_;
  assign new_D5712_ = new_D5653_ & ~new_D5667_;
  assign new_D5713_ = new_D5653_ & ~new_D5667_;
  assign new_D5714_ = ~new_D5653_ & new_D5667_;
  assign new_D5715_ = new_E3834_;
  assign new_D5716_ = new_E3901_;
  assign new_D5717_ = new_E3968_;
  assign new_D5718_ = new_E4035_;
  assign new_D5719_ = new_E4102_;
  assign new_D5720_ = new_E4169_;
  assign new_D5721_ = new_D5728_ & new_D5727_;
  assign new_D5722_ = new_D5730_ | new_D5729_;
  assign new_D5723_ = new_D5732_ | new_D5731_;
  assign new_D5724_ = new_D5734_ & new_D5733_;
  assign new_D5725_ = new_D5734_ & new_D5735_;
  assign new_D5726_ = new_D5727_ | new_D5736_;
  assign new_D5727_ = new_D5716_ | new_D5739_;
  assign new_D5728_ = new_D5738_ | new_D5737_;
  assign new_D5729_ = new_D5743_ & new_D5742_;
  assign new_D5730_ = new_D5741_ & new_D5740_;
  assign new_D5731_ = new_D5746_ | new_D5745_;
  assign new_D5732_ = new_D5741_ & new_D5744_;
  assign new_D5733_ = new_D5716_ | new_D5749_;
  assign new_D5734_ = new_D5748_ | new_D5747_;
  assign new_D5735_ = new_D5751_ | new_D5750_;
  assign new_D5736_ = ~new_D5727_ & new_D5753_;
  assign new_D5737_ = ~new_D5729_ & new_D5741_;
  assign new_D5738_ = new_D5729_ & ~new_D5741_;
  assign new_D5739_ = new_D5715_ & ~new_D5716_;
  assign new_D5740_ = ~new_D5762_ | ~new_D5763_;
  assign new_D5741_ = new_D5755_ | new_D5757_;
  assign new_D5742_ = new_D5765_ | new_D5764_;
  assign new_D5743_ = new_D5759_ | new_D5758_;
  assign new_D5744_ = ~new_D5767_ | ~new_D5766_;
  assign new_D5745_ = ~new_D5768_ & new_D5769_;
  assign new_D5746_ = new_D5768_ & ~new_D5769_;
  assign new_D5747_ = ~new_D5715_ & new_D5716_;
  assign new_D5748_ = new_D5715_ & ~new_D5716_;
  assign new_D5749_ = ~new_D5731_ | new_D5741_;
  assign new_D5750_ = new_D5731_ & new_D5741_;
  assign new_D5751_ = ~new_D5731_ & ~new_D5741_;
  assign new_D5752_ = new_D5773_ | new_D5772_;
  assign new_D5753_ = new_D5719_ | new_D5752_;
  assign new_D5754_ = new_D5777_ | new_D5776_;
  assign new_D5755_ = ~new_D5719_ & new_D5754_;
  assign new_D5756_ = new_D5775_ | new_D5774_;
  assign new_D5757_ = new_D5719_ & new_D5756_;
  assign new_D5758_ = new_D5717_ & ~new_D5727_;
  assign new_D5759_ = ~new_D5717_ & new_D5727_;
  assign new_D5760_ = ~new_D5716_ | ~new_D5741_;
  assign new_D5761_ = new_D5727_ & new_D5760_;
  assign new_D5762_ = ~new_D5727_ & ~new_D5761_;
  assign new_D5763_ = new_D5727_ | new_D5760_;
  assign new_D5764_ = ~new_D5717_ & new_D5718_;
  assign new_D5765_ = new_D5717_ & ~new_D5718_;
  assign new_D5766_ = new_D5734_ | new_D5771_;
  assign new_D5767_ = ~new_D5734_ & ~new_D5770_;
  assign new_D5768_ = new_D5717_ | new_D5734_;
  assign new_D5769_ = new_D5717_ | new_D5718_;
  assign new_D5770_ = new_D5734_ & new_D5771_;
  assign new_D5771_ = ~new_D5716_ | ~new_D5741_;
  assign new_D5772_ = new_D5749_ & new_D5769_;
  assign new_D5773_ = ~new_D5749_ & ~new_D5769_;
  assign new_D5774_ = new_D5778_ | new_D5779_;
  assign new_D5775_ = ~new_D5720_ & new_D5734_;
  assign new_D5776_ = new_D5780_ | new_D5781_;
  assign new_D5777_ = new_D5720_ & new_D5734_;
  assign new_D5778_ = ~new_D5720_ & ~new_D5734_;
  assign new_D5779_ = new_D5720_ & ~new_D5734_;
  assign new_D5780_ = new_D5720_ & ~new_D5734_;
  assign new_D5781_ = ~new_D5720_ & new_D5734_;
  assign new_D5782_ = new_E4236_;
  assign new_D5783_ = new_E4303_;
  assign new_D5784_ = new_E4370_;
  assign new_D5785_ = new_E4437_;
  assign new_D5786_ = new_E4504_;
  assign new_D5787_ = new_E4571_;
  assign new_D5788_ = new_D5795_ & new_D5794_;
  assign new_D5789_ = new_D5797_ | new_D5796_;
  assign new_D5790_ = new_D5799_ | new_D5798_;
  assign new_D5791_ = new_D5801_ & new_D5800_;
  assign new_D5792_ = new_D5801_ & new_D5802_;
  assign new_D5793_ = new_D5794_ | new_D5803_;
  assign new_D5794_ = new_D5783_ | new_D5806_;
  assign new_D5795_ = new_D5805_ | new_D5804_;
  assign new_D5796_ = new_D5810_ & new_D5809_;
  assign new_D5797_ = new_D5808_ & new_D5807_;
  assign new_D5798_ = new_D5813_ | new_D5812_;
  assign new_D5799_ = new_D5808_ & new_D5811_;
  assign new_D5800_ = new_D5783_ | new_D5816_;
  assign new_D5801_ = new_D5815_ | new_D5814_;
  assign new_D5802_ = new_D5818_ | new_D5817_;
  assign new_D5803_ = ~new_D5794_ & new_D5820_;
  assign new_D5804_ = ~new_D5796_ & new_D5808_;
  assign new_D5805_ = new_D5796_ & ~new_D5808_;
  assign new_D5806_ = new_D5782_ & ~new_D5783_;
  assign new_D5807_ = ~new_D5829_ | ~new_D5830_;
  assign new_D5808_ = new_D5822_ | new_D5824_;
  assign new_D5809_ = new_D5832_ | new_D5831_;
  assign new_D5810_ = new_D5826_ | new_D5825_;
  assign new_D5811_ = ~new_D5834_ | ~new_D5833_;
  assign new_D5812_ = ~new_D5835_ & new_D5836_;
  assign new_D5813_ = new_D5835_ & ~new_D5836_;
  assign new_D5814_ = ~new_D5782_ & new_D5783_;
  assign new_D5815_ = new_D5782_ & ~new_D5783_;
  assign new_D5816_ = ~new_D5798_ | new_D5808_;
  assign new_D5817_ = new_D5798_ & new_D5808_;
  assign new_D5818_ = ~new_D5798_ & ~new_D5808_;
  assign new_D5819_ = new_D5840_ | new_D5839_;
  assign new_D5820_ = new_D5786_ | new_D5819_;
  assign new_D5821_ = new_D5844_ | new_D5843_;
  assign new_D5822_ = ~new_D5786_ & new_D5821_;
  assign new_D5823_ = new_D5842_ | new_D5841_;
  assign new_D5824_ = new_D5786_ & new_D5823_;
  assign new_D5825_ = new_D5784_ & ~new_D5794_;
  assign new_D5826_ = ~new_D5784_ & new_D5794_;
  assign new_D5827_ = ~new_D5783_ | ~new_D5808_;
  assign new_D5828_ = new_D5794_ & new_D5827_;
  assign new_D5829_ = ~new_D5794_ & ~new_D5828_;
  assign new_D5830_ = new_D5794_ | new_D5827_;
  assign new_D5831_ = ~new_D5784_ & new_D5785_;
  assign new_D5832_ = new_D5784_ & ~new_D5785_;
  assign new_D5833_ = new_D5801_ | new_D5838_;
  assign new_D5834_ = ~new_D5801_ & ~new_D5837_;
  assign new_D5835_ = new_D5784_ | new_D5801_;
  assign new_D5836_ = new_D5784_ | new_D5785_;
  assign new_D5837_ = new_D5801_ & new_D5838_;
  assign new_D5838_ = ~new_D5783_ | ~new_D5808_;
  assign new_D5839_ = new_D5816_ & new_D5836_;
  assign new_D5840_ = ~new_D5816_ & ~new_D5836_;
  assign new_D5841_ = new_D5845_ | new_D5846_;
  assign new_D5842_ = ~new_D5787_ & new_D5801_;
  assign new_D5843_ = new_D5847_ | new_D5848_;
  assign new_D5844_ = new_D5787_ & new_D5801_;
  assign new_D5845_ = ~new_D5787_ & ~new_D5801_;
  assign new_D5846_ = new_D5787_ & ~new_D5801_;
  assign new_D5847_ = new_D5787_ & ~new_D5801_;
  assign new_D5848_ = ~new_D5787_ & new_D5801_;
  assign new_D5849_ = new_E4638_;
  assign new_D5850_ = new_E4705_;
  assign new_D5851_ = new_E4772_;
  assign new_D5852_ = new_E4839_;
  assign new_D5853_ = new_E4906_;
  assign new_D5854_ = new_E4973_;
  assign new_D5855_ = new_D5862_ & new_D5861_;
  assign new_D5856_ = new_D5864_ | new_D5863_;
  assign new_D5857_ = new_D5866_ | new_D5865_;
  assign new_D5858_ = new_D5868_ & new_D5867_;
  assign new_D5859_ = new_D5868_ & new_D5869_;
  assign new_D5860_ = new_D5861_ | new_D5870_;
  assign new_D5861_ = new_D5850_ | new_D5873_;
  assign new_D5862_ = new_D5872_ | new_D5871_;
  assign new_D5863_ = new_D5877_ & new_D5876_;
  assign new_D5864_ = new_D5875_ & new_D5874_;
  assign new_D5865_ = new_D5880_ | new_D5879_;
  assign new_D5866_ = new_D5875_ & new_D5878_;
  assign new_D5867_ = new_D5850_ | new_D5883_;
  assign new_D5868_ = new_D5882_ | new_D5881_;
  assign new_D5869_ = new_D5885_ | new_D5884_;
  assign new_D5870_ = ~new_D5861_ & new_D5887_;
  assign new_D5871_ = ~new_D5863_ & new_D5875_;
  assign new_D5872_ = new_D5863_ & ~new_D5875_;
  assign new_D5873_ = new_D5849_ & ~new_D5850_;
  assign new_D5874_ = ~new_D5896_ | ~new_D5897_;
  assign new_D5875_ = new_D5889_ | new_D5891_;
  assign new_D5876_ = new_D5899_ | new_D5898_;
  assign new_D5877_ = new_D5893_ | new_D5892_;
  assign new_D5878_ = ~new_D5901_ | ~new_D5900_;
  assign new_D5879_ = ~new_D5902_ & new_D5903_;
  assign new_D5880_ = new_D5902_ & ~new_D5903_;
  assign new_D5881_ = ~new_D5849_ & new_D5850_;
  assign new_D5882_ = new_D5849_ & ~new_D5850_;
  assign new_D5883_ = ~new_D5865_ | new_D5875_;
  assign new_D5884_ = new_D5865_ & new_D5875_;
  assign new_D5885_ = ~new_D5865_ & ~new_D5875_;
  assign new_D5886_ = new_D5907_ | new_D5906_;
  assign new_D5887_ = new_D5853_ | new_D5886_;
  assign new_D5888_ = new_D5911_ | new_D5910_;
  assign new_D5889_ = ~new_D5853_ & new_D5888_;
  assign new_D5890_ = new_D5909_ | new_D5908_;
  assign new_D5891_ = new_D5853_ & new_D5890_;
  assign new_D5892_ = new_D5851_ & ~new_D5861_;
  assign new_D5893_ = ~new_D5851_ & new_D5861_;
  assign new_D5894_ = ~new_D5850_ | ~new_D5875_;
  assign new_D5895_ = new_D5861_ & new_D5894_;
  assign new_D5896_ = ~new_D5861_ & ~new_D5895_;
  assign new_D5897_ = new_D5861_ | new_D5894_;
  assign new_D5898_ = ~new_D5851_ & new_D5852_;
  assign new_D5899_ = new_D5851_ & ~new_D5852_;
  assign new_D5900_ = new_D5868_ | new_D5905_;
  assign new_D5901_ = ~new_D5868_ & ~new_D5904_;
  assign new_D5902_ = new_D5851_ | new_D5868_;
  assign new_D5903_ = new_D5851_ | new_D5852_;
  assign new_D5904_ = new_D5868_ & new_D5905_;
  assign new_D5905_ = ~new_D5850_ | ~new_D5875_;
  assign new_D5906_ = new_D5883_ & new_D5903_;
  assign new_D5907_ = ~new_D5883_ & ~new_D5903_;
  assign new_D5908_ = new_D5912_ | new_D5913_;
  assign new_D5909_ = ~new_D5854_ & new_D5868_;
  assign new_D5910_ = new_D5914_ | new_D5915_;
  assign new_D5911_ = new_D5854_ & new_D5868_;
  assign new_D5912_ = ~new_D5854_ & ~new_D5868_;
  assign new_D5913_ = new_D5854_ & ~new_D5868_;
  assign new_D5914_ = new_D5854_ & ~new_D5868_;
  assign new_D5915_ = ~new_D5854_ & new_D5868_;
  assign new_D5916_ = new_E5040_;
  assign new_D5917_ = new_E5107_;
  assign new_D5918_ = new_E5174_;
  assign new_D5919_ = new_E5241_;
  assign new_D5920_ = new_E5308_;
  assign new_D5921_ = new_E5375_;
  assign new_D5922_ = new_D5929_ & new_D5928_;
  assign new_D5923_ = new_D5931_ | new_D5930_;
  assign new_D5924_ = new_D5933_ | new_D5932_;
  assign new_D5925_ = new_D5935_ & new_D5934_;
  assign new_D5926_ = new_D5935_ & new_D5936_;
  assign new_D5927_ = new_D5928_ | new_D5937_;
  assign new_D5928_ = new_D5917_ | new_D5940_;
  assign new_D5929_ = new_D5939_ | new_D5938_;
  assign new_D5930_ = new_D5944_ & new_D5943_;
  assign new_D5931_ = new_D5942_ & new_D5941_;
  assign new_D5932_ = new_D5947_ | new_D5946_;
  assign new_D5933_ = new_D5942_ & new_D5945_;
  assign new_D5934_ = new_D5917_ | new_D5950_;
  assign new_D5935_ = new_D5949_ | new_D5948_;
  assign new_D5936_ = new_D5952_ | new_D5951_;
  assign new_D5937_ = ~new_D5928_ & new_D5954_;
  assign new_D5938_ = ~new_D5930_ & new_D5942_;
  assign new_D5939_ = new_D5930_ & ~new_D5942_;
  assign new_D5940_ = new_D5916_ & ~new_D5917_;
  assign new_D5941_ = ~new_D5963_ | ~new_D5964_;
  assign new_D5942_ = new_D5956_ | new_D5958_;
  assign new_D5943_ = new_D5966_ | new_D5965_;
  assign new_D5944_ = new_D5960_ | new_D5959_;
  assign new_D5945_ = ~new_D5968_ | ~new_D5967_;
  assign new_D5946_ = ~new_D5969_ & new_D5970_;
  assign new_D5947_ = new_D5969_ & ~new_D5970_;
  assign new_D5948_ = ~new_D5916_ & new_D5917_;
  assign new_D5949_ = new_D5916_ & ~new_D5917_;
  assign new_D5950_ = ~new_D5932_ | new_D5942_;
  assign new_D5951_ = new_D5932_ & new_D5942_;
  assign new_D5952_ = ~new_D5932_ & ~new_D5942_;
  assign new_D5953_ = new_D5974_ | new_D5973_;
  assign new_D5954_ = new_D5920_ | new_D5953_;
  assign new_D5955_ = new_D5978_ | new_D5977_;
  assign new_D5956_ = ~new_D5920_ & new_D5955_;
  assign new_D5957_ = new_D5976_ | new_D5975_;
  assign new_D5958_ = new_D5920_ & new_D5957_;
  assign new_D5959_ = new_D5918_ & ~new_D5928_;
  assign new_D5960_ = ~new_D5918_ & new_D5928_;
  assign new_D5961_ = ~new_D5917_ | ~new_D5942_;
  assign new_D5962_ = new_D5928_ & new_D5961_;
  assign new_D5963_ = ~new_D5928_ & ~new_D5962_;
  assign new_D5964_ = new_D5928_ | new_D5961_;
  assign new_D5965_ = ~new_D5918_ & new_D5919_;
  assign new_D5966_ = new_D5918_ & ~new_D5919_;
  assign new_D5967_ = new_D5935_ | new_D5972_;
  assign new_D5968_ = ~new_D5935_ & ~new_D5971_;
  assign new_D5969_ = new_D5918_ | new_D5935_;
  assign new_D5970_ = new_D5918_ | new_D5919_;
  assign new_D5971_ = new_D5935_ & new_D5972_;
  assign new_D5972_ = ~new_D5917_ | ~new_D5942_;
  assign new_D5973_ = new_D5950_ & new_D5970_;
  assign new_D5974_ = ~new_D5950_ & ~new_D5970_;
  assign new_D5975_ = new_D5979_ | new_D5980_;
  assign new_D5976_ = ~new_D5921_ & new_D5935_;
  assign new_D5977_ = new_D5981_ | new_D5982_;
  assign new_D5978_ = new_D5921_ & new_D5935_;
  assign new_D5979_ = ~new_D5921_ & ~new_D5935_;
  assign new_D5980_ = new_D5921_ & ~new_D5935_;
  assign new_D5981_ = new_D5921_ & ~new_D5935_;
  assign new_D5982_ = ~new_D5921_ & new_D5935_;
  assign new_D5983_ = new_E5442_;
  assign new_D5984_ = new_E5509_;
  assign new_D5985_ = new_E5576_;
  assign new_D5986_ = new_E5643_;
  assign new_D5987_ = new_E5710_;
  assign new_D5988_ = new_E5777_;
  assign new_D5989_ = new_D5996_ & new_D5995_;
  assign new_D5990_ = new_D5998_ | new_D5997_;
  assign new_D5991_ = new_D6000_ | new_D5999_;
  assign new_D5992_ = new_D6002_ & new_D6001_;
  assign new_D5993_ = new_D6002_ & new_D6003_;
  assign new_D5994_ = new_D5995_ | new_D6004_;
  assign new_D5995_ = new_D5984_ | new_D6007_;
  assign new_D5996_ = new_D6006_ | new_D6005_;
  assign new_D5997_ = new_D6011_ & new_D6010_;
  assign new_D5998_ = new_D6009_ & new_D6008_;
  assign new_D5999_ = new_D6014_ | new_D6013_;
  assign new_D6000_ = new_D6009_ & new_D6012_;
  assign new_D6001_ = new_D5984_ | new_D6017_;
  assign new_D6002_ = new_D6016_ | new_D6015_;
  assign new_D6003_ = new_D6019_ | new_D6018_;
  assign new_D6004_ = ~new_D5995_ & new_D6021_;
  assign new_D6005_ = ~new_D5997_ & new_D6009_;
  assign new_D6006_ = new_D5997_ & ~new_D6009_;
  assign new_D6007_ = new_D5983_ & ~new_D5984_;
  assign new_D6008_ = ~new_D6030_ | ~new_D6031_;
  assign new_D6009_ = new_D6023_ | new_D6025_;
  assign new_D6010_ = new_D6033_ | new_D6032_;
  assign new_D6011_ = new_D6027_ | new_D6026_;
  assign new_D6012_ = ~new_D6035_ | ~new_D6034_;
  assign new_D6013_ = ~new_D6036_ & new_D6037_;
  assign new_D6014_ = new_D6036_ & ~new_D6037_;
  assign new_D6015_ = ~new_D5983_ & new_D5984_;
  assign new_D6016_ = new_D5983_ & ~new_D5984_;
  assign new_D6017_ = ~new_D5999_ | new_D6009_;
  assign new_D6018_ = new_D5999_ & new_D6009_;
  assign new_D6019_ = ~new_D5999_ & ~new_D6009_;
  assign new_D6020_ = new_D6041_ | new_D6040_;
  assign new_D6021_ = new_D5987_ | new_D6020_;
  assign new_D6022_ = new_D6045_ | new_D6044_;
  assign new_D6023_ = ~new_D5987_ & new_D6022_;
  assign new_D6024_ = new_D6043_ | new_D6042_;
  assign new_D6025_ = new_D5987_ & new_D6024_;
  assign new_D6026_ = new_D5985_ & ~new_D5995_;
  assign new_D6027_ = ~new_D5985_ & new_D5995_;
  assign new_D6028_ = ~new_D5984_ | ~new_D6009_;
  assign new_D6029_ = new_D5995_ & new_D6028_;
  assign new_D6030_ = ~new_D5995_ & ~new_D6029_;
  assign new_D6031_ = new_D5995_ | new_D6028_;
  assign new_D6032_ = ~new_D5985_ & new_D5986_;
  assign new_D6033_ = new_D5985_ & ~new_D5986_;
  assign new_D6034_ = new_D6002_ | new_D6039_;
  assign new_D6035_ = ~new_D6002_ & ~new_D6038_;
  assign new_D6036_ = new_D5985_ | new_D6002_;
  assign new_D6037_ = new_D5985_ | new_D5986_;
  assign new_D6038_ = new_D6002_ & new_D6039_;
  assign new_D6039_ = ~new_D5984_ | ~new_D6009_;
  assign new_D6040_ = new_D6017_ & new_D6037_;
  assign new_D6041_ = ~new_D6017_ & ~new_D6037_;
  assign new_D6042_ = new_D6046_ | new_D6047_;
  assign new_D6043_ = ~new_D5988_ & new_D6002_;
  assign new_D6044_ = new_D6048_ | new_D6049_;
  assign new_D6045_ = new_D5988_ & new_D6002_;
  assign new_D6046_ = ~new_D5988_ & ~new_D6002_;
  assign new_D6047_ = new_D5988_ & ~new_D6002_;
  assign new_D6048_ = new_D5988_ & ~new_D6002_;
  assign new_D6049_ = ~new_D5988_ & new_D6002_;
  assign new_D6050_ = new_E5844_;
  assign new_D6051_ = new_E5911_;
  assign new_D6052_ = new_E5978_;
  assign new_D6053_ = new_E6045_;
  assign new_D6054_ = new_E6112_;
  assign new_D6055_ = new_E6179_;
  assign new_D6056_ = new_D6063_ & new_D6062_;
  assign new_D6057_ = new_D6065_ | new_D6064_;
  assign new_D6058_ = new_D6067_ | new_D6066_;
  assign new_D6059_ = new_D6069_ & new_D6068_;
  assign new_D6060_ = new_D6069_ & new_D6070_;
  assign new_D6061_ = new_D6062_ | new_D6071_;
  assign new_D6062_ = new_D6051_ | new_D6074_;
  assign new_D6063_ = new_D6073_ | new_D6072_;
  assign new_D6064_ = new_D6078_ & new_D6077_;
  assign new_D6065_ = new_D6076_ & new_D6075_;
  assign new_D6066_ = new_D6081_ | new_D6080_;
  assign new_D6067_ = new_D6076_ & new_D6079_;
  assign new_D6068_ = new_D6051_ | new_D6084_;
  assign new_D6069_ = new_D6083_ | new_D6082_;
  assign new_D6070_ = new_D6086_ | new_D6085_;
  assign new_D6071_ = ~new_D6062_ & new_D6088_;
  assign new_D6072_ = ~new_D6064_ & new_D6076_;
  assign new_D6073_ = new_D6064_ & ~new_D6076_;
  assign new_D6074_ = new_D6050_ & ~new_D6051_;
  assign new_D6075_ = ~new_D6097_ | ~new_D6098_;
  assign new_D6076_ = new_D6090_ | new_D6092_;
  assign new_D6077_ = new_D6100_ | new_D6099_;
  assign new_D6078_ = new_D6094_ | new_D6093_;
  assign new_D6079_ = ~new_D6102_ | ~new_D6101_;
  assign new_D6080_ = ~new_D6103_ & new_D6104_;
  assign new_D6081_ = new_D6103_ & ~new_D6104_;
  assign new_D6082_ = ~new_D6050_ & new_D6051_;
  assign new_D6083_ = new_D6050_ & ~new_D6051_;
  assign new_D6084_ = ~new_D6066_ | new_D6076_;
  assign new_D6085_ = new_D6066_ & new_D6076_;
  assign new_D6086_ = ~new_D6066_ & ~new_D6076_;
  assign new_D6087_ = new_D6108_ | new_D6107_;
  assign new_D6088_ = new_D6054_ | new_D6087_;
  assign new_D6089_ = new_D6112_ | new_D6111_;
  assign new_D6090_ = ~new_D6054_ & new_D6089_;
  assign new_D6091_ = new_D6110_ | new_D6109_;
  assign new_D6092_ = new_D6054_ & new_D6091_;
  assign new_D6093_ = new_D6052_ & ~new_D6062_;
  assign new_D6094_ = ~new_D6052_ & new_D6062_;
  assign new_D6095_ = ~new_D6051_ | ~new_D6076_;
  assign new_D6096_ = new_D6062_ & new_D6095_;
  assign new_D6097_ = ~new_D6062_ & ~new_D6096_;
  assign new_D6098_ = new_D6062_ | new_D6095_;
  assign new_D6099_ = ~new_D6052_ & new_D6053_;
  assign new_D6100_ = new_D6052_ & ~new_D6053_;
  assign new_D6101_ = new_D6069_ | new_D6106_;
  assign new_D6102_ = ~new_D6069_ & ~new_D6105_;
  assign new_D6103_ = new_D6052_ | new_D6069_;
  assign new_D6104_ = new_D6052_ | new_D6053_;
  assign new_D6105_ = new_D6069_ & new_D6106_;
  assign new_D6106_ = ~new_D6051_ | ~new_D6076_;
  assign new_D6107_ = new_D6084_ & new_D6104_;
  assign new_D6108_ = ~new_D6084_ & ~new_D6104_;
  assign new_D6109_ = new_D6113_ | new_D6114_;
  assign new_D6110_ = ~new_D6055_ & new_D6069_;
  assign new_D6111_ = new_D6115_ | new_D6116_;
  assign new_D6112_ = new_D6055_ & new_D6069_;
  assign new_D6113_ = ~new_D6055_ & ~new_D6069_;
  assign new_D6114_ = new_D6055_ & ~new_D6069_;
  assign new_D6115_ = new_D6055_ & ~new_D6069_;
  assign new_D6116_ = ~new_D6055_ & new_D6069_;
  assign new_D6117_ = new_E6246_;
  assign new_D6118_ = new_E6313_;
  assign new_D6119_ = new_E6380_;
  assign new_D6120_ = new_E6447_;
  assign new_D6121_ = new_E6514_;
  assign new_D6122_ = new_E6581_;
  assign new_D6123_ = new_D6130_ & new_D6129_;
  assign new_D6124_ = new_D6132_ | new_D6131_;
  assign new_D6125_ = new_D6134_ | new_D6133_;
  assign new_D6126_ = new_D6136_ & new_D6135_;
  assign new_D6127_ = new_D6136_ & new_D6137_;
  assign new_D6128_ = new_D6129_ | new_D6138_;
  assign new_D6129_ = new_D6118_ | new_D6141_;
  assign new_D6130_ = new_D6140_ | new_D6139_;
  assign new_D6131_ = new_D6145_ & new_D6144_;
  assign new_D6132_ = new_D6143_ & new_D6142_;
  assign new_D6133_ = new_D6148_ | new_D6147_;
  assign new_D6134_ = new_D6143_ & new_D6146_;
  assign new_D6135_ = new_D6118_ | new_D6151_;
  assign new_D6136_ = new_D6150_ | new_D6149_;
  assign new_D6137_ = new_D6153_ | new_D6152_;
  assign new_D6138_ = ~new_D6129_ & new_D6155_;
  assign new_D6139_ = ~new_D6131_ & new_D6143_;
  assign new_D6140_ = new_D6131_ & ~new_D6143_;
  assign new_D6141_ = new_D6117_ & ~new_D6118_;
  assign new_D6142_ = ~new_D6164_ | ~new_D6165_;
  assign new_D6143_ = new_D6157_ | new_D6159_;
  assign new_D6144_ = new_D6167_ | new_D6166_;
  assign new_D6145_ = new_D6161_ | new_D6160_;
  assign new_D6146_ = ~new_D6169_ | ~new_D6168_;
  assign new_D6147_ = ~new_D6170_ & new_D6171_;
  assign new_D6148_ = new_D6170_ & ~new_D6171_;
  assign new_D6149_ = ~new_D6117_ & new_D6118_;
  assign new_D6150_ = new_D6117_ & ~new_D6118_;
  assign new_D6151_ = ~new_D6133_ | new_D6143_;
  assign new_D6152_ = new_D6133_ & new_D6143_;
  assign new_D6153_ = ~new_D6133_ & ~new_D6143_;
  assign new_D6154_ = new_D6175_ | new_D6174_;
  assign new_D6155_ = new_D6121_ | new_D6154_;
  assign new_D6156_ = new_D6179_ | new_D6178_;
  assign new_D6157_ = ~new_D6121_ & new_D6156_;
  assign new_D6158_ = new_D6177_ | new_D6176_;
  assign new_D6159_ = new_D6121_ & new_D6158_;
  assign new_D6160_ = new_D6119_ & ~new_D6129_;
  assign new_D6161_ = ~new_D6119_ & new_D6129_;
  assign new_D6162_ = ~new_D6118_ | ~new_D6143_;
  assign new_D6163_ = new_D6129_ & new_D6162_;
  assign new_D6164_ = ~new_D6129_ & ~new_D6163_;
  assign new_D6165_ = new_D6129_ | new_D6162_;
  assign new_D6166_ = ~new_D6119_ & new_D6120_;
  assign new_D6167_ = new_D6119_ & ~new_D6120_;
  assign new_D6168_ = new_D6136_ | new_D6173_;
  assign new_D6169_ = ~new_D6136_ & ~new_D6172_;
  assign new_D6170_ = new_D6119_ | new_D6136_;
  assign new_D6171_ = new_D6119_ | new_D6120_;
  assign new_D6172_ = new_D6136_ & new_D6173_;
  assign new_D6173_ = ~new_D6118_ | ~new_D6143_;
  assign new_D6174_ = new_D6151_ & new_D6171_;
  assign new_D6175_ = ~new_D6151_ & ~new_D6171_;
  assign new_D6176_ = new_D6180_ | new_D6181_;
  assign new_D6177_ = ~new_D6122_ & new_D6136_;
  assign new_D6178_ = new_D6182_ | new_D6183_;
  assign new_D6179_ = new_D6122_ & new_D6136_;
  assign new_D6180_ = ~new_D6122_ & ~new_D6136_;
  assign new_D6181_ = new_D6122_ & ~new_D6136_;
  assign new_D6182_ = new_D6122_ & ~new_D6136_;
  assign new_D6183_ = ~new_D6122_ & new_D6136_;
  assign new_D6184_ = new_E6648_;
  assign new_D6185_ = new_E6715_;
  assign new_D6186_ = new_E6782_;
  assign new_D6187_ = new_E6849_;
  assign new_D6188_ = new_E6916_;
  assign new_D6189_ = new_E6983_;
  assign new_D6190_ = new_D6197_ & new_D6196_;
  assign new_D6191_ = new_D6199_ | new_D6198_;
  assign new_D6192_ = new_D6201_ | new_D6200_;
  assign new_D6193_ = new_D6203_ & new_D6202_;
  assign new_D6194_ = new_D6203_ & new_D6204_;
  assign new_D6195_ = new_D6196_ | new_D6205_;
  assign new_D6196_ = new_D6185_ | new_D6208_;
  assign new_D6197_ = new_D6207_ | new_D6206_;
  assign new_D6198_ = new_D6212_ & new_D6211_;
  assign new_D6199_ = new_D6210_ & new_D6209_;
  assign new_D6200_ = new_D6215_ | new_D6214_;
  assign new_D6201_ = new_D6210_ & new_D6213_;
  assign new_D6202_ = new_D6185_ | new_D6218_;
  assign new_D6203_ = new_D6217_ | new_D6216_;
  assign new_D6204_ = new_D6220_ | new_D6219_;
  assign new_D6205_ = ~new_D6196_ & new_D6222_;
  assign new_D6206_ = ~new_D6198_ & new_D6210_;
  assign new_D6207_ = new_D6198_ & ~new_D6210_;
  assign new_D6208_ = new_D6184_ & ~new_D6185_;
  assign new_D6209_ = ~new_D6231_ | ~new_D6232_;
  assign new_D6210_ = new_D6224_ | new_D6226_;
  assign new_D6211_ = new_D6234_ | new_D6233_;
  assign new_D6212_ = new_D6228_ | new_D6227_;
  assign new_D6213_ = ~new_D6236_ | ~new_D6235_;
  assign new_D6214_ = ~new_D6237_ & new_D6238_;
  assign new_D6215_ = new_D6237_ & ~new_D6238_;
  assign new_D6216_ = ~new_D6184_ & new_D6185_;
  assign new_D6217_ = new_D6184_ & ~new_D6185_;
  assign new_D6218_ = ~new_D6200_ | new_D6210_;
  assign new_D6219_ = new_D6200_ & new_D6210_;
  assign new_D6220_ = ~new_D6200_ & ~new_D6210_;
  assign new_D6221_ = new_D6242_ | new_D6241_;
  assign new_D6222_ = new_D6188_ | new_D6221_;
  assign new_D6223_ = new_D6246_ | new_D6245_;
  assign new_D6224_ = ~new_D6188_ & new_D6223_;
  assign new_D6225_ = new_D6244_ | new_D6243_;
  assign new_D6226_ = new_D6188_ & new_D6225_;
  assign new_D6227_ = new_D6186_ & ~new_D6196_;
  assign new_D6228_ = ~new_D6186_ & new_D6196_;
  assign new_D6229_ = ~new_D6185_ | ~new_D6210_;
  assign new_D6230_ = new_D6196_ & new_D6229_;
  assign new_D6231_ = ~new_D6196_ & ~new_D6230_;
  assign new_D6232_ = new_D6196_ | new_D6229_;
  assign new_D6233_ = ~new_D6186_ & new_D6187_;
  assign new_D6234_ = new_D6186_ & ~new_D6187_;
  assign new_D6235_ = new_D6203_ | new_D6240_;
  assign new_D6236_ = ~new_D6203_ & ~new_D6239_;
  assign new_D6237_ = new_D6186_ | new_D6203_;
  assign new_D6238_ = new_D6186_ | new_D6187_;
  assign new_D6239_ = new_D6203_ & new_D6240_;
  assign new_D6240_ = ~new_D6185_ | ~new_D6210_;
  assign new_D6241_ = new_D6218_ & new_D6238_;
  assign new_D6242_ = ~new_D6218_ & ~new_D6238_;
  assign new_D6243_ = new_D6247_ | new_D6248_;
  assign new_D6244_ = ~new_D6189_ & new_D6203_;
  assign new_D6245_ = new_D6249_ | new_D6250_;
  assign new_D6246_ = new_D6189_ & new_D6203_;
  assign new_D6247_ = ~new_D6189_ & ~new_D6203_;
  assign new_D6248_ = new_D6189_ & ~new_D6203_;
  assign new_D6249_ = new_D6189_ & ~new_D6203_;
  assign new_D6250_ = ~new_D6189_ & new_D6203_;
  assign new_D6251_ = new_E7050_;
  assign new_D6252_ = new_E7117_;
  assign new_D6253_ = new_E7184_;
  assign new_D6254_ = new_E7251_;
  assign new_D6255_ = new_E7318_;
  assign new_D6256_ = new_E7385_;
  assign new_D6257_ = new_D6264_ & new_D6263_;
  assign new_D6258_ = new_D6266_ | new_D6265_;
  assign new_D6259_ = new_D6268_ | new_D6267_;
  assign new_D6260_ = new_D6270_ & new_D6269_;
  assign new_D6261_ = new_D6270_ & new_D6271_;
  assign new_D6262_ = new_D6263_ | new_D6272_;
  assign new_D6263_ = new_D6252_ | new_D6275_;
  assign new_D6264_ = new_D6274_ | new_D6273_;
  assign new_D6265_ = new_D6279_ & new_D6278_;
  assign new_D6266_ = new_D6277_ & new_D6276_;
  assign new_D6267_ = new_D6282_ | new_D6281_;
  assign new_D6268_ = new_D6277_ & new_D6280_;
  assign new_D6269_ = new_D6252_ | new_D6285_;
  assign new_D6270_ = new_D6284_ | new_D6283_;
  assign new_D6271_ = new_D6287_ | new_D6286_;
  assign new_D6272_ = ~new_D6263_ & new_D6289_;
  assign new_D6273_ = ~new_D6265_ & new_D6277_;
  assign new_D6274_ = new_D6265_ & ~new_D6277_;
  assign new_D6275_ = new_D6251_ & ~new_D6252_;
  assign new_D6276_ = ~new_D6298_ | ~new_D6299_;
  assign new_D6277_ = new_D6291_ | new_D6293_;
  assign new_D6278_ = new_D6301_ | new_D6300_;
  assign new_D6279_ = new_D6295_ | new_D6294_;
  assign new_D6280_ = ~new_D6303_ | ~new_D6302_;
  assign new_D6281_ = ~new_D6304_ & new_D6305_;
  assign new_D6282_ = new_D6304_ & ~new_D6305_;
  assign new_D6283_ = ~new_D6251_ & new_D6252_;
  assign new_D6284_ = new_D6251_ & ~new_D6252_;
  assign new_D6285_ = ~new_D6267_ | new_D6277_;
  assign new_D6286_ = new_D6267_ & new_D6277_;
  assign new_D6287_ = ~new_D6267_ & ~new_D6277_;
  assign new_D6288_ = new_D6309_ | new_D6308_;
  assign new_D6289_ = new_D6255_ | new_D6288_;
  assign new_D6290_ = new_D6313_ | new_D6312_;
  assign new_D6291_ = ~new_D6255_ & new_D6290_;
  assign new_D6292_ = new_D6311_ | new_D6310_;
  assign new_D6293_ = new_D6255_ & new_D6292_;
  assign new_D6294_ = new_D6253_ & ~new_D6263_;
  assign new_D6295_ = ~new_D6253_ & new_D6263_;
  assign new_D6296_ = ~new_D6252_ | ~new_D6277_;
  assign new_D6297_ = new_D6263_ & new_D6296_;
  assign new_D6298_ = ~new_D6263_ & ~new_D6297_;
  assign new_D6299_ = new_D6263_ | new_D6296_;
  assign new_D6300_ = ~new_D6253_ & new_D6254_;
  assign new_D6301_ = new_D6253_ & ~new_D6254_;
  assign new_D6302_ = new_D6270_ | new_D6307_;
  assign new_D6303_ = ~new_D6270_ & ~new_D6306_;
  assign new_D6304_ = new_D6253_ | new_D6270_;
  assign new_D6305_ = new_D6253_ | new_D6254_;
  assign new_D6306_ = new_D6270_ & new_D6307_;
  assign new_D6307_ = ~new_D6252_ | ~new_D6277_;
  assign new_D6308_ = new_D6285_ & new_D6305_;
  assign new_D6309_ = ~new_D6285_ & ~new_D6305_;
  assign new_D6310_ = new_D6314_ | new_D6315_;
  assign new_D6311_ = ~new_D6256_ & new_D6270_;
  assign new_D6312_ = new_D6316_ | new_D6317_;
  assign new_D6313_ = new_D6256_ & new_D6270_;
  assign new_D6314_ = ~new_D6256_ & ~new_D6270_;
  assign new_D6315_ = new_D6256_ & ~new_D6270_;
  assign new_D6316_ = new_D6256_ & ~new_D6270_;
  assign new_D6317_ = ~new_D6256_ & new_D6270_;
  assign new_D6318_ = new_E7452_;
  assign new_D6319_ = new_E7519_;
  assign new_D6320_ = new_E7586_;
  assign new_D6321_ = new_E7653_;
  assign new_D6322_ = new_E7720_;
  assign new_D6323_ = new_E7787_;
  assign new_D6324_ = new_D6331_ & new_D6330_;
  assign new_D6325_ = new_D6333_ | new_D6332_;
  assign new_D6326_ = new_D6335_ | new_D6334_;
  assign new_D6327_ = new_D6337_ & new_D6336_;
  assign new_D6328_ = new_D6337_ & new_D6338_;
  assign new_D6329_ = new_D6330_ | new_D6339_;
  assign new_D6330_ = new_D6319_ | new_D6342_;
  assign new_D6331_ = new_D6341_ | new_D6340_;
  assign new_D6332_ = new_D6346_ & new_D6345_;
  assign new_D6333_ = new_D6344_ & new_D6343_;
  assign new_D6334_ = new_D6349_ | new_D6348_;
  assign new_D6335_ = new_D6344_ & new_D6347_;
  assign new_D6336_ = new_D6319_ | new_D6352_;
  assign new_D6337_ = new_D6351_ | new_D6350_;
  assign new_D6338_ = new_D6354_ | new_D6353_;
  assign new_D6339_ = ~new_D6330_ & new_D6356_;
  assign new_D6340_ = ~new_D6332_ & new_D6344_;
  assign new_D6341_ = new_D6332_ & ~new_D6344_;
  assign new_D6342_ = new_D6318_ & ~new_D6319_;
  assign new_D6343_ = ~new_D6365_ | ~new_D6366_;
  assign new_D6344_ = new_D6358_ | new_D6360_;
  assign new_D6345_ = new_D6368_ | new_D6367_;
  assign new_D6346_ = new_D6362_ | new_D6361_;
  assign new_D6347_ = ~new_D6370_ | ~new_D6369_;
  assign new_D6348_ = ~new_D6371_ & new_D6372_;
  assign new_D6349_ = new_D6371_ & ~new_D6372_;
  assign new_D6350_ = ~new_D6318_ & new_D6319_;
  assign new_D6351_ = new_D6318_ & ~new_D6319_;
  assign new_D6352_ = ~new_D6334_ | new_D6344_;
  assign new_D6353_ = new_D6334_ & new_D6344_;
  assign new_D6354_ = ~new_D6334_ & ~new_D6344_;
  assign new_D6355_ = new_D6376_ | new_D6375_;
  assign new_D6356_ = new_D6322_ | new_D6355_;
  assign new_D6357_ = new_D6380_ | new_D6379_;
  assign new_D6358_ = ~new_D6322_ & new_D6357_;
  assign new_D6359_ = new_D6378_ | new_D6377_;
  assign new_D6360_ = new_D6322_ & new_D6359_;
  assign new_D6361_ = new_D6320_ & ~new_D6330_;
  assign new_D6362_ = ~new_D6320_ & new_D6330_;
  assign new_D6363_ = ~new_D6319_ | ~new_D6344_;
  assign new_D6364_ = new_D6330_ & new_D6363_;
  assign new_D6365_ = ~new_D6330_ & ~new_D6364_;
  assign new_D6366_ = new_D6330_ | new_D6363_;
  assign new_D6367_ = ~new_D6320_ & new_D6321_;
  assign new_D6368_ = new_D6320_ & ~new_D6321_;
  assign new_D6369_ = new_D6337_ | new_D6374_;
  assign new_D6370_ = ~new_D6337_ & ~new_D6373_;
  assign new_D6371_ = new_D6320_ | new_D6337_;
  assign new_D6372_ = new_D6320_ | new_D6321_;
  assign new_D6373_ = new_D6337_ & new_D6374_;
  assign new_D6374_ = ~new_D6319_ | ~new_D6344_;
  assign new_D6375_ = new_D6352_ & new_D6372_;
  assign new_D6376_ = ~new_D6352_ & ~new_D6372_;
  assign new_D6377_ = new_D6381_ | new_D6382_;
  assign new_D6378_ = ~new_D6323_ & new_D6337_;
  assign new_D6379_ = new_D6383_ | new_D6384_;
  assign new_D6380_ = new_D6323_ & new_D6337_;
  assign new_D6381_ = ~new_D6323_ & ~new_D6337_;
  assign new_D6382_ = new_D6323_ & ~new_D6337_;
  assign new_D6383_ = new_D6323_ & ~new_D6337_;
  assign new_D6384_ = ~new_D6323_ & new_D6337_;
  assign new_D6385_ = new_E7854_;
  assign new_D6386_ = new_E7921_;
  assign new_D6387_ = new_E7988_;
  assign new_D6388_ = new_E8055_;
  assign new_D6389_ = new_E8122_;
  assign new_D6390_ = new_E8189_;
  assign new_D6391_ = new_D6398_ & new_D6397_;
  assign new_D6392_ = new_D6400_ | new_D6399_;
  assign new_D6393_ = new_D6402_ | new_D6401_;
  assign new_D6394_ = new_D6404_ & new_D6403_;
  assign new_D6395_ = new_D6404_ & new_D6405_;
  assign new_D6396_ = new_D6397_ | new_D6406_;
  assign new_D6397_ = new_D6386_ | new_D6409_;
  assign new_D6398_ = new_D6408_ | new_D6407_;
  assign new_D6399_ = new_D6413_ & new_D6412_;
  assign new_D6400_ = new_D6411_ & new_D6410_;
  assign new_D6401_ = new_D6416_ | new_D6415_;
  assign new_D6402_ = new_D6411_ & new_D6414_;
  assign new_D6403_ = new_D6386_ | new_D6419_;
  assign new_D6404_ = new_D6418_ | new_D6417_;
  assign new_D6405_ = new_D6421_ | new_D6420_;
  assign new_D6406_ = ~new_D6397_ & new_D6423_;
  assign new_D6407_ = ~new_D6399_ & new_D6411_;
  assign new_D6408_ = new_D6399_ & ~new_D6411_;
  assign new_D6409_ = new_D6385_ & ~new_D6386_;
  assign new_D6410_ = ~new_D6432_ | ~new_D6433_;
  assign new_D6411_ = new_D6425_ | new_D6427_;
  assign new_D6412_ = new_D6435_ | new_D6434_;
  assign new_D6413_ = new_D6429_ | new_D6428_;
  assign new_D6414_ = ~new_D6437_ | ~new_D6436_;
  assign new_D6415_ = ~new_D6438_ & new_D6439_;
  assign new_D6416_ = new_D6438_ & ~new_D6439_;
  assign new_D6417_ = ~new_D6385_ & new_D6386_;
  assign new_D6418_ = new_D6385_ & ~new_D6386_;
  assign new_D6419_ = ~new_D6401_ | new_D6411_;
  assign new_D6420_ = new_D6401_ & new_D6411_;
  assign new_D6421_ = ~new_D6401_ & ~new_D6411_;
  assign new_D6422_ = new_D6443_ | new_D6442_;
  assign new_D6423_ = new_D6389_ | new_D6422_;
  assign new_D6424_ = new_D6447_ | new_D6446_;
  assign new_D6425_ = ~new_D6389_ & new_D6424_;
  assign new_D6426_ = new_D6445_ | new_D6444_;
  assign new_D6427_ = new_D6389_ & new_D6426_;
  assign new_D6428_ = new_D6387_ & ~new_D6397_;
  assign new_D6429_ = ~new_D6387_ & new_D6397_;
  assign new_D6430_ = ~new_D6386_ | ~new_D6411_;
  assign new_D6431_ = new_D6397_ & new_D6430_;
  assign new_D6432_ = ~new_D6397_ & ~new_D6431_;
  assign new_D6433_ = new_D6397_ | new_D6430_;
  assign new_D6434_ = ~new_D6387_ & new_D6388_;
  assign new_D6435_ = new_D6387_ & ~new_D6388_;
  assign new_D6436_ = new_D6404_ | new_D6441_;
  assign new_D6437_ = ~new_D6404_ & ~new_D6440_;
  assign new_D6438_ = new_D6387_ | new_D6404_;
  assign new_D6439_ = new_D6387_ | new_D6388_;
  assign new_D6440_ = new_D6404_ & new_D6441_;
  assign new_D6441_ = ~new_D6386_ | ~new_D6411_;
  assign new_D6442_ = new_D6419_ & new_D6439_;
  assign new_D6443_ = ~new_D6419_ & ~new_D6439_;
  assign new_D6444_ = new_D6448_ | new_D6449_;
  assign new_D6445_ = ~new_D6390_ & new_D6404_;
  assign new_D6446_ = new_D6450_ | new_D6451_;
  assign new_D6447_ = new_D6390_ & new_D6404_;
  assign new_D6448_ = ~new_D6390_ & ~new_D6404_;
  assign new_D6449_ = new_D6390_ & ~new_D6404_;
  assign new_D6450_ = new_D6390_ & ~new_D6404_;
  assign new_D6451_ = ~new_D6390_ & new_D6404_;
  assign new_D6452_ = new_E8256_;
  assign new_D6453_ = new_E8323_;
  assign new_D6454_ = new_E8390_;
  assign new_D6455_ = new_E8457_;
  assign new_D6456_ = new_E8524_;
  assign new_D6457_ = new_E8591_;
  assign new_D6458_ = new_D6465_ & new_D6464_;
  assign new_D6459_ = new_D6467_ | new_D6466_;
  assign new_D6460_ = new_D6469_ | new_D6468_;
  assign new_D6461_ = new_D6471_ & new_D6470_;
  assign new_D6462_ = new_D6471_ & new_D6472_;
  assign new_D6463_ = new_D6464_ | new_D6473_;
  assign new_D6464_ = new_D6453_ | new_D6476_;
  assign new_D6465_ = new_D6475_ | new_D6474_;
  assign new_D6466_ = new_D6480_ & new_D6479_;
  assign new_D6467_ = new_D6478_ & new_D6477_;
  assign new_D6468_ = new_D6483_ | new_D6482_;
  assign new_D6469_ = new_D6478_ & new_D6481_;
  assign new_D6470_ = new_D6453_ | new_D6486_;
  assign new_D6471_ = new_D6485_ | new_D6484_;
  assign new_D6472_ = new_D6488_ | new_D6487_;
  assign new_D6473_ = ~new_D6464_ & new_D6490_;
  assign new_D6474_ = ~new_D6466_ & new_D6478_;
  assign new_D6475_ = new_D6466_ & ~new_D6478_;
  assign new_D6476_ = new_D6452_ & ~new_D6453_;
  assign new_D6477_ = ~new_D6499_ | ~new_D6500_;
  assign new_D6478_ = new_D6492_ | new_D6494_;
  assign new_D6479_ = new_D6502_ | new_D6501_;
  assign new_D6480_ = new_D6496_ | new_D6495_;
  assign new_D6481_ = ~new_D6504_ | ~new_D6503_;
  assign new_D6482_ = ~new_D6505_ & new_D6506_;
  assign new_D6483_ = new_D6505_ & ~new_D6506_;
  assign new_D6484_ = ~new_D6452_ & new_D6453_;
  assign new_D6485_ = new_D6452_ & ~new_D6453_;
  assign new_D6486_ = ~new_D6468_ | new_D6478_;
  assign new_D6487_ = new_D6468_ & new_D6478_;
  assign new_D6488_ = ~new_D6468_ & ~new_D6478_;
  assign new_D6489_ = new_D6510_ | new_D6509_;
  assign new_D6490_ = new_D6456_ | new_D6489_;
  assign new_D6491_ = new_D6514_ | new_D6513_;
  assign new_D6492_ = ~new_D6456_ & new_D6491_;
  assign new_D6493_ = new_D6512_ | new_D6511_;
  assign new_D6494_ = new_D6456_ & new_D6493_;
  assign new_D6495_ = new_D6454_ & ~new_D6464_;
  assign new_D6496_ = ~new_D6454_ & new_D6464_;
  assign new_D6497_ = ~new_D6453_ | ~new_D6478_;
  assign new_D6498_ = new_D6464_ & new_D6497_;
  assign new_D6499_ = ~new_D6464_ & ~new_D6498_;
  assign new_D6500_ = new_D6464_ | new_D6497_;
  assign new_D6501_ = ~new_D6454_ & new_D6455_;
  assign new_D6502_ = new_D6454_ & ~new_D6455_;
  assign new_D6503_ = new_D6471_ | new_D6508_;
  assign new_D6504_ = ~new_D6471_ & ~new_D6507_;
  assign new_D6505_ = new_D6454_ | new_D6471_;
  assign new_D6506_ = new_D6454_ | new_D6455_;
  assign new_D6507_ = new_D6471_ & new_D6508_;
  assign new_D6508_ = ~new_D6453_ | ~new_D6478_;
  assign new_D6509_ = new_D6486_ & new_D6506_;
  assign new_D6510_ = ~new_D6486_ & ~new_D6506_;
  assign new_D6511_ = new_D6515_ | new_D6516_;
  assign new_D6512_ = ~new_D6457_ & new_D6471_;
  assign new_D6513_ = new_D6517_ | new_D6518_;
  assign new_D6514_ = new_D6457_ & new_D6471_;
  assign new_D6515_ = ~new_D6457_ & ~new_D6471_;
  assign new_D6516_ = new_D6457_ & ~new_D6471_;
  assign new_D6517_ = new_D6457_ & ~new_D6471_;
  assign new_D6518_ = ~new_D6457_ & new_D6471_;
  assign new_D6519_ = new_E8658_;
  assign new_D6520_ = new_E8725_;
  assign new_D6521_ = new_E8792_;
  assign new_D6522_ = new_E8859_;
  assign new_D6523_ = new_E8926_;
  assign new_D6524_ = new_E8993_;
  assign new_D6525_ = new_D6532_ & new_D6531_;
  assign new_D6526_ = new_D6534_ | new_D6533_;
  assign new_D6527_ = new_D6536_ | new_D6535_;
  assign new_D6528_ = new_D6538_ & new_D6537_;
  assign new_D6529_ = new_D6538_ & new_D6539_;
  assign new_D6530_ = new_D6531_ | new_D6540_;
  assign new_D6531_ = new_D6520_ | new_D6543_;
  assign new_D6532_ = new_D6542_ | new_D6541_;
  assign new_D6533_ = new_D6547_ & new_D6546_;
  assign new_D6534_ = new_D6545_ & new_D6544_;
  assign new_D6535_ = new_D6550_ | new_D6549_;
  assign new_D6536_ = new_D6545_ & new_D6548_;
  assign new_D6537_ = new_D6520_ | new_D6553_;
  assign new_D6538_ = new_D6552_ | new_D6551_;
  assign new_D6539_ = new_D6555_ | new_D6554_;
  assign new_D6540_ = ~new_D6531_ & new_D6557_;
  assign new_D6541_ = ~new_D6533_ & new_D6545_;
  assign new_D6542_ = new_D6533_ & ~new_D6545_;
  assign new_D6543_ = new_D6519_ & ~new_D6520_;
  assign new_D6544_ = ~new_D6566_ | ~new_D6567_;
  assign new_D6545_ = new_D6559_ | new_D6561_;
  assign new_D6546_ = new_D6569_ | new_D6568_;
  assign new_D6547_ = new_D6563_ | new_D6562_;
  assign new_D6548_ = ~new_D6571_ | ~new_D6570_;
  assign new_D6549_ = ~new_D6572_ & new_D6573_;
  assign new_D6550_ = new_D6572_ & ~new_D6573_;
  assign new_D6551_ = ~new_D6519_ & new_D6520_;
  assign new_D6552_ = new_D6519_ & ~new_D6520_;
  assign new_D6553_ = ~new_D6535_ | new_D6545_;
  assign new_D6554_ = new_D6535_ & new_D6545_;
  assign new_D6555_ = ~new_D6535_ & ~new_D6545_;
  assign new_D6556_ = new_D6577_ | new_D6576_;
  assign new_D6557_ = new_D6523_ | new_D6556_;
  assign new_D6558_ = new_D6581_ | new_D6580_;
  assign new_D6559_ = ~new_D6523_ & new_D6558_;
  assign new_D6560_ = new_D6579_ | new_D6578_;
  assign new_D6561_ = new_D6523_ & new_D6560_;
  assign new_D6562_ = new_D6521_ & ~new_D6531_;
  assign new_D6563_ = ~new_D6521_ & new_D6531_;
  assign new_D6564_ = ~new_D6520_ | ~new_D6545_;
  assign new_D6565_ = new_D6531_ & new_D6564_;
  assign new_D6566_ = ~new_D6531_ & ~new_D6565_;
  assign new_D6567_ = new_D6531_ | new_D6564_;
  assign new_D6568_ = ~new_D6521_ & new_D6522_;
  assign new_D6569_ = new_D6521_ & ~new_D6522_;
  assign new_D6570_ = new_D6538_ | new_D6575_;
  assign new_D6571_ = ~new_D6538_ & ~new_D6574_;
  assign new_D6572_ = new_D6521_ | new_D6538_;
  assign new_D6573_ = new_D6521_ | new_D6522_;
  assign new_D6574_ = new_D6538_ & new_D6575_;
  assign new_D6575_ = ~new_D6520_ | ~new_D6545_;
  assign new_D6576_ = new_D6553_ & new_D6573_;
  assign new_D6577_ = ~new_D6553_ & ~new_D6573_;
  assign new_D6578_ = new_D6582_ | new_D6583_;
  assign new_D6579_ = ~new_D6524_ & new_D6538_;
  assign new_D6580_ = new_D6584_ | new_D6585_;
  assign new_D6581_ = new_D6524_ & new_D6538_;
  assign new_D6582_ = ~new_D6524_ & ~new_D6538_;
  assign new_D6583_ = new_D6524_ & ~new_D6538_;
  assign new_D6584_ = new_D6524_ & ~new_D6538_;
  assign new_D6585_ = ~new_D6524_ & new_D6538_;
  assign new_D6586_ = new_E9060_;
  assign new_D6587_ = new_E9127_;
  assign new_D6588_ = new_E9194_;
  assign new_D6589_ = new_E9261_;
  assign new_D6590_ = new_E9328_;
  assign new_D6591_ = new_E9395_;
  assign new_D6592_ = new_D6599_ & new_D6598_;
  assign new_D6593_ = new_D6601_ | new_D6600_;
  assign new_D6594_ = new_D6603_ | new_D6602_;
  assign new_D6595_ = new_D6605_ & new_D6604_;
  assign new_D6596_ = new_D6605_ & new_D6606_;
  assign new_D6597_ = new_D6598_ | new_D6607_;
  assign new_D6598_ = new_D6587_ | new_D6610_;
  assign new_D6599_ = new_D6609_ | new_D6608_;
  assign new_D6600_ = new_D6614_ & new_D6613_;
  assign new_D6601_ = new_D6612_ & new_D6611_;
  assign new_D6602_ = new_D6617_ | new_D6616_;
  assign new_D6603_ = new_D6612_ & new_D6615_;
  assign new_D6604_ = new_D6587_ | new_D6620_;
  assign new_D6605_ = new_D6619_ | new_D6618_;
  assign new_D6606_ = new_D6622_ | new_D6621_;
  assign new_D6607_ = ~new_D6598_ & new_D6624_;
  assign new_D6608_ = ~new_D6600_ & new_D6612_;
  assign new_D6609_ = new_D6600_ & ~new_D6612_;
  assign new_D6610_ = new_D6586_ & ~new_D6587_;
  assign new_D6611_ = ~new_D6633_ | ~new_D6634_;
  assign new_D6612_ = new_D6626_ | new_D6628_;
  assign new_D6613_ = new_D6636_ | new_D6635_;
  assign new_D6614_ = new_D6630_ | new_D6629_;
  assign new_D6615_ = ~new_D6638_ | ~new_D6637_;
  assign new_D6616_ = ~new_D6639_ & new_D6640_;
  assign new_D6617_ = new_D6639_ & ~new_D6640_;
  assign new_D6618_ = ~new_D6586_ & new_D6587_;
  assign new_D6619_ = new_D6586_ & ~new_D6587_;
  assign new_D6620_ = ~new_D6602_ | new_D6612_;
  assign new_D6621_ = new_D6602_ & new_D6612_;
  assign new_D6622_ = ~new_D6602_ & ~new_D6612_;
  assign new_D6623_ = new_D6644_ | new_D6643_;
  assign new_D6624_ = new_D6590_ | new_D6623_;
  assign new_D6625_ = new_D6648_ | new_D6647_;
  assign new_D6626_ = ~new_D6590_ & new_D6625_;
  assign new_D6627_ = new_D6646_ | new_D6645_;
  assign new_D6628_ = new_D6590_ & new_D6627_;
  assign new_D6629_ = new_D6588_ & ~new_D6598_;
  assign new_D6630_ = ~new_D6588_ & new_D6598_;
  assign new_D6631_ = ~new_D6587_ | ~new_D6612_;
  assign new_D6632_ = new_D6598_ & new_D6631_;
  assign new_D6633_ = ~new_D6598_ & ~new_D6632_;
  assign new_D6634_ = new_D6598_ | new_D6631_;
  assign new_D6635_ = ~new_D6588_ & new_D6589_;
  assign new_D6636_ = new_D6588_ & ~new_D6589_;
  assign new_D6637_ = new_D6605_ | new_D6642_;
  assign new_D6638_ = ~new_D6605_ & ~new_D6641_;
  assign new_D6639_ = new_D6588_ | new_D6605_;
  assign new_D6640_ = new_D6588_ | new_D6589_;
  assign new_D6641_ = new_D6605_ & new_D6642_;
  assign new_D6642_ = ~new_D6587_ | ~new_D6612_;
  assign new_D6643_ = new_D6620_ & new_D6640_;
  assign new_D6644_ = ~new_D6620_ & ~new_D6640_;
  assign new_D6645_ = new_D6649_ | new_D6650_;
  assign new_D6646_ = ~new_D6591_ & new_D6605_;
  assign new_D6647_ = new_D6651_ | new_D6652_;
  assign new_D6648_ = new_D6591_ & new_D6605_;
  assign new_D6649_ = ~new_D6591_ & ~new_D6605_;
  assign new_D6650_ = new_D6591_ & ~new_D6605_;
  assign new_D6651_ = new_D6591_ & ~new_D6605_;
  assign new_D6652_ = ~new_D6591_ & new_D6605_;
  assign new_D6653_ = new_E9462_;
  assign new_D6654_ = new_E9529_;
  assign new_D6655_ = new_E9596_;
  assign new_D6656_ = new_E9663_;
  assign new_D6657_ = new_E9730_;
  assign new_D6658_ = new_E9797_;
  assign new_D6659_ = new_D6666_ & new_D6665_;
  assign new_D6660_ = new_D6668_ | new_D6667_;
  assign new_D6661_ = new_D6670_ | new_D6669_;
  assign new_D6662_ = new_D6672_ & new_D6671_;
  assign new_D6663_ = new_D6672_ & new_D6673_;
  assign new_D6664_ = new_D6665_ | new_D6674_;
  assign new_D6665_ = new_D6654_ | new_D6677_;
  assign new_D6666_ = new_D6676_ | new_D6675_;
  assign new_D6667_ = new_D6681_ & new_D6680_;
  assign new_D6668_ = new_D6679_ & new_D6678_;
  assign new_D6669_ = new_D6684_ | new_D6683_;
  assign new_D6670_ = new_D6679_ & new_D6682_;
  assign new_D6671_ = new_D6654_ | new_D6687_;
  assign new_D6672_ = new_D6686_ | new_D6685_;
  assign new_D6673_ = new_D6689_ | new_D6688_;
  assign new_D6674_ = ~new_D6665_ & new_D6691_;
  assign new_D6675_ = ~new_D6667_ & new_D6679_;
  assign new_D6676_ = new_D6667_ & ~new_D6679_;
  assign new_D6677_ = new_D6653_ & ~new_D6654_;
  assign new_D6678_ = ~new_D6700_ | ~new_D6701_;
  assign new_D6679_ = new_D6693_ | new_D6695_;
  assign new_D6680_ = new_D6703_ | new_D6702_;
  assign new_D6681_ = new_D6697_ | new_D6696_;
  assign new_D6682_ = ~new_D6705_ | ~new_D6704_;
  assign new_D6683_ = ~new_D6706_ & new_D6707_;
  assign new_D6684_ = new_D6706_ & ~new_D6707_;
  assign new_D6685_ = ~new_D6653_ & new_D6654_;
  assign new_D6686_ = new_D6653_ & ~new_D6654_;
  assign new_D6687_ = ~new_D6669_ | new_D6679_;
  assign new_D6688_ = new_D6669_ & new_D6679_;
  assign new_D6689_ = ~new_D6669_ & ~new_D6679_;
  assign new_D6690_ = new_D6711_ | new_D6710_;
  assign new_D6691_ = new_D6657_ | new_D6690_;
  assign new_D6692_ = new_D6715_ | new_D6714_;
  assign new_D6693_ = ~new_D6657_ & new_D6692_;
  assign new_D6694_ = new_D6713_ | new_D6712_;
  assign new_D6695_ = new_D6657_ & new_D6694_;
  assign new_D6696_ = new_D6655_ & ~new_D6665_;
  assign new_D6697_ = ~new_D6655_ & new_D6665_;
  assign new_D6698_ = ~new_D6654_ | ~new_D6679_;
  assign new_D6699_ = new_D6665_ & new_D6698_;
  assign new_D6700_ = ~new_D6665_ & ~new_D6699_;
  assign new_D6701_ = new_D6665_ | new_D6698_;
  assign new_D6702_ = ~new_D6655_ & new_D6656_;
  assign new_D6703_ = new_D6655_ & ~new_D6656_;
  assign new_D6704_ = new_D6672_ | new_D6709_;
  assign new_D6705_ = ~new_D6672_ & ~new_D6708_;
  assign new_D6706_ = new_D6655_ | new_D6672_;
  assign new_D6707_ = new_D6655_ | new_D6656_;
  assign new_D6708_ = new_D6672_ & new_D6709_;
  assign new_D6709_ = ~new_D6654_ | ~new_D6679_;
  assign new_D6710_ = new_D6687_ & new_D6707_;
  assign new_D6711_ = ~new_D6687_ & ~new_D6707_;
  assign new_D6712_ = new_D6716_ | new_D6717_;
  assign new_D6713_ = ~new_D6658_ & new_D6672_;
  assign new_D6714_ = new_D6718_ | new_D6719_;
  assign new_D6715_ = new_D6658_ & new_D6672_;
  assign new_D6716_ = ~new_D6658_ & ~new_D6672_;
  assign new_D6717_ = new_D6658_ & ~new_D6672_;
  assign new_D6718_ = new_D6658_ & ~new_D6672_;
  assign new_D6719_ = ~new_D6658_ & new_D6672_;
  assign new_D6720_ = new_E9864_;
  assign new_D6721_ = new_E9931_;
  assign new_D6722_ = new_E9998_;
  assign new_D6723_ = new_F66_;
  assign new_D6724_ = new_F133_;
  assign new_D6725_ = new_F200_;
  assign new_D6726_ = new_D6733_ & new_D6732_;
  assign new_D6727_ = new_D6735_ | new_D6734_;
  assign new_D6728_ = new_D6737_ | new_D6736_;
  assign new_D6729_ = new_D6739_ & new_D6738_;
  assign new_D6730_ = new_D6739_ & new_D6740_;
  assign new_D6731_ = new_D6732_ | new_D6741_;
  assign new_D6732_ = new_D6721_ | new_D6744_;
  assign new_D6733_ = new_D6743_ | new_D6742_;
  assign new_D6734_ = new_D6748_ & new_D6747_;
  assign new_D6735_ = new_D6746_ & new_D6745_;
  assign new_D6736_ = new_D6751_ | new_D6750_;
  assign new_D6737_ = new_D6746_ & new_D6749_;
  assign new_D6738_ = new_D6721_ | new_D6754_;
  assign new_D6739_ = new_D6753_ | new_D6752_;
  assign new_D6740_ = new_D6756_ | new_D6755_;
  assign new_D6741_ = ~new_D6732_ & new_D6758_;
  assign new_D6742_ = ~new_D6734_ & new_D6746_;
  assign new_D6743_ = new_D6734_ & ~new_D6746_;
  assign new_D6744_ = new_D6720_ & ~new_D6721_;
  assign new_D6745_ = ~new_D6767_ | ~new_D6768_;
  assign new_D6746_ = new_D6760_ | new_D6762_;
  assign new_D6747_ = new_D6770_ | new_D6769_;
  assign new_D6748_ = new_D6764_ | new_D6763_;
  assign new_D6749_ = ~new_D6772_ | ~new_D6771_;
  assign new_D6750_ = ~new_D6773_ & new_D6774_;
  assign new_D6751_ = new_D6773_ & ~new_D6774_;
  assign new_D6752_ = ~new_D6720_ & new_D6721_;
  assign new_D6753_ = new_D6720_ & ~new_D6721_;
  assign new_D6754_ = ~new_D6736_ | new_D6746_;
  assign new_D6755_ = new_D6736_ & new_D6746_;
  assign new_D6756_ = ~new_D6736_ & ~new_D6746_;
  assign new_D6757_ = new_D6778_ | new_D6777_;
  assign new_D6758_ = new_D6724_ | new_D6757_;
  assign new_D6759_ = new_D6782_ | new_D6781_;
  assign new_D6760_ = ~new_D6724_ & new_D6759_;
  assign new_D6761_ = new_D6780_ | new_D6779_;
  assign new_D6762_ = new_D6724_ & new_D6761_;
  assign new_D6763_ = new_D6722_ & ~new_D6732_;
  assign new_D6764_ = ~new_D6722_ & new_D6732_;
  assign new_D6765_ = ~new_D6721_ | ~new_D6746_;
  assign new_D6766_ = new_D6732_ & new_D6765_;
  assign new_D6767_ = ~new_D6732_ & ~new_D6766_;
  assign new_D6768_ = new_D6732_ | new_D6765_;
  assign new_D6769_ = ~new_D6722_ & new_D6723_;
  assign new_D6770_ = new_D6722_ & ~new_D6723_;
  assign new_D6771_ = new_D6739_ | new_D6776_;
  assign new_D6772_ = ~new_D6739_ & ~new_D6775_;
  assign new_D6773_ = new_D6722_ | new_D6739_;
  assign new_D6774_ = new_D6722_ | new_D6723_;
  assign new_D6775_ = new_D6739_ & new_D6776_;
  assign new_D6776_ = ~new_D6721_ | ~new_D6746_;
  assign new_D6777_ = new_D6754_ & new_D6774_;
  assign new_D6778_ = ~new_D6754_ & ~new_D6774_;
  assign new_D6779_ = new_D6783_ | new_D6784_;
  assign new_D6780_ = ~new_D6725_ & new_D6739_;
  assign new_D6781_ = new_D6785_ | new_D6786_;
  assign new_D6782_ = new_D6725_ & new_D6739_;
  assign new_D6783_ = ~new_D6725_ & ~new_D6739_;
  assign new_D6784_ = new_D6725_ & ~new_D6739_;
  assign new_D6785_ = new_D6725_ & ~new_D6739_;
  assign new_D6786_ = ~new_D6725_ & new_D6739_;
  assign new_D6787_ = new_F267_;
  assign new_D6788_ = new_F334_;
  assign new_D6789_ = new_F401_;
  assign new_D6790_ = new_F468_;
  assign new_D6791_ = new_F535_;
  assign new_D6792_ = new_F602_;
  assign new_D6793_ = new_D6800_ & new_D6799_;
  assign new_D6794_ = new_D6802_ | new_D6801_;
  assign new_D6795_ = new_D6804_ | new_D6803_;
  assign new_D6796_ = new_D6806_ & new_D6805_;
  assign new_D6797_ = new_D6806_ & new_D6807_;
  assign new_D6798_ = new_D6799_ | new_D6808_;
  assign new_D6799_ = new_D6788_ | new_D6811_;
  assign new_D6800_ = new_D6810_ | new_D6809_;
  assign new_D6801_ = new_D6815_ & new_D6814_;
  assign new_D6802_ = new_D6813_ & new_D6812_;
  assign new_D6803_ = new_D6818_ | new_D6817_;
  assign new_D6804_ = new_D6813_ & new_D6816_;
  assign new_D6805_ = new_D6788_ | new_D6821_;
  assign new_D6806_ = new_D6820_ | new_D6819_;
  assign new_D6807_ = new_D6823_ | new_D6822_;
  assign new_D6808_ = ~new_D6799_ & new_D6825_;
  assign new_D6809_ = ~new_D6801_ & new_D6813_;
  assign new_D6810_ = new_D6801_ & ~new_D6813_;
  assign new_D6811_ = new_D6787_ & ~new_D6788_;
  assign new_D6812_ = ~new_D6834_ | ~new_D6835_;
  assign new_D6813_ = new_D6827_ | new_D6829_;
  assign new_D6814_ = new_D6837_ | new_D6836_;
  assign new_D6815_ = new_D6831_ | new_D6830_;
  assign new_D6816_ = ~new_D6839_ | ~new_D6838_;
  assign new_D6817_ = ~new_D6840_ & new_D6841_;
  assign new_D6818_ = new_D6840_ & ~new_D6841_;
  assign new_D6819_ = ~new_D6787_ & new_D6788_;
  assign new_D6820_ = new_D6787_ & ~new_D6788_;
  assign new_D6821_ = ~new_D6803_ | new_D6813_;
  assign new_D6822_ = new_D6803_ & new_D6813_;
  assign new_D6823_ = ~new_D6803_ & ~new_D6813_;
  assign new_D6824_ = new_D6845_ | new_D6844_;
  assign new_D6825_ = new_D6791_ | new_D6824_;
  assign new_D6826_ = new_D6849_ | new_D6848_;
  assign new_D6827_ = ~new_D6791_ & new_D6826_;
  assign new_D6828_ = new_D6847_ | new_D6846_;
  assign new_D6829_ = new_D6791_ & new_D6828_;
  assign new_D6830_ = new_D6789_ & ~new_D6799_;
  assign new_D6831_ = ~new_D6789_ & new_D6799_;
  assign new_D6832_ = ~new_D6788_ | ~new_D6813_;
  assign new_D6833_ = new_D6799_ & new_D6832_;
  assign new_D6834_ = ~new_D6799_ & ~new_D6833_;
  assign new_D6835_ = new_D6799_ | new_D6832_;
  assign new_D6836_ = ~new_D6789_ & new_D6790_;
  assign new_D6837_ = new_D6789_ & ~new_D6790_;
  assign new_D6838_ = new_D6806_ | new_D6843_;
  assign new_D6839_ = ~new_D6806_ & ~new_D6842_;
  assign new_D6840_ = new_D6789_ | new_D6806_;
  assign new_D6841_ = new_D6789_ | new_D6790_;
  assign new_D6842_ = new_D6806_ & new_D6843_;
  assign new_D6843_ = ~new_D6788_ | ~new_D6813_;
  assign new_D6844_ = new_D6821_ & new_D6841_;
  assign new_D6845_ = ~new_D6821_ & ~new_D6841_;
  assign new_D6846_ = new_D6850_ | new_D6851_;
  assign new_D6847_ = ~new_D6792_ & new_D6806_;
  assign new_D6848_ = new_D6852_ | new_D6853_;
  assign new_D6849_ = new_D6792_ & new_D6806_;
  assign new_D6850_ = ~new_D6792_ & ~new_D6806_;
  assign new_D6851_ = new_D6792_ & ~new_D6806_;
  assign new_D6852_ = new_D6792_ & ~new_D6806_;
  assign new_D6853_ = ~new_D6792_ & new_D6806_;
  assign new_D6854_ = new_F669_;
  assign new_D6855_ = new_F736_;
  assign new_D6856_ = new_F803_;
  assign new_D6857_ = new_F870_;
  assign new_D6858_ = new_F937_;
  assign new_D6859_ = new_F1004_;
  assign new_D6860_ = new_D6867_ & new_D6866_;
  assign new_D6861_ = new_D6869_ | new_D6868_;
  assign new_D6862_ = new_D6871_ | new_D6870_;
  assign new_D6863_ = new_D6873_ & new_D6872_;
  assign new_D6864_ = new_D6873_ & new_D6874_;
  assign new_D6865_ = new_D6866_ | new_D6875_;
  assign new_D6866_ = new_D6855_ | new_D6878_;
  assign new_D6867_ = new_D6877_ | new_D6876_;
  assign new_D6868_ = new_D6882_ & new_D6881_;
  assign new_D6869_ = new_D6880_ & new_D6879_;
  assign new_D6870_ = new_D6885_ | new_D6884_;
  assign new_D6871_ = new_D6880_ & new_D6883_;
  assign new_D6872_ = new_D6855_ | new_D6888_;
  assign new_D6873_ = new_D6887_ | new_D6886_;
  assign new_D6874_ = new_D6890_ | new_D6889_;
  assign new_D6875_ = ~new_D6866_ & new_D6892_;
  assign new_D6876_ = ~new_D6868_ & new_D6880_;
  assign new_D6877_ = new_D6868_ & ~new_D6880_;
  assign new_D6878_ = new_D6854_ & ~new_D6855_;
  assign new_D6879_ = ~new_D6901_ | ~new_D6902_;
  assign new_D6880_ = new_D6894_ | new_D6896_;
  assign new_D6881_ = new_D6904_ | new_D6903_;
  assign new_D6882_ = new_D6898_ | new_D6897_;
  assign new_D6883_ = ~new_D6906_ | ~new_D6905_;
  assign new_D6884_ = ~new_D6907_ & new_D6908_;
  assign new_D6885_ = new_D6907_ & ~new_D6908_;
  assign new_D6886_ = ~new_D6854_ & new_D6855_;
  assign new_D6887_ = new_D6854_ & ~new_D6855_;
  assign new_D6888_ = ~new_D6870_ | new_D6880_;
  assign new_D6889_ = new_D6870_ & new_D6880_;
  assign new_D6890_ = ~new_D6870_ & ~new_D6880_;
  assign new_D6891_ = new_D6912_ | new_D6911_;
  assign new_D6892_ = new_D6858_ | new_D6891_;
  assign new_D6893_ = new_D6916_ | new_D6915_;
  assign new_D6894_ = ~new_D6858_ & new_D6893_;
  assign new_D6895_ = new_D6914_ | new_D6913_;
  assign new_D6896_ = new_D6858_ & new_D6895_;
  assign new_D6897_ = new_D6856_ & ~new_D6866_;
  assign new_D6898_ = ~new_D6856_ & new_D6866_;
  assign new_D6899_ = ~new_D6855_ | ~new_D6880_;
  assign new_D6900_ = new_D6866_ & new_D6899_;
  assign new_D6901_ = ~new_D6866_ & ~new_D6900_;
  assign new_D6902_ = new_D6866_ | new_D6899_;
  assign new_D6903_ = ~new_D6856_ & new_D6857_;
  assign new_D6904_ = new_D6856_ & ~new_D6857_;
  assign new_D6905_ = new_D6873_ | new_D6910_;
  assign new_D6906_ = ~new_D6873_ & ~new_D6909_;
  assign new_D6907_ = new_D6856_ | new_D6873_;
  assign new_D6908_ = new_D6856_ | new_D6857_;
  assign new_D6909_ = new_D6873_ & new_D6910_;
  assign new_D6910_ = ~new_D6855_ | ~new_D6880_;
  assign new_D6911_ = new_D6888_ & new_D6908_;
  assign new_D6912_ = ~new_D6888_ & ~new_D6908_;
  assign new_D6913_ = new_D6917_ | new_D6918_;
  assign new_D6914_ = ~new_D6859_ & new_D6873_;
  assign new_D6915_ = new_D6919_ | new_D6920_;
  assign new_D6916_ = new_D6859_ & new_D6873_;
  assign new_D6917_ = ~new_D6859_ & ~new_D6873_;
  assign new_D6918_ = new_D6859_ & ~new_D6873_;
  assign new_D6919_ = new_D6859_ & ~new_D6873_;
  assign new_D6920_ = ~new_D6859_ & new_D6873_;
  assign new_D6921_ = new_F1071_;
  assign new_D6922_ = new_F1138_;
  assign new_D6923_ = new_F1205_;
  assign new_D6924_ = new_F1272_;
  assign new_D6925_ = new_F1339_;
  assign new_D6926_ = new_F1406_;
  assign new_D6927_ = new_D6934_ & new_D6933_;
  assign new_D6928_ = new_D6936_ | new_D6935_;
  assign new_D6929_ = new_D6938_ | new_D6937_;
  assign new_D6930_ = new_D6940_ & new_D6939_;
  assign new_D6931_ = new_D6940_ & new_D6941_;
  assign new_D6932_ = new_D6933_ | new_D6942_;
  assign new_D6933_ = new_D6922_ | new_D6945_;
  assign new_D6934_ = new_D6944_ | new_D6943_;
  assign new_D6935_ = new_D6949_ & new_D6948_;
  assign new_D6936_ = new_D6947_ & new_D6946_;
  assign new_D6937_ = new_D6952_ | new_D6951_;
  assign new_D6938_ = new_D6947_ & new_D6950_;
  assign new_D6939_ = new_D6922_ | new_D6955_;
  assign new_D6940_ = new_D6954_ | new_D6953_;
  assign new_D6941_ = new_D6957_ | new_D6956_;
  assign new_D6942_ = ~new_D6933_ & new_D6959_;
  assign new_D6943_ = ~new_D6935_ & new_D6947_;
  assign new_D6944_ = new_D6935_ & ~new_D6947_;
  assign new_D6945_ = new_D6921_ & ~new_D6922_;
  assign new_D6946_ = ~new_D6968_ | ~new_D6969_;
  assign new_D6947_ = new_D6961_ | new_D6963_;
  assign new_D6948_ = new_D6971_ | new_D6970_;
  assign new_D6949_ = new_D6965_ | new_D6964_;
  assign new_D6950_ = ~new_D6973_ | ~new_D6972_;
  assign new_D6951_ = ~new_D6974_ & new_D6975_;
  assign new_D6952_ = new_D6974_ & ~new_D6975_;
  assign new_D6953_ = ~new_D6921_ & new_D6922_;
  assign new_D6954_ = new_D6921_ & ~new_D6922_;
  assign new_D6955_ = ~new_D6937_ | new_D6947_;
  assign new_D6956_ = new_D6937_ & new_D6947_;
  assign new_D6957_ = ~new_D6937_ & ~new_D6947_;
  assign new_D6958_ = new_D6979_ | new_D6978_;
  assign new_D6959_ = new_D6925_ | new_D6958_;
  assign new_D6960_ = new_D6983_ | new_D6982_;
  assign new_D6961_ = ~new_D6925_ & new_D6960_;
  assign new_D6962_ = new_D6981_ | new_D6980_;
  assign new_D6963_ = new_D6925_ & new_D6962_;
  assign new_D6964_ = new_D6923_ & ~new_D6933_;
  assign new_D6965_ = ~new_D6923_ & new_D6933_;
  assign new_D6966_ = ~new_D6922_ | ~new_D6947_;
  assign new_D6967_ = new_D6933_ & new_D6966_;
  assign new_D6968_ = ~new_D6933_ & ~new_D6967_;
  assign new_D6969_ = new_D6933_ | new_D6966_;
  assign new_D6970_ = ~new_D6923_ & new_D6924_;
  assign new_D6971_ = new_D6923_ & ~new_D6924_;
  assign new_D6972_ = new_D6940_ | new_D6977_;
  assign new_D6973_ = ~new_D6940_ & ~new_D6976_;
  assign new_D6974_ = new_D6923_ | new_D6940_;
  assign new_D6975_ = new_D6923_ | new_D6924_;
  assign new_D6976_ = new_D6940_ & new_D6977_;
  assign new_D6977_ = ~new_D6922_ | ~new_D6947_;
  assign new_D6978_ = new_D6955_ & new_D6975_;
  assign new_D6979_ = ~new_D6955_ & ~new_D6975_;
  assign new_D6980_ = new_D6984_ | new_D6985_;
  assign new_D6981_ = ~new_D6926_ & new_D6940_;
  assign new_D6982_ = new_D6986_ | new_D6987_;
  assign new_D6983_ = new_D6926_ & new_D6940_;
  assign new_D6984_ = ~new_D6926_ & ~new_D6940_;
  assign new_D6985_ = new_D6926_ & ~new_D6940_;
  assign new_D6986_ = new_D6926_ & ~new_D6940_;
  assign new_D6987_ = ~new_D6926_ & new_D6940_;
  assign new_C2514_ = ~new_C2453_ & new_C2467_;
  assign new_C2513_ = new_C2453_ & ~new_C2467_;
  assign new_C2512_ = new_C2453_ & ~new_C2467_;
  assign new_C2511_ = ~new_C2453_ & ~new_C2467_;
  assign new_C2510_ = new_C2453_ & new_C2467_;
  assign new_C2509_ = new_C2513_ | new_C2514_;
  assign new_C2508_ = ~new_C2453_ & new_C2467_;
  assign new_C2507_ = new_C2511_ | new_C2512_;
  assign new_C2506_ = ~new_C2482_ & ~new_C2502_;
  assign new_C2505_ = new_C2482_ & new_C2502_;
  assign new_C2504_ = ~new_C2449_ | ~new_C2474_;
  assign new_C2503_ = new_C2467_ & new_C2504_;
  assign new_C2502_ = new_C2450_ | new_C2451_;
  assign new_C2501_ = new_C2450_ | new_C2467_;
  assign new_C2500_ = ~new_C2467_ & ~new_C2503_;
  assign new_C2499_ = new_C2467_ | new_C2504_;
  assign new_C2498_ = new_C2450_ & ~new_C2451_;
  assign new_C2497_ = ~new_C2450_ & new_C2451_;
  assign new_C2496_ = new_C2460_ | new_C2493_;
  assign new_C2495_ = ~new_C2460_ & ~new_C2494_;
  assign new_C2494_ = new_C2460_ & new_C2493_;
  assign new_C2493_ = ~new_C2449_ | ~new_C2474_;
  assign new_C2492_ = ~new_C2450_ & new_C2460_;
  assign new_C2491_ = new_C2450_ & ~new_C2460_;
  assign new_C2490_ = new_C2452_ & new_C2489_;
  assign new_C2489_ = new_C2508_ | new_C2507_;
  assign new_C2488_ = ~new_C2452_ & new_C2487_;
  assign new_C2487_ = new_C2510_ | new_C2509_;
  assign new_C2486_ = new_C2452_ | new_C2485_;
  assign new_C2485_ = new_C2506_ | new_C2505_;
  assign new_C2484_ = ~new_C2464_ & ~new_C2474_;
  assign new_C2483_ = new_C2464_ & new_C2474_;
  assign new_C2482_ = ~new_C2464_ | new_C2474_;
  assign new_C2481_ = new_C2448_ & ~new_C2449_;
  assign new_C2480_ = ~new_C2448_ & new_C2449_;
  assign new_C2479_ = new_C2501_ & ~new_C2502_;
  assign new_C2478_ = ~new_C2501_ & new_C2502_;
  assign new_C2477_ = ~new_C2500_ | ~new_C2499_;
  assign new_C2476_ = new_C2492_ | new_C2491_;
  assign new_C2475_ = new_C2498_ | new_C2497_;
  assign new_C2474_ = new_C2488_ | new_C2490_;
  assign new_C2473_ = ~new_C2495_ | ~new_C2496_;
  assign new_C2472_ = new_C2448_ & ~new_C2449_;
  assign new_C2471_ = new_C2462_ & ~new_C2474_;
  assign new_C2470_ = ~new_C2462_ & new_C2474_;
  assign new_C2469_ = ~new_C2460_ & new_C2486_;
  assign new_C2468_ = new_C2484_ | new_C2483_;
  assign new_C2467_ = new_C2481_ | new_C2480_;
  assign new_C2466_ = new_C2449_ | new_C2482_;
  assign new_C2465_ = new_C2474_ & new_C2477_;
  assign new_C2464_ = new_C2479_ | new_C2478_;
  assign new_C2463_ = new_C2474_ & new_C2473_;
  assign new_C2462_ = new_C2476_ & new_C2475_;
  assign new_C2461_ = new_C2471_ | new_C2470_;
  assign new_C2460_ = new_C2449_ | new_C2472_;
  assign C2459 = new_C2460_ | new_C2469_;
  assign C2458 = new_C2467_ & new_C2468_;
  assign C2457 = new_C2467_ & new_C2466_;
  assign C2456 = new_C2465_ | new_C2464_;
  assign C2455 = new_C2463_ | new_C2462_;
  assign C2454 = new_C2461_ & new_C2460_;
  assign new_C2453_ = new_D6932_;
  assign new_C2452_ = new_D6865_;
  assign new_C2451_ = new_D6798_;
  assign new_C2450_ = new_D6731_;
  assign new_C2449_ = new_D6664_;
  assign new_C2448_ = new_D6597_;
  assign new_C2447_ = ~new_C2386_ & new_C2400_;
  assign new_C2446_ = new_C2386_ & ~new_C2400_;
  assign new_C2445_ = new_C2386_ & ~new_C2400_;
  assign new_C2444_ = ~new_C2386_ & ~new_C2400_;
  assign new_C2443_ = new_C2386_ & new_C2400_;
  assign new_C2442_ = new_C2446_ | new_C2447_;
  assign new_C2441_ = ~new_C2386_ & new_C2400_;
  assign new_C2440_ = new_C2444_ | new_C2445_;
  assign new_C2439_ = ~new_C2415_ & ~new_C2435_;
  assign new_C2438_ = new_C2415_ & new_C2435_;
  assign new_C2437_ = ~new_C2382_ | ~new_C2407_;
  assign new_C2436_ = new_C2400_ & new_C2437_;
  assign new_C2435_ = new_C2383_ | new_C2384_;
  assign new_C2434_ = new_C2383_ | new_C2400_;
  assign new_C2433_ = ~new_C2400_ & ~new_C2436_;
  assign new_C2432_ = new_C2400_ | new_C2437_;
  assign new_C2431_ = new_C2383_ & ~new_C2384_;
  assign new_C2430_ = ~new_C2383_ & new_C2384_;
  assign new_C2429_ = new_C2393_ | new_C2426_;
  assign new_C2428_ = ~new_C2393_ & ~new_C2427_;
  assign new_C2427_ = new_C2393_ & new_C2426_;
  assign new_C2426_ = ~new_C2382_ | ~new_C2407_;
  assign new_C2425_ = ~new_C2383_ & new_C2393_;
  assign new_C2424_ = new_C2383_ & ~new_C2393_;
  assign new_C2423_ = new_C2385_ & new_C2422_;
  assign new_C2422_ = new_C2441_ | new_C2440_;
  assign new_C2421_ = ~new_C2385_ & new_C2420_;
  assign new_C2420_ = new_C2443_ | new_C2442_;
  assign new_C2419_ = new_C2385_ | new_C2418_;
  assign new_C2418_ = new_C2439_ | new_C2438_;
  assign new_C2417_ = ~new_C2397_ & ~new_C2407_;
  assign new_C2416_ = new_C2397_ & new_C2407_;
  assign new_C2415_ = ~new_C2397_ | new_C2407_;
  assign new_C2414_ = new_C2381_ & ~new_C2382_;
  assign new_C2413_ = ~new_C2381_ & new_C2382_;
  assign new_C2412_ = new_C2434_ & ~new_C2435_;
  assign new_C2411_ = ~new_C2434_ & new_C2435_;
  assign new_C2410_ = ~new_C2433_ | ~new_C2432_;
  assign new_C2409_ = new_C2425_ | new_C2424_;
  assign new_C2408_ = new_C2431_ | new_C2430_;
  assign new_C2407_ = new_C2421_ | new_C2423_;
  assign new_C2406_ = ~new_C2428_ | ~new_C2429_;
  assign new_C2405_ = new_C2381_ & ~new_C2382_;
  assign new_C2404_ = new_C2395_ & ~new_C2407_;
  assign new_C2403_ = ~new_C2395_ & new_C2407_;
  assign new_C2402_ = ~new_C2393_ & new_C2419_;
  assign new_C2401_ = new_C2417_ | new_C2416_;
  assign new_C2400_ = new_C2414_ | new_C2413_;
  assign new_C2399_ = new_C2382_ | new_C2415_;
  assign new_C2398_ = new_C2407_ & new_C2410_;
  assign new_C2397_ = new_C2412_ | new_C2411_;
  assign new_C2396_ = new_C2407_ & new_C2406_;
  assign new_C2395_ = new_C2409_ & new_C2408_;
  assign new_C2394_ = new_C2404_ | new_C2403_;
  assign new_C2393_ = new_C2382_ | new_C2405_;
  assign C2392 = new_C2393_ | new_C2402_;
  assign C2391 = new_C2400_ & new_C2401_;
  assign C2390 = new_C2400_ & new_C2399_;
  assign C2389 = new_C2398_ | new_C2397_;
  assign C2388 = new_C2396_ | new_C2395_;
  assign C2387 = new_C2394_ & new_C2393_;
  assign new_C2386_ = new_D6530_;
  assign new_C2385_ = new_D6463_;
  assign new_C2384_ = new_D6396_;
  assign new_C2383_ = new_D6329_;
  assign new_C2382_ = new_D6262_;
  assign new_C2381_ = new_D6195_;
  assign new_C2380_ = ~new_C2319_ & new_C2333_;
  assign new_C2379_ = new_C2319_ & ~new_C2333_;
  assign new_C2378_ = new_C2319_ & ~new_C2333_;
  assign new_C2377_ = ~new_C2319_ & ~new_C2333_;
  assign new_C2376_ = new_C2319_ & new_C2333_;
  assign new_C2375_ = new_C2379_ | new_C2380_;
  assign new_C2374_ = ~new_C2319_ & new_C2333_;
  assign new_C2373_ = new_C2377_ | new_C2378_;
  assign new_C2372_ = ~new_C2348_ & ~new_C2368_;
  assign new_C2371_ = new_C2348_ & new_C2368_;
  assign new_C2370_ = ~new_C2315_ | ~new_C2340_;
  assign new_C2369_ = new_C2333_ & new_C2370_;
  assign new_C2368_ = new_C2316_ | new_C2317_;
  assign new_C2367_ = new_C2316_ | new_C2333_;
  assign new_C2366_ = ~new_C2333_ & ~new_C2369_;
  assign new_C2365_ = new_C2333_ | new_C2370_;
  assign new_C2364_ = new_C2316_ & ~new_C2317_;
  assign new_C2363_ = ~new_C2316_ & new_C2317_;
  assign new_C2362_ = new_C2326_ | new_C2359_;
  assign new_C2361_ = ~new_C2326_ & ~new_C2360_;
  assign new_C2360_ = new_C2326_ & new_C2359_;
  assign new_C2359_ = ~new_C2315_ | ~new_C2340_;
  assign new_C2358_ = ~new_C2316_ & new_C2326_;
  assign new_C2357_ = new_C2316_ & ~new_C2326_;
  assign new_C2356_ = new_C2318_ & new_C2355_;
  assign new_C2355_ = new_C2374_ | new_C2373_;
  assign new_C2354_ = ~new_C2318_ & new_C2353_;
  assign new_C2353_ = new_C2376_ | new_C2375_;
  assign new_C2352_ = new_C2318_ | new_C2351_;
  assign new_C2351_ = new_C2372_ | new_C2371_;
  assign new_C2350_ = ~new_C2330_ & ~new_C2340_;
  assign new_C2349_ = new_C2330_ & new_C2340_;
  assign new_C2348_ = ~new_C2330_ | new_C2340_;
  assign new_C2347_ = new_C2314_ & ~new_C2315_;
  assign new_C2346_ = ~new_C2314_ & new_C2315_;
  assign new_C2345_ = new_C2367_ & ~new_C2368_;
  assign new_C2344_ = ~new_C2367_ & new_C2368_;
  assign new_C2343_ = ~new_C2366_ | ~new_C2365_;
  assign new_C2342_ = new_C2358_ | new_C2357_;
  assign new_C2341_ = new_C2364_ | new_C2363_;
  assign new_C2340_ = new_C2354_ | new_C2356_;
  assign new_C2339_ = ~new_C2361_ | ~new_C2362_;
  assign new_C2338_ = new_C2314_ & ~new_C2315_;
  assign new_C2337_ = new_C2328_ & ~new_C2340_;
  assign new_C2336_ = ~new_C2328_ & new_C2340_;
  assign new_C2335_ = ~new_C2326_ & new_C2352_;
  assign new_C2334_ = new_C2350_ | new_C2349_;
  assign new_C2333_ = new_C2347_ | new_C2346_;
  assign new_C2332_ = new_C2315_ | new_C2348_;
  assign new_C2331_ = new_C2340_ & new_C2343_;
  assign new_C2330_ = new_C2345_ | new_C2344_;
  assign new_C2329_ = new_C2340_ & new_C2339_;
  assign new_C2328_ = new_C2342_ & new_C2341_;
  assign new_C2327_ = new_C2337_ | new_C2336_;
  assign new_C2326_ = new_C2315_ | new_C2338_;
  assign C2325 = new_C2326_ | new_C2335_;
  assign C2324 = new_C2333_ & new_C2334_;
  assign C2323 = new_C2333_ & new_C2332_;
  assign C2322 = new_C2331_ | new_C2330_;
  assign C2321 = new_C2329_ | new_C2328_;
  assign C2320 = new_C2327_ & new_C2326_;
  assign new_C2319_ = new_D6128_;
  assign new_C2318_ = new_D6061_;
  assign new_C2317_ = new_D5994_;
  assign new_C2316_ = new_D5927_;
  assign new_C2315_ = new_D5860_;
  assign new_C2314_ = new_D5793_;
  assign new_C2313_ = ~new_C2252_ & new_C2266_;
  assign new_C2312_ = new_C2252_ & ~new_C2266_;
  assign new_C2311_ = new_C2252_ & ~new_C2266_;
  assign new_C2310_ = ~new_C2252_ & ~new_C2266_;
  assign new_C2309_ = new_C2252_ & new_C2266_;
  assign new_C2308_ = new_C2312_ | new_C2313_;
  assign new_C2307_ = ~new_C2252_ & new_C2266_;
  assign new_C2306_ = new_C2310_ | new_C2311_;
  assign new_C2305_ = ~new_C2281_ & ~new_C2301_;
  assign new_C2304_ = new_C2281_ & new_C2301_;
  assign new_C2303_ = ~new_C2248_ | ~new_C2273_;
  assign new_C2302_ = new_C2266_ & new_C2303_;
  assign new_C2301_ = new_C2249_ | new_C2250_;
  assign new_C2300_ = new_C2249_ | new_C2266_;
  assign new_C2299_ = ~new_C2266_ & ~new_C2302_;
  assign new_C2298_ = new_C2266_ | new_C2303_;
  assign new_C2297_ = new_C2249_ & ~new_C2250_;
  assign new_C2296_ = ~new_C2249_ & new_C2250_;
  assign new_C2295_ = new_C2259_ | new_C2292_;
  assign new_C2294_ = ~new_C2259_ & ~new_C2293_;
  assign new_C2293_ = new_C2259_ & new_C2292_;
  assign new_C2292_ = ~new_C2248_ | ~new_C2273_;
  assign new_C2291_ = ~new_C2249_ & new_C2259_;
  assign new_C2290_ = new_C2249_ & ~new_C2259_;
  assign new_C2289_ = new_C2251_ & new_C2288_;
  assign new_C2288_ = new_C2307_ | new_C2306_;
  assign new_C2287_ = ~new_C2251_ & new_C2286_;
  assign new_C2286_ = new_C2309_ | new_C2308_;
  assign new_C2285_ = new_C2251_ | new_C2284_;
  assign new_C2284_ = new_C2305_ | new_C2304_;
  assign new_C2283_ = ~new_C2263_ & ~new_C2273_;
  assign new_C2282_ = new_C2263_ & new_C2273_;
  assign new_C2281_ = ~new_C2263_ | new_C2273_;
  assign new_C2280_ = new_C2247_ & ~new_C2248_;
  assign new_C2279_ = ~new_C2247_ & new_C2248_;
  assign new_C2278_ = new_C2300_ & ~new_C2301_;
  assign new_C2277_ = ~new_C2300_ & new_C2301_;
  assign new_C2276_ = ~new_C2299_ | ~new_C2298_;
  assign new_C2275_ = new_C2291_ | new_C2290_;
  assign new_C2274_ = new_C2297_ | new_C2296_;
  assign new_C2273_ = new_C2287_ | new_C2289_;
  assign new_C2272_ = ~new_C2294_ | ~new_C2295_;
  assign new_C2271_ = new_C2247_ & ~new_C2248_;
  assign new_C2270_ = new_C2261_ & ~new_C2273_;
  assign new_C2269_ = ~new_C2261_ & new_C2273_;
  assign new_C2268_ = ~new_C2259_ & new_C2285_;
  assign new_C2267_ = new_C2283_ | new_C2282_;
  assign new_C2266_ = new_C2280_ | new_C2279_;
  assign new_C2265_ = new_C2248_ | new_C2281_;
  assign new_C2264_ = new_C2273_ & new_C2276_;
  assign new_C2263_ = new_C2278_ | new_C2277_;
  assign new_C2262_ = new_C2273_ & new_C2272_;
  assign new_C2261_ = new_C2275_ & new_C2274_;
  assign new_C2260_ = new_C2270_ | new_C2269_;
  assign new_C2259_ = new_C2248_ | new_C2271_;
  assign C2258 = new_C2259_ | new_C2268_;
  assign C2257 = new_C2266_ & new_C2267_;
  assign C2256 = new_C2266_ & new_C2265_;
  assign C2255 = new_C2264_ | new_C2263_;
  assign C2254 = new_C2262_ | new_C2261_;
  assign C2253 = new_C2260_ & new_C2259_;
  assign new_C2252_ = new_D5726_;
  assign new_C2251_ = new_D5659_;
  assign new_C2250_ = new_D5592_;
  assign new_C2249_ = new_D5525_;
  assign new_C2248_ = new_D5458_;
  assign new_C2247_ = new_D5391_;
  assign new_C2246_ = ~new_C2185_ & new_C2199_;
  assign new_C2245_ = new_C2185_ & ~new_C2199_;
  assign new_C2244_ = new_C2185_ & ~new_C2199_;
  assign new_C2243_ = ~new_C2185_ & ~new_C2199_;
  assign new_C2242_ = new_C2185_ & new_C2199_;
  assign new_C2241_ = new_C2245_ | new_C2246_;
  assign new_C2240_ = ~new_C2185_ & new_C2199_;
  assign new_C2239_ = new_C2243_ | new_C2244_;
  assign new_C2238_ = ~new_C2214_ & ~new_C2234_;
  assign new_C2237_ = new_C2214_ & new_C2234_;
  assign new_C2236_ = ~new_C2181_ | ~new_C2206_;
  assign new_C2235_ = new_C2199_ & new_C2236_;
  assign new_C2234_ = new_C2182_ | new_C2183_;
  assign new_C2233_ = new_C2182_ | new_C2199_;
  assign new_C2232_ = ~new_C2199_ & ~new_C2235_;
  assign new_C2231_ = new_C2199_ | new_C2236_;
  assign new_C2230_ = new_C2182_ & ~new_C2183_;
  assign new_C2229_ = ~new_C2182_ & new_C2183_;
  assign new_C2228_ = new_C2192_ | new_C2225_;
  assign new_C2227_ = ~new_C2192_ & ~new_C2226_;
  assign new_C2226_ = new_C2192_ & new_C2225_;
  assign new_C2225_ = ~new_C2181_ | ~new_C2206_;
  assign new_C2224_ = ~new_C2182_ & new_C2192_;
  assign new_C2223_ = new_C2182_ & ~new_C2192_;
  assign new_C2222_ = new_C2184_ & new_C2221_;
  assign new_C2221_ = new_C2240_ | new_C2239_;
  assign new_C2220_ = ~new_C2184_ & new_C2219_;
  assign new_C2219_ = new_C2242_ | new_C2241_;
  assign new_C2218_ = new_C2184_ | new_C2217_;
  assign new_C2217_ = new_C2238_ | new_C2237_;
  assign new_C2216_ = ~new_C2196_ & ~new_C2206_;
  assign new_C2215_ = new_C2196_ & new_C2206_;
  assign new_C2214_ = ~new_C2196_ | new_C2206_;
  assign new_C2213_ = new_C2180_ & ~new_C2181_;
  assign new_C2212_ = ~new_C2180_ & new_C2181_;
  assign new_C2211_ = new_C2233_ & ~new_C2234_;
  assign new_C2210_ = ~new_C2233_ & new_C2234_;
  assign new_C2209_ = ~new_C2232_ | ~new_C2231_;
  assign new_C2208_ = new_C2224_ | new_C2223_;
  assign new_C2207_ = new_C2230_ | new_C2229_;
  assign new_C2206_ = new_C2220_ | new_C2222_;
  assign new_C2205_ = ~new_C2227_ | ~new_C2228_;
  assign new_C2204_ = new_C2180_ & ~new_C2181_;
  assign new_C2203_ = new_C2194_ & ~new_C2206_;
  assign new_C2202_ = ~new_C2194_ & new_C2206_;
  assign new_C2201_ = ~new_C2192_ & new_C2218_;
  assign new_C2200_ = new_C2216_ | new_C2215_;
  assign new_C2199_ = new_C2213_ | new_C2212_;
  assign new_C2198_ = new_C2181_ | new_C2214_;
  assign new_C2197_ = new_C2206_ & new_C2209_;
  assign new_C2196_ = new_C2211_ | new_C2210_;
  assign new_C2195_ = new_C2206_ & new_C2205_;
  assign new_C2194_ = new_C2208_ & new_C2207_;
  assign new_C2193_ = new_C2203_ | new_C2202_;
  assign new_C2192_ = new_C2181_ | new_C2204_;
  assign C2191 = new_C2192_ | new_C2201_;
  assign C2190 = new_C2199_ & new_C2200_;
  assign C2189 = new_C2199_ & new_C2198_;
  assign C2188 = new_C2197_ | new_C2196_;
  assign C2187 = new_C2195_ | new_C2194_;
  assign C2186 = new_C2193_ & new_C2192_;
  assign new_C2185_ = new_D5324_;
  assign new_C2184_ = new_D5257_;
  assign new_C2183_ = new_D5190_;
  assign new_C2182_ = new_D5123_;
  assign new_C2181_ = new_D5056_;
  assign new_C2180_ = new_D4989_;
  assign new_C2179_ = ~new_C2118_ & new_C2132_;
  assign new_C2178_ = new_C2118_ & ~new_C2132_;
  assign new_C2177_ = new_C2118_ & ~new_C2132_;
  assign new_C2176_ = ~new_C2118_ & ~new_C2132_;
  assign new_C2175_ = new_C2118_ & new_C2132_;
  assign new_C2174_ = new_C2178_ | new_C2179_;
  assign new_C2173_ = ~new_C2118_ & new_C2132_;
  assign new_C2172_ = new_C2176_ | new_C2177_;
  assign new_C2171_ = ~new_C2147_ & ~new_C2167_;
  assign new_C2170_ = new_C2147_ & new_C2167_;
  assign new_C2169_ = ~new_C2114_ | ~new_C2139_;
  assign new_C2168_ = new_C2132_ & new_C2169_;
  assign new_C2167_ = new_C2115_ | new_C2116_;
  assign new_C2166_ = new_C2115_ | new_C2132_;
  assign new_C2165_ = ~new_C2132_ & ~new_C2168_;
  assign new_C2164_ = new_C2132_ | new_C2169_;
  assign new_C2163_ = new_C2115_ & ~new_C2116_;
  assign new_C2162_ = ~new_C2115_ & new_C2116_;
  assign new_C2161_ = new_C2125_ | new_C2158_;
  assign new_C2160_ = ~new_C2125_ & ~new_C2159_;
  assign new_C2159_ = new_C2125_ & new_C2158_;
  assign new_C2158_ = ~new_C2114_ | ~new_C2139_;
  assign new_C2157_ = ~new_C2115_ & new_C2125_;
  assign new_C2156_ = new_C2115_ & ~new_C2125_;
  assign new_C2155_ = new_C2117_ & new_C2154_;
  assign new_C2154_ = new_C2173_ | new_C2172_;
  assign new_C2153_ = ~new_C2117_ & new_C2152_;
  assign new_C2152_ = new_C2175_ | new_C2174_;
  assign new_C2151_ = new_C2117_ | new_C2150_;
  assign new_C2150_ = new_C2171_ | new_C2170_;
  assign new_C2149_ = ~new_C2129_ & ~new_C2139_;
  assign new_C2148_ = new_C2129_ & new_C2139_;
  assign new_C2147_ = ~new_C2129_ | new_C2139_;
  assign new_C2146_ = new_C2113_ & ~new_C2114_;
  assign new_C2145_ = ~new_C2113_ & new_C2114_;
  assign new_C2144_ = new_C2166_ & ~new_C2167_;
  assign new_C2143_ = ~new_C2166_ & new_C2167_;
  assign new_C2142_ = ~new_C2165_ | ~new_C2164_;
  assign new_C2141_ = new_C2157_ | new_C2156_;
  assign new_C2140_ = new_C2163_ | new_C2162_;
  assign new_C2139_ = new_C2153_ | new_C2155_;
  assign new_C2138_ = ~new_C2160_ | ~new_C2161_;
  assign new_C2137_ = new_C2113_ & ~new_C2114_;
  assign new_C2136_ = new_C2127_ & ~new_C2139_;
  assign new_C2135_ = ~new_C2127_ & new_C2139_;
  assign new_C2134_ = ~new_C2125_ & new_C2151_;
  assign new_C2133_ = new_C2149_ | new_C2148_;
  assign new_C2132_ = new_C2146_ | new_C2145_;
  assign new_C2131_ = new_C2114_ | new_C2147_;
  assign new_C2130_ = new_C2139_ & new_C2142_;
  assign new_C2129_ = new_C2144_ | new_C2143_;
  assign new_C2128_ = new_C2139_ & new_C2138_;
  assign new_C2127_ = new_C2141_ & new_C2140_;
  assign new_C2126_ = new_C2136_ | new_C2135_;
  assign new_C2125_ = new_C2114_ | new_C2137_;
  assign C2124 = new_C2125_ | new_C2134_;
  assign C2123 = new_C2132_ & new_C2133_;
  assign C2122 = new_C2132_ & new_C2131_;
  assign C2121 = new_C2130_ | new_C2129_;
  assign C2120 = new_C2128_ | new_C2127_;
  assign C2119 = new_C2126_ & new_C2125_;
  assign new_C2118_ = new_D4922_;
  assign new_C2117_ = new_D4855_;
  assign new_C2116_ = new_D4788_;
  assign new_C2115_ = new_D4721_;
  assign new_C2114_ = new_D4654_;
  assign new_C2113_ = new_D4587_;
  assign new_C2112_ = ~new_C2051_ & new_C2065_;
  assign new_C2111_ = new_C2051_ & ~new_C2065_;
  assign new_C2110_ = new_C2051_ & ~new_C2065_;
  assign new_C2109_ = ~new_C2051_ & ~new_C2065_;
  assign new_C2108_ = new_C2051_ & new_C2065_;
  assign new_C2107_ = new_C2111_ | new_C2112_;
  assign new_C2106_ = ~new_C2051_ & new_C2065_;
  assign new_C2105_ = new_C2109_ | new_C2110_;
  assign new_C2104_ = ~new_C2080_ & ~new_C2100_;
  assign new_C2103_ = new_C2080_ & new_C2100_;
  assign new_C2102_ = ~new_C2047_ | ~new_C2072_;
  assign new_C2101_ = new_C2065_ & new_C2102_;
  assign new_C2100_ = new_C2048_ | new_C2049_;
  assign new_C2099_ = new_C2048_ | new_C2065_;
  assign new_C2098_ = ~new_C2065_ & ~new_C2101_;
  assign new_C2097_ = new_C2065_ | new_C2102_;
  assign new_C2096_ = new_C2048_ & ~new_C2049_;
  assign new_C2095_ = ~new_C2048_ & new_C2049_;
  assign new_C2094_ = new_C2058_ | new_C2091_;
  assign new_C2093_ = ~new_C2058_ & ~new_C2092_;
  assign new_C2092_ = new_C2058_ & new_C2091_;
  assign new_C2091_ = ~new_C2047_ | ~new_C2072_;
  assign new_C2090_ = ~new_C2048_ & new_C2058_;
  assign new_C2089_ = new_C2048_ & ~new_C2058_;
  assign new_C2088_ = new_C2050_ & new_C2087_;
  assign new_C2087_ = new_C2106_ | new_C2105_;
  assign new_C2086_ = ~new_C2050_ & new_C2085_;
  assign new_C2085_ = new_C2108_ | new_C2107_;
  assign new_C2084_ = new_C2050_ | new_C2083_;
  assign new_C2083_ = new_C2104_ | new_C2103_;
  assign new_C2082_ = ~new_C2062_ & ~new_C2072_;
  assign new_C2081_ = new_C2062_ & new_C2072_;
  assign new_C2080_ = ~new_C2062_ | new_C2072_;
  assign new_C2079_ = new_C2046_ & ~new_C2047_;
  assign new_C2078_ = ~new_C2046_ & new_C2047_;
  assign new_C2077_ = new_C2099_ & ~new_C2100_;
  assign new_C2076_ = ~new_C2099_ & new_C2100_;
  assign new_C2075_ = ~new_C2098_ | ~new_C2097_;
  assign new_C2074_ = new_C2090_ | new_C2089_;
  assign new_C2073_ = new_C2096_ | new_C2095_;
  assign new_C2072_ = new_C2086_ | new_C2088_;
  assign new_C2071_ = ~new_C2093_ | ~new_C2094_;
  assign new_C2070_ = new_C2046_ & ~new_C2047_;
  assign new_C2069_ = new_C2060_ & ~new_C2072_;
  assign new_C2068_ = ~new_C2060_ & new_C2072_;
  assign new_C2067_ = ~new_C2058_ & new_C2084_;
  assign new_C2066_ = new_C2082_ | new_C2081_;
  assign new_C2065_ = new_C2079_ | new_C2078_;
  assign new_C2064_ = new_C2047_ | new_C2080_;
  assign new_C2063_ = new_C2072_ & new_C2075_;
  assign new_C2062_ = new_C2077_ | new_C2076_;
  assign new_C2061_ = new_C2072_ & new_C2071_;
  assign new_C2060_ = new_C2074_ & new_C2073_;
  assign new_C2059_ = new_C2069_ | new_C2068_;
  assign new_C2058_ = new_C2047_ | new_C2070_;
  assign C2057 = new_C2058_ | new_C2067_;
  assign C2056 = new_C2065_ & new_C2066_;
  assign C2055 = new_C2065_ & new_C2064_;
  assign C2054 = new_C2063_ | new_C2062_;
  assign C2053 = new_C2061_ | new_C2060_;
  assign C2052 = new_C2059_ & new_C2058_;
  assign new_C2051_ = new_D4520_;
  assign new_C2050_ = new_D4453_;
  assign new_C2049_ = new_D4386_;
  assign new_C2048_ = new_D4319_;
  assign new_C2047_ = new_D4252_;
  assign new_C2046_ = new_D4185_;
  assign new_C2045_ = ~new_C1984_ & new_C1998_;
  assign new_C2044_ = new_C1984_ & ~new_C1998_;
  assign new_C2043_ = new_C1984_ & ~new_C1998_;
  assign new_C2042_ = ~new_C1984_ & ~new_C1998_;
  assign new_C2041_ = new_C1984_ & new_C1998_;
  assign new_C2040_ = new_C2044_ | new_C2045_;
  assign new_C2039_ = ~new_C1984_ & new_C1998_;
  assign new_C2038_ = new_C2042_ | new_C2043_;
  assign new_C2037_ = ~new_C2013_ & ~new_C2033_;
  assign new_C2036_ = new_C2013_ & new_C2033_;
  assign new_C2035_ = ~new_C1980_ | ~new_C2005_;
  assign new_C2034_ = new_C1998_ & new_C2035_;
  assign new_C2033_ = new_C1981_ | new_C1982_;
  assign new_C2032_ = new_C1981_ | new_C1998_;
  assign new_C2031_ = ~new_C1998_ & ~new_C2034_;
  assign new_C2030_ = new_C1998_ | new_C2035_;
  assign new_C2029_ = new_C1981_ & ~new_C1982_;
  assign new_C2028_ = ~new_C1981_ & new_C1982_;
  assign new_C2027_ = new_C1991_ | new_C2024_;
  assign new_C2026_ = ~new_C1991_ & ~new_C2025_;
  assign new_C2025_ = new_C1991_ & new_C2024_;
  assign new_C2024_ = ~new_C1980_ | ~new_C2005_;
  assign new_C2023_ = ~new_C1981_ & new_C1991_;
  assign new_C2022_ = new_C1981_ & ~new_C1991_;
  assign new_C2021_ = new_C1983_ & new_C2020_;
  assign new_C2020_ = new_C2039_ | new_C2038_;
  assign new_C2019_ = ~new_C1983_ & new_C2018_;
  assign new_C2018_ = new_C2041_ | new_C2040_;
  assign new_C2017_ = new_C1983_ | new_C2016_;
  assign new_C2016_ = new_C2037_ | new_C2036_;
  assign new_C2015_ = ~new_C1995_ & ~new_C2005_;
  assign new_C2014_ = new_C1995_ & new_C2005_;
  assign new_C2013_ = ~new_C1995_ | new_C2005_;
  assign new_C2012_ = new_C1979_ & ~new_C1980_;
  assign new_C2011_ = ~new_C1979_ & new_C1980_;
  assign new_C2010_ = new_C2032_ & ~new_C2033_;
  assign new_C2009_ = ~new_C2032_ & new_C2033_;
  assign new_C2008_ = ~new_C2031_ | ~new_C2030_;
  assign new_C2007_ = new_C2023_ | new_C2022_;
  assign new_C2006_ = new_C2029_ | new_C2028_;
  assign new_C2005_ = new_C2019_ | new_C2021_;
  assign new_C2004_ = ~new_C2026_ | ~new_C2027_;
  assign new_C2003_ = new_C1979_ & ~new_C1980_;
  assign new_C2002_ = new_C1993_ & ~new_C2005_;
  assign new_C2001_ = ~new_C1993_ & new_C2005_;
  assign new_C2000_ = ~new_C1991_ & new_C2017_;
  assign new_C1999_ = new_C2015_ | new_C2014_;
  assign new_C1998_ = new_C2012_ | new_C2011_;
  assign new_C1997_ = new_C1980_ | new_C2013_;
  assign new_C1996_ = new_C2005_ & new_C2008_;
  assign new_C1995_ = new_C2010_ | new_C2009_;
  assign new_C1994_ = new_C2005_ & new_C2004_;
  assign new_C1993_ = new_C2007_ & new_C2006_;
  assign new_C1992_ = new_C2002_ | new_C2001_;
  assign new_C1991_ = new_C1980_ | new_C2003_;
  assign C1990 = new_C1991_ | new_C2000_;
  assign C1989 = new_C1998_ & new_C1999_;
  assign C1988 = new_C1998_ & new_C1997_;
  assign C1987 = new_C1996_ | new_C1995_;
  assign C1986 = new_C1994_ | new_C1993_;
  assign C1985 = new_C1992_ & new_C1991_;
  assign new_C1984_ = new_D4118_;
  assign new_C1983_ = new_D4051_;
  assign new_C1982_ = new_D3984_;
  assign new_C1981_ = new_D3917_;
  assign new_C1980_ = new_D3850_;
  assign new_C1979_ = new_D3783_;
  assign new_C1978_ = ~new_C1917_ & new_C1931_;
  assign new_C1977_ = new_C1917_ & ~new_C1931_;
  assign new_C1976_ = new_C1917_ & ~new_C1931_;
  assign new_C1975_ = ~new_C1917_ & ~new_C1931_;
  assign new_C1974_ = new_C1917_ & new_C1931_;
  assign new_C1973_ = new_C1977_ | new_C1978_;
  assign new_C1972_ = ~new_C1917_ & new_C1931_;
  assign new_C1971_ = new_C1975_ | new_C1976_;
  assign new_C1970_ = ~new_C1946_ & ~new_C1966_;
  assign new_C1969_ = new_C1946_ & new_C1966_;
  assign new_C1968_ = ~new_C1913_ | ~new_C1938_;
  assign new_C1967_ = new_C1931_ & new_C1968_;
  assign new_C1966_ = new_C1914_ | new_C1915_;
  assign new_C1965_ = new_C1914_ | new_C1931_;
  assign new_C1964_ = ~new_C1931_ & ~new_C1967_;
  assign new_C1963_ = new_C1931_ | new_C1968_;
  assign new_C1962_ = new_C1914_ & ~new_C1915_;
  assign new_C1961_ = ~new_C1914_ & new_C1915_;
  assign new_C1960_ = new_C1924_ | new_C1957_;
  assign new_C1959_ = ~new_C1924_ & ~new_C1958_;
  assign new_C1958_ = new_C1924_ & new_C1957_;
  assign new_C1957_ = ~new_C1913_ | ~new_C1938_;
  assign new_C1956_ = ~new_C1914_ & new_C1924_;
  assign new_C1955_ = new_C1914_ & ~new_C1924_;
  assign new_C1954_ = new_C1916_ & new_C1953_;
  assign new_C1953_ = new_C1972_ | new_C1971_;
  assign new_C1952_ = ~new_C1916_ & new_C1951_;
  assign new_C1951_ = new_C1974_ | new_C1973_;
  assign new_C1950_ = new_C1916_ | new_C1949_;
  assign new_C1949_ = new_C1970_ | new_C1969_;
  assign new_C1948_ = ~new_C1928_ & ~new_C1938_;
  assign new_C1947_ = new_C1928_ & new_C1938_;
  assign new_C1946_ = ~new_C1928_ | new_C1938_;
  assign new_C1945_ = new_C1912_ & ~new_C1913_;
  assign new_C1944_ = ~new_C1912_ & new_C1913_;
  assign new_C1943_ = new_C1965_ & ~new_C1966_;
  assign new_C1942_ = ~new_C1965_ & new_C1966_;
  assign new_C1941_ = ~new_C1964_ | ~new_C1963_;
  assign new_C1940_ = new_C1956_ | new_C1955_;
  assign new_C1939_ = new_C1962_ | new_C1961_;
  assign new_C1938_ = new_C1952_ | new_C1954_;
  assign new_C1937_ = ~new_C1959_ | ~new_C1960_;
  assign new_C1936_ = new_C1912_ & ~new_C1913_;
  assign new_C1935_ = new_C1926_ & ~new_C1938_;
  assign new_C1934_ = ~new_C1926_ & new_C1938_;
  assign new_C1933_ = ~new_C1924_ & new_C1950_;
  assign new_C1932_ = new_C1948_ | new_C1947_;
  assign new_C1931_ = new_C1945_ | new_C1944_;
  assign new_C1930_ = new_C1913_ | new_C1946_;
  assign new_C1929_ = new_C1938_ & new_C1941_;
  assign new_C1928_ = new_C1943_ | new_C1942_;
  assign new_C1927_ = new_C1938_ & new_C1937_;
  assign new_C1926_ = new_C1940_ & new_C1939_;
  assign new_C1925_ = new_C1935_ | new_C1934_;
  assign new_C1924_ = new_C1913_ | new_C1936_;
  assign C1923 = new_C1924_ | new_C1933_;
  assign C1922 = new_C1931_ & new_C1932_;
  assign C1921 = new_C1931_ & new_C1930_;
  assign C1920 = new_C1929_ | new_C1928_;
  assign C1919 = new_C1927_ | new_C1926_;
  assign C1918 = new_C1925_ & new_C1924_;
  assign new_C1917_ = new_D3716_;
  assign new_C1916_ = new_D3649_;
  assign new_C1915_ = new_D3582_;
  assign new_C1914_ = new_D3515_;
  assign new_C1913_ = new_D3448_;
  assign new_C1912_ = new_D3381_;
  assign new_C1911_ = ~new_C1850_ & new_C1864_;
  assign new_C1910_ = new_C1850_ & ~new_C1864_;
  assign new_C1909_ = new_C1850_ & ~new_C1864_;
  assign new_C1908_ = ~new_C1850_ & ~new_C1864_;
  assign new_C1907_ = new_C1850_ & new_C1864_;
  assign new_C1906_ = new_C1910_ | new_C1911_;
  assign new_C1905_ = ~new_C1850_ & new_C1864_;
  assign new_C1904_ = new_C1908_ | new_C1909_;
  assign new_C1903_ = ~new_C1879_ & ~new_C1899_;
  assign new_C1902_ = new_C1879_ & new_C1899_;
  assign new_C1901_ = ~new_C1846_ | ~new_C1871_;
  assign new_C1900_ = new_C1864_ & new_C1901_;
  assign new_C1899_ = new_C1847_ | new_C1848_;
  assign new_C1898_ = new_C1847_ | new_C1864_;
  assign new_C1897_ = ~new_C1864_ & ~new_C1900_;
  assign new_C1896_ = new_C1864_ | new_C1901_;
  assign new_C1895_ = new_C1847_ & ~new_C1848_;
  assign new_C1894_ = ~new_C1847_ & new_C1848_;
  assign new_C1893_ = new_C1857_ | new_C1890_;
  assign new_C1892_ = ~new_C1857_ & ~new_C1891_;
  assign new_C1891_ = new_C1857_ & new_C1890_;
  assign new_C1890_ = ~new_C1846_ | ~new_C1871_;
  assign new_C1889_ = ~new_C1847_ & new_C1857_;
  assign new_C1888_ = new_C1847_ & ~new_C1857_;
  assign new_C1887_ = new_C1849_ & new_C1886_;
  assign new_C1886_ = new_C1905_ | new_C1904_;
  assign new_C1885_ = ~new_C1849_ & new_C1884_;
  assign new_C1884_ = new_C1907_ | new_C1906_;
  assign new_C1883_ = new_C1849_ | new_C1882_;
  assign new_C1882_ = new_C1903_ | new_C1902_;
  assign new_C1881_ = ~new_C1861_ & ~new_C1871_;
  assign new_C1880_ = new_C1861_ & new_C1871_;
  assign new_C1879_ = ~new_C1861_ | new_C1871_;
  assign new_C1878_ = new_C1845_ & ~new_C1846_;
  assign new_C1877_ = ~new_C1845_ & new_C1846_;
  assign new_C1876_ = new_C1898_ & ~new_C1899_;
  assign new_C1875_ = ~new_C1898_ & new_C1899_;
  assign new_C1874_ = ~new_C1897_ | ~new_C1896_;
  assign new_C1873_ = new_C1889_ | new_C1888_;
  assign new_C1872_ = new_C1895_ | new_C1894_;
  assign new_C1871_ = new_C1885_ | new_C1887_;
  assign new_C1870_ = ~new_C1892_ | ~new_C1893_;
  assign new_C1869_ = new_C1845_ & ~new_C1846_;
  assign new_C1868_ = new_C1859_ & ~new_C1871_;
  assign new_C1867_ = ~new_C1859_ & new_C1871_;
  assign new_C1866_ = ~new_C1857_ & new_C1883_;
  assign new_C1865_ = new_C1881_ | new_C1880_;
  assign new_C1864_ = new_C1878_ | new_C1877_;
  assign new_C1863_ = new_C1846_ | new_C1879_;
  assign new_C1862_ = new_C1871_ & new_C1874_;
  assign new_C1861_ = new_C1876_ | new_C1875_;
  assign new_C1860_ = new_C1871_ & new_C1870_;
  assign new_C1859_ = new_C1873_ & new_C1872_;
  assign new_C1858_ = new_C1868_ | new_C1867_;
  assign new_C1857_ = new_C1846_ | new_C1869_;
  assign C1856 = new_C1857_ | new_C1866_;
  assign C1855 = new_C1864_ & new_C1865_;
  assign C1854 = new_C1864_ & new_C1863_;
  assign C1853 = new_C1862_ | new_C1861_;
  assign C1852 = new_C1860_ | new_C1859_;
  assign C1851 = new_C1858_ & new_C1857_;
  assign new_C1850_ = new_D3314_;
  assign new_C1849_ = new_D3247_;
  assign new_C1848_ = new_D3180_;
  assign new_C1847_ = new_D3113_;
  assign new_C1846_ = new_D3046_;
  assign new_C1845_ = new_D2979_;
  assign new_C1844_ = ~new_C1783_ & new_C1797_;
  assign new_C1843_ = new_C1783_ & ~new_C1797_;
  assign new_C1842_ = new_C1783_ & ~new_C1797_;
  assign new_C1841_ = ~new_C1783_ & ~new_C1797_;
  assign new_C1840_ = new_C1783_ & new_C1797_;
  assign new_C1839_ = new_C1843_ | new_C1844_;
  assign new_C1838_ = ~new_C1783_ & new_C1797_;
  assign new_C1837_ = new_C1841_ | new_C1842_;
  assign new_C1836_ = ~new_C1812_ & ~new_C1832_;
  assign new_C1835_ = new_C1812_ & new_C1832_;
  assign new_C1834_ = ~new_C1779_ | ~new_C1804_;
  assign new_C1833_ = new_C1797_ & new_C1834_;
  assign new_C1832_ = new_C1780_ | new_C1781_;
  assign new_C1831_ = new_C1780_ | new_C1797_;
  assign new_C1830_ = ~new_C1797_ & ~new_C1833_;
  assign new_C1829_ = new_C1797_ | new_C1834_;
  assign new_C1828_ = new_C1780_ & ~new_C1781_;
  assign new_C1827_ = ~new_C1780_ & new_C1781_;
  assign new_C1826_ = new_C1790_ | new_C1823_;
  assign new_C1825_ = ~new_C1790_ & ~new_C1824_;
  assign new_C1824_ = new_C1790_ & new_C1823_;
  assign new_C1823_ = ~new_C1779_ | ~new_C1804_;
  assign new_C1822_ = ~new_C1780_ & new_C1790_;
  assign new_C1821_ = new_C1780_ & ~new_C1790_;
  assign new_C1820_ = new_C1782_ & new_C1819_;
  assign new_C1819_ = new_C1838_ | new_C1837_;
  assign new_C1818_ = ~new_C1782_ & new_C1817_;
  assign new_C1817_ = new_C1840_ | new_C1839_;
  assign new_C1816_ = new_C1782_ | new_C1815_;
  assign new_C1815_ = new_C1836_ | new_C1835_;
  assign new_C1814_ = ~new_C1794_ & ~new_C1804_;
  assign new_C1813_ = new_C1794_ & new_C1804_;
  assign new_C1812_ = ~new_C1794_ | new_C1804_;
  assign new_C1811_ = new_C1778_ & ~new_C1779_;
  assign new_C1810_ = ~new_C1778_ & new_C1779_;
  assign new_C1809_ = new_C1831_ & ~new_C1832_;
  assign new_C1808_ = ~new_C1831_ & new_C1832_;
  assign new_C1807_ = ~new_C1830_ | ~new_C1829_;
  assign new_C1806_ = new_C1822_ | new_C1821_;
  assign new_C1805_ = new_C1828_ | new_C1827_;
  assign new_C1804_ = new_C1818_ | new_C1820_;
  assign new_C1803_ = ~new_C1825_ | ~new_C1826_;
  assign new_C1802_ = new_C1778_ & ~new_C1779_;
  assign new_C1801_ = new_C1792_ & ~new_C1804_;
  assign new_C1800_ = ~new_C1792_ & new_C1804_;
  assign new_C1799_ = ~new_C1790_ & new_C1816_;
  assign new_C1798_ = new_C1814_ | new_C1813_;
  assign new_C1797_ = new_C1811_ | new_C1810_;
  assign new_C1796_ = new_C1779_ | new_C1812_;
  assign new_C1795_ = new_C1804_ & new_C1807_;
  assign new_C1794_ = new_C1809_ | new_C1808_;
  assign new_C1793_ = new_C1804_ & new_C1803_;
  assign new_C1792_ = new_C1806_ & new_C1805_;
  assign new_C1791_ = new_C1801_ | new_C1800_;
  assign new_C1790_ = new_C1779_ | new_C1802_;
  assign C1789 = new_C1790_ | new_C1799_;
  assign C1788 = new_C1797_ & new_C1798_;
  assign C1787 = new_C1797_ & new_C1796_;
  assign C1786 = new_C1795_ | new_C1794_;
  assign C1785 = new_C1793_ | new_C1792_;
  assign C1784 = new_C1791_ & new_C1790_;
  assign new_C1783_ = new_D2912_;
  assign new_C1782_ = new_D2845_;
  assign new_C1781_ = new_D2778_;
  assign new_C1780_ = new_D2711_;
  assign new_C1779_ = new_D2644_;
  assign new_C1778_ = new_D2577_;
  assign new_C1777_ = ~new_C1716_ & new_C1730_;
  assign new_C1776_ = new_C1716_ & ~new_C1730_;
  assign new_C1775_ = new_C1716_ & ~new_C1730_;
  assign new_C1774_ = ~new_C1716_ & ~new_C1730_;
  assign new_C1773_ = new_C1716_ & new_C1730_;
  assign new_C1772_ = new_C1776_ | new_C1777_;
  assign new_C1771_ = ~new_C1716_ & new_C1730_;
  assign new_C1770_ = new_C1774_ | new_C1775_;
  assign new_C1769_ = ~new_C1745_ & ~new_C1765_;
  assign new_C1768_ = new_C1745_ & new_C1765_;
  assign new_C1767_ = ~new_C1712_ | ~new_C1737_;
  assign new_C1766_ = new_C1730_ & new_C1767_;
  assign new_C1765_ = new_C1713_ | new_C1714_;
  assign new_C1764_ = new_C1713_ | new_C1730_;
  assign new_C1763_ = ~new_C1730_ & ~new_C1766_;
  assign new_C1762_ = new_C1730_ | new_C1767_;
  assign new_C1761_ = new_C1713_ & ~new_C1714_;
  assign new_C1760_ = ~new_C1713_ & new_C1714_;
  assign new_C1759_ = new_C1723_ | new_C1756_;
  assign new_C1758_ = ~new_C1723_ & ~new_C1757_;
  assign new_C1757_ = new_C1723_ & new_C1756_;
  assign new_C1756_ = ~new_C1712_ | ~new_C1737_;
  assign new_C1755_ = ~new_C1713_ & new_C1723_;
  assign new_C1754_ = new_C1713_ & ~new_C1723_;
  assign new_C1753_ = new_C1715_ & new_C1752_;
  assign new_C1752_ = new_C1771_ | new_C1770_;
  assign new_C1751_ = ~new_C1715_ & new_C1750_;
  assign new_C1750_ = new_C1773_ | new_C1772_;
  assign new_C1749_ = new_C1715_ | new_C1748_;
  assign new_C1748_ = new_C1769_ | new_C1768_;
  assign new_C1747_ = ~new_C1727_ & ~new_C1737_;
  assign new_C1746_ = new_C1727_ & new_C1737_;
  assign new_C1745_ = ~new_C1727_ | new_C1737_;
  assign new_C1744_ = new_C1711_ & ~new_C1712_;
  assign new_C1743_ = ~new_C1711_ & new_C1712_;
  assign new_C1742_ = new_C1764_ & ~new_C1765_;
  assign new_C1741_ = ~new_C1764_ & new_C1765_;
  assign new_C1740_ = ~new_C1763_ | ~new_C1762_;
  assign new_C1739_ = new_C1755_ | new_C1754_;
  assign new_C1738_ = new_C1761_ | new_C1760_;
  assign new_C1737_ = new_C1751_ | new_C1753_;
  assign new_C1736_ = ~new_C1758_ | ~new_C1759_;
  assign new_C1735_ = new_C1711_ & ~new_C1712_;
  assign new_C1734_ = new_C1725_ & ~new_C1737_;
  assign new_C1733_ = ~new_C1725_ & new_C1737_;
  assign new_C1732_ = ~new_C1723_ & new_C1749_;
  assign new_C1731_ = new_C1747_ | new_C1746_;
  assign new_C1730_ = new_C1744_ | new_C1743_;
  assign new_C1729_ = new_C1712_ | new_C1745_;
  assign new_C1728_ = new_C1737_ & new_C1740_;
  assign new_C1727_ = new_C1742_ | new_C1741_;
  assign new_C1726_ = new_C1737_ & new_C1736_;
  assign new_C1725_ = new_C1739_ & new_C1738_;
  assign new_C1724_ = new_C1734_ | new_C1733_;
  assign new_C1723_ = new_C1712_ | new_C1735_;
  assign C1722 = new_C1723_ | new_C1732_;
  assign C1721 = new_C1730_ & new_C1731_;
  assign C1720 = new_C1730_ & new_C1729_;
  assign C1719 = new_C1728_ | new_C1727_;
  assign C1718 = new_C1726_ | new_C1725_;
  assign C1717 = new_C1724_ & new_C1723_;
  assign new_C1716_ = new_D2510_;
  assign new_C1715_ = new_D2443_;
  assign new_C1714_ = new_D2376_;
  assign new_C1713_ = new_D2309_;
  assign new_C1712_ = new_D2242_;
  assign new_C1711_ = new_D2175_;
  assign new_C1710_ = ~new_C1649_ & new_C1663_;
  assign new_C1709_ = new_C1649_ & ~new_C1663_;
  assign new_C1708_ = new_C1649_ & ~new_C1663_;
  assign new_C1707_ = ~new_C1649_ & ~new_C1663_;
  assign new_C1706_ = new_C1649_ & new_C1663_;
  assign new_C1705_ = new_C1709_ | new_C1710_;
  assign new_C1704_ = ~new_C1649_ & new_C1663_;
  assign new_C1703_ = new_C1707_ | new_C1708_;
  assign new_C1702_ = ~new_C1678_ & ~new_C1698_;
  assign new_C1701_ = new_C1678_ & new_C1698_;
  assign new_C1700_ = ~new_C1645_ | ~new_C1670_;
  assign new_C1699_ = new_C1663_ & new_C1700_;
  assign new_C1698_ = new_C1646_ | new_C1647_;
  assign new_C1697_ = new_C1646_ | new_C1663_;
  assign new_C1696_ = ~new_C1663_ & ~new_C1699_;
  assign new_C1695_ = new_C1663_ | new_C1700_;
  assign new_C1694_ = new_C1646_ & ~new_C1647_;
  assign new_C1693_ = ~new_C1646_ & new_C1647_;
  assign new_C1692_ = new_C1656_ | new_C1689_;
  assign new_C1691_ = ~new_C1656_ & ~new_C1690_;
  assign new_C1690_ = new_C1656_ & new_C1689_;
  assign new_C1689_ = ~new_C1645_ | ~new_C1670_;
  assign new_C1688_ = ~new_C1646_ & new_C1656_;
  assign new_C1687_ = new_C1646_ & ~new_C1656_;
  assign new_C1686_ = new_C1648_ & new_C1685_;
  assign new_C1685_ = new_C1704_ | new_C1703_;
  assign new_C1684_ = ~new_C1648_ & new_C1683_;
  assign new_C1683_ = new_C1706_ | new_C1705_;
  assign new_C1682_ = new_C1648_ | new_C1681_;
  assign new_C1681_ = new_C1702_ | new_C1701_;
  assign new_C1680_ = ~new_C1660_ & ~new_C1670_;
  assign new_C1679_ = new_C1660_ & new_C1670_;
  assign new_C1678_ = ~new_C1660_ | new_C1670_;
  assign new_C1677_ = new_C1644_ & ~new_C1645_;
  assign new_C1676_ = ~new_C1644_ & new_C1645_;
  assign new_C1675_ = new_C1697_ & ~new_C1698_;
  assign new_C1674_ = ~new_C1697_ & new_C1698_;
  assign new_C1673_ = ~new_C1696_ | ~new_C1695_;
  assign new_C1672_ = new_C1688_ | new_C1687_;
  assign new_C1671_ = new_C1694_ | new_C1693_;
  assign new_C1670_ = new_C1684_ | new_C1686_;
  assign new_C1669_ = ~new_C1691_ | ~new_C1692_;
  assign new_C1668_ = new_C1644_ & ~new_C1645_;
  assign new_C1667_ = new_C1658_ & ~new_C1670_;
  assign new_C1666_ = ~new_C1658_ & new_C1670_;
  assign new_C1665_ = ~new_C1656_ & new_C1682_;
  assign new_C1664_ = new_C1680_ | new_C1679_;
  assign new_C1663_ = new_C1677_ | new_C1676_;
  assign new_C1662_ = new_C1645_ | new_C1678_;
  assign new_C1661_ = new_C1670_ & new_C1673_;
  assign new_C1660_ = new_C1675_ | new_C1674_;
  assign new_C1659_ = new_C1670_ & new_C1669_;
  assign new_C1658_ = new_C1672_ & new_C1671_;
  assign new_C1657_ = new_C1667_ | new_C1666_;
  assign new_C1656_ = new_C1645_ | new_C1668_;
  assign C1655 = new_C1656_ | new_C1665_;
  assign C1654 = new_C1663_ & new_C1664_;
  assign C1653 = new_C1663_ & new_C1662_;
  assign C1652 = new_C1661_ | new_C1660_;
  assign C1651 = new_C1659_ | new_C1658_;
  assign C1650 = new_C1657_ & new_C1656_;
  assign new_C1649_ = new_D2108_;
  assign new_C1648_ = new_D2041_;
  assign new_C1647_ = new_D1974_;
  assign new_C1646_ = new_D1907_;
  assign new_C1645_ = new_D1840_;
  assign new_C1644_ = new_D1773_;
  assign new_C1643_ = ~new_C1582_ & new_C1596_;
  assign new_C1642_ = new_C1582_ & ~new_C1596_;
  assign new_C1641_ = new_C1582_ & ~new_C1596_;
  assign new_C1640_ = ~new_C1582_ & ~new_C1596_;
  assign new_C1639_ = new_C1582_ & new_C1596_;
  assign new_C1638_ = new_C1642_ | new_C1643_;
  assign new_C1637_ = ~new_C1582_ & new_C1596_;
  assign new_C1636_ = new_C1640_ | new_C1641_;
  assign new_C1635_ = ~new_C1611_ & ~new_C1631_;
  assign new_C1634_ = new_C1611_ & new_C1631_;
  assign new_C1633_ = ~new_C1578_ | ~new_C1603_;
  assign new_C1632_ = new_C1596_ & new_C1633_;
  assign new_C1631_ = new_C1579_ | new_C1580_;
  assign new_C1630_ = new_C1579_ | new_C1596_;
  assign new_C1629_ = ~new_C1596_ & ~new_C1632_;
  assign new_C1628_ = new_C1596_ | new_C1633_;
  assign new_C1627_ = new_C1579_ & ~new_C1580_;
  assign new_C1626_ = ~new_C1579_ & new_C1580_;
  assign new_C1625_ = new_C1589_ | new_C1622_;
  assign new_C1624_ = ~new_C1589_ & ~new_C1623_;
  assign new_C1623_ = new_C1589_ & new_C1622_;
  assign new_C1622_ = ~new_C1578_ | ~new_C1603_;
  assign new_C1621_ = ~new_C1579_ & new_C1589_;
  assign new_C1620_ = new_C1579_ & ~new_C1589_;
  assign new_C1619_ = new_C1581_ & new_C1618_;
  assign new_C1618_ = new_C1637_ | new_C1636_;
  assign new_C1617_ = ~new_C1581_ & new_C1616_;
  assign new_C1616_ = new_C1639_ | new_C1638_;
  assign new_C1615_ = new_C1581_ | new_C1614_;
  assign new_C1614_ = new_C1635_ | new_C1634_;
  assign new_C1613_ = ~new_C1593_ & ~new_C1603_;
  assign new_C1612_ = new_C1593_ & new_C1603_;
  assign new_C1611_ = ~new_C1593_ | new_C1603_;
  assign new_C1610_ = new_C1577_ & ~new_C1578_;
  assign new_C1609_ = ~new_C1577_ & new_C1578_;
  assign new_C1608_ = new_C1630_ & ~new_C1631_;
  assign new_C1607_ = ~new_C1630_ & new_C1631_;
  assign new_C1606_ = ~new_C1629_ | ~new_C1628_;
  assign new_C1605_ = new_C1621_ | new_C1620_;
  assign new_C1604_ = new_C1627_ | new_C1626_;
  assign new_C1603_ = new_C1617_ | new_C1619_;
  assign new_C1602_ = ~new_C1624_ | ~new_C1625_;
  assign new_C1601_ = new_C1577_ & ~new_C1578_;
  assign new_C1600_ = new_C1591_ & ~new_C1603_;
  assign new_C1599_ = ~new_C1591_ & new_C1603_;
  assign new_C1598_ = ~new_C1589_ & new_C1615_;
  assign new_C1597_ = new_C1613_ | new_C1612_;
  assign new_C1596_ = new_C1610_ | new_C1609_;
  assign new_C1595_ = new_C1578_ | new_C1611_;
  assign new_C1594_ = new_C1603_ & new_C1606_;
  assign new_C1593_ = new_C1608_ | new_C1607_;
  assign new_C1592_ = new_C1603_ & new_C1602_;
  assign new_C1591_ = new_C1605_ & new_C1604_;
  assign new_C1590_ = new_C1600_ | new_C1599_;
  assign new_C1589_ = new_C1578_ | new_C1601_;
  assign C1588 = new_C1589_ | new_C1598_;
  assign C1587 = new_C1596_ & new_C1597_;
  assign C1586 = new_C1596_ & new_C1595_;
  assign C1585 = new_C1594_ | new_C1593_;
  assign C1584 = new_C1592_ | new_C1591_;
  assign C1583 = new_C1590_ & new_C1589_;
  assign new_C1582_ = new_D1706_;
  assign new_C1581_ = new_D1639_;
  assign new_C1580_ = new_D1572_;
  assign new_C1579_ = new_D1505_;
  assign new_C1578_ = new_D1438_;
  assign new_C1577_ = new_D1371_;
  assign new_C1576_ = ~new_C1515_ & new_C1529_;
  assign new_C1575_ = new_C1515_ & ~new_C1529_;
  assign new_C1574_ = new_C1515_ & ~new_C1529_;
  assign new_C1573_ = ~new_C1515_ & ~new_C1529_;
  assign new_C1572_ = new_C1515_ & new_C1529_;
  assign new_C1571_ = new_C1575_ | new_C1576_;
  assign new_C1570_ = ~new_C1515_ & new_C1529_;
  assign new_C1569_ = new_C1573_ | new_C1574_;
  assign new_C1568_ = ~new_C1544_ & ~new_C1564_;
  assign new_C1567_ = new_C1544_ & new_C1564_;
  assign new_C1566_ = ~new_C1511_ | ~new_C1536_;
  assign new_C1565_ = new_C1529_ & new_C1566_;
  assign new_C1564_ = new_C1512_ | new_C1513_;
  assign new_C1563_ = new_C1512_ | new_C1529_;
  assign new_C1562_ = ~new_C1529_ & ~new_C1565_;
  assign new_C1561_ = new_C1529_ | new_C1566_;
  assign new_C1560_ = new_C1512_ & ~new_C1513_;
  assign new_C1559_ = ~new_C1512_ & new_C1513_;
  assign new_C1558_ = new_C1522_ | new_C1555_;
  assign new_C1557_ = ~new_C1522_ & ~new_C1556_;
  assign new_C1556_ = new_C1522_ & new_C1555_;
  assign new_C1555_ = ~new_C1511_ | ~new_C1536_;
  assign new_C1554_ = ~new_C1512_ & new_C1522_;
  assign new_C1553_ = new_C1512_ & ~new_C1522_;
  assign new_C1552_ = new_C1514_ & new_C1551_;
  assign new_C1551_ = new_C1570_ | new_C1569_;
  assign new_C1550_ = ~new_C1514_ & new_C1549_;
  assign new_C1549_ = new_C1572_ | new_C1571_;
  assign new_C1548_ = new_C1514_ | new_C1547_;
  assign new_C1547_ = new_C1568_ | new_C1567_;
  assign new_C1546_ = ~new_C1526_ & ~new_C1536_;
  assign new_C1545_ = new_C1526_ & new_C1536_;
  assign new_C1544_ = ~new_C1526_ | new_C1536_;
  assign new_C1543_ = new_C1510_ & ~new_C1511_;
  assign new_C1542_ = ~new_C1510_ & new_C1511_;
  assign new_C1541_ = new_C1563_ & ~new_C1564_;
  assign new_C1540_ = ~new_C1563_ & new_C1564_;
  assign new_C1539_ = ~new_C1562_ | ~new_C1561_;
  assign new_C1538_ = new_C1554_ | new_C1553_;
  assign new_C1537_ = new_C1560_ | new_C1559_;
  assign new_C1536_ = new_C1550_ | new_C1552_;
  assign new_C1535_ = ~new_C1557_ | ~new_C1558_;
  assign new_C1534_ = new_C1510_ & ~new_C1511_;
  assign new_C1533_ = new_C1524_ & ~new_C1536_;
  assign new_C1532_ = ~new_C1524_ & new_C1536_;
  assign new_C1531_ = ~new_C1522_ & new_C1548_;
  assign new_C1530_ = new_C1546_ | new_C1545_;
  assign new_C1529_ = new_C1543_ | new_C1542_;
  assign new_C1528_ = new_C1511_ | new_C1544_;
  assign new_C1527_ = new_C1536_ & new_C1539_;
  assign new_C1526_ = new_C1541_ | new_C1540_;
  assign new_C1525_ = new_C1536_ & new_C1535_;
  assign new_C1524_ = new_C1538_ & new_C1537_;
  assign new_C1523_ = new_C1533_ | new_C1532_;
  assign new_C1522_ = new_C1511_ | new_C1534_;
  assign C1521 = new_C1522_ | new_C1531_;
  assign C1520 = new_C1529_ & new_C1530_;
  assign C1519 = new_C1529_ & new_C1528_;
  assign C1518 = new_C1527_ | new_C1526_;
  assign C1517 = new_C1525_ | new_C1524_;
  assign C1516 = new_C1523_ & new_C1522_;
  assign new_C1515_ = new_D1304_;
  assign new_C1514_ = new_D1237_;
  assign new_C1513_ = new_D1170_;
  assign new_C1512_ = new_D1103_;
  assign new_C1511_ = new_D1036_;
  assign new_C1510_ = new_D969_;
  assign new_C1509_ = ~new_C1448_ & new_C1462_;
  assign new_C1508_ = new_C1448_ & ~new_C1462_;
  assign new_C1507_ = new_C1448_ & ~new_C1462_;
  assign new_C1506_ = ~new_C1448_ & ~new_C1462_;
  assign new_C1505_ = new_C1448_ & new_C1462_;
  assign new_C1504_ = new_C1508_ | new_C1509_;
  assign new_C1503_ = ~new_C1448_ & new_C1462_;
  assign new_C1502_ = new_C1506_ | new_C1507_;
  assign new_C1501_ = ~new_C1477_ & ~new_C1497_;
  assign new_C1500_ = new_C1477_ & new_C1497_;
  assign new_C1499_ = ~new_C1444_ | ~new_C1469_;
  assign new_C1498_ = new_C1462_ & new_C1499_;
  assign new_C1497_ = new_C1445_ | new_C1446_;
  assign new_C1496_ = new_C1445_ | new_C1462_;
  assign new_C1495_ = ~new_C1462_ & ~new_C1498_;
  assign new_C1494_ = new_C1462_ | new_C1499_;
  assign new_C1493_ = new_C1445_ & ~new_C1446_;
  assign new_C1492_ = ~new_C1445_ & new_C1446_;
  assign new_C1491_ = new_C1455_ | new_C1488_;
  assign new_C1490_ = ~new_C1455_ & ~new_C1489_;
  assign new_C1489_ = new_C1455_ & new_C1488_;
  assign new_C1488_ = ~new_C1444_ | ~new_C1469_;
  assign new_C1487_ = ~new_C1445_ & new_C1455_;
  assign new_C1486_ = new_C1445_ & ~new_C1455_;
  assign new_C1485_ = new_C1447_ & new_C1484_;
  assign new_C1484_ = new_C1503_ | new_C1502_;
  assign new_C1483_ = ~new_C1447_ & new_C1482_;
  assign new_C1482_ = new_C1505_ | new_C1504_;
  assign new_C1481_ = new_C1447_ | new_C1480_;
  assign new_C1480_ = new_C1501_ | new_C1500_;
  assign new_C1479_ = ~new_C1459_ & ~new_C1469_;
  assign new_C1478_ = new_C1459_ & new_C1469_;
  assign new_C1477_ = ~new_C1459_ | new_C1469_;
  assign new_C1476_ = new_C1443_ & ~new_C1444_;
  assign new_C1475_ = ~new_C1443_ & new_C1444_;
  assign new_C1474_ = new_C1496_ & ~new_C1497_;
  assign new_C1473_ = ~new_C1496_ & new_C1497_;
  assign new_C1472_ = ~new_C1495_ | ~new_C1494_;
  assign new_C1471_ = new_C1487_ | new_C1486_;
  assign new_C1470_ = new_C1493_ | new_C1492_;
  assign new_C1469_ = new_C1483_ | new_C1485_;
  assign new_C1468_ = ~new_C1490_ | ~new_C1491_;
  assign new_C1467_ = new_C1443_ & ~new_C1444_;
  assign new_C1466_ = new_C1457_ & ~new_C1469_;
  assign new_C1465_ = ~new_C1457_ & new_C1469_;
  assign new_C1464_ = ~new_C1455_ & new_C1481_;
  assign new_C1463_ = new_C1479_ | new_C1478_;
  assign new_C1462_ = new_C1476_ | new_C1475_;
  assign new_C1461_ = new_C1444_ | new_C1477_;
  assign new_C1460_ = new_C1469_ & new_C1472_;
  assign new_C1459_ = new_C1474_ | new_C1473_;
  assign new_C1458_ = new_C1469_ & new_C1468_;
  assign new_C1457_ = new_C1471_ & new_C1470_;
  assign new_C1456_ = new_C1466_ | new_C1465_;
  assign new_C1455_ = new_C1444_ | new_C1467_;
  assign C1454 = new_C1455_ | new_C1464_;
  assign C1453 = new_C1462_ & new_C1463_;
  assign C1452 = new_C1462_ & new_C1461_;
  assign C1451 = new_C1460_ | new_C1459_;
  assign C1450 = new_C1458_ | new_C1457_;
  assign C1449 = new_C1456_ & new_C1455_;
  assign new_C1448_ = new_D902_;
  assign new_C1447_ = new_D835_;
  assign new_C1446_ = new_D768_;
  assign new_C1445_ = new_D701_;
  assign new_C1444_ = new_D634_;
  assign new_C1443_ = new_D567_;
  assign new_C1442_ = ~new_C1381_ & new_C1395_;
  assign new_C1441_ = new_C1381_ & ~new_C1395_;
  assign new_C1440_ = new_C1381_ & ~new_C1395_;
  assign new_C1439_ = ~new_C1381_ & ~new_C1395_;
  assign new_C1438_ = new_C1381_ & new_C1395_;
  assign new_C1437_ = new_C1441_ | new_C1442_;
  assign new_C1436_ = ~new_C1381_ & new_C1395_;
  assign new_C1435_ = new_C1439_ | new_C1440_;
  assign new_C1434_ = ~new_C1410_ & ~new_C1430_;
  assign new_C1433_ = new_C1410_ & new_C1430_;
  assign new_C1432_ = ~new_C1377_ | ~new_C1402_;
  assign new_C1431_ = new_C1395_ & new_C1432_;
  assign new_C1430_ = new_C1378_ | new_C1379_;
  assign new_C1429_ = new_C1378_ | new_C1395_;
  assign new_C1428_ = ~new_C1395_ & ~new_C1431_;
  assign new_C1427_ = new_C1395_ | new_C1432_;
  assign new_C1426_ = new_C1378_ & ~new_C1379_;
  assign new_C1425_ = ~new_C1378_ & new_C1379_;
  assign new_C1424_ = new_C1388_ | new_C1421_;
  assign new_C1423_ = ~new_C1388_ & ~new_C1422_;
  assign new_C1422_ = new_C1388_ & new_C1421_;
  assign new_C1421_ = ~new_C1377_ | ~new_C1402_;
  assign new_C1420_ = ~new_C1378_ & new_C1388_;
  assign new_C1419_ = new_C1378_ & ~new_C1388_;
  assign new_C1418_ = new_C1380_ & new_C1417_;
  assign new_C1417_ = new_C1436_ | new_C1435_;
  assign new_C1416_ = ~new_C1380_ & new_C1415_;
  assign new_C1415_ = new_C1438_ | new_C1437_;
  assign new_C1414_ = new_C1380_ | new_C1413_;
  assign new_C1413_ = new_C1434_ | new_C1433_;
  assign new_C1412_ = ~new_C1392_ & ~new_C1402_;
  assign new_C1411_ = new_C1392_ & new_C1402_;
  assign new_C1410_ = ~new_C1392_ | new_C1402_;
  assign new_C1409_ = new_C1376_ & ~new_C1377_;
  assign new_C1408_ = ~new_C1376_ & new_C1377_;
  assign new_C1407_ = new_C1429_ & ~new_C1430_;
  assign new_C1406_ = ~new_C1429_ & new_C1430_;
  assign new_C1405_ = ~new_C1428_ | ~new_C1427_;
  assign new_C1404_ = new_C1420_ | new_C1419_;
  assign new_C1403_ = new_C1426_ | new_C1425_;
  assign new_C1402_ = new_C1416_ | new_C1418_;
  assign new_C1401_ = ~new_C1423_ | ~new_C1424_;
  assign new_C1400_ = new_C1376_ & ~new_C1377_;
  assign new_C1399_ = new_C1390_ & ~new_C1402_;
  assign new_C1398_ = ~new_C1390_ & new_C1402_;
  assign new_C1397_ = ~new_C1388_ & new_C1414_;
  assign new_C1396_ = new_C1412_ | new_C1411_;
  assign new_C1395_ = new_C1409_ | new_C1408_;
  assign new_C1394_ = new_C1377_ | new_C1410_;
  assign new_C1393_ = new_C1402_ & new_C1405_;
  assign new_C1392_ = new_C1407_ | new_C1406_;
  assign new_C1391_ = new_C1402_ & new_C1401_;
  assign new_C1390_ = new_C1404_ & new_C1403_;
  assign new_C1389_ = new_C1399_ | new_C1398_;
  assign new_C1388_ = new_C1377_ | new_C1400_;
  assign C1387 = new_C1388_ | new_C1397_;
  assign C1386 = new_C1395_ & new_C1396_;
  assign C1385 = new_C1395_ & new_C1394_;
  assign C1384 = new_C1393_ | new_C1392_;
  assign C1383 = new_C1391_ | new_C1390_;
  assign C1382 = new_C1389_ & new_C1388_;
  assign new_C1381_ = new_D500_;
  assign new_C1380_ = new_D433_;
  assign new_C1379_ = new_D366_;
  assign new_C1378_ = new_D299_;
  assign new_C1377_ = new_D232_;
  assign new_C1376_ = new_D165_;
  assign new_C1375_ = ~new_C1314_ & new_C1328_;
  assign new_C1374_ = new_C1314_ & ~new_C1328_;
  assign new_C1373_ = new_C1314_ & ~new_C1328_;
  assign new_C1372_ = ~new_C1314_ & ~new_C1328_;
  assign new_C1371_ = new_C1314_ & new_C1328_;
  assign new_C1370_ = new_C1374_ | new_C1375_;
  assign new_C1369_ = ~new_C1314_ & new_C1328_;
  assign new_C1368_ = new_C1372_ | new_C1373_;
  assign new_C1367_ = ~new_C1343_ & ~new_C1363_;
  assign new_C1366_ = new_C1343_ & new_C1363_;
  assign new_C1365_ = ~new_C1310_ | ~new_C1335_;
  assign new_C1364_ = new_C1328_ & new_C1365_;
  assign new_C1363_ = new_C1311_ | new_C1312_;
  assign new_C1362_ = new_C1311_ | new_C1328_;
  assign new_C1361_ = ~new_C1328_ & ~new_C1364_;
  assign new_C1360_ = new_C1328_ | new_C1365_;
  assign new_C1359_ = new_C1311_ & ~new_C1312_;
  assign new_C1358_ = ~new_C1311_ & new_C1312_;
  assign new_C1357_ = new_C1321_ | new_C1354_;
  assign new_C1356_ = ~new_C1321_ & ~new_C1355_;
  assign new_C1355_ = new_C1321_ & new_C1354_;
  assign new_C1354_ = ~new_C1310_ | ~new_C1335_;
  assign new_C1353_ = ~new_C1311_ & new_C1321_;
  assign new_C1352_ = new_C1311_ & ~new_C1321_;
  assign new_C1351_ = new_C1313_ & new_C1350_;
  assign new_C1350_ = new_C1369_ | new_C1368_;
  assign new_C1349_ = ~new_C1313_ & new_C1348_;
  assign new_C1348_ = new_C1371_ | new_C1370_;
  assign new_C1347_ = new_C1313_ | new_C1346_;
  assign new_C1346_ = new_C1367_ | new_C1366_;
  assign new_C1345_ = ~new_C1325_ & ~new_C1335_;
  assign new_C1344_ = new_C1325_ & new_C1335_;
  assign new_C1343_ = ~new_C1325_ | new_C1335_;
  assign new_C1342_ = new_C1309_ & ~new_C1310_;
  assign new_C1341_ = ~new_C1309_ & new_C1310_;
  assign new_C1340_ = new_C1362_ & ~new_C1363_;
  assign new_C1339_ = ~new_C1362_ & new_C1363_;
  assign new_C1338_ = ~new_C1361_ | ~new_C1360_;
  assign new_C1337_ = new_C1353_ | new_C1352_;
  assign new_C1336_ = new_C1359_ | new_C1358_;
  assign new_C1335_ = new_C1349_ | new_C1351_;
  assign new_C1334_ = ~new_C1356_ | ~new_C1357_;
  assign new_C1333_ = new_C1309_ & ~new_C1310_;
  assign new_C1332_ = new_C1323_ & ~new_C1335_;
  assign new_C1331_ = ~new_C1323_ & new_C1335_;
  assign new_C1330_ = ~new_C1321_ & new_C1347_;
  assign new_C1329_ = new_C1345_ | new_C1344_;
  assign new_C1328_ = new_C1342_ | new_C1341_;
  assign new_C1327_ = new_C1310_ | new_C1343_;
  assign new_C1326_ = new_C1335_ & new_C1338_;
  assign new_C1325_ = new_C1340_ | new_C1339_;
  assign new_C1324_ = new_C1335_ & new_C1334_;
  assign new_C1323_ = new_C1337_ & new_C1336_;
  assign new_C1322_ = new_C1332_ | new_C1331_;
  assign new_C1321_ = new_C1310_ | new_C1333_;
  assign C1320 = new_C1321_ | new_C1330_;
  assign C1319 = new_C1328_ & new_C1329_;
  assign C1318 = new_C1328_ & new_C1327_;
  assign C1317 = new_C1326_ | new_C1325_;
  assign C1316 = new_C1324_ | new_C1323_;
  assign C1315 = new_C1322_ & new_C1321_;
  assign new_C1314_ = new_D98_;
  assign new_C1313_ = new_D31_;
  assign new_C1312_ = new_C9963_;
  assign new_C1311_ = new_C9896_;
  assign new_C1310_ = new_C9829_;
  assign new_C1309_ = new_C9762_;
  assign new_C1308_ = ~new_C1247_ & new_C1261_;
  assign new_C1307_ = new_C1247_ & ~new_C1261_;
  assign new_C1306_ = new_C1247_ & ~new_C1261_;
  assign new_C1305_ = ~new_C1247_ & ~new_C1261_;
  assign new_C1304_ = new_C1247_ & new_C1261_;
  assign new_C1303_ = new_C1307_ | new_C1308_;
  assign new_C1302_ = ~new_C1247_ & new_C1261_;
  assign new_C1301_ = new_C1305_ | new_C1306_;
  assign new_C1300_ = ~new_C1276_ & ~new_C1296_;
  assign new_C1299_ = new_C1276_ & new_C1296_;
  assign new_C1298_ = ~new_C1243_ | ~new_C1268_;
  assign new_C1297_ = new_C1261_ & new_C1298_;
  assign new_C1296_ = new_C1244_ | new_C1245_;
  assign new_C1295_ = new_C1244_ | new_C1261_;
  assign new_C1294_ = ~new_C1261_ & ~new_C1297_;
  assign new_C1293_ = new_C1261_ | new_C1298_;
  assign new_C1292_ = new_C1244_ & ~new_C1245_;
  assign new_C1291_ = ~new_C1244_ & new_C1245_;
  assign new_C1290_ = new_C1254_ | new_C1287_;
  assign new_C1289_ = ~new_C1254_ & ~new_C1288_;
  assign new_C1288_ = new_C1254_ & new_C1287_;
  assign new_C1287_ = ~new_C1243_ | ~new_C1268_;
  assign new_C1286_ = ~new_C1244_ & new_C1254_;
  assign new_C1285_ = new_C1244_ & ~new_C1254_;
  assign new_C1284_ = new_C1246_ & new_C1283_;
  assign new_C1283_ = new_C1302_ | new_C1301_;
  assign new_C1282_ = ~new_C1246_ & new_C1281_;
  assign new_C1281_ = new_C1304_ | new_C1303_;
  assign new_C1280_ = new_C1246_ | new_C1279_;
  assign new_C1279_ = new_C1300_ | new_C1299_;
  assign new_C1278_ = ~new_C1258_ & ~new_C1268_;
  assign new_C1277_ = new_C1258_ & new_C1268_;
  assign new_C1276_ = ~new_C1258_ | new_C1268_;
  assign new_C1275_ = new_C1242_ & ~new_C1243_;
  assign new_C1274_ = ~new_C1242_ & new_C1243_;
  assign new_C1273_ = new_C1295_ & ~new_C1296_;
  assign new_C1272_ = ~new_C1295_ & new_C1296_;
  assign new_C1271_ = ~new_C1294_ | ~new_C1293_;
  assign new_C1270_ = new_C1286_ | new_C1285_;
  assign new_C1269_ = new_C1292_ | new_C1291_;
  assign new_C1268_ = new_C1282_ | new_C1284_;
  assign new_C1267_ = ~new_C1289_ | ~new_C1290_;
  assign new_C1266_ = new_C1242_ & ~new_C1243_;
  assign new_C1265_ = new_C1256_ & ~new_C1268_;
  assign new_C1264_ = ~new_C1256_ & new_C1268_;
  assign new_C1263_ = ~new_C1254_ & new_C1280_;
  assign new_C1262_ = new_C1278_ | new_C1277_;
  assign new_C1261_ = new_C1275_ | new_C1274_;
  assign new_C1260_ = new_C1243_ | new_C1276_;
  assign new_C1259_ = new_C1268_ & new_C1271_;
  assign new_C1258_ = new_C1273_ | new_C1272_;
  assign new_C1257_ = new_C1268_ & new_C1267_;
  assign new_C1256_ = new_C1270_ & new_C1269_;
  assign new_C1255_ = new_C1265_ | new_C1264_;
  assign new_C1254_ = new_C1243_ | new_C1266_;
  assign C1253 = new_C1254_ | new_C1263_;
  assign C1252 = new_C1261_ & new_C1262_;
  assign C1251 = new_C1261_ & new_C1260_;
  assign C1250 = new_C1259_ | new_C1258_;
  assign C1249 = new_C1257_ | new_C1256_;
  assign C1248 = new_C1255_ & new_C1254_;
  assign new_C1247_ = new_C9695_;
  assign new_C1246_ = new_C9628_;
  assign new_C1245_ = new_C9561_;
  assign new_C1244_ = new_C9494_;
  assign new_C1243_ = new_C9427_;
  assign new_C1242_ = new_C9360_;
  assign new_C1241_ = ~new_C1180_ & new_C1194_;
  assign new_C1240_ = new_C1180_ & ~new_C1194_;
  assign new_C1239_ = new_C1180_ & ~new_C1194_;
  assign new_C1238_ = ~new_C1180_ & ~new_C1194_;
  assign new_C1237_ = new_C1180_ & new_C1194_;
  assign new_C1236_ = new_C1240_ | new_C1241_;
  assign new_C1235_ = ~new_C1180_ & new_C1194_;
  assign new_C1234_ = new_C1238_ | new_C1239_;
  assign new_C1233_ = ~new_C1209_ & ~new_C1229_;
  assign new_C1232_ = new_C1209_ & new_C1229_;
  assign new_C1231_ = ~new_C1176_ | ~new_C1201_;
  assign new_C1230_ = new_C1194_ & new_C1231_;
  assign new_C1229_ = new_C1177_ | new_C1178_;
  assign new_C1228_ = new_C1177_ | new_C1194_;
  assign new_C1227_ = ~new_C1194_ & ~new_C1230_;
  assign new_C1226_ = new_C1194_ | new_C1231_;
  assign new_C1225_ = new_C1177_ & ~new_C1178_;
  assign new_C1224_ = ~new_C1177_ & new_C1178_;
  assign new_C1223_ = new_C1187_ | new_C1220_;
  assign new_C1222_ = ~new_C1187_ & ~new_C1221_;
  assign new_C1221_ = new_C1187_ & new_C1220_;
  assign new_C1220_ = ~new_C1176_ | ~new_C1201_;
  assign new_C1219_ = ~new_C1177_ & new_C1187_;
  assign new_C1218_ = new_C1177_ & ~new_C1187_;
  assign new_C1217_ = new_C1179_ & new_C1216_;
  assign new_C1216_ = new_C1235_ | new_C1234_;
  assign new_C1215_ = ~new_C1179_ & new_C1214_;
  assign new_C1214_ = new_C1237_ | new_C1236_;
  assign new_C1213_ = new_C1179_ | new_C1212_;
  assign new_C1212_ = new_C1233_ | new_C1232_;
  assign new_C1211_ = ~new_C1191_ & ~new_C1201_;
  assign new_C1210_ = new_C1191_ & new_C1201_;
  assign new_C1209_ = ~new_C1191_ | new_C1201_;
  assign new_C1208_ = new_C1175_ & ~new_C1176_;
  assign new_C1207_ = ~new_C1175_ & new_C1176_;
  assign new_C1206_ = new_C1228_ & ~new_C1229_;
  assign new_C1205_ = ~new_C1228_ & new_C1229_;
  assign new_C1204_ = ~new_C1227_ | ~new_C1226_;
  assign new_C1203_ = new_C1219_ | new_C1218_;
  assign new_C1202_ = new_C1225_ | new_C1224_;
  assign new_C1201_ = new_C1215_ | new_C1217_;
  assign new_C1200_ = ~new_C1222_ | ~new_C1223_;
  assign new_C1199_ = new_C1175_ & ~new_C1176_;
  assign new_C1198_ = new_C1189_ & ~new_C1201_;
  assign new_C1197_ = ~new_C1189_ & new_C1201_;
  assign new_C1196_ = ~new_C1187_ & new_C1213_;
  assign new_C1195_ = new_C1211_ | new_C1210_;
  assign new_C1194_ = new_C1208_ | new_C1207_;
  assign new_C1193_ = new_C1176_ | new_C1209_;
  assign new_C1192_ = new_C1201_ & new_C1204_;
  assign new_C1191_ = new_C1206_ | new_C1205_;
  assign new_C1190_ = new_C1201_ & new_C1200_;
  assign new_C1189_ = new_C1203_ & new_C1202_;
  assign new_C1188_ = new_C1198_ | new_C1197_;
  assign new_C1187_ = new_C1176_ | new_C1199_;
  assign C1186 = new_C1187_ | new_C1196_;
  assign C1185 = new_C1194_ & new_C1195_;
  assign C1184 = new_C1194_ & new_C1193_;
  assign C1183 = new_C1192_ | new_C1191_;
  assign C1182 = new_C1190_ | new_C1189_;
  assign C1181 = new_C1188_ & new_C1187_;
  assign new_C1180_ = new_C9293_;
  assign new_C1179_ = new_C9226_;
  assign new_C1178_ = new_C9159_;
  assign new_C1177_ = new_C9092_;
  assign new_C1176_ = new_C9025_;
  assign new_C1175_ = new_C8958_;
  assign new_C1174_ = ~new_C1113_ & new_C1127_;
  assign new_C1173_ = new_C1113_ & ~new_C1127_;
  assign new_C1172_ = new_C1113_ & ~new_C1127_;
  assign new_C1171_ = ~new_C1113_ & ~new_C1127_;
  assign new_C1170_ = new_C1113_ & new_C1127_;
  assign new_C1169_ = new_C1173_ | new_C1174_;
  assign new_C1168_ = ~new_C1113_ & new_C1127_;
  assign new_C1167_ = new_C1171_ | new_C1172_;
  assign new_C1166_ = ~new_C1142_ & ~new_C1162_;
  assign new_C1165_ = new_C1142_ & new_C1162_;
  assign new_C1164_ = ~new_C1109_ | ~new_C1134_;
  assign new_C1163_ = new_C1127_ & new_C1164_;
  assign new_C1162_ = new_C1110_ | new_C1111_;
  assign new_C1161_ = new_C1110_ | new_C1127_;
  assign new_C1160_ = ~new_C1127_ & ~new_C1163_;
  assign new_C1159_ = new_C1127_ | new_C1164_;
  assign new_C1158_ = new_C1110_ & ~new_C1111_;
  assign new_C1157_ = ~new_C1110_ & new_C1111_;
  assign new_C1156_ = new_C1120_ | new_C1153_;
  assign new_C1155_ = ~new_C1120_ & ~new_C1154_;
  assign new_C1154_ = new_C1120_ & new_C1153_;
  assign new_C1153_ = ~new_C1109_ | ~new_C1134_;
  assign new_C1152_ = ~new_C1110_ & new_C1120_;
  assign new_C1151_ = new_C1110_ & ~new_C1120_;
  assign new_C1150_ = new_C1112_ & new_C1149_;
  assign new_C1149_ = new_C1168_ | new_C1167_;
  assign new_C1148_ = ~new_C1112_ & new_C1147_;
  assign new_C1147_ = new_C1170_ | new_C1169_;
  assign new_C1146_ = new_C1112_ | new_C1145_;
  assign new_C1145_ = new_C1166_ | new_C1165_;
  assign new_C1144_ = ~new_C1124_ & ~new_C1134_;
  assign new_C1143_ = new_C1124_ & new_C1134_;
  assign new_C1142_ = ~new_C1124_ | new_C1134_;
  assign new_C1141_ = new_C1108_ & ~new_C1109_;
  assign new_C1140_ = ~new_C1108_ & new_C1109_;
  assign new_C1139_ = new_C1161_ & ~new_C1162_;
  assign new_C1138_ = ~new_C1161_ & new_C1162_;
  assign new_C1137_ = ~new_C1160_ | ~new_C1159_;
  assign new_C1136_ = new_C1152_ | new_C1151_;
  assign new_C1135_ = new_C1158_ | new_C1157_;
  assign new_C1134_ = new_C1148_ | new_C1150_;
  assign new_C1133_ = ~new_C1155_ | ~new_C1156_;
  assign new_C1132_ = new_C1108_ & ~new_C1109_;
  assign new_C1131_ = new_C1122_ & ~new_C1134_;
  assign new_C1130_ = ~new_C1122_ & new_C1134_;
  assign new_C1129_ = ~new_C1120_ & new_C1146_;
  assign new_C1128_ = new_C1144_ | new_C1143_;
  assign new_C1127_ = new_C1141_ | new_C1140_;
  assign new_C1126_ = new_C1109_ | new_C1142_;
  assign new_C1125_ = new_C1134_ & new_C1137_;
  assign new_C1124_ = new_C1139_ | new_C1138_;
  assign new_C1123_ = new_C1134_ & new_C1133_;
  assign new_C1122_ = new_C1136_ & new_C1135_;
  assign new_C1121_ = new_C1131_ | new_C1130_;
  assign new_C1120_ = new_C1109_ | new_C1132_;
  assign C1119 = new_C1120_ | new_C1129_;
  assign C1118 = new_C1127_ & new_C1128_;
  assign C1117 = new_C1127_ & new_C1126_;
  assign C1116 = new_C1125_ | new_C1124_;
  assign C1115 = new_C1123_ | new_C1122_;
  assign C1114 = new_C1121_ & new_C1120_;
  assign new_C1113_ = new_C8891_;
  assign new_C1112_ = new_C8824_;
  assign new_C1111_ = new_C8757_;
  assign new_C1110_ = new_C8690_;
  assign new_C1109_ = new_C8623_;
  assign new_C1108_ = new_C8556_;
  assign new_C1107_ = ~new_C1046_ & new_C1060_;
  assign new_C1106_ = new_C1046_ & ~new_C1060_;
  assign new_C1105_ = new_C1046_ & ~new_C1060_;
  assign new_C1104_ = ~new_C1046_ & ~new_C1060_;
  assign new_C1103_ = new_C1046_ & new_C1060_;
  assign new_C1102_ = new_C1106_ | new_C1107_;
  assign new_C1101_ = ~new_C1046_ & new_C1060_;
  assign new_C1100_ = new_C1104_ | new_C1105_;
  assign new_C1099_ = ~new_C1075_ & ~new_C1095_;
  assign new_C1098_ = new_C1075_ & new_C1095_;
  assign new_C1097_ = ~new_C1042_ | ~new_C1067_;
  assign new_C1096_ = new_C1060_ & new_C1097_;
  assign new_C1095_ = new_C1043_ | new_C1044_;
  assign new_C1094_ = new_C1043_ | new_C1060_;
  assign new_C1093_ = ~new_C1060_ & ~new_C1096_;
  assign new_C1092_ = new_C1060_ | new_C1097_;
  assign new_C1091_ = new_C1043_ & ~new_C1044_;
  assign new_C1090_ = ~new_C1043_ & new_C1044_;
  assign new_C1089_ = new_C1053_ | new_C1086_;
  assign new_C1088_ = ~new_C1053_ & ~new_C1087_;
  assign new_C1087_ = new_C1053_ & new_C1086_;
  assign new_C1086_ = ~new_C1042_ | ~new_C1067_;
  assign new_C1085_ = ~new_C1043_ & new_C1053_;
  assign new_C1084_ = new_C1043_ & ~new_C1053_;
  assign new_C1083_ = new_C1045_ & new_C1082_;
  assign new_C1082_ = new_C1101_ | new_C1100_;
  assign new_C1081_ = ~new_C1045_ & new_C1080_;
  assign new_C1080_ = new_C1103_ | new_C1102_;
  assign new_C1079_ = new_C1045_ | new_C1078_;
  assign new_C1078_ = new_C1099_ | new_C1098_;
  assign new_C1077_ = ~new_C1057_ & ~new_C1067_;
  assign new_C1076_ = new_C1057_ & new_C1067_;
  assign new_C1075_ = ~new_C1057_ | new_C1067_;
  assign new_C1074_ = new_C1041_ & ~new_C1042_;
  assign new_C1073_ = ~new_C1041_ & new_C1042_;
  assign new_C1072_ = new_C1094_ & ~new_C1095_;
  assign new_C1071_ = ~new_C1094_ & new_C1095_;
  assign new_C1070_ = ~new_C1093_ | ~new_C1092_;
  assign new_C1069_ = new_C1085_ | new_C1084_;
  assign new_C1068_ = new_C1091_ | new_C1090_;
  assign new_C1067_ = new_C1081_ | new_C1083_;
  assign new_C1066_ = ~new_C1088_ | ~new_C1089_;
  assign new_C1065_ = new_C1041_ & ~new_C1042_;
  assign new_C1064_ = new_C1055_ & ~new_C1067_;
  assign new_C1063_ = ~new_C1055_ & new_C1067_;
  assign new_C1062_ = ~new_C1053_ & new_C1079_;
  assign new_C1061_ = new_C1077_ | new_C1076_;
  assign new_C1060_ = new_C1074_ | new_C1073_;
  assign new_C1059_ = new_C1042_ | new_C1075_;
  assign new_C1058_ = new_C1067_ & new_C1070_;
  assign new_C1057_ = new_C1072_ | new_C1071_;
  assign new_C1056_ = new_C1067_ & new_C1066_;
  assign new_C1055_ = new_C1069_ & new_C1068_;
  assign new_C1054_ = new_C1064_ | new_C1063_;
  assign new_C1053_ = new_C1042_ | new_C1065_;
  assign C1052 = new_C1053_ | new_C1062_;
  assign C1051 = new_C1060_ & new_C1061_;
  assign C1050 = new_C1060_ & new_C1059_;
  assign C1049 = new_C1058_ | new_C1057_;
  assign C1048 = new_C1056_ | new_C1055_;
  assign C1047 = new_C1054_ & new_C1053_;
  assign new_C1046_ = new_C8489_;
  assign new_C1045_ = new_C8422_;
  assign new_C1044_ = new_C8355_;
  assign new_C1043_ = new_C8288_;
  assign new_C1042_ = new_C8221_;
  assign new_C1041_ = new_C8154_;
  assign new_C1040_ = ~new_C979_ & new_C993_;
  assign new_C1039_ = new_C979_ & ~new_C993_;
  assign new_C1038_ = new_C979_ & ~new_C993_;
  assign new_C1037_ = ~new_C979_ & ~new_C993_;
  assign new_C1036_ = new_C979_ & new_C993_;
  assign new_C1035_ = new_C1039_ | new_C1040_;
  assign new_C1034_ = ~new_C979_ & new_C993_;
  assign new_C1033_ = new_C1037_ | new_C1038_;
  assign new_C1032_ = ~new_C1008_ & ~new_C1028_;
  assign new_C1031_ = new_C1008_ & new_C1028_;
  assign new_C1030_ = ~new_C975_ | ~new_C1000_;
  assign new_C1029_ = new_C993_ & new_C1030_;
  assign new_C1028_ = new_C976_ | new_C977_;
  assign new_C1027_ = new_C976_ | new_C993_;
  assign new_C1026_ = ~new_C993_ & ~new_C1029_;
  assign new_C1025_ = new_C993_ | new_C1030_;
  assign new_C1024_ = new_C976_ & ~new_C977_;
  assign new_C1023_ = ~new_C976_ & new_C977_;
  assign new_C1022_ = new_C986_ | new_C1019_;
  assign new_C1021_ = ~new_C986_ & ~new_C1020_;
  assign new_C1020_ = new_C986_ & new_C1019_;
  assign new_C1019_ = ~new_C975_ | ~new_C1000_;
  assign new_C1018_ = ~new_C976_ & new_C986_;
  assign new_C1017_ = new_C976_ & ~new_C986_;
  assign new_C1016_ = new_C978_ & new_C1015_;
  assign new_C1015_ = new_C1034_ | new_C1033_;
  assign new_C1014_ = ~new_C978_ & new_C1013_;
  assign new_C1013_ = new_C1036_ | new_C1035_;
  assign new_C1012_ = new_C978_ | new_C1011_;
  assign new_C1011_ = new_C1032_ | new_C1031_;
  assign new_C1010_ = ~new_C990_ & ~new_C1000_;
  assign new_C1009_ = new_C990_ & new_C1000_;
  assign new_C1008_ = ~new_C990_ | new_C1000_;
  assign new_C1007_ = new_C974_ & ~new_C975_;
  assign new_C1006_ = ~new_C974_ & new_C975_;
  assign new_C1005_ = new_C1027_ & ~new_C1028_;
  assign new_C1004_ = ~new_C1027_ & new_C1028_;
  assign new_C1003_ = ~new_C1026_ | ~new_C1025_;
  assign new_C1002_ = new_C1018_ | new_C1017_;
  assign new_C1001_ = new_C1024_ | new_C1023_;
  assign new_C1000_ = new_C1014_ | new_C1016_;
  assign new_C999_ = ~new_C1021_ | ~new_C1022_;
  assign new_C998_ = new_C974_ & ~new_C975_;
  assign new_C997_ = new_C988_ & ~new_C1000_;
  assign new_C996_ = ~new_C988_ & new_C1000_;
  assign new_C995_ = ~new_C986_ & new_C1012_;
  assign new_C994_ = new_C1010_ | new_C1009_;
  assign new_C993_ = new_C1007_ | new_C1006_;
  assign new_C992_ = new_C975_ | new_C1008_;
  assign new_C991_ = new_C1000_ & new_C1003_;
  assign new_C990_ = new_C1005_ | new_C1004_;
  assign new_C989_ = new_C1000_ & new_C999_;
  assign new_C988_ = new_C1002_ & new_C1001_;
  assign new_C987_ = new_C997_ | new_C996_;
  assign new_C986_ = new_C975_ | new_C998_;
  assign C985 = new_C986_ | new_C995_;
  assign C984 = new_C993_ & new_C994_;
  assign C983 = new_C993_ & new_C992_;
  assign C982 = new_C991_ | new_C990_;
  assign C981 = new_C989_ | new_C988_;
  assign C980 = new_C987_ & new_C986_;
  assign new_C979_ = new_C8087_;
  assign new_C978_ = new_C8020_;
  assign new_C977_ = new_C7953_;
  assign new_C976_ = new_C7886_;
  assign new_C975_ = new_C7819_;
  assign new_C974_ = new_C7752_;
  assign new_C973_ = ~new_C912_ & new_C926_;
  assign new_C972_ = new_C912_ & ~new_C926_;
  assign new_C971_ = new_C912_ & ~new_C926_;
  assign new_C970_ = ~new_C912_ & ~new_C926_;
  assign new_C969_ = new_C912_ & new_C926_;
  assign new_C968_ = new_C972_ | new_C973_;
  assign new_C967_ = ~new_C912_ & new_C926_;
  assign new_C966_ = new_C970_ | new_C971_;
  assign new_C965_ = ~new_C941_ & ~new_C961_;
  assign new_C964_ = new_C941_ & new_C961_;
  assign new_C963_ = ~new_C908_ | ~new_C933_;
  assign new_C962_ = new_C926_ & new_C963_;
  assign new_C961_ = new_C909_ | new_C910_;
  assign new_C960_ = new_C909_ | new_C926_;
  assign new_C959_ = ~new_C926_ & ~new_C962_;
  assign new_C958_ = new_C926_ | new_C963_;
  assign new_C957_ = new_C909_ & ~new_C910_;
  assign new_C956_ = ~new_C909_ & new_C910_;
  assign new_C955_ = new_C919_ | new_C952_;
  assign new_C954_ = ~new_C919_ & ~new_C953_;
  assign new_C953_ = new_C919_ & new_C952_;
  assign new_C952_ = ~new_C908_ | ~new_C933_;
  assign new_C951_ = ~new_C909_ & new_C919_;
  assign new_C950_ = new_C909_ & ~new_C919_;
  assign new_C949_ = new_C911_ & new_C948_;
  assign new_C948_ = new_C967_ | new_C966_;
  assign new_C947_ = ~new_C911_ & new_C946_;
  assign new_C946_ = new_C969_ | new_C968_;
  assign new_C945_ = new_C911_ | new_C944_;
  assign new_C944_ = new_C965_ | new_C964_;
  assign new_C943_ = ~new_C923_ & ~new_C933_;
  assign new_C942_ = new_C923_ & new_C933_;
  assign new_C941_ = ~new_C923_ | new_C933_;
  assign new_C940_ = new_C907_ & ~new_C908_;
  assign new_C939_ = ~new_C907_ & new_C908_;
  assign new_C938_ = new_C960_ & ~new_C961_;
  assign new_C937_ = ~new_C960_ & new_C961_;
  assign new_C936_ = ~new_C959_ | ~new_C958_;
  assign new_C935_ = new_C951_ | new_C950_;
  assign new_C934_ = new_C957_ | new_C956_;
  assign new_C933_ = new_C947_ | new_C949_;
  assign new_C932_ = ~new_C954_ | ~new_C955_;
  assign new_C931_ = new_C907_ & ~new_C908_;
  assign new_C930_ = new_C921_ & ~new_C933_;
  assign new_C929_ = ~new_C921_ & new_C933_;
  assign new_C928_ = ~new_C919_ & new_C945_;
  assign new_C927_ = new_C943_ | new_C942_;
  assign new_C926_ = new_C940_ | new_C939_;
  assign new_C925_ = new_C908_ | new_C941_;
  assign new_C924_ = new_C933_ & new_C936_;
  assign new_C923_ = new_C938_ | new_C937_;
  assign new_C922_ = new_C933_ & new_C932_;
  assign new_C921_ = new_C935_ & new_C934_;
  assign new_C920_ = new_C930_ | new_C929_;
  assign new_C919_ = new_C908_ | new_C931_;
  assign C918 = new_C919_ | new_C928_;
  assign C917 = new_C926_ & new_C927_;
  assign C916 = new_C926_ & new_C925_;
  assign C915 = new_C924_ | new_C923_;
  assign C914 = new_C922_ | new_C921_;
  assign C913 = new_C920_ & new_C919_;
  assign new_C912_ = new_C7685_;
  assign new_C911_ = new_C7618_;
  assign new_C910_ = new_C7551_;
  assign new_C909_ = new_C7484_;
  assign new_C908_ = new_C7417_;
  assign new_C907_ = new_C7350_;
  assign new_C906_ = ~new_C845_ & new_C859_;
  assign new_C905_ = new_C845_ & ~new_C859_;
  assign new_C904_ = new_C845_ & ~new_C859_;
  assign new_C903_ = ~new_C845_ & ~new_C859_;
  assign new_C902_ = new_C845_ & new_C859_;
  assign new_C901_ = new_C905_ | new_C906_;
  assign new_C900_ = ~new_C845_ & new_C859_;
  assign new_C899_ = new_C903_ | new_C904_;
  assign new_C898_ = ~new_C874_ & ~new_C894_;
  assign new_C897_ = new_C874_ & new_C894_;
  assign new_C896_ = ~new_C841_ | ~new_C866_;
  assign new_C895_ = new_C859_ & new_C896_;
  assign new_C894_ = new_C842_ | new_C843_;
  assign new_C893_ = new_C842_ | new_C859_;
  assign new_C892_ = ~new_C859_ & ~new_C895_;
  assign new_C891_ = new_C859_ | new_C896_;
  assign new_C890_ = new_C842_ & ~new_C843_;
  assign new_C889_ = ~new_C842_ & new_C843_;
  assign new_C888_ = new_C852_ | new_C885_;
  assign new_C887_ = ~new_C852_ & ~new_C886_;
  assign new_C886_ = new_C852_ & new_C885_;
  assign new_C885_ = ~new_C841_ | ~new_C866_;
  assign new_C884_ = ~new_C842_ & new_C852_;
  assign new_C883_ = new_C842_ & ~new_C852_;
  assign new_C882_ = new_C844_ & new_C881_;
  assign new_C881_ = new_C900_ | new_C899_;
  assign new_C880_ = ~new_C844_ & new_C879_;
  assign new_C879_ = new_C902_ | new_C901_;
  assign new_C878_ = new_C844_ | new_C877_;
  assign new_C877_ = new_C898_ | new_C897_;
  assign new_C876_ = ~new_C856_ & ~new_C866_;
  assign new_C875_ = new_C856_ & new_C866_;
  assign new_C874_ = ~new_C856_ | new_C866_;
  assign new_C873_ = new_C840_ & ~new_C841_;
  assign new_C872_ = ~new_C840_ & new_C841_;
  assign new_C871_ = new_C893_ & ~new_C894_;
  assign new_C870_ = ~new_C893_ & new_C894_;
  assign new_C869_ = ~new_C892_ | ~new_C891_;
  assign new_C868_ = new_C884_ | new_C883_;
  assign new_C867_ = new_C890_ | new_C889_;
  assign new_C866_ = new_C880_ | new_C882_;
  assign new_C865_ = ~new_C887_ | ~new_C888_;
  assign new_C864_ = new_C840_ & ~new_C841_;
  assign new_C863_ = new_C854_ & ~new_C866_;
  assign new_C862_ = ~new_C854_ & new_C866_;
  assign new_C861_ = ~new_C852_ & new_C878_;
  assign new_C860_ = new_C876_ | new_C875_;
  assign new_C859_ = new_C873_ | new_C872_;
  assign new_C858_ = new_C841_ | new_C874_;
  assign new_C857_ = new_C866_ & new_C869_;
  assign new_C856_ = new_C871_ | new_C870_;
  assign new_C855_ = new_C866_ & new_C865_;
  assign new_C854_ = new_C868_ & new_C867_;
  assign new_C853_ = new_C863_ | new_C862_;
  assign new_C852_ = new_C841_ | new_C864_;
  assign C851 = new_C852_ | new_C861_;
  assign C850 = new_C859_ & new_C860_;
  assign C849 = new_C859_ & new_C858_;
  assign C848 = new_C857_ | new_C856_;
  assign C847 = new_C855_ | new_C854_;
  assign C846 = new_C853_ & new_C852_;
  assign new_C845_ = new_C7283_;
  assign new_C844_ = new_C7216_;
  assign new_C843_ = new_C7149_;
  assign new_C842_ = new_C7082_;
  assign new_C841_ = new_C7015_;
  assign new_C840_ = new_C6948_;
  assign new_C839_ = ~new_C778_ & new_C792_;
  assign new_C838_ = new_C778_ & ~new_C792_;
  assign new_C837_ = new_C778_ & ~new_C792_;
  assign new_C836_ = ~new_C778_ & ~new_C792_;
  assign new_C835_ = new_C778_ & new_C792_;
  assign new_C834_ = new_C838_ | new_C839_;
  assign new_C833_ = ~new_C778_ & new_C792_;
  assign new_C832_ = new_C836_ | new_C837_;
  assign new_C831_ = ~new_C807_ & ~new_C827_;
  assign new_C830_ = new_C807_ & new_C827_;
  assign new_C829_ = ~new_C774_ | ~new_C799_;
  assign new_C828_ = new_C792_ & new_C829_;
  assign new_C827_ = new_C775_ | new_C776_;
  assign new_C826_ = new_C775_ | new_C792_;
  assign new_C825_ = ~new_C792_ & ~new_C828_;
  assign new_C824_ = new_C792_ | new_C829_;
  assign new_C823_ = new_C775_ & ~new_C776_;
  assign new_C822_ = ~new_C775_ & new_C776_;
  assign new_C821_ = new_C785_ | new_C818_;
  assign new_C820_ = ~new_C785_ & ~new_C819_;
  assign new_C819_ = new_C785_ & new_C818_;
  assign new_C818_ = ~new_C774_ | ~new_C799_;
  assign new_C817_ = ~new_C775_ & new_C785_;
  assign new_C816_ = new_C775_ & ~new_C785_;
  assign new_C815_ = new_C777_ & new_C814_;
  assign new_C814_ = new_C833_ | new_C832_;
  assign new_C813_ = ~new_C777_ & new_C812_;
  assign new_C812_ = new_C835_ | new_C834_;
  assign new_C811_ = new_C777_ | new_C810_;
  assign new_C810_ = new_C831_ | new_C830_;
  assign new_C809_ = ~new_C789_ & ~new_C799_;
  assign new_C808_ = new_C789_ & new_C799_;
  assign new_C807_ = ~new_C789_ | new_C799_;
  assign new_C806_ = new_C773_ & ~new_C774_;
  assign new_C805_ = ~new_C773_ & new_C774_;
  assign new_C804_ = new_C826_ & ~new_C827_;
  assign new_C803_ = ~new_C826_ & new_C827_;
  assign new_C802_ = ~new_C825_ | ~new_C824_;
  assign new_C801_ = new_C817_ | new_C816_;
  assign new_C800_ = new_C823_ | new_C822_;
  assign new_C799_ = new_C813_ | new_C815_;
  assign new_C798_ = ~new_C820_ | ~new_C821_;
  assign new_C797_ = new_C773_ & ~new_C774_;
  assign new_C796_ = new_C787_ & ~new_C799_;
  assign new_C795_ = ~new_C787_ & new_C799_;
  assign new_C794_ = ~new_C785_ & new_C811_;
  assign new_C793_ = new_C809_ | new_C808_;
  assign new_C792_ = new_C806_ | new_C805_;
  assign new_C791_ = new_C774_ | new_C807_;
  assign new_C790_ = new_C799_ & new_C802_;
  assign new_C789_ = new_C804_ | new_C803_;
  assign new_C788_ = new_C799_ & new_C798_;
  assign new_C787_ = new_C801_ & new_C800_;
  assign new_C786_ = new_C796_ | new_C795_;
  assign new_C785_ = new_C774_ | new_C797_;
  assign C784 = new_C785_ | new_C794_;
  assign C783 = new_C792_ & new_C793_;
  assign C782 = new_C792_ & new_C791_;
  assign C781 = new_C790_ | new_C789_;
  assign C780 = new_C788_ | new_C787_;
  assign C779 = new_C786_ & new_C785_;
  assign new_C778_ = new_C6881_;
  assign new_C777_ = new_C6814_;
  assign new_C776_ = new_C6747_;
  assign new_C775_ = new_C6680_;
  assign new_C774_ = new_C6613_;
  assign new_C773_ = new_C6546_;
  assign new_C772_ = ~new_C711_ & new_C725_;
  assign new_C771_ = new_C711_ & ~new_C725_;
  assign new_C770_ = new_C711_ & ~new_C725_;
  assign new_C769_ = ~new_C711_ & ~new_C725_;
  assign new_C768_ = new_C711_ & new_C725_;
  assign new_C767_ = new_C771_ | new_C772_;
  assign new_C766_ = ~new_C711_ & new_C725_;
  assign new_C765_ = new_C769_ | new_C770_;
  assign new_C764_ = ~new_C740_ & ~new_C760_;
  assign new_C763_ = new_C740_ & new_C760_;
  assign new_C762_ = ~new_C707_ | ~new_C732_;
  assign new_C761_ = new_C725_ & new_C762_;
  assign new_C760_ = new_C708_ | new_C709_;
  assign new_C759_ = new_C708_ | new_C725_;
  assign new_C758_ = ~new_C725_ & ~new_C761_;
  assign new_C757_ = new_C725_ | new_C762_;
  assign new_C756_ = new_C708_ & ~new_C709_;
  assign new_C755_ = ~new_C708_ & new_C709_;
  assign new_C754_ = new_C718_ | new_C751_;
  assign new_C753_ = ~new_C718_ & ~new_C752_;
  assign new_C752_ = new_C718_ & new_C751_;
  assign new_C751_ = ~new_C707_ | ~new_C732_;
  assign new_C750_ = ~new_C708_ & new_C718_;
  assign new_C749_ = new_C708_ & ~new_C718_;
  assign new_C748_ = new_C710_ & new_C747_;
  assign new_C747_ = new_C766_ | new_C765_;
  assign new_C746_ = ~new_C710_ & new_C745_;
  assign new_C745_ = new_C768_ | new_C767_;
  assign new_C744_ = new_C710_ | new_C743_;
  assign new_C743_ = new_C764_ | new_C763_;
  assign new_C742_ = ~new_C722_ & ~new_C732_;
  assign new_C741_ = new_C722_ & new_C732_;
  assign new_C740_ = ~new_C722_ | new_C732_;
  assign new_C739_ = new_C706_ & ~new_C707_;
  assign new_C738_ = ~new_C706_ & new_C707_;
  assign new_C737_ = new_C759_ & ~new_C760_;
  assign new_C736_ = ~new_C759_ & new_C760_;
  assign new_C735_ = ~new_C758_ | ~new_C757_;
  assign new_C734_ = new_C750_ | new_C749_;
  assign new_C733_ = new_C756_ | new_C755_;
  assign new_C732_ = new_C746_ | new_C748_;
  assign new_C731_ = ~new_C753_ | ~new_C754_;
  assign new_C730_ = new_C706_ & ~new_C707_;
  assign new_C729_ = new_C720_ & ~new_C732_;
  assign new_C728_ = ~new_C720_ & new_C732_;
  assign new_C727_ = ~new_C718_ & new_C744_;
  assign new_C726_ = new_C742_ | new_C741_;
  assign new_C725_ = new_C739_ | new_C738_;
  assign new_C724_ = new_C707_ | new_C740_;
  assign new_C723_ = new_C732_ & new_C735_;
  assign new_C722_ = new_C737_ | new_C736_;
  assign new_C721_ = new_C732_ & new_C731_;
  assign new_C720_ = new_C734_ & new_C733_;
  assign new_C719_ = new_C729_ | new_C728_;
  assign new_C718_ = new_C707_ | new_C730_;
  assign C717 = new_C718_ | new_C727_;
  assign C716 = new_C725_ & new_C726_;
  assign C715 = new_C725_ & new_C724_;
  assign C714 = new_C723_ | new_C722_;
  assign C713 = new_C721_ | new_C720_;
  assign C712 = new_C719_ & new_C718_;
  assign new_C711_ = new_C6479_;
  assign new_C710_ = new_C6412_;
  assign new_C709_ = new_C6345_;
  assign new_C708_ = new_C6278_;
  assign new_C707_ = new_C6211_;
  assign new_C706_ = new_C6144_;
  assign new_C705_ = ~new_C644_ & new_C658_;
  assign new_C704_ = new_C644_ & ~new_C658_;
  assign new_C703_ = new_C644_ & ~new_C658_;
  assign new_C702_ = ~new_C644_ & ~new_C658_;
  assign new_C701_ = new_C644_ & new_C658_;
  assign new_C700_ = new_C704_ | new_C705_;
  assign new_C699_ = ~new_C644_ & new_C658_;
  assign new_C698_ = new_C702_ | new_C703_;
  assign new_C697_ = ~new_C673_ & ~new_C693_;
  assign new_C696_ = new_C673_ & new_C693_;
  assign new_C695_ = ~new_C640_ | ~new_C665_;
  assign new_C694_ = new_C658_ & new_C695_;
  assign new_C693_ = new_C641_ | new_C642_;
  assign new_C692_ = new_C641_ | new_C658_;
  assign new_C691_ = ~new_C658_ & ~new_C694_;
  assign new_C690_ = new_C658_ | new_C695_;
  assign new_C689_ = new_C641_ & ~new_C642_;
  assign new_C688_ = ~new_C641_ & new_C642_;
  assign new_C687_ = new_C651_ | new_C684_;
  assign new_C686_ = ~new_C651_ & ~new_C685_;
  assign new_C685_ = new_C651_ & new_C684_;
  assign new_C684_ = ~new_C640_ | ~new_C665_;
  assign new_C683_ = ~new_C641_ & new_C651_;
  assign new_C682_ = new_C641_ & ~new_C651_;
  assign new_C681_ = new_C643_ & new_C680_;
  assign new_C680_ = new_C699_ | new_C698_;
  assign new_C679_ = ~new_C643_ & new_C678_;
  assign new_C678_ = new_C701_ | new_C700_;
  assign new_C677_ = new_C643_ | new_C676_;
  assign new_C676_ = new_C697_ | new_C696_;
  assign new_C675_ = ~new_C655_ & ~new_C665_;
  assign new_C674_ = new_C655_ & new_C665_;
  assign new_C673_ = ~new_C655_ | new_C665_;
  assign new_C672_ = new_C639_ & ~new_C640_;
  assign new_C671_ = ~new_C639_ & new_C640_;
  assign new_C670_ = new_C692_ & ~new_C693_;
  assign new_C669_ = ~new_C692_ & new_C693_;
  assign new_C668_ = ~new_C691_ | ~new_C690_;
  assign new_C667_ = new_C683_ | new_C682_;
  assign new_C666_ = new_C689_ | new_C688_;
  assign new_C665_ = new_C679_ | new_C681_;
  assign new_C664_ = ~new_C686_ | ~new_C687_;
  assign new_C663_ = new_C639_ & ~new_C640_;
  assign new_C662_ = new_C653_ & ~new_C665_;
  assign new_C661_ = ~new_C653_ & new_C665_;
  assign new_C660_ = ~new_C651_ & new_C677_;
  assign new_C659_ = new_C675_ | new_C674_;
  assign new_C658_ = new_C672_ | new_C671_;
  assign new_C657_ = new_C640_ | new_C673_;
  assign new_C656_ = new_C665_ & new_C668_;
  assign new_C655_ = new_C670_ | new_C669_;
  assign new_C654_ = new_C665_ & new_C664_;
  assign new_C653_ = new_C667_ & new_C666_;
  assign new_C652_ = new_C662_ | new_C661_;
  assign new_C651_ = new_C640_ | new_C663_;
  assign C650 = new_C651_ | new_C660_;
  assign C649 = new_C658_ & new_C659_;
  assign C648 = new_C658_ & new_C657_;
  assign C647 = new_C656_ | new_C655_;
  assign C646 = new_C654_ | new_C653_;
  assign C645 = new_C652_ & new_C651_;
  assign new_C644_ = new_C6077_;
  assign new_C643_ = new_C6010_;
  assign new_C642_ = new_C5943_;
  assign new_C641_ = new_C5876_;
  assign new_C640_ = new_C5809_;
  assign new_C639_ = new_C5742_;
  assign new_C638_ = ~new_C577_ & new_C591_;
  assign new_C637_ = new_C577_ & ~new_C591_;
  assign new_C636_ = new_C577_ & ~new_C591_;
  assign new_C635_ = ~new_C577_ & ~new_C591_;
  assign new_C634_ = new_C577_ & new_C591_;
  assign new_C633_ = new_C637_ | new_C638_;
  assign new_C632_ = ~new_C577_ & new_C591_;
  assign new_C631_ = new_C635_ | new_C636_;
  assign new_C630_ = ~new_C606_ & ~new_C626_;
  assign new_C629_ = new_C606_ & new_C626_;
  assign new_C628_ = ~new_C573_ | ~new_C598_;
  assign new_C627_ = new_C591_ & new_C628_;
  assign new_C626_ = new_C574_ | new_C575_;
  assign new_C625_ = new_C574_ | new_C591_;
  assign new_C624_ = ~new_C591_ & ~new_C627_;
  assign new_C623_ = new_C591_ | new_C628_;
  assign new_C622_ = new_C574_ & ~new_C575_;
  assign new_C621_ = ~new_C574_ & new_C575_;
  assign new_C620_ = new_C584_ | new_C617_;
  assign new_C619_ = ~new_C584_ & ~new_C618_;
  assign new_C618_ = new_C584_ & new_C617_;
  assign new_C617_ = ~new_C573_ | ~new_C598_;
  assign new_C616_ = ~new_C574_ & new_C584_;
  assign new_C615_ = new_C574_ & ~new_C584_;
  assign new_C614_ = new_C576_ & new_C613_;
  assign new_C613_ = new_C632_ | new_C631_;
  assign new_C612_ = ~new_C576_ & new_C611_;
  assign new_C611_ = new_C634_ | new_C633_;
  assign new_C610_ = new_C576_ | new_C609_;
  assign new_C609_ = new_C630_ | new_C629_;
  assign new_C608_ = ~new_C588_ & ~new_C598_;
  assign new_C607_ = new_C588_ & new_C598_;
  assign new_C606_ = ~new_C588_ | new_C598_;
  assign new_C605_ = new_C572_ & ~new_C573_;
  assign new_C604_ = ~new_C572_ & new_C573_;
  assign new_C603_ = new_C625_ & ~new_C626_;
  assign new_C602_ = ~new_C625_ & new_C626_;
  assign new_C601_ = ~new_C624_ | ~new_C623_;
  assign new_C600_ = new_C616_ | new_C615_;
  assign new_C599_ = new_C622_ | new_C621_;
  assign new_C598_ = new_C612_ | new_C614_;
  assign new_C597_ = ~new_C619_ | ~new_C620_;
  assign new_C596_ = new_C572_ & ~new_C573_;
  assign new_C595_ = new_C586_ & ~new_C598_;
  assign new_C594_ = ~new_C586_ & new_C598_;
  assign new_C593_ = ~new_C584_ & new_C610_;
  assign new_C592_ = new_C608_ | new_C607_;
  assign new_C591_ = new_C605_ | new_C604_;
  assign new_C590_ = new_C573_ | new_C606_;
  assign new_C589_ = new_C598_ & new_C601_;
  assign new_C588_ = new_C603_ | new_C602_;
  assign new_C587_ = new_C598_ & new_C597_;
  assign new_C586_ = new_C600_ & new_C599_;
  assign new_C585_ = new_C595_ | new_C594_;
  assign new_C584_ = new_C573_ | new_C596_;
  assign C583 = new_C584_ | new_C593_;
  assign C582 = new_C591_ & new_C592_;
  assign C581 = new_C591_ & new_C590_;
  assign C580 = new_C589_ | new_C588_;
  assign C579 = new_C587_ | new_C586_;
  assign C578 = new_C585_ & new_C584_;
  assign new_C577_ = new_C5675_;
  assign new_C576_ = new_C5608_;
  assign new_C575_ = new_C5541_;
  assign new_C574_ = new_C5474_;
  assign new_C573_ = new_C5407_;
  assign new_C572_ = new_C5340_;
  assign new_C571_ = ~new_C510_ & new_C524_;
  assign new_C570_ = new_C510_ & ~new_C524_;
  assign new_C569_ = new_C510_ & ~new_C524_;
  assign new_C568_ = ~new_C510_ & ~new_C524_;
  assign new_C567_ = new_C510_ & new_C524_;
  assign new_C566_ = new_C570_ | new_C571_;
  assign new_C565_ = ~new_C510_ & new_C524_;
  assign new_C564_ = new_C568_ | new_C569_;
  assign new_C563_ = ~new_C539_ & ~new_C559_;
  assign new_C562_ = new_C539_ & new_C559_;
  assign new_C561_ = ~new_C506_ | ~new_C531_;
  assign new_C560_ = new_C524_ & new_C561_;
  assign new_C559_ = new_C507_ | new_C508_;
  assign new_C558_ = new_C507_ | new_C524_;
  assign new_C557_ = ~new_C524_ & ~new_C560_;
  assign new_C556_ = new_C524_ | new_C561_;
  assign new_C555_ = new_C507_ & ~new_C508_;
  assign new_C554_ = ~new_C507_ & new_C508_;
  assign new_C553_ = new_C517_ | new_C550_;
  assign new_C552_ = ~new_C517_ & ~new_C551_;
  assign new_C551_ = new_C517_ & new_C550_;
  assign new_C550_ = ~new_C506_ | ~new_C531_;
  assign new_C549_ = ~new_C507_ & new_C517_;
  assign new_C548_ = new_C507_ & ~new_C517_;
  assign new_C547_ = new_C509_ & new_C546_;
  assign new_C546_ = new_C565_ | new_C564_;
  assign new_C545_ = ~new_C509_ & new_C544_;
  assign new_C544_ = new_C567_ | new_C566_;
  assign new_C543_ = new_C509_ | new_C542_;
  assign new_C542_ = new_C563_ | new_C562_;
  assign new_C541_ = ~new_C521_ & ~new_C531_;
  assign new_C540_ = new_C521_ & new_C531_;
  assign new_C539_ = ~new_C521_ | new_C531_;
  assign new_C538_ = new_C505_ & ~new_C506_;
  assign new_C537_ = ~new_C505_ & new_C506_;
  assign new_C536_ = new_C558_ & ~new_C559_;
  assign new_C535_ = ~new_C558_ & new_C559_;
  assign new_C534_ = ~new_C557_ | ~new_C556_;
  assign new_C533_ = new_C549_ | new_C548_;
  assign new_C532_ = new_C555_ | new_C554_;
  assign new_C531_ = new_C545_ | new_C547_;
  assign new_C530_ = ~new_C552_ | ~new_C553_;
  assign new_C529_ = new_C505_ & ~new_C506_;
  assign new_C528_ = new_C519_ & ~new_C531_;
  assign new_C527_ = ~new_C519_ & new_C531_;
  assign new_C526_ = ~new_C517_ & new_C543_;
  assign new_C525_ = new_C541_ | new_C540_;
  assign new_C524_ = new_C538_ | new_C537_;
  assign new_C523_ = new_C506_ | new_C539_;
  assign new_C522_ = new_C531_ & new_C534_;
  assign new_C521_ = new_C536_ | new_C535_;
  assign new_C520_ = new_C531_ & new_C530_;
  assign new_C519_ = new_C533_ & new_C532_;
  assign new_C518_ = new_C528_ | new_C527_;
  assign new_C517_ = new_C506_ | new_C529_;
  assign C516 = new_C517_ | new_C526_;
  assign C515 = new_C524_ & new_C525_;
  assign C514 = new_C524_ & new_C523_;
  assign C513 = new_C522_ | new_C521_;
  assign C512 = new_C520_ | new_C519_;
  assign C511 = new_C518_ & new_C517_;
  assign new_C510_ = new_C5273_;
  assign new_C509_ = new_C5206_;
  assign new_C508_ = new_C5139_;
  assign new_C507_ = new_C5072_;
  assign new_C506_ = new_C5005_;
  assign new_C505_ = new_C4938_;
  assign new_C504_ = ~new_C443_ & new_C457_;
  assign new_C503_ = new_C443_ & ~new_C457_;
  assign new_C502_ = new_C443_ & ~new_C457_;
  assign new_C501_ = ~new_C443_ & ~new_C457_;
  assign new_C500_ = new_C443_ & new_C457_;
  assign new_C499_ = new_C503_ | new_C504_;
  assign new_C498_ = ~new_C443_ & new_C457_;
  assign new_C497_ = new_C501_ | new_C502_;
  assign new_C496_ = ~new_C472_ & ~new_C492_;
  assign new_C495_ = new_C472_ & new_C492_;
  assign new_C494_ = ~new_C439_ | ~new_C464_;
  assign new_C493_ = new_C457_ & new_C494_;
  assign new_C492_ = new_C440_ | new_C441_;
  assign new_C491_ = new_C440_ | new_C457_;
  assign new_C490_ = ~new_C457_ & ~new_C493_;
  assign new_C489_ = new_C457_ | new_C494_;
  assign new_C488_ = new_C440_ & ~new_C441_;
  assign new_C487_ = ~new_C440_ & new_C441_;
  assign new_C486_ = new_C450_ | new_C483_;
  assign new_C485_ = ~new_C450_ & ~new_C484_;
  assign new_C484_ = new_C450_ & new_C483_;
  assign new_C483_ = ~new_C439_ | ~new_C464_;
  assign new_C482_ = ~new_C440_ & new_C450_;
  assign new_C481_ = new_C440_ & ~new_C450_;
  assign new_C480_ = new_C442_ & new_C479_;
  assign new_C479_ = new_C498_ | new_C497_;
  assign new_C478_ = ~new_C442_ & new_C477_;
  assign new_C477_ = new_C500_ | new_C499_;
  assign new_C476_ = new_C442_ | new_C475_;
  assign new_C475_ = new_C496_ | new_C495_;
  assign new_C474_ = ~new_C454_ & ~new_C464_;
  assign new_C473_ = new_C454_ & new_C464_;
  assign new_C472_ = ~new_C454_ | new_C464_;
  assign new_C471_ = new_C438_ & ~new_C439_;
  assign new_C470_ = ~new_C438_ & new_C439_;
  assign new_C469_ = new_C491_ & ~new_C492_;
  assign new_C468_ = ~new_C491_ & new_C492_;
  assign new_C467_ = ~new_C490_ | ~new_C489_;
  assign new_C466_ = new_C482_ | new_C481_;
  assign new_C465_ = new_C488_ | new_C487_;
  assign new_C464_ = new_C478_ | new_C480_;
  assign new_C463_ = ~new_C485_ | ~new_C486_;
  assign new_C462_ = new_C438_ & ~new_C439_;
  assign new_C461_ = new_C452_ & ~new_C464_;
  assign new_C460_ = ~new_C452_ & new_C464_;
  assign new_C459_ = ~new_C450_ & new_C476_;
  assign new_C458_ = new_C474_ | new_C473_;
  assign new_C457_ = new_C471_ | new_C470_;
  assign new_C456_ = new_C439_ | new_C472_;
  assign new_C455_ = new_C464_ & new_C467_;
  assign new_C454_ = new_C469_ | new_C468_;
  assign new_C453_ = new_C464_ & new_C463_;
  assign new_C452_ = new_C466_ & new_C465_;
  assign new_C451_ = new_C461_ | new_C460_;
  assign new_C450_ = new_C439_ | new_C462_;
  assign C449 = new_C450_ | new_C459_;
  assign C448 = new_C457_ & new_C458_;
  assign C447 = new_C457_ & new_C456_;
  assign C446 = new_C455_ | new_C454_;
  assign C445 = new_C453_ | new_C452_;
  assign C444 = new_C451_ & new_C450_;
  assign new_C443_ = new_C4871_;
  assign new_C442_ = new_C4804_;
  assign new_C441_ = new_C4737_;
  assign new_C440_ = new_C4670_;
  assign new_C439_ = new_C4603_;
  assign new_C438_ = new_C4536_;
  assign new_C437_ = ~new_C376_ & new_C390_;
  assign new_C436_ = new_C376_ & ~new_C390_;
  assign new_C435_ = new_C376_ & ~new_C390_;
  assign new_C434_ = ~new_C376_ & ~new_C390_;
  assign new_C433_ = new_C376_ & new_C390_;
  assign new_C432_ = new_C436_ | new_C437_;
  assign new_C431_ = ~new_C376_ & new_C390_;
  assign new_C430_ = new_C434_ | new_C435_;
  assign new_C429_ = ~new_C405_ & ~new_C425_;
  assign new_C428_ = new_C405_ & new_C425_;
  assign new_C427_ = ~new_C372_ | ~new_C397_;
  assign new_C426_ = new_C390_ & new_C427_;
  assign new_C425_ = new_C373_ | new_C374_;
  assign new_C424_ = new_C373_ | new_C390_;
  assign new_C423_ = ~new_C390_ & ~new_C426_;
  assign new_C422_ = new_C390_ | new_C427_;
  assign new_C421_ = new_C373_ & ~new_C374_;
  assign new_C420_ = ~new_C373_ & new_C374_;
  assign new_C419_ = new_C383_ | new_C416_;
  assign new_C418_ = ~new_C383_ & ~new_C417_;
  assign new_C417_ = new_C383_ & new_C416_;
  assign new_C416_ = ~new_C372_ | ~new_C397_;
  assign new_C415_ = ~new_C373_ & new_C383_;
  assign new_C414_ = new_C373_ & ~new_C383_;
  assign new_C413_ = new_C375_ & new_C412_;
  assign new_C412_ = new_C431_ | new_C430_;
  assign new_C411_ = ~new_C375_ & new_C410_;
  assign new_C410_ = new_C433_ | new_C432_;
  assign new_C409_ = new_C375_ | new_C408_;
  assign new_C408_ = new_C429_ | new_C428_;
  assign new_C407_ = ~new_C387_ & ~new_C397_;
  assign new_C406_ = new_C387_ & new_C397_;
  assign new_C405_ = ~new_C387_ | new_C397_;
  assign new_C404_ = new_C371_ & ~new_C372_;
  assign new_C403_ = ~new_C371_ & new_C372_;
  assign new_C402_ = new_C424_ & ~new_C425_;
  assign new_C401_ = ~new_C424_ & new_C425_;
  assign new_C400_ = ~new_C423_ | ~new_C422_;
  assign new_C399_ = new_C415_ | new_C414_;
  assign new_C398_ = new_C421_ | new_C420_;
  assign new_C397_ = new_C411_ | new_C413_;
  assign new_C396_ = ~new_C418_ | ~new_C419_;
  assign new_C395_ = new_C371_ & ~new_C372_;
  assign new_C394_ = new_C385_ & ~new_C397_;
  assign new_C393_ = ~new_C385_ & new_C397_;
  assign new_C392_ = ~new_C383_ & new_C409_;
  assign new_C391_ = new_C407_ | new_C406_;
  assign new_C390_ = new_C404_ | new_C403_;
  assign new_C389_ = new_C372_ | new_C405_;
  assign new_C388_ = new_C397_ & new_C400_;
  assign new_C387_ = new_C402_ | new_C401_;
  assign new_C386_ = new_C397_ & new_C396_;
  assign new_C385_ = new_C399_ & new_C398_;
  assign new_C384_ = new_C394_ | new_C393_;
  assign new_C383_ = new_C372_ | new_C395_;
  assign C382 = new_C383_ | new_C392_;
  assign C381 = new_C390_ & new_C391_;
  assign C380 = new_C390_ & new_C389_;
  assign C379 = new_C388_ | new_C387_;
  assign C378 = new_C386_ | new_C385_;
  assign C377 = new_C384_ & new_C383_;
  assign new_C376_ = new_C4469_;
  assign new_C375_ = new_C4402_;
  assign new_C374_ = new_C4335_;
  assign new_C373_ = new_C4268_;
  assign new_C372_ = new_C4201_;
  assign new_C371_ = new_C4134_;
  assign new_C370_ = ~new_C309_ & new_C323_;
  assign new_C369_ = new_C309_ & ~new_C323_;
  assign new_C368_ = new_C309_ & ~new_C323_;
  assign new_C367_ = ~new_C309_ & ~new_C323_;
  assign new_C366_ = new_C309_ & new_C323_;
  assign new_C365_ = new_C369_ | new_C370_;
  assign new_C364_ = ~new_C309_ & new_C323_;
  assign new_C363_ = new_C367_ | new_C368_;
  assign new_C362_ = ~new_C338_ & ~new_C358_;
  assign new_C361_ = new_C338_ & new_C358_;
  assign new_C360_ = ~new_C305_ | ~new_C330_;
  assign new_C359_ = new_C323_ & new_C360_;
  assign new_C358_ = new_C306_ | new_C307_;
  assign new_C357_ = new_C306_ | new_C323_;
  assign new_C356_ = ~new_C323_ & ~new_C359_;
  assign new_C355_ = new_C323_ | new_C360_;
  assign new_C354_ = new_C306_ & ~new_C307_;
  assign new_C353_ = ~new_C306_ & new_C307_;
  assign new_C352_ = new_C316_ | new_C349_;
  assign new_C351_ = ~new_C316_ & ~new_C350_;
  assign new_C350_ = new_C316_ & new_C349_;
  assign new_C349_ = ~new_C305_ | ~new_C330_;
  assign new_C348_ = ~new_C306_ & new_C316_;
  assign new_C347_ = new_C306_ & ~new_C316_;
  assign new_C346_ = new_C308_ & new_C345_;
  assign new_C345_ = new_C364_ | new_C363_;
  assign new_C344_ = ~new_C308_ & new_C343_;
  assign new_C343_ = new_C366_ | new_C365_;
  assign new_C342_ = new_C308_ | new_C341_;
  assign new_C341_ = new_C362_ | new_C361_;
  assign new_C340_ = ~new_C320_ & ~new_C330_;
  assign new_C339_ = new_C320_ & new_C330_;
  assign new_C338_ = ~new_C320_ | new_C330_;
  assign new_C337_ = new_C304_ & ~new_C305_;
  assign new_C336_ = ~new_C304_ & new_C305_;
  assign new_C335_ = new_C357_ & ~new_C358_;
  assign new_C334_ = ~new_C357_ & new_C358_;
  assign new_C333_ = ~new_C356_ | ~new_C355_;
  assign new_C332_ = new_C348_ | new_C347_;
  assign new_C331_ = new_C354_ | new_C353_;
  assign new_C330_ = new_C344_ | new_C346_;
  assign new_C329_ = ~new_C351_ | ~new_C352_;
  assign new_C328_ = new_C304_ & ~new_C305_;
  assign new_C327_ = new_C318_ & ~new_C330_;
  assign new_C326_ = ~new_C318_ & new_C330_;
  assign new_C325_ = ~new_C316_ & new_C342_;
  assign new_C324_ = new_C340_ | new_C339_;
  assign new_C323_ = new_C337_ | new_C336_;
  assign new_C322_ = new_C305_ | new_C338_;
  assign new_C321_ = new_C330_ & new_C333_;
  assign new_C320_ = new_C335_ | new_C334_;
  assign new_C319_ = new_C330_ & new_C329_;
  assign new_C318_ = new_C332_ & new_C331_;
  assign new_C317_ = new_C327_ | new_C326_;
  assign new_C316_ = new_C305_ | new_C328_;
  assign C315 = new_C316_ | new_C325_;
  assign C314 = new_C323_ & new_C324_;
  assign C313 = new_C323_ & new_C322_;
  assign C312 = new_C321_ | new_C320_;
  assign C311 = new_C319_ | new_C318_;
  assign C310 = new_C317_ & new_C316_;
  assign new_C309_ = new_C4067_;
  assign new_C308_ = new_C4000_;
  assign new_C307_ = new_C3933_;
  assign new_C306_ = new_C3866_;
  assign new_C305_ = new_C3799_;
  assign new_C304_ = new_C3732_;
  assign new_C303_ = ~new_C242_ & new_C256_;
  assign new_C302_ = new_C242_ & ~new_C256_;
  assign new_C301_ = new_C242_ & ~new_C256_;
  assign new_C300_ = ~new_C242_ & ~new_C256_;
  assign new_C299_ = new_C242_ & new_C256_;
  assign new_C298_ = new_C302_ | new_C303_;
  assign new_C297_ = ~new_C242_ & new_C256_;
  assign new_C296_ = new_C300_ | new_C301_;
  assign new_C295_ = ~new_C271_ & ~new_C291_;
  assign new_C294_ = new_C271_ & new_C291_;
  assign new_C293_ = ~new_C238_ | ~new_C263_;
  assign new_C292_ = new_C256_ & new_C293_;
  assign new_C291_ = new_C239_ | new_C240_;
  assign new_C290_ = new_C239_ | new_C256_;
  assign new_C289_ = ~new_C256_ & ~new_C292_;
  assign new_C288_ = new_C256_ | new_C293_;
  assign new_C287_ = new_C239_ & ~new_C240_;
  assign new_C286_ = ~new_C239_ & new_C240_;
  assign new_C285_ = new_C249_ | new_C282_;
  assign new_C284_ = ~new_C249_ & ~new_C283_;
  assign new_C283_ = new_C249_ & new_C282_;
  assign new_C282_ = ~new_C238_ | ~new_C263_;
  assign new_C281_ = ~new_C239_ & new_C249_;
  assign new_C280_ = new_C239_ & ~new_C249_;
  assign new_C279_ = new_C241_ & new_C278_;
  assign new_C278_ = new_C297_ | new_C296_;
  assign new_C277_ = ~new_C241_ & new_C276_;
  assign new_C276_ = new_C299_ | new_C298_;
  assign new_C275_ = new_C241_ | new_C274_;
  assign new_C274_ = new_C295_ | new_C294_;
  assign new_C273_ = ~new_C253_ & ~new_C263_;
  assign new_C272_ = new_C253_ & new_C263_;
  assign new_C271_ = ~new_C253_ | new_C263_;
  assign new_C270_ = new_C237_ & ~new_C238_;
  assign new_C269_ = ~new_C237_ & new_C238_;
  assign new_C268_ = new_C290_ & ~new_C291_;
  assign new_C267_ = ~new_C290_ & new_C291_;
  assign new_C266_ = ~new_C289_ | ~new_C288_;
  assign new_C265_ = new_C281_ | new_C280_;
  assign new_C264_ = new_C287_ | new_C286_;
  assign new_C263_ = new_C277_ | new_C279_;
  assign new_C262_ = ~new_C284_ | ~new_C285_;
  assign new_C261_ = new_C237_ & ~new_C238_;
  assign new_C260_ = new_C251_ & ~new_C263_;
  assign new_C259_ = ~new_C251_ & new_C263_;
  assign new_C258_ = ~new_C249_ & new_C275_;
  assign new_C257_ = new_C273_ | new_C272_;
  assign new_C256_ = new_C270_ | new_C269_;
  assign new_C255_ = new_C238_ | new_C271_;
  assign new_C254_ = new_C263_ & new_C266_;
  assign new_C253_ = new_C268_ | new_C267_;
  assign new_C252_ = new_C263_ & new_C262_;
  assign new_C251_ = new_C265_ & new_C264_;
  assign new_C250_ = new_C260_ | new_C259_;
  assign new_C249_ = new_C238_ | new_C261_;
  assign C248 = new_C249_ | new_C258_;
  assign C247 = new_C256_ & new_C257_;
  assign C246 = new_C256_ & new_C255_;
  assign C245 = new_C254_ | new_C253_;
  assign C244 = new_C252_ | new_C251_;
  assign C243 = new_C250_ & new_C249_;
  assign new_C242_ = new_C3665_;
  assign new_C241_ = new_C3598_;
  assign new_C240_ = new_C3531_;
  assign new_C239_ = new_C3464_;
  assign new_C238_ = new_C3397_;
  assign new_C237_ = new_C3330_;
  assign new_C236_ = ~new_C175_ & new_C189_;
  assign new_C235_ = new_C175_ & ~new_C189_;
  assign new_C234_ = new_C175_ & ~new_C189_;
  assign new_C233_ = ~new_C175_ & ~new_C189_;
  assign new_C232_ = new_C175_ & new_C189_;
  assign new_C231_ = new_C235_ | new_C236_;
  assign new_C230_ = ~new_C175_ & new_C189_;
  assign new_C229_ = new_C233_ | new_C234_;
  assign new_C228_ = ~new_C204_ & ~new_C224_;
  assign new_C227_ = new_C204_ & new_C224_;
  assign new_C226_ = ~new_C171_ | ~new_C196_;
  assign new_C225_ = new_C189_ & new_C226_;
  assign new_C224_ = new_C172_ | new_C173_;
  assign new_C223_ = new_C172_ | new_C189_;
  assign new_C222_ = ~new_C189_ & ~new_C225_;
  assign new_C221_ = new_C189_ | new_C226_;
  assign new_C220_ = new_C172_ & ~new_C173_;
  assign new_C219_ = ~new_C172_ & new_C173_;
  assign new_C218_ = new_C182_ | new_C215_;
  assign new_C217_ = ~new_C182_ & ~new_C216_;
  assign new_C216_ = new_C182_ & new_C215_;
  assign new_C215_ = ~new_C171_ | ~new_C196_;
  assign new_C214_ = ~new_C172_ & new_C182_;
  assign new_C213_ = new_C172_ & ~new_C182_;
  assign new_C212_ = new_C174_ & new_C211_;
  assign new_C211_ = new_C230_ | new_C229_;
  assign new_C210_ = ~new_C174_ & new_C209_;
  assign new_C209_ = new_C232_ | new_C231_;
  assign new_C208_ = new_C174_ | new_C207_;
  assign new_C207_ = new_C228_ | new_C227_;
  assign new_C206_ = ~new_C186_ & ~new_C196_;
  assign new_C205_ = new_C186_ & new_C196_;
  assign new_C204_ = ~new_C186_ | new_C196_;
  assign new_C203_ = new_C170_ & ~new_C171_;
  assign new_C202_ = ~new_C170_ & new_C171_;
  assign new_C201_ = new_C223_ & ~new_C224_;
  assign new_C200_ = ~new_C223_ & new_C224_;
  assign new_C199_ = ~new_C222_ | ~new_C221_;
  assign new_C198_ = new_C214_ | new_C213_;
  assign new_C197_ = new_C220_ | new_C219_;
  assign new_C196_ = new_C210_ | new_C212_;
  assign new_C195_ = ~new_C217_ | ~new_C218_;
  assign new_C194_ = new_C170_ & ~new_C171_;
  assign new_C193_ = new_C184_ & ~new_C196_;
  assign new_C192_ = ~new_C184_ & new_C196_;
  assign new_C191_ = ~new_C182_ & new_C208_;
  assign new_C190_ = new_C206_ | new_C205_;
  assign new_C189_ = new_C203_ | new_C202_;
  assign new_C188_ = new_C171_ | new_C204_;
  assign new_C187_ = new_C196_ & new_C199_;
  assign new_C186_ = new_C201_ | new_C200_;
  assign new_C185_ = new_C196_ & new_C195_;
  assign new_C184_ = new_C198_ & new_C197_;
  assign new_C183_ = new_C193_ | new_C192_;
  assign new_C182_ = new_C171_ | new_C194_;
  assign C181 = new_C182_ | new_C191_;
  assign C180 = new_C189_ & new_C190_;
  assign C179 = new_C189_ & new_C188_;
  assign C178 = new_C187_ | new_C186_;
  assign C177 = new_C185_ | new_C184_;
  assign C176 = new_C183_ & new_C182_;
  assign new_C175_ = new_C3263_;
  assign new_C174_ = new_C3196_;
  assign new_C173_ = new_C3129_;
  assign new_C172_ = new_C3062_;
  assign new_C171_ = new_C2995_;
  assign new_C170_ = new_C2928_;
  assign new_C169_ = ~new_C108_ & new_C122_;
  assign new_C168_ = new_C108_ & ~new_C122_;
  assign new_C167_ = new_C108_ & ~new_C122_;
  assign new_C166_ = ~new_C108_ & ~new_C122_;
  assign new_C165_ = new_C108_ & new_C122_;
  assign new_C164_ = new_C168_ | new_C169_;
  assign new_C163_ = ~new_C108_ & new_C122_;
  assign new_C162_ = new_C166_ | new_C167_;
  assign new_C161_ = ~new_C137_ & ~new_C157_;
  assign new_C160_ = new_C137_ & new_C157_;
  assign new_C159_ = ~new_C104_ | ~new_C129_;
  assign new_C158_ = new_C122_ & new_C159_;
  assign new_C157_ = new_C105_ | new_C106_;
  assign new_C156_ = new_C105_ | new_C122_;
  assign new_C155_ = ~new_C122_ & ~new_C158_;
  assign new_C154_ = new_C122_ | new_C159_;
  assign new_C153_ = new_C105_ & ~new_C106_;
  assign new_C152_ = ~new_C105_ & new_C106_;
  assign new_C151_ = new_C115_ | new_C148_;
  assign new_C150_ = ~new_C115_ & ~new_C149_;
  assign new_C149_ = new_C115_ & new_C148_;
  assign new_C148_ = ~new_C104_ | ~new_C129_;
  assign new_C147_ = ~new_C105_ & new_C115_;
  assign new_C146_ = new_C105_ & ~new_C115_;
  assign new_C145_ = new_C107_ & new_C144_;
  assign new_C144_ = new_C163_ | new_C162_;
  assign new_C143_ = ~new_C107_ & new_C142_;
  assign new_C142_ = new_C165_ | new_C164_;
  assign new_C141_ = new_C107_ | new_C140_;
  assign new_C140_ = new_C161_ | new_C160_;
  assign new_C139_ = ~new_C119_ & ~new_C129_;
  assign new_C138_ = new_C119_ & new_C129_;
  assign new_C137_ = ~new_C119_ | new_C129_;
  assign new_C136_ = new_C103_ & ~new_C104_;
  assign new_C135_ = ~new_C103_ & new_C104_;
  assign new_C134_ = new_C156_ & ~new_C157_;
  assign new_C133_ = ~new_C156_ & new_C157_;
  assign new_C132_ = ~new_C155_ | ~new_C154_;
  assign new_C131_ = new_C147_ | new_C146_;
  assign new_C130_ = new_C153_ | new_C152_;
  assign new_C129_ = new_C143_ | new_C145_;
  assign new_C128_ = ~new_C150_ | ~new_C151_;
  assign new_C127_ = new_C103_ & ~new_C104_;
  assign new_C126_ = new_C117_ & ~new_C129_;
  assign new_C125_ = ~new_C117_ & new_C129_;
  assign new_C124_ = ~new_C115_ & new_C141_;
  assign new_C123_ = new_C139_ | new_C138_;
  assign new_C122_ = new_C136_ | new_C135_;
  assign new_C121_ = new_C104_ | new_C137_;
  assign new_C120_ = new_C129_ & new_C132_;
  assign new_C119_ = new_C134_ | new_C133_;
  assign new_C118_ = new_C129_ & new_C128_;
  assign new_C117_ = new_C131_ & new_C130_;
  assign new_C116_ = new_C126_ | new_C125_;
  assign new_C115_ = new_C104_ | new_C127_;
  assign C114 = new_C115_ | new_C124_;
  assign C113 = new_C122_ & new_C123_;
  assign C112 = new_C122_ & new_C121_;
  assign C111 = new_C120_ | new_C119_;
  assign C110 = new_C118_ | new_C117_;
  assign C109 = new_C116_ & new_C115_;
  assign new_C108_ = new_C2861_;
  assign new_C107_ = new_C2794_;
  assign new_C106_ = new_C2727_;
  assign new_C105_ = new_C2660_;
  assign new_C104_ = new_C2593_;
  assign new_C103_ = new_C2521_;
  assign new_C102_ = ~new_C41_ & new_C55_;
  assign new_C101_ = new_C41_ & ~new_C55_;
  assign new_C100_ = new_C41_ & ~new_C55_;
  assign new_C99_ = ~new_C41_ & ~new_C55_;
  assign new_C98_ = new_C41_ & new_C55_;
  assign new_C97_ = new_C101_ | new_C102_;
  assign new_C96_ = ~new_C41_ & new_C55_;
  assign new_C95_ = new_C99_ | new_C100_;
  assign new_C94_ = ~new_C70_ & ~new_C90_;
  assign new_C93_ = new_C70_ & new_C90_;
  assign new_C92_ = ~new_C37_ | ~new_C62_;
  assign new_C91_ = new_C55_ & new_C92_;
  assign new_C90_ = new_C38_ | new_C39_;
  assign new_C89_ = new_C38_ | new_C55_;
  assign new_C88_ = ~new_C55_ & ~new_C91_;
  assign new_C87_ = new_C55_ | new_C92_;
  assign new_C86_ = new_C38_ & ~new_C39_;
  assign new_C85_ = ~new_C38_ & new_C39_;
  assign new_C84_ = new_C48_ | new_C81_;
  assign new_C83_ = ~new_C48_ & ~new_C82_;
  assign new_C82_ = new_C48_ & new_C81_;
  assign new_C81_ = ~new_C37_ | ~new_C62_;
  assign new_C80_ = ~new_C38_ & new_C48_;
  assign new_C79_ = new_C38_ & ~new_C48_;
  assign new_C78_ = new_C40_ & new_C77_;
  assign new_C77_ = new_C96_ | new_C95_;
  assign new_C76_ = ~new_C40_ & new_C75_;
  assign new_C75_ = new_C98_ | new_C97_;
  assign new_C74_ = new_C40_ | new_C73_;
  assign new_C73_ = new_C94_ | new_C93_;
  assign new_C72_ = ~new_C52_ & ~new_C62_;
  assign new_C71_ = new_C52_ & new_C62_;
  assign new_C70_ = ~new_C52_ | new_C62_;
  assign new_C69_ = new_C36_ & ~new_C37_;
  assign new_C68_ = ~new_C36_ & new_C37_;
  assign new_C67_ = new_C89_ & ~new_C90_;
  assign new_C66_ = ~new_C89_ & new_C90_;
  assign new_C65_ = ~new_C88_ | ~new_C87_;
  assign new_C64_ = new_C80_ | new_C79_;
  assign new_C63_ = new_C86_ | new_C85_;
  assign new_C62_ = new_C76_ | new_C78_;
  assign new_C61_ = ~new_C83_ | ~new_C84_;
  assign new_C60_ = new_C36_ & ~new_C37_;
  assign new_C59_ = new_C50_ & ~new_C62_;
  assign new_C58_ = ~new_C50_ & new_C62_;
  assign new_C57_ = ~new_C48_ & new_C74_;
  assign new_C56_ = new_C72_ | new_C71_;
  assign new_C55_ = new_C69_ | new_C68_;
  assign new_C54_ = new_C37_ | new_C70_;
  assign new_C53_ = new_C62_ & new_C65_;
  assign new_C52_ = new_C67_ | new_C66_;
  assign new_C51_ = new_C62_ & new_C61_;
  assign new_C50_ = new_C64_ & new_C63_;
  assign new_C49_ = new_C59_ | new_C58_;
  assign new_C48_ = new_C37_ | new_C60_;
  assign C47 = new_C48_ | new_C57_;
  assign C46 = new_C55_ & new_C56_;
  assign C45 = new_C55_ & new_C54_;
  assign C44 = new_C53_ | new_C52_;
  assign C43 = new_C51_ | new_C50_;
  assign C42 = new_C49_ & new_C48_;
  assign new_C41_ = new_D6931_;
  assign new_C40_ = new_D6864_;
  assign new_C39_ = new_D6797_;
  assign new_C38_ = new_D6730_;
  assign new_C37_ = new_D6663_;
  assign new_C36_ = new_D6596_;
  assign new_C35_ = ~new_B9973_ & new_B9987_;
  assign new_C34_ = new_B9973_ & ~new_B9987_;
  assign new_C33_ = new_B9973_ & ~new_B9987_;
  assign new_C32_ = ~new_B9973_ & ~new_B9987_;
  assign new_C31_ = new_B9973_ & new_B9987_;
  assign new_C30_ = new_C34_ | new_C35_;
  assign new_C29_ = ~new_B9973_ & new_B9987_;
  assign new_C28_ = new_C32_ | new_C33_;
  assign new_C27_ = ~new_C3_ & ~new_C23_;
  assign new_C26_ = new_C3_ & new_C23_;
  assign new_C25_ = ~new_B9969_ | ~new_B9994_;
  assign new_C24_ = new_B9987_ & new_C25_;
  assign new_C23_ = new_B9970_ | new_B9971_;
  assign new_C22_ = new_B9970_ | new_B9987_;
  assign new_C21_ = ~new_B9987_ & ~new_C24_;
  assign new_C20_ = new_B9987_ | new_C25_;
  assign new_C19_ = new_B9970_ & ~new_B9971_;
  assign new_C18_ = ~new_B9970_ & new_B9971_;
  assign new_C17_ = new_B9980_ | new_C14_;
  assign new_C16_ = ~new_B9980_ & ~new_C15_;
  assign new_C15_ = new_B9980_ & new_C14_;
  assign new_C14_ = ~new_B9969_ | ~new_B9994_;
  assign new_C13_ = ~new_B9970_ & new_B9980_;
  assign new_C12_ = new_B9970_ & ~new_B9980_;
  assign new_C11_ = new_B9972_ & new_C10_;
  assign new_C10_ = new_C29_ | new_C28_;
  assign new_C9_ = ~new_B9972_ & new_C8_;
  assign new_C8_ = new_C31_ | new_C30_;
  assign new_C7_ = new_B9972_ | new_C6_;
  assign new_C6_ = new_C27_ | new_C26_;
  assign new_C5_ = ~new_B9984_ & ~new_B9994_;
  assign new_C4_ = new_B9984_ & new_B9994_;
  assign new_C3_ = ~new_B9984_ | new_B9994_;
  assign new_C2_ = new_B9968_ & ~new_B9969_;
  assign new_C1_ = ~new_B9968_ & new_B9969_;
  assign new_B9999_ = new_C22_ & ~new_C23_;
  assign new_B9998_ = ~new_C22_ & new_C23_;
  assign new_B9997_ = ~new_C21_ | ~new_C20_;
  assign new_B9996_ = new_C13_ | new_C12_;
  assign new_B9995_ = new_C19_ | new_C18_;
  assign new_B9994_ = new_C9_ | new_C11_;
  assign new_B9993_ = ~new_C16_ | ~new_C17_;
  assign new_B9992_ = new_B9968_ & ~new_B9969_;
  assign new_B9991_ = new_B9982_ & ~new_B9994_;
  assign new_B9990_ = ~new_B9982_ & new_B9994_;
  assign new_B9989_ = ~new_B9980_ & new_C7_;
  assign new_B9988_ = new_C5_ | new_C4_;
  assign new_B9987_ = new_C2_ | new_C1_;
  assign new_B9986_ = new_B9969_ | new_C3_;
  assign new_B9985_ = new_B9994_ & new_B9997_;
  assign new_B9984_ = new_B9999_ | new_B9998_;
  assign new_B9983_ = new_B9994_ & new_B9993_;
  assign new_B9982_ = new_B9996_ & new_B9995_;
  assign new_B9981_ = new_B9991_ | new_B9990_;
  assign new_B9980_ = new_B9969_ | new_B9992_;
  assign B9979 = new_B9980_ | new_B9989_;
  assign B9978 = new_B9987_ & new_B9988_;
  assign B9977 = new_B9987_ & new_B9986_;
  assign B9976 = new_B9985_ | new_B9984_;
  assign B9975 = new_B9983_ | new_B9982_;
  assign B9974 = new_B9981_ & new_B9980_;
  assign new_B9973_ = new_D6529_;
  assign new_B9972_ = new_D6462_;
  assign new_B9971_ = new_D6395_;
  assign new_B9970_ = new_D6328_;
  assign new_B9969_ = new_D6261_;
  assign new_B9968_ = new_D6194_;
  assign new_B9967_ = ~new_B9906_ & new_B9920_;
  assign new_B9966_ = new_B9906_ & ~new_B9920_;
  assign new_B9965_ = new_B9906_ & ~new_B9920_;
  assign new_B9964_ = ~new_B9906_ & ~new_B9920_;
  assign new_B9963_ = new_B9906_ & new_B9920_;
  assign new_B9962_ = new_B9966_ | new_B9967_;
  assign new_B9961_ = ~new_B9906_ & new_B9920_;
  assign new_B9960_ = new_B9964_ | new_B9965_;
  assign new_B9959_ = ~new_B9935_ & ~new_B9955_;
  assign new_B9958_ = new_B9935_ & new_B9955_;
  assign new_B9957_ = ~new_B9902_ | ~new_B9927_;
  assign new_B9956_ = new_B9920_ & new_B9957_;
  assign new_B9955_ = new_B9903_ | new_B9904_;
  assign new_B9954_ = new_B9903_ | new_B9920_;
  assign new_B9953_ = ~new_B9920_ & ~new_B9956_;
  assign new_B9952_ = new_B9920_ | new_B9957_;
  assign new_B9951_ = new_B9903_ & ~new_B9904_;
  assign new_B9950_ = ~new_B9903_ & new_B9904_;
  assign new_B9949_ = new_B9913_ | new_B9946_;
  assign new_B9948_ = ~new_B9913_ & ~new_B9947_;
  assign new_B9947_ = new_B9913_ & new_B9946_;
  assign new_B9946_ = ~new_B9902_ | ~new_B9927_;
  assign new_B9945_ = ~new_B9903_ & new_B9913_;
  assign new_B9944_ = new_B9903_ & ~new_B9913_;
  assign new_B9943_ = new_B9905_ & new_B9942_;
  assign new_B9942_ = new_B9961_ | new_B9960_;
  assign new_B9941_ = ~new_B9905_ & new_B9940_;
  assign new_B9940_ = new_B9963_ | new_B9962_;
  assign new_B9939_ = new_B9905_ | new_B9938_;
  assign new_B9938_ = new_B9959_ | new_B9958_;
  assign new_B9937_ = ~new_B9917_ & ~new_B9927_;
  assign new_B9936_ = new_B9917_ & new_B9927_;
  assign new_B9935_ = ~new_B9917_ | new_B9927_;
  assign new_B9934_ = new_B9901_ & ~new_B9902_;
  assign new_B9933_ = ~new_B9901_ & new_B9902_;
  assign new_B9932_ = new_B9954_ & ~new_B9955_;
  assign new_B9931_ = ~new_B9954_ & new_B9955_;
  assign new_B9930_ = ~new_B9953_ | ~new_B9952_;
  assign new_B9929_ = new_B9945_ | new_B9944_;
  assign new_B9928_ = new_B9951_ | new_B9950_;
  assign new_B9927_ = new_B9941_ | new_B9943_;
  assign new_B9926_ = ~new_B9948_ | ~new_B9949_;
  assign new_B9925_ = new_B9901_ & ~new_B9902_;
  assign new_B9924_ = new_B9915_ & ~new_B9927_;
  assign new_B9923_ = ~new_B9915_ & new_B9927_;
  assign new_B9922_ = ~new_B9913_ & new_B9939_;
  assign new_B9921_ = new_B9937_ | new_B9936_;
  assign new_B9920_ = new_B9934_ | new_B9933_;
  assign new_B9919_ = new_B9902_ | new_B9935_;
  assign new_B9918_ = new_B9927_ & new_B9930_;
  assign new_B9917_ = new_B9932_ | new_B9931_;
  assign new_B9916_ = new_B9927_ & new_B9926_;
  assign new_B9915_ = new_B9929_ & new_B9928_;
  assign new_B9914_ = new_B9924_ | new_B9923_;
  assign new_B9913_ = new_B9902_ | new_B9925_;
  assign B9912 = new_B9913_ | new_B9922_;
  assign B9911 = new_B9920_ & new_B9921_;
  assign B9910 = new_B9920_ & new_B9919_;
  assign B9909 = new_B9918_ | new_B9917_;
  assign B9908 = new_B9916_ | new_B9915_;
  assign B9907 = new_B9914_ & new_B9913_;
  assign new_B9906_ = new_D6127_;
  assign new_B9905_ = new_D6060_;
  assign new_B9904_ = new_D5993_;
  assign new_B9903_ = new_D5926_;
  assign new_B9902_ = new_D5859_;
  assign new_B9901_ = new_D5792_;
  assign new_B9900_ = ~new_B9839_ & new_B9853_;
  assign new_B9899_ = new_B9839_ & ~new_B9853_;
  assign new_B9898_ = new_B9839_ & ~new_B9853_;
  assign new_B9897_ = ~new_B9839_ & ~new_B9853_;
  assign new_B9896_ = new_B9839_ & new_B9853_;
  assign new_B9895_ = new_B9899_ | new_B9900_;
  assign new_B9894_ = ~new_B9839_ & new_B9853_;
  assign new_B9893_ = new_B9897_ | new_B9898_;
  assign new_B9892_ = ~new_B9868_ & ~new_B9888_;
  assign new_B9891_ = new_B9868_ & new_B9888_;
  assign new_B9890_ = ~new_B9835_ | ~new_B9860_;
  assign new_B9889_ = new_B9853_ & new_B9890_;
  assign new_B9888_ = new_B9836_ | new_B9837_;
  assign new_B9887_ = new_B9836_ | new_B9853_;
  assign new_B9886_ = ~new_B9853_ & ~new_B9889_;
  assign new_B9885_ = new_B9853_ | new_B9890_;
  assign new_B9884_ = new_B9836_ & ~new_B9837_;
  assign new_B9883_ = ~new_B9836_ & new_B9837_;
  assign new_B9882_ = new_B9846_ | new_B9879_;
  assign new_B9881_ = ~new_B9846_ & ~new_B9880_;
  assign new_B9880_ = new_B9846_ & new_B9879_;
  assign new_B9879_ = ~new_B9835_ | ~new_B9860_;
  assign new_B9878_ = ~new_B9836_ & new_B9846_;
  assign new_B9877_ = new_B9836_ & ~new_B9846_;
  assign new_B9876_ = new_B9838_ & new_B9875_;
  assign new_B9875_ = new_B9894_ | new_B9893_;
  assign new_B9874_ = ~new_B9838_ & new_B9873_;
  assign new_B9873_ = new_B9896_ | new_B9895_;
  assign new_B9872_ = new_B9838_ | new_B9871_;
  assign new_B9871_ = new_B9892_ | new_B9891_;
  assign new_B9870_ = ~new_B9850_ & ~new_B9860_;
  assign new_B9869_ = new_B9850_ & new_B9860_;
  assign new_B9868_ = ~new_B9850_ | new_B9860_;
  assign new_B9867_ = new_B9834_ & ~new_B9835_;
  assign new_B9866_ = ~new_B9834_ & new_B9835_;
  assign new_B9865_ = new_B9887_ & ~new_B9888_;
  assign new_B9864_ = ~new_B9887_ & new_B9888_;
  assign new_B9863_ = ~new_B9886_ | ~new_B9885_;
  assign new_B9862_ = new_B9878_ | new_B9877_;
  assign new_B9861_ = new_B9884_ | new_B9883_;
  assign new_B9860_ = new_B9874_ | new_B9876_;
  assign new_B9859_ = ~new_B9881_ | ~new_B9882_;
  assign new_B9858_ = new_B9834_ & ~new_B9835_;
  assign new_B9857_ = new_B9848_ & ~new_B9860_;
  assign new_B9856_ = ~new_B9848_ & new_B9860_;
  assign new_B9855_ = ~new_B9846_ & new_B9872_;
  assign new_B9854_ = new_B9870_ | new_B9869_;
  assign new_B9853_ = new_B9867_ | new_B9866_;
  assign new_B9852_ = new_B9835_ | new_B9868_;
  assign new_B9851_ = new_B9860_ & new_B9863_;
  assign new_B9850_ = new_B9865_ | new_B9864_;
  assign new_B9849_ = new_B9860_ & new_B9859_;
  assign new_B9848_ = new_B9862_ & new_B9861_;
  assign new_B9847_ = new_B9857_ | new_B9856_;
  assign new_B9846_ = new_B9835_ | new_B9858_;
  assign B9845 = new_B9846_ | new_B9855_;
  assign B9844 = new_B9853_ & new_B9854_;
  assign B9843 = new_B9853_ & new_B9852_;
  assign B9842 = new_B9851_ | new_B9850_;
  assign B9841 = new_B9849_ | new_B9848_;
  assign B9840 = new_B9847_ & new_B9846_;
  assign new_B9839_ = new_D5725_;
  assign new_B9838_ = new_D5658_;
  assign new_B9837_ = new_D5591_;
  assign new_B9836_ = new_D5524_;
  assign new_B9835_ = new_D5457_;
  assign new_B9834_ = new_D5390_;
  assign new_B9833_ = ~new_B9772_ & new_B9786_;
  assign new_B9832_ = new_B9772_ & ~new_B9786_;
  assign new_B9831_ = new_B9772_ & ~new_B9786_;
  assign new_B9830_ = ~new_B9772_ & ~new_B9786_;
  assign new_B9829_ = new_B9772_ & new_B9786_;
  assign new_B9828_ = new_B9832_ | new_B9833_;
  assign new_B9827_ = ~new_B9772_ & new_B9786_;
  assign new_B9826_ = new_B9830_ | new_B9831_;
  assign new_B9825_ = ~new_B9801_ & ~new_B9821_;
  assign new_B9824_ = new_B9801_ & new_B9821_;
  assign new_B9823_ = ~new_B9768_ | ~new_B9793_;
  assign new_B9822_ = new_B9786_ & new_B9823_;
  assign new_B9821_ = new_B9769_ | new_B9770_;
  assign new_B9820_ = new_B9769_ | new_B9786_;
  assign new_B9819_ = ~new_B9786_ & ~new_B9822_;
  assign new_B9818_ = new_B9786_ | new_B9823_;
  assign new_B9817_ = new_B9769_ & ~new_B9770_;
  assign new_B9816_ = ~new_B9769_ & new_B9770_;
  assign new_B9815_ = new_B9779_ | new_B9812_;
  assign new_B9814_ = ~new_B9779_ & ~new_B9813_;
  assign new_B9813_ = new_B9779_ & new_B9812_;
  assign new_B9812_ = ~new_B9768_ | ~new_B9793_;
  assign new_B9811_ = ~new_B9769_ & new_B9779_;
  assign new_B9810_ = new_B9769_ & ~new_B9779_;
  assign new_B9809_ = new_B9771_ & new_B9808_;
  assign new_B9808_ = new_B9827_ | new_B9826_;
  assign new_B9807_ = ~new_B9771_ & new_B9806_;
  assign new_B9806_ = new_B9829_ | new_B9828_;
  assign new_B9805_ = new_B9771_ | new_B9804_;
  assign new_B9804_ = new_B9825_ | new_B9824_;
  assign new_B9803_ = ~new_B9783_ & ~new_B9793_;
  assign new_B9802_ = new_B9783_ & new_B9793_;
  assign new_B9801_ = ~new_B9783_ | new_B9793_;
  assign new_B9800_ = new_B9767_ & ~new_B9768_;
  assign new_B9799_ = ~new_B9767_ & new_B9768_;
  assign new_B9798_ = new_B9820_ & ~new_B9821_;
  assign new_B9797_ = ~new_B9820_ & new_B9821_;
  assign new_B9796_ = ~new_B9819_ | ~new_B9818_;
  assign new_B9795_ = new_B9811_ | new_B9810_;
  assign new_B9794_ = new_B9817_ | new_B9816_;
  assign new_B9793_ = new_B9807_ | new_B9809_;
  assign new_B9792_ = ~new_B9814_ | ~new_B9815_;
  assign new_B9791_ = new_B9767_ & ~new_B9768_;
  assign new_B9790_ = new_B9781_ & ~new_B9793_;
  assign new_B9789_ = ~new_B9781_ & new_B9793_;
  assign new_B9788_ = ~new_B9779_ & new_B9805_;
  assign new_B9787_ = new_B9803_ | new_B9802_;
  assign new_B9786_ = new_B9800_ | new_B9799_;
  assign new_B9785_ = new_B9768_ | new_B9801_;
  assign new_B9784_ = new_B9793_ & new_B9796_;
  assign new_B9783_ = new_B9798_ | new_B9797_;
  assign new_B9782_ = new_B9793_ & new_B9792_;
  assign new_B9781_ = new_B9795_ & new_B9794_;
  assign new_B9780_ = new_B9790_ | new_B9789_;
  assign new_B9779_ = new_B9768_ | new_B9791_;
  assign B9778 = new_B9779_ | new_B9788_;
  assign B9777 = new_B9786_ & new_B9787_;
  assign B9776 = new_B9786_ & new_B9785_;
  assign B9775 = new_B9784_ | new_B9783_;
  assign B9774 = new_B9782_ | new_B9781_;
  assign B9773 = new_B9780_ & new_B9779_;
  assign new_B9772_ = new_D5323_;
  assign new_B9771_ = new_D5256_;
  assign new_B9770_ = new_D5189_;
  assign new_B9769_ = new_D5122_;
  assign new_B9768_ = new_D5055_;
  assign new_B9767_ = new_D4988_;
  assign new_B9766_ = ~new_B9705_ & new_B9719_;
  assign new_B9765_ = new_B9705_ & ~new_B9719_;
  assign new_B9764_ = new_B9705_ & ~new_B9719_;
  assign new_B9763_ = ~new_B9705_ & ~new_B9719_;
  assign new_B9762_ = new_B9705_ & new_B9719_;
  assign new_B9761_ = new_B9765_ | new_B9766_;
  assign new_B9760_ = ~new_B9705_ & new_B9719_;
  assign new_B9759_ = new_B9763_ | new_B9764_;
  assign new_B9758_ = ~new_B9734_ & ~new_B9754_;
  assign new_B9757_ = new_B9734_ & new_B9754_;
  assign new_B9756_ = ~new_B9701_ | ~new_B9726_;
  assign new_B9755_ = new_B9719_ & new_B9756_;
  assign new_B9754_ = new_B9702_ | new_B9703_;
  assign new_B9753_ = new_B9702_ | new_B9719_;
  assign new_B9752_ = ~new_B9719_ & ~new_B9755_;
  assign new_B9751_ = new_B9719_ | new_B9756_;
  assign new_B9750_ = new_B9702_ & ~new_B9703_;
  assign new_B9749_ = ~new_B9702_ & new_B9703_;
  assign new_B9748_ = new_B9712_ | new_B9745_;
  assign new_B9747_ = ~new_B9712_ & ~new_B9746_;
  assign new_B9746_ = new_B9712_ & new_B9745_;
  assign new_B9745_ = ~new_B9701_ | ~new_B9726_;
  assign new_B9744_ = ~new_B9702_ & new_B9712_;
  assign new_B9743_ = new_B9702_ & ~new_B9712_;
  assign new_B9742_ = new_B9704_ & new_B9741_;
  assign new_B9741_ = new_B9760_ | new_B9759_;
  assign new_B9740_ = ~new_B9704_ & new_B9739_;
  assign new_B9739_ = new_B9762_ | new_B9761_;
  assign new_B9738_ = new_B9704_ | new_B9737_;
  assign new_B9737_ = new_B9758_ | new_B9757_;
  assign new_B9736_ = ~new_B9716_ & ~new_B9726_;
  assign new_B9735_ = new_B9716_ & new_B9726_;
  assign new_B9734_ = ~new_B9716_ | new_B9726_;
  assign new_B9733_ = new_B9700_ & ~new_B9701_;
  assign new_B9732_ = ~new_B9700_ & new_B9701_;
  assign new_B9731_ = new_B9753_ & ~new_B9754_;
  assign new_B9730_ = ~new_B9753_ & new_B9754_;
  assign new_B9729_ = ~new_B9752_ | ~new_B9751_;
  assign new_B9728_ = new_B9744_ | new_B9743_;
  assign new_B9727_ = new_B9750_ | new_B9749_;
  assign new_B9726_ = new_B9740_ | new_B9742_;
  assign new_B9725_ = ~new_B9747_ | ~new_B9748_;
  assign new_B9724_ = new_B9700_ & ~new_B9701_;
  assign new_B9723_ = new_B9714_ & ~new_B9726_;
  assign new_B9722_ = ~new_B9714_ & new_B9726_;
  assign new_B9721_ = ~new_B9712_ & new_B9738_;
  assign new_B9720_ = new_B9736_ | new_B9735_;
  assign new_B9719_ = new_B9733_ | new_B9732_;
  assign new_B9718_ = new_B9701_ | new_B9734_;
  assign new_B9717_ = new_B9726_ & new_B9729_;
  assign new_B9716_ = new_B9731_ | new_B9730_;
  assign new_B9715_ = new_B9726_ & new_B9725_;
  assign new_B9714_ = new_B9728_ & new_B9727_;
  assign new_B9713_ = new_B9723_ | new_B9722_;
  assign new_B9712_ = new_B9701_ | new_B9724_;
  assign B9711 = new_B9712_ | new_B9721_;
  assign B9710 = new_B9719_ & new_B9720_;
  assign B9709 = new_B9719_ & new_B9718_;
  assign B9708 = new_B9717_ | new_B9716_;
  assign B9707 = new_B9715_ | new_B9714_;
  assign B9706 = new_B9713_ & new_B9712_;
  assign new_B9705_ = new_D4921_;
  assign new_B9704_ = new_D4854_;
  assign new_B9703_ = new_D4787_;
  assign new_B9702_ = new_D4720_;
  assign new_B9701_ = new_D4653_;
  assign new_B9700_ = new_D4586_;
  assign new_B9699_ = ~new_B9638_ & new_B9652_;
  assign new_B9698_ = new_B9638_ & ~new_B9652_;
  assign new_B9697_ = new_B9638_ & ~new_B9652_;
  assign new_B9696_ = ~new_B9638_ & ~new_B9652_;
  assign new_B9695_ = new_B9638_ & new_B9652_;
  assign new_B9694_ = new_B9698_ | new_B9699_;
  assign new_B9693_ = ~new_B9638_ & new_B9652_;
  assign new_B9692_ = new_B9696_ | new_B9697_;
  assign new_B9691_ = ~new_B9667_ & ~new_B9687_;
  assign new_B9690_ = new_B9667_ & new_B9687_;
  assign new_B9689_ = ~new_B9634_ | ~new_B9659_;
  assign new_B9688_ = new_B9652_ & new_B9689_;
  assign new_B9687_ = new_B9635_ | new_B9636_;
  assign new_B9686_ = new_B9635_ | new_B9652_;
  assign new_B9685_ = ~new_B9652_ & ~new_B9688_;
  assign new_B9684_ = new_B9652_ | new_B9689_;
  assign new_B9683_ = new_B9635_ & ~new_B9636_;
  assign new_B9682_ = ~new_B9635_ & new_B9636_;
  assign new_B9681_ = new_B9645_ | new_B9678_;
  assign new_B9680_ = ~new_B9645_ & ~new_B9679_;
  assign new_B9679_ = new_B9645_ & new_B9678_;
  assign new_B9678_ = ~new_B9634_ | ~new_B9659_;
  assign new_B9677_ = ~new_B9635_ & new_B9645_;
  assign new_B9676_ = new_B9635_ & ~new_B9645_;
  assign new_B9675_ = new_B9637_ & new_B9674_;
  assign new_B9674_ = new_B9693_ | new_B9692_;
  assign new_B9673_ = ~new_B9637_ & new_B9672_;
  assign new_B9672_ = new_B9695_ | new_B9694_;
  assign new_B9671_ = new_B9637_ | new_B9670_;
  assign new_B9670_ = new_B9691_ | new_B9690_;
  assign new_B9669_ = ~new_B9649_ & ~new_B9659_;
  assign new_B9668_ = new_B9649_ & new_B9659_;
  assign new_B9667_ = ~new_B9649_ | new_B9659_;
  assign new_B9666_ = new_B9633_ & ~new_B9634_;
  assign new_B9665_ = ~new_B9633_ & new_B9634_;
  assign new_B9664_ = new_B9686_ & ~new_B9687_;
  assign new_B9663_ = ~new_B9686_ & new_B9687_;
  assign new_B9662_ = ~new_B9685_ | ~new_B9684_;
  assign new_B9661_ = new_B9677_ | new_B9676_;
  assign new_B9660_ = new_B9683_ | new_B9682_;
  assign new_B9659_ = new_B9673_ | new_B9675_;
  assign new_B9658_ = ~new_B9680_ | ~new_B9681_;
  assign new_B9657_ = new_B9633_ & ~new_B9634_;
  assign new_B9656_ = new_B9647_ & ~new_B9659_;
  assign new_B9655_ = ~new_B9647_ & new_B9659_;
  assign new_B9654_ = ~new_B9645_ & new_B9671_;
  assign new_B9653_ = new_B9669_ | new_B9668_;
  assign new_B9652_ = new_B9666_ | new_B9665_;
  assign new_B9651_ = new_B9634_ | new_B9667_;
  assign new_B9650_ = new_B9659_ & new_B9662_;
  assign new_B9649_ = new_B9664_ | new_B9663_;
  assign new_B9648_ = new_B9659_ & new_B9658_;
  assign new_B9647_ = new_B9661_ & new_B9660_;
  assign new_B9646_ = new_B9656_ | new_B9655_;
  assign new_B9645_ = new_B9634_ | new_B9657_;
  assign B9644 = new_B9645_ | new_B9654_;
  assign B9643 = new_B9652_ & new_B9653_;
  assign B9642 = new_B9652_ & new_B9651_;
  assign B9641 = new_B9650_ | new_B9649_;
  assign B9640 = new_B9648_ | new_B9647_;
  assign B9639 = new_B9646_ & new_B9645_;
  assign new_B9638_ = new_D4519_;
  assign new_B9637_ = new_D4452_;
  assign new_B9636_ = new_D4385_;
  assign new_B9635_ = new_D4318_;
  assign new_B9634_ = new_D4251_;
  assign new_B9633_ = new_D4184_;
  assign new_B9632_ = ~new_B9571_ & new_B9585_;
  assign new_B9631_ = new_B9571_ & ~new_B9585_;
  assign new_B9630_ = new_B9571_ & ~new_B9585_;
  assign new_B9629_ = ~new_B9571_ & ~new_B9585_;
  assign new_B9628_ = new_B9571_ & new_B9585_;
  assign new_B9627_ = new_B9631_ | new_B9632_;
  assign new_B9626_ = ~new_B9571_ & new_B9585_;
  assign new_B9625_ = new_B9629_ | new_B9630_;
  assign new_B9624_ = ~new_B9600_ & ~new_B9620_;
  assign new_B9623_ = new_B9600_ & new_B9620_;
  assign new_B9622_ = ~new_B9567_ | ~new_B9592_;
  assign new_B9621_ = new_B9585_ & new_B9622_;
  assign new_B9620_ = new_B9568_ | new_B9569_;
  assign new_B9619_ = new_B9568_ | new_B9585_;
  assign new_B9618_ = ~new_B9585_ & ~new_B9621_;
  assign new_B9617_ = new_B9585_ | new_B9622_;
  assign new_B9616_ = new_B9568_ & ~new_B9569_;
  assign new_B9615_ = ~new_B9568_ & new_B9569_;
  assign new_B9614_ = new_B9578_ | new_B9611_;
  assign new_B9613_ = ~new_B9578_ & ~new_B9612_;
  assign new_B9612_ = new_B9578_ & new_B9611_;
  assign new_B9611_ = ~new_B9567_ | ~new_B9592_;
  assign new_B9610_ = ~new_B9568_ & new_B9578_;
  assign new_B9609_ = new_B9568_ & ~new_B9578_;
  assign new_B9608_ = new_B9570_ & new_B9607_;
  assign new_B9607_ = new_B9626_ | new_B9625_;
  assign new_B9606_ = ~new_B9570_ & new_B9605_;
  assign new_B9605_ = new_B9628_ | new_B9627_;
  assign new_B9604_ = new_B9570_ | new_B9603_;
  assign new_B9603_ = new_B9624_ | new_B9623_;
  assign new_B9602_ = ~new_B9582_ & ~new_B9592_;
  assign new_B9601_ = new_B9582_ & new_B9592_;
  assign new_B9600_ = ~new_B9582_ | new_B9592_;
  assign new_B9599_ = new_B9566_ & ~new_B9567_;
  assign new_B9598_ = ~new_B9566_ & new_B9567_;
  assign new_B9597_ = new_B9619_ & ~new_B9620_;
  assign new_B9596_ = ~new_B9619_ & new_B9620_;
  assign new_B9595_ = ~new_B9618_ | ~new_B9617_;
  assign new_B9594_ = new_B9610_ | new_B9609_;
  assign new_B9593_ = new_B9616_ | new_B9615_;
  assign new_B9592_ = new_B9606_ | new_B9608_;
  assign new_B9591_ = ~new_B9613_ | ~new_B9614_;
  assign new_B9590_ = new_B9566_ & ~new_B9567_;
  assign new_B9589_ = new_B9580_ & ~new_B9592_;
  assign new_B9588_ = ~new_B9580_ & new_B9592_;
  assign new_B9587_ = ~new_B9578_ & new_B9604_;
  assign new_B9586_ = new_B9602_ | new_B9601_;
  assign new_B9585_ = new_B9599_ | new_B9598_;
  assign new_B9584_ = new_B9567_ | new_B9600_;
  assign new_B9583_ = new_B9592_ & new_B9595_;
  assign new_B9582_ = new_B9597_ | new_B9596_;
  assign new_B9581_ = new_B9592_ & new_B9591_;
  assign new_B9580_ = new_B9594_ & new_B9593_;
  assign new_B9579_ = new_B9589_ | new_B9588_;
  assign new_B9578_ = new_B9567_ | new_B9590_;
  assign B9577 = new_B9578_ | new_B9587_;
  assign B9576 = new_B9585_ & new_B9586_;
  assign B9575 = new_B9585_ & new_B9584_;
  assign B9574 = new_B9583_ | new_B9582_;
  assign B9573 = new_B9581_ | new_B9580_;
  assign B9572 = new_B9579_ & new_B9578_;
  assign new_B9571_ = new_D4117_;
  assign new_B9570_ = new_D4050_;
  assign new_B9569_ = new_D3983_;
  assign new_B9568_ = new_D3916_;
  assign new_B9567_ = new_D3849_;
  assign new_B9566_ = new_D3782_;
  assign new_B9565_ = ~new_B9504_ & new_B9518_;
  assign new_B9564_ = new_B9504_ & ~new_B9518_;
  assign new_B9563_ = new_B9504_ & ~new_B9518_;
  assign new_B9562_ = ~new_B9504_ & ~new_B9518_;
  assign new_B9561_ = new_B9504_ & new_B9518_;
  assign new_B9560_ = new_B9564_ | new_B9565_;
  assign new_B9559_ = ~new_B9504_ & new_B9518_;
  assign new_B9558_ = new_B9562_ | new_B9563_;
  assign new_B9557_ = ~new_B9533_ & ~new_B9553_;
  assign new_B9556_ = new_B9533_ & new_B9553_;
  assign new_B9555_ = ~new_B9500_ | ~new_B9525_;
  assign new_B9554_ = new_B9518_ & new_B9555_;
  assign new_B9553_ = new_B9501_ | new_B9502_;
  assign new_B9552_ = new_B9501_ | new_B9518_;
  assign new_B9551_ = ~new_B9518_ & ~new_B9554_;
  assign new_B9550_ = new_B9518_ | new_B9555_;
  assign new_B9549_ = new_B9501_ & ~new_B9502_;
  assign new_B9548_ = ~new_B9501_ & new_B9502_;
  assign new_B9547_ = new_B9511_ | new_B9544_;
  assign new_B9546_ = ~new_B9511_ & ~new_B9545_;
  assign new_B9545_ = new_B9511_ & new_B9544_;
  assign new_B9544_ = ~new_B9500_ | ~new_B9525_;
  assign new_B9543_ = ~new_B9501_ & new_B9511_;
  assign new_B9542_ = new_B9501_ & ~new_B9511_;
  assign new_B9541_ = new_B9503_ & new_B9540_;
  assign new_B9540_ = new_B9559_ | new_B9558_;
  assign new_B9539_ = ~new_B9503_ & new_B9538_;
  assign new_B9538_ = new_B9561_ | new_B9560_;
  assign new_B9537_ = new_B9503_ | new_B9536_;
  assign new_B9536_ = new_B9557_ | new_B9556_;
  assign new_B9535_ = ~new_B9515_ & ~new_B9525_;
  assign new_B9534_ = new_B9515_ & new_B9525_;
  assign new_B9533_ = ~new_B9515_ | new_B9525_;
  assign new_B9532_ = new_B9499_ & ~new_B9500_;
  assign new_B9531_ = ~new_B9499_ & new_B9500_;
  assign new_B9530_ = new_B9552_ & ~new_B9553_;
  assign new_B9529_ = ~new_B9552_ & new_B9553_;
  assign new_B9528_ = ~new_B9551_ | ~new_B9550_;
  assign new_B9527_ = new_B9543_ | new_B9542_;
  assign new_B9526_ = new_B9549_ | new_B9548_;
  assign new_B9525_ = new_B9539_ | new_B9541_;
  assign new_B9524_ = ~new_B9546_ | ~new_B9547_;
  assign new_B9523_ = new_B9499_ & ~new_B9500_;
  assign new_B9522_ = new_B9513_ & ~new_B9525_;
  assign new_B9521_ = ~new_B9513_ & new_B9525_;
  assign new_B9520_ = ~new_B9511_ & new_B9537_;
  assign new_B9519_ = new_B9535_ | new_B9534_;
  assign new_B9518_ = new_B9532_ | new_B9531_;
  assign new_B9517_ = new_B9500_ | new_B9533_;
  assign new_B9516_ = new_B9525_ & new_B9528_;
  assign new_B9515_ = new_B9530_ | new_B9529_;
  assign new_B9514_ = new_B9525_ & new_B9524_;
  assign new_B9513_ = new_B9527_ & new_B9526_;
  assign new_B9512_ = new_B9522_ | new_B9521_;
  assign new_B9511_ = new_B9500_ | new_B9523_;
  assign B9510 = new_B9511_ | new_B9520_;
  assign B9509 = new_B9518_ & new_B9519_;
  assign B9508 = new_B9518_ & new_B9517_;
  assign B9507 = new_B9516_ | new_B9515_;
  assign B9506 = new_B9514_ | new_B9513_;
  assign B9505 = new_B9512_ & new_B9511_;
  assign new_B9504_ = new_D3715_;
  assign new_B9503_ = new_D3648_;
  assign new_B9502_ = new_D3581_;
  assign new_B9501_ = new_D3514_;
  assign new_B9500_ = new_D3447_;
  assign new_B9499_ = new_D3380_;
  assign new_B9498_ = ~new_B9437_ & new_B9451_;
  assign new_B9497_ = new_B9437_ & ~new_B9451_;
  assign new_B9496_ = new_B9437_ & ~new_B9451_;
  assign new_B9495_ = ~new_B9437_ & ~new_B9451_;
  assign new_B9494_ = new_B9437_ & new_B9451_;
  assign new_B9493_ = new_B9497_ | new_B9498_;
  assign new_B9492_ = ~new_B9437_ & new_B9451_;
  assign new_B9491_ = new_B9495_ | new_B9496_;
  assign new_B9490_ = ~new_B9466_ & ~new_B9486_;
  assign new_B9489_ = new_B9466_ & new_B9486_;
  assign new_B9488_ = ~new_B9433_ | ~new_B9458_;
  assign new_B9487_ = new_B9451_ & new_B9488_;
  assign new_B9486_ = new_B9434_ | new_B9435_;
  assign new_B9485_ = new_B9434_ | new_B9451_;
  assign new_B9484_ = ~new_B9451_ & ~new_B9487_;
  assign new_B9483_ = new_B9451_ | new_B9488_;
  assign new_B9482_ = new_B9434_ & ~new_B9435_;
  assign new_B9481_ = ~new_B9434_ & new_B9435_;
  assign new_B9480_ = new_B9444_ | new_B9477_;
  assign new_B9479_ = ~new_B9444_ & ~new_B9478_;
  assign new_B9478_ = new_B9444_ & new_B9477_;
  assign new_B9477_ = ~new_B9433_ | ~new_B9458_;
  assign new_B9476_ = ~new_B9434_ & new_B9444_;
  assign new_B9475_ = new_B9434_ & ~new_B9444_;
  assign new_B9474_ = new_B9436_ & new_B9473_;
  assign new_B9473_ = new_B9492_ | new_B9491_;
  assign new_B9472_ = ~new_B9436_ & new_B9471_;
  assign new_B9471_ = new_B9494_ | new_B9493_;
  assign new_B9470_ = new_B9436_ | new_B9469_;
  assign new_B9469_ = new_B9490_ | new_B9489_;
  assign new_B9468_ = ~new_B9448_ & ~new_B9458_;
  assign new_B9467_ = new_B9448_ & new_B9458_;
  assign new_B9466_ = ~new_B9448_ | new_B9458_;
  assign new_B9465_ = new_B9432_ & ~new_B9433_;
  assign new_B9464_ = ~new_B9432_ & new_B9433_;
  assign new_B9463_ = new_B9485_ & ~new_B9486_;
  assign new_B9462_ = ~new_B9485_ & new_B9486_;
  assign new_B9461_ = ~new_B9484_ | ~new_B9483_;
  assign new_B9460_ = new_B9476_ | new_B9475_;
  assign new_B9459_ = new_B9482_ | new_B9481_;
  assign new_B9458_ = new_B9472_ | new_B9474_;
  assign new_B9457_ = ~new_B9479_ | ~new_B9480_;
  assign new_B9456_ = new_B9432_ & ~new_B9433_;
  assign new_B9455_ = new_B9446_ & ~new_B9458_;
  assign new_B9454_ = ~new_B9446_ & new_B9458_;
  assign new_B9453_ = ~new_B9444_ & new_B9470_;
  assign new_B9452_ = new_B9468_ | new_B9467_;
  assign new_B9451_ = new_B9465_ | new_B9464_;
  assign new_B9450_ = new_B9433_ | new_B9466_;
  assign new_B9449_ = new_B9458_ & new_B9461_;
  assign new_B9448_ = new_B9463_ | new_B9462_;
  assign new_B9447_ = new_B9458_ & new_B9457_;
  assign new_B9446_ = new_B9460_ & new_B9459_;
  assign new_B9445_ = new_B9455_ | new_B9454_;
  assign new_B9444_ = new_B9433_ | new_B9456_;
  assign B9443 = new_B9444_ | new_B9453_;
  assign B9442 = new_B9451_ & new_B9452_;
  assign B9441 = new_B9451_ & new_B9450_;
  assign B9440 = new_B9449_ | new_B9448_;
  assign B9439 = new_B9447_ | new_B9446_;
  assign B9438 = new_B9445_ & new_B9444_;
  assign new_B9437_ = new_D3313_;
  assign new_B9436_ = new_D3246_;
  assign new_B9435_ = new_D3179_;
  assign new_B9434_ = new_D3112_;
  assign new_B9433_ = new_D3045_;
  assign new_B9432_ = new_D2978_;
  assign new_B9431_ = ~new_B9370_ & new_B9384_;
  assign new_B9430_ = new_B9370_ & ~new_B9384_;
  assign new_B9429_ = new_B9370_ & ~new_B9384_;
  assign new_B9428_ = ~new_B9370_ & ~new_B9384_;
  assign new_B9427_ = new_B9370_ & new_B9384_;
  assign new_B9426_ = new_B9430_ | new_B9431_;
  assign new_B9425_ = ~new_B9370_ & new_B9384_;
  assign new_B9424_ = new_B9428_ | new_B9429_;
  assign new_B9423_ = ~new_B9399_ & ~new_B9419_;
  assign new_B9422_ = new_B9399_ & new_B9419_;
  assign new_B9421_ = ~new_B9366_ | ~new_B9391_;
  assign new_B9420_ = new_B9384_ & new_B9421_;
  assign new_B9419_ = new_B9367_ | new_B9368_;
  assign new_B9418_ = new_B9367_ | new_B9384_;
  assign new_B9417_ = ~new_B9384_ & ~new_B9420_;
  assign new_B9416_ = new_B9384_ | new_B9421_;
  assign new_B9415_ = new_B9367_ & ~new_B9368_;
  assign new_B9414_ = ~new_B9367_ & new_B9368_;
  assign new_B9413_ = new_B9377_ | new_B9410_;
  assign new_B9412_ = ~new_B9377_ & ~new_B9411_;
  assign new_B9411_ = new_B9377_ & new_B9410_;
  assign new_B9410_ = ~new_B9366_ | ~new_B9391_;
  assign new_B9409_ = ~new_B9367_ & new_B9377_;
  assign new_B9408_ = new_B9367_ & ~new_B9377_;
  assign new_B9407_ = new_B9369_ & new_B9406_;
  assign new_B9406_ = new_B9425_ | new_B9424_;
  assign new_B9405_ = ~new_B9369_ & new_B9404_;
  assign new_B9404_ = new_B9427_ | new_B9426_;
  assign new_B9403_ = new_B9369_ | new_B9402_;
  assign new_B9402_ = new_B9423_ | new_B9422_;
  assign new_B9401_ = ~new_B9381_ & ~new_B9391_;
  assign new_B9400_ = new_B9381_ & new_B9391_;
  assign new_B9399_ = ~new_B9381_ | new_B9391_;
  assign new_B9398_ = new_B9365_ & ~new_B9366_;
  assign new_B9397_ = ~new_B9365_ & new_B9366_;
  assign new_B9396_ = new_B9418_ & ~new_B9419_;
  assign new_B9395_ = ~new_B9418_ & new_B9419_;
  assign new_B9394_ = ~new_B9417_ | ~new_B9416_;
  assign new_B9393_ = new_B9409_ | new_B9408_;
  assign new_B9392_ = new_B9415_ | new_B9414_;
  assign new_B9391_ = new_B9405_ | new_B9407_;
  assign new_B9390_ = ~new_B9412_ | ~new_B9413_;
  assign new_B9389_ = new_B9365_ & ~new_B9366_;
  assign new_B9388_ = new_B9379_ & ~new_B9391_;
  assign new_B9387_ = ~new_B9379_ & new_B9391_;
  assign new_B9386_ = ~new_B9377_ & new_B9403_;
  assign new_B9385_ = new_B9401_ | new_B9400_;
  assign new_B9384_ = new_B9398_ | new_B9397_;
  assign new_B9383_ = new_B9366_ | new_B9399_;
  assign new_B9382_ = new_B9391_ & new_B9394_;
  assign new_B9381_ = new_B9396_ | new_B9395_;
  assign new_B9380_ = new_B9391_ & new_B9390_;
  assign new_B9379_ = new_B9393_ & new_B9392_;
  assign new_B9378_ = new_B9388_ | new_B9387_;
  assign new_B9377_ = new_B9366_ | new_B9389_;
  assign B9376 = new_B9377_ | new_B9386_;
  assign B9375 = new_B9384_ & new_B9385_;
  assign B9374 = new_B9384_ & new_B9383_;
  assign B9373 = new_B9382_ | new_B9381_;
  assign B9372 = new_B9380_ | new_B9379_;
  assign B9371 = new_B9378_ & new_B9377_;
  assign new_B9370_ = new_D2911_;
  assign new_B9369_ = new_D2844_;
  assign new_B9368_ = new_D2777_;
  assign new_B9367_ = new_D2710_;
  assign new_B9366_ = new_D2643_;
  assign new_B9365_ = new_D2576_;
  assign new_B9364_ = ~new_B9303_ & new_B9317_;
  assign new_B9363_ = new_B9303_ & ~new_B9317_;
  assign new_B9362_ = new_B9303_ & ~new_B9317_;
  assign new_B9361_ = ~new_B9303_ & ~new_B9317_;
  assign new_B9360_ = new_B9303_ & new_B9317_;
  assign new_B9359_ = new_B9363_ | new_B9364_;
  assign new_B9358_ = ~new_B9303_ & new_B9317_;
  assign new_B9357_ = new_B9361_ | new_B9362_;
  assign new_B9356_ = ~new_B9332_ & ~new_B9352_;
  assign new_B9355_ = new_B9332_ & new_B9352_;
  assign new_B9354_ = ~new_B9299_ | ~new_B9324_;
  assign new_B9353_ = new_B9317_ & new_B9354_;
  assign new_B9352_ = new_B9300_ | new_B9301_;
  assign new_B9351_ = new_B9300_ | new_B9317_;
  assign new_B9350_ = ~new_B9317_ & ~new_B9353_;
  assign new_B9349_ = new_B9317_ | new_B9354_;
  assign new_B9348_ = new_B9300_ & ~new_B9301_;
  assign new_B9347_ = ~new_B9300_ & new_B9301_;
  assign new_B9346_ = new_B9310_ | new_B9343_;
  assign new_B9345_ = ~new_B9310_ & ~new_B9344_;
  assign new_B9344_ = new_B9310_ & new_B9343_;
  assign new_B9343_ = ~new_B9299_ | ~new_B9324_;
  assign new_B9342_ = ~new_B9300_ & new_B9310_;
  assign new_B9341_ = new_B9300_ & ~new_B9310_;
  assign new_B9340_ = new_B9302_ & new_B9339_;
  assign new_B9339_ = new_B9358_ | new_B9357_;
  assign new_B9338_ = ~new_B9302_ & new_B9337_;
  assign new_B9337_ = new_B9360_ | new_B9359_;
  assign new_B9336_ = new_B9302_ | new_B9335_;
  assign new_B9335_ = new_B9356_ | new_B9355_;
  assign new_B9334_ = ~new_B9314_ & ~new_B9324_;
  assign new_B9333_ = new_B9314_ & new_B9324_;
  assign new_B9332_ = ~new_B9314_ | new_B9324_;
  assign new_B9331_ = new_B9298_ & ~new_B9299_;
  assign new_B9330_ = ~new_B9298_ & new_B9299_;
  assign new_B9329_ = new_B9351_ & ~new_B9352_;
  assign new_B9328_ = ~new_B9351_ & new_B9352_;
  assign new_B9327_ = ~new_B9350_ | ~new_B9349_;
  assign new_B9326_ = new_B9342_ | new_B9341_;
  assign new_B9325_ = new_B9348_ | new_B9347_;
  assign new_B9324_ = new_B9338_ | new_B9340_;
  assign new_B9323_ = ~new_B9345_ | ~new_B9346_;
  assign new_B9322_ = new_B9298_ & ~new_B9299_;
  assign new_B9321_ = new_B9312_ & ~new_B9324_;
  assign new_B9320_ = ~new_B9312_ & new_B9324_;
  assign new_B9319_ = ~new_B9310_ & new_B9336_;
  assign new_B9318_ = new_B9334_ | new_B9333_;
  assign new_B9317_ = new_B9331_ | new_B9330_;
  assign new_B9316_ = new_B9299_ | new_B9332_;
  assign new_B9315_ = new_B9324_ & new_B9327_;
  assign new_B9314_ = new_B9329_ | new_B9328_;
  assign new_B9313_ = new_B9324_ & new_B9323_;
  assign new_B9312_ = new_B9326_ & new_B9325_;
  assign new_B9311_ = new_B9321_ | new_B9320_;
  assign new_B9310_ = new_B9299_ | new_B9322_;
  assign B9309 = new_B9310_ | new_B9319_;
  assign B9308 = new_B9317_ & new_B9318_;
  assign B9307 = new_B9317_ & new_B9316_;
  assign B9306 = new_B9315_ | new_B9314_;
  assign B9305 = new_B9313_ | new_B9312_;
  assign B9304 = new_B9311_ & new_B9310_;
  assign new_B9303_ = new_D2509_;
  assign new_B9302_ = new_D2442_;
  assign new_B9301_ = new_D2375_;
  assign new_B9300_ = new_D2308_;
  assign new_B9299_ = new_D2241_;
  assign new_B9298_ = new_D2174_;
  assign new_B9297_ = ~new_B9236_ & new_B9250_;
  assign new_B9296_ = new_B9236_ & ~new_B9250_;
  assign new_B9295_ = new_B9236_ & ~new_B9250_;
  assign new_B9294_ = ~new_B9236_ & ~new_B9250_;
  assign new_B9293_ = new_B9236_ & new_B9250_;
  assign new_B9292_ = new_B9296_ | new_B9297_;
  assign new_B9291_ = ~new_B9236_ & new_B9250_;
  assign new_B9290_ = new_B9294_ | new_B9295_;
  assign new_B9289_ = ~new_B9265_ & ~new_B9285_;
  assign new_B9288_ = new_B9265_ & new_B9285_;
  assign new_B9287_ = ~new_B9232_ | ~new_B9257_;
  assign new_B9286_ = new_B9250_ & new_B9287_;
  assign new_B9285_ = new_B9233_ | new_B9234_;
  assign new_B9284_ = new_B9233_ | new_B9250_;
  assign new_B9283_ = ~new_B9250_ & ~new_B9286_;
  assign new_B9282_ = new_B9250_ | new_B9287_;
  assign new_B9281_ = new_B9233_ & ~new_B9234_;
  assign new_B9280_ = ~new_B9233_ & new_B9234_;
  assign new_B9279_ = new_B9243_ | new_B9276_;
  assign new_B9278_ = ~new_B9243_ & ~new_B9277_;
  assign new_B9277_ = new_B9243_ & new_B9276_;
  assign new_B9276_ = ~new_B9232_ | ~new_B9257_;
  assign new_B9275_ = ~new_B9233_ & new_B9243_;
  assign new_B9274_ = new_B9233_ & ~new_B9243_;
  assign new_B9273_ = new_B9235_ & new_B9272_;
  assign new_B9272_ = new_B9291_ | new_B9290_;
  assign new_B9271_ = ~new_B9235_ & new_B9270_;
  assign new_B9270_ = new_B9293_ | new_B9292_;
  assign new_B9269_ = new_B9235_ | new_B9268_;
  assign new_B9268_ = new_B9289_ | new_B9288_;
  assign new_B9267_ = ~new_B9247_ & ~new_B9257_;
  assign new_B9266_ = new_B9247_ & new_B9257_;
  assign new_B9265_ = ~new_B9247_ | new_B9257_;
  assign new_B9264_ = new_B9231_ & ~new_B9232_;
  assign new_B9263_ = ~new_B9231_ & new_B9232_;
  assign new_B9262_ = new_B9284_ & ~new_B9285_;
  assign new_B9261_ = ~new_B9284_ & new_B9285_;
  assign new_B9260_ = ~new_B9283_ | ~new_B9282_;
  assign new_B9259_ = new_B9275_ | new_B9274_;
  assign new_B9258_ = new_B9281_ | new_B9280_;
  assign new_B9257_ = new_B9271_ | new_B9273_;
  assign new_B9256_ = ~new_B9278_ | ~new_B9279_;
  assign new_B9255_ = new_B9231_ & ~new_B9232_;
  assign new_B9254_ = new_B9245_ & ~new_B9257_;
  assign new_B9253_ = ~new_B9245_ & new_B9257_;
  assign new_B9252_ = ~new_B9243_ & new_B9269_;
  assign new_B9251_ = new_B9267_ | new_B9266_;
  assign new_B9250_ = new_B9264_ | new_B9263_;
  assign new_B9249_ = new_B9232_ | new_B9265_;
  assign new_B9248_ = new_B9257_ & new_B9260_;
  assign new_B9247_ = new_B9262_ | new_B9261_;
  assign new_B9246_ = new_B9257_ & new_B9256_;
  assign new_B9245_ = new_B9259_ & new_B9258_;
  assign new_B9244_ = new_B9254_ | new_B9253_;
  assign new_B9243_ = new_B9232_ | new_B9255_;
  assign B9242 = new_B9243_ | new_B9252_;
  assign B9241 = new_B9250_ & new_B9251_;
  assign B9240 = new_B9250_ & new_B9249_;
  assign B9239 = new_B9248_ | new_B9247_;
  assign B9238 = new_B9246_ | new_B9245_;
  assign B9237 = new_B9244_ & new_B9243_;
  assign new_B9236_ = new_D2107_;
  assign new_B9235_ = new_D2040_;
  assign new_B9234_ = new_D1973_;
  assign new_B9233_ = new_D1906_;
  assign new_B9232_ = new_D1839_;
  assign new_B9231_ = new_D1772_;
  assign new_B9230_ = ~new_B9169_ & new_B9183_;
  assign new_B9229_ = new_B9169_ & ~new_B9183_;
  assign new_B9228_ = new_B9169_ & ~new_B9183_;
  assign new_B9227_ = ~new_B9169_ & ~new_B9183_;
  assign new_B9226_ = new_B9169_ & new_B9183_;
  assign new_B9225_ = new_B9229_ | new_B9230_;
  assign new_B9224_ = ~new_B9169_ & new_B9183_;
  assign new_B9223_ = new_B9227_ | new_B9228_;
  assign new_B9222_ = ~new_B9198_ & ~new_B9218_;
  assign new_B9221_ = new_B9198_ & new_B9218_;
  assign new_B9220_ = ~new_B9165_ | ~new_B9190_;
  assign new_B9219_ = new_B9183_ & new_B9220_;
  assign new_B9218_ = new_B9166_ | new_B9167_;
  assign new_B9217_ = new_B9166_ | new_B9183_;
  assign new_B9216_ = ~new_B9183_ & ~new_B9219_;
  assign new_B9215_ = new_B9183_ | new_B9220_;
  assign new_B9214_ = new_B9166_ & ~new_B9167_;
  assign new_B9213_ = ~new_B9166_ & new_B9167_;
  assign new_B9212_ = new_B9176_ | new_B9209_;
  assign new_B9211_ = ~new_B9176_ & ~new_B9210_;
  assign new_B9210_ = new_B9176_ & new_B9209_;
  assign new_B9209_ = ~new_B9165_ | ~new_B9190_;
  assign new_B9208_ = ~new_B9166_ & new_B9176_;
  assign new_B9207_ = new_B9166_ & ~new_B9176_;
  assign new_B9206_ = new_B9168_ & new_B9205_;
  assign new_B9205_ = new_B9224_ | new_B9223_;
  assign new_B9204_ = ~new_B9168_ & new_B9203_;
  assign new_B9203_ = new_B9226_ | new_B9225_;
  assign new_B9202_ = new_B9168_ | new_B9201_;
  assign new_B9201_ = new_B9222_ | new_B9221_;
  assign new_B9200_ = ~new_B9180_ & ~new_B9190_;
  assign new_B9199_ = new_B9180_ & new_B9190_;
  assign new_B9198_ = ~new_B9180_ | new_B9190_;
  assign new_B9197_ = new_B9164_ & ~new_B9165_;
  assign new_B9196_ = ~new_B9164_ & new_B9165_;
  assign new_B9195_ = new_B9217_ & ~new_B9218_;
  assign new_B9194_ = ~new_B9217_ & new_B9218_;
  assign new_B9193_ = ~new_B9216_ | ~new_B9215_;
  assign new_B9192_ = new_B9208_ | new_B9207_;
  assign new_B9191_ = new_B9214_ | new_B9213_;
  assign new_B9190_ = new_B9204_ | new_B9206_;
  assign new_B9189_ = ~new_B9211_ | ~new_B9212_;
  assign new_B9188_ = new_B9164_ & ~new_B9165_;
  assign new_B9187_ = new_B9178_ & ~new_B9190_;
  assign new_B9186_ = ~new_B9178_ & new_B9190_;
  assign new_B9185_ = ~new_B9176_ & new_B9202_;
  assign new_B9184_ = new_B9200_ | new_B9199_;
  assign new_B9183_ = new_B9197_ | new_B9196_;
  assign new_B9182_ = new_B9165_ | new_B9198_;
  assign new_B9181_ = new_B9190_ & new_B9193_;
  assign new_B9180_ = new_B9195_ | new_B9194_;
  assign new_B9179_ = new_B9190_ & new_B9189_;
  assign new_B9178_ = new_B9192_ & new_B9191_;
  assign new_B9177_ = new_B9187_ | new_B9186_;
  assign new_B9176_ = new_B9165_ | new_B9188_;
  assign B9175 = new_B9176_ | new_B9185_;
  assign B9174 = new_B9183_ & new_B9184_;
  assign B9173 = new_B9183_ & new_B9182_;
  assign B9172 = new_B9181_ | new_B9180_;
  assign B9171 = new_B9179_ | new_B9178_;
  assign B9170 = new_B9177_ & new_B9176_;
  assign new_B9169_ = new_D1705_;
  assign new_B9168_ = new_D1638_;
  assign new_B9167_ = new_D1571_;
  assign new_B9166_ = new_D1504_;
  assign new_B9165_ = new_D1437_;
  assign new_B9164_ = new_D1370_;
  assign new_B9163_ = ~new_B9102_ & new_B9116_;
  assign new_B9162_ = new_B9102_ & ~new_B9116_;
  assign new_B9161_ = new_B9102_ & ~new_B9116_;
  assign new_B9160_ = ~new_B9102_ & ~new_B9116_;
  assign new_B9159_ = new_B9102_ & new_B9116_;
  assign new_B9158_ = new_B9162_ | new_B9163_;
  assign new_B9157_ = ~new_B9102_ & new_B9116_;
  assign new_B9156_ = new_B9160_ | new_B9161_;
  assign new_B9155_ = ~new_B9131_ & ~new_B9151_;
  assign new_B9154_ = new_B9131_ & new_B9151_;
  assign new_B9153_ = ~new_B9098_ | ~new_B9123_;
  assign new_B9152_ = new_B9116_ & new_B9153_;
  assign new_B9151_ = new_B9099_ | new_B9100_;
  assign new_B9150_ = new_B9099_ | new_B9116_;
  assign new_B9149_ = ~new_B9116_ & ~new_B9152_;
  assign new_B9148_ = new_B9116_ | new_B9153_;
  assign new_B9147_ = new_B9099_ & ~new_B9100_;
  assign new_B9146_ = ~new_B9099_ & new_B9100_;
  assign new_B9145_ = new_B9109_ | new_B9142_;
  assign new_B9144_ = ~new_B9109_ & ~new_B9143_;
  assign new_B9143_ = new_B9109_ & new_B9142_;
  assign new_B9142_ = ~new_B9098_ | ~new_B9123_;
  assign new_B9141_ = ~new_B9099_ & new_B9109_;
  assign new_B9140_ = new_B9099_ & ~new_B9109_;
  assign new_B9139_ = new_B9101_ & new_B9138_;
  assign new_B9138_ = new_B9157_ | new_B9156_;
  assign new_B9137_ = ~new_B9101_ & new_B9136_;
  assign new_B9136_ = new_B9159_ | new_B9158_;
  assign new_B9135_ = new_B9101_ | new_B9134_;
  assign new_B9134_ = new_B9155_ | new_B9154_;
  assign new_B9133_ = ~new_B9113_ & ~new_B9123_;
  assign new_B9132_ = new_B9113_ & new_B9123_;
  assign new_B9131_ = ~new_B9113_ | new_B9123_;
  assign new_B9130_ = new_B9097_ & ~new_B9098_;
  assign new_B9129_ = ~new_B9097_ & new_B9098_;
  assign new_B9128_ = new_B9150_ & ~new_B9151_;
  assign new_B9127_ = ~new_B9150_ & new_B9151_;
  assign new_B9126_ = ~new_B9149_ | ~new_B9148_;
  assign new_B9125_ = new_B9141_ | new_B9140_;
  assign new_B9124_ = new_B9147_ | new_B9146_;
  assign new_B9123_ = new_B9137_ | new_B9139_;
  assign new_B9122_ = ~new_B9144_ | ~new_B9145_;
  assign new_B9121_ = new_B9097_ & ~new_B9098_;
  assign new_B9120_ = new_B9111_ & ~new_B9123_;
  assign new_B9119_ = ~new_B9111_ & new_B9123_;
  assign new_B9118_ = ~new_B9109_ & new_B9135_;
  assign new_B9117_ = new_B9133_ | new_B9132_;
  assign new_B9116_ = new_B9130_ | new_B9129_;
  assign new_B9115_ = new_B9098_ | new_B9131_;
  assign new_B9114_ = new_B9123_ & new_B9126_;
  assign new_B9113_ = new_B9128_ | new_B9127_;
  assign new_B9112_ = new_B9123_ & new_B9122_;
  assign new_B9111_ = new_B9125_ & new_B9124_;
  assign new_B9110_ = new_B9120_ | new_B9119_;
  assign new_B9109_ = new_B9098_ | new_B9121_;
  assign B9108 = new_B9109_ | new_B9118_;
  assign B9107 = new_B9116_ & new_B9117_;
  assign B9106 = new_B9116_ & new_B9115_;
  assign B9105 = new_B9114_ | new_B9113_;
  assign B9104 = new_B9112_ | new_B9111_;
  assign B9103 = new_B9110_ & new_B9109_;
  assign new_B9102_ = new_D1303_;
  assign new_B9101_ = new_D1236_;
  assign new_B9100_ = new_D1169_;
  assign new_B9099_ = new_D1102_;
  assign new_B9098_ = new_D1035_;
  assign new_B9097_ = new_D968_;
  assign new_B9096_ = ~new_B9035_ & new_B9049_;
  assign new_B9095_ = new_B9035_ & ~new_B9049_;
  assign new_B9094_ = new_B9035_ & ~new_B9049_;
  assign new_B9093_ = ~new_B9035_ & ~new_B9049_;
  assign new_B9092_ = new_B9035_ & new_B9049_;
  assign new_B9091_ = new_B9095_ | new_B9096_;
  assign new_B9090_ = ~new_B9035_ & new_B9049_;
  assign new_B9089_ = new_B9093_ | new_B9094_;
  assign new_B9088_ = ~new_B9064_ & ~new_B9084_;
  assign new_B9087_ = new_B9064_ & new_B9084_;
  assign new_B9086_ = ~new_B9031_ | ~new_B9056_;
  assign new_B9085_ = new_B9049_ & new_B9086_;
  assign new_B9084_ = new_B9032_ | new_B9033_;
  assign new_B9083_ = new_B9032_ | new_B9049_;
  assign new_B9082_ = ~new_B9049_ & ~new_B9085_;
  assign new_B9081_ = new_B9049_ | new_B9086_;
  assign new_B9080_ = new_B9032_ & ~new_B9033_;
  assign new_B9079_ = ~new_B9032_ & new_B9033_;
  assign new_B9078_ = new_B9042_ | new_B9075_;
  assign new_B9077_ = ~new_B9042_ & ~new_B9076_;
  assign new_B9076_ = new_B9042_ & new_B9075_;
  assign new_B9075_ = ~new_B9031_ | ~new_B9056_;
  assign new_B9074_ = ~new_B9032_ & new_B9042_;
  assign new_B9073_ = new_B9032_ & ~new_B9042_;
  assign new_B9072_ = new_B9034_ & new_B9071_;
  assign new_B9071_ = new_B9090_ | new_B9089_;
  assign new_B9070_ = ~new_B9034_ & new_B9069_;
  assign new_B9069_ = new_B9092_ | new_B9091_;
  assign new_B9068_ = new_B9034_ | new_B9067_;
  assign new_B9067_ = new_B9088_ | new_B9087_;
  assign new_B9066_ = ~new_B9046_ & ~new_B9056_;
  assign new_B9065_ = new_B9046_ & new_B9056_;
  assign new_B9064_ = ~new_B9046_ | new_B9056_;
  assign new_B9063_ = new_B9030_ & ~new_B9031_;
  assign new_B9062_ = ~new_B9030_ & new_B9031_;
  assign new_B9061_ = new_B9083_ & ~new_B9084_;
  assign new_B9060_ = ~new_B9083_ & new_B9084_;
  assign new_B9059_ = ~new_B9082_ | ~new_B9081_;
  assign new_B9058_ = new_B9074_ | new_B9073_;
  assign new_B9057_ = new_B9080_ | new_B9079_;
  assign new_B9056_ = new_B9070_ | new_B9072_;
  assign new_B9055_ = ~new_B9077_ | ~new_B9078_;
  assign new_B9054_ = new_B9030_ & ~new_B9031_;
  assign new_B9053_ = new_B9044_ & ~new_B9056_;
  assign new_B9052_ = ~new_B9044_ & new_B9056_;
  assign new_B9051_ = ~new_B9042_ & new_B9068_;
  assign new_B9050_ = new_B9066_ | new_B9065_;
  assign new_B9049_ = new_B9063_ | new_B9062_;
  assign new_B9048_ = new_B9031_ | new_B9064_;
  assign new_B9047_ = new_B9056_ & new_B9059_;
  assign new_B9046_ = new_B9061_ | new_B9060_;
  assign new_B9045_ = new_B9056_ & new_B9055_;
  assign new_B9044_ = new_B9058_ & new_B9057_;
  assign new_B9043_ = new_B9053_ | new_B9052_;
  assign new_B9042_ = new_B9031_ | new_B9054_;
  assign B9041 = new_B9042_ | new_B9051_;
  assign B9040 = new_B9049_ & new_B9050_;
  assign B9039 = new_B9049_ & new_B9048_;
  assign B9038 = new_B9047_ | new_B9046_;
  assign B9037 = new_B9045_ | new_B9044_;
  assign B9036 = new_B9043_ & new_B9042_;
  assign new_B9035_ = new_D901_;
  assign new_B9034_ = new_D834_;
  assign new_B9033_ = new_D767_;
  assign new_B9032_ = new_D700_;
  assign new_B9031_ = new_D633_;
  assign new_B9030_ = new_D566_;
  assign new_B9029_ = ~new_B8968_ & new_B8982_;
  assign new_B9028_ = new_B8968_ & ~new_B8982_;
  assign new_B9027_ = new_B8968_ & ~new_B8982_;
  assign new_B9026_ = ~new_B8968_ & ~new_B8982_;
  assign new_B9025_ = new_B8968_ & new_B8982_;
  assign new_B9024_ = new_B9028_ | new_B9029_;
  assign new_B9023_ = ~new_B8968_ & new_B8982_;
  assign new_B9022_ = new_B9026_ | new_B9027_;
  assign new_B9021_ = ~new_B8997_ & ~new_B9017_;
  assign new_B9020_ = new_B8997_ & new_B9017_;
  assign new_B9019_ = ~new_B8964_ | ~new_B8989_;
  assign new_B9018_ = new_B8982_ & new_B9019_;
  assign new_B9017_ = new_B8965_ | new_B8966_;
  assign new_B9016_ = new_B8965_ | new_B8982_;
  assign new_B9015_ = ~new_B8982_ & ~new_B9018_;
  assign new_B9014_ = new_B8982_ | new_B9019_;
  assign new_B9013_ = new_B8965_ & ~new_B8966_;
  assign new_B9012_ = ~new_B8965_ & new_B8966_;
  assign new_B9011_ = new_B8975_ | new_B9008_;
  assign new_B9010_ = ~new_B8975_ & ~new_B9009_;
  assign new_B9009_ = new_B8975_ & new_B9008_;
  assign new_B9008_ = ~new_B8964_ | ~new_B8989_;
  assign new_B9007_ = ~new_B8965_ & new_B8975_;
  assign new_B9006_ = new_B8965_ & ~new_B8975_;
  assign new_B9005_ = new_B8967_ & new_B9004_;
  assign new_B9004_ = new_B9023_ | new_B9022_;
  assign new_B9003_ = ~new_B8967_ & new_B9002_;
  assign new_B9002_ = new_B9025_ | new_B9024_;
  assign new_B9001_ = new_B8967_ | new_B9000_;
  assign new_B9000_ = new_B9021_ | new_B9020_;
  assign new_B8999_ = ~new_B8979_ & ~new_B8989_;
  assign new_B8998_ = new_B8979_ & new_B8989_;
  assign new_B8997_ = ~new_B8979_ | new_B8989_;
  assign new_B8996_ = new_B8963_ & ~new_B8964_;
  assign new_B8995_ = ~new_B8963_ & new_B8964_;
  assign new_B8994_ = new_B9016_ & ~new_B9017_;
  assign new_B8993_ = ~new_B9016_ & new_B9017_;
  assign new_B8992_ = ~new_B9015_ | ~new_B9014_;
  assign new_B8991_ = new_B9007_ | new_B9006_;
  assign new_B8990_ = new_B9013_ | new_B9012_;
  assign new_B8989_ = new_B9003_ | new_B9005_;
  assign new_B8988_ = ~new_B9010_ | ~new_B9011_;
  assign new_B8987_ = new_B8963_ & ~new_B8964_;
  assign new_B8986_ = new_B8977_ & ~new_B8989_;
  assign new_B8985_ = ~new_B8977_ & new_B8989_;
  assign new_B8984_ = ~new_B8975_ & new_B9001_;
  assign new_B8983_ = new_B8999_ | new_B8998_;
  assign new_B8982_ = new_B8996_ | new_B8995_;
  assign new_B8981_ = new_B8964_ | new_B8997_;
  assign new_B8980_ = new_B8989_ & new_B8992_;
  assign new_B8979_ = new_B8994_ | new_B8993_;
  assign new_B8978_ = new_B8989_ & new_B8988_;
  assign new_B8977_ = new_B8991_ & new_B8990_;
  assign new_B8976_ = new_B8986_ | new_B8985_;
  assign new_B8975_ = new_B8964_ | new_B8987_;
  assign B8974 = new_B8975_ | new_B8984_;
  assign B8973 = new_B8982_ & new_B8983_;
  assign B8972 = new_B8982_ & new_B8981_;
  assign B8971 = new_B8980_ | new_B8979_;
  assign B8970 = new_B8978_ | new_B8977_;
  assign B8969 = new_B8976_ & new_B8975_;
  assign new_B8968_ = new_D499_;
  assign new_B8967_ = new_D432_;
  assign new_B8966_ = new_D365_;
  assign new_B8965_ = new_D298_;
  assign new_B8964_ = new_D231_;
  assign new_B8963_ = new_D164_;
  assign new_B8962_ = ~new_B8901_ & new_B8915_;
  assign new_B8961_ = new_B8901_ & ~new_B8915_;
  assign new_B8960_ = new_B8901_ & ~new_B8915_;
  assign new_B8959_ = ~new_B8901_ & ~new_B8915_;
  assign new_B8958_ = new_B8901_ & new_B8915_;
  assign new_B8957_ = new_B8961_ | new_B8962_;
  assign new_B8956_ = ~new_B8901_ & new_B8915_;
  assign new_B8955_ = new_B8959_ | new_B8960_;
  assign new_B8954_ = ~new_B8930_ & ~new_B8950_;
  assign new_B8953_ = new_B8930_ & new_B8950_;
  assign new_B8952_ = ~new_B8897_ | ~new_B8922_;
  assign new_B8951_ = new_B8915_ & new_B8952_;
  assign new_B8950_ = new_B8898_ | new_B8899_;
  assign new_B8949_ = new_B8898_ | new_B8915_;
  assign new_B8948_ = ~new_B8915_ & ~new_B8951_;
  assign new_B8947_ = new_B8915_ | new_B8952_;
  assign new_B8946_ = new_B8898_ & ~new_B8899_;
  assign new_B8945_ = ~new_B8898_ & new_B8899_;
  assign new_B8944_ = new_B8908_ | new_B8941_;
  assign new_B8943_ = ~new_B8908_ & ~new_B8942_;
  assign new_B8942_ = new_B8908_ & new_B8941_;
  assign new_B8941_ = ~new_B8897_ | ~new_B8922_;
  assign new_B8940_ = ~new_B8898_ & new_B8908_;
  assign new_B8939_ = new_B8898_ & ~new_B8908_;
  assign new_B8938_ = new_B8900_ & new_B8937_;
  assign new_B8937_ = new_B8956_ | new_B8955_;
  assign new_B8936_ = ~new_B8900_ & new_B8935_;
  assign new_B8935_ = new_B8958_ | new_B8957_;
  assign new_B8934_ = new_B8900_ | new_B8933_;
  assign new_B8933_ = new_B8954_ | new_B8953_;
  assign new_B8932_ = ~new_B8912_ & ~new_B8922_;
  assign new_B8931_ = new_B8912_ & new_B8922_;
  assign new_B8930_ = ~new_B8912_ | new_B8922_;
  assign new_B8929_ = new_B8896_ & ~new_B8897_;
  assign new_B8928_ = ~new_B8896_ & new_B8897_;
  assign new_B8927_ = new_B8949_ & ~new_B8950_;
  assign new_B8926_ = ~new_B8949_ & new_B8950_;
  assign new_B8925_ = ~new_B8948_ | ~new_B8947_;
  assign new_B8924_ = new_B8940_ | new_B8939_;
  assign new_B8923_ = new_B8946_ | new_B8945_;
  assign new_B8922_ = new_B8936_ | new_B8938_;
  assign new_B8921_ = ~new_B8943_ | ~new_B8944_;
  assign new_B8920_ = new_B8896_ & ~new_B8897_;
  assign new_B8919_ = new_B8910_ & ~new_B8922_;
  assign new_B8918_ = ~new_B8910_ & new_B8922_;
  assign new_B8917_ = ~new_B8908_ & new_B8934_;
  assign new_B8916_ = new_B8932_ | new_B8931_;
  assign new_B8915_ = new_B8929_ | new_B8928_;
  assign new_B8914_ = new_B8897_ | new_B8930_;
  assign new_B8913_ = new_B8922_ & new_B8925_;
  assign new_B8912_ = new_B8927_ | new_B8926_;
  assign new_B8911_ = new_B8922_ & new_B8921_;
  assign new_B8910_ = new_B8924_ & new_B8923_;
  assign new_B8909_ = new_B8919_ | new_B8918_;
  assign new_B8908_ = new_B8897_ | new_B8920_;
  assign B8907 = new_B8908_ | new_B8917_;
  assign B8906 = new_B8915_ & new_B8916_;
  assign B8905 = new_B8915_ & new_B8914_;
  assign B8904 = new_B8913_ | new_B8912_;
  assign B8903 = new_B8911_ | new_B8910_;
  assign B8902 = new_B8909_ & new_B8908_;
  assign new_B8901_ = new_D97_;
  assign new_B8900_ = new_D30_;
  assign new_B8899_ = new_C9962_;
  assign new_B8898_ = new_C9895_;
  assign new_B8897_ = new_C9828_;
  assign new_B8896_ = new_C9761_;
  assign new_B8895_ = ~new_B8834_ & new_B8848_;
  assign new_B8894_ = new_B8834_ & ~new_B8848_;
  assign new_B8893_ = new_B8834_ & ~new_B8848_;
  assign new_B8892_ = ~new_B8834_ & ~new_B8848_;
  assign new_B8891_ = new_B8834_ & new_B8848_;
  assign new_B8890_ = new_B8894_ | new_B8895_;
  assign new_B8889_ = ~new_B8834_ & new_B8848_;
  assign new_B8888_ = new_B8892_ | new_B8893_;
  assign new_B8887_ = ~new_B8863_ & ~new_B8883_;
  assign new_B8886_ = new_B8863_ & new_B8883_;
  assign new_B8885_ = ~new_B8830_ | ~new_B8855_;
  assign new_B8884_ = new_B8848_ & new_B8885_;
  assign new_B8883_ = new_B8831_ | new_B8832_;
  assign new_B8882_ = new_B8831_ | new_B8848_;
  assign new_B8881_ = ~new_B8848_ & ~new_B8884_;
  assign new_B8880_ = new_B8848_ | new_B8885_;
  assign new_B8879_ = new_B8831_ & ~new_B8832_;
  assign new_B8878_ = ~new_B8831_ & new_B8832_;
  assign new_B8877_ = new_B8841_ | new_B8874_;
  assign new_B8876_ = ~new_B8841_ & ~new_B8875_;
  assign new_B8875_ = new_B8841_ & new_B8874_;
  assign new_B8874_ = ~new_B8830_ | ~new_B8855_;
  assign new_B8873_ = ~new_B8831_ & new_B8841_;
  assign new_B8872_ = new_B8831_ & ~new_B8841_;
  assign new_B8871_ = new_B8833_ & new_B8870_;
  assign new_B8870_ = new_B8889_ | new_B8888_;
  assign new_B8869_ = ~new_B8833_ & new_B8868_;
  assign new_B8868_ = new_B8891_ | new_B8890_;
  assign new_B8867_ = new_B8833_ | new_B8866_;
  assign new_B8866_ = new_B8887_ | new_B8886_;
  assign new_B8865_ = ~new_B8845_ & ~new_B8855_;
  assign new_B8864_ = new_B8845_ & new_B8855_;
  assign new_B8863_ = ~new_B8845_ | new_B8855_;
  assign new_B8862_ = new_B8829_ & ~new_B8830_;
  assign new_B8861_ = ~new_B8829_ & new_B8830_;
  assign new_B8860_ = new_B8882_ & ~new_B8883_;
  assign new_B8859_ = ~new_B8882_ & new_B8883_;
  assign new_B8858_ = ~new_B8881_ | ~new_B8880_;
  assign new_B8857_ = new_B8873_ | new_B8872_;
  assign new_B8856_ = new_B8879_ | new_B8878_;
  assign new_B8855_ = new_B8869_ | new_B8871_;
  assign new_B8854_ = ~new_B8876_ | ~new_B8877_;
  assign new_B8853_ = new_B8829_ & ~new_B8830_;
  assign new_B8852_ = new_B8843_ & ~new_B8855_;
  assign new_B8851_ = ~new_B8843_ & new_B8855_;
  assign new_B8850_ = ~new_B8841_ & new_B8867_;
  assign new_B8849_ = new_B8865_ | new_B8864_;
  assign new_B8848_ = new_B8862_ | new_B8861_;
  assign new_B8847_ = new_B8830_ | new_B8863_;
  assign new_B8846_ = new_B8855_ & new_B8858_;
  assign new_B8845_ = new_B8860_ | new_B8859_;
  assign new_B8844_ = new_B8855_ & new_B8854_;
  assign new_B8843_ = new_B8857_ & new_B8856_;
  assign new_B8842_ = new_B8852_ | new_B8851_;
  assign new_B8841_ = new_B8830_ | new_B8853_;
  assign B8840 = new_B8841_ | new_B8850_;
  assign B8839 = new_B8848_ & new_B8849_;
  assign B8838 = new_B8848_ & new_B8847_;
  assign B8837 = new_B8846_ | new_B8845_;
  assign B8836 = new_B8844_ | new_B8843_;
  assign B8835 = new_B8842_ & new_B8841_;
  assign new_B8834_ = new_C9694_;
  assign new_B8833_ = new_C9627_;
  assign new_B8832_ = new_C9560_;
  assign new_B8831_ = new_C9493_;
  assign new_B8830_ = new_C9426_;
  assign new_B8829_ = new_C9359_;
  assign new_B8828_ = ~new_B8767_ & new_B8781_;
  assign new_B8827_ = new_B8767_ & ~new_B8781_;
  assign new_B8826_ = new_B8767_ & ~new_B8781_;
  assign new_B8825_ = ~new_B8767_ & ~new_B8781_;
  assign new_B8824_ = new_B8767_ & new_B8781_;
  assign new_B8823_ = new_B8827_ | new_B8828_;
  assign new_B8822_ = ~new_B8767_ & new_B8781_;
  assign new_B8821_ = new_B8825_ | new_B8826_;
  assign new_B8820_ = ~new_B8796_ & ~new_B8816_;
  assign new_B8819_ = new_B8796_ & new_B8816_;
  assign new_B8818_ = ~new_B8763_ | ~new_B8788_;
  assign new_B8817_ = new_B8781_ & new_B8818_;
  assign new_B8816_ = new_B8764_ | new_B8765_;
  assign new_B8815_ = new_B8764_ | new_B8781_;
  assign new_B8814_ = ~new_B8781_ & ~new_B8817_;
  assign new_B8813_ = new_B8781_ | new_B8818_;
  assign new_B8812_ = new_B8764_ & ~new_B8765_;
  assign new_B8811_ = ~new_B8764_ & new_B8765_;
  assign new_B8810_ = new_B8774_ | new_B8807_;
  assign new_B8809_ = ~new_B8774_ & ~new_B8808_;
  assign new_B8808_ = new_B8774_ & new_B8807_;
  assign new_B8807_ = ~new_B8763_ | ~new_B8788_;
  assign new_B8806_ = ~new_B8764_ & new_B8774_;
  assign new_B8805_ = new_B8764_ & ~new_B8774_;
  assign new_B8804_ = new_B8766_ & new_B8803_;
  assign new_B8803_ = new_B8822_ | new_B8821_;
  assign new_B8802_ = ~new_B8766_ & new_B8801_;
  assign new_B8801_ = new_B8824_ | new_B8823_;
  assign new_B8800_ = new_B8766_ | new_B8799_;
  assign new_B8799_ = new_B8820_ | new_B8819_;
  assign new_B8798_ = ~new_B8778_ & ~new_B8788_;
  assign new_B8797_ = new_B8778_ & new_B8788_;
  assign new_B8796_ = ~new_B8778_ | new_B8788_;
  assign new_B8795_ = new_B8762_ & ~new_B8763_;
  assign new_B8794_ = ~new_B8762_ & new_B8763_;
  assign new_B8793_ = new_B8815_ & ~new_B8816_;
  assign new_B8792_ = ~new_B8815_ & new_B8816_;
  assign new_B8791_ = ~new_B8814_ | ~new_B8813_;
  assign new_B8790_ = new_B8806_ | new_B8805_;
  assign new_B8789_ = new_B8812_ | new_B8811_;
  assign new_B8788_ = new_B8802_ | new_B8804_;
  assign new_B8787_ = ~new_B8809_ | ~new_B8810_;
  assign new_B8786_ = new_B8762_ & ~new_B8763_;
  assign new_B8785_ = new_B8776_ & ~new_B8788_;
  assign new_B8784_ = ~new_B8776_ & new_B8788_;
  assign new_B8783_ = ~new_B8774_ & new_B8800_;
  assign new_B8782_ = new_B8798_ | new_B8797_;
  assign new_B8781_ = new_B8795_ | new_B8794_;
  assign new_B8780_ = new_B8763_ | new_B8796_;
  assign new_B8779_ = new_B8788_ & new_B8791_;
  assign new_B8778_ = new_B8793_ | new_B8792_;
  assign new_B8777_ = new_B8788_ & new_B8787_;
  assign new_B8776_ = new_B8790_ & new_B8789_;
  assign new_B8775_ = new_B8785_ | new_B8784_;
  assign new_B8774_ = new_B8763_ | new_B8786_;
  assign B8773 = new_B8774_ | new_B8783_;
  assign B8772 = new_B8781_ & new_B8782_;
  assign B8771 = new_B8781_ & new_B8780_;
  assign B8770 = new_B8779_ | new_B8778_;
  assign B8769 = new_B8777_ | new_B8776_;
  assign B8768 = new_B8775_ & new_B8774_;
  assign new_B8767_ = new_C9292_;
  assign new_B8766_ = new_C9225_;
  assign new_B8765_ = new_C9158_;
  assign new_B8764_ = new_C9091_;
  assign new_B8763_ = new_C9024_;
  assign new_B8762_ = new_C8957_;
  assign new_B8761_ = ~new_B8700_ & new_B8714_;
  assign new_B8760_ = new_B8700_ & ~new_B8714_;
  assign new_B8759_ = new_B8700_ & ~new_B8714_;
  assign new_B8758_ = ~new_B8700_ & ~new_B8714_;
  assign new_B8757_ = new_B8700_ & new_B8714_;
  assign new_B8756_ = new_B8760_ | new_B8761_;
  assign new_B8755_ = ~new_B8700_ & new_B8714_;
  assign new_B8754_ = new_B8758_ | new_B8759_;
  assign new_B8753_ = ~new_B8729_ & ~new_B8749_;
  assign new_B8752_ = new_B8729_ & new_B8749_;
  assign new_B8751_ = ~new_B8696_ | ~new_B8721_;
  assign new_B8750_ = new_B8714_ & new_B8751_;
  assign new_B8749_ = new_B8697_ | new_B8698_;
  assign new_B8748_ = new_B8697_ | new_B8714_;
  assign new_B8747_ = ~new_B8714_ & ~new_B8750_;
  assign new_B8746_ = new_B8714_ | new_B8751_;
  assign new_B8745_ = new_B8697_ & ~new_B8698_;
  assign new_B8744_ = ~new_B8697_ & new_B8698_;
  assign new_B8743_ = new_B8707_ | new_B8740_;
  assign new_B8742_ = ~new_B8707_ & ~new_B8741_;
  assign new_B8741_ = new_B8707_ & new_B8740_;
  assign new_B8740_ = ~new_B8696_ | ~new_B8721_;
  assign new_B8739_ = ~new_B8697_ & new_B8707_;
  assign new_B8738_ = new_B8697_ & ~new_B8707_;
  assign new_B8737_ = new_B8699_ & new_B8736_;
  assign new_B8736_ = new_B8755_ | new_B8754_;
  assign new_B8735_ = ~new_B8699_ & new_B8734_;
  assign new_B8734_ = new_B8757_ | new_B8756_;
  assign new_B8733_ = new_B8699_ | new_B8732_;
  assign new_B8732_ = new_B8753_ | new_B8752_;
  assign new_B8731_ = ~new_B8711_ & ~new_B8721_;
  assign new_B8730_ = new_B8711_ & new_B8721_;
  assign new_B8729_ = ~new_B8711_ | new_B8721_;
  assign new_B8728_ = new_B8695_ & ~new_B8696_;
  assign new_B8727_ = ~new_B8695_ & new_B8696_;
  assign new_B8726_ = new_B8748_ & ~new_B8749_;
  assign new_B8725_ = ~new_B8748_ & new_B8749_;
  assign new_B8724_ = ~new_B8747_ | ~new_B8746_;
  assign new_B8723_ = new_B8739_ | new_B8738_;
  assign new_B8722_ = new_B8745_ | new_B8744_;
  assign new_B8721_ = new_B8735_ | new_B8737_;
  assign new_B8720_ = ~new_B8742_ | ~new_B8743_;
  assign new_B8719_ = new_B8695_ & ~new_B8696_;
  assign new_B8718_ = new_B8709_ & ~new_B8721_;
  assign new_B8717_ = ~new_B8709_ & new_B8721_;
  assign new_B8716_ = ~new_B8707_ & new_B8733_;
  assign new_B8715_ = new_B8731_ | new_B8730_;
  assign new_B8714_ = new_B8728_ | new_B8727_;
  assign new_B8713_ = new_B8696_ | new_B8729_;
  assign new_B8712_ = new_B8721_ & new_B8724_;
  assign new_B8711_ = new_B8726_ | new_B8725_;
  assign new_B8710_ = new_B8721_ & new_B8720_;
  assign new_B8709_ = new_B8723_ & new_B8722_;
  assign new_B8708_ = new_B8718_ | new_B8717_;
  assign new_B8707_ = new_B8696_ | new_B8719_;
  assign B8706 = new_B8707_ | new_B8716_;
  assign B8705 = new_B8714_ & new_B8715_;
  assign B8704 = new_B8714_ & new_B8713_;
  assign B8703 = new_B8712_ | new_B8711_;
  assign B8702 = new_B8710_ | new_B8709_;
  assign B8701 = new_B8708_ & new_B8707_;
  assign new_B8700_ = new_C8890_;
  assign new_B8699_ = new_C8823_;
  assign new_B8698_ = new_C8756_;
  assign new_B8697_ = new_C8689_;
  assign new_B8696_ = new_C8622_;
  assign new_B8695_ = new_C8555_;
  assign new_B8694_ = ~new_B8633_ & new_B8647_;
  assign new_B8693_ = new_B8633_ & ~new_B8647_;
  assign new_B8692_ = new_B8633_ & ~new_B8647_;
  assign new_B8691_ = ~new_B8633_ & ~new_B8647_;
  assign new_B8690_ = new_B8633_ & new_B8647_;
  assign new_B8689_ = new_B8693_ | new_B8694_;
  assign new_B8688_ = ~new_B8633_ & new_B8647_;
  assign new_B8687_ = new_B8691_ | new_B8692_;
  assign new_B8686_ = ~new_B8662_ & ~new_B8682_;
  assign new_B8685_ = new_B8662_ & new_B8682_;
  assign new_B8684_ = ~new_B8629_ | ~new_B8654_;
  assign new_B8683_ = new_B8647_ & new_B8684_;
  assign new_B8682_ = new_B8630_ | new_B8631_;
  assign new_B8681_ = new_B8630_ | new_B8647_;
  assign new_B8680_ = ~new_B8647_ & ~new_B8683_;
  assign new_B8679_ = new_B8647_ | new_B8684_;
  assign new_B8678_ = new_B8630_ & ~new_B8631_;
  assign new_B8677_ = ~new_B8630_ & new_B8631_;
  assign new_B8676_ = new_B8640_ | new_B8673_;
  assign new_B8675_ = ~new_B8640_ & ~new_B8674_;
  assign new_B8674_ = new_B8640_ & new_B8673_;
  assign new_B8673_ = ~new_B8629_ | ~new_B8654_;
  assign new_B8672_ = ~new_B8630_ & new_B8640_;
  assign new_B8671_ = new_B8630_ & ~new_B8640_;
  assign new_B8670_ = new_B8632_ & new_B8669_;
  assign new_B8669_ = new_B8688_ | new_B8687_;
  assign new_B8668_ = ~new_B8632_ & new_B8667_;
  assign new_B8667_ = new_B8690_ | new_B8689_;
  assign new_B8666_ = new_B8632_ | new_B8665_;
  assign new_B8665_ = new_B8686_ | new_B8685_;
  assign new_B8664_ = ~new_B8644_ & ~new_B8654_;
  assign new_B8663_ = new_B8644_ & new_B8654_;
  assign new_B8662_ = ~new_B8644_ | new_B8654_;
  assign new_B8661_ = new_B8628_ & ~new_B8629_;
  assign new_B8660_ = ~new_B8628_ & new_B8629_;
  assign new_B8659_ = new_B8681_ & ~new_B8682_;
  assign new_B8658_ = ~new_B8681_ & new_B8682_;
  assign new_B8657_ = ~new_B8680_ | ~new_B8679_;
  assign new_B8656_ = new_B8672_ | new_B8671_;
  assign new_B8655_ = new_B8678_ | new_B8677_;
  assign new_B8654_ = new_B8668_ | new_B8670_;
  assign new_B8653_ = ~new_B8675_ | ~new_B8676_;
  assign new_B8652_ = new_B8628_ & ~new_B8629_;
  assign new_B8651_ = new_B8642_ & ~new_B8654_;
  assign new_B8650_ = ~new_B8642_ & new_B8654_;
  assign new_B8649_ = ~new_B8640_ & new_B8666_;
  assign new_B8648_ = new_B8664_ | new_B8663_;
  assign new_B8647_ = new_B8661_ | new_B8660_;
  assign new_B8646_ = new_B8629_ | new_B8662_;
  assign new_B8645_ = new_B8654_ & new_B8657_;
  assign new_B8644_ = new_B8659_ | new_B8658_;
  assign new_B8643_ = new_B8654_ & new_B8653_;
  assign new_B8642_ = new_B8656_ & new_B8655_;
  assign new_B8641_ = new_B8651_ | new_B8650_;
  assign new_B8640_ = new_B8629_ | new_B8652_;
  assign B8639 = new_B8640_ | new_B8649_;
  assign B8638 = new_B8647_ & new_B8648_;
  assign B8637 = new_B8647_ & new_B8646_;
  assign B8636 = new_B8645_ | new_B8644_;
  assign B8635 = new_B8643_ | new_B8642_;
  assign B8634 = new_B8641_ & new_B8640_;
  assign new_B8633_ = new_C8488_;
  assign new_B8632_ = new_C8421_;
  assign new_B8631_ = new_C8354_;
  assign new_B8630_ = new_C8287_;
  assign new_B8629_ = new_C8220_;
  assign new_B8628_ = new_C8153_;
  assign new_B8627_ = ~new_B8566_ & new_B8580_;
  assign new_B8626_ = new_B8566_ & ~new_B8580_;
  assign new_B8625_ = new_B8566_ & ~new_B8580_;
  assign new_B8624_ = ~new_B8566_ & ~new_B8580_;
  assign new_B8623_ = new_B8566_ & new_B8580_;
  assign new_B8622_ = new_B8626_ | new_B8627_;
  assign new_B8621_ = ~new_B8566_ & new_B8580_;
  assign new_B8620_ = new_B8624_ | new_B8625_;
  assign new_B8619_ = ~new_B8595_ & ~new_B8615_;
  assign new_B8618_ = new_B8595_ & new_B8615_;
  assign new_B8617_ = ~new_B8562_ | ~new_B8587_;
  assign new_B8616_ = new_B8580_ & new_B8617_;
  assign new_B8615_ = new_B8563_ | new_B8564_;
  assign new_B8614_ = new_B8563_ | new_B8580_;
  assign new_B8613_ = ~new_B8580_ & ~new_B8616_;
  assign new_B8612_ = new_B8580_ | new_B8617_;
  assign new_B8611_ = new_B8563_ & ~new_B8564_;
  assign new_B8610_ = ~new_B8563_ & new_B8564_;
  assign new_B8609_ = new_B8573_ | new_B8606_;
  assign new_B8608_ = ~new_B8573_ & ~new_B8607_;
  assign new_B8607_ = new_B8573_ & new_B8606_;
  assign new_B8606_ = ~new_B8562_ | ~new_B8587_;
  assign new_B8605_ = ~new_B8563_ & new_B8573_;
  assign new_B8604_ = new_B8563_ & ~new_B8573_;
  assign new_B8603_ = new_B8565_ & new_B8602_;
  assign new_B8602_ = new_B8621_ | new_B8620_;
  assign new_B8601_ = ~new_B8565_ & new_B8600_;
  assign new_B8600_ = new_B8623_ | new_B8622_;
  assign new_B8599_ = new_B8565_ | new_B8598_;
  assign new_B8598_ = new_B8619_ | new_B8618_;
  assign new_B8597_ = ~new_B8577_ & ~new_B8587_;
  assign new_B8596_ = new_B8577_ & new_B8587_;
  assign new_B8595_ = ~new_B8577_ | new_B8587_;
  assign new_B8594_ = new_B8561_ & ~new_B8562_;
  assign new_B8593_ = ~new_B8561_ & new_B8562_;
  assign new_B8592_ = new_B8614_ & ~new_B8615_;
  assign new_B8591_ = ~new_B8614_ & new_B8615_;
  assign new_B8590_ = ~new_B8613_ | ~new_B8612_;
  assign new_B8589_ = new_B8605_ | new_B8604_;
  assign new_B8588_ = new_B8611_ | new_B8610_;
  assign new_B8587_ = new_B8601_ | new_B8603_;
  assign new_B8586_ = ~new_B8608_ | ~new_B8609_;
  assign new_B8585_ = new_B8561_ & ~new_B8562_;
  assign new_B8584_ = new_B8575_ & ~new_B8587_;
  assign new_B8583_ = ~new_B8575_ & new_B8587_;
  assign new_B8582_ = ~new_B8573_ & new_B8599_;
  assign new_B8581_ = new_B8597_ | new_B8596_;
  assign new_B8580_ = new_B8594_ | new_B8593_;
  assign new_B8579_ = new_B8562_ | new_B8595_;
  assign new_B8578_ = new_B8587_ & new_B8590_;
  assign new_B8577_ = new_B8592_ | new_B8591_;
  assign new_B8576_ = new_B8587_ & new_B8586_;
  assign new_B8575_ = new_B8589_ & new_B8588_;
  assign new_B8574_ = new_B8584_ | new_B8583_;
  assign new_B8573_ = new_B8562_ | new_B8585_;
  assign B8572 = new_B8573_ | new_B8582_;
  assign B8571 = new_B8580_ & new_B8581_;
  assign B8570 = new_B8580_ & new_B8579_;
  assign B8569 = new_B8578_ | new_B8577_;
  assign B8568 = new_B8576_ | new_B8575_;
  assign B8567 = new_B8574_ & new_B8573_;
  assign new_B8566_ = new_C8086_;
  assign new_B8565_ = new_C8019_;
  assign new_B8564_ = new_C7952_;
  assign new_B8563_ = new_C7885_;
  assign new_B8562_ = new_C7818_;
  assign new_B8561_ = new_C7751_;
  assign new_B8560_ = ~new_B8499_ & new_B8513_;
  assign new_B8559_ = new_B8499_ & ~new_B8513_;
  assign new_B8558_ = new_B8499_ & ~new_B8513_;
  assign new_B8557_ = ~new_B8499_ & ~new_B8513_;
  assign new_B8556_ = new_B8499_ & new_B8513_;
  assign new_B8555_ = new_B8559_ | new_B8560_;
  assign new_B8554_ = ~new_B8499_ & new_B8513_;
  assign new_B8553_ = new_B8557_ | new_B8558_;
  assign new_B8552_ = ~new_B8528_ & ~new_B8548_;
  assign new_B8551_ = new_B8528_ & new_B8548_;
  assign new_B8550_ = ~new_B8495_ | ~new_B8520_;
  assign new_B8549_ = new_B8513_ & new_B8550_;
  assign new_B8548_ = new_B8496_ | new_B8497_;
  assign new_B8547_ = new_B8496_ | new_B8513_;
  assign new_B8546_ = ~new_B8513_ & ~new_B8549_;
  assign new_B8545_ = new_B8513_ | new_B8550_;
  assign new_B8544_ = new_B8496_ & ~new_B8497_;
  assign new_B8543_ = ~new_B8496_ & new_B8497_;
  assign new_B8542_ = new_B8506_ | new_B8539_;
  assign new_B8541_ = ~new_B8506_ & ~new_B8540_;
  assign new_B8540_ = new_B8506_ & new_B8539_;
  assign new_B8539_ = ~new_B8495_ | ~new_B8520_;
  assign new_B8538_ = ~new_B8496_ & new_B8506_;
  assign new_B8537_ = new_B8496_ & ~new_B8506_;
  assign new_B8536_ = new_B8498_ & new_B8535_;
  assign new_B8535_ = new_B8554_ | new_B8553_;
  assign new_B8534_ = ~new_B8498_ & new_B8533_;
  assign new_B8533_ = new_B8556_ | new_B8555_;
  assign new_B8532_ = new_B8498_ | new_B8531_;
  assign new_B8531_ = new_B8552_ | new_B8551_;
  assign new_B8530_ = ~new_B8510_ & ~new_B8520_;
  assign new_B8529_ = new_B8510_ & new_B8520_;
  assign new_B8528_ = ~new_B8510_ | new_B8520_;
  assign new_B8527_ = new_B8494_ & ~new_B8495_;
  assign new_B8526_ = ~new_B8494_ & new_B8495_;
  assign new_B8525_ = new_B8547_ & ~new_B8548_;
  assign new_B8524_ = ~new_B8547_ & new_B8548_;
  assign new_B8523_ = ~new_B8546_ | ~new_B8545_;
  assign new_B8522_ = new_B8538_ | new_B8537_;
  assign new_B8521_ = new_B8544_ | new_B8543_;
  assign new_B8520_ = new_B8534_ | new_B8536_;
  assign new_B8519_ = ~new_B8541_ | ~new_B8542_;
  assign new_B8518_ = new_B8494_ & ~new_B8495_;
  assign new_B8517_ = new_B8508_ & ~new_B8520_;
  assign new_B8516_ = ~new_B8508_ & new_B8520_;
  assign new_B8515_ = ~new_B8506_ & new_B8532_;
  assign new_B8514_ = new_B8530_ | new_B8529_;
  assign new_B8513_ = new_B8527_ | new_B8526_;
  assign new_B8512_ = new_B8495_ | new_B8528_;
  assign new_B8511_ = new_B8520_ & new_B8523_;
  assign new_B8510_ = new_B8525_ | new_B8524_;
  assign new_B8509_ = new_B8520_ & new_B8519_;
  assign new_B8508_ = new_B8522_ & new_B8521_;
  assign new_B8507_ = new_B8517_ | new_B8516_;
  assign new_B8506_ = new_B8495_ | new_B8518_;
  assign B8505 = new_B8506_ | new_B8515_;
  assign B8504 = new_B8513_ & new_B8514_;
  assign B8503 = new_B8513_ & new_B8512_;
  assign B8502 = new_B8511_ | new_B8510_;
  assign B8501 = new_B8509_ | new_B8508_;
  assign B8500 = new_B8507_ & new_B8506_;
  assign new_B8499_ = new_C7684_;
  assign new_B8498_ = new_C7617_;
  assign new_B8497_ = new_C7550_;
  assign new_B8496_ = new_C7483_;
  assign new_B8495_ = new_C7416_;
  assign new_B8494_ = new_C7349_;
  assign new_B8493_ = ~new_B8432_ & new_B8446_;
  assign new_B8492_ = new_B8432_ & ~new_B8446_;
  assign new_B8491_ = new_B8432_ & ~new_B8446_;
  assign new_B8490_ = ~new_B8432_ & ~new_B8446_;
  assign new_B8489_ = new_B8432_ & new_B8446_;
  assign new_B8488_ = new_B8492_ | new_B8493_;
  assign new_B8487_ = ~new_B8432_ & new_B8446_;
  assign new_B8486_ = new_B8490_ | new_B8491_;
  assign new_B8485_ = ~new_B8461_ & ~new_B8481_;
  assign new_B8484_ = new_B8461_ & new_B8481_;
  assign new_B8483_ = ~new_B8428_ | ~new_B8453_;
  assign new_B8482_ = new_B8446_ & new_B8483_;
  assign new_B8481_ = new_B8429_ | new_B8430_;
  assign new_B8480_ = new_B8429_ | new_B8446_;
  assign new_B8479_ = ~new_B8446_ & ~new_B8482_;
  assign new_B8478_ = new_B8446_ | new_B8483_;
  assign new_B8477_ = new_B8429_ & ~new_B8430_;
  assign new_B8476_ = ~new_B8429_ & new_B8430_;
  assign new_B8475_ = new_B8439_ | new_B8472_;
  assign new_B8474_ = ~new_B8439_ & ~new_B8473_;
  assign new_B8473_ = new_B8439_ & new_B8472_;
  assign new_B8472_ = ~new_B8428_ | ~new_B8453_;
  assign new_B8471_ = ~new_B8429_ & new_B8439_;
  assign new_B8470_ = new_B8429_ & ~new_B8439_;
  assign new_B8469_ = new_B8431_ & new_B8468_;
  assign new_B8468_ = new_B8487_ | new_B8486_;
  assign new_B8467_ = ~new_B8431_ & new_B8466_;
  assign new_B8466_ = new_B8489_ | new_B8488_;
  assign new_B8465_ = new_B8431_ | new_B8464_;
  assign new_B8464_ = new_B8485_ | new_B8484_;
  assign new_B8463_ = ~new_B8443_ & ~new_B8453_;
  assign new_B8462_ = new_B8443_ & new_B8453_;
  assign new_B8461_ = ~new_B8443_ | new_B8453_;
  assign new_B8460_ = new_B8427_ & ~new_B8428_;
  assign new_B8459_ = ~new_B8427_ & new_B8428_;
  assign new_B8458_ = new_B8480_ & ~new_B8481_;
  assign new_B8457_ = ~new_B8480_ & new_B8481_;
  assign new_B8456_ = ~new_B8479_ | ~new_B8478_;
  assign new_B8455_ = new_B8471_ | new_B8470_;
  assign new_B8454_ = new_B8477_ | new_B8476_;
  assign new_B8453_ = new_B8467_ | new_B8469_;
  assign new_B8452_ = ~new_B8474_ | ~new_B8475_;
  assign new_B8451_ = new_B8427_ & ~new_B8428_;
  assign new_B8450_ = new_B8441_ & ~new_B8453_;
  assign new_B8449_ = ~new_B8441_ & new_B8453_;
  assign new_B8448_ = ~new_B8439_ & new_B8465_;
  assign new_B8447_ = new_B8463_ | new_B8462_;
  assign new_B8446_ = new_B8460_ | new_B8459_;
  assign new_B8445_ = new_B8428_ | new_B8461_;
  assign new_B8444_ = new_B8453_ & new_B8456_;
  assign new_B8443_ = new_B8458_ | new_B8457_;
  assign new_B8442_ = new_B8453_ & new_B8452_;
  assign new_B8441_ = new_B8455_ & new_B8454_;
  assign new_B8440_ = new_B8450_ | new_B8449_;
  assign new_B8439_ = new_B8428_ | new_B8451_;
  assign B8438 = new_B8439_ | new_B8448_;
  assign B8437 = new_B8446_ & new_B8447_;
  assign B8436 = new_B8446_ & new_B8445_;
  assign B8435 = new_B8444_ | new_B8443_;
  assign B8434 = new_B8442_ | new_B8441_;
  assign B8433 = new_B8440_ & new_B8439_;
  assign new_B8432_ = new_C7282_;
  assign new_B8431_ = new_C7215_;
  assign new_B8430_ = new_C7148_;
  assign new_B8429_ = new_C7081_;
  assign new_B8428_ = new_C7014_;
  assign new_B8427_ = new_C6947_;
  assign new_B8426_ = ~new_B8365_ & new_B8379_;
  assign new_B8425_ = new_B8365_ & ~new_B8379_;
  assign new_B8424_ = new_B8365_ & ~new_B8379_;
  assign new_B8423_ = ~new_B8365_ & ~new_B8379_;
  assign new_B8422_ = new_B8365_ & new_B8379_;
  assign new_B8421_ = new_B8425_ | new_B8426_;
  assign new_B8420_ = ~new_B8365_ & new_B8379_;
  assign new_B8419_ = new_B8423_ | new_B8424_;
  assign new_B8418_ = ~new_B8394_ & ~new_B8414_;
  assign new_B8417_ = new_B8394_ & new_B8414_;
  assign new_B8416_ = ~new_B8361_ | ~new_B8386_;
  assign new_B8415_ = new_B8379_ & new_B8416_;
  assign new_B8414_ = new_B8362_ | new_B8363_;
  assign new_B8413_ = new_B8362_ | new_B8379_;
  assign new_B8412_ = ~new_B8379_ & ~new_B8415_;
  assign new_B8411_ = new_B8379_ | new_B8416_;
  assign new_B8410_ = new_B8362_ & ~new_B8363_;
  assign new_B8409_ = ~new_B8362_ & new_B8363_;
  assign new_B8408_ = new_B8372_ | new_B8405_;
  assign new_B8407_ = ~new_B8372_ & ~new_B8406_;
  assign new_B8406_ = new_B8372_ & new_B8405_;
  assign new_B8405_ = ~new_B8361_ | ~new_B8386_;
  assign new_B8404_ = ~new_B8362_ & new_B8372_;
  assign new_B8403_ = new_B8362_ & ~new_B8372_;
  assign new_B8402_ = new_B8364_ & new_B8401_;
  assign new_B8401_ = new_B8420_ | new_B8419_;
  assign new_B8400_ = ~new_B8364_ & new_B8399_;
  assign new_B8399_ = new_B8422_ | new_B8421_;
  assign new_B8398_ = new_B8364_ | new_B8397_;
  assign new_B8397_ = new_B8418_ | new_B8417_;
  assign new_B8396_ = ~new_B8376_ & ~new_B8386_;
  assign new_B8395_ = new_B8376_ & new_B8386_;
  assign new_B8394_ = ~new_B8376_ | new_B8386_;
  assign new_B8393_ = new_B8360_ & ~new_B8361_;
  assign new_B8392_ = ~new_B8360_ & new_B8361_;
  assign new_B8391_ = new_B8413_ & ~new_B8414_;
  assign new_B8390_ = ~new_B8413_ & new_B8414_;
  assign new_B8389_ = ~new_B8412_ | ~new_B8411_;
  assign new_B8388_ = new_B8404_ | new_B8403_;
  assign new_B8387_ = new_B8410_ | new_B8409_;
  assign new_B8386_ = new_B8400_ | new_B8402_;
  assign new_B8385_ = ~new_B8407_ | ~new_B8408_;
  assign new_B8384_ = new_B8360_ & ~new_B8361_;
  assign new_B8383_ = new_B8374_ & ~new_B8386_;
  assign new_B8382_ = ~new_B8374_ & new_B8386_;
  assign new_B8381_ = ~new_B8372_ & new_B8398_;
  assign new_B8380_ = new_B8396_ | new_B8395_;
  assign new_B8379_ = new_B8393_ | new_B8392_;
  assign new_B8378_ = new_B8361_ | new_B8394_;
  assign new_B8377_ = new_B8386_ & new_B8389_;
  assign new_B8376_ = new_B8391_ | new_B8390_;
  assign new_B8375_ = new_B8386_ & new_B8385_;
  assign new_B8374_ = new_B8388_ & new_B8387_;
  assign new_B8373_ = new_B8383_ | new_B8382_;
  assign new_B8372_ = new_B8361_ | new_B8384_;
  assign B8371 = new_B8372_ | new_B8381_;
  assign B8370 = new_B8379_ & new_B8380_;
  assign B8369 = new_B8379_ & new_B8378_;
  assign B8368 = new_B8377_ | new_B8376_;
  assign B8367 = new_B8375_ | new_B8374_;
  assign B8366 = new_B8373_ & new_B8372_;
  assign new_B8365_ = new_C6880_;
  assign new_B8364_ = new_C6813_;
  assign new_B8363_ = new_C6746_;
  assign new_B8362_ = new_C6679_;
  assign new_B8361_ = new_C6612_;
  assign new_B8360_ = new_C6545_;
  assign new_B8359_ = ~new_B8298_ & new_B8312_;
  assign new_B8358_ = new_B8298_ & ~new_B8312_;
  assign new_B8357_ = new_B8298_ & ~new_B8312_;
  assign new_B8356_ = ~new_B8298_ & ~new_B8312_;
  assign new_B8355_ = new_B8298_ & new_B8312_;
  assign new_B8354_ = new_B8358_ | new_B8359_;
  assign new_B8353_ = ~new_B8298_ & new_B8312_;
  assign new_B8352_ = new_B8356_ | new_B8357_;
  assign new_B8351_ = ~new_B8327_ & ~new_B8347_;
  assign new_B8350_ = new_B8327_ & new_B8347_;
  assign new_B8349_ = ~new_B8294_ | ~new_B8319_;
  assign new_B8348_ = new_B8312_ & new_B8349_;
  assign new_B8347_ = new_B8295_ | new_B8296_;
  assign new_B8346_ = new_B8295_ | new_B8312_;
  assign new_B8345_ = ~new_B8312_ & ~new_B8348_;
  assign new_B8344_ = new_B8312_ | new_B8349_;
  assign new_B8343_ = new_B8295_ & ~new_B8296_;
  assign new_B8342_ = ~new_B8295_ & new_B8296_;
  assign new_B8341_ = new_B8305_ | new_B8338_;
  assign new_B8340_ = ~new_B8305_ & ~new_B8339_;
  assign new_B8339_ = new_B8305_ & new_B8338_;
  assign new_B8338_ = ~new_B8294_ | ~new_B8319_;
  assign new_B8337_ = ~new_B8295_ & new_B8305_;
  assign new_B8336_ = new_B8295_ & ~new_B8305_;
  assign new_B8335_ = new_B8297_ & new_B8334_;
  assign new_B8334_ = new_B8353_ | new_B8352_;
  assign new_B8333_ = ~new_B8297_ & new_B8332_;
  assign new_B8332_ = new_B8355_ | new_B8354_;
  assign new_B8331_ = new_B8297_ | new_B8330_;
  assign new_B8330_ = new_B8351_ | new_B8350_;
  assign new_B8329_ = ~new_B8309_ & ~new_B8319_;
  assign new_B8328_ = new_B8309_ & new_B8319_;
  assign new_B8327_ = ~new_B8309_ | new_B8319_;
  assign new_B8326_ = new_B8293_ & ~new_B8294_;
  assign new_B8325_ = ~new_B8293_ & new_B8294_;
  assign new_B8324_ = new_B8346_ & ~new_B8347_;
  assign new_B8323_ = ~new_B8346_ & new_B8347_;
  assign new_B8322_ = ~new_B8345_ | ~new_B8344_;
  assign new_B8321_ = new_B8337_ | new_B8336_;
  assign new_B8320_ = new_B8343_ | new_B8342_;
  assign new_B8319_ = new_B8333_ | new_B8335_;
  assign new_B8318_ = ~new_B8340_ | ~new_B8341_;
  assign new_B8317_ = new_B8293_ & ~new_B8294_;
  assign new_B8316_ = new_B8307_ & ~new_B8319_;
  assign new_B8315_ = ~new_B8307_ & new_B8319_;
  assign new_B8314_ = ~new_B8305_ & new_B8331_;
  assign new_B8313_ = new_B8329_ | new_B8328_;
  assign new_B8312_ = new_B8326_ | new_B8325_;
  assign new_B8311_ = new_B8294_ | new_B8327_;
  assign new_B8310_ = new_B8319_ & new_B8322_;
  assign new_B8309_ = new_B8324_ | new_B8323_;
  assign new_B8308_ = new_B8319_ & new_B8318_;
  assign new_B8307_ = new_B8321_ & new_B8320_;
  assign new_B8306_ = new_B8316_ | new_B8315_;
  assign new_B8305_ = new_B8294_ | new_B8317_;
  assign B8304 = new_B8305_ | new_B8314_;
  assign B8303 = new_B8312_ & new_B8313_;
  assign B8302 = new_B8312_ & new_B8311_;
  assign B8301 = new_B8310_ | new_B8309_;
  assign B8300 = new_B8308_ | new_B8307_;
  assign B8299 = new_B8306_ & new_B8305_;
  assign new_B8298_ = new_C6478_;
  assign new_B8297_ = new_C6411_;
  assign new_B8296_ = new_C6344_;
  assign new_B8295_ = new_C6277_;
  assign new_B8294_ = new_C6210_;
  assign new_B8293_ = new_C6143_;
  assign new_B8292_ = ~new_B8231_ & new_B8245_;
  assign new_B8291_ = new_B8231_ & ~new_B8245_;
  assign new_B8290_ = new_B8231_ & ~new_B8245_;
  assign new_B8289_ = ~new_B8231_ & ~new_B8245_;
  assign new_B8288_ = new_B8231_ & new_B8245_;
  assign new_B8287_ = new_B8291_ | new_B8292_;
  assign new_B8286_ = ~new_B8231_ & new_B8245_;
  assign new_B8285_ = new_B8289_ | new_B8290_;
  assign new_B8284_ = ~new_B8260_ & ~new_B8280_;
  assign new_B8283_ = new_B8260_ & new_B8280_;
  assign new_B8282_ = ~new_B8227_ | ~new_B8252_;
  assign new_B8281_ = new_B8245_ & new_B8282_;
  assign new_B8280_ = new_B8228_ | new_B8229_;
  assign new_B8279_ = new_B8228_ | new_B8245_;
  assign new_B8278_ = ~new_B8245_ & ~new_B8281_;
  assign new_B8277_ = new_B8245_ | new_B8282_;
  assign new_B8276_ = new_B8228_ & ~new_B8229_;
  assign new_B8275_ = ~new_B8228_ & new_B8229_;
  assign new_B8274_ = new_B8238_ | new_B8271_;
  assign new_B8273_ = ~new_B8238_ & ~new_B8272_;
  assign new_B8272_ = new_B8238_ & new_B8271_;
  assign new_B8271_ = ~new_B8227_ | ~new_B8252_;
  assign new_B8270_ = ~new_B8228_ & new_B8238_;
  assign new_B8269_ = new_B8228_ & ~new_B8238_;
  assign new_B8268_ = new_B8230_ & new_B8267_;
  assign new_B8267_ = new_B8286_ | new_B8285_;
  assign new_B8266_ = ~new_B8230_ & new_B8265_;
  assign new_B8265_ = new_B8288_ | new_B8287_;
  assign new_B8264_ = new_B8230_ | new_B8263_;
  assign new_B8263_ = new_B8284_ | new_B8283_;
  assign new_B8262_ = ~new_B8242_ & ~new_B8252_;
  assign new_B8261_ = new_B8242_ & new_B8252_;
  assign new_B8260_ = ~new_B8242_ | new_B8252_;
  assign new_B8259_ = new_B8226_ & ~new_B8227_;
  assign new_B8258_ = ~new_B8226_ & new_B8227_;
  assign new_B8257_ = new_B8279_ & ~new_B8280_;
  assign new_B8256_ = ~new_B8279_ & new_B8280_;
  assign new_B8255_ = ~new_B8278_ | ~new_B8277_;
  assign new_B8254_ = new_B8270_ | new_B8269_;
  assign new_B8253_ = new_B8276_ | new_B8275_;
  assign new_B8252_ = new_B8266_ | new_B8268_;
  assign new_B8251_ = ~new_B8273_ | ~new_B8274_;
  assign new_B8250_ = new_B8226_ & ~new_B8227_;
  assign new_B8249_ = new_B8240_ & ~new_B8252_;
  assign new_B8248_ = ~new_B8240_ & new_B8252_;
  assign new_B8247_ = ~new_B8238_ & new_B8264_;
  assign new_B8246_ = new_B8262_ | new_B8261_;
  assign new_B8245_ = new_B8259_ | new_B8258_;
  assign new_B8244_ = new_B8227_ | new_B8260_;
  assign new_B8243_ = new_B8252_ & new_B8255_;
  assign new_B8242_ = new_B8257_ | new_B8256_;
  assign new_B8241_ = new_B8252_ & new_B8251_;
  assign new_B8240_ = new_B8254_ & new_B8253_;
  assign new_B8239_ = new_B8249_ | new_B8248_;
  assign new_B8238_ = new_B8227_ | new_B8250_;
  assign B8237 = new_B8238_ | new_B8247_;
  assign B8236 = new_B8245_ & new_B8246_;
  assign B8235 = new_B8245_ & new_B8244_;
  assign B8234 = new_B8243_ | new_B8242_;
  assign B8233 = new_B8241_ | new_B8240_;
  assign B8232 = new_B8239_ & new_B8238_;
  assign new_B8231_ = new_C6076_;
  assign new_B8230_ = new_C6009_;
  assign new_B8229_ = new_C5942_;
  assign new_B8228_ = new_C5875_;
  assign new_B8227_ = new_C5808_;
  assign new_B8226_ = new_C5741_;
  assign new_B8225_ = ~new_B8164_ & new_B8178_;
  assign new_B8224_ = new_B8164_ & ~new_B8178_;
  assign new_B8223_ = new_B8164_ & ~new_B8178_;
  assign new_B8222_ = ~new_B8164_ & ~new_B8178_;
  assign new_B8221_ = new_B8164_ & new_B8178_;
  assign new_B8220_ = new_B8224_ | new_B8225_;
  assign new_B8219_ = ~new_B8164_ & new_B8178_;
  assign new_B8218_ = new_B8222_ | new_B8223_;
  assign new_B8217_ = ~new_B8193_ & ~new_B8213_;
  assign new_B8216_ = new_B8193_ & new_B8213_;
  assign new_B8215_ = ~new_B8160_ | ~new_B8185_;
  assign new_B8214_ = new_B8178_ & new_B8215_;
  assign new_B8213_ = new_B8161_ | new_B8162_;
  assign new_B8212_ = new_B8161_ | new_B8178_;
  assign new_B8211_ = ~new_B8178_ & ~new_B8214_;
  assign new_B8210_ = new_B8178_ | new_B8215_;
  assign new_B8209_ = new_B8161_ & ~new_B8162_;
  assign new_B8208_ = ~new_B8161_ & new_B8162_;
  assign new_B8207_ = new_B8171_ | new_B8204_;
  assign new_B8206_ = ~new_B8171_ & ~new_B8205_;
  assign new_B8205_ = new_B8171_ & new_B8204_;
  assign new_B8204_ = ~new_B8160_ | ~new_B8185_;
  assign new_B8203_ = ~new_B8161_ & new_B8171_;
  assign new_B8202_ = new_B8161_ & ~new_B8171_;
  assign new_B8201_ = new_B8163_ & new_B8200_;
  assign new_B8200_ = new_B8219_ | new_B8218_;
  assign new_B8199_ = ~new_B8163_ & new_B8198_;
  assign new_B8198_ = new_B8221_ | new_B8220_;
  assign new_B8197_ = new_B8163_ | new_B8196_;
  assign new_B8196_ = new_B8217_ | new_B8216_;
  assign new_B8195_ = ~new_B8175_ & ~new_B8185_;
  assign new_B8194_ = new_B8175_ & new_B8185_;
  assign new_B8193_ = ~new_B8175_ | new_B8185_;
  assign new_B8192_ = new_B8159_ & ~new_B8160_;
  assign new_B8191_ = ~new_B8159_ & new_B8160_;
  assign new_B8190_ = new_B8212_ & ~new_B8213_;
  assign new_B8189_ = ~new_B8212_ & new_B8213_;
  assign new_B8188_ = ~new_B8211_ | ~new_B8210_;
  assign new_B8187_ = new_B8203_ | new_B8202_;
  assign new_B8186_ = new_B8209_ | new_B8208_;
  assign new_B8185_ = new_B8199_ | new_B8201_;
  assign new_B8184_ = ~new_B8206_ | ~new_B8207_;
  assign new_B8183_ = new_B8159_ & ~new_B8160_;
  assign new_B8182_ = new_B8173_ & ~new_B8185_;
  assign new_B8181_ = ~new_B8173_ & new_B8185_;
  assign new_B8180_ = ~new_B8171_ & new_B8197_;
  assign new_B8179_ = new_B8195_ | new_B8194_;
  assign new_B8178_ = new_B8192_ | new_B8191_;
  assign new_B8177_ = new_B8160_ | new_B8193_;
  assign new_B8176_ = new_B8185_ & new_B8188_;
  assign new_B8175_ = new_B8190_ | new_B8189_;
  assign new_B8174_ = new_B8185_ & new_B8184_;
  assign new_B8173_ = new_B8187_ & new_B8186_;
  assign new_B8172_ = new_B8182_ | new_B8181_;
  assign new_B8171_ = new_B8160_ | new_B8183_;
  assign B8170 = new_B8171_ | new_B8180_;
  assign B8169 = new_B8178_ & new_B8179_;
  assign B8168 = new_B8178_ & new_B8177_;
  assign B8167 = new_B8176_ | new_B8175_;
  assign B8166 = new_B8174_ | new_B8173_;
  assign B8165 = new_B8172_ & new_B8171_;
  assign new_B8164_ = new_C5674_;
  assign new_B8163_ = new_C5607_;
  assign new_B8162_ = new_C5540_;
  assign new_B8161_ = new_C5473_;
  assign new_B8160_ = new_C5406_;
  assign new_B8159_ = new_C5339_;
  assign new_B8158_ = ~new_B8097_ & new_B8111_;
  assign new_B8157_ = new_B8097_ & ~new_B8111_;
  assign new_B8156_ = new_B8097_ & ~new_B8111_;
  assign new_B8155_ = ~new_B8097_ & ~new_B8111_;
  assign new_B8154_ = new_B8097_ & new_B8111_;
  assign new_B8153_ = new_B8157_ | new_B8158_;
  assign new_B8152_ = ~new_B8097_ & new_B8111_;
  assign new_B8151_ = new_B8155_ | new_B8156_;
  assign new_B8150_ = ~new_B8126_ & ~new_B8146_;
  assign new_B8149_ = new_B8126_ & new_B8146_;
  assign new_B8148_ = ~new_B8093_ | ~new_B8118_;
  assign new_B8147_ = new_B8111_ & new_B8148_;
  assign new_B8146_ = new_B8094_ | new_B8095_;
  assign new_B8145_ = new_B8094_ | new_B8111_;
  assign new_B8144_ = ~new_B8111_ & ~new_B8147_;
  assign new_B8143_ = new_B8111_ | new_B8148_;
  assign new_B8142_ = new_B8094_ & ~new_B8095_;
  assign new_B8141_ = ~new_B8094_ & new_B8095_;
  assign new_B8140_ = new_B8104_ | new_B8137_;
  assign new_B8139_ = ~new_B8104_ & ~new_B8138_;
  assign new_B8138_ = new_B8104_ & new_B8137_;
  assign new_B8137_ = ~new_B8093_ | ~new_B8118_;
  assign new_B8136_ = ~new_B8094_ & new_B8104_;
  assign new_B8135_ = new_B8094_ & ~new_B8104_;
  assign new_B8134_ = new_B8096_ & new_B8133_;
  assign new_B8133_ = new_B8152_ | new_B8151_;
  assign new_B8132_ = ~new_B8096_ & new_B8131_;
  assign new_B8131_ = new_B8154_ | new_B8153_;
  assign new_B8130_ = new_B8096_ | new_B8129_;
  assign new_B8129_ = new_B8150_ | new_B8149_;
  assign new_B8128_ = ~new_B8108_ & ~new_B8118_;
  assign new_B8127_ = new_B8108_ & new_B8118_;
  assign new_B8126_ = ~new_B8108_ | new_B8118_;
  assign new_B8125_ = new_B8092_ & ~new_B8093_;
  assign new_B8124_ = ~new_B8092_ & new_B8093_;
  assign new_B8123_ = new_B8145_ & ~new_B8146_;
  assign new_B8122_ = ~new_B8145_ & new_B8146_;
  assign new_B8121_ = ~new_B8144_ | ~new_B8143_;
  assign new_B8120_ = new_B8136_ | new_B8135_;
  assign new_B8119_ = new_B8142_ | new_B8141_;
  assign new_B8118_ = new_B8132_ | new_B8134_;
  assign new_B8117_ = ~new_B8139_ | ~new_B8140_;
  assign new_B8116_ = new_B8092_ & ~new_B8093_;
  assign new_B8115_ = new_B8106_ & ~new_B8118_;
  assign new_B8114_ = ~new_B8106_ & new_B8118_;
  assign new_B8113_ = ~new_B8104_ & new_B8130_;
  assign new_B8112_ = new_B8128_ | new_B8127_;
  assign new_B8111_ = new_B8125_ | new_B8124_;
  assign new_B8110_ = new_B8093_ | new_B8126_;
  assign new_B8109_ = new_B8118_ & new_B8121_;
  assign new_B8108_ = new_B8123_ | new_B8122_;
  assign new_B8107_ = new_B8118_ & new_B8117_;
  assign new_B8106_ = new_B8120_ & new_B8119_;
  assign new_B8105_ = new_B8115_ | new_B8114_;
  assign new_B8104_ = new_B8093_ | new_B8116_;
  assign B8103 = new_B8104_ | new_B8113_;
  assign B8102 = new_B8111_ & new_B8112_;
  assign B8101 = new_B8111_ & new_B8110_;
  assign B8100 = new_B8109_ | new_B8108_;
  assign B8099 = new_B8107_ | new_B8106_;
  assign B8098 = new_B8105_ & new_B8104_;
  assign new_B8097_ = new_C5272_;
  assign new_B8096_ = new_C5205_;
  assign new_B8095_ = new_C5138_;
  assign new_B8094_ = new_C5071_;
  assign new_B8093_ = new_C5004_;
  assign new_B8092_ = new_C4937_;
  assign new_B8091_ = ~new_B8030_ & new_B8044_;
  assign new_B8090_ = new_B8030_ & ~new_B8044_;
  assign new_B8089_ = new_B8030_ & ~new_B8044_;
  assign new_B8088_ = ~new_B8030_ & ~new_B8044_;
  assign new_B8087_ = new_B8030_ & new_B8044_;
  assign new_B8086_ = new_B8090_ | new_B8091_;
  assign new_B8085_ = ~new_B8030_ & new_B8044_;
  assign new_B8084_ = new_B8088_ | new_B8089_;
  assign new_B8083_ = ~new_B8059_ & ~new_B8079_;
  assign new_B8082_ = new_B8059_ & new_B8079_;
  assign new_B8081_ = ~new_B8026_ | ~new_B8051_;
  assign new_B8080_ = new_B8044_ & new_B8081_;
  assign new_B8079_ = new_B8027_ | new_B8028_;
  assign new_B8078_ = new_B8027_ | new_B8044_;
  assign new_B8077_ = ~new_B8044_ & ~new_B8080_;
  assign new_B8076_ = new_B8044_ | new_B8081_;
  assign new_B8075_ = new_B8027_ & ~new_B8028_;
  assign new_B8074_ = ~new_B8027_ & new_B8028_;
  assign new_B8073_ = new_B8037_ | new_B8070_;
  assign new_B8072_ = ~new_B8037_ & ~new_B8071_;
  assign new_B8071_ = new_B8037_ & new_B8070_;
  assign new_B8070_ = ~new_B8026_ | ~new_B8051_;
  assign new_B8069_ = ~new_B8027_ & new_B8037_;
  assign new_B8068_ = new_B8027_ & ~new_B8037_;
  assign new_B8067_ = new_B8029_ & new_B8066_;
  assign new_B8066_ = new_B8085_ | new_B8084_;
  assign new_B8065_ = ~new_B8029_ & new_B8064_;
  assign new_B8064_ = new_B8087_ | new_B8086_;
  assign new_B8063_ = new_B8029_ | new_B8062_;
  assign new_B8062_ = new_B8083_ | new_B8082_;
  assign new_B8061_ = ~new_B8041_ & ~new_B8051_;
  assign new_B8060_ = new_B8041_ & new_B8051_;
  assign new_B8059_ = ~new_B8041_ | new_B8051_;
  assign new_B8058_ = new_B8025_ & ~new_B8026_;
  assign new_B8057_ = ~new_B8025_ & new_B8026_;
  assign new_B8056_ = new_B8078_ & ~new_B8079_;
  assign new_B8055_ = ~new_B8078_ & new_B8079_;
  assign new_B8054_ = ~new_B8077_ | ~new_B8076_;
  assign new_B8053_ = new_B8069_ | new_B8068_;
  assign new_B8052_ = new_B8075_ | new_B8074_;
  assign new_B8051_ = new_B8065_ | new_B8067_;
  assign new_B8050_ = ~new_B8072_ | ~new_B8073_;
  assign new_B8049_ = new_B8025_ & ~new_B8026_;
  assign new_B8048_ = new_B8039_ & ~new_B8051_;
  assign new_B8047_ = ~new_B8039_ & new_B8051_;
  assign new_B8046_ = ~new_B8037_ & new_B8063_;
  assign new_B8045_ = new_B8061_ | new_B8060_;
  assign new_B8044_ = new_B8058_ | new_B8057_;
  assign new_B8043_ = new_B8026_ | new_B8059_;
  assign new_B8042_ = new_B8051_ & new_B8054_;
  assign new_B8041_ = new_B8056_ | new_B8055_;
  assign new_B8040_ = new_B8051_ & new_B8050_;
  assign new_B8039_ = new_B8053_ & new_B8052_;
  assign new_B8038_ = new_B8048_ | new_B8047_;
  assign new_B8037_ = new_B8026_ | new_B8049_;
  assign B8036 = new_B8037_ | new_B8046_;
  assign B8035 = new_B8044_ & new_B8045_;
  assign B8034 = new_B8044_ & new_B8043_;
  assign B8033 = new_B8042_ | new_B8041_;
  assign B8032 = new_B8040_ | new_B8039_;
  assign B8031 = new_B8038_ & new_B8037_;
  assign new_B8030_ = new_C4870_;
  assign new_B8029_ = new_C4803_;
  assign new_B8028_ = new_C4736_;
  assign new_B8027_ = new_C4669_;
  assign new_B8026_ = new_C4602_;
  assign new_B8025_ = new_C4535_;
  assign new_B8024_ = ~new_B7963_ & new_B7977_;
  assign new_B8023_ = new_B7963_ & ~new_B7977_;
  assign new_B8022_ = new_B7963_ & ~new_B7977_;
  assign new_B8021_ = ~new_B7963_ & ~new_B7977_;
  assign new_B8020_ = new_B7963_ & new_B7977_;
  assign new_B8019_ = new_B8023_ | new_B8024_;
  assign new_B8018_ = ~new_B7963_ & new_B7977_;
  assign new_B8017_ = new_B8021_ | new_B8022_;
  assign new_B8016_ = ~new_B7992_ & ~new_B8012_;
  assign new_B8015_ = new_B7992_ & new_B8012_;
  assign new_B8014_ = ~new_B7959_ | ~new_B7984_;
  assign new_B8013_ = new_B7977_ & new_B8014_;
  assign new_B8012_ = new_B7960_ | new_B7961_;
  assign new_B8011_ = new_B7960_ | new_B7977_;
  assign new_B8010_ = ~new_B7977_ & ~new_B8013_;
  assign new_B8009_ = new_B7977_ | new_B8014_;
  assign new_B8008_ = new_B7960_ & ~new_B7961_;
  assign new_B8007_ = ~new_B7960_ & new_B7961_;
  assign new_B8006_ = new_B7970_ | new_B8003_;
  assign new_B8005_ = ~new_B7970_ & ~new_B8004_;
  assign new_B8004_ = new_B7970_ & new_B8003_;
  assign new_B8003_ = ~new_B7959_ | ~new_B7984_;
  assign new_B8002_ = ~new_B7960_ & new_B7970_;
  assign new_B8001_ = new_B7960_ & ~new_B7970_;
  assign new_B8000_ = new_B7962_ & new_B7999_;
  assign new_B7999_ = new_B8018_ | new_B8017_;
  assign new_B7998_ = ~new_B7962_ & new_B7997_;
  assign new_B7997_ = new_B8020_ | new_B8019_;
  assign new_B7996_ = new_B7962_ | new_B7995_;
  assign new_B7995_ = new_B8016_ | new_B8015_;
  assign new_B7994_ = ~new_B7974_ & ~new_B7984_;
  assign new_B7993_ = new_B7974_ & new_B7984_;
  assign new_B7992_ = ~new_B7974_ | new_B7984_;
  assign new_B7991_ = new_B7958_ & ~new_B7959_;
  assign new_B7990_ = ~new_B7958_ & new_B7959_;
  assign new_B7989_ = new_B8011_ & ~new_B8012_;
  assign new_B7988_ = ~new_B8011_ & new_B8012_;
  assign new_B7987_ = ~new_B8010_ | ~new_B8009_;
  assign new_B7986_ = new_B8002_ | new_B8001_;
  assign new_B7985_ = new_B8008_ | new_B8007_;
  assign new_B7984_ = new_B7998_ | new_B8000_;
  assign new_B7983_ = ~new_B8005_ | ~new_B8006_;
  assign new_B7982_ = new_B7958_ & ~new_B7959_;
  assign new_B7981_ = new_B7972_ & ~new_B7984_;
  assign new_B7980_ = ~new_B7972_ & new_B7984_;
  assign new_B7979_ = ~new_B7970_ & new_B7996_;
  assign new_B7978_ = new_B7994_ | new_B7993_;
  assign new_B7977_ = new_B7991_ | new_B7990_;
  assign new_B7976_ = new_B7959_ | new_B7992_;
  assign new_B7975_ = new_B7984_ & new_B7987_;
  assign new_B7974_ = new_B7989_ | new_B7988_;
  assign new_B7973_ = new_B7984_ & new_B7983_;
  assign new_B7972_ = new_B7986_ & new_B7985_;
  assign new_B7971_ = new_B7981_ | new_B7980_;
  assign new_B7970_ = new_B7959_ | new_B7982_;
  assign B7969 = new_B7970_ | new_B7979_;
  assign B7968 = new_B7977_ & new_B7978_;
  assign B7967 = new_B7977_ & new_B7976_;
  assign B7966 = new_B7975_ | new_B7974_;
  assign B7965 = new_B7973_ | new_B7972_;
  assign B7964 = new_B7971_ & new_B7970_;
  assign new_B7963_ = new_C4468_;
  assign new_B7962_ = new_C4401_;
  assign new_B7961_ = new_C4334_;
  assign new_B7960_ = new_C4267_;
  assign new_B7959_ = new_C4200_;
  assign new_B7958_ = new_C4133_;
  assign new_B7957_ = ~new_B7896_ & new_B7910_;
  assign new_B7956_ = new_B7896_ & ~new_B7910_;
  assign new_B7955_ = new_B7896_ & ~new_B7910_;
  assign new_B7954_ = ~new_B7896_ & ~new_B7910_;
  assign new_B7953_ = new_B7896_ & new_B7910_;
  assign new_B7952_ = new_B7956_ | new_B7957_;
  assign new_B7951_ = ~new_B7896_ & new_B7910_;
  assign new_B7950_ = new_B7954_ | new_B7955_;
  assign new_B7949_ = ~new_B7925_ & ~new_B7945_;
  assign new_B7948_ = new_B7925_ & new_B7945_;
  assign new_B7947_ = ~new_B7892_ | ~new_B7917_;
  assign new_B7946_ = new_B7910_ & new_B7947_;
  assign new_B7945_ = new_B7893_ | new_B7894_;
  assign new_B7944_ = new_B7893_ | new_B7910_;
  assign new_B7943_ = ~new_B7910_ & ~new_B7946_;
  assign new_B7942_ = new_B7910_ | new_B7947_;
  assign new_B7941_ = new_B7893_ & ~new_B7894_;
  assign new_B7940_ = ~new_B7893_ & new_B7894_;
  assign new_B7939_ = new_B7903_ | new_B7936_;
  assign new_B7938_ = ~new_B7903_ & ~new_B7937_;
  assign new_B7937_ = new_B7903_ & new_B7936_;
  assign new_B7936_ = ~new_B7892_ | ~new_B7917_;
  assign new_B7935_ = ~new_B7893_ & new_B7903_;
  assign new_B7934_ = new_B7893_ & ~new_B7903_;
  assign new_B7933_ = new_B7895_ & new_B7932_;
  assign new_B7932_ = new_B7951_ | new_B7950_;
  assign new_B7931_ = ~new_B7895_ & new_B7930_;
  assign new_B7930_ = new_B7953_ | new_B7952_;
  assign new_B7929_ = new_B7895_ | new_B7928_;
  assign new_B7928_ = new_B7949_ | new_B7948_;
  assign new_B7927_ = ~new_B7907_ & ~new_B7917_;
  assign new_B7926_ = new_B7907_ & new_B7917_;
  assign new_B7925_ = ~new_B7907_ | new_B7917_;
  assign new_B7924_ = new_B7891_ & ~new_B7892_;
  assign new_B7923_ = ~new_B7891_ & new_B7892_;
  assign new_B7922_ = new_B7944_ & ~new_B7945_;
  assign new_B7921_ = ~new_B7944_ & new_B7945_;
  assign new_B7920_ = ~new_B7943_ | ~new_B7942_;
  assign new_B7919_ = new_B7935_ | new_B7934_;
  assign new_B7918_ = new_B7941_ | new_B7940_;
  assign new_B7917_ = new_B7931_ | new_B7933_;
  assign new_B7916_ = ~new_B7938_ | ~new_B7939_;
  assign new_B7915_ = new_B7891_ & ~new_B7892_;
  assign new_B7914_ = new_B7905_ & ~new_B7917_;
  assign new_B7913_ = ~new_B7905_ & new_B7917_;
  assign new_B7912_ = ~new_B7903_ & new_B7929_;
  assign new_B7911_ = new_B7927_ | new_B7926_;
  assign new_B7910_ = new_B7924_ | new_B7923_;
  assign new_B7909_ = new_B7892_ | new_B7925_;
  assign new_B7908_ = new_B7917_ & new_B7920_;
  assign new_B7907_ = new_B7922_ | new_B7921_;
  assign new_B7906_ = new_B7917_ & new_B7916_;
  assign new_B7905_ = new_B7919_ & new_B7918_;
  assign new_B7904_ = new_B7914_ | new_B7913_;
  assign new_B7903_ = new_B7892_ | new_B7915_;
  assign B7902 = new_B7903_ | new_B7912_;
  assign B7901 = new_B7910_ & new_B7911_;
  assign B7900 = new_B7910_ & new_B7909_;
  assign B7899 = new_B7908_ | new_B7907_;
  assign B7898 = new_B7906_ | new_B7905_;
  assign B7897 = new_B7904_ & new_B7903_;
  assign new_B7896_ = new_C4066_;
  assign new_B7895_ = new_C3999_;
  assign new_B7894_ = new_C3932_;
  assign new_B7893_ = new_C3865_;
  assign new_B7892_ = new_C3798_;
  assign new_B7891_ = new_C3731_;
  assign new_B7890_ = ~new_B7829_ & new_B7843_;
  assign new_B7889_ = new_B7829_ & ~new_B7843_;
  assign new_B7888_ = new_B7829_ & ~new_B7843_;
  assign new_B7887_ = ~new_B7829_ & ~new_B7843_;
  assign new_B7886_ = new_B7829_ & new_B7843_;
  assign new_B7885_ = new_B7889_ | new_B7890_;
  assign new_B7884_ = ~new_B7829_ & new_B7843_;
  assign new_B7883_ = new_B7887_ | new_B7888_;
  assign new_B7882_ = ~new_B7858_ & ~new_B7878_;
  assign new_B7881_ = new_B7858_ & new_B7878_;
  assign new_B7880_ = ~new_B7825_ | ~new_B7850_;
  assign new_B7879_ = new_B7843_ & new_B7880_;
  assign new_B7878_ = new_B7826_ | new_B7827_;
  assign new_B7877_ = new_B7826_ | new_B7843_;
  assign new_B7876_ = ~new_B7843_ & ~new_B7879_;
  assign new_B7875_ = new_B7843_ | new_B7880_;
  assign new_B7874_ = new_B7826_ & ~new_B7827_;
  assign new_B7873_ = ~new_B7826_ & new_B7827_;
  assign new_B7872_ = new_B7836_ | new_B7869_;
  assign new_B7871_ = ~new_B7836_ & ~new_B7870_;
  assign new_B7870_ = new_B7836_ & new_B7869_;
  assign new_B7869_ = ~new_B7825_ | ~new_B7850_;
  assign new_B7868_ = ~new_B7826_ & new_B7836_;
  assign new_B7867_ = new_B7826_ & ~new_B7836_;
  assign new_B7866_ = new_B7828_ & new_B7865_;
  assign new_B7865_ = new_B7884_ | new_B7883_;
  assign new_B7864_ = ~new_B7828_ & new_B7863_;
  assign new_B7863_ = new_B7886_ | new_B7885_;
  assign new_B7862_ = new_B7828_ | new_B7861_;
  assign new_B7861_ = new_B7882_ | new_B7881_;
  assign new_B7860_ = ~new_B7840_ & ~new_B7850_;
  assign new_B7859_ = new_B7840_ & new_B7850_;
  assign new_B7858_ = ~new_B7840_ | new_B7850_;
  assign new_B7857_ = new_B7824_ & ~new_B7825_;
  assign new_B7856_ = ~new_B7824_ & new_B7825_;
  assign new_B7855_ = new_B7877_ & ~new_B7878_;
  assign new_B7854_ = ~new_B7877_ & new_B7878_;
  assign new_B7853_ = ~new_B7876_ | ~new_B7875_;
  assign new_B7852_ = new_B7868_ | new_B7867_;
  assign new_B7851_ = new_B7874_ | new_B7873_;
  assign new_B7850_ = new_B7864_ | new_B7866_;
  assign new_B7849_ = ~new_B7871_ | ~new_B7872_;
  assign new_B7848_ = new_B7824_ & ~new_B7825_;
  assign new_B7847_ = new_B7838_ & ~new_B7850_;
  assign new_B7846_ = ~new_B7838_ & new_B7850_;
  assign new_B7845_ = ~new_B7836_ & new_B7862_;
  assign new_B7844_ = new_B7860_ | new_B7859_;
  assign new_B7843_ = new_B7857_ | new_B7856_;
  assign new_B7842_ = new_B7825_ | new_B7858_;
  assign new_B7841_ = new_B7850_ & new_B7853_;
  assign new_B7840_ = new_B7855_ | new_B7854_;
  assign new_B7839_ = new_B7850_ & new_B7849_;
  assign new_B7838_ = new_B7852_ & new_B7851_;
  assign new_B7837_ = new_B7847_ | new_B7846_;
  assign new_B7836_ = new_B7825_ | new_B7848_;
  assign B7835 = new_B7836_ | new_B7845_;
  assign B7834 = new_B7843_ & new_B7844_;
  assign B7833 = new_B7843_ & new_B7842_;
  assign B7832 = new_B7841_ | new_B7840_;
  assign B7831 = new_B7839_ | new_B7838_;
  assign B7830 = new_B7837_ & new_B7836_;
  assign new_B7829_ = new_C3664_;
  assign new_B7828_ = new_C3597_;
  assign new_B7827_ = new_C3530_;
  assign new_B7826_ = new_C3463_;
  assign new_B7825_ = new_C3396_;
  assign new_B7824_ = new_C3329_;
  assign new_B7823_ = ~new_B7762_ & new_B7776_;
  assign new_B7822_ = new_B7762_ & ~new_B7776_;
  assign new_B7821_ = new_B7762_ & ~new_B7776_;
  assign new_B7820_ = ~new_B7762_ & ~new_B7776_;
  assign new_B7819_ = new_B7762_ & new_B7776_;
  assign new_B7818_ = new_B7822_ | new_B7823_;
  assign new_B7817_ = ~new_B7762_ & new_B7776_;
  assign new_B7816_ = new_B7820_ | new_B7821_;
  assign new_B7815_ = ~new_B7791_ & ~new_B7811_;
  assign new_B7814_ = new_B7791_ & new_B7811_;
  assign new_B7813_ = ~new_B7758_ | ~new_B7783_;
  assign new_B7812_ = new_B7776_ & new_B7813_;
  assign new_B7811_ = new_B7759_ | new_B7760_;
  assign new_B7810_ = new_B7759_ | new_B7776_;
  assign new_B7809_ = ~new_B7776_ & ~new_B7812_;
  assign new_B7808_ = new_B7776_ | new_B7813_;
  assign new_B7807_ = new_B7759_ & ~new_B7760_;
  assign new_B7806_ = ~new_B7759_ & new_B7760_;
  assign new_B7805_ = new_B7769_ | new_B7802_;
  assign new_B7804_ = ~new_B7769_ & ~new_B7803_;
  assign new_B7803_ = new_B7769_ & new_B7802_;
  assign new_B7802_ = ~new_B7758_ | ~new_B7783_;
  assign new_B7801_ = ~new_B7759_ & new_B7769_;
  assign new_B7800_ = new_B7759_ & ~new_B7769_;
  assign new_B7799_ = new_B7761_ & new_B7798_;
  assign new_B7798_ = new_B7817_ | new_B7816_;
  assign new_B7797_ = ~new_B7761_ & new_B7796_;
  assign new_B7796_ = new_B7819_ | new_B7818_;
  assign new_B7795_ = new_B7761_ | new_B7794_;
  assign new_B7794_ = new_B7815_ | new_B7814_;
  assign new_B7793_ = ~new_B7773_ & ~new_B7783_;
  assign new_B7792_ = new_B7773_ & new_B7783_;
  assign new_B7791_ = ~new_B7773_ | new_B7783_;
  assign new_B7790_ = new_B7757_ & ~new_B7758_;
  assign new_B7789_ = ~new_B7757_ & new_B7758_;
  assign new_B7788_ = new_B7810_ & ~new_B7811_;
  assign new_B7787_ = ~new_B7810_ & new_B7811_;
  assign new_B7786_ = ~new_B7809_ | ~new_B7808_;
  assign new_B7785_ = new_B7801_ | new_B7800_;
  assign new_B7784_ = new_B7807_ | new_B7806_;
  assign new_B7783_ = new_B7797_ | new_B7799_;
  assign new_B7782_ = ~new_B7804_ | ~new_B7805_;
  assign new_B7781_ = new_B7757_ & ~new_B7758_;
  assign new_B7780_ = new_B7771_ & ~new_B7783_;
  assign new_B7779_ = ~new_B7771_ & new_B7783_;
  assign new_B7778_ = ~new_B7769_ & new_B7795_;
  assign new_B7777_ = new_B7793_ | new_B7792_;
  assign new_B7776_ = new_B7790_ | new_B7789_;
  assign new_B7775_ = new_B7758_ | new_B7791_;
  assign new_B7774_ = new_B7783_ & new_B7786_;
  assign new_B7773_ = new_B7788_ | new_B7787_;
  assign new_B7772_ = new_B7783_ & new_B7782_;
  assign new_B7771_ = new_B7785_ & new_B7784_;
  assign new_B7770_ = new_B7780_ | new_B7779_;
  assign new_B7769_ = new_B7758_ | new_B7781_;
  assign B7768 = new_B7769_ | new_B7778_;
  assign B7767 = new_B7776_ & new_B7777_;
  assign B7766 = new_B7776_ & new_B7775_;
  assign B7765 = new_B7774_ | new_B7773_;
  assign B7764 = new_B7772_ | new_B7771_;
  assign B7763 = new_B7770_ & new_B7769_;
  assign new_B7762_ = new_C3262_;
  assign new_B7761_ = new_C3195_;
  assign new_B7760_ = new_C3128_;
  assign new_B7759_ = new_C3061_;
  assign new_B7758_ = new_C2994_;
  assign new_B7757_ = new_C2927_;
  assign new_B7756_ = ~new_B7695_ & new_B7709_;
  assign new_B7755_ = new_B7695_ & ~new_B7709_;
  assign new_B7754_ = new_B7695_ & ~new_B7709_;
  assign new_B7753_ = ~new_B7695_ & ~new_B7709_;
  assign new_B7752_ = new_B7695_ & new_B7709_;
  assign new_B7751_ = new_B7755_ | new_B7756_;
  assign new_B7750_ = ~new_B7695_ & new_B7709_;
  assign new_B7749_ = new_B7753_ | new_B7754_;
  assign new_B7748_ = ~new_B7724_ & ~new_B7744_;
  assign new_B7747_ = new_B7724_ & new_B7744_;
  assign new_B7746_ = ~new_B7691_ | ~new_B7716_;
  assign new_B7745_ = new_B7709_ & new_B7746_;
  assign new_B7744_ = new_B7692_ | new_B7693_;
  assign new_B7743_ = new_B7692_ | new_B7709_;
  assign new_B7742_ = ~new_B7709_ & ~new_B7745_;
  assign new_B7741_ = new_B7709_ | new_B7746_;
  assign new_B7740_ = new_B7692_ & ~new_B7693_;
  assign new_B7739_ = ~new_B7692_ & new_B7693_;
  assign new_B7738_ = new_B7702_ | new_B7735_;
  assign new_B7737_ = ~new_B7702_ & ~new_B7736_;
  assign new_B7736_ = new_B7702_ & new_B7735_;
  assign new_B7735_ = ~new_B7691_ | ~new_B7716_;
  assign new_B7734_ = ~new_B7692_ & new_B7702_;
  assign new_B7733_ = new_B7692_ & ~new_B7702_;
  assign new_B7732_ = new_B7694_ & new_B7731_;
  assign new_B7731_ = new_B7750_ | new_B7749_;
  assign new_B7730_ = ~new_B7694_ & new_B7729_;
  assign new_B7729_ = new_B7752_ | new_B7751_;
  assign new_B7728_ = new_B7694_ | new_B7727_;
  assign new_B7727_ = new_B7748_ | new_B7747_;
  assign new_B7726_ = ~new_B7706_ & ~new_B7716_;
  assign new_B7725_ = new_B7706_ & new_B7716_;
  assign new_B7724_ = ~new_B7706_ | new_B7716_;
  assign new_B7723_ = new_B7690_ & ~new_B7691_;
  assign new_B7722_ = ~new_B7690_ & new_B7691_;
  assign new_B7721_ = new_B7743_ & ~new_B7744_;
  assign new_B7720_ = ~new_B7743_ & new_B7744_;
  assign new_B7719_ = ~new_B7742_ | ~new_B7741_;
  assign new_B7718_ = new_B7734_ | new_B7733_;
  assign new_B7717_ = new_B7740_ | new_B7739_;
  assign new_B7716_ = new_B7730_ | new_B7732_;
  assign new_B7715_ = ~new_B7737_ | ~new_B7738_;
  assign new_B7714_ = new_B7690_ & ~new_B7691_;
  assign new_B7713_ = new_B7704_ & ~new_B7716_;
  assign new_B7712_ = ~new_B7704_ & new_B7716_;
  assign new_B7711_ = ~new_B7702_ & new_B7728_;
  assign new_B7710_ = new_B7726_ | new_B7725_;
  assign new_B7709_ = new_B7723_ | new_B7722_;
  assign new_B7708_ = new_B7691_ | new_B7724_;
  assign new_B7707_ = new_B7716_ & new_B7719_;
  assign new_B7706_ = new_B7721_ | new_B7720_;
  assign new_B7705_ = new_B7716_ & new_B7715_;
  assign new_B7704_ = new_B7718_ & new_B7717_;
  assign new_B7703_ = new_B7713_ | new_B7712_;
  assign new_B7702_ = new_B7691_ | new_B7714_;
  assign B7701 = new_B7702_ | new_B7711_;
  assign B7700 = new_B7709_ & new_B7710_;
  assign B7699 = new_B7709_ & new_B7708_;
  assign B7698 = new_B7707_ | new_B7706_;
  assign B7697 = new_B7705_ | new_B7704_;
  assign B7696 = new_B7703_ & new_B7702_;
  assign new_B7695_ = new_C2860_;
  assign new_B7694_ = new_C2793_;
  assign new_B7693_ = new_C2726_;
  assign new_B7692_ = new_C2659_;
  assign new_B7691_ = new_C2592_;
  assign new_B7690_ = new_C2522_;
  assign new_B7689_ = ~new_B7628_ & new_B7642_;
  assign new_B7688_ = new_B7628_ & ~new_B7642_;
  assign new_B7687_ = new_B7628_ & ~new_B7642_;
  assign new_B7686_ = ~new_B7628_ & ~new_B7642_;
  assign new_B7685_ = new_B7628_ & new_B7642_;
  assign new_B7684_ = new_B7688_ | new_B7689_;
  assign new_B7683_ = ~new_B7628_ & new_B7642_;
  assign new_B7682_ = new_B7686_ | new_B7687_;
  assign new_B7681_ = ~new_B7657_ & ~new_B7677_;
  assign new_B7680_ = new_B7657_ & new_B7677_;
  assign new_B7679_ = ~new_B7624_ | ~new_B7649_;
  assign new_B7678_ = new_B7642_ & new_B7679_;
  assign new_B7677_ = new_B7625_ | new_B7626_;
  assign new_B7676_ = new_B7625_ | new_B7642_;
  assign new_B7675_ = ~new_B7642_ & ~new_B7678_;
  assign new_B7674_ = new_B7642_ | new_B7679_;
  assign new_B7673_ = new_B7625_ & ~new_B7626_;
  assign new_B7672_ = ~new_B7625_ & new_B7626_;
  assign new_B7671_ = new_B7635_ | new_B7668_;
  assign new_B7670_ = ~new_B7635_ & ~new_B7669_;
  assign new_B7669_ = new_B7635_ & new_B7668_;
  assign new_B7668_ = ~new_B7624_ | ~new_B7649_;
  assign new_B7667_ = ~new_B7625_ & new_B7635_;
  assign new_B7666_ = new_B7625_ & ~new_B7635_;
  assign new_B7665_ = new_B7627_ & new_B7664_;
  assign new_B7664_ = new_B7683_ | new_B7682_;
  assign new_B7663_ = ~new_B7627_ & new_B7662_;
  assign new_B7662_ = new_B7685_ | new_B7684_;
  assign new_B7661_ = new_B7627_ | new_B7660_;
  assign new_B7660_ = new_B7681_ | new_B7680_;
  assign new_B7659_ = ~new_B7639_ & ~new_B7649_;
  assign new_B7658_ = new_B7639_ & new_B7649_;
  assign new_B7657_ = ~new_B7639_ | new_B7649_;
  assign new_B7656_ = new_B7623_ & ~new_B7624_;
  assign new_B7655_ = ~new_B7623_ & new_B7624_;
  assign new_B7654_ = new_B7676_ & ~new_B7677_;
  assign new_B7653_ = ~new_B7676_ & new_B7677_;
  assign new_B7652_ = ~new_B7675_ | ~new_B7674_;
  assign new_B7651_ = new_B7667_ | new_B7666_;
  assign new_B7650_ = new_B7673_ | new_B7672_;
  assign new_B7649_ = new_B7663_ | new_B7665_;
  assign new_B7648_ = ~new_B7670_ | ~new_B7671_;
  assign new_B7647_ = new_B7623_ & ~new_B7624_;
  assign new_B7646_ = new_B7637_ & ~new_B7649_;
  assign new_B7645_ = ~new_B7637_ & new_B7649_;
  assign new_B7644_ = ~new_B7635_ & new_B7661_;
  assign new_B7643_ = new_B7659_ | new_B7658_;
  assign new_B7642_ = new_B7656_ | new_B7655_;
  assign new_B7641_ = new_B7624_ | new_B7657_;
  assign new_B7640_ = new_B7649_ & new_B7652_;
  assign new_B7639_ = new_B7654_ | new_B7653_;
  assign new_B7638_ = new_B7649_ & new_B7648_;
  assign new_B7637_ = new_B7651_ & new_B7650_;
  assign new_B7636_ = new_B7646_ | new_B7645_;
  assign new_B7635_ = new_B7624_ | new_B7647_;
  assign B7634 = new_B7635_ | new_B7644_;
  assign B7633 = new_B7642_ & new_B7643_;
  assign B7632 = new_B7642_ & new_B7641_;
  assign B7631 = new_B7640_ | new_B7639_;
  assign B7630 = new_B7638_ | new_B7637_;
  assign B7629 = new_B7636_ & new_B7635_;
  assign new_B7628_ = new_D6930_;
  assign new_B7627_ = new_D6863_;
  assign new_B7626_ = new_D6796_;
  assign new_B7625_ = new_D6729_;
  assign new_B7624_ = new_D6662_;
  assign new_B7623_ = new_D6595_;
  assign new_B7622_ = ~new_B7561_ & new_B7575_;
  assign new_B7621_ = new_B7561_ & ~new_B7575_;
  assign new_B7620_ = new_B7561_ & ~new_B7575_;
  assign new_B7619_ = ~new_B7561_ & ~new_B7575_;
  assign new_B7618_ = new_B7561_ & new_B7575_;
  assign new_B7617_ = new_B7621_ | new_B7622_;
  assign new_B7616_ = ~new_B7561_ & new_B7575_;
  assign new_B7615_ = new_B7619_ | new_B7620_;
  assign new_B7614_ = ~new_B7590_ & ~new_B7610_;
  assign new_B7613_ = new_B7590_ & new_B7610_;
  assign new_B7612_ = ~new_B7557_ | ~new_B7582_;
  assign new_B7611_ = new_B7575_ & new_B7612_;
  assign new_B7610_ = new_B7558_ | new_B7559_;
  assign new_B7609_ = new_B7558_ | new_B7575_;
  assign new_B7608_ = ~new_B7575_ & ~new_B7611_;
  assign new_B7607_ = new_B7575_ | new_B7612_;
  assign new_B7606_ = new_B7558_ & ~new_B7559_;
  assign new_B7605_ = ~new_B7558_ & new_B7559_;
  assign new_B7604_ = new_B7568_ | new_B7601_;
  assign new_B7603_ = ~new_B7568_ & ~new_B7602_;
  assign new_B7602_ = new_B7568_ & new_B7601_;
  assign new_B7601_ = ~new_B7557_ | ~new_B7582_;
  assign new_B7600_ = ~new_B7558_ & new_B7568_;
  assign new_B7599_ = new_B7558_ & ~new_B7568_;
  assign new_B7598_ = new_B7560_ & new_B7597_;
  assign new_B7597_ = new_B7616_ | new_B7615_;
  assign new_B7596_ = ~new_B7560_ & new_B7595_;
  assign new_B7595_ = new_B7618_ | new_B7617_;
  assign new_B7594_ = new_B7560_ | new_B7593_;
  assign new_B7593_ = new_B7614_ | new_B7613_;
  assign new_B7592_ = ~new_B7572_ & ~new_B7582_;
  assign new_B7591_ = new_B7572_ & new_B7582_;
  assign new_B7590_ = ~new_B7572_ | new_B7582_;
  assign new_B7589_ = new_B7556_ & ~new_B7557_;
  assign new_B7588_ = ~new_B7556_ & new_B7557_;
  assign new_B7587_ = new_B7609_ & ~new_B7610_;
  assign new_B7586_ = ~new_B7609_ & new_B7610_;
  assign new_B7585_ = ~new_B7608_ | ~new_B7607_;
  assign new_B7584_ = new_B7600_ | new_B7599_;
  assign new_B7583_ = new_B7606_ | new_B7605_;
  assign new_B7582_ = new_B7596_ | new_B7598_;
  assign new_B7581_ = ~new_B7603_ | ~new_B7604_;
  assign new_B7580_ = new_B7556_ & ~new_B7557_;
  assign new_B7579_ = new_B7570_ & ~new_B7582_;
  assign new_B7578_ = ~new_B7570_ & new_B7582_;
  assign new_B7577_ = ~new_B7568_ & new_B7594_;
  assign new_B7576_ = new_B7592_ | new_B7591_;
  assign new_B7575_ = new_B7589_ | new_B7588_;
  assign new_B7574_ = new_B7557_ | new_B7590_;
  assign new_B7573_ = new_B7582_ & new_B7585_;
  assign new_B7572_ = new_B7587_ | new_B7586_;
  assign new_B7571_ = new_B7582_ & new_B7581_;
  assign new_B7570_ = new_B7584_ & new_B7583_;
  assign new_B7569_ = new_B7579_ | new_B7578_;
  assign new_B7568_ = new_B7557_ | new_B7580_;
  assign B7567 = new_B7568_ | new_B7577_;
  assign B7566 = new_B7575_ & new_B7576_;
  assign B7565 = new_B7575_ & new_B7574_;
  assign B7564 = new_B7573_ | new_B7572_;
  assign B7563 = new_B7571_ | new_B7570_;
  assign B7562 = new_B7569_ & new_B7568_;
  assign new_B7561_ = new_D6528_;
  assign new_B7560_ = new_D6461_;
  assign new_B7559_ = new_D6394_;
  assign new_B7558_ = new_D6327_;
  assign new_B7557_ = new_D6260_;
  assign new_B7556_ = new_D6193_;
  assign new_B7555_ = ~new_B7494_ & new_B7508_;
  assign new_B7554_ = new_B7494_ & ~new_B7508_;
  assign new_B7553_ = new_B7494_ & ~new_B7508_;
  assign new_B7552_ = ~new_B7494_ & ~new_B7508_;
  assign new_B7551_ = new_B7494_ & new_B7508_;
  assign new_B7550_ = new_B7554_ | new_B7555_;
  assign new_B7549_ = ~new_B7494_ & new_B7508_;
  assign new_B7548_ = new_B7552_ | new_B7553_;
  assign new_B7547_ = ~new_B7523_ & ~new_B7543_;
  assign new_B7546_ = new_B7523_ & new_B7543_;
  assign new_B7545_ = ~new_B7490_ | ~new_B7515_;
  assign new_B7544_ = new_B7508_ & new_B7545_;
  assign new_B7543_ = new_B7491_ | new_B7492_;
  assign new_B7542_ = new_B7491_ | new_B7508_;
  assign new_B7541_ = ~new_B7508_ & ~new_B7544_;
  assign new_B7540_ = new_B7508_ | new_B7545_;
  assign new_B7539_ = new_B7491_ & ~new_B7492_;
  assign new_B7538_ = ~new_B7491_ & new_B7492_;
  assign new_B7537_ = new_B7501_ | new_B7534_;
  assign new_B7536_ = ~new_B7501_ & ~new_B7535_;
  assign new_B7535_ = new_B7501_ & new_B7534_;
  assign new_B7534_ = ~new_B7490_ | ~new_B7515_;
  assign new_B7533_ = ~new_B7491_ & new_B7501_;
  assign new_B7532_ = new_B7491_ & ~new_B7501_;
  assign new_B7531_ = new_B7493_ & new_B7530_;
  assign new_B7530_ = new_B7549_ | new_B7548_;
  assign new_B7529_ = ~new_B7493_ & new_B7528_;
  assign new_B7528_ = new_B7551_ | new_B7550_;
  assign new_B7527_ = new_B7493_ | new_B7526_;
  assign new_B7526_ = new_B7547_ | new_B7546_;
  assign new_B7525_ = ~new_B7505_ & ~new_B7515_;
  assign new_B7524_ = new_B7505_ & new_B7515_;
  assign new_B7523_ = ~new_B7505_ | new_B7515_;
  assign new_B7522_ = new_B7489_ & ~new_B7490_;
  assign new_B7521_ = ~new_B7489_ & new_B7490_;
  assign new_B7520_ = new_B7542_ & ~new_B7543_;
  assign new_B7519_ = ~new_B7542_ & new_B7543_;
  assign new_B7518_ = ~new_B7541_ | ~new_B7540_;
  assign new_B7517_ = new_B7533_ | new_B7532_;
  assign new_B7516_ = new_B7539_ | new_B7538_;
  assign new_B7515_ = new_B7529_ | new_B7531_;
  assign new_B7514_ = ~new_B7536_ | ~new_B7537_;
  assign new_B7513_ = new_B7489_ & ~new_B7490_;
  assign new_B7512_ = new_B7503_ & ~new_B7515_;
  assign new_B7511_ = ~new_B7503_ & new_B7515_;
  assign new_B7510_ = ~new_B7501_ & new_B7527_;
  assign new_B7509_ = new_B7525_ | new_B7524_;
  assign new_B7508_ = new_B7522_ | new_B7521_;
  assign new_B7507_ = new_B7490_ | new_B7523_;
  assign new_B7506_ = new_B7515_ & new_B7518_;
  assign new_B7505_ = new_B7520_ | new_B7519_;
  assign new_B7504_ = new_B7515_ & new_B7514_;
  assign new_B7503_ = new_B7517_ & new_B7516_;
  assign new_B7502_ = new_B7512_ | new_B7511_;
  assign new_B7501_ = new_B7490_ | new_B7513_;
  assign B7500 = new_B7501_ | new_B7510_;
  assign B7499 = new_B7508_ & new_B7509_;
  assign B7498 = new_B7508_ & new_B7507_;
  assign B7497 = new_B7506_ | new_B7505_;
  assign B7496 = new_B7504_ | new_B7503_;
  assign B7495 = new_B7502_ & new_B7501_;
  assign new_B7494_ = new_D6126_;
  assign new_B7493_ = new_D6059_;
  assign new_B7492_ = new_D5992_;
  assign new_B7491_ = new_D5925_;
  assign new_B7490_ = new_D5858_;
  assign new_B7489_ = new_D5791_;
  assign new_B7488_ = ~new_B7427_ & new_B7441_;
  assign new_B7487_ = new_B7427_ & ~new_B7441_;
  assign new_B7486_ = new_B7427_ & ~new_B7441_;
  assign new_B7485_ = ~new_B7427_ & ~new_B7441_;
  assign new_B7484_ = new_B7427_ & new_B7441_;
  assign new_B7483_ = new_B7487_ | new_B7488_;
  assign new_B7482_ = ~new_B7427_ & new_B7441_;
  assign new_B7481_ = new_B7485_ | new_B7486_;
  assign new_B7480_ = ~new_B7456_ & ~new_B7476_;
  assign new_B7479_ = new_B7456_ & new_B7476_;
  assign new_B7478_ = ~new_B7423_ | ~new_B7448_;
  assign new_B7477_ = new_B7441_ & new_B7478_;
  assign new_B7476_ = new_B7424_ | new_B7425_;
  assign new_B7475_ = new_B7424_ | new_B7441_;
  assign new_B7474_ = ~new_B7441_ & ~new_B7477_;
  assign new_B7473_ = new_B7441_ | new_B7478_;
  assign new_B7472_ = new_B7424_ & ~new_B7425_;
  assign new_B7471_ = ~new_B7424_ & new_B7425_;
  assign new_B7470_ = new_B7434_ | new_B7467_;
  assign new_B7469_ = ~new_B7434_ & ~new_B7468_;
  assign new_B7468_ = new_B7434_ & new_B7467_;
  assign new_B7467_ = ~new_B7423_ | ~new_B7448_;
  assign new_B7466_ = ~new_B7424_ & new_B7434_;
  assign new_B7465_ = new_B7424_ & ~new_B7434_;
  assign new_B7464_ = new_B7426_ & new_B7463_;
  assign new_B7463_ = new_B7482_ | new_B7481_;
  assign new_B7462_ = ~new_B7426_ & new_B7461_;
  assign new_B7461_ = new_B7484_ | new_B7483_;
  assign new_B7460_ = new_B7426_ | new_B7459_;
  assign new_B7459_ = new_B7480_ | new_B7479_;
  assign new_B7458_ = ~new_B7438_ & ~new_B7448_;
  assign new_B7457_ = new_B7438_ & new_B7448_;
  assign new_B7456_ = ~new_B7438_ | new_B7448_;
  assign new_B7455_ = new_B7422_ & ~new_B7423_;
  assign new_B7454_ = ~new_B7422_ & new_B7423_;
  assign new_B7453_ = new_B7475_ & ~new_B7476_;
  assign new_B7452_ = ~new_B7475_ & new_B7476_;
  assign new_B7451_ = ~new_B7474_ | ~new_B7473_;
  assign new_B7450_ = new_B7466_ | new_B7465_;
  assign new_B7449_ = new_B7472_ | new_B7471_;
  assign new_B7448_ = new_B7462_ | new_B7464_;
  assign new_B7447_ = ~new_B7469_ | ~new_B7470_;
  assign new_B7446_ = new_B7422_ & ~new_B7423_;
  assign new_B7445_ = new_B7436_ & ~new_B7448_;
  assign new_B7444_ = ~new_B7436_ & new_B7448_;
  assign new_B7443_ = ~new_B7434_ & new_B7460_;
  assign new_B7442_ = new_B7458_ | new_B7457_;
  assign new_B7441_ = new_B7455_ | new_B7454_;
  assign new_B7440_ = new_B7423_ | new_B7456_;
  assign new_B7439_ = new_B7448_ & new_B7451_;
  assign new_B7438_ = new_B7453_ | new_B7452_;
  assign new_B7437_ = new_B7448_ & new_B7447_;
  assign new_B7436_ = new_B7450_ & new_B7449_;
  assign new_B7435_ = new_B7445_ | new_B7444_;
  assign new_B7434_ = new_B7423_ | new_B7446_;
  assign B7433 = new_B7434_ | new_B7443_;
  assign B7432 = new_B7441_ & new_B7442_;
  assign B7431 = new_B7441_ & new_B7440_;
  assign B7430 = new_B7439_ | new_B7438_;
  assign B7429 = new_B7437_ | new_B7436_;
  assign B7428 = new_B7435_ & new_B7434_;
  assign new_B7427_ = new_D5724_;
  assign new_B7426_ = new_D5657_;
  assign new_B7425_ = new_D5590_;
  assign new_B7424_ = new_D5523_;
  assign new_B7423_ = new_D5456_;
  assign new_B7422_ = new_D5389_;
  assign new_B7421_ = ~new_B7360_ & new_B7374_;
  assign new_B7420_ = new_B7360_ & ~new_B7374_;
  assign new_B7419_ = new_B7360_ & ~new_B7374_;
  assign new_B7418_ = ~new_B7360_ & ~new_B7374_;
  assign new_B7417_ = new_B7360_ & new_B7374_;
  assign new_B7416_ = new_B7420_ | new_B7421_;
  assign new_B7415_ = ~new_B7360_ & new_B7374_;
  assign new_B7414_ = new_B7418_ | new_B7419_;
  assign new_B7413_ = ~new_B7389_ & ~new_B7409_;
  assign new_B7412_ = new_B7389_ & new_B7409_;
  assign new_B7411_ = ~new_B7356_ | ~new_B7381_;
  assign new_B7410_ = new_B7374_ & new_B7411_;
  assign new_B7409_ = new_B7357_ | new_B7358_;
  assign new_B7408_ = new_B7357_ | new_B7374_;
  assign new_B7407_ = ~new_B7374_ & ~new_B7410_;
  assign new_B7406_ = new_B7374_ | new_B7411_;
  assign new_B7405_ = new_B7357_ & ~new_B7358_;
  assign new_B7404_ = ~new_B7357_ & new_B7358_;
  assign new_B7403_ = new_B7367_ | new_B7400_;
  assign new_B7402_ = ~new_B7367_ & ~new_B7401_;
  assign new_B7401_ = new_B7367_ & new_B7400_;
  assign new_B7400_ = ~new_B7356_ | ~new_B7381_;
  assign new_B7399_ = ~new_B7357_ & new_B7367_;
  assign new_B7398_ = new_B7357_ & ~new_B7367_;
  assign new_B7397_ = new_B7359_ & new_B7396_;
  assign new_B7396_ = new_B7415_ | new_B7414_;
  assign new_B7395_ = ~new_B7359_ & new_B7394_;
  assign new_B7394_ = new_B7417_ | new_B7416_;
  assign new_B7393_ = new_B7359_ | new_B7392_;
  assign new_B7392_ = new_B7413_ | new_B7412_;
  assign new_B7391_ = ~new_B7371_ & ~new_B7381_;
  assign new_B7390_ = new_B7371_ & new_B7381_;
  assign new_B7389_ = ~new_B7371_ | new_B7381_;
  assign new_B7388_ = new_B7355_ & ~new_B7356_;
  assign new_B7387_ = ~new_B7355_ & new_B7356_;
  assign new_B7386_ = new_B7408_ & ~new_B7409_;
  assign new_B7385_ = ~new_B7408_ & new_B7409_;
  assign new_B7384_ = ~new_B7407_ | ~new_B7406_;
  assign new_B7383_ = new_B7399_ | new_B7398_;
  assign new_B7382_ = new_B7405_ | new_B7404_;
  assign new_B7381_ = new_B7395_ | new_B7397_;
  assign new_B7380_ = ~new_B7402_ | ~new_B7403_;
  assign new_B7379_ = new_B7355_ & ~new_B7356_;
  assign new_B7378_ = new_B7369_ & ~new_B7381_;
  assign new_B7377_ = ~new_B7369_ & new_B7381_;
  assign new_B7376_ = ~new_B7367_ & new_B7393_;
  assign new_B7375_ = new_B7391_ | new_B7390_;
  assign new_B7374_ = new_B7388_ | new_B7387_;
  assign new_B7373_ = new_B7356_ | new_B7389_;
  assign new_B7372_ = new_B7381_ & new_B7384_;
  assign new_B7371_ = new_B7386_ | new_B7385_;
  assign new_B7370_ = new_B7381_ & new_B7380_;
  assign new_B7369_ = new_B7383_ & new_B7382_;
  assign new_B7368_ = new_B7378_ | new_B7377_;
  assign new_B7367_ = new_B7356_ | new_B7379_;
  assign B7366 = new_B7367_ | new_B7376_;
  assign B7365 = new_B7374_ & new_B7375_;
  assign B7364 = new_B7374_ & new_B7373_;
  assign B7363 = new_B7372_ | new_B7371_;
  assign B7362 = new_B7370_ | new_B7369_;
  assign B7361 = new_B7368_ & new_B7367_;
  assign new_B7360_ = new_D5322_;
  assign new_B7359_ = new_D5255_;
  assign new_B7358_ = new_D5188_;
  assign new_B7357_ = new_D5121_;
  assign new_B7356_ = new_D5054_;
  assign new_B7355_ = new_D4987_;
  assign new_B7354_ = ~new_B7293_ & new_B7307_;
  assign new_B7353_ = new_B7293_ & ~new_B7307_;
  assign new_B7352_ = new_B7293_ & ~new_B7307_;
  assign new_B7351_ = ~new_B7293_ & ~new_B7307_;
  assign new_B7350_ = new_B7293_ & new_B7307_;
  assign new_B7349_ = new_B7353_ | new_B7354_;
  assign new_B7348_ = ~new_B7293_ & new_B7307_;
  assign new_B7347_ = new_B7351_ | new_B7352_;
  assign new_B7346_ = ~new_B7322_ & ~new_B7342_;
  assign new_B7345_ = new_B7322_ & new_B7342_;
  assign new_B7344_ = ~new_B7289_ | ~new_B7314_;
  assign new_B7343_ = new_B7307_ & new_B7344_;
  assign new_B7342_ = new_B7290_ | new_B7291_;
  assign new_B7341_ = new_B7290_ | new_B7307_;
  assign new_B7340_ = ~new_B7307_ & ~new_B7343_;
  assign new_B7339_ = new_B7307_ | new_B7344_;
  assign new_B7338_ = new_B7290_ & ~new_B7291_;
  assign new_B7337_ = ~new_B7290_ & new_B7291_;
  assign new_B7336_ = new_B7300_ | new_B7333_;
  assign new_B7335_ = ~new_B7300_ & ~new_B7334_;
  assign new_B7334_ = new_B7300_ & new_B7333_;
  assign new_B7333_ = ~new_B7289_ | ~new_B7314_;
  assign new_B7332_ = ~new_B7290_ & new_B7300_;
  assign new_B7331_ = new_B7290_ & ~new_B7300_;
  assign new_B7330_ = new_B7292_ & new_B7329_;
  assign new_B7329_ = new_B7348_ | new_B7347_;
  assign new_B7328_ = ~new_B7292_ & new_B7327_;
  assign new_B7327_ = new_B7350_ | new_B7349_;
  assign new_B7326_ = new_B7292_ | new_B7325_;
  assign new_B7325_ = new_B7346_ | new_B7345_;
  assign new_B7324_ = ~new_B7304_ & ~new_B7314_;
  assign new_B7323_ = new_B7304_ & new_B7314_;
  assign new_B7322_ = ~new_B7304_ | new_B7314_;
  assign new_B7321_ = new_B7288_ & ~new_B7289_;
  assign new_B7320_ = ~new_B7288_ & new_B7289_;
  assign new_B7319_ = new_B7341_ & ~new_B7342_;
  assign new_B7318_ = ~new_B7341_ & new_B7342_;
  assign new_B7317_ = ~new_B7340_ | ~new_B7339_;
  assign new_B7316_ = new_B7332_ | new_B7331_;
  assign new_B7315_ = new_B7338_ | new_B7337_;
  assign new_B7314_ = new_B7328_ | new_B7330_;
  assign new_B7313_ = ~new_B7335_ | ~new_B7336_;
  assign new_B7312_ = new_B7288_ & ~new_B7289_;
  assign new_B7311_ = new_B7302_ & ~new_B7314_;
  assign new_B7310_ = ~new_B7302_ & new_B7314_;
  assign new_B7309_ = ~new_B7300_ & new_B7326_;
  assign new_B7308_ = new_B7324_ | new_B7323_;
  assign new_B7307_ = new_B7321_ | new_B7320_;
  assign new_B7306_ = new_B7289_ | new_B7322_;
  assign new_B7305_ = new_B7314_ & new_B7317_;
  assign new_B7304_ = new_B7319_ | new_B7318_;
  assign new_B7303_ = new_B7314_ & new_B7313_;
  assign new_B7302_ = new_B7316_ & new_B7315_;
  assign new_B7301_ = new_B7311_ | new_B7310_;
  assign new_B7300_ = new_B7289_ | new_B7312_;
  assign B7299 = new_B7300_ | new_B7309_;
  assign B7298 = new_B7307_ & new_B7308_;
  assign B7297 = new_B7307_ & new_B7306_;
  assign B7296 = new_B7305_ | new_B7304_;
  assign B7295 = new_B7303_ | new_B7302_;
  assign B7294 = new_B7301_ & new_B7300_;
  assign new_B7293_ = new_D4920_;
  assign new_B7292_ = new_D4853_;
  assign new_B7291_ = new_D4786_;
  assign new_B7290_ = new_D4719_;
  assign new_B7289_ = new_D4652_;
  assign new_B7288_ = new_D4585_;
  assign new_B7287_ = ~new_B7226_ & new_B7240_;
  assign new_B7286_ = new_B7226_ & ~new_B7240_;
  assign new_B7285_ = new_B7226_ & ~new_B7240_;
  assign new_B7284_ = ~new_B7226_ & ~new_B7240_;
  assign new_B7283_ = new_B7226_ & new_B7240_;
  assign new_B7282_ = new_B7286_ | new_B7287_;
  assign new_B7281_ = ~new_B7226_ & new_B7240_;
  assign new_B7280_ = new_B7284_ | new_B7285_;
  assign new_B7279_ = ~new_B7255_ & ~new_B7275_;
  assign new_B7278_ = new_B7255_ & new_B7275_;
  assign new_B7277_ = ~new_B7222_ | ~new_B7247_;
  assign new_B7276_ = new_B7240_ & new_B7277_;
  assign new_B7275_ = new_B7223_ | new_B7224_;
  assign new_B7274_ = new_B7223_ | new_B7240_;
  assign new_B7273_ = ~new_B7240_ & ~new_B7276_;
  assign new_B7272_ = new_B7240_ | new_B7277_;
  assign new_B7271_ = new_B7223_ & ~new_B7224_;
  assign new_B7270_ = ~new_B7223_ & new_B7224_;
  assign new_B7269_ = new_B7233_ | new_B7266_;
  assign new_B7268_ = ~new_B7233_ & ~new_B7267_;
  assign new_B7267_ = new_B7233_ & new_B7266_;
  assign new_B7266_ = ~new_B7222_ | ~new_B7247_;
  assign new_B7265_ = ~new_B7223_ & new_B7233_;
  assign new_B7264_ = new_B7223_ & ~new_B7233_;
  assign new_B7263_ = new_B7225_ & new_B7262_;
  assign new_B7262_ = new_B7281_ | new_B7280_;
  assign new_B7261_ = ~new_B7225_ & new_B7260_;
  assign new_B7260_ = new_B7283_ | new_B7282_;
  assign new_B7259_ = new_B7225_ | new_B7258_;
  assign new_B7258_ = new_B7279_ | new_B7278_;
  assign new_B7257_ = ~new_B7237_ & ~new_B7247_;
  assign new_B7256_ = new_B7237_ & new_B7247_;
  assign new_B7255_ = ~new_B7237_ | new_B7247_;
  assign new_B7254_ = new_B7221_ & ~new_B7222_;
  assign new_B7253_ = ~new_B7221_ & new_B7222_;
  assign new_B7252_ = new_B7274_ & ~new_B7275_;
  assign new_B7251_ = ~new_B7274_ & new_B7275_;
  assign new_B7250_ = ~new_B7273_ | ~new_B7272_;
  assign new_B7249_ = new_B7265_ | new_B7264_;
  assign new_B7248_ = new_B7271_ | new_B7270_;
  assign new_B7247_ = new_B7261_ | new_B7263_;
  assign new_B7246_ = ~new_B7268_ | ~new_B7269_;
  assign new_B7245_ = new_B7221_ & ~new_B7222_;
  assign new_B7244_ = new_B7235_ & ~new_B7247_;
  assign new_B7243_ = ~new_B7235_ & new_B7247_;
  assign new_B7242_ = ~new_B7233_ & new_B7259_;
  assign new_B7241_ = new_B7257_ | new_B7256_;
  assign new_B7240_ = new_B7254_ | new_B7253_;
  assign new_B7239_ = new_B7222_ | new_B7255_;
  assign new_B7238_ = new_B7247_ & new_B7250_;
  assign new_B7237_ = new_B7252_ | new_B7251_;
  assign new_B7236_ = new_B7247_ & new_B7246_;
  assign new_B7235_ = new_B7249_ & new_B7248_;
  assign new_B7234_ = new_B7244_ | new_B7243_;
  assign new_B7233_ = new_B7222_ | new_B7245_;
  assign B7232 = new_B7233_ | new_B7242_;
  assign B7231 = new_B7240_ & new_B7241_;
  assign B7230 = new_B7240_ & new_B7239_;
  assign B7229 = new_B7238_ | new_B7237_;
  assign B7228 = new_B7236_ | new_B7235_;
  assign B7227 = new_B7234_ & new_B7233_;
  assign new_B7226_ = new_D4518_;
  assign new_B7225_ = new_D4451_;
  assign new_B7224_ = new_D4384_;
  assign new_B7223_ = new_D4317_;
  assign new_B7222_ = new_D4250_;
  assign new_B7221_ = new_D4183_;
  assign new_B7220_ = ~new_B7159_ & new_B7173_;
  assign new_B7219_ = new_B7159_ & ~new_B7173_;
  assign new_B7218_ = new_B7159_ & ~new_B7173_;
  assign new_B7217_ = ~new_B7159_ & ~new_B7173_;
  assign new_B7216_ = new_B7159_ & new_B7173_;
  assign new_B7215_ = new_B7219_ | new_B7220_;
  assign new_B7214_ = ~new_B7159_ & new_B7173_;
  assign new_B7213_ = new_B7217_ | new_B7218_;
  assign new_B7212_ = ~new_B7188_ & ~new_B7208_;
  assign new_B7211_ = new_B7188_ & new_B7208_;
  assign new_B7210_ = ~new_B7155_ | ~new_B7180_;
  assign new_B7209_ = new_B7173_ & new_B7210_;
  assign new_B7208_ = new_B7156_ | new_B7157_;
  assign new_B7207_ = new_B7156_ | new_B7173_;
  assign new_B7206_ = ~new_B7173_ & ~new_B7209_;
  assign new_B7205_ = new_B7173_ | new_B7210_;
  assign new_B7204_ = new_B7156_ & ~new_B7157_;
  assign new_B7203_ = ~new_B7156_ & new_B7157_;
  assign new_B7202_ = new_B7166_ | new_B7199_;
  assign new_B7201_ = ~new_B7166_ & ~new_B7200_;
  assign new_B7200_ = new_B7166_ & new_B7199_;
  assign new_B7199_ = ~new_B7155_ | ~new_B7180_;
  assign new_B7198_ = ~new_B7156_ & new_B7166_;
  assign new_B7197_ = new_B7156_ & ~new_B7166_;
  assign new_B7196_ = new_B7158_ & new_B7195_;
  assign new_B7195_ = new_B7214_ | new_B7213_;
  assign new_B7194_ = ~new_B7158_ & new_B7193_;
  assign new_B7193_ = new_B7216_ | new_B7215_;
  assign new_B7192_ = new_B7158_ | new_B7191_;
  assign new_B7191_ = new_B7212_ | new_B7211_;
  assign new_B7190_ = ~new_B7170_ & ~new_B7180_;
  assign new_B7189_ = new_B7170_ & new_B7180_;
  assign new_B7188_ = ~new_B7170_ | new_B7180_;
  assign new_B7187_ = new_B7154_ & ~new_B7155_;
  assign new_B7186_ = ~new_B7154_ & new_B7155_;
  assign new_B7185_ = new_B7207_ & ~new_B7208_;
  assign new_B7184_ = ~new_B7207_ & new_B7208_;
  assign new_B7183_ = ~new_B7206_ | ~new_B7205_;
  assign new_B7182_ = new_B7198_ | new_B7197_;
  assign new_B7181_ = new_B7204_ | new_B7203_;
  assign new_B7180_ = new_B7194_ | new_B7196_;
  assign new_B7179_ = ~new_B7201_ | ~new_B7202_;
  assign new_B7178_ = new_B7154_ & ~new_B7155_;
  assign new_B7177_ = new_B7168_ & ~new_B7180_;
  assign new_B7176_ = ~new_B7168_ & new_B7180_;
  assign new_B7175_ = ~new_B7166_ & new_B7192_;
  assign new_B7174_ = new_B7190_ | new_B7189_;
  assign new_B7173_ = new_B7187_ | new_B7186_;
  assign new_B7172_ = new_B7155_ | new_B7188_;
  assign new_B7171_ = new_B7180_ & new_B7183_;
  assign new_B7170_ = new_B7185_ | new_B7184_;
  assign new_B7169_ = new_B7180_ & new_B7179_;
  assign new_B7168_ = new_B7182_ & new_B7181_;
  assign new_B7167_ = new_B7177_ | new_B7176_;
  assign new_B7166_ = new_B7155_ | new_B7178_;
  assign B7165 = new_B7166_ | new_B7175_;
  assign B7164 = new_B7173_ & new_B7174_;
  assign B7163 = new_B7173_ & new_B7172_;
  assign B7162 = new_B7171_ | new_B7170_;
  assign B7161 = new_B7169_ | new_B7168_;
  assign B7160 = new_B7167_ & new_B7166_;
  assign new_B7159_ = new_D4116_;
  assign new_B7158_ = new_D4049_;
  assign new_B7157_ = new_D3982_;
  assign new_B7156_ = new_D3915_;
  assign new_B7155_ = new_D3848_;
  assign new_B7154_ = new_D3781_;
  assign new_B7153_ = ~new_B7092_ & new_B7106_;
  assign new_B7152_ = new_B7092_ & ~new_B7106_;
  assign new_B7151_ = new_B7092_ & ~new_B7106_;
  assign new_B7150_ = ~new_B7092_ & ~new_B7106_;
  assign new_B7149_ = new_B7092_ & new_B7106_;
  assign new_B7148_ = new_B7152_ | new_B7153_;
  assign new_B7147_ = ~new_B7092_ & new_B7106_;
  assign new_B7146_ = new_B7150_ | new_B7151_;
  assign new_B7145_ = ~new_B7121_ & ~new_B7141_;
  assign new_B7144_ = new_B7121_ & new_B7141_;
  assign new_B7143_ = ~new_B7088_ | ~new_B7113_;
  assign new_B7142_ = new_B7106_ & new_B7143_;
  assign new_B7141_ = new_B7089_ | new_B7090_;
  assign new_B7140_ = new_B7089_ | new_B7106_;
  assign new_B7139_ = ~new_B7106_ & ~new_B7142_;
  assign new_B7138_ = new_B7106_ | new_B7143_;
  assign new_B7137_ = new_B7089_ & ~new_B7090_;
  assign new_B7136_ = ~new_B7089_ & new_B7090_;
  assign new_B7135_ = new_B7099_ | new_B7132_;
  assign new_B7134_ = ~new_B7099_ & ~new_B7133_;
  assign new_B7133_ = new_B7099_ & new_B7132_;
  assign new_B7132_ = ~new_B7088_ | ~new_B7113_;
  assign new_B7131_ = ~new_B7089_ & new_B7099_;
  assign new_B7130_ = new_B7089_ & ~new_B7099_;
  assign new_B7129_ = new_B7091_ & new_B7128_;
  assign new_B7128_ = new_B7147_ | new_B7146_;
  assign new_B7127_ = ~new_B7091_ & new_B7126_;
  assign new_B7126_ = new_B7149_ | new_B7148_;
  assign new_B7125_ = new_B7091_ | new_B7124_;
  assign new_B7124_ = new_B7145_ | new_B7144_;
  assign new_B7123_ = ~new_B7103_ & ~new_B7113_;
  assign new_B7122_ = new_B7103_ & new_B7113_;
  assign new_B7121_ = ~new_B7103_ | new_B7113_;
  assign new_B7120_ = new_B7087_ & ~new_B7088_;
  assign new_B7119_ = ~new_B7087_ & new_B7088_;
  assign new_B7118_ = new_B7140_ & ~new_B7141_;
  assign new_B7117_ = ~new_B7140_ & new_B7141_;
  assign new_B7116_ = ~new_B7139_ | ~new_B7138_;
  assign new_B7115_ = new_B7131_ | new_B7130_;
  assign new_B7114_ = new_B7137_ | new_B7136_;
  assign new_B7113_ = new_B7127_ | new_B7129_;
  assign new_B7112_ = ~new_B7134_ | ~new_B7135_;
  assign new_B7111_ = new_B7087_ & ~new_B7088_;
  assign new_B7110_ = new_B7101_ & ~new_B7113_;
  assign new_B7109_ = ~new_B7101_ & new_B7113_;
  assign new_B7108_ = ~new_B7099_ & new_B7125_;
  assign new_B7107_ = new_B7123_ | new_B7122_;
  assign new_B7106_ = new_B7120_ | new_B7119_;
  assign new_B7105_ = new_B7088_ | new_B7121_;
  assign new_B7104_ = new_B7113_ & new_B7116_;
  assign new_B7103_ = new_B7118_ | new_B7117_;
  assign new_B7102_ = new_B7113_ & new_B7112_;
  assign new_B7101_ = new_B7115_ & new_B7114_;
  assign new_B7100_ = new_B7110_ | new_B7109_;
  assign new_B7099_ = new_B7088_ | new_B7111_;
  assign B7098 = new_B7099_ | new_B7108_;
  assign B7097 = new_B7106_ & new_B7107_;
  assign B7096 = new_B7106_ & new_B7105_;
  assign B7095 = new_B7104_ | new_B7103_;
  assign B7094 = new_B7102_ | new_B7101_;
  assign B7093 = new_B7100_ & new_B7099_;
  assign new_B7092_ = new_D3714_;
  assign new_B7091_ = new_D3647_;
  assign new_B7090_ = new_D3580_;
  assign new_B7089_ = new_D3513_;
  assign new_B7088_ = new_D3446_;
  assign new_B7087_ = new_D3379_;
  assign new_B7086_ = ~new_B7025_ & new_B7039_;
  assign new_B7085_ = new_B7025_ & ~new_B7039_;
  assign new_B7084_ = new_B7025_ & ~new_B7039_;
  assign new_B7083_ = ~new_B7025_ & ~new_B7039_;
  assign new_B7082_ = new_B7025_ & new_B7039_;
  assign new_B7081_ = new_B7085_ | new_B7086_;
  assign new_B7080_ = ~new_B7025_ & new_B7039_;
  assign new_B7079_ = new_B7083_ | new_B7084_;
  assign new_B7078_ = ~new_B7054_ & ~new_B7074_;
  assign new_B7077_ = new_B7054_ & new_B7074_;
  assign new_B7076_ = ~new_B7021_ | ~new_B7046_;
  assign new_B7075_ = new_B7039_ & new_B7076_;
  assign new_B7074_ = new_B7022_ | new_B7023_;
  assign new_B7073_ = new_B7022_ | new_B7039_;
  assign new_B7072_ = ~new_B7039_ & ~new_B7075_;
  assign new_B7071_ = new_B7039_ | new_B7076_;
  assign new_B7070_ = new_B7022_ & ~new_B7023_;
  assign new_B7069_ = ~new_B7022_ & new_B7023_;
  assign new_B7068_ = new_B7032_ | new_B7065_;
  assign new_B7067_ = ~new_B7032_ & ~new_B7066_;
  assign new_B7066_ = new_B7032_ & new_B7065_;
  assign new_B7065_ = ~new_B7021_ | ~new_B7046_;
  assign new_B7064_ = ~new_B7022_ & new_B7032_;
  assign new_B7063_ = new_B7022_ & ~new_B7032_;
  assign new_B7062_ = new_B7024_ & new_B7061_;
  assign new_B7061_ = new_B7080_ | new_B7079_;
  assign new_B7060_ = ~new_B7024_ & new_B7059_;
  assign new_B7059_ = new_B7082_ | new_B7081_;
  assign new_B7058_ = new_B7024_ | new_B7057_;
  assign new_B7057_ = new_B7078_ | new_B7077_;
  assign new_B7056_ = ~new_B7036_ & ~new_B7046_;
  assign new_B7055_ = new_B7036_ & new_B7046_;
  assign new_B7054_ = ~new_B7036_ | new_B7046_;
  assign new_B7053_ = new_B7020_ & ~new_B7021_;
  assign new_B7052_ = ~new_B7020_ & new_B7021_;
  assign new_B7051_ = new_B7073_ & ~new_B7074_;
  assign new_B7050_ = ~new_B7073_ & new_B7074_;
  assign new_B7049_ = ~new_B7072_ | ~new_B7071_;
  assign new_B7048_ = new_B7064_ | new_B7063_;
  assign new_B7047_ = new_B7070_ | new_B7069_;
  assign new_B7046_ = new_B7060_ | new_B7062_;
  assign new_B7045_ = ~new_B7067_ | ~new_B7068_;
  assign new_B7044_ = new_B7020_ & ~new_B7021_;
  assign new_B7043_ = new_B7034_ & ~new_B7046_;
  assign new_B7042_ = ~new_B7034_ & new_B7046_;
  assign new_B7041_ = ~new_B7032_ & new_B7058_;
  assign new_B7040_ = new_B7056_ | new_B7055_;
  assign new_B7039_ = new_B7053_ | new_B7052_;
  assign new_B7038_ = new_B7021_ | new_B7054_;
  assign new_B7037_ = new_B7046_ & new_B7049_;
  assign new_B7036_ = new_B7051_ | new_B7050_;
  assign new_B7035_ = new_B7046_ & new_B7045_;
  assign new_B7034_ = new_B7048_ & new_B7047_;
  assign new_B7033_ = new_B7043_ | new_B7042_;
  assign new_B7032_ = new_B7021_ | new_B7044_;
  assign B7031 = new_B7032_ | new_B7041_;
  assign B7030 = new_B7039_ & new_B7040_;
  assign B7029 = new_B7039_ & new_B7038_;
  assign B7028 = new_B7037_ | new_B7036_;
  assign B7027 = new_B7035_ | new_B7034_;
  assign B7026 = new_B7033_ & new_B7032_;
  assign new_B7025_ = new_D3312_;
  assign new_B7024_ = new_D3245_;
  assign new_B7023_ = new_D3178_;
  assign new_B7022_ = new_D3111_;
  assign new_B7021_ = new_D3044_;
  assign new_B7020_ = new_D2977_;
  assign new_B7019_ = ~new_B6958_ & new_B6972_;
  assign new_B7018_ = new_B6958_ & ~new_B6972_;
  assign new_B7017_ = new_B6958_ & ~new_B6972_;
  assign new_B7016_ = ~new_B6958_ & ~new_B6972_;
  assign new_B7015_ = new_B6958_ & new_B6972_;
  assign new_B7014_ = new_B7018_ | new_B7019_;
  assign new_B7013_ = ~new_B6958_ & new_B6972_;
  assign new_B7012_ = new_B7016_ | new_B7017_;
  assign new_B7011_ = ~new_B6987_ & ~new_B7007_;
  assign new_B7010_ = new_B6987_ & new_B7007_;
  assign new_B7009_ = ~new_B6954_ | ~new_B6979_;
  assign new_B7008_ = new_B6972_ & new_B7009_;
  assign new_B7007_ = new_B6955_ | new_B6956_;
  assign new_B7006_ = new_B6955_ | new_B6972_;
  assign new_B7005_ = ~new_B6972_ & ~new_B7008_;
  assign new_B7004_ = new_B6972_ | new_B7009_;
  assign new_B7003_ = new_B6955_ & ~new_B6956_;
  assign new_B7002_ = ~new_B6955_ & new_B6956_;
  assign new_B7001_ = new_B6965_ | new_B6998_;
  assign new_B7000_ = ~new_B6965_ & ~new_B6999_;
  assign new_B6999_ = new_B6965_ & new_B6998_;
  assign new_B6998_ = ~new_B6954_ | ~new_B6979_;
  assign new_B6997_ = ~new_B6955_ & new_B6965_;
  assign new_B6996_ = new_B6955_ & ~new_B6965_;
  assign new_B6995_ = new_B6957_ & new_B6994_;
  assign new_B6994_ = new_B7013_ | new_B7012_;
  assign new_B6993_ = ~new_B6957_ & new_B6992_;
  assign new_B6992_ = new_B7015_ | new_B7014_;
  assign new_B6991_ = new_B6957_ | new_B6990_;
  assign new_B6990_ = new_B7011_ | new_B7010_;
  assign new_B6989_ = ~new_B6969_ & ~new_B6979_;
  assign new_B6988_ = new_B6969_ & new_B6979_;
  assign new_B6987_ = ~new_B6969_ | new_B6979_;
  assign new_B6986_ = new_B6953_ & ~new_B6954_;
  assign new_B6985_ = ~new_B6953_ & new_B6954_;
  assign new_B6984_ = new_B7006_ & ~new_B7007_;
  assign new_B6983_ = ~new_B7006_ & new_B7007_;
  assign new_B6982_ = ~new_B7005_ | ~new_B7004_;
  assign new_B6981_ = new_B6997_ | new_B6996_;
  assign new_B6980_ = new_B7003_ | new_B7002_;
  assign new_B6979_ = new_B6993_ | new_B6995_;
  assign new_B6978_ = ~new_B7000_ | ~new_B7001_;
  assign new_B6977_ = new_B6953_ & ~new_B6954_;
  assign new_B6976_ = new_B6967_ & ~new_B6979_;
  assign new_B6975_ = ~new_B6967_ & new_B6979_;
  assign new_B6974_ = ~new_B6965_ & new_B6991_;
  assign new_B6973_ = new_B6989_ | new_B6988_;
  assign new_B6972_ = new_B6986_ | new_B6985_;
  assign new_B6971_ = new_B6954_ | new_B6987_;
  assign new_B6970_ = new_B6979_ & new_B6982_;
  assign new_B6969_ = new_B6984_ | new_B6983_;
  assign new_B6968_ = new_B6979_ & new_B6978_;
  assign new_B6967_ = new_B6981_ & new_B6980_;
  assign new_B6966_ = new_B6976_ | new_B6975_;
  assign new_B6965_ = new_B6954_ | new_B6977_;
  assign B6964 = new_B6965_ | new_B6974_;
  assign B6963 = new_B6972_ & new_B6973_;
  assign B6962 = new_B6972_ & new_B6971_;
  assign B6961 = new_B6970_ | new_B6969_;
  assign B6960 = new_B6968_ | new_B6967_;
  assign B6959 = new_B6966_ & new_B6965_;
  assign new_B6958_ = new_D2910_;
  assign new_B6957_ = new_D2843_;
  assign new_B6956_ = new_D2776_;
  assign new_B6955_ = new_D2709_;
  assign new_B6954_ = new_D2642_;
  assign new_B6953_ = new_D2575_;
  assign new_B6952_ = ~new_B6891_ & new_B6905_;
  assign new_B6951_ = new_B6891_ & ~new_B6905_;
  assign new_B6950_ = new_B6891_ & ~new_B6905_;
  assign new_B6949_ = ~new_B6891_ & ~new_B6905_;
  assign new_B6948_ = new_B6891_ & new_B6905_;
  assign new_B6947_ = new_B6951_ | new_B6952_;
  assign new_B6946_ = ~new_B6891_ & new_B6905_;
  assign new_B6945_ = new_B6949_ | new_B6950_;
  assign new_B6944_ = ~new_B6920_ & ~new_B6940_;
  assign new_B6943_ = new_B6920_ & new_B6940_;
  assign new_B6942_ = ~new_B6887_ | ~new_B6912_;
  assign new_B6941_ = new_B6905_ & new_B6942_;
  assign new_B6940_ = new_B6888_ | new_B6889_;
  assign new_B6939_ = new_B6888_ | new_B6905_;
  assign new_B6938_ = ~new_B6905_ & ~new_B6941_;
  assign new_B6937_ = new_B6905_ | new_B6942_;
  assign new_B6936_ = new_B6888_ & ~new_B6889_;
  assign new_B6935_ = ~new_B6888_ & new_B6889_;
  assign new_B6934_ = new_B6898_ | new_B6931_;
  assign new_B6933_ = ~new_B6898_ & ~new_B6932_;
  assign new_B6932_ = new_B6898_ & new_B6931_;
  assign new_B6931_ = ~new_B6887_ | ~new_B6912_;
  assign new_B6930_ = ~new_B6888_ & new_B6898_;
  assign new_B6929_ = new_B6888_ & ~new_B6898_;
  assign new_B6928_ = new_B6890_ & new_B6927_;
  assign new_B6927_ = new_B6946_ | new_B6945_;
  assign new_B6926_ = ~new_B6890_ & new_B6925_;
  assign new_B6925_ = new_B6948_ | new_B6947_;
  assign new_B6924_ = new_B6890_ | new_B6923_;
  assign new_B6923_ = new_B6944_ | new_B6943_;
  assign new_B6922_ = ~new_B6902_ & ~new_B6912_;
  assign new_B6921_ = new_B6902_ & new_B6912_;
  assign new_B6920_ = ~new_B6902_ | new_B6912_;
  assign new_B6919_ = new_B6886_ & ~new_B6887_;
  assign new_B6918_ = ~new_B6886_ & new_B6887_;
  assign new_B6917_ = new_B6939_ & ~new_B6940_;
  assign new_B6916_ = ~new_B6939_ & new_B6940_;
  assign new_B6915_ = ~new_B6938_ | ~new_B6937_;
  assign new_B6914_ = new_B6930_ | new_B6929_;
  assign new_B6913_ = new_B6936_ | new_B6935_;
  assign new_B6912_ = new_B6926_ | new_B6928_;
  assign new_B6911_ = ~new_B6933_ | ~new_B6934_;
  assign new_B6910_ = new_B6886_ & ~new_B6887_;
  assign new_B6909_ = new_B6900_ & ~new_B6912_;
  assign new_B6908_ = ~new_B6900_ & new_B6912_;
  assign new_B6907_ = ~new_B6898_ & new_B6924_;
  assign new_B6906_ = new_B6922_ | new_B6921_;
  assign new_B6905_ = new_B6919_ | new_B6918_;
  assign new_B6904_ = new_B6887_ | new_B6920_;
  assign new_B6903_ = new_B6912_ & new_B6915_;
  assign new_B6902_ = new_B6917_ | new_B6916_;
  assign new_B6901_ = new_B6912_ & new_B6911_;
  assign new_B6900_ = new_B6914_ & new_B6913_;
  assign new_B6899_ = new_B6909_ | new_B6908_;
  assign new_B6898_ = new_B6887_ | new_B6910_;
  assign B6897 = new_B6898_ | new_B6907_;
  assign B6896 = new_B6905_ & new_B6906_;
  assign B6895 = new_B6905_ & new_B6904_;
  assign B6894 = new_B6903_ | new_B6902_;
  assign B6893 = new_B6901_ | new_B6900_;
  assign B6892 = new_B6899_ & new_B6898_;
  assign new_B6891_ = new_D2508_;
  assign new_B6890_ = new_D2441_;
  assign new_B6889_ = new_D2374_;
  assign new_B6888_ = new_D2307_;
  assign new_B6887_ = new_D2240_;
  assign new_B6886_ = new_D2173_;
  assign new_B6885_ = ~new_B6824_ & new_B6838_;
  assign new_B6884_ = new_B6824_ & ~new_B6838_;
  assign new_B6883_ = new_B6824_ & ~new_B6838_;
  assign new_B6882_ = ~new_B6824_ & ~new_B6838_;
  assign new_B6881_ = new_B6824_ & new_B6838_;
  assign new_B6880_ = new_B6884_ | new_B6885_;
  assign new_B6879_ = ~new_B6824_ & new_B6838_;
  assign new_B6878_ = new_B6882_ | new_B6883_;
  assign new_B6877_ = ~new_B6853_ & ~new_B6873_;
  assign new_B6876_ = new_B6853_ & new_B6873_;
  assign new_B6875_ = ~new_B6820_ | ~new_B6845_;
  assign new_B6874_ = new_B6838_ & new_B6875_;
  assign new_B6873_ = new_B6821_ | new_B6822_;
  assign new_B6872_ = new_B6821_ | new_B6838_;
  assign new_B6871_ = ~new_B6838_ & ~new_B6874_;
  assign new_B6870_ = new_B6838_ | new_B6875_;
  assign new_B6869_ = new_B6821_ & ~new_B6822_;
  assign new_B6868_ = ~new_B6821_ & new_B6822_;
  assign new_B6867_ = new_B6831_ | new_B6864_;
  assign new_B6866_ = ~new_B6831_ & ~new_B6865_;
  assign new_B6865_ = new_B6831_ & new_B6864_;
  assign new_B6864_ = ~new_B6820_ | ~new_B6845_;
  assign new_B6863_ = ~new_B6821_ & new_B6831_;
  assign new_B6862_ = new_B6821_ & ~new_B6831_;
  assign new_B6861_ = new_B6823_ & new_B6860_;
  assign new_B6860_ = new_B6879_ | new_B6878_;
  assign new_B6859_ = ~new_B6823_ & new_B6858_;
  assign new_B6858_ = new_B6881_ | new_B6880_;
  assign new_B6857_ = new_B6823_ | new_B6856_;
  assign new_B6856_ = new_B6877_ | new_B6876_;
  assign new_B6855_ = ~new_B6835_ & ~new_B6845_;
  assign new_B6854_ = new_B6835_ & new_B6845_;
  assign new_B6853_ = ~new_B6835_ | new_B6845_;
  assign new_B6852_ = new_B6819_ & ~new_B6820_;
  assign new_B6851_ = ~new_B6819_ & new_B6820_;
  assign new_B6850_ = new_B6872_ & ~new_B6873_;
  assign new_B6849_ = ~new_B6872_ & new_B6873_;
  assign new_B6848_ = ~new_B6871_ | ~new_B6870_;
  assign new_B6847_ = new_B6863_ | new_B6862_;
  assign new_B6846_ = new_B6869_ | new_B6868_;
  assign new_B6845_ = new_B6859_ | new_B6861_;
  assign new_B6844_ = ~new_B6866_ | ~new_B6867_;
  assign new_B6843_ = new_B6819_ & ~new_B6820_;
  assign new_B6842_ = new_B6833_ & ~new_B6845_;
  assign new_B6841_ = ~new_B6833_ & new_B6845_;
  assign new_B6840_ = ~new_B6831_ & new_B6857_;
  assign new_B6839_ = new_B6855_ | new_B6854_;
  assign new_B6838_ = new_B6852_ | new_B6851_;
  assign new_B6837_ = new_B6820_ | new_B6853_;
  assign new_B6836_ = new_B6845_ & new_B6848_;
  assign new_B6835_ = new_B6850_ | new_B6849_;
  assign new_B6834_ = new_B6845_ & new_B6844_;
  assign new_B6833_ = new_B6847_ & new_B6846_;
  assign new_B6832_ = new_B6842_ | new_B6841_;
  assign new_B6831_ = new_B6820_ | new_B6843_;
  assign B6830 = new_B6831_ | new_B6840_;
  assign B6829 = new_B6838_ & new_B6839_;
  assign B6828 = new_B6838_ & new_B6837_;
  assign B6827 = new_B6836_ | new_B6835_;
  assign B6826 = new_B6834_ | new_B6833_;
  assign B6825 = new_B6832_ & new_B6831_;
  assign new_B6824_ = new_D2106_;
  assign new_B6823_ = new_D2039_;
  assign new_B6822_ = new_D1972_;
  assign new_B6821_ = new_D1905_;
  assign new_B6820_ = new_D1838_;
  assign new_B6819_ = new_D1771_;
  assign new_B6818_ = ~new_B6757_ & new_B6771_;
  assign new_B6817_ = new_B6757_ & ~new_B6771_;
  assign new_B6816_ = new_B6757_ & ~new_B6771_;
  assign new_B6815_ = ~new_B6757_ & ~new_B6771_;
  assign new_B6814_ = new_B6757_ & new_B6771_;
  assign new_B6813_ = new_B6817_ | new_B6818_;
  assign new_B6812_ = ~new_B6757_ & new_B6771_;
  assign new_B6811_ = new_B6815_ | new_B6816_;
  assign new_B6810_ = ~new_B6786_ & ~new_B6806_;
  assign new_B6809_ = new_B6786_ & new_B6806_;
  assign new_B6808_ = ~new_B6753_ | ~new_B6778_;
  assign new_B6807_ = new_B6771_ & new_B6808_;
  assign new_B6806_ = new_B6754_ | new_B6755_;
  assign new_B6805_ = new_B6754_ | new_B6771_;
  assign new_B6804_ = ~new_B6771_ & ~new_B6807_;
  assign new_B6803_ = new_B6771_ | new_B6808_;
  assign new_B6802_ = new_B6754_ & ~new_B6755_;
  assign new_B6801_ = ~new_B6754_ & new_B6755_;
  assign new_B6800_ = new_B6764_ | new_B6797_;
  assign new_B6799_ = ~new_B6764_ & ~new_B6798_;
  assign new_B6798_ = new_B6764_ & new_B6797_;
  assign new_B6797_ = ~new_B6753_ | ~new_B6778_;
  assign new_B6796_ = ~new_B6754_ & new_B6764_;
  assign new_B6795_ = new_B6754_ & ~new_B6764_;
  assign new_B6794_ = new_B6756_ & new_B6793_;
  assign new_B6793_ = new_B6812_ | new_B6811_;
  assign new_B6792_ = ~new_B6756_ & new_B6791_;
  assign new_B6791_ = new_B6814_ | new_B6813_;
  assign new_B6790_ = new_B6756_ | new_B6789_;
  assign new_B6789_ = new_B6810_ | new_B6809_;
  assign new_B6788_ = ~new_B6768_ & ~new_B6778_;
  assign new_B6787_ = new_B6768_ & new_B6778_;
  assign new_B6786_ = ~new_B6768_ | new_B6778_;
  assign new_B6785_ = new_B6752_ & ~new_B6753_;
  assign new_B6784_ = ~new_B6752_ & new_B6753_;
  assign new_B6783_ = new_B6805_ & ~new_B6806_;
  assign new_B6782_ = ~new_B6805_ & new_B6806_;
  assign new_B6781_ = ~new_B6804_ | ~new_B6803_;
  assign new_B6780_ = new_B6796_ | new_B6795_;
  assign new_B6779_ = new_B6802_ | new_B6801_;
  assign new_B6778_ = new_B6792_ | new_B6794_;
  assign new_B6777_ = ~new_B6799_ | ~new_B6800_;
  assign new_B6776_ = new_B6752_ & ~new_B6753_;
  assign new_B6775_ = new_B6766_ & ~new_B6778_;
  assign new_B6774_ = ~new_B6766_ & new_B6778_;
  assign new_B6773_ = ~new_B6764_ & new_B6790_;
  assign new_B6772_ = new_B6788_ | new_B6787_;
  assign new_B6771_ = new_B6785_ | new_B6784_;
  assign new_B6770_ = new_B6753_ | new_B6786_;
  assign new_B6769_ = new_B6778_ & new_B6781_;
  assign new_B6768_ = new_B6783_ | new_B6782_;
  assign new_B6767_ = new_B6778_ & new_B6777_;
  assign new_B6766_ = new_B6780_ & new_B6779_;
  assign new_B6765_ = new_B6775_ | new_B6774_;
  assign new_B6764_ = new_B6753_ | new_B6776_;
  assign B6763 = new_B6764_ | new_B6773_;
  assign B6762 = new_B6771_ & new_B6772_;
  assign B6761 = new_B6771_ & new_B6770_;
  assign B6760 = new_B6769_ | new_B6768_;
  assign B6759 = new_B6767_ | new_B6766_;
  assign B6758 = new_B6765_ & new_B6764_;
  assign new_B6757_ = new_D1704_;
  assign new_B6756_ = new_D1637_;
  assign new_B6755_ = new_D1570_;
  assign new_B6754_ = new_D1503_;
  assign new_B6753_ = new_D1436_;
  assign new_B6752_ = new_D1369_;
  assign new_B6751_ = ~new_B6690_ & new_B6704_;
  assign new_B6750_ = new_B6690_ & ~new_B6704_;
  assign new_B6749_ = new_B6690_ & ~new_B6704_;
  assign new_B6748_ = ~new_B6690_ & ~new_B6704_;
  assign new_B6747_ = new_B6690_ & new_B6704_;
  assign new_B6746_ = new_B6750_ | new_B6751_;
  assign new_B6745_ = ~new_B6690_ & new_B6704_;
  assign new_B6744_ = new_B6748_ | new_B6749_;
  assign new_B6743_ = ~new_B6719_ & ~new_B6739_;
  assign new_B6742_ = new_B6719_ & new_B6739_;
  assign new_B6741_ = ~new_B6686_ | ~new_B6711_;
  assign new_B6740_ = new_B6704_ & new_B6741_;
  assign new_B6739_ = new_B6687_ | new_B6688_;
  assign new_B6738_ = new_B6687_ | new_B6704_;
  assign new_B6737_ = ~new_B6704_ & ~new_B6740_;
  assign new_B6736_ = new_B6704_ | new_B6741_;
  assign new_B6735_ = new_B6687_ & ~new_B6688_;
  assign new_B6734_ = ~new_B6687_ & new_B6688_;
  assign new_B6733_ = new_B6697_ | new_B6730_;
  assign new_B6732_ = ~new_B6697_ & ~new_B6731_;
  assign new_B6731_ = new_B6697_ & new_B6730_;
  assign new_B6730_ = ~new_B6686_ | ~new_B6711_;
  assign new_B6729_ = ~new_B6687_ & new_B6697_;
  assign new_B6728_ = new_B6687_ & ~new_B6697_;
  assign new_B6727_ = new_B6689_ & new_B6726_;
  assign new_B6726_ = new_B6745_ | new_B6744_;
  assign new_B6725_ = ~new_B6689_ & new_B6724_;
  assign new_B6724_ = new_B6747_ | new_B6746_;
  assign new_B6723_ = new_B6689_ | new_B6722_;
  assign new_B6722_ = new_B6743_ | new_B6742_;
  assign new_B6721_ = ~new_B6701_ & ~new_B6711_;
  assign new_B6720_ = new_B6701_ & new_B6711_;
  assign new_B6719_ = ~new_B6701_ | new_B6711_;
  assign new_B6718_ = new_B6685_ & ~new_B6686_;
  assign new_B6717_ = ~new_B6685_ & new_B6686_;
  assign new_B6716_ = new_B6738_ & ~new_B6739_;
  assign new_B6715_ = ~new_B6738_ & new_B6739_;
  assign new_B6714_ = ~new_B6737_ | ~new_B6736_;
  assign new_B6713_ = new_B6729_ | new_B6728_;
  assign new_B6712_ = new_B6735_ | new_B6734_;
  assign new_B6711_ = new_B6725_ | new_B6727_;
  assign new_B6710_ = ~new_B6732_ | ~new_B6733_;
  assign new_B6709_ = new_B6685_ & ~new_B6686_;
  assign new_B6708_ = new_B6699_ & ~new_B6711_;
  assign new_B6707_ = ~new_B6699_ & new_B6711_;
  assign new_B6706_ = ~new_B6697_ & new_B6723_;
  assign new_B6705_ = new_B6721_ | new_B6720_;
  assign new_B6704_ = new_B6718_ | new_B6717_;
  assign new_B6703_ = new_B6686_ | new_B6719_;
  assign new_B6702_ = new_B6711_ & new_B6714_;
  assign new_B6701_ = new_B6716_ | new_B6715_;
  assign new_B6700_ = new_B6711_ & new_B6710_;
  assign new_B6699_ = new_B6713_ & new_B6712_;
  assign new_B6698_ = new_B6708_ | new_B6707_;
  assign new_B6697_ = new_B6686_ | new_B6709_;
  assign B6696 = new_B6697_ | new_B6706_;
  assign B6695 = new_B6704_ & new_B6705_;
  assign B6694 = new_B6704_ & new_B6703_;
  assign B6693 = new_B6702_ | new_B6701_;
  assign B6692 = new_B6700_ | new_B6699_;
  assign B6691 = new_B6698_ & new_B6697_;
  assign new_B6690_ = new_D1302_;
  assign new_B6689_ = new_D1235_;
  assign new_B6688_ = new_D1168_;
  assign new_B6687_ = new_D1101_;
  assign new_B6686_ = new_D1034_;
  assign new_B6685_ = new_D967_;
  assign new_B6684_ = ~new_B6623_ & new_B6637_;
  assign new_B6683_ = new_B6623_ & ~new_B6637_;
  assign new_B6682_ = new_B6623_ & ~new_B6637_;
  assign new_B6681_ = ~new_B6623_ & ~new_B6637_;
  assign new_B6680_ = new_B6623_ & new_B6637_;
  assign new_B6679_ = new_B6683_ | new_B6684_;
  assign new_B6678_ = ~new_B6623_ & new_B6637_;
  assign new_B6677_ = new_B6681_ | new_B6682_;
  assign new_B6676_ = ~new_B6652_ & ~new_B6672_;
  assign new_B6675_ = new_B6652_ & new_B6672_;
  assign new_B6674_ = ~new_B6619_ | ~new_B6644_;
  assign new_B6673_ = new_B6637_ & new_B6674_;
  assign new_B6672_ = new_B6620_ | new_B6621_;
  assign new_B6671_ = new_B6620_ | new_B6637_;
  assign new_B6670_ = ~new_B6637_ & ~new_B6673_;
  assign new_B6669_ = new_B6637_ | new_B6674_;
  assign new_B6668_ = new_B6620_ & ~new_B6621_;
  assign new_B6667_ = ~new_B6620_ & new_B6621_;
  assign new_B6666_ = new_B6630_ | new_B6663_;
  assign new_B6665_ = ~new_B6630_ & ~new_B6664_;
  assign new_B6664_ = new_B6630_ & new_B6663_;
  assign new_B6663_ = ~new_B6619_ | ~new_B6644_;
  assign new_B6662_ = ~new_B6620_ & new_B6630_;
  assign new_B6661_ = new_B6620_ & ~new_B6630_;
  assign new_B6660_ = new_B6622_ & new_B6659_;
  assign new_B6659_ = new_B6678_ | new_B6677_;
  assign new_B6658_ = ~new_B6622_ & new_B6657_;
  assign new_B6657_ = new_B6680_ | new_B6679_;
  assign new_B6656_ = new_B6622_ | new_B6655_;
  assign new_B6655_ = new_B6676_ | new_B6675_;
  assign new_B6654_ = ~new_B6634_ & ~new_B6644_;
  assign new_B6653_ = new_B6634_ & new_B6644_;
  assign new_B6652_ = ~new_B6634_ | new_B6644_;
  assign new_B6651_ = new_B6618_ & ~new_B6619_;
  assign new_B6650_ = ~new_B6618_ & new_B6619_;
  assign new_B6649_ = new_B6671_ & ~new_B6672_;
  assign new_B6648_ = ~new_B6671_ & new_B6672_;
  assign new_B6647_ = ~new_B6670_ | ~new_B6669_;
  assign new_B6646_ = new_B6662_ | new_B6661_;
  assign new_B6645_ = new_B6668_ | new_B6667_;
  assign new_B6644_ = new_B6658_ | new_B6660_;
  assign new_B6643_ = ~new_B6665_ | ~new_B6666_;
  assign new_B6642_ = new_B6618_ & ~new_B6619_;
  assign new_B6641_ = new_B6632_ & ~new_B6644_;
  assign new_B6640_ = ~new_B6632_ & new_B6644_;
  assign new_B6639_ = ~new_B6630_ & new_B6656_;
  assign new_B6638_ = new_B6654_ | new_B6653_;
  assign new_B6637_ = new_B6651_ | new_B6650_;
  assign new_B6636_ = new_B6619_ | new_B6652_;
  assign new_B6635_ = new_B6644_ & new_B6647_;
  assign new_B6634_ = new_B6649_ | new_B6648_;
  assign new_B6633_ = new_B6644_ & new_B6643_;
  assign new_B6632_ = new_B6646_ & new_B6645_;
  assign new_B6631_ = new_B6641_ | new_B6640_;
  assign new_B6630_ = new_B6619_ | new_B6642_;
  assign B6629 = new_B6630_ | new_B6639_;
  assign B6628 = new_B6637_ & new_B6638_;
  assign B6627 = new_B6637_ & new_B6636_;
  assign B6626 = new_B6635_ | new_B6634_;
  assign B6625 = new_B6633_ | new_B6632_;
  assign B6624 = new_B6631_ & new_B6630_;
  assign new_B6623_ = new_D900_;
  assign new_B6622_ = new_D833_;
  assign new_B6621_ = new_D766_;
  assign new_B6620_ = new_D699_;
  assign new_B6619_ = new_D632_;
  assign new_B6618_ = new_D565_;
  assign new_B6617_ = ~new_B6556_ & new_B6570_;
  assign new_B6616_ = new_B6556_ & ~new_B6570_;
  assign new_B6615_ = new_B6556_ & ~new_B6570_;
  assign new_B6614_ = ~new_B6556_ & ~new_B6570_;
  assign new_B6613_ = new_B6556_ & new_B6570_;
  assign new_B6612_ = new_B6616_ | new_B6617_;
  assign new_B6611_ = ~new_B6556_ & new_B6570_;
  assign new_B6610_ = new_B6614_ | new_B6615_;
  assign new_B6609_ = ~new_B6585_ & ~new_B6605_;
  assign new_B6608_ = new_B6585_ & new_B6605_;
  assign new_B6607_ = ~new_B6552_ | ~new_B6577_;
  assign new_B6606_ = new_B6570_ & new_B6607_;
  assign new_B6605_ = new_B6553_ | new_B6554_;
  assign new_B6604_ = new_B6553_ | new_B6570_;
  assign new_B6603_ = ~new_B6570_ & ~new_B6606_;
  assign new_B6602_ = new_B6570_ | new_B6607_;
  assign new_B6601_ = new_B6553_ & ~new_B6554_;
  assign new_B6600_ = ~new_B6553_ & new_B6554_;
  assign new_B6599_ = new_B6563_ | new_B6596_;
  assign new_B6598_ = ~new_B6563_ & ~new_B6597_;
  assign new_B6597_ = new_B6563_ & new_B6596_;
  assign new_B6596_ = ~new_B6552_ | ~new_B6577_;
  assign new_B6595_ = ~new_B6553_ & new_B6563_;
  assign new_B6594_ = new_B6553_ & ~new_B6563_;
  assign new_B6593_ = new_B6555_ & new_B6592_;
  assign new_B6592_ = new_B6611_ | new_B6610_;
  assign new_B6591_ = ~new_B6555_ & new_B6590_;
  assign new_B6590_ = new_B6613_ | new_B6612_;
  assign new_B6589_ = new_B6555_ | new_B6588_;
  assign new_B6588_ = new_B6609_ | new_B6608_;
  assign new_B6587_ = ~new_B6567_ & ~new_B6577_;
  assign new_B6586_ = new_B6567_ & new_B6577_;
  assign new_B6585_ = ~new_B6567_ | new_B6577_;
  assign new_B6584_ = new_B6551_ & ~new_B6552_;
  assign new_B6583_ = ~new_B6551_ & new_B6552_;
  assign new_B6582_ = new_B6604_ & ~new_B6605_;
  assign new_B6581_ = ~new_B6604_ & new_B6605_;
  assign new_B6580_ = ~new_B6603_ | ~new_B6602_;
  assign new_B6579_ = new_B6595_ | new_B6594_;
  assign new_B6578_ = new_B6601_ | new_B6600_;
  assign new_B6577_ = new_B6591_ | new_B6593_;
  assign new_B6576_ = ~new_B6598_ | ~new_B6599_;
  assign new_B6575_ = new_B6551_ & ~new_B6552_;
  assign new_B6574_ = new_B6565_ & ~new_B6577_;
  assign new_B6573_ = ~new_B6565_ & new_B6577_;
  assign new_B6572_ = ~new_B6563_ & new_B6589_;
  assign new_B6571_ = new_B6587_ | new_B6586_;
  assign new_B6570_ = new_B6584_ | new_B6583_;
  assign new_B6569_ = new_B6552_ | new_B6585_;
  assign new_B6568_ = new_B6577_ & new_B6580_;
  assign new_B6567_ = new_B6582_ | new_B6581_;
  assign new_B6566_ = new_B6577_ & new_B6576_;
  assign new_B6565_ = new_B6579_ & new_B6578_;
  assign new_B6564_ = new_B6574_ | new_B6573_;
  assign new_B6563_ = new_B6552_ | new_B6575_;
  assign B6562 = new_B6563_ | new_B6572_;
  assign B6561 = new_B6570_ & new_B6571_;
  assign B6560 = new_B6570_ & new_B6569_;
  assign B6559 = new_B6568_ | new_B6567_;
  assign B6558 = new_B6566_ | new_B6565_;
  assign B6557 = new_B6564_ & new_B6563_;
  assign new_B6556_ = new_D498_;
  assign new_B6555_ = new_D431_;
  assign new_B6554_ = new_D364_;
  assign new_B6553_ = new_D297_;
  assign new_B6552_ = new_D230_;
  assign new_B6551_ = new_D163_;
  assign new_B6550_ = ~new_B6489_ & new_B6503_;
  assign new_B6549_ = new_B6489_ & ~new_B6503_;
  assign new_B6548_ = new_B6489_ & ~new_B6503_;
  assign new_B6547_ = ~new_B6489_ & ~new_B6503_;
  assign new_B6546_ = new_B6489_ & new_B6503_;
  assign new_B6545_ = new_B6549_ | new_B6550_;
  assign new_B6544_ = ~new_B6489_ & new_B6503_;
  assign new_B6543_ = new_B6547_ | new_B6548_;
  assign new_B6542_ = ~new_B6518_ & ~new_B6538_;
  assign new_B6541_ = new_B6518_ & new_B6538_;
  assign new_B6540_ = ~new_B6485_ | ~new_B6510_;
  assign new_B6539_ = new_B6503_ & new_B6540_;
  assign new_B6538_ = new_B6486_ | new_B6487_;
  assign new_B6537_ = new_B6486_ | new_B6503_;
  assign new_B6536_ = ~new_B6503_ & ~new_B6539_;
  assign new_B6535_ = new_B6503_ | new_B6540_;
  assign new_B6534_ = new_B6486_ & ~new_B6487_;
  assign new_B6533_ = ~new_B6486_ & new_B6487_;
  assign new_B6532_ = new_B6496_ | new_B6529_;
  assign new_B6531_ = ~new_B6496_ & ~new_B6530_;
  assign new_B6530_ = new_B6496_ & new_B6529_;
  assign new_B6529_ = ~new_B6485_ | ~new_B6510_;
  assign new_B6528_ = ~new_B6486_ & new_B6496_;
  assign new_B6527_ = new_B6486_ & ~new_B6496_;
  assign new_B6526_ = new_B6488_ & new_B6525_;
  assign new_B6525_ = new_B6544_ | new_B6543_;
  assign new_B6524_ = ~new_B6488_ & new_B6523_;
  assign new_B6523_ = new_B6546_ | new_B6545_;
  assign new_B6522_ = new_B6488_ | new_B6521_;
  assign new_B6521_ = new_B6542_ | new_B6541_;
  assign new_B6520_ = ~new_B6500_ & ~new_B6510_;
  assign new_B6519_ = new_B6500_ & new_B6510_;
  assign new_B6518_ = ~new_B6500_ | new_B6510_;
  assign new_B6517_ = new_B6484_ & ~new_B6485_;
  assign new_B6516_ = ~new_B6484_ & new_B6485_;
  assign new_B6515_ = new_B6537_ & ~new_B6538_;
  assign new_B6514_ = ~new_B6537_ & new_B6538_;
  assign new_B6513_ = ~new_B6536_ | ~new_B6535_;
  assign new_B6512_ = new_B6528_ | new_B6527_;
  assign new_B6511_ = new_B6534_ | new_B6533_;
  assign new_B6510_ = new_B6524_ | new_B6526_;
  assign new_B6509_ = ~new_B6531_ | ~new_B6532_;
  assign new_B6508_ = new_B6484_ & ~new_B6485_;
  assign new_B6507_ = new_B6498_ & ~new_B6510_;
  assign new_B6506_ = ~new_B6498_ & new_B6510_;
  assign new_B6505_ = ~new_B6496_ & new_B6522_;
  assign new_B6504_ = new_B6520_ | new_B6519_;
  assign new_B6503_ = new_B6517_ | new_B6516_;
  assign new_B6502_ = new_B6485_ | new_B6518_;
  assign new_B6501_ = new_B6510_ & new_B6513_;
  assign new_B6500_ = new_B6515_ | new_B6514_;
  assign new_B6499_ = new_B6510_ & new_B6509_;
  assign new_B6498_ = new_B6512_ & new_B6511_;
  assign new_B6497_ = new_B6507_ | new_B6506_;
  assign new_B6496_ = new_B6485_ | new_B6508_;
  assign B6495 = new_B6496_ | new_B6505_;
  assign B6494 = new_B6503_ & new_B6504_;
  assign B6493 = new_B6503_ & new_B6502_;
  assign B6492 = new_B6501_ | new_B6500_;
  assign B6491 = new_B6499_ | new_B6498_;
  assign B6490 = new_B6497_ & new_B6496_;
  assign new_B6489_ = new_D96_;
  assign new_B6488_ = new_D29_;
  assign new_B6487_ = new_C9961_;
  assign new_B6486_ = new_C9894_;
  assign new_B6485_ = new_C9827_;
  assign new_B6484_ = new_C9760_;
  assign new_B6483_ = ~new_B6422_ & new_B6436_;
  assign new_B6482_ = new_B6422_ & ~new_B6436_;
  assign new_B6481_ = new_B6422_ & ~new_B6436_;
  assign new_B6480_ = ~new_B6422_ & ~new_B6436_;
  assign new_B6479_ = new_B6422_ & new_B6436_;
  assign new_B6478_ = new_B6482_ | new_B6483_;
  assign new_B6477_ = ~new_B6422_ & new_B6436_;
  assign new_B6476_ = new_B6480_ | new_B6481_;
  assign new_B6475_ = ~new_B6451_ & ~new_B6471_;
  assign new_B6474_ = new_B6451_ & new_B6471_;
  assign new_B6473_ = ~new_B6418_ | ~new_B6443_;
  assign new_B6472_ = new_B6436_ & new_B6473_;
  assign new_B6471_ = new_B6419_ | new_B6420_;
  assign new_B6470_ = new_B6419_ | new_B6436_;
  assign new_B6469_ = ~new_B6436_ & ~new_B6472_;
  assign new_B6468_ = new_B6436_ | new_B6473_;
  assign new_B6467_ = new_B6419_ & ~new_B6420_;
  assign new_B6466_ = ~new_B6419_ & new_B6420_;
  assign new_B6465_ = new_B6429_ | new_B6462_;
  assign new_B6464_ = ~new_B6429_ & ~new_B6463_;
  assign new_B6463_ = new_B6429_ & new_B6462_;
  assign new_B6462_ = ~new_B6418_ | ~new_B6443_;
  assign new_B6461_ = ~new_B6419_ & new_B6429_;
  assign new_B6460_ = new_B6419_ & ~new_B6429_;
  assign new_B6459_ = new_B6421_ & new_B6458_;
  assign new_B6458_ = new_B6477_ | new_B6476_;
  assign new_B6457_ = ~new_B6421_ & new_B6456_;
  assign new_B6456_ = new_B6479_ | new_B6478_;
  assign new_B6455_ = new_B6421_ | new_B6454_;
  assign new_B6454_ = new_B6475_ | new_B6474_;
  assign new_B6453_ = ~new_B6433_ & ~new_B6443_;
  assign new_B6452_ = new_B6433_ & new_B6443_;
  assign new_B6451_ = ~new_B6433_ | new_B6443_;
  assign new_B6450_ = new_B6417_ & ~new_B6418_;
  assign new_B6449_ = ~new_B6417_ & new_B6418_;
  assign new_B6448_ = new_B6470_ & ~new_B6471_;
  assign new_B6447_ = ~new_B6470_ & new_B6471_;
  assign new_B6446_ = ~new_B6469_ | ~new_B6468_;
  assign new_B6445_ = new_B6461_ | new_B6460_;
  assign new_B6444_ = new_B6467_ | new_B6466_;
  assign new_B6443_ = new_B6457_ | new_B6459_;
  assign new_B6442_ = ~new_B6464_ | ~new_B6465_;
  assign new_B6441_ = new_B6417_ & ~new_B6418_;
  assign new_B6440_ = new_B6431_ & ~new_B6443_;
  assign new_B6439_ = ~new_B6431_ & new_B6443_;
  assign new_B6438_ = ~new_B6429_ & new_B6455_;
  assign new_B6437_ = new_B6453_ | new_B6452_;
  assign new_B6436_ = new_B6450_ | new_B6449_;
  assign new_B6435_ = new_B6418_ | new_B6451_;
  assign new_B6434_ = new_B6443_ & new_B6446_;
  assign new_B6433_ = new_B6448_ | new_B6447_;
  assign new_B6432_ = new_B6443_ & new_B6442_;
  assign new_B6431_ = new_B6445_ & new_B6444_;
  assign new_B6430_ = new_B6440_ | new_B6439_;
  assign new_B6429_ = new_B6418_ | new_B6441_;
  assign B6428 = new_B6429_ | new_B6438_;
  assign B6427 = new_B6436_ & new_B6437_;
  assign B6426 = new_B6436_ & new_B6435_;
  assign B6425 = new_B6434_ | new_B6433_;
  assign B6424 = new_B6432_ | new_B6431_;
  assign B6423 = new_B6430_ & new_B6429_;
  assign new_B6422_ = new_C9693_;
  assign new_B6421_ = new_C9626_;
  assign new_B6420_ = new_C9559_;
  assign new_B6419_ = new_C9492_;
  assign new_B6418_ = new_C9425_;
  assign new_B6417_ = new_C9358_;
  assign new_B6416_ = ~new_B6355_ & new_B6369_;
  assign new_B6415_ = new_B6355_ & ~new_B6369_;
  assign new_B6414_ = new_B6355_ & ~new_B6369_;
  assign new_B6413_ = ~new_B6355_ & ~new_B6369_;
  assign new_B6412_ = new_B6355_ & new_B6369_;
  assign new_B6411_ = new_B6415_ | new_B6416_;
  assign new_B6410_ = ~new_B6355_ & new_B6369_;
  assign new_B6409_ = new_B6413_ | new_B6414_;
  assign new_B6408_ = ~new_B6384_ & ~new_B6404_;
  assign new_B6407_ = new_B6384_ & new_B6404_;
  assign new_B6406_ = ~new_B6351_ | ~new_B6376_;
  assign new_B6405_ = new_B6369_ & new_B6406_;
  assign new_B6404_ = new_B6352_ | new_B6353_;
  assign new_B6403_ = new_B6352_ | new_B6369_;
  assign new_B6402_ = ~new_B6369_ & ~new_B6405_;
  assign new_B6401_ = new_B6369_ | new_B6406_;
  assign new_B6400_ = new_B6352_ & ~new_B6353_;
  assign new_B6399_ = ~new_B6352_ & new_B6353_;
  assign new_B6398_ = new_B6362_ | new_B6395_;
  assign new_B6397_ = ~new_B6362_ & ~new_B6396_;
  assign new_B6396_ = new_B6362_ & new_B6395_;
  assign new_B6395_ = ~new_B6351_ | ~new_B6376_;
  assign new_B6394_ = ~new_B6352_ & new_B6362_;
  assign new_B6393_ = new_B6352_ & ~new_B6362_;
  assign new_B6392_ = new_B6354_ & new_B6391_;
  assign new_B6391_ = new_B6410_ | new_B6409_;
  assign new_B6390_ = ~new_B6354_ & new_B6389_;
  assign new_B6389_ = new_B6412_ | new_B6411_;
  assign new_B6388_ = new_B6354_ | new_B6387_;
  assign new_B6387_ = new_B6408_ | new_B6407_;
  assign new_B6386_ = ~new_B6366_ & ~new_B6376_;
  assign new_B6385_ = new_B6366_ & new_B6376_;
  assign new_B6384_ = ~new_B6366_ | new_B6376_;
  assign new_B6383_ = new_B6350_ & ~new_B6351_;
  assign new_B6382_ = ~new_B6350_ & new_B6351_;
  assign new_B6381_ = new_B6403_ & ~new_B6404_;
  assign new_B6380_ = ~new_B6403_ & new_B6404_;
  assign new_B6379_ = ~new_B6402_ | ~new_B6401_;
  assign new_B6378_ = new_B6394_ | new_B6393_;
  assign new_B6377_ = new_B6400_ | new_B6399_;
  assign new_B6376_ = new_B6390_ | new_B6392_;
  assign new_B6375_ = ~new_B6397_ | ~new_B6398_;
  assign new_B6374_ = new_B6350_ & ~new_B6351_;
  assign new_B6373_ = new_B6364_ & ~new_B6376_;
  assign new_B6372_ = ~new_B6364_ & new_B6376_;
  assign new_B6371_ = ~new_B6362_ & new_B6388_;
  assign new_B6370_ = new_B6386_ | new_B6385_;
  assign new_B6369_ = new_B6383_ | new_B6382_;
  assign new_B6368_ = new_B6351_ | new_B6384_;
  assign new_B6367_ = new_B6376_ & new_B6379_;
  assign new_B6366_ = new_B6381_ | new_B6380_;
  assign new_B6365_ = new_B6376_ & new_B6375_;
  assign new_B6364_ = new_B6378_ & new_B6377_;
  assign new_B6363_ = new_B6373_ | new_B6372_;
  assign new_B6362_ = new_B6351_ | new_B6374_;
  assign B6361 = new_B6362_ | new_B6371_;
  assign B6360 = new_B6369_ & new_B6370_;
  assign B6359 = new_B6369_ & new_B6368_;
  assign B6358 = new_B6367_ | new_B6366_;
  assign B6357 = new_B6365_ | new_B6364_;
  assign B6356 = new_B6363_ & new_B6362_;
  assign new_B6355_ = new_C9291_;
  assign new_B6354_ = new_C9224_;
  assign new_B6353_ = new_C9157_;
  assign new_B6352_ = new_C9090_;
  assign new_B6351_ = new_C9023_;
  assign new_B6350_ = new_C8956_;
  assign new_B6349_ = ~new_B6288_ & new_B6302_;
  assign new_B6348_ = new_B6288_ & ~new_B6302_;
  assign new_B6347_ = new_B6288_ & ~new_B6302_;
  assign new_B6346_ = ~new_B6288_ & ~new_B6302_;
  assign new_B6345_ = new_B6288_ & new_B6302_;
  assign new_B6344_ = new_B6348_ | new_B6349_;
  assign new_B6343_ = ~new_B6288_ & new_B6302_;
  assign new_B6342_ = new_B6346_ | new_B6347_;
  assign new_B6341_ = ~new_B6317_ & ~new_B6337_;
  assign new_B6340_ = new_B6317_ & new_B6337_;
  assign new_B6339_ = ~new_B6284_ | ~new_B6309_;
  assign new_B6338_ = new_B6302_ & new_B6339_;
  assign new_B6337_ = new_B6285_ | new_B6286_;
  assign new_B6336_ = new_B6285_ | new_B6302_;
  assign new_B6335_ = ~new_B6302_ & ~new_B6338_;
  assign new_B6334_ = new_B6302_ | new_B6339_;
  assign new_B6333_ = new_B6285_ & ~new_B6286_;
  assign new_B6332_ = ~new_B6285_ & new_B6286_;
  assign new_B6331_ = new_B6295_ | new_B6328_;
  assign new_B6330_ = ~new_B6295_ & ~new_B6329_;
  assign new_B6329_ = new_B6295_ & new_B6328_;
  assign new_B6328_ = ~new_B6284_ | ~new_B6309_;
  assign new_B6327_ = ~new_B6285_ & new_B6295_;
  assign new_B6326_ = new_B6285_ & ~new_B6295_;
  assign new_B6325_ = new_B6287_ & new_B6324_;
  assign new_B6324_ = new_B6343_ | new_B6342_;
  assign new_B6323_ = ~new_B6287_ & new_B6322_;
  assign new_B6322_ = new_B6345_ | new_B6344_;
  assign new_B6321_ = new_B6287_ | new_B6320_;
  assign new_B6320_ = new_B6341_ | new_B6340_;
  assign new_B6319_ = ~new_B6299_ & ~new_B6309_;
  assign new_B6318_ = new_B6299_ & new_B6309_;
  assign new_B6317_ = ~new_B6299_ | new_B6309_;
  assign new_B6316_ = new_B6283_ & ~new_B6284_;
  assign new_B6315_ = ~new_B6283_ & new_B6284_;
  assign new_B6314_ = new_B6336_ & ~new_B6337_;
  assign new_B6313_ = ~new_B6336_ & new_B6337_;
  assign new_B6312_ = ~new_B6335_ | ~new_B6334_;
  assign new_B6311_ = new_B6327_ | new_B6326_;
  assign new_B6310_ = new_B6333_ | new_B6332_;
  assign new_B6309_ = new_B6323_ | new_B6325_;
  assign new_B6308_ = ~new_B6330_ | ~new_B6331_;
  assign new_B6307_ = new_B6283_ & ~new_B6284_;
  assign new_B6306_ = new_B6297_ & ~new_B6309_;
  assign new_B6305_ = ~new_B6297_ & new_B6309_;
  assign new_B6304_ = ~new_B6295_ & new_B6321_;
  assign new_B6303_ = new_B6319_ | new_B6318_;
  assign new_B6302_ = new_B6316_ | new_B6315_;
  assign new_B6301_ = new_B6284_ | new_B6317_;
  assign new_B6300_ = new_B6309_ & new_B6312_;
  assign new_B6299_ = new_B6314_ | new_B6313_;
  assign new_B6298_ = new_B6309_ & new_B6308_;
  assign new_B6297_ = new_B6311_ & new_B6310_;
  assign new_B6296_ = new_B6306_ | new_B6305_;
  assign new_B6295_ = new_B6284_ | new_B6307_;
  assign B6294 = new_B6295_ | new_B6304_;
  assign B6293 = new_B6302_ & new_B6303_;
  assign B6292 = new_B6302_ & new_B6301_;
  assign B6291 = new_B6300_ | new_B6299_;
  assign B6290 = new_B6298_ | new_B6297_;
  assign B6289 = new_B6296_ & new_B6295_;
  assign new_B6288_ = new_C8889_;
  assign new_B6287_ = new_C8822_;
  assign new_B6286_ = new_C8755_;
  assign new_B6285_ = new_C8688_;
  assign new_B6284_ = new_C8621_;
  assign new_B6283_ = new_C8554_;
  assign new_B6282_ = ~new_B6221_ & new_B6235_;
  assign new_B6281_ = new_B6221_ & ~new_B6235_;
  assign new_B6280_ = new_B6221_ & ~new_B6235_;
  assign new_B6279_ = ~new_B6221_ & ~new_B6235_;
  assign new_B6278_ = new_B6221_ & new_B6235_;
  assign new_B6277_ = new_B6281_ | new_B6282_;
  assign new_B6276_ = ~new_B6221_ & new_B6235_;
  assign new_B6275_ = new_B6279_ | new_B6280_;
  assign new_B6274_ = ~new_B6250_ & ~new_B6270_;
  assign new_B6273_ = new_B6250_ & new_B6270_;
  assign new_B6272_ = ~new_B6217_ | ~new_B6242_;
  assign new_B6271_ = new_B6235_ & new_B6272_;
  assign new_B6270_ = new_B6218_ | new_B6219_;
  assign new_B6269_ = new_B6218_ | new_B6235_;
  assign new_B6268_ = ~new_B6235_ & ~new_B6271_;
  assign new_B6267_ = new_B6235_ | new_B6272_;
  assign new_B6266_ = new_B6218_ & ~new_B6219_;
  assign new_B6265_ = ~new_B6218_ & new_B6219_;
  assign new_B6264_ = new_B6228_ | new_B6261_;
  assign new_B6263_ = ~new_B6228_ & ~new_B6262_;
  assign new_B6262_ = new_B6228_ & new_B6261_;
  assign new_B6261_ = ~new_B6217_ | ~new_B6242_;
  assign new_B6260_ = ~new_B6218_ & new_B6228_;
  assign new_B6259_ = new_B6218_ & ~new_B6228_;
  assign new_B6258_ = new_B6220_ & new_B6257_;
  assign new_B6257_ = new_B6276_ | new_B6275_;
  assign new_B6256_ = ~new_B6220_ & new_B6255_;
  assign new_B6255_ = new_B6278_ | new_B6277_;
  assign new_B6254_ = new_B6220_ | new_B6253_;
  assign new_B6253_ = new_B6274_ | new_B6273_;
  assign new_B6252_ = ~new_B6232_ & ~new_B6242_;
  assign new_B6251_ = new_B6232_ & new_B6242_;
  assign new_B6250_ = ~new_B6232_ | new_B6242_;
  assign new_B6249_ = new_B6216_ & ~new_B6217_;
  assign new_B6248_ = ~new_B6216_ & new_B6217_;
  assign new_B6247_ = new_B6269_ & ~new_B6270_;
  assign new_B6246_ = ~new_B6269_ & new_B6270_;
  assign new_B6245_ = ~new_B6268_ | ~new_B6267_;
  assign new_B6244_ = new_B6260_ | new_B6259_;
  assign new_B6243_ = new_B6266_ | new_B6265_;
  assign new_B6242_ = new_B6256_ | new_B6258_;
  assign new_B6241_ = ~new_B6263_ | ~new_B6264_;
  assign new_B6240_ = new_B6216_ & ~new_B6217_;
  assign new_B6239_ = new_B6230_ & ~new_B6242_;
  assign new_B6238_ = ~new_B6230_ & new_B6242_;
  assign new_B6237_ = ~new_B6228_ & new_B6254_;
  assign new_B6236_ = new_B6252_ | new_B6251_;
  assign new_B6235_ = new_B6249_ | new_B6248_;
  assign new_B6234_ = new_B6217_ | new_B6250_;
  assign new_B6233_ = new_B6242_ & new_B6245_;
  assign new_B6232_ = new_B6247_ | new_B6246_;
  assign new_B6231_ = new_B6242_ & new_B6241_;
  assign new_B6230_ = new_B6244_ & new_B6243_;
  assign new_B6229_ = new_B6239_ | new_B6238_;
  assign new_B6228_ = new_B6217_ | new_B6240_;
  assign B6227 = new_B6228_ | new_B6237_;
  assign B6226 = new_B6235_ & new_B6236_;
  assign B6225 = new_B6235_ & new_B6234_;
  assign B6224 = new_B6233_ | new_B6232_;
  assign B6223 = new_B6231_ | new_B6230_;
  assign B6222 = new_B6229_ & new_B6228_;
  assign new_B6221_ = new_C8487_;
  assign new_B6220_ = new_C8420_;
  assign new_B6219_ = new_C8353_;
  assign new_B6218_ = new_C8286_;
  assign new_B6217_ = new_C8219_;
  assign new_B6216_ = new_C8152_;
  assign new_B6215_ = ~new_B6154_ & new_B6168_;
  assign new_B6214_ = new_B6154_ & ~new_B6168_;
  assign new_B6213_ = new_B6154_ & ~new_B6168_;
  assign new_B6212_ = ~new_B6154_ & ~new_B6168_;
  assign new_B6211_ = new_B6154_ & new_B6168_;
  assign new_B6210_ = new_B6214_ | new_B6215_;
  assign new_B6209_ = ~new_B6154_ & new_B6168_;
  assign new_B6208_ = new_B6212_ | new_B6213_;
  assign new_B6207_ = ~new_B6183_ & ~new_B6203_;
  assign new_B6206_ = new_B6183_ & new_B6203_;
  assign new_B6205_ = ~new_B6150_ | ~new_B6175_;
  assign new_B6204_ = new_B6168_ & new_B6205_;
  assign new_B6203_ = new_B6151_ | new_B6152_;
  assign new_B6202_ = new_B6151_ | new_B6168_;
  assign new_B6201_ = ~new_B6168_ & ~new_B6204_;
  assign new_B6200_ = new_B6168_ | new_B6205_;
  assign new_B6199_ = new_B6151_ & ~new_B6152_;
  assign new_B6198_ = ~new_B6151_ & new_B6152_;
  assign new_B6197_ = new_B6161_ | new_B6194_;
  assign new_B6196_ = ~new_B6161_ & ~new_B6195_;
  assign new_B6195_ = new_B6161_ & new_B6194_;
  assign new_B6194_ = ~new_B6150_ | ~new_B6175_;
  assign new_B6193_ = ~new_B6151_ & new_B6161_;
  assign new_B6192_ = new_B6151_ & ~new_B6161_;
  assign new_B6191_ = new_B6153_ & new_B6190_;
  assign new_B6190_ = new_B6209_ | new_B6208_;
  assign new_B6189_ = ~new_B6153_ & new_B6188_;
  assign new_B6188_ = new_B6211_ | new_B6210_;
  assign new_B6187_ = new_B6153_ | new_B6186_;
  assign new_B6186_ = new_B6207_ | new_B6206_;
  assign new_B6185_ = ~new_B6165_ & ~new_B6175_;
  assign new_B6184_ = new_B6165_ & new_B6175_;
  assign new_B6183_ = ~new_B6165_ | new_B6175_;
  assign new_B6182_ = new_B6149_ & ~new_B6150_;
  assign new_B6181_ = ~new_B6149_ & new_B6150_;
  assign new_B6180_ = new_B6202_ & ~new_B6203_;
  assign new_B6179_ = ~new_B6202_ & new_B6203_;
  assign new_B6178_ = ~new_B6201_ | ~new_B6200_;
  assign new_B6177_ = new_B6193_ | new_B6192_;
  assign new_B6176_ = new_B6199_ | new_B6198_;
  assign new_B6175_ = new_B6189_ | new_B6191_;
  assign new_B6174_ = ~new_B6196_ | ~new_B6197_;
  assign new_B6173_ = new_B6149_ & ~new_B6150_;
  assign new_B6172_ = new_B6163_ & ~new_B6175_;
  assign new_B6171_ = ~new_B6163_ & new_B6175_;
  assign new_B6170_ = ~new_B6161_ & new_B6187_;
  assign new_B6169_ = new_B6185_ | new_B6184_;
  assign new_B6168_ = new_B6182_ | new_B6181_;
  assign new_B6167_ = new_B6150_ | new_B6183_;
  assign new_B6166_ = new_B6175_ & new_B6178_;
  assign new_B6165_ = new_B6180_ | new_B6179_;
  assign new_B6164_ = new_B6175_ & new_B6174_;
  assign new_B6163_ = new_B6177_ & new_B6176_;
  assign new_B6162_ = new_B6172_ | new_B6171_;
  assign new_B6161_ = new_B6150_ | new_B6173_;
  assign B6160 = new_B6161_ | new_B6170_;
  assign B6159 = new_B6168_ & new_B6169_;
  assign B6158 = new_B6168_ & new_B6167_;
  assign B6157 = new_B6166_ | new_B6165_;
  assign B6156 = new_B6164_ | new_B6163_;
  assign B6155 = new_B6162_ & new_B6161_;
  assign new_B6154_ = new_C8085_;
  assign new_B6153_ = new_C8018_;
  assign new_B6152_ = new_C7951_;
  assign new_B6151_ = new_C7884_;
  assign new_B6150_ = new_C7817_;
  assign new_B6149_ = new_C7750_;
  assign new_B6148_ = ~new_B6087_ & new_B6101_;
  assign new_B6147_ = new_B6087_ & ~new_B6101_;
  assign new_B6146_ = new_B6087_ & ~new_B6101_;
  assign new_B6145_ = ~new_B6087_ & ~new_B6101_;
  assign new_B6144_ = new_B6087_ & new_B6101_;
  assign new_B6143_ = new_B6147_ | new_B6148_;
  assign new_B6142_ = ~new_B6087_ & new_B6101_;
  assign new_B6141_ = new_B6145_ | new_B6146_;
  assign new_B6140_ = ~new_B6116_ & ~new_B6136_;
  assign new_B6139_ = new_B6116_ & new_B6136_;
  assign new_B6138_ = ~new_B6083_ | ~new_B6108_;
  assign new_B6137_ = new_B6101_ & new_B6138_;
  assign new_B6136_ = new_B6084_ | new_B6085_;
  assign new_B6135_ = new_B6084_ | new_B6101_;
  assign new_B6134_ = ~new_B6101_ & ~new_B6137_;
  assign new_B6133_ = new_B6101_ | new_B6138_;
  assign new_B6132_ = new_B6084_ & ~new_B6085_;
  assign new_B6131_ = ~new_B6084_ & new_B6085_;
  assign new_B6130_ = new_B6094_ | new_B6127_;
  assign new_B6129_ = ~new_B6094_ & ~new_B6128_;
  assign new_B6128_ = new_B6094_ & new_B6127_;
  assign new_B6127_ = ~new_B6083_ | ~new_B6108_;
  assign new_B6126_ = ~new_B6084_ & new_B6094_;
  assign new_B6125_ = new_B6084_ & ~new_B6094_;
  assign new_B6124_ = new_B6086_ & new_B6123_;
  assign new_B6123_ = new_B6142_ | new_B6141_;
  assign new_B6122_ = ~new_B6086_ & new_B6121_;
  assign new_B6121_ = new_B6144_ | new_B6143_;
  assign new_B6120_ = new_B6086_ | new_B6119_;
  assign new_B6119_ = new_B6140_ | new_B6139_;
  assign new_B6118_ = ~new_B6098_ & ~new_B6108_;
  assign new_B6117_ = new_B6098_ & new_B6108_;
  assign new_B6116_ = ~new_B6098_ | new_B6108_;
  assign new_B6115_ = new_B6082_ & ~new_B6083_;
  assign new_B6114_ = ~new_B6082_ & new_B6083_;
  assign new_B6113_ = new_B6135_ & ~new_B6136_;
  assign new_B6112_ = ~new_B6135_ & new_B6136_;
  assign new_B6111_ = ~new_B6134_ | ~new_B6133_;
  assign new_B6110_ = new_B6126_ | new_B6125_;
  assign new_B6109_ = new_B6132_ | new_B6131_;
  assign new_B6108_ = new_B6122_ | new_B6124_;
  assign new_B6107_ = ~new_B6129_ | ~new_B6130_;
  assign new_B6106_ = new_B6082_ & ~new_B6083_;
  assign new_B6105_ = new_B6096_ & ~new_B6108_;
  assign new_B6104_ = ~new_B6096_ & new_B6108_;
  assign new_B6103_ = ~new_B6094_ & new_B6120_;
  assign new_B6102_ = new_B6118_ | new_B6117_;
  assign new_B6101_ = new_B6115_ | new_B6114_;
  assign new_B6100_ = new_B6083_ | new_B6116_;
  assign new_B6099_ = new_B6108_ & new_B6111_;
  assign new_B6098_ = new_B6113_ | new_B6112_;
  assign new_B6097_ = new_B6108_ & new_B6107_;
  assign new_B6096_ = new_B6110_ & new_B6109_;
  assign new_B6095_ = new_B6105_ | new_B6104_;
  assign new_B6094_ = new_B6083_ | new_B6106_;
  assign B6093 = new_B6094_ | new_B6103_;
  assign B6092 = new_B6101_ & new_B6102_;
  assign B6091 = new_B6101_ & new_B6100_;
  assign B6090 = new_B6099_ | new_B6098_;
  assign B6089 = new_B6097_ | new_B6096_;
  assign B6088 = new_B6095_ & new_B6094_;
  assign new_B6087_ = new_C7683_;
  assign new_B6086_ = new_C7616_;
  assign new_B6085_ = new_C7549_;
  assign new_B6084_ = new_C7482_;
  assign new_B6083_ = new_C7415_;
  assign new_B6082_ = new_C7348_;
  assign new_B6081_ = ~new_B6020_ & new_B6034_;
  assign new_B6080_ = new_B6020_ & ~new_B6034_;
  assign new_B6079_ = new_B6020_ & ~new_B6034_;
  assign new_B6078_ = ~new_B6020_ & ~new_B6034_;
  assign new_B6077_ = new_B6020_ & new_B6034_;
  assign new_B6076_ = new_B6080_ | new_B6081_;
  assign new_B6075_ = ~new_B6020_ & new_B6034_;
  assign new_B6074_ = new_B6078_ | new_B6079_;
  assign new_B6073_ = ~new_B6049_ & ~new_B6069_;
  assign new_B6072_ = new_B6049_ & new_B6069_;
  assign new_B6071_ = ~new_B6016_ | ~new_B6041_;
  assign new_B6070_ = new_B6034_ & new_B6071_;
  assign new_B6069_ = new_B6017_ | new_B6018_;
  assign new_B6068_ = new_B6017_ | new_B6034_;
  assign new_B6067_ = ~new_B6034_ & ~new_B6070_;
  assign new_B6066_ = new_B6034_ | new_B6071_;
  assign new_B6065_ = new_B6017_ & ~new_B6018_;
  assign new_B6064_ = ~new_B6017_ & new_B6018_;
  assign new_B6063_ = new_B6027_ | new_B6060_;
  assign new_B6062_ = ~new_B6027_ & ~new_B6061_;
  assign new_B6061_ = new_B6027_ & new_B6060_;
  assign new_B6060_ = ~new_B6016_ | ~new_B6041_;
  assign new_B6059_ = ~new_B6017_ & new_B6027_;
  assign new_B6058_ = new_B6017_ & ~new_B6027_;
  assign new_B6057_ = new_B6019_ & new_B6056_;
  assign new_B6056_ = new_B6075_ | new_B6074_;
  assign new_B6055_ = ~new_B6019_ & new_B6054_;
  assign new_B6054_ = new_B6077_ | new_B6076_;
  assign new_B6053_ = new_B6019_ | new_B6052_;
  assign new_B6052_ = new_B6073_ | new_B6072_;
  assign new_B6051_ = ~new_B6031_ & ~new_B6041_;
  assign new_B6050_ = new_B6031_ & new_B6041_;
  assign new_B6049_ = ~new_B6031_ | new_B6041_;
  assign new_B6048_ = new_B6015_ & ~new_B6016_;
  assign new_B6047_ = ~new_B6015_ & new_B6016_;
  assign new_B6046_ = new_B6068_ & ~new_B6069_;
  assign new_B6045_ = ~new_B6068_ & new_B6069_;
  assign new_B6044_ = ~new_B6067_ | ~new_B6066_;
  assign new_B6043_ = new_B6059_ | new_B6058_;
  assign new_B6042_ = new_B6065_ | new_B6064_;
  assign new_B6041_ = new_B6055_ | new_B6057_;
  assign new_B6040_ = ~new_B6062_ | ~new_B6063_;
  assign new_B6039_ = new_B6015_ & ~new_B6016_;
  assign new_B6038_ = new_B6029_ & ~new_B6041_;
  assign new_B6037_ = ~new_B6029_ & new_B6041_;
  assign new_B6036_ = ~new_B6027_ & new_B6053_;
  assign new_B6035_ = new_B6051_ | new_B6050_;
  assign new_B6034_ = new_B6048_ | new_B6047_;
  assign new_B6033_ = new_B6016_ | new_B6049_;
  assign new_B6032_ = new_B6041_ & new_B6044_;
  assign new_B6031_ = new_B6046_ | new_B6045_;
  assign new_B6030_ = new_B6041_ & new_B6040_;
  assign new_B6029_ = new_B6043_ & new_B6042_;
  assign new_B6028_ = new_B6038_ | new_B6037_;
  assign new_B6027_ = new_B6016_ | new_B6039_;
  assign B6026 = new_B6027_ | new_B6036_;
  assign B6025 = new_B6034_ & new_B6035_;
  assign B6024 = new_B6034_ & new_B6033_;
  assign B6023 = new_B6032_ | new_B6031_;
  assign B6022 = new_B6030_ | new_B6029_;
  assign B6021 = new_B6028_ & new_B6027_;
  assign new_B6020_ = new_C7281_;
  assign new_B6019_ = new_C7214_;
  assign new_B6018_ = new_C7147_;
  assign new_B6017_ = new_C7080_;
  assign new_B6016_ = new_C7013_;
  assign new_B6015_ = new_C6946_;
  assign new_B6014_ = ~new_B5953_ & new_B5967_;
  assign new_B6013_ = new_B5953_ & ~new_B5967_;
  assign new_B6012_ = new_B5953_ & ~new_B5967_;
  assign new_B6011_ = ~new_B5953_ & ~new_B5967_;
  assign new_B6010_ = new_B5953_ & new_B5967_;
  assign new_B6009_ = new_B6013_ | new_B6014_;
  assign new_B6008_ = ~new_B5953_ & new_B5967_;
  assign new_B6007_ = new_B6011_ | new_B6012_;
  assign new_B6006_ = ~new_B5982_ & ~new_B6002_;
  assign new_B6005_ = new_B5982_ & new_B6002_;
  assign new_B6004_ = ~new_B5949_ | ~new_B5974_;
  assign new_B6003_ = new_B5967_ & new_B6004_;
  assign new_B6002_ = new_B5950_ | new_B5951_;
  assign new_B6001_ = new_B5950_ | new_B5967_;
  assign new_B6000_ = ~new_B5967_ & ~new_B6003_;
  assign new_B5999_ = new_B5967_ | new_B6004_;
  assign new_B5998_ = new_B5950_ & ~new_B5951_;
  assign new_B5997_ = ~new_B5950_ & new_B5951_;
  assign new_B5996_ = new_B5960_ | new_B5993_;
  assign new_B5995_ = ~new_B5960_ & ~new_B5994_;
  assign new_B5994_ = new_B5960_ & new_B5993_;
  assign new_B5993_ = ~new_B5949_ | ~new_B5974_;
  assign new_B5992_ = ~new_B5950_ & new_B5960_;
  assign new_B5991_ = new_B5950_ & ~new_B5960_;
  assign new_B5990_ = new_B5952_ & new_B5989_;
  assign new_B5989_ = new_B6008_ | new_B6007_;
  assign new_B5988_ = ~new_B5952_ & new_B5987_;
  assign new_B5987_ = new_B6010_ | new_B6009_;
  assign new_B5986_ = new_B5952_ | new_B5985_;
  assign new_B5985_ = new_B6006_ | new_B6005_;
  assign new_B5984_ = ~new_B5964_ & ~new_B5974_;
  assign new_B5983_ = new_B5964_ & new_B5974_;
  assign new_B5982_ = ~new_B5964_ | new_B5974_;
  assign new_B5981_ = new_B5948_ & ~new_B5949_;
  assign new_B5980_ = ~new_B5948_ & new_B5949_;
  assign new_B5979_ = new_B6001_ & ~new_B6002_;
  assign new_B5978_ = ~new_B6001_ & new_B6002_;
  assign new_B5977_ = ~new_B6000_ | ~new_B5999_;
  assign new_B5976_ = new_B5992_ | new_B5991_;
  assign new_B5975_ = new_B5998_ | new_B5997_;
  assign new_B5974_ = new_B5988_ | new_B5990_;
  assign new_B5973_ = ~new_B5995_ | ~new_B5996_;
  assign new_B5972_ = new_B5948_ & ~new_B5949_;
  assign new_B5971_ = new_B5962_ & ~new_B5974_;
  assign new_B5970_ = ~new_B5962_ & new_B5974_;
  assign new_B5969_ = ~new_B5960_ & new_B5986_;
  assign new_B5968_ = new_B5984_ | new_B5983_;
  assign new_B5967_ = new_B5981_ | new_B5980_;
  assign new_B5966_ = new_B5949_ | new_B5982_;
  assign new_B5965_ = new_B5974_ & new_B5977_;
  assign new_B5964_ = new_B5979_ | new_B5978_;
  assign new_B5963_ = new_B5974_ & new_B5973_;
  assign new_B5962_ = new_B5976_ & new_B5975_;
  assign new_B5961_ = new_B5971_ | new_B5970_;
  assign new_B5960_ = new_B5949_ | new_B5972_;
  assign B5959 = new_B5960_ | new_B5969_;
  assign B5958 = new_B5967_ & new_B5968_;
  assign B5957 = new_B5967_ & new_B5966_;
  assign B5956 = new_B5965_ | new_B5964_;
  assign B5955 = new_B5963_ | new_B5962_;
  assign B5954 = new_B5961_ & new_B5960_;
  assign new_B5953_ = new_C6879_;
  assign new_B5952_ = new_C6812_;
  assign new_B5951_ = new_C6745_;
  assign new_B5950_ = new_C6678_;
  assign new_B5949_ = new_C6611_;
  assign new_B5948_ = new_C6544_;
  assign new_B5947_ = ~new_B5886_ & new_B5900_;
  assign new_B5946_ = new_B5886_ & ~new_B5900_;
  assign new_B5945_ = new_B5886_ & ~new_B5900_;
  assign new_B5944_ = ~new_B5886_ & ~new_B5900_;
  assign new_B5943_ = new_B5886_ & new_B5900_;
  assign new_B5942_ = new_B5946_ | new_B5947_;
  assign new_B5941_ = ~new_B5886_ & new_B5900_;
  assign new_B5940_ = new_B5944_ | new_B5945_;
  assign new_B5939_ = ~new_B5915_ & ~new_B5935_;
  assign new_B5938_ = new_B5915_ & new_B5935_;
  assign new_B5937_ = ~new_B5882_ | ~new_B5907_;
  assign new_B5936_ = new_B5900_ & new_B5937_;
  assign new_B5935_ = new_B5883_ | new_B5884_;
  assign new_B5934_ = new_B5883_ | new_B5900_;
  assign new_B5933_ = ~new_B5900_ & ~new_B5936_;
  assign new_B5932_ = new_B5900_ | new_B5937_;
  assign new_B5931_ = new_B5883_ & ~new_B5884_;
  assign new_B5930_ = ~new_B5883_ & new_B5884_;
  assign new_B5929_ = new_B5893_ | new_B5926_;
  assign new_B5928_ = ~new_B5893_ & ~new_B5927_;
  assign new_B5927_ = new_B5893_ & new_B5926_;
  assign new_B5926_ = ~new_B5882_ | ~new_B5907_;
  assign new_B5925_ = ~new_B5883_ & new_B5893_;
  assign new_B5924_ = new_B5883_ & ~new_B5893_;
  assign new_B5923_ = new_B5885_ & new_B5922_;
  assign new_B5922_ = new_B5941_ | new_B5940_;
  assign new_B5921_ = ~new_B5885_ & new_B5920_;
  assign new_B5920_ = new_B5943_ | new_B5942_;
  assign new_B5919_ = new_B5885_ | new_B5918_;
  assign new_B5918_ = new_B5939_ | new_B5938_;
  assign new_B5917_ = ~new_B5897_ & ~new_B5907_;
  assign new_B5916_ = new_B5897_ & new_B5907_;
  assign new_B5915_ = ~new_B5897_ | new_B5907_;
  assign new_B5914_ = new_B5881_ & ~new_B5882_;
  assign new_B5913_ = ~new_B5881_ & new_B5882_;
  assign new_B5912_ = new_B5934_ & ~new_B5935_;
  assign new_B5911_ = ~new_B5934_ & new_B5935_;
  assign new_B5910_ = ~new_B5933_ | ~new_B5932_;
  assign new_B5909_ = new_B5925_ | new_B5924_;
  assign new_B5908_ = new_B5931_ | new_B5930_;
  assign new_B5907_ = new_B5921_ | new_B5923_;
  assign new_B5906_ = ~new_B5928_ | ~new_B5929_;
  assign new_B5905_ = new_B5881_ & ~new_B5882_;
  assign new_B5904_ = new_B5895_ & ~new_B5907_;
  assign new_B5903_ = ~new_B5895_ & new_B5907_;
  assign new_B5902_ = ~new_B5893_ & new_B5919_;
  assign new_B5901_ = new_B5917_ | new_B5916_;
  assign new_B5900_ = new_B5914_ | new_B5913_;
  assign new_B5899_ = new_B5882_ | new_B5915_;
  assign new_B5898_ = new_B5907_ & new_B5910_;
  assign new_B5897_ = new_B5912_ | new_B5911_;
  assign new_B5896_ = new_B5907_ & new_B5906_;
  assign new_B5895_ = new_B5909_ & new_B5908_;
  assign new_B5894_ = new_B5904_ | new_B5903_;
  assign new_B5893_ = new_B5882_ | new_B5905_;
  assign B5892 = new_B5893_ | new_B5902_;
  assign B5891 = new_B5900_ & new_B5901_;
  assign B5890 = new_B5900_ & new_B5899_;
  assign B5889 = new_B5898_ | new_B5897_;
  assign B5888 = new_B5896_ | new_B5895_;
  assign B5887 = new_B5894_ & new_B5893_;
  assign new_B5886_ = new_C6477_;
  assign new_B5885_ = new_C6410_;
  assign new_B5884_ = new_C6343_;
  assign new_B5883_ = new_C6276_;
  assign new_B5882_ = new_C6209_;
  assign new_B5881_ = new_C6142_;
  assign new_B5880_ = ~new_B5819_ & new_B5833_;
  assign new_B5879_ = new_B5819_ & ~new_B5833_;
  assign new_B5878_ = new_B5819_ & ~new_B5833_;
  assign new_B5877_ = ~new_B5819_ & ~new_B5833_;
  assign new_B5876_ = new_B5819_ & new_B5833_;
  assign new_B5875_ = new_B5879_ | new_B5880_;
  assign new_B5874_ = ~new_B5819_ & new_B5833_;
  assign new_B5873_ = new_B5877_ | new_B5878_;
  assign new_B5872_ = ~new_B5848_ & ~new_B5868_;
  assign new_B5871_ = new_B5848_ & new_B5868_;
  assign new_B5870_ = ~new_B5815_ | ~new_B5840_;
  assign new_B5869_ = new_B5833_ & new_B5870_;
  assign new_B5868_ = new_B5816_ | new_B5817_;
  assign new_B5867_ = new_B5816_ | new_B5833_;
  assign new_B5866_ = ~new_B5833_ & ~new_B5869_;
  assign new_B5865_ = new_B5833_ | new_B5870_;
  assign new_B5864_ = new_B5816_ & ~new_B5817_;
  assign new_B5863_ = ~new_B5816_ & new_B5817_;
  assign new_B5862_ = new_B5826_ | new_B5859_;
  assign new_B5861_ = ~new_B5826_ & ~new_B5860_;
  assign new_B5860_ = new_B5826_ & new_B5859_;
  assign new_B5859_ = ~new_B5815_ | ~new_B5840_;
  assign new_B5858_ = ~new_B5816_ & new_B5826_;
  assign new_B5857_ = new_B5816_ & ~new_B5826_;
  assign new_B5856_ = new_B5818_ & new_B5855_;
  assign new_B5855_ = new_B5874_ | new_B5873_;
  assign new_B5854_ = ~new_B5818_ & new_B5853_;
  assign new_B5853_ = new_B5876_ | new_B5875_;
  assign new_B5852_ = new_B5818_ | new_B5851_;
  assign new_B5851_ = new_B5872_ | new_B5871_;
  assign new_B5850_ = ~new_B5830_ & ~new_B5840_;
  assign new_B5849_ = new_B5830_ & new_B5840_;
  assign new_B5848_ = ~new_B5830_ | new_B5840_;
  assign new_B5847_ = new_B5814_ & ~new_B5815_;
  assign new_B5846_ = ~new_B5814_ & new_B5815_;
  assign new_B5845_ = new_B5867_ & ~new_B5868_;
  assign new_B5844_ = ~new_B5867_ & new_B5868_;
  assign new_B5843_ = ~new_B5866_ | ~new_B5865_;
  assign new_B5842_ = new_B5858_ | new_B5857_;
  assign new_B5841_ = new_B5864_ | new_B5863_;
  assign new_B5840_ = new_B5854_ | new_B5856_;
  assign new_B5839_ = ~new_B5861_ | ~new_B5862_;
  assign new_B5838_ = new_B5814_ & ~new_B5815_;
  assign new_B5837_ = new_B5828_ & ~new_B5840_;
  assign new_B5836_ = ~new_B5828_ & new_B5840_;
  assign new_B5835_ = ~new_B5826_ & new_B5852_;
  assign new_B5834_ = new_B5850_ | new_B5849_;
  assign new_B5833_ = new_B5847_ | new_B5846_;
  assign new_B5832_ = new_B5815_ | new_B5848_;
  assign new_B5831_ = new_B5840_ & new_B5843_;
  assign new_B5830_ = new_B5845_ | new_B5844_;
  assign new_B5829_ = new_B5840_ & new_B5839_;
  assign new_B5828_ = new_B5842_ & new_B5841_;
  assign new_B5827_ = new_B5837_ | new_B5836_;
  assign new_B5826_ = new_B5815_ | new_B5838_;
  assign B5825 = new_B5826_ | new_B5835_;
  assign B5824 = new_B5833_ & new_B5834_;
  assign B5823 = new_B5833_ & new_B5832_;
  assign B5822 = new_B5831_ | new_B5830_;
  assign B5821 = new_B5829_ | new_B5828_;
  assign B5820 = new_B5827_ & new_B5826_;
  assign new_B5819_ = new_C6075_;
  assign new_B5818_ = new_C6008_;
  assign new_B5817_ = new_C5941_;
  assign new_B5816_ = new_C5874_;
  assign new_B5815_ = new_C5807_;
  assign new_B5814_ = new_C5740_;
  assign new_B5813_ = ~new_B5752_ & new_B5766_;
  assign new_B5812_ = new_B5752_ & ~new_B5766_;
  assign new_B5811_ = new_B5752_ & ~new_B5766_;
  assign new_B5810_ = ~new_B5752_ & ~new_B5766_;
  assign new_B5809_ = new_B5752_ & new_B5766_;
  assign new_B5808_ = new_B5812_ | new_B5813_;
  assign new_B5807_ = ~new_B5752_ & new_B5766_;
  assign new_B5806_ = new_B5810_ | new_B5811_;
  assign new_B5805_ = ~new_B5781_ & ~new_B5801_;
  assign new_B5804_ = new_B5781_ & new_B5801_;
  assign new_B5803_ = ~new_B5748_ | ~new_B5773_;
  assign new_B5802_ = new_B5766_ & new_B5803_;
  assign new_B5801_ = new_B5749_ | new_B5750_;
  assign new_B5800_ = new_B5749_ | new_B5766_;
  assign new_B5799_ = ~new_B5766_ & ~new_B5802_;
  assign new_B5798_ = new_B5766_ | new_B5803_;
  assign new_B5797_ = new_B5749_ & ~new_B5750_;
  assign new_B5796_ = ~new_B5749_ & new_B5750_;
  assign new_B5795_ = new_B5759_ | new_B5792_;
  assign new_B5794_ = ~new_B5759_ & ~new_B5793_;
  assign new_B5793_ = new_B5759_ & new_B5792_;
  assign new_B5792_ = ~new_B5748_ | ~new_B5773_;
  assign new_B5791_ = ~new_B5749_ & new_B5759_;
  assign new_B5790_ = new_B5749_ & ~new_B5759_;
  assign new_B5789_ = new_B5751_ & new_B5788_;
  assign new_B5788_ = new_B5807_ | new_B5806_;
  assign new_B5787_ = ~new_B5751_ & new_B5786_;
  assign new_B5786_ = new_B5809_ | new_B5808_;
  assign new_B5785_ = new_B5751_ | new_B5784_;
  assign new_B5784_ = new_B5805_ | new_B5804_;
  assign new_B5783_ = ~new_B5763_ & ~new_B5773_;
  assign new_B5782_ = new_B5763_ & new_B5773_;
  assign new_B5781_ = ~new_B5763_ | new_B5773_;
  assign new_B5780_ = new_B5747_ & ~new_B5748_;
  assign new_B5779_ = ~new_B5747_ & new_B5748_;
  assign new_B5778_ = new_B5800_ & ~new_B5801_;
  assign new_B5777_ = ~new_B5800_ & new_B5801_;
  assign new_B5776_ = ~new_B5799_ | ~new_B5798_;
  assign new_B5775_ = new_B5791_ | new_B5790_;
  assign new_B5774_ = new_B5797_ | new_B5796_;
  assign new_B5773_ = new_B5787_ | new_B5789_;
  assign new_B5772_ = ~new_B5794_ | ~new_B5795_;
  assign new_B5771_ = new_B5747_ & ~new_B5748_;
  assign new_B5770_ = new_B5761_ & ~new_B5773_;
  assign new_B5769_ = ~new_B5761_ & new_B5773_;
  assign new_B5768_ = ~new_B5759_ & new_B5785_;
  assign new_B5767_ = new_B5783_ | new_B5782_;
  assign new_B5766_ = new_B5780_ | new_B5779_;
  assign new_B5765_ = new_B5748_ | new_B5781_;
  assign new_B5764_ = new_B5773_ & new_B5776_;
  assign new_B5763_ = new_B5778_ | new_B5777_;
  assign new_B5762_ = new_B5773_ & new_B5772_;
  assign new_B5761_ = new_B5775_ & new_B5774_;
  assign new_B5760_ = new_B5770_ | new_B5769_;
  assign new_B5759_ = new_B5748_ | new_B5771_;
  assign B5758 = new_B5759_ | new_B5768_;
  assign B5757 = new_B5766_ & new_B5767_;
  assign B5756 = new_B5766_ & new_B5765_;
  assign B5755 = new_B5764_ | new_B5763_;
  assign B5754 = new_B5762_ | new_B5761_;
  assign B5753 = new_B5760_ & new_B5759_;
  assign new_B5752_ = new_C5673_;
  assign new_B5751_ = new_C5606_;
  assign new_B5750_ = new_C5539_;
  assign new_B5749_ = new_C5472_;
  assign new_B5748_ = new_C5405_;
  assign new_B5747_ = new_C5338_;
  assign new_B5746_ = ~new_B5685_ & new_B5699_;
  assign new_B5745_ = new_B5685_ & ~new_B5699_;
  assign new_B5744_ = new_B5685_ & ~new_B5699_;
  assign new_B5743_ = ~new_B5685_ & ~new_B5699_;
  assign new_B5742_ = new_B5685_ & new_B5699_;
  assign new_B5741_ = new_B5745_ | new_B5746_;
  assign new_B5740_ = ~new_B5685_ & new_B5699_;
  assign new_B5739_ = new_B5743_ | new_B5744_;
  assign new_B5738_ = ~new_B5714_ & ~new_B5734_;
  assign new_B5737_ = new_B5714_ & new_B5734_;
  assign new_B5736_ = ~new_B5681_ | ~new_B5706_;
  assign new_B5735_ = new_B5699_ & new_B5736_;
  assign new_B5734_ = new_B5682_ | new_B5683_;
  assign new_B5733_ = new_B5682_ | new_B5699_;
  assign new_B5732_ = ~new_B5699_ & ~new_B5735_;
  assign new_B5731_ = new_B5699_ | new_B5736_;
  assign new_B5730_ = new_B5682_ & ~new_B5683_;
  assign new_B5729_ = ~new_B5682_ & new_B5683_;
  assign new_B5728_ = new_B5692_ | new_B5725_;
  assign new_B5727_ = ~new_B5692_ & ~new_B5726_;
  assign new_B5726_ = new_B5692_ & new_B5725_;
  assign new_B5725_ = ~new_B5681_ | ~new_B5706_;
  assign new_B5724_ = ~new_B5682_ & new_B5692_;
  assign new_B5723_ = new_B5682_ & ~new_B5692_;
  assign new_B5722_ = new_B5684_ & new_B5721_;
  assign new_B5721_ = new_B5740_ | new_B5739_;
  assign new_B5720_ = ~new_B5684_ & new_B5719_;
  assign new_B5719_ = new_B5742_ | new_B5741_;
  assign new_B5718_ = new_B5684_ | new_B5717_;
  assign new_B5717_ = new_B5738_ | new_B5737_;
  assign new_B5716_ = ~new_B5696_ & ~new_B5706_;
  assign new_B5715_ = new_B5696_ & new_B5706_;
  assign new_B5714_ = ~new_B5696_ | new_B5706_;
  assign new_B5713_ = new_B5680_ & ~new_B5681_;
  assign new_B5712_ = ~new_B5680_ & new_B5681_;
  assign new_B5711_ = new_B5733_ & ~new_B5734_;
  assign new_B5710_ = ~new_B5733_ & new_B5734_;
  assign new_B5709_ = ~new_B5732_ | ~new_B5731_;
  assign new_B5708_ = new_B5724_ | new_B5723_;
  assign new_B5707_ = new_B5730_ | new_B5729_;
  assign new_B5706_ = new_B5720_ | new_B5722_;
  assign new_B5705_ = ~new_B5727_ | ~new_B5728_;
  assign new_B5704_ = new_B5680_ & ~new_B5681_;
  assign new_B5703_ = new_B5694_ & ~new_B5706_;
  assign new_B5702_ = ~new_B5694_ & new_B5706_;
  assign new_B5701_ = ~new_B5692_ & new_B5718_;
  assign new_B5700_ = new_B5716_ | new_B5715_;
  assign new_B5699_ = new_B5713_ | new_B5712_;
  assign new_B5698_ = new_B5681_ | new_B5714_;
  assign new_B5697_ = new_B5706_ & new_B5709_;
  assign new_B5696_ = new_B5711_ | new_B5710_;
  assign new_B5695_ = new_B5706_ & new_B5705_;
  assign new_B5694_ = new_B5708_ & new_B5707_;
  assign new_B5693_ = new_B5703_ | new_B5702_;
  assign new_B5692_ = new_B5681_ | new_B5704_;
  assign B5691 = new_B5692_ | new_B5701_;
  assign B5690 = new_B5699_ & new_B5700_;
  assign B5689 = new_B5699_ & new_B5698_;
  assign B5688 = new_B5697_ | new_B5696_;
  assign B5687 = new_B5695_ | new_B5694_;
  assign B5686 = new_B5693_ & new_B5692_;
  assign new_B5685_ = new_C5271_;
  assign new_B5684_ = new_C5204_;
  assign new_B5683_ = new_C5137_;
  assign new_B5682_ = new_C5070_;
  assign new_B5681_ = new_C5003_;
  assign new_B5680_ = new_C4936_;
  assign new_B5679_ = ~new_B5618_ & new_B5632_;
  assign new_B5678_ = new_B5618_ & ~new_B5632_;
  assign new_B5677_ = new_B5618_ & ~new_B5632_;
  assign new_B5676_ = ~new_B5618_ & ~new_B5632_;
  assign new_B5675_ = new_B5618_ & new_B5632_;
  assign new_B5674_ = new_B5678_ | new_B5679_;
  assign new_B5673_ = ~new_B5618_ & new_B5632_;
  assign new_B5672_ = new_B5676_ | new_B5677_;
  assign new_B5671_ = ~new_B5647_ & ~new_B5667_;
  assign new_B5670_ = new_B5647_ & new_B5667_;
  assign new_B5669_ = ~new_B5614_ | ~new_B5639_;
  assign new_B5668_ = new_B5632_ & new_B5669_;
  assign new_B5667_ = new_B5615_ | new_B5616_;
  assign new_B5666_ = new_B5615_ | new_B5632_;
  assign new_B5665_ = ~new_B5632_ & ~new_B5668_;
  assign new_B5664_ = new_B5632_ | new_B5669_;
  assign new_B5663_ = new_B5615_ & ~new_B5616_;
  assign new_B5662_ = ~new_B5615_ & new_B5616_;
  assign new_B5661_ = new_B5625_ | new_B5658_;
  assign new_B5660_ = ~new_B5625_ & ~new_B5659_;
  assign new_B5659_ = new_B5625_ & new_B5658_;
  assign new_B5658_ = ~new_B5614_ | ~new_B5639_;
  assign new_B5657_ = ~new_B5615_ & new_B5625_;
  assign new_B5656_ = new_B5615_ & ~new_B5625_;
  assign new_B5655_ = new_B5617_ & new_B5654_;
  assign new_B5654_ = new_B5673_ | new_B5672_;
  assign new_B5653_ = ~new_B5617_ & new_B5652_;
  assign new_B5652_ = new_B5675_ | new_B5674_;
  assign new_B5651_ = new_B5617_ | new_B5650_;
  assign new_B5650_ = new_B5671_ | new_B5670_;
  assign new_B5649_ = ~new_B5629_ & ~new_B5639_;
  assign new_B5648_ = new_B5629_ & new_B5639_;
  assign new_B5647_ = ~new_B5629_ | new_B5639_;
  assign new_B5646_ = new_B5613_ & ~new_B5614_;
  assign new_B5645_ = ~new_B5613_ & new_B5614_;
  assign new_B5644_ = new_B5666_ & ~new_B5667_;
  assign new_B5643_ = ~new_B5666_ & new_B5667_;
  assign new_B5642_ = ~new_B5665_ | ~new_B5664_;
  assign new_B5641_ = new_B5657_ | new_B5656_;
  assign new_B5640_ = new_B5663_ | new_B5662_;
  assign new_B5639_ = new_B5653_ | new_B5655_;
  assign new_B5638_ = ~new_B5660_ | ~new_B5661_;
  assign new_B5637_ = new_B5613_ & ~new_B5614_;
  assign new_B5636_ = new_B5627_ & ~new_B5639_;
  assign new_B5635_ = ~new_B5627_ & new_B5639_;
  assign new_B5634_ = ~new_B5625_ & new_B5651_;
  assign new_B5633_ = new_B5649_ | new_B5648_;
  assign new_B5632_ = new_B5646_ | new_B5645_;
  assign new_B5631_ = new_B5614_ | new_B5647_;
  assign new_B5630_ = new_B5639_ & new_B5642_;
  assign new_B5629_ = new_B5644_ | new_B5643_;
  assign new_B5628_ = new_B5639_ & new_B5638_;
  assign new_B5627_ = new_B5641_ & new_B5640_;
  assign new_B5626_ = new_B5636_ | new_B5635_;
  assign new_B5625_ = new_B5614_ | new_B5637_;
  assign B5624 = new_B5625_ | new_B5634_;
  assign B5623 = new_B5632_ & new_B5633_;
  assign B5622 = new_B5632_ & new_B5631_;
  assign B5621 = new_B5630_ | new_B5629_;
  assign B5620 = new_B5628_ | new_B5627_;
  assign B5619 = new_B5626_ & new_B5625_;
  assign new_B5618_ = new_C4869_;
  assign new_B5617_ = new_C4802_;
  assign new_B5616_ = new_C4735_;
  assign new_B5615_ = new_C4668_;
  assign new_B5614_ = new_C4601_;
  assign new_B5613_ = new_C4534_;
  assign new_B5612_ = ~new_B5551_ & new_B5565_;
  assign new_B5611_ = new_B5551_ & ~new_B5565_;
  assign new_B5610_ = new_B5551_ & ~new_B5565_;
  assign new_B5609_ = ~new_B5551_ & ~new_B5565_;
  assign new_B5608_ = new_B5551_ & new_B5565_;
  assign new_B5607_ = new_B5611_ | new_B5612_;
  assign new_B5606_ = ~new_B5551_ & new_B5565_;
  assign new_B5605_ = new_B5609_ | new_B5610_;
  assign new_B5604_ = ~new_B5580_ & ~new_B5600_;
  assign new_B5603_ = new_B5580_ & new_B5600_;
  assign new_B5602_ = ~new_B5547_ | ~new_B5572_;
  assign new_B5601_ = new_B5565_ & new_B5602_;
  assign new_B5600_ = new_B5548_ | new_B5549_;
  assign new_B5599_ = new_B5548_ | new_B5565_;
  assign new_B5598_ = ~new_B5565_ & ~new_B5601_;
  assign new_B5597_ = new_B5565_ | new_B5602_;
  assign new_B5596_ = new_B5548_ & ~new_B5549_;
  assign new_B5595_ = ~new_B5548_ & new_B5549_;
  assign new_B5594_ = new_B5558_ | new_B5591_;
  assign new_B5593_ = ~new_B5558_ & ~new_B5592_;
  assign new_B5592_ = new_B5558_ & new_B5591_;
  assign new_B5591_ = ~new_B5547_ | ~new_B5572_;
  assign new_B5590_ = ~new_B5548_ & new_B5558_;
  assign new_B5589_ = new_B5548_ & ~new_B5558_;
  assign new_B5588_ = new_B5550_ & new_B5587_;
  assign new_B5587_ = new_B5606_ | new_B5605_;
  assign new_B5586_ = ~new_B5550_ & new_B5585_;
  assign new_B5585_ = new_B5608_ | new_B5607_;
  assign new_B5584_ = new_B5550_ | new_B5583_;
  assign new_B5583_ = new_B5604_ | new_B5603_;
  assign new_B5582_ = ~new_B5562_ & ~new_B5572_;
  assign new_B5581_ = new_B5562_ & new_B5572_;
  assign new_B5580_ = ~new_B5562_ | new_B5572_;
  assign new_B5579_ = new_B5546_ & ~new_B5547_;
  assign new_B5578_ = ~new_B5546_ & new_B5547_;
  assign new_B5577_ = new_B5599_ & ~new_B5600_;
  assign new_B5576_ = ~new_B5599_ & new_B5600_;
  assign new_B5575_ = ~new_B5598_ | ~new_B5597_;
  assign new_B5574_ = new_B5590_ | new_B5589_;
  assign new_B5573_ = new_B5596_ | new_B5595_;
  assign new_B5572_ = new_B5586_ | new_B5588_;
  assign new_B5571_ = ~new_B5593_ | ~new_B5594_;
  assign new_B5570_ = new_B5546_ & ~new_B5547_;
  assign new_B5569_ = new_B5560_ & ~new_B5572_;
  assign new_B5568_ = ~new_B5560_ & new_B5572_;
  assign new_B5567_ = ~new_B5558_ & new_B5584_;
  assign new_B5566_ = new_B5582_ | new_B5581_;
  assign new_B5565_ = new_B5579_ | new_B5578_;
  assign new_B5564_ = new_B5547_ | new_B5580_;
  assign new_B5563_ = new_B5572_ & new_B5575_;
  assign new_B5562_ = new_B5577_ | new_B5576_;
  assign new_B5561_ = new_B5572_ & new_B5571_;
  assign new_B5560_ = new_B5574_ & new_B5573_;
  assign new_B5559_ = new_B5569_ | new_B5568_;
  assign new_B5558_ = new_B5547_ | new_B5570_;
  assign B5557 = new_B5558_ | new_B5567_;
  assign B5556 = new_B5565_ & new_B5566_;
  assign B5555 = new_B5565_ & new_B5564_;
  assign B5554 = new_B5563_ | new_B5562_;
  assign B5553 = new_B5561_ | new_B5560_;
  assign B5552 = new_B5559_ & new_B5558_;
  assign new_B5551_ = new_C4467_;
  assign new_B5550_ = new_C4400_;
  assign new_B5549_ = new_C4333_;
  assign new_B5548_ = new_C4266_;
  assign new_B5547_ = new_C4199_;
  assign new_B5546_ = new_C4132_;
  assign new_B5545_ = ~new_B5484_ & new_B5498_;
  assign new_B5544_ = new_B5484_ & ~new_B5498_;
  assign new_B5543_ = new_B5484_ & ~new_B5498_;
  assign new_B5542_ = ~new_B5484_ & ~new_B5498_;
  assign new_B5541_ = new_B5484_ & new_B5498_;
  assign new_B5540_ = new_B5544_ | new_B5545_;
  assign new_B5539_ = ~new_B5484_ & new_B5498_;
  assign new_B5538_ = new_B5542_ | new_B5543_;
  assign new_B5537_ = ~new_B5513_ & ~new_B5533_;
  assign new_B5536_ = new_B5513_ & new_B5533_;
  assign new_B5535_ = ~new_B5480_ | ~new_B5505_;
  assign new_B5534_ = new_B5498_ & new_B5535_;
  assign new_B5533_ = new_B5481_ | new_B5482_;
  assign new_B5532_ = new_B5481_ | new_B5498_;
  assign new_B5531_ = ~new_B5498_ & ~new_B5534_;
  assign new_B5530_ = new_B5498_ | new_B5535_;
  assign new_B5529_ = new_B5481_ & ~new_B5482_;
  assign new_B5528_ = ~new_B5481_ & new_B5482_;
  assign new_B5527_ = new_B5491_ | new_B5524_;
  assign new_B5526_ = ~new_B5491_ & ~new_B5525_;
  assign new_B5525_ = new_B5491_ & new_B5524_;
  assign new_B5524_ = ~new_B5480_ | ~new_B5505_;
  assign new_B5523_ = ~new_B5481_ & new_B5491_;
  assign new_B5522_ = new_B5481_ & ~new_B5491_;
  assign new_B5521_ = new_B5483_ & new_B5520_;
  assign new_B5520_ = new_B5539_ | new_B5538_;
  assign new_B5519_ = ~new_B5483_ & new_B5518_;
  assign new_B5518_ = new_B5541_ | new_B5540_;
  assign new_B5517_ = new_B5483_ | new_B5516_;
  assign new_B5516_ = new_B5537_ | new_B5536_;
  assign new_B5515_ = ~new_B5495_ & ~new_B5505_;
  assign new_B5514_ = new_B5495_ & new_B5505_;
  assign new_B5513_ = ~new_B5495_ | new_B5505_;
  assign new_B5512_ = new_B5479_ & ~new_B5480_;
  assign new_B5511_ = ~new_B5479_ & new_B5480_;
  assign new_B5510_ = new_B5532_ & ~new_B5533_;
  assign new_B5509_ = ~new_B5532_ & new_B5533_;
  assign new_B5508_ = ~new_B5531_ | ~new_B5530_;
  assign new_B5507_ = new_B5523_ | new_B5522_;
  assign new_B5506_ = new_B5529_ | new_B5528_;
  assign new_B5505_ = new_B5519_ | new_B5521_;
  assign new_B5504_ = ~new_B5526_ | ~new_B5527_;
  assign new_B5503_ = new_B5479_ & ~new_B5480_;
  assign new_B5502_ = new_B5493_ & ~new_B5505_;
  assign new_B5501_ = ~new_B5493_ & new_B5505_;
  assign new_B5500_ = ~new_B5491_ & new_B5517_;
  assign new_B5499_ = new_B5515_ | new_B5514_;
  assign new_B5498_ = new_B5512_ | new_B5511_;
  assign new_B5497_ = new_B5480_ | new_B5513_;
  assign new_B5496_ = new_B5505_ & new_B5508_;
  assign new_B5495_ = new_B5510_ | new_B5509_;
  assign new_B5494_ = new_B5505_ & new_B5504_;
  assign new_B5493_ = new_B5507_ & new_B5506_;
  assign new_B5492_ = new_B5502_ | new_B5501_;
  assign new_B5491_ = new_B5480_ | new_B5503_;
  assign B5490 = new_B5491_ | new_B5500_;
  assign B5489 = new_B5498_ & new_B5499_;
  assign B5488 = new_B5498_ & new_B5497_;
  assign B5487 = new_B5496_ | new_B5495_;
  assign B5486 = new_B5494_ | new_B5493_;
  assign B5485 = new_B5492_ & new_B5491_;
  assign new_B5484_ = new_C4065_;
  assign new_B5483_ = new_C3998_;
  assign new_B5482_ = new_C3931_;
  assign new_B5481_ = new_C3864_;
  assign new_B5480_ = new_C3797_;
  assign new_B5479_ = new_C3730_;
  assign new_B5478_ = ~new_B5417_ & new_B5431_;
  assign new_B5477_ = new_B5417_ & ~new_B5431_;
  assign new_B5476_ = new_B5417_ & ~new_B5431_;
  assign new_B5475_ = ~new_B5417_ & ~new_B5431_;
  assign new_B5474_ = new_B5417_ & new_B5431_;
  assign new_B5473_ = new_B5477_ | new_B5478_;
  assign new_B5472_ = ~new_B5417_ & new_B5431_;
  assign new_B5471_ = new_B5475_ | new_B5476_;
  assign new_B5470_ = ~new_B5446_ & ~new_B5466_;
  assign new_B5469_ = new_B5446_ & new_B5466_;
  assign new_B5468_ = ~new_B5413_ | ~new_B5438_;
  assign new_B5467_ = new_B5431_ & new_B5468_;
  assign new_B5466_ = new_B5414_ | new_B5415_;
  assign new_B5465_ = new_B5414_ | new_B5431_;
  assign new_B5464_ = ~new_B5431_ & ~new_B5467_;
  assign new_B5463_ = new_B5431_ | new_B5468_;
  assign new_B5462_ = new_B5414_ & ~new_B5415_;
  assign new_B5461_ = ~new_B5414_ & new_B5415_;
  assign new_B5460_ = new_B5424_ | new_B5457_;
  assign new_B5459_ = ~new_B5424_ & ~new_B5458_;
  assign new_B5458_ = new_B5424_ & new_B5457_;
  assign new_B5457_ = ~new_B5413_ | ~new_B5438_;
  assign new_B5456_ = ~new_B5414_ & new_B5424_;
  assign new_B5455_ = new_B5414_ & ~new_B5424_;
  assign new_B5454_ = new_B5416_ & new_B5453_;
  assign new_B5453_ = new_B5472_ | new_B5471_;
  assign new_B5452_ = ~new_B5416_ & new_B5451_;
  assign new_B5451_ = new_B5474_ | new_B5473_;
  assign new_B5450_ = new_B5416_ | new_B5449_;
  assign new_B5449_ = new_B5470_ | new_B5469_;
  assign new_B5448_ = ~new_B5428_ & ~new_B5438_;
  assign new_B5447_ = new_B5428_ & new_B5438_;
  assign new_B5446_ = ~new_B5428_ | new_B5438_;
  assign new_B5445_ = new_B5412_ & ~new_B5413_;
  assign new_B5444_ = ~new_B5412_ & new_B5413_;
  assign new_B5443_ = new_B5465_ & ~new_B5466_;
  assign new_B5442_ = ~new_B5465_ & new_B5466_;
  assign new_B5441_ = ~new_B5464_ | ~new_B5463_;
  assign new_B5440_ = new_B5456_ | new_B5455_;
  assign new_B5439_ = new_B5462_ | new_B5461_;
  assign new_B5438_ = new_B5452_ | new_B5454_;
  assign new_B5437_ = ~new_B5459_ | ~new_B5460_;
  assign new_B5436_ = new_B5412_ & ~new_B5413_;
  assign new_B5435_ = new_B5426_ & ~new_B5438_;
  assign new_B5434_ = ~new_B5426_ & new_B5438_;
  assign new_B5433_ = ~new_B5424_ & new_B5450_;
  assign new_B5432_ = new_B5448_ | new_B5447_;
  assign new_B5431_ = new_B5445_ | new_B5444_;
  assign new_B5430_ = new_B5413_ | new_B5446_;
  assign new_B5429_ = new_B5438_ & new_B5441_;
  assign new_B5428_ = new_B5443_ | new_B5442_;
  assign new_B5427_ = new_B5438_ & new_B5437_;
  assign new_B5426_ = new_B5440_ & new_B5439_;
  assign new_B5425_ = new_B5435_ | new_B5434_;
  assign new_B5424_ = new_B5413_ | new_B5436_;
  assign B5423 = new_B5424_ | new_B5433_;
  assign B5422 = new_B5431_ & new_B5432_;
  assign B5421 = new_B5431_ & new_B5430_;
  assign B5420 = new_B5429_ | new_B5428_;
  assign B5419 = new_B5427_ | new_B5426_;
  assign B5418 = new_B5425_ & new_B5424_;
  assign new_B5417_ = new_C3663_;
  assign new_B5416_ = new_C3596_;
  assign new_B5415_ = new_C3529_;
  assign new_B5414_ = new_C3462_;
  assign new_B5413_ = new_C3395_;
  assign new_B5412_ = new_C3328_;
  assign new_B5411_ = ~new_B5350_ & new_B5364_;
  assign new_B5410_ = new_B5350_ & ~new_B5364_;
  assign new_B5409_ = new_B5350_ & ~new_B5364_;
  assign new_B5408_ = ~new_B5350_ & ~new_B5364_;
  assign new_B5407_ = new_B5350_ & new_B5364_;
  assign new_B5406_ = new_B5410_ | new_B5411_;
  assign new_B5405_ = ~new_B5350_ & new_B5364_;
  assign new_B5404_ = new_B5408_ | new_B5409_;
  assign new_B5403_ = ~new_B5379_ & ~new_B5399_;
  assign new_B5402_ = new_B5379_ & new_B5399_;
  assign new_B5401_ = ~new_B5346_ | ~new_B5371_;
  assign new_B5400_ = new_B5364_ & new_B5401_;
  assign new_B5399_ = new_B5347_ | new_B5348_;
  assign new_B5398_ = new_B5347_ | new_B5364_;
  assign new_B5397_ = ~new_B5364_ & ~new_B5400_;
  assign new_B5396_ = new_B5364_ | new_B5401_;
  assign new_B5395_ = new_B5347_ & ~new_B5348_;
  assign new_B5394_ = ~new_B5347_ & new_B5348_;
  assign new_B5393_ = new_B5357_ | new_B5390_;
  assign new_B5392_ = ~new_B5357_ & ~new_B5391_;
  assign new_B5391_ = new_B5357_ & new_B5390_;
  assign new_B5390_ = ~new_B5346_ | ~new_B5371_;
  assign new_B5389_ = ~new_B5347_ & new_B5357_;
  assign new_B5388_ = new_B5347_ & ~new_B5357_;
  assign new_B5387_ = new_B5349_ & new_B5386_;
  assign new_B5386_ = new_B5405_ | new_B5404_;
  assign new_B5385_ = ~new_B5349_ & new_B5384_;
  assign new_B5384_ = new_B5407_ | new_B5406_;
  assign new_B5383_ = new_B5349_ | new_B5382_;
  assign new_B5382_ = new_B5403_ | new_B5402_;
  assign new_B5381_ = ~new_B5361_ & ~new_B5371_;
  assign new_B5380_ = new_B5361_ & new_B5371_;
  assign new_B5379_ = ~new_B5361_ | new_B5371_;
  assign new_B5378_ = new_B5345_ & ~new_B5346_;
  assign new_B5377_ = ~new_B5345_ & new_B5346_;
  assign new_B5376_ = new_B5398_ & ~new_B5399_;
  assign new_B5375_ = ~new_B5398_ & new_B5399_;
  assign new_B5374_ = ~new_B5397_ | ~new_B5396_;
  assign new_B5373_ = new_B5389_ | new_B5388_;
  assign new_B5372_ = new_B5395_ | new_B5394_;
  assign new_B5371_ = new_B5385_ | new_B5387_;
  assign new_B5370_ = ~new_B5392_ | ~new_B5393_;
  assign new_B5369_ = new_B5345_ & ~new_B5346_;
  assign new_B5368_ = new_B5359_ & ~new_B5371_;
  assign new_B5367_ = ~new_B5359_ & new_B5371_;
  assign new_B5366_ = ~new_B5357_ & new_B5383_;
  assign new_B5365_ = new_B5381_ | new_B5380_;
  assign new_B5364_ = new_B5378_ | new_B5377_;
  assign new_B5363_ = new_B5346_ | new_B5379_;
  assign new_B5362_ = new_B5371_ & new_B5374_;
  assign new_B5361_ = new_B5376_ | new_B5375_;
  assign new_B5360_ = new_B5371_ & new_B5370_;
  assign new_B5359_ = new_B5373_ & new_B5372_;
  assign new_B5358_ = new_B5368_ | new_B5367_;
  assign new_B5357_ = new_B5346_ | new_B5369_;
  assign B5356 = new_B5357_ | new_B5366_;
  assign B5355 = new_B5364_ & new_B5365_;
  assign B5354 = new_B5364_ & new_B5363_;
  assign B5353 = new_B5362_ | new_B5361_;
  assign B5352 = new_B5360_ | new_B5359_;
  assign B5351 = new_B5358_ & new_B5357_;
  assign new_B5350_ = new_C3261_;
  assign new_B5349_ = new_C3194_;
  assign new_B5348_ = new_C3127_;
  assign new_B5347_ = new_C3060_;
  assign new_B5346_ = new_C2993_;
  assign new_B5345_ = new_C2926_;
  assign new_B5344_ = ~new_B5283_ & new_B5297_;
  assign new_B5343_ = new_B5283_ & ~new_B5297_;
  assign new_B5342_ = new_B5283_ & ~new_B5297_;
  assign new_B5341_ = ~new_B5283_ & ~new_B5297_;
  assign new_B5340_ = new_B5283_ & new_B5297_;
  assign new_B5339_ = new_B5343_ | new_B5344_;
  assign new_B5338_ = ~new_B5283_ & new_B5297_;
  assign new_B5337_ = new_B5341_ | new_B5342_;
  assign new_B5336_ = ~new_B5312_ & ~new_B5332_;
  assign new_B5335_ = new_B5312_ & new_B5332_;
  assign new_B5334_ = ~new_B5279_ | ~new_B5304_;
  assign new_B5333_ = new_B5297_ & new_B5334_;
  assign new_B5332_ = new_B5280_ | new_B5281_;
  assign new_B5331_ = new_B5280_ | new_B5297_;
  assign new_B5330_ = ~new_B5297_ & ~new_B5333_;
  assign new_B5329_ = new_B5297_ | new_B5334_;
  assign new_B5328_ = new_B5280_ & ~new_B5281_;
  assign new_B5327_ = ~new_B5280_ & new_B5281_;
  assign new_B5326_ = new_B5290_ | new_B5323_;
  assign new_B5325_ = ~new_B5290_ & ~new_B5324_;
  assign new_B5324_ = new_B5290_ & new_B5323_;
  assign new_B5323_ = ~new_B5279_ | ~new_B5304_;
  assign new_B5322_ = ~new_B5280_ & new_B5290_;
  assign new_B5321_ = new_B5280_ & ~new_B5290_;
  assign new_B5320_ = new_B5282_ & new_B5319_;
  assign new_B5319_ = new_B5338_ | new_B5337_;
  assign new_B5318_ = ~new_B5282_ & new_B5317_;
  assign new_B5317_ = new_B5340_ | new_B5339_;
  assign new_B5316_ = new_B5282_ | new_B5315_;
  assign new_B5315_ = new_B5336_ | new_B5335_;
  assign new_B5314_ = ~new_B5294_ & ~new_B5304_;
  assign new_B5313_ = new_B5294_ & new_B5304_;
  assign new_B5312_ = ~new_B5294_ | new_B5304_;
  assign new_B5311_ = new_B5278_ & ~new_B5279_;
  assign new_B5310_ = ~new_B5278_ & new_B5279_;
  assign new_B5309_ = new_B5331_ & ~new_B5332_;
  assign new_B5308_ = ~new_B5331_ & new_B5332_;
  assign new_B5307_ = ~new_B5330_ | ~new_B5329_;
  assign new_B5306_ = new_B5322_ | new_B5321_;
  assign new_B5305_ = new_B5328_ | new_B5327_;
  assign new_B5304_ = new_B5318_ | new_B5320_;
  assign new_B5303_ = ~new_B5325_ | ~new_B5326_;
  assign new_B5302_ = new_B5278_ & ~new_B5279_;
  assign new_B5301_ = new_B5292_ & ~new_B5304_;
  assign new_B5300_ = ~new_B5292_ & new_B5304_;
  assign new_B5299_ = ~new_B5290_ & new_B5316_;
  assign new_B5298_ = new_B5314_ | new_B5313_;
  assign new_B5297_ = new_B5311_ | new_B5310_;
  assign new_B5296_ = new_B5279_ | new_B5312_;
  assign new_B5295_ = new_B5304_ & new_B5307_;
  assign new_B5294_ = new_B5309_ | new_B5308_;
  assign new_B5293_ = new_B5304_ & new_B5303_;
  assign new_B5292_ = new_B5306_ & new_B5305_;
  assign new_B5291_ = new_B5301_ | new_B5300_;
  assign new_B5290_ = new_B5279_ | new_B5302_;
  assign B5289 = new_B5290_ | new_B5299_;
  assign B5288 = new_B5297_ & new_B5298_;
  assign B5287 = new_B5297_ & new_B5296_;
  assign B5286 = new_B5295_ | new_B5294_;
  assign B5285 = new_B5293_ | new_B5292_;
  assign B5284 = new_B5291_ & new_B5290_;
  assign new_B5283_ = new_C2859_;
  assign new_B5282_ = new_C2792_;
  assign new_B5281_ = new_C2725_;
  assign new_B5280_ = new_C2658_;
  assign new_B5279_ = new_C2591_;
  assign new_B5278_ = new_C2523_;
  assign new_B5277_ = ~new_B5216_ & new_B5230_;
  assign new_B5276_ = new_B5216_ & ~new_B5230_;
  assign new_B5275_ = new_B5216_ & ~new_B5230_;
  assign new_B5274_ = ~new_B5216_ & ~new_B5230_;
  assign new_B5273_ = new_B5216_ & new_B5230_;
  assign new_B5272_ = new_B5276_ | new_B5277_;
  assign new_B5271_ = ~new_B5216_ & new_B5230_;
  assign new_B5270_ = new_B5274_ | new_B5275_;
  assign new_B5269_ = ~new_B5245_ & ~new_B5265_;
  assign new_B5268_ = new_B5245_ & new_B5265_;
  assign new_B5267_ = ~new_B5212_ | ~new_B5237_;
  assign new_B5266_ = new_B5230_ & new_B5267_;
  assign new_B5265_ = new_B5213_ | new_B5214_;
  assign new_B5264_ = new_B5213_ | new_B5230_;
  assign new_B5263_ = ~new_B5230_ & ~new_B5266_;
  assign new_B5262_ = new_B5230_ | new_B5267_;
  assign new_B5261_ = new_B5213_ & ~new_B5214_;
  assign new_B5260_ = ~new_B5213_ & new_B5214_;
  assign new_B5259_ = new_B5223_ | new_B5256_;
  assign new_B5258_ = ~new_B5223_ & ~new_B5257_;
  assign new_B5257_ = new_B5223_ & new_B5256_;
  assign new_B5256_ = ~new_B5212_ | ~new_B5237_;
  assign new_B5255_ = ~new_B5213_ & new_B5223_;
  assign new_B5254_ = new_B5213_ & ~new_B5223_;
  assign new_B5253_ = new_B5215_ & new_B5252_;
  assign new_B5252_ = new_B5271_ | new_B5270_;
  assign new_B5251_ = ~new_B5215_ & new_B5250_;
  assign new_B5250_ = new_B5273_ | new_B5272_;
  assign new_B5249_ = new_B5215_ | new_B5248_;
  assign new_B5248_ = new_B5269_ | new_B5268_;
  assign new_B5247_ = ~new_B5227_ & ~new_B5237_;
  assign new_B5246_ = new_B5227_ & new_B5237_;
  assign new_B5245_ = ~new_B5227_ | new_B5237_;
  assign new_B5244_ = new_B5211_ & ~new_B5212_;
  assign new_B5243_ = ~new_B5211_ & new_B5212_;
  assign new_B5242_ = new_B5264_ & ~new_B5265_;
  assign new_B5241_ = ~new_B5264_ & new_B5265_;
  assign new_B5240_ = ~new_B5263_ | ~new_B5262_;
  assign new_B5239_ = new_B5255_ | new_B5254_;
  assign new_B5238_ = new_B5261_ | new_B5260_;
  assign new_B5237_ = new_B5251_ | new_B5253_;
  assign new_B5236_ = ~new_B5258_ | ~new_B5259_;
  assign new_B5235_ = new_B5211_ & ~new_B5212_;
  assign new_B5234_ = new_B5225_ & ~new_B5237_;
  assign new_B5233_ = ~new_B5225_ & new_B5237_;
  assign new_B5232_ = ~new_B5223_ & new_B5249_;
  assign new_B5231_ = new_B5247_ | new_B5246_;
  assign new_B5230_ = new_B5244_ | new_B5243_;
  assign new_B5229_ = new_B5212_ | new_B5245_;
  assign new_B5228_ = new_B5237_ & new_B5240_;
  assign new_B5227_ = new_B5242_ | new_B5241_;
  assign new_B5226_ = new_B5237_ & new_B5236_;
  assign new_B5225_ = new_B5239_ & new_B5238_;
  assign new_B5224_ = new_B5234_ | new_B5233_;
  assign new_B5223_ = new_B5212_ | new_B5235_;
  assign B5222 = new_B5223_ | new_B5232_;
  assign B5221 = new_B5230_ & new_B5231_;
  assign B5220 = new_B5230_ & new_B5229_;
  assign B5219 = new_B5228_ | new_B5227_;
  assign B5218 = new_B5226_ | new_B5225_;
  assign B5217 = new_B5224_ & new_B5223_;
  assign new_B5216_ = new_D6929_;
  assign new_B5215_ = new_D6862_;
  assign new_B5214_ = new_D6795_;
  assign new_B5213_ = new_D6728_;
  assign new_B5212_ = new_D6661_;
  assign new_B5211_ = new_D6594_;
  assign new_B5210_ = ~new_B5149_ & new_B5163_;
  assign new_B5209_ = new_B5149_ & ~new_B5163_;
  assign new_B5208_ = new_B5149_ & ~new_B5163_;
  assign new_B5207_ = ~new_B5149_ & ~new_B5163_;
  assign new_B5206_ = new_B5149_ & new_B5163_;
  assign new_B5205_ = new_B5209_ | new_B5210_;
  assign new_B5204_ = ~new_B5149_ & new_B5163_;
  assign new_B5203_ = new_B5207_ | new_B5208_;
  assign new_B5202_ = ~new_B5178_ & ~new_B5198_;
  assign new_B5201_ = new_B5178_ & new_B5198_;
  assign new_B5200_ = ~new_B5145_ | ~new_B5170_;
  assign new_B5199_ = new_B5163_ & new_B5200_;
  assign new_B5198_ = new_B5146_ | new_B5147_;
  assign new_B5197_ = new_B5146_ | new_B5163_;
  assign new_B5196_ = ~new_B5163_ & ~new_B5199_;
  assign new_B5195_ = new_B5163_ | new_B5200_;
  assign new_B5194_ = new_B5146_ & ~new_B5147_;
  assign new_B5193_ = ~new_B5146_ & new_B5147_;
  assign new_B5192_ = new_B5156_ | new_B5189_;
  assign new_B5191_ = ~new_B5156_ & ~new_B5190_;
  assign new_B5190_ = new_B5156_ & new_B5189_;
  assign new_B5189_ = ~new_B5145_ | ~new_B5170_;
  assign new_B5188_ = ~new_B5146_ & new_B5156_;
  assign new_B5187_ = new_B5146_ & ~new_B5156_;
  assign new_B5186_ = new_B5148_ & new_B5185_;
  assign new_B5185_ = new_B5204_ | new_B5203_;
  assign new_B5184_ = ~new_B5148_ & new_B5183_;
  assign new_B5183_ = new_B5206_ | new_B5205_;
  assign new_B5182_ = new_B5148_ | new_B5181_;
  assign new_B5181_ = new_B5202_ | new_B5201_;
  assign new_B5180_ = ~new_B5160_ & ~new_B5170_;
  assign new_B5179_ = new_B5160_ & new_B5170_;
  assign new_B5178_ = ~new_B5160_ | new_B5170_;
  assign new_B5177_ = new_B5144_ & ~new_B5145_;
  assign new_B5176_ = ~new_B5144_ & new_B5145_;
  assign new_B5175_ = new_B5197_ & ~new_B5198_;
  assign new_B5174_ = ~new_B5197_ & new_B5198_;
  assign new_B5173_ = ~new_B5196_ | ~new_B5195_;
  assign new_B5172_ = new_B5188_ | new_B5187_;
  assign new_B5171_ = new_B5194_ | new_B5193_;
  assign new_B5170_ = new_B5184_ | new_B5186_;
  assign new_B5169_ = ~new_B5191_ | ~new_B5192_;
  assign new_B5168_ = new_B5144_ & ~new_B5145_;
  assign new_B5167_ = new_B5158_ & ~new_B5170_;
  assign new_B5166_ = ~new_B5158_ & new_B5170_;
  assign new_B5165_ = ~new_B5156_ & new_B5182_;
  assign new_B5164_ = new_B5180_ | new_B5179_;
  assign new_B5163_ = new_B5177_ | new_B5176_;
  assign new_B5162_ = new_B5145_ | new_B5178_;
  assign new_B5161_ = new_B5170_ & new_B5173_;
  assign new_B5160_ = new_B5175_ | new_B5174_;
  assign new_B5159_ = new_B5170_ & new_B5169_;
  assign new_B5158_ = new_B5172_ & new_B5171_;
  assign new_B5157_ = new_B5167_ | new_B5166_;
  assign new_B5156_ = new_B5145_ | new_B5168_;
  assign B5155 = new_B5156_ | new_B5165_;
  assign B5154 = new_B5163_ & new_B5164_;
  assign B5153 = new_B5163_ & new_B5162_;
  assign B5152 = new_B5161_ | new_B5160_;
  assign B5151 = new_B5159_ | new_B5158_;
  assign B5150 = new_B5157_ & new_B5156_;
  assign new_B5149_ = new_D6527_;
  assign new_B5148_ = new_D6460_;
  assign new_B5147_ = new_D6393_;
  assign new_B5146_ = new_D6326_;
  assign new_B5145_ = new_D6259_;
  assign new_B5144_ = new_D6192_;
  assign new_B5143_ = ~new_B5082_ & new_B5096_;
  assign new_B5142_ = new_B5082_ & ~new_B5096_;
  assign new_B5141_ = new_B5082_ & ~new_B5096_;
  assign new_B5140_ = ~new_B5082_ & ~new_B5096_;
  assign new_B5139_ = new_B5082_ & new_B5096_;
  assign new_B5138_ = new_B5142_ | new_B5143_;
  assign new_B5137_ = ~new_B5082_ & new_B5096_;
  assign new_B5136_ = new_B5140_ | new_B5141_;
  assign new_B5135_ = ~new_B5111_ & ~new_B5131_;
  assign new_B5134_ = new_B5111_ & new_B5131_;
  assign new_B5133_ = ~new_B5078_ | ~new_B5103_;
  assign new_B5132_ = new_B5096_ & new_B5133_;
  assign new_B5131_ = new_B5079_ | new_B5080_;
  assign new_B5130_ = new_B5079_ | new_B5096_;
  assign new_B5129_ = ~new_B5096_ & ~new_B5132_;
  assign new_B5128_ = new_B5096_ | new_B5133_;
  assign new_B5127_ = new_B5079_ & ~new_B5080_;
  assign new_B5126_ = ~new_B5079_ & new_B5080_;
  assign new_B5125_ = new_B5089_ | new_B5122_;
  assign new_B5124_ = ~new_B5089_ & ~new_B5123_;
  assign new_B5123_ = new_B5089_ & new_B5122_;
  assign new_B5122_ = ~new_B5078_ | ~new_B5103_;
  assign new_B5121_ = ~new_B5079_ & new_B5089_;
  assign new_B5120_ = new_B5079_ & ~new_B5089_;
  assign new_B5119_ = new_B5081_ & new_B5118_;
  assign new_B5118_ = new_B5137_ | new_B5136_;
  assign new_B5117_ = ~new_B5081_ & new_B5116_;
  assign new_B5116_ = new_B5139_ | new_B5138_;
  assign new_B5115_ = new_B5081_ | new_B5114_;
  assign new_B5114_ = new_B5135_ | new_B5134_;
  assign new_B5113_ = ~new_B5093_ & ~new_B5103_;
  assign new_B5112_ = new_B5093_ & new_B5103_;
  assign new_B5111_ = ~new_B5093_ | new_B5103_;
  assign new_B5110_ = new_B5077_ & ~new_B5078_;
  assign new_B5109_ = ~new_B5077_ & new_B5078_;
  assign new_B5108_ = new_B5130_ & ~new_B5131_;
  assign new_B5107_ = ~new_B5130_ & new_B5131_;
  assign new_B5106_ = ~new_B5129_ | ~new_B5128_;
  assign new_B5105_ = new_B5121_ | new_B5120_;
  assign new_B5104_ = new_B5127_ | new_B5126_;
  assign new_B5103_ = new_B5117_ | new_B5119_;
  assign new_B5102_ = ~new_B5124_ | ~new_B5125_;
  assign new_B5101_ = new_B5077_ & ~new_B5078_;
  assign new_B5100_ = new_B5091_ & ~new_B5103_;
  assign new_B5099_ = ~new_B5091_ & new_B5103_;
  assign new_B5098_ = ~new_B5089_ & new_B5115_;
  assign new_B5097_ = new_B5113_ | new_B5112_;
  assign new_B5096_ = new_B5110_ | new_B5109_;
  assign new_B5095_ = new_B5078_ | new_B5111_;
  assign new_B5094_ = new_B5103_ & new_B5106_;
  assign new_B5093_ = new_B5108_ | new_B5107_;
  assign new_B5092_ = new_B5103_ & new_B5102_;
  assign new_B5091_ = new_B5105_ & new_B5104_;
  assign new_B5090_ = new_B5100_ | new_B5099_;
  assign new_B5089_ = new_B5078_ | new_B5101_;
  assign B5088 = new_B5089_ | new_B5098_;
  assign B5087 = new_B5096_ & new_B5097_;
  assign B5086 = new_B5096_ & new_B5095_;
  assign B5085 = new_B5094_ | new_B5093_;
  assign B5084 = new_B5092_ | new_B5091_;
  assign B5083 = new_B5090_ & new_B5089_;
  assign new_B5082_ = new_D6125_;
  assign new_B5081_ = new_D6058_;
  assign new_B5080_ = new_D5991_;
  assign new_B5079_ = new_D5924_;
  assign new_B5078_ = new_D5857_;
  assign new_B5077_ = new_D5790_;
  assign new_B5076_ = ~new_B5015_ & new_B5029_;
  assign new_B5075_ = new_B5015_ & ~new_B5029_;
  assign new_B5074_ = new_B5015_ & ~new_B5029_;
  assign new_B5073_ = ~new_B5015_ & ~new_B5029_;
  assign new_B5072_ = new_B5015_ & new_B5029_;
  assign new_B5071_ = new_B5075_ | new_B5076_;
  assign new_B5070_ = ~new_B5015_ & new_B5029_;
  assign new_B5069_ = new_B5073_ | new_B5074_;
  assign new_B5068_ = ~new_B5044_ & ~new_B5064_;
  assign new_B5067_ = new_B5044_ & new_B5064_;
  assign new_B5066_ = ~new_B5011_ | ~new_B5036_;
  assign new_B5065_ = new_B5029_ & new_B5066_;
  assign new_B5064_ = new_B5012_ | new_B5013_;
  assign new_B5063_ = new_B5012_ | new_B5029_;
  assign new_B5062_ = ~new_B5029_ & ~new_B5065_;
  assign new_B5061_ = new_B5029_ | new_B5066_;
  assign new_B5060_ = new_B5012_ & ~new_B5013_;
  assign new_B5059_ = ~new_B5012_ & new_B5013_;
  assign new_B5058_ = new_B5022_ | new_B5055_;
  assign new_B5057_ = ~new_B5022_ & ~new_B5056_;
  assign new_B5056_ = new_B5022_ & new_B5055_;
  assign new_B5055_ = ~new_B5011_ | ~new_B5036_;
  assign new_B5054_ = ~new_B5012_ & new_B5022_;
  assign new_B5053_ = new_B5012_ & ~new_B5022_;
  assign new_B5052_ = new_B5014_ & new_B5051_;
  assign new_B5051_ = new_B5070_ | new_B5069_;
  assign new_B5050_ = ~new_B5014_ & new_B5049_;
  assign new_B5049_ = new_B5072_ | new_B5071_;
  assign new_B5048_ = new_B5014_ | new_B5047_;
  assign new_B5047_ = new_B5068_ | new_B5067_;
  assign new_B5046_ = ~new_B5026_ & ~new_B5036_;
  assign new_B5045_ = new_B5026_ & new_B5036_;
  assign new_B5044_ = ~new_B5026_ | new_B5036_;
  assign new_B5043_ = new_B5010_ & ~new_B5011_;
  assign new_B5042_ = ~new_B5010_ & new_B5011_;
  assign new_B5041_ = new_B5063_ & ~new_B5064_;
  assign new_B5040_ = ~new_B5063_ & new_B5064_;
  assign new_B5039_ = ~new_B5062_ | ~new_B5061_;
  assign new_B5038_ = new_B5054_ | new_B5053_;
  assign new_B5037_ = new_B5060_ | new_B5059_;
  assign new_B5036_ = new_B5050_ | new_B5052_;
  assign new_B5035_ = ~new_B5057_ | ~new_B5058_;
  assign new_B5034_ = new_B5010_ & ~new_B5011_;
  assign new_B5033_ = new_B5024_ & ~new_B5036_;
  assign new_B5032_ = ~new_B5024_ & new_B5036_;
  assign new_B5031_ = ~new_B5022_ & new_B5048_;
  assign new_B5030_ = new_B5046_ | new_B5045_;
  assign new_B5029_ = new_B5043_ | new_B5042_;
  assign new_B5028_ = new_B5011_ | new_B5044_;
  assign new_B5027_ = new_B5036_ & new_B5039_;
  assign new_B5026_ = new_B5041_ | new_B5040_;
  assign new_B5025_ = new_B5036_ & new_B5035_;
  assign new_B5024_ = new_B5038_ & new_B5037_;
  assign new_B5023_ = new_B5033_ | new_B5032_;
  assign new_B5022_ = new_B5011_ | new_B5034_;
  assign B5021 = new_B5022_ | new_B5031_;
  assign B5020 = new_B5029_ & new_B5030_;
  assign B5019 = new_B5029_ & new_B5028_;
  assign B5018 = new_B5027_ | new_B5026_;
  assign B5017 = new_B5025_ | new_B5024_;
  assign B5016 = new_B5023_ & new_B5022_;
  assign new_B5015_ = new_D5723_;
  assign new_B5014_ = new_D5656_;
  assign new_B5013_ = new_D5589_;
  assign new_B5012_ = new_D5522_;
  assign new_B5011_ = new_D5455_;
  assign new_B5010_ = new_D5388_;
  assign new_B5009_ = ~new_B4948_ & new_B4962_;
  assign new_B5008_ = new_B4948_ & ~new_B4962_;
  assign new_B5007_ = new_B4948_ & ~new_B4962_;
  assign new_B5006_ = ~new_B4948_ & ~new_B4962_;
  assign new_B5005_ = new_B4948_ & new_B4962_;
  assign new_B5004_ = new_B5008_ | new_B5009_;
  assign new_B5003_ = ~new_B4948_ & new_B4962_;
  assign new_B5002_ = new_B5006_ | new_B5007_;
  assign new_B5001_ = ~new_B4977_ & ~new_B4997_;
  assign new_B5000_ = new_B4977_ & new_B4997_;
  assign new_B4999_ = ~new_B4944_ | ~new_B4969_;
  assign new_B4998_ = new_B4962_ & new_B4999_;
  assign new_B4997_ = new_B4945_ | new_B4946_;
  assign new_B4996_ = new_B4945_ | new_B4962_;
  assign new_B4995_ = ~new_B4962_ & ~new_B4998_;
  assign new_B4994_ = new_B4962_ | new_B4999_;
  assign new_B4993_ = new_B4945_ & ~new_B4946_;
  assign new_B4992_ = ~new_B4945_ & new_B4946_;
  assign new_B4991_ = new_B4955_ | new_B4988_;
  assign new_B4990_ = ~new_B4955_ & ~new_B4989_;
  assign new_B4989_ = new_B4955_ & new_B4988_;
  assign new_B4988_ = ~new_B4944_ | ~new_B4969_;
  assign new_B4987_ = ~new_B4945_ & new_B4955_;
  assign new_B4986_ = new_B4945_ & ~new_B4955_;
  assign new_B4985_ = new_B4947_ & new_B4984_;
  assign new_B4984_ = new_B5003_ | new_B5002_;
  assign new_B4983_ = ~new_B4947_ & new_B4982_;
  assign new_B4982_ = new_B5005_ | new_B5004_;
  assign new_B4981_ = new_B4947_ | new_B4980_;
  assign new_B4980_ = new_B5001_ | new_B5000_;
  assign new_B4979_ = ~new_B4959_ & ~new_B4969_;
  assign new_B4978_ = new_B4959_ & new_B4969_;
  assign new_B4977_ = ~new_B4959_ | new_B4969_;
  assign new_B4976_ = new_B4943_ & ~new_B4944_;
  assign new_B4975_ = ~new_B4943_ & new_B4944_;
  assign new_B4974_ = new_B4996_ & ~new_B4997_;
  assign new_B4973_ = ~new_B4996_ & new_B4997_;
  assign new_B4972_ = ~new_B4995_ | ~new_B4994_;
  assign new_B4971_ = new_B4987_ | new_B4986_;
  assign new_B4970_ = new_B4993_ | new_B4992_;
  assign new_B4969_ = new_B4983_ | new_B4985_;
  assign new_B4968_ = ~new_B4990_ | ~new_B4991_;
  assign new_B4967_ = new_B4943_ & ~new_B4944_;
  assign new_B4966_ = new_B4957_ & ~new_B4969_;
  assign new_B4965_ = ~new_B4957_ & new_B4969_;
  assign new_B4964_ = ~new_B4955_ & new_B4981_;
  assign new_B4963_ = new_B4979_ | new_B4978_;
  assign new_B4962_ = new_B4976_ | new_B4975_;
  assign new_B4961_ = new_B4944_ | new_B4977_;
  assign new_B4960_ = new_B4969_ & new_B4972_;
  assign new_B4959_ = new_B4974_ | new_B4973_;
  assign new_B4958_ = new_B4969_ & new_B4968_;
  assign new_B4957_ = new_B4971_ & new_B4970_;
  assign new_B4956_ = new_B4966_ | new_B4965_;
  assign new_B4955_ = new_B4944_ | new_B4967_;
  assign B4954 = new_B4955_ | new_B4964_;
  assign B4953 = new_B4962_ & new_B4963_;
  assign B4952 = new_B4962_ & new_B4961_;
  assign B4951 = new_B4960_ | new_B4959_;
  assign B4950 = new_B4958_ | new_B4957_;
  assign B4949 = new_B4956_ & new_B4955_;
  assign new_B4948_ = new_D5321_;
  assign new_B4947_ = new_D5254_;
  assign new_B4946_ = new_D5187_;
  assign new_B4945_ = new_D5120_;
  assign new_B4944_ = new_D5053_;
  assign new_B4943_ = new_D4986_;
  assign new_B4942_ = ~new_B4881_ & new_B4895_;
  assign new_B4941_ = new_B4881_ & ~new_B4895_;
  assign new_B4940_ = new_B4881_ & ~new_B4895_;
  assign new_B4939_ = ~new_B4881_ & ~new_B4895_;
  assign new_B4938_ = new_B4881_ & new_B4895_;
  assign new_B4937_ = new_B4941_ | new_B4942_;
  assign new_B4936_ = ~new_B4881_ & new_B4895_;
  assign new_B4935_ = new_B4939_ | new_B4940_;
  assign new_B4934_ = ~new_B4910_ & ~new_B4930_;
  assign new_B4933_ = new_B4910_ & new_B4930_;
  assign new_B4932_ = ~new_B4877_ | ~new_B4902_;
  assign new_B4931_ = new_B4895_ & new_B4932_;
  assign new_B4930_ = new_B4878_ | new_B4879_;
  assign new_B4929_ = new_B4878_ | new_B4895_;
  assign new_B4928_ = ~new_B4895_ & ~new_B4931_;
  assign new_B4927_ = new_B4895_ | new_B4932_;
  assign new_B4926_ = new_B4878_ & ~new_B4879_;
  assign new_B4925_ = ~new_B4878_ & new_B4879_;
  assign new_B4924_ = new_B4888_ | new_B4921_;
  assign new_B4923_ = ~new_B4888_ & ~new_B4922_;
  assign new_B4922_ = new_B4888_ & new_B4921_;
  assign new_B4921_ = ~new_B4877_ | ~new_B4902_;
  assign new_B4920_ = ~new_B4878_ & new_B4888_;
  assign new_B4919_ = new_B4878_ & ~new_B4888_;
  assign new_B4918_ = new_B4880_ & new_B4917_;
  assign new_B4917_ = new_B4936_ | new_B4935_;
  assign new_B4916_ = ~new_B4880_ & new_B4915_;
  assign new_B4915_ = new_B4938_ | new_B4937_;
  assign new_B4914_ = new_B4880_ | new_B4913_;
  assign new_B4913_ = new_B4934_ | new_B4933_;
  assign new_B4912_ = ~new_B4892_ & ~new_B4902_;
  assign new_B4911_ = new_B4892_ & new_B4902_;
  assign new_B4910_ = ~new_B4892_ | new_B4902_;
  assign new_B4909_ = new_B4876_ & ~new_B4877_;
  assign new_B4908_ = ~new_B4876_ & new_B4877_;
  assign new_B4907_ = new_B4929_ & ~new_B4930_;
  assign new_B4906_ = ~new_B4929_ & new_B4930_;
  assign new_B4905_ = ~new_B4928_ | ~new_B4927_;
  assign new_B4904_ = new_B4920_ | new_B4919_;
  assign new_B4903_ = new_B4926_ | new_B4925_;
  assign new_B4902_ = new_B4916_ | new_B4918_;
  assign new_B4901_ = ~new_B4923_ | ~new_B4924_;
  assign new_B4900_ = new_B4876_ & ~new_B4877_;
  assign new_B4899_ = new_B4890_ & ~new_B4902_;
  assign new_B4898_ = ~new_B4890_ & new_B4902_;
  assign new_B4897_ = ~new_B4888_ & new_B4914_;
  assign new_B4896_ = new_B4912_ | new_B4911_;
  assign new_B4895_ = new_B4909_ | new_B4908_;
  assign new_B4894_ = new_B4877_ | new_B4910_;
  assign new_B4893_ = new_B4902_ & new_B4905_;
  assign new_B4892_ = new_B4907_ | new_B4906_;
  assign new_B4891_ = new_B4902_ & new_B4901_;
  assign new_B4890_ = new_B4904_ & new_B4903_;
  assign new_B4889_ = new_B4899_ | new_B4898_;
  assign new_B4888_ = new_B4877_ | new_B4900_;
  assign B4887 = new_B4888_ | new_B4897_;
  assign B4886 = new_B4895_ & new_B4896_;
  assign B4885 = new_B4895_ & new_B4894_;
  assign B4884 = new_B4893_ | new_B4892_;
  assign B4883 = new_B4891_ | new_B4890_;
  assign B4882 = new_B4889_ & new_B4888_;
  assign new_B4881_ = new_D4919_;
  assign new_B4880_ = new_D4852_;
  assign new_B4879_ = new_D4785_;
  assign new_B4878_ = new_D4718_;
  assign new_B4877_ = new_D4651_;
  assign new_B4876_ = new_D4584_;
  assign new_B4875_ = ~new_B4814_ & new_B4828_;
  assign new_B4874_ = new_B4814_ & ~new_B4828_;
  assign new_B4873_ = new_B4814_ & ~new_B4828_;
  assign new_B4872_ = ~new_B4814_ & ~new_B4828_;
  assign new_B4871_ = new_B4814_ & new_B4828_;
  assign new_B4870_ = new_B4874_ | new_B4875_;
  assign new_B4869_ = ~new_B4814_ & new_B4828_;
  assign new_B4868_ = new_B4872_ | new_B4873_;
  assign new_B4867_ = ~new_B4843_ & ~new_B4863_;
  assign new_B4866_ = new_B4843_ & new_B4863_;
  assign new_B4865_ = ~new_B4810_ | ~new_B4835_;
  assign new_B4864_ = new_B4828_ & new_B4865_;
  assign new_B4863_ = new_B4811_ | new_B4812_;
  assign new_B4862_ = new_B4811_ | new_B4828_;
  assign new_B4861_ = ~new_B4828_ & ~new_B4864_;
  assign new_B4860_ = new_B4828_ | new_B4865_;
  assign new_B4859_ = new_B4811_ & ~new_B4812_;
  assign new_B4858_ = ~new_B4811_ & new_B4812_;
  assign new_B4857_ = new_B4821_ | new_B4854_;
  assign new_B4856_ = ~new_B4821_ & ~new_B4855_;
  assign new_B4855_ = new_B4821_ & new_B4854_;
  assign new_B4854_ = ~new_B4810_ | ~new_B4835_;
  assign new_B4853_ = ~new_B4811_ & new_B4821_;
  assign new_B4852_ = new_B4811_ & ~new_B4821_;
  assign new_B4851_ = new_B4813_ & new_B4850_;
  assign new_B4850_ = new_B4869_ | new_B4868_;
  assign new_B4849_ = ~new_B4813_ & new_B4848_;
  assign new_B4848_ = new_B4871_ | new_B4870_;
  assign new_B4847_ = new_B4813_ | new_B4846_;
  assign new_B4846_ = new_B4867_ | new_B4866_;
  assign new_B4845_ = ~new_B4825_ & ~new_B4835_;
  assign new_B4844_ = new_B4825_ & new_B4835_;
  assign new_B4843_ = ~new_B4825_ | new_B4835_;
  assign new_B4842_ = new_B4809_ & ~new_B4810_;
  assign new_B4841_ = ~new_B4809_ & new_B4810_;
  assign new_B4840_ = new_B4862_ & ~new_B4863_;
  assign new_B4839_ = ~new_B4862_ & new_B4863_;
  assign new_B4838_ = ~new_B4861_ | ~new_B4860_;
  assign new_B4837_ = new_B4853_ | new_B4852_;
  assign new_B4836_ = new_B4859_ | new_B4858_;
  assign new_B4835_ = new_B4849_ | new_B4851_;
  assign new_B4834_ = ~new_B4856_ | ~new_B4857_;
  assign new_B4833_ = new_B4809_ & ~new_B4810_;
  assign new_B4832_ = new_B4823_ & ~new_B4835_;
  assign new_B4831_ = ~new_B4823_ & new_B4835_;
  assign new_B4830_ = ~new_B4821_ & new_B4847_;
  assign new_B4829_ = new_B4845_ | new_B4844_;
  assign new_B4828_ = new_B4842_ | new_B4841_;
  assign new_B4827_ = new_B4810_ | new_B4843_;
  assign new_B4826_ = new_B4835_ & new_B4838_;
  assign new_B4825_ = new_B4840_ | new_B4839_;
  assign new_B4824_ = new_B4835_ & new_B4834_;
  assign new_B4823_ = new_B4837_ & new_B4836_;
  assign new_B4822_ = new_B4832_ | new_B4831_;
  assign new_B4821_ = new_B4810_ | new_B4833_;
  assign B4820 = new_B4821_ | new_B4830_;
  assign B4819 = new_B4828_ & new_B4829_;
  assign B4818 = new_B4828_ & new_B4827_;
  assign B4817 = new_B4826_ | new_B4825_;
  assign B4816 = new_B4824_ | new_B4823_;
  assign B4815 = new_B4822_ & new_B4821_;
  assign new_B4814_ = new_D4517_;
  assign new_B4813_ = new_D4450_;
  assign new_B4812_ = new_D4383_;
  assign new_B4811_ = new_D4316_;
  assign new_B4810_ = new_D4249_;
  assign new_B4809_ = new_D4182_;
  assign new_B4808_ = ~new_B4747_ & new_B4761_;
  assign new_B4807_ = new_B4747_ & ~new_B4761_;
  assign new_B4806_ = new_B4747_ & ~new_B4761_;
  assign new_B4805_ = ~new_B4747_ & ~new_B4761_;
  assign new_B4804_ = new_B4747_ & new_B4761_;
  assign new_B4803_ = new_B4807_ | new_B4808_;
  assign new_B4802_ = ~new_B4747_ & new_B4761_;
  assign new_B4801_ = new_B4805_ | new_B4806_;
  assign new_B4800_ = ~new_B4776_ & ~new_B4796_;
  assign new_B4799_ = new_B4776_ & new_B4796_;
  assign new_B4798_ = ~new_B4743_ | ~new_B4768_;
  assign new_B4797_ = new_B4761_ & new_B4798_;
  assign new_B4796_ = new_B4744_ | new_B4745_;
  assign new_B4795_ = new_B4744_ | new_B4761_;
  assign new_B4794_ = ~new_B4761_ & ~new_B4797_;
  assign new_B4793_ = new_B4761_ | new_B4798_;
  assign new_B4792_ = new_B4744_ & ~new_B4745_;
  assign new_B4791_ = ~new_B4744_ & new_B4745_;
  assign new_B4790_ = new_B4754_ | new_B4787_;
  assign new_B4789_ = ~new_B4754_ & ~new_B4788_;
  assign new_B4788_ = new_B4754_ & new_B4787_;
  assign new_B4787_ = ~new_B4743_ | ~new_B4768_;
  assign new_B4786_ = ~new_B4744_ & new_B4754_;
  assign new_B4785_ = new_B4744_ & ~new_B4754_;
  assign new_B4784_ = new_B4746_ & new_B4783_;
  assign new_B4783_ = new_B4802_ | new_B4801_;
  assign new_B4782_ = ~new_B4746_ & new_B4781_;
  assign new_B4781_ = new_B4804_ | new_B4803_;
  assign new_B4780_ = new_B4746_ | new_B4779_;
  assign new_B4779_ = new_B4800_ | new_B4799_;
  assign new_B4778_ = ~new_B4758_ & ~new_B4768_;
  assign new_B4777_ = new_B4758_ & new_B4768_;
  assign new_B4776_ = ~new_B4758_ | new_B4768_;
  assign new_B4775_ = new_B4742_ & ~new_B4743_;
  assign new_B4774_ = ~new_B4742_ & new_B4743_;
  assign new_B4773_ = new_B4795_ & ~new_B4796_;
  assign new_B4772_ = ~new_B4795_ & new_B4796_;
  assign new_B4771_ = ~new_B4794_ | ~new_B4793_;
  assign new_B4770_ = new_B4786_ | new_B4785_;
  assign new_B4769_ = new_B4792_ | new_B4791_;
  assign new_B4768_ = new_B4782_ | new_B4784_;
  assign new_B4767_ = ~new_B4789_ | ~new_B4790_;
  assign new_B4766_ = new_B4742_ & ~new_B4743_;
  assign new_B4765_ = new_B4756_ & ~new_B4768_;
  assign new_B4764_ = ~new_B4756_ & new_B4768_;
  assign new_B4763_ = ~new_B4754_ & new_B4780_;
  assign new_B4762_ = new_B4778_ | new_B4777_;
  assign new_B4761_ = new_B4775_ | new_B4774_;
  assign new_B4760_ = new_B4743_ | new_B4776_;
  assign new_B4759_ = new_B4768_ & new_B4771_;
  assign new_B4758_ = new_B4773_ | new_B4772_;
  assign new_B4757_ = new_B4768_ & new_B4767_;
  assign new_B4756_ = new_B4770_ & new_B4769_;
  assign new_B4755_ = new_B4765_ | new_B4764_;
  assign new_B4754_ = new_B4743_ | new_B4766_;
  assign B4753 = new_B4754_ | new_B4763_;
  assign B4752 = new_B4761_ & new_B4762_;
  assign B4751 = new_B4761_ & new_B4760_;
  assign B4750 = new_B4759_ | new_B4758_;
  assign B4749 = new_B4757_ | new_B4756_;
  assign B4748 = new_B4755_ & new_B4754_;
  assign new_B4747_ = new_D4115_;
  assign new_B4746_ = new_D4048_;
  assign new_B4745_ = new_D3981_;
  assign new_B4744_ = new_D3914_;
  assign new_B4743_ = new_D3847_;
  assign new_B4742_ = new_D3780_;
  assign new_B4741_ = ~new_B4680_ & new_B4694_;
  assign new_B4740_ = new_B4680_ & ~new_B4694_;
  assign new_B4739_ = new_B4680_ & ~new_B4694_;
  assign new_B4738_ = ~new_B4680_ & ~new_B4694_;
  assign new_B4737_ = new_B4680_ & new_B4694_;
  assign new_B4736_ = new_B4740_ | new_B4741_;
  assign new_B4735_ = ~new_B4680_ & new_B4694_;
  assign new_B4734_ = new_B4738_ | new_B4739_;
  assign new_B4733_ = ~new_B4709_ & ~new_B4729_;
  assign new_B4732_ = new_B4709_ & new_B4729_;
  assign new_B4731_ = ~new_B4676_ | ~new_B4701_;
  assign new_B4730_ = new_B4694_ & new_B4731_;
  assign new_B4729_ = new_B4677_ | new_B4678_;
  assign new_B4728_ = new_B4677_ | new_B4694_;
  assign new_B4727_ = ~new_B4694_ & ~new_B4730_;
  assign new_B4726_ = new_B4694_ | new_B4731_;
  assign new_B4725_ = new_B4677_ & ~new_B4678_;
  assign new_B4724_ = ~new_B4677_ & new_B4678_;
  assign new_B4723_ = new_B4687_ | new_B4720_;
  assign new_B4722_ = ~new_B4687_ & ~new_B4721_;
  assign new_B4721_ = new_B4687_ & new_B4720_;
  assign new_B4720_ = ~new_B4676_ | ~new_B4701_;
  assign new_B4719_ = ~new_B4677_ & new_B4687_;
  assign new_B4718_ = new_B4677_ & ~new_B4687_;
  assign new_B4717_ = new_B4679_ & new_B4716_;
  assign new_B4716_ = new_B4735_ | new_B4734_;
  assign new_B4715_ = ~new_B4679_ & new_B4714_;
  assign new_B4714_ = new_B4737_ | new_B4736_;
  assign new_B4713_ = new_B4679_ | new_B4712_;
  assign new_B4712_ = new_B4733_ | new_B4732_;
  assign new_B4711_ = ~new_B4691_ & ~new_B4701_;
  assign new_B4710_ = new_B4691_ & new_B4701_;
  assign new_B4709_ = ~new_B4691_ | new_B4701_;
  assign new_B4708_ = new_B4675_ & ~new_B4676_;
  assign new_B4707_ = ~new_B4675_ & new_B4676_;
  assign new_B4706_ = new_B4728_ & ~new_B4729_;
  assign new_B4705_ = ~new_B4728_ & new_B4729_;
  assign new_B4704_ = ~new_B4727_ | ~new_B4726_;
  assign new_B4703_ = new_B4719_ | new_B4718_;
  assign new_B4702_ = new_B4725_ | new_B4724_;
  assign new_B4701_ = new_B4715_ | new_B4717_;
  assign new_B4700_ = ~new_B4722_ | ~new_B4723_;
  assign new_B4699_ = new_B4675_ & ~new_B4676_;
  assign new_B4698_ = new_B4689_ & ~new_B4701_;
  assign new_B4697_ = ~new_B4689_ & new_B4701_;
  assign new_B4696_ = ~new_B4687_ & new_B4713_;
  assign new_B4695_ = new_B4711_ | new_B4710_;
  assign new_B4694_ = new_B4708_ | new_B4707_;
  assign new_B4693_ = new_B4676_ | new_B4709_;
  assign new_B4692_ = new_B4701_ & new_B4704_;
  assign new_B4691_ = new_B4706_ | new_B4705_;
  assign new_B4690_ = new_B4701_ & new_B4700_;
  assign new_B4689_ = new_B4703_ & new_B4702_;
  assign new_B4688_ = new_B4698_ | new_B4697_;
  assign new_B4687_ = new_B4676_ | new_B4699_;
  assign B4686 = new_B4687_ | new_B4696_;
  assign B4685 = new_B4694_ & new_B4695_;
  assign B4684 = new_B4694_ & new_B4693_;
  assign B4683 = new_B4692_ | new_B4691_;
  assign B4682 = new_B4690_ | new_B4689_;
  assign B4681 = new_B4688_ & new_B4687_;
  assign new_B4680_ = new_D3713_;
  assign new_B4679_ = new_D3646_;
  assign new_B4678_ = new_D3579_;
  assign new_B4677_ = new_D3512_;
  assign new_B4676_ = new_D3445_;
  assign new_B4675_ = new_D3378_;
  assign new_B4674_ = ~new_B4613_ & new_B4627_;
  assign new_B4673_ = new_B4613_ & ~new_B4627_;
  assign new_B4672_ = new_B4613_ & ~new_B4627_;
  assign new_B4671_ = ~new_B4613_ & ~new_B4627_;
  assign new_B4670_ = new_B4613_ & new_B4627_;
  assign new_B4669_ = new_B4673_ | new_B4674_;
  assign new_B4668_ = ~new_B4613_ & new_B4627_;
  assign new_B4667_ = new_B4671_ | new_B4672_;
  assign new_B4666_ = ~new_B4642_ & ~new_B4662_;
  assign new_B4665_ = new_B4642_ & new_B4662_;
  assign new_B4664_ = ~new_B4609_ | ~new_B4634_;
  assign new_B4663_ = new_B4627_ & new_B4664_;
  assign new_B4662_ = new_B4610_ | new_B4611_;
  assign new_B4661_ = new_B4610_ | new_B4627_;
  assign new_B4660_ = ~new_B4627_ & ~new_B4663_;
  assign new_B4659_ = new_B4627_ | new_B4664_;
  assign new_B4658_ = new_B4610_ & ~new_B4611_;
  assign new_B4657_ = ~new_B4610_ & new_B4611_;
  assign new_B4656_ = new_B4620_ | new_B4653_;
  assign new_B4655_ = ~new_B4620_ & ~new_B4654_;
  assign new_B4654_ = new_B4620_ & new_B4653_;
  assign new_B4653_ = ~new_B4609_ | ~new_B4634_;
  assign new_B4652_ = ~new_B4610_ & new_B4620_;
  assign new_B4651_ = new_B4610_ & ~new_B4620_;
  assign new_B4650_ = new_B4612_ & new_B4649_;
  assign new_B4649_ = new_B4668_ | new_B4667_;
  assign new_B4648_ = ~new_B4612_ & new_B4647_;
  assign new_B4647_ = new_B4670_ | new_B4669_;
  assign new_B4646_ = new_B4612_ | new_B4645_;
  assign new_B4645_ = new_B4666_ | new_B4665_;
  assign new_B4644_ = ~new_B4624_ & ~new_B4634_;
  assign new_B4643_ = new_B4624_ & new_B4634_;
  assign new_B4642_ = ~new_B4624_ | new_B4634_;
  assign new_B4641_ = new_B4608_ & ~new_B4609_;
  assign new_B4640_ = ~new_B4608_ & new_B4609_;
  assign new_B4639_ = new_B4661_ & ~new_B4662_;
  assign new_B4638_ = ~new_B4661_ & new_B4662_;
  assign new_B4637_ = ~new_B4660_ | ~new_B4659_;
  assign new_B4636_ = new_B4652_ | new_B4651_;
  assign new_B4635_ = new_B4658_ | new_B4657_;
  assign new_B4634_ = new_B4648_ | new_B4650_;
  assign new_B4633_ = ~new_B4655_ | ~new_B4656_;
  assign new_B4632_ = new_B4608_ & ~new_B4609_;
  assign new_B4631_ = new_B4622_ & ~new_B4634_;
  assign new_B4630_ = ~new_B4622_ & new_B4634_;
  assign new_B4629_ = ~new_B4620_ & new_B4646_;
  assign new_B4628_ = new_B4644_ | new_B4643_;
  assign new_B4627_ = new_B4641_ | new_B4640_;
  assign new_B4626_ = new_B4609_ | new_B4642_;
  assign new_B4625_ = new_B4634_ & new_B4637_;
  assign new_B4624_ = new_B4639_ | new_B4638_;
  assign new_B4623_ = new_B4634_ & new_B4633_;
  assign new_B4622_ = new_B4636_ & new_B4635_;
  assign new_B4621_ = new_B4631_ | new_B4630_;
  assign new_B4620_ = new_B4609_ | new_B4632_;
  assign B4619 = new_B4620_ | new_B4629_;
  assign B4618 = new_B4627_ & new_B4628_;
  assign B4617 = new_B4627_ & new_B4626_;
  assign B4616 = new_B4625_ | new_B4624_;
  assign B4615 = new_B4623_ | new_B4622_;
  assign B4614 = new_B4621_ & new_B4620_;
  assign new_B4613_ = new_D3311_;
  assign new_B4612_ = new_D3244_;
  assign new_B4611_ = new_D3177_;
  assign new_B4610_ = new_D3110_;
  assign new_B4609_ = new_D3043_;
  assign new_B4608_ = new_D2976_;
  assign new_B4607_ = ~new_B4546_ & new_B4560_;
  assign new_B4606_ = new_B4546_ & ~new_B4560_;
  assign new_B4605_ = new_B4546_ & ~new_B4560_;
  assign new_B4604_ = ~new_B4546_ & ~new_B4560_;
  assign new_B4603_ = new_B4546_ & new_B4560_;
  assign new_B4602_ = new_B4606_ | new_B4607_;
  assign new_B4601_ = ~new_B4546_ & new_B4560_;
  assign new_B4600_ = new_B4604_ | new_B4605_;
  assign new_B4599_ = ~new_B4575_ & ~new_B4595_;
  assign new_B4598_ = new_B4575_ & new_B4595_;
  assign new_B4597_ = ~new_B4542_ | ~new_B4567_;
  assign new_B4596_ = new_B4560_ & new_B4597_;
  assign new_B4595_ = new_B4543_ | new_B4544_;
  assign new_B4594_ = new_B4543_ | new_B4560_;
  assign new_B4593_ = ~new_B4560_ & ~new_B4596_;
  assign new_B4592_ = new_B4560_ | new_B4597_;
  assign new_B4591_ = new_B4543_ & ~new_B4544_;
  assign new_B4590_ = ~new_B4543_ & new_B4544_;
  assign new_B4589_ = new_B4553_ | new_B4586_;
  assign new_B4588_ = ~new_B4553_ & ~new_B4587_;
  assign new_B4587_ = new_B4553_ & new_B4586_;
  assign new_B4586_ = ~new_B4542_ | ~new_B4567_;
  assign new_B4585_ = ~new_B4543_ & new_B4553_;
  assign new_B4584_ = new_B4543_ & ~new_B4553_;
  assign new_B4583_ = new_B4545_ & new_B4582_;
  assign new_B4582_ = new_B4601_ | new_B4600_;
  assign new_B4581_ = ~new_B4545_ & new_B4580_;
  assign new_B4580_ = new_B4603_ | new_B4602_;
  assign new_B4579_ = new_B4545_ | new_B4578_;
  assign new_B4578_ = new_B4599_ | new_B4598_;
  assign new_B4577_ = ~new_B4557_ & ~new_B4567_;
  assign new_B4576_ = new_B4557_ & new_B4567_;
  assign new_B4575_ = ~new_B4557_ | new_B4567_;
  assign new_B4574_ = new_B4541_ & ~new_B4542_;
  assign new_B4573_ = ~new_B4541_ & new_B4542_;
  assign new_B4572_ = new_B4594_ & ~new_B4595_;
  assign new_B4571_ = ~new_B4594_ & new_B4595_;
  assign new_B4570_ = ~new_B4593_ | ~new_B4592_;
  assign new_B4569_ = new_B4585_ | new_B4584_;
  assign new_B4568_ = new_B4591_ | new_B4590_;
  assign new_B4567_ = new_B4581_ | new_B4583_;
  assign new_B4566_ = ~new_B4588_ | ~new_B4589_;
  assign new_B4565_ = new_B4541_ & ~new_B4542_;
  assign new_B4564_ = new_B4555_ & ~new_B4567_;
  assign new_B4563_ = ~new_B4555_ & new_B4567_;
  assign new_B4562_ = ~new_B4553_ & new_B4579_;
  assign new_B4561_ = new_B4577_ | new_B4576_;
  assign new_B4560_ = new_B4574_ | new_B4573_;
  assign new_B4559_ = new_B4542_ | new_B4575_;
  assign new_B4558_ = new_B4567_ & new_B4570_;
  assign new_B4557_ = new_B4572_ | new_B4571_;
  assign new_B4556_ = new_B4567_ & new_B4566_;
  assign new_B4555_ = new_B4569_ & new_B4568_;
  assign new_B4554_ = new_B4564_ | new_B4563_;
  assign new_B4553_ = new_B4542_ | new_B4565_;
  assign B4552 = new_B4553_ | new_B4562_;
  assign B4551 = new_B4560_ & new_B4561_;
  assign B4550 = new_B4560_ & new_B4559_;
  assign B4549 = new_B4558_ | new_B4557_;
  assign B4548 = new_B4556_ | new_B4555_;
  assign B4547 = new_B4554_ & new_B4553_;
  assign new_B4546_ = new_D2909_;
  assign new_B4545_ = new_D2842_;
  assign new_B4544_ = new_D2775_;
  assign new_B4543_ = new_D2708_;
  assign new_B4542_ = new_D2641_;
  assign new_B4541_ = new_D2574_;
  assign new_B4540_ = ~new_B4479_ & new_B4493_;
  assign new_B4539_ = new_B4479_ & ~new_B4493_;
  assign new_B4538_ = new_B4479_ & ~new_B4493_;
  assign new_B4537_ = ~new_B4479_ & ~new_B4493_;
  assign new_B4536_ = new_B4479_ & new_B4493_;
  assign new_B4535_ = new_B4539_ | new_B4540_;
  assign new_B4534_ = ~new_B4479_ & new_B4493_;
  assign new_B4533_ = new_B4537_ | new_B4538_;
  assign new_B4532_ = ~new_B4508_ & ~new_B4528_;
  assign new_B4531_ = new_B4508_ & new_B4528_;
  assign new_B4530_ = ~new_B4475_ | ~new_B4500_;
  assign new_B4529_ = new_B4493_ & new_B4530_;
  assign new_B4528_ = new_B4476_ | new_B4477_;
  assign new_B4527_ = new_B4476_ | new_B4493_;
  assign new_B4526_ = ~new_B4493_ & ~new_B4529_;
  assign new_B4525_ = new_B4493_ | new_B4530_;
  assign new_B4524_ = new_B4476_ & ~new_B4477_;
  assign new_B4523_ = ~new_B4476_ & new_B4477_;
  assign new_B4522_ = new_B4486_ | new_B4519_;
  assign new_B4521_ = ~new_B4486_ & ~new_B4520_;
  assign new_B4520_ = new_B4486_ & new_B4519_;
  assign new_B4519_ = ~new_B4475_ | ~new_B4500_;
  assign new_B4518_ = ~new_B4476_ & new_B4486_;
  assign new_B4517_ = new_B4476_ & ~new_B4486_;
  assign new_B4516_ = new_B4478_ & new_B4515_;
  assign new_B4515_ = new_B4534_ | new_B4533_;
  assign new_B4514_ = ~new_B4478_ & new_B4513_;
  assign new_B4513_ = new_B4536_ | new_B4535_;
  assign new_B4512_ = new_B4478_ | new_B4511_;
  assign new_B4511_ = new_B4532_ | new_B4531_;
  assign new_B4510_ = ~new_B4490_ & ~new_B4500_;
  assign new_B4509_ = new_B4490_ & new_B4500_;
  assign new_B4508_ = ~new_B4490_ | new_B4500_;
  assign new_B4507_ = new_B4474_ & ~new_B4475_;
  assign new_B4506_ = ~new_B4474_ & new_B4475_;
  assign new_B4505_ = new_B4527_ & ~new_B4528_;
  assign new_B4504_ = ~new_B4527_ & new_B4528_;
  assign new_B4503_ = ~new_B4526_ | ~new_B4525_;
  assign new_B4502_ = new_B4518_ | new_B4517_;
  assign new_B4501_ = new_B4524_ | new_B4523_;
  assign new_B4500_ = new_B4514_ | new_B4516_;
  assign new_B4499_ = ~new_B4521_ | ~new_B4522_;
  assign new_B4498_ = new_B4474_ & ~new_B4475_;
  assign new_B4497_ = new_B4488_ & ~new_B4500_;
  assign new_B4496_ = ~new_B4488_ & new_B4500_;
  assign new_B4495_ = ~new_B4486_ & new_B4512_;
  assign new_B4494_ = new_B4510_ | new_B4509_;
  assign new_B4493_ = new_B4507_ | new_B4506_;
  assign new_B4492_ = new_B4475_ | new_B4508_;
  assign new_B4491_ = new_B4500_ & new_B4503_;
  assign new_B4490_ = new_B4505_ | new_B4504_;
  assign new_B4489_ = new_B4500_ & new_B4499_;
  assign new_B4488_ = new_B4502_ & new_B4501_;
  assign new_B4487_ = new_B4497_ | new_B4496_;
  assign new_B4486_ = new_B4475_ | new_B4498_;
  assign B4485 = new_B4486_ | new_B4495_;
  assign B4484 = new_B4493_ & new_B4494_;
  assign B4483 = new_B4493_ & new_B4492_;
  assign B4482 = new_B4491_ | new_B4490_;
  assign B4481 = new_B4489_ | new_B4488_;
  assign B4480 = new_B4487_ & new_B4486_;
  assign new_B4479_ = new_D2507_;
  assign new_B4478_ = new_D2440_;
  assign new_B4477_ = new_D2373_;
  assign new_B4476_ = new_D2306_;
  assign new_B4475_ = new_D2239_;
  assign new_B4474_ = new_D2172_;
  assign new_B4473_ = ~new_B4412_ & new_B4426_;
  assign new_B4472_ = new_B4412_ & ~new_B4426_;
  assign new_B4471_ = new_B4412_ & ~new_B4426_;
  assign new_B4470_ = ~new_B4412_ & ~new_B4426_;
  assign new_B4469_ = new_B4412_ & new_B4426_;
  assign new_B4468_ = new_B4472_ | new_B4473_;
  assign new_B4467_ = ~new_B4412_ & new_B4426_;
  assign new_B4466_ = new_B4470_ | new_B4471_;
  assign new_B4465_ = ~new_B4441_ & ~new_B4461_;
  assign new_B4464_ = new_B4441_ & new_B4461_;
  assign new_B4463_ = ~new_B4408_ | ~new_B4433_;
  assign new_B4462_ = new_B4426_ & new_B4463_;
  assign new_B4461_ = new_B4409_ | new_B4410_;
  assign new_B4460_ = new_B4409_ | new_B4426_;
  assign new_B4459_ = ~new_B4426_ & ~new_B4462_;
  assign new_B4458_ = new_B4426_ | new_B4463_;
  assign new_B4457_ = new_B4409_ & ~new_B4410_;
  assign new_B4456_ = ~new_B4409_ & new_B4410_;
  assign new_B4455_ = new_B4419_ | new_B4452_;
  assign new_B4454_ = ~new_B4419_ & ~new_B4453_;
  assign new_B4453_ = new_B4419_ & new_B4452_;
  assign new_B4452_ = ~new_B4408_ | ~new_B4433_;
  assign new_B4451_ = ~new_B4409_ & new_B4419_;
  assign new_B4450_ = new_B4409_ & ~new_B4419_;
  assign new_B4449_ = new_B4411_ & new_B4448_;
  assign new_B4448_ = new_B4467_ | new_B4466_;
  assign new_B4447_ = ~new_B4411_ & new_B4446_;
  assign new_B4446_ = new_B4469_ | new_B4468_;
  assign new_B4445_ = new_B4411_ | new_B4444_;
  assign new_B4444_ = new_B4465_ | new_B4464_;
  assign new_B4443_ = ~new_B4423_ & ~new_B4433_;
  assign new_B4442_ = new_B4423_ & new_B4433_;
  assign new_B4441_ = ~new_B4423_ | new_B4433_;
  assign new_B4440_ = new_B4407_ & ~new_B4408_;
  assign new_B4439_ = ~new_B4407_ & new_B4408_;
  assign new_B4438_ = new_B4460_ & ~new_B4461_;
  assign new_B4437_ = ~new_B4460_ & new_B4461_;
  assign new_B4436_ = ~new_B4459_ | ~new_B4458_;
  assign new_B4435_ = new_B4451_ | new_B4450_;
  assign new_B4434_ = new_B4457_ | new_B4456_;
  assign new_B4433_ = new_B4447_ | new_B4449_;
  assign new_B4432_ = ~new_B4454_ | ~new_B4455_;
  assign new_B4431_ = new_B4407_ & ~new_B4408_;
  assign new_B4430_ = new_B4421_ & ~new_B4433_;
  assign new_B4429_ = ~new_B4421_ & new_B4433_;
  assign new_B4428_ = ~new_B4419_ & new_B4445_;
  assign new_B4427_ = new_B4443_ | new_B4442_;
  assign new_B4426_ = new_B4440_ | new_B4439_;
  assign new_B4425_ = new_B4408_ | new_B4441_;
  assign new_B4424_ = new_B4433_ & new_B4436_;
  assign new_B4423_ = new_B4438_ | new_B4437_;
  assign new_B4422_ = new_B4433_ & new_B4432_;
  assign new_B4421_ = new_B4435_ & new_B4434_;
  assign new_B4420_ = new_B4430_ | new_B4429_;
  assign new_B4419_ = new_B4408_ | new_B4431_;
  assign B4418 = new_B4419_ | new_B4428_;
  assign B4417 = new_B4426_ & new_B4427_;
  assign B4416 = new_B4426_ & new_B4425_;
  assign B4415 = new_B4424_ | new_B4423_;
  assign B4414 = new_B4422_ | new_B4421_;
  assign B4413 = new_B4420_ & new_B4419_;
  assign new_B4412_ = new_D2105_;
  assign new_B4411_ = new_D2038_;
  assign new_B4410_ = new_D1971_;
  assign new_B4409_ = new_D1904_;
  assign new_B4408_ = new_D1837_;
  assign new_B4407_ = new_D1770_;
  assign new_B4406_ = ~new_B4345_ & new_B4359_;
  assign new_B4405_ = new_B4345_ & ~new_B4359_;
  assign new_B4404_ = new_B4345_ & ~new_B4359_;
  assign new_B4403_ = ~new_B4345_ & ~new_B4359_;
  assign new_B4402_ = new_B4345_ & new_B4359_;
  assign new_B4401_ = new_B4405_ | new_B4406_;
  assign new_B4400_ = ~new_B4345_ & new_B4359_;
  assign new_B4399_ = new_B4403_ | new_B4404_;
  assign new_B4398_ = ~new_B4374_ & ~new_B4394_;
  assign new_B4397_ = new_B4374_ & new_B4394_;
  assign new_B4396_ = ~new_B4341_ | ~new_B4366_;
  assign new_B4395_ = new_B4359_ & new_B4396_;
  assign new_B4394_ = new_B4342_ | new_B4343_;
  assign new_B4393_ = new_B4342_ | new_B4359_;
  assign new_B4392_ = ~new_B4359_ & ~new_B4395_;
  assign new_B4391_ = new_B4359_ | new_B4396_;
  assign new_B4390_ = new_B4342_ & ~new_B4343_;
  assign new_B4389_ = ~new_B4342_ & new_B4343_;
  assign new_B4388_ = new_B4352_ | new_B4385_;
  assign new_B4387_ = ~new_B4352_ & ~new_B4386_;
  assign new_B4386_ = new_B4352_ & new_B4385_;
  assign new_B4385_ = ~new_B4341_ | ~new_B4366_;
  assign new_B4384_ = ~new_B4342_ & new_B4352_;
  assign new_B4383_ = new_B4342_ & ~new_B4352_;
  assign new_B4382_ = new_B4344_ & new_B4381_;
  assign new_B4381_ = new_B4400_ | new_B4399_;
  assign new_B4380_ = ~new_B4344_ & new_B4379_;
  assign new_B4379_ = new_B4402_ | new_B4401_;
  assign new_B4378_ = new_B4344_ | new_B4377_;
  assign new_B4377_ = new_B4398_ | new_B4397_;
  assign new_B4376_ = ~new_B4356_ & ~new_B4366_;
  assign new_B4375_ = new_B4356_ & new_B4366_;
  assign new_B4374_ = ~new_B4356_ | new_B4366_;
  assign new_B4373_ = new_B4340_ & ~new_B4341_;
  assign new_B4372_ = ~new_B4340_ & new_B4341_;
  assign new_B4371_ = new_B4393_ & ~new_B4394_;
  assign new_B4370_ = ~new_B4393_ & new_B4394_;
  assign new_B4369_ = ~new_B4392_ | ~new_B4391_;
  assign new_B4368_ = new_B4384_ | new_B4383_;
  assign new_B4367_ = new_B4390_ | new_B4389_;
  assign new_B4366_ = new_B4380_ | new_B4382_;
  assign new_B4365_ = ~new_B4387_ | ~new_B4388_;
  assign new_B4364_ = new_B4340_ & ~new_B4341_;
  assign new_B4363_ = new_B4354_ & ~new_B4366_;
  assign new_B4362_ = ~new_B4354_ & new_B4366_;
  assign new_B4361_ = ~new_B4352_ & new_B4378_;
  assign new_B4360_ = new_B4376_ | new_B4375_;
  assign new_B4359_ = new_B4373_ | new_B4372_;
  assign new_B4358_ = new_B4341_ | new_B4374_;
  assign new_B4357_ = new_B4366_ & new_B4369_;
  assign new_B4356_ = new_B4371_ | new_B4370_;
  assign new_B4355_ = new_B4366_ & new_B4365_;
  assign new_B4354_ = new_B4368_ & new_B4367_;
  assign new_B4353_ = new_B4363_ | new_B4362_;
  assign new_B4352_ = new_B4341_ | new_B4364_;
  assign B4351 = new_B4352_ | new_B4361_;
  assign B4350 = new_B4359_ & new_B4360_;
  assign B4349 = new_B4359_ & new_B4358_;
  assign B4348 = new_B4357_ | new_B4356_;
  assign B4347 = new_B4355_ | new_B4354_;
  assign B4346 = new_B4353_ & new_B4352_;
  assign new_B4345_ = new_D1703_;
  assign new_B4344_ = new_D1636_;
  assign new_B4343_ = new_D1569_;
  assign new_B4342_ = new_D1502_;
  assign new_B4341_ = new_D1435_;
  assign new_B4340_ = new_D1368_;
  assign new_B4339_ = ~new_B4278_ & new_B4292_;
  assign new_B4338_ = new_B4278_ & ~new_B4292_;
  assign new_B4337_ = new_B4278_ & ~new_B4292_;
  assign new_B4336_ = ~new_B4278_ & ~new_B4292_;
  assign new_B4335_ = new_B4278_ & new_B4292_;
  assign new_B4334_ = new_B4338_ | new_B4339_;
  assign new_B4333_ = ~new_B4278_ & new_B4292_;
  assign new_B4332_ = new_B4336_ | new_B4337_;
  assign new_B4331_ = ~new_B4307_ & ~new_B4327_;
  assign new_B4330_ = new_B4307_ & new_B4327_;
  assign new_B4329_ = ~new_B4274_ | ~new_B4299_;
  assign new_B4328_ = new_B4292_ & new_B4329_;
  assign new_B4327_ = new_B4275_ | new_B4276_;
  assign new_B4326_ = new_B4275_ | new_B4292_;
  assign new_B4325_ = ~new_B4292_ & ~new_B4328_;
  assign new_B4324_ = new_B4292_ | new_B4329_;
  assign new_B4323_ = new_B4275_ & ~new_B4276_;
  assign new_B4322_ = ~new_B4275_ & new_B4276_;
  assign new_B4321_ = new_B4285_ | new_B4318_;
  assign new_B4320_ = ~new_B4285_ & ~new_B4319_;
  assign new_B4319_ = new_B4285_ & new_B4318_;
  assign new_B4318_ = ~new_B4274_ | ~new_B4299_;
  assign new_B4317_ = ~new_B4275_ & new_B4285_;
  assign new_B4316_ = new_B4275_ & ~new_B4285_;
  assign new_B4315_ = new_B4277_ & new_B4314_;
  assign new_B4314_ = new_B4333_ | new_B4332_;
  assign new_B4313_ = ~new_B4277_ & new_B4312_;
  assign new_B4312_ = new_B4335_ | new_B4334_;
  assign new_B4311_ = new_B4277_ | new_B4310_;
  assign new_B4310_ = new_B4331_ | new_B4330_;
  assign new_B4309_ = ~new_B4289_ & ~new_B4299_;
  assign new_B4308_ = new_B4289_ & new_B4299_;
  assign new_B4307_ = ~new_B4289_ | new_B4299_;
  assign new_B4306_ = new_B4273_ & ~new_B4274_;
  assign new_B4305_ = ~new_B4273_ & new_B4274_;
  assign new_B4304_ = new_B4326_ & ~new_B4327_;
  assign new_B4303_ = ~new_B4326_ & new_B4327_;
  assign new_B4302_ = ~new_B4325_ | ~new_B4324_;
  assign new_B4301_ = new_B4317_ | new_B4316_;
  assign new_B4300_ = new_B4323_ | new_B4322_;
  assign new_B4299_ = new_B4313_ | new_B4315_;
  assign new_B4298_ = ~new_B4320_ | ~new_B4321_;
  assign new_B4297_ = new_B4273_ & ~new_B4274_;
  assign new_B4296_ = new_B4287_ & ~new_B4299_;
  assign new_B4295_ = ~new_B4287_ & new_B4299_;
  assign new_B4294_ = ~new_B4285_ & new_B4311_;
  assign new_B4293_ = new_B4309_ | new_B4308_;
  assign new_B4292_ = new_B4306_ | new_B4305_;
  assign new_B4291_ = new_B4274_ | new_B4307_;
  assign new_B4290_ = new_B4299_ & new_B4302_;
  assign new_B4289_ = new_B4304_ | new_B4303_;
  assign new_B4288_ = new_B4299_ & new_B4298_;
  assign new_B4287_ = new_B4301_ & new_B4300_;
  assign new_B4286_ = new_B4296_ | new_B4295_;
  assign new_B4285_ = new_B4274_ | new_B4297_;
  assign B4284 = new_B4285_ | new_B4294_;
  assign B4283 = new_B4292_ & new_B4293_;
  assign B4282 = new_B4292_ & new_B4291_;
  assign B4281 = new_B4290_ | new_B4289_;
  assign B4280 = new_B4288_ | new_B4287_;
  assign B4279 = new_B4286_ & new_B4285_;
  assign new_B4278_ = new_D1301_;
  assign new_B4277_ = new_D1234_;
  assign new_B4276_ = new_D1167_;
  assign new_B4275_ = new_D1100_;
  assign new_B4274_ = new_D1033_;
  assign new_B4273_ = new_D966_;
  assign new_B4272_ = ~new_B4211_ & new_B4225_;
  assign new_B4271_ = new_B4211_ & ~new_B4225_;
  assign new_B4270_ = new_B4211_ & ~new_B4225_;
  assign new_B4269_ = ~new_B4211_ & ~new_B4225_;
  assign new_B4268_ = new_B4211_ & new_B4225_;
  assign new_B4267_ = new_B4271_ | new_B4272_;
  assign new_B4266_ = ~new_B4211_ & new_B4225_;
  assign new_B4265_ = new_B4269_ | new_B4270_;
  assign new_B4264_ = ~new_B4240_ & ~new_B4260_;
  assign new_B4263_ = new_B4240_ & new_B4260_;
  assign new_B4262_ = ~new_B4207_ | ~new_B4232_;
  assign new_B4261_ = new_B4225_ & new_B4262_;
  assign new_B4260_ = new_B4208_ | new_B4209_;
  assign new_B4259_ = new_B4208_ | new_B4225_;
  assign new_B4258_ = ~new_B4225_ & ~new_B4261_;
  assign new_B4257_ = new_B4225_ | new_B4262_;
  assign new_B4256_ = new_B4208_ & ~new_B4209_;
  assign new_B4255_ = ~new_B4208_ & new_B4209_;
  assign new_B4254_ = new_B4218_ | new_B4251_;
  assign new_B4253_ = ~new_B4218_ & ~new_B4252_;
  assign new_B4252_ = new_B4218_ & new_B4251_;
  assign new_B4251_ = ~new_B4207_ | ~new_B4232_;
  assign new_B4250_ = ~new_B4208_ & new_B4218_;
  assign new_B4249_ = new_B4208_ & ~new_B4218_;
  assign new_B4248_ = new_B4210_ & new_B4247_;
  assign new_B4247_ = new_B4266_ | new_B4265_;
  assign new_B4246_ = ~new_B4210_ & new_B4245_;
  assign new_B4245_ = new_B4268_ | new_B4267_;
  assign new_B4244_ = new_B4210_ | new_B4243_;
  assign new_B4243_ = new_B4264_ | new_B4263_;
  assign new_B4242_ = ~new_B4222_ & ~new_B4232_;
  assign new_B4241_ = new_B4222_ & new_B4232_;
  assign new_B4240_ = ~new_B4222_ | new_B4232_;
  assign new_B4239_ = new_B4206_ & ~new_B4207_;
  assign new_B4238_ = ~new_B4206_ & new_B4207_;
  assign new_B4237_ = new_B4259_ & ~new_B4260_;
  assign new_B4236_ = ~new_B4259_ & new_B4260_;
  assign new_B4235_ = ~new_B4258_ | ~new_B4257_;
  assign new_B4234_ = new_B4250_ | new_B4249_;
  assign new_B4233_ = new_B4256_ | new_B4255_;
  assign new_B4232_ = new_B4246_ | new_B4248_;
  assign new_B4231_ = ~new_B4253_ | ~new_B4254_;
  assign new_B4230_ = new_B4206_ & ~new_B4207_;
  assign new_B4229_ = new_B4220_ & ~new_B4232_;
  assign new_B4228_ = ~new_B4220_ & new_B4232_;
  assign new_B4227_ = ~new_B4218_ & new_B4244_;
  assign new_B4226_ = new_B4242_ | new_B4241_;
  assign new_B4225_ = new_B4239_ | new_B4238_;
  assign new_B4224_ = new_B4207_ | new_B4240_;
  assign new_B4223_ = new_B4232_ & new_B4235_;
  assign new_B4222_ = new_B4237_ | new_B4236_;
  assign new_B4221_ = new_B4232_ & new_B4231_;
  assign new_B4220_ = new_B4234_ & new_B4233_;
  assign new_B4219_ = new_B4229_ | new_B4228_;
  assign new_B4218_ = new_B4207_ | new_B4230_;
  assign B4217 = new_B4218_ | new_B4227_;
  assign B4216 = new_B4225_ & new_B4226_;
  assign B4215 = new_B4225_ & new_B4224_;
  assign B4214 = new_B4223_ | new_B4222_;
  assign B4213 = new_B4221_ | new_B4220_;
  assign B4212 = new_B4219_ & new_B4218_;
  assign new_B4211_ = new_D899_;
  assign new_B4210_ = new_D832_;
  assign new_B4209_ = new_D765_;
  assign new_B4208_ = new_D698_;
  assign new_B4207_ = new_D631_;
  assign new_B4206_ = new_D564_;
  assign new_B4205_ = ~new_B4144_ & new_B4158_;
  assign new_B4204_ = new_B4144_ & ~new_B4158_;
  assign new_B4203_ = new_B4144_ & ~new_B4158_;
  assign new_B4202_ = ~new_B4144_ & ~new_B4158_;
  assign new_B4201_ = new_B4144_ & new_B4158_;
  assign new_B4200_ = new_B4204_ | new_B4205_;
  assign new_B4199_ = ~new_B4144_ & new_B4158_;
  assign new_B4198_ = new_B4202_ | new_B4203_;
  assign new_B4197_ = ~new_B4173_ & ~new_B4193_;
  assign new_B4196_ = new_B4173_ & new_B4193_;
  assign new_B4195_ = ~new_B4140_ | ~new_B4165_;
  assign new_B4194_ = new_B4158_ & new_B4195_;
  assign new_B4193_ = new_B4141_ | new_B4142_;
  assign new_B4192_ = new_B4141_ | new_B4158_;
  assign new_B4191_ = ~new_B4158_ & ~new_B4194_;
  assign new_B4190_ = new_B4158_ | new_B4195_;
  assign new_B4189_ = new_B4141_ & ~new_B4142_;
  assign new_B4188_ = ~new_B4141_ & new_B4142_;
  assign new_B4187_ = new_B4151_ | new_B4184_;
  assign new_B4186_ = ~new_B4151_ & ~new_B4185_;
  assign new_B4185_ = new_B4151_ & new_B4184_;
  assign new_B4184_ = ~new_B4140_ | ~new_B4165_;
  assign new_B4183_ = ~new_B4141_ & new_B4151_;
  assign new_B4182_ = new_B4141_ & ~new_B4151_;
  assign new_B4181_ = new_B4143_ & new_B4180_;
  assign new_B4180_ = new_B4199_ | new_B4198_;
  assign new_B4179_ = ~new_B4143_ & new_B4178_;
  assign new_B4178_ = new_B4201_ | new_B4200_;
  assign new_B4177_ = new_B4143_ | new_B4176_;
  assign new_B4176_ = new_B4197_ | new_B4196_;
  assign new_B4175_ = ~new_B4155_ & ~new_B4165_;
  assign new_B4174_ = new_B4155_ & new_B4165_;
  assign new_B4173_ = ~new_B4155_ | new_B4165_;
  assign new_B4172_ = new_B4139_ & ~new_B4140_;
  assign new_B4171_ = ~new_B4139_ & new_B4140_;
  assign new_B4170_ = new_B4192_ & ~new_B4193_;
  assign new_B4169_ = ~new_B4192_ & new_B4193_;
  assign new_B4168_ = ~new_B4191_ | ~new_B4190_;
  assign new_B4167_ = new_B4183_ | new_B4182_;
  assign new_B4166_ = new_B4189_ | new_B4188_;
  assign new_B4165_ = new_B4179_ | new_B4181_;
  assign new_B4164_ = ~new_B4186_ | ~new_B4187_;
  assign new_B4163_ = new_B4139_ & ~new_B4140_;
  assign new_B4162_ = new_B4153_ & ~new_B4165_;
  assign new_B4161_ = ~new_B4153_ & new_B4165_;
  assign new_B4160_ = ~new_B4151_ & new_B4177_;
  assign new_B4159_ = new_B4175_ | new_B4174_;
  assign new_B4158_ = new_B4172_ | new_B4171_;
  assign new_B4157_ = new_B4140_ | new_B4173_;
  assign new_B4156_ = new_B4165_ & new_B4168_;
  assign new_B4155_ = new_B4170_ | new_B4169_;
  assign new_B4154_ = new_B4165_ & new_B4164_;
  assign new_B4153_ = new_B4167_ & new_B4166_;
  assign new_B4152_ = new_B4162_ | new_B4161_;
  assign new_B4151_ = new_B4140_ | new_B4163_;
  assign B4150 = new_B4151_ | new_B4160_;
  assign B4149 = new_B4158_ & new_B4159_;
  assign B4148 = new_B4158_ & new_B4157_;
  assign B4147 = new_B4156_ | new_B4155_;
  assign B4146 = new_B4154_ | new_B4153_;
  assign B4145 = new_B4152_ & new_B4151_;
  assign new_B4144_ = new_D497_;
  assign new_B4143_ = new_D430_;
  assign new_B4142_ = new_D363_;
  assign new_B4141_ = new_D296_;
  assign new_B4140_ = new_D229_;
  assign new_B4139_ = new_D162_;
  assign new_B4138_ = ~new_B4077_ & new_B4091_;
  assign new_B4137_ = new_B4077_ & ~new_B4091_;
  assign new_B4136_ = new_B4077_ & ~new_B4091_;
  assign new_B4135_ = ~new_B4077_ & ~new_B4091_;
  assign new_B4134_ = new_B4077_ & new_B4091_;
  assign new_B4133_ = new_B4137_ | new_B4138_;
  assign new_B4132_ = ~new_B4077_ & new_B4091_;
  assign new_B4131_ = new_B4135_ | new_B4136_;
  assign new_B4130_ = ~new_B4106_ & ~new_B4126_;
  assign new_B4129_ = new_B4106_ & new_B4126_;
  assign new_B4128_ = ~new_B4073_ | ~new_B4098_;
  assign new_B4127_ = new_B4091_ & new_B4128_;
  assign new_B4126_ = new_B4074_ | new_B4075_;
  assign new_B4125_ = new_B4074_ | new_B4091_;
  assign new_B4124_ = ~new_B4091_ & ~new_B4127_;
  assign new_B4123_ = new_B4091_ | new_B4128_;
  assign new_B4122_ = new_B4074_ & ~new_B4075_;
  assign new_B4121_ = ~new_B4074_ & new_B4075_;
  assign new_B4120_ = new_B4084_ | new_B4117_;
  assign new_B4119_ = ~new_B4084_ & ~new_B4118_;
  assign new_B4118_ = new_B4084_ & new_B4117_;
  assign new_B4117_ = ~new_B4073_ | ~new_B4098_;
  assign new_B4116_ = ~new_B4074_ & new_B4084_;
  assign new_B4115_ = new_B4074_ & ~new_B4084_;
  assign new_B4114_ = new_B4076_ & new_B4113_;
  assign new_B4113_ = new_B4132_ | new_B4131_;
  assign new_B4112_ = ~new_B4076_ & new_B4111_;
  assign new_B4111_ = new_B4134_ | new_B4133_;
  assign new_B4110_ = new_B4076_ | new_B4109_;
  assign new_B4109_ = new_B4130_ | new_B4129_;
  assign new_B4108_ = ~new_B4088_ & ~new_B4098_;
  assign new_B4107_ = new_B4088_ & new_B4098_;
  assign new_B4106_ = ~new_B4088_ | new_B4098_;
  assign new_B4105_ = new_B4072_ & ~new_B4073_;
  assign new_B4104_ = ~new_B4072_ & new_B4073_;
  assign new_B4103_ = new_B4125_ & ~new_B4126_;
  assign new_B4102_ = ~new_B4125_ & new_B4126_;
  assign new_B4101_ = ~new_B4124_ | ~new_B4123_;
  assign new_B4100_ = new_B4116_ | new_B4115_;
  assign new_B4099_ = new_B4122_ | new_B4121_;
  assign new_B4098_ = new_B4112_ | new_B4114_;
  assign new_B4097_ = ~new_B4119_ | ~new_B4120_;
  assign new_B4096_ = new_B4072_ & ~new_B4073_;
  assign new_B4095_ = new_B4086_ & ~new_B4098_;
  assign new_B4094_ = ~new_B4086_ & new_B4098_;
  assign new_B4093_ = ~new_B4084_ & new_B4110_;
  assign new_B4092_ = new_B4108_ | new_B4107_;
  assign new_B4091_ = new_B4105_ | new_B4104_;
  assign new_B4090_ = new_B4073_ | new_B4106_;
  assign new_B4089_ = new_B4098_ & new_B4101_;
  assign new_B4088_ = new_B4103_ | new_B4102_;
  assign new_B4087_ = new_B4098_ & new_B4097_;
  assign new_B4086_ = new_B4100_ & new_B4099_;
  assign new_B4085_ = new_B4095_ | new_B4094_;
  assign new_B4084_ = new_B4073_ | new_B4096_;
  assign B4083 = new_B4084_ | new_B4093_;
  assign B4082 = new_B4091_ & new_B4092_;
  assign B4081 = new_B4091_ & new_B4090_;
  assign B4080 = new_B4089_ | new_B4088_;
  assign B4079 = new_B4087_ | new_B4086_;
  assign B4078 = new_B4085_ & new_B4084_;
  assign new_B4077_ = new_D95_;
  assign new_B4076_ = new_D28_;
  assign new_B4075_ = new_C9960_;
  assign new_B4074_ = new_C9893_;
  assign new_B4073_ = new_C9826_;
  assign new_B4072_ = new_C9759_;
  assign new_B4071_ = ~new_B4010_ & new_B4024_;
  assign new_B4070_ = new_B4010_ & ~new_B4024_;
  assign new_B4069_ = new_B4010_ & ~new_B4024_;
  assign new_B4068_ = ~new_B4010_ & ~new_B4024_;
  assign new_B4067_ = new_B4010_ & new_B4024_;
  assign new_B4066_ = new_B4070_ | new_B4071_;
  assign new_B4065_ = ~new_B4010_ & new_B4024_;
  assign new_B4064_ = new_B4068_ | new_B4069_;
  assign new_B4063_ = ~new_B4039_ & ~new_B4059_;
  assign new_B4062_ = new_B4039_ & new_B4059_;
  assign new_B4061_ = ~new_B4006_ | ~new_B4031_;
  assign new_B4060_ = new_B4024_ & new_B4061_;
  assign new_B4059_ = new_B4007_ | new_B4008_;
  assign new_B4058_ = new_B4007_ | new_B4024_;
  assign new_B4057_ = ~new_B4024_ & ~new_B4060_;
  assign new_B4056_ = new_B4024_ | new_B4061_;
  assign new_B4055_ = new_B4007_ & ~new_B4008_;
  assign new_B4054_ = ~new_B4007_ & new_B4008_;
  assign new_B4053_ = new_B4017_ | new_B4050_;
  assign new_B4052_ = ~new_B4017_ & ~new_B4051_;
  assign new_B4051_ = new_B4017_ & new_B4050_;
  assign new_B4050_ = ~new_B4006_ | ~new_B4031_;
  assign new_B4049_ = ~new_B4007_ & new_B4017_;
  assign new_B4048_ = new_B4007_ & ~new_B4017_;
  assign new_B4047_ = new_B4009_ & new_B4046_;
  assign new_B4046_ = new_B4065_ | new_B4064_;
  assign new_B4045_ = ~new_B4009_ & new_B4044_;
  assign new_B4044_ = new_B4067_ | new_B4066_;
  assign new_B4043_ = new_B4009_ | new_B4042_;
  assign new_B4042_ = new_B4063_ | new_B4062_;
  assign new_B4041_ = ~new_B4021_ & ~new_B4031_;
  assign new_B4040_ = new_B4021_ & new_B4031_;
  assign new_B4039_ = ~new_B4021_ | new_B4031_;
  assign new_B4038_ = new_B4005_ & ~new_B4006_;
  assign new_B4037_ = ~new_B4005_ & new_B4006_;
  assign new_B4036_ = new_B4058_ & ~new_B4059_;
  assign new_B4035_ = ~new_B4058_ & new_B4059_;
  assign new_B4034_ = ~new_B4057_ | ~new_B4056_;
  assign new_B4033_ = new_B4049_ | new_B4048_;
  assign new_B4032_ = new_B4055_ | new_B4054_;
  assign new_B4031_ = new_B4045_ | new_B4047_;
  assign new_B4030_ = ~new_B4052_ | ~new_B4053_;
  assign new_B4029_ = new_B4005_ & ~new_B4006_;
  assign new_B4028_ = new_B4019_ & ~new_B4031_;
  assign new_B4027_ = ~new_B4019_ & new_B4031_;
  assign new_B4026_ = ~new_B4017_ & new_B4043_;
  assign new_B4025_ = new_B4041_ | new_B4040_;
  assign new_B4024_ = new_B4038_ | new_B4037_;
  assign new_B4023_ = new_B4006_ | new_B4039_;
  assign new_B4022_ = new_B4031_ & new_B4034_;
  assign new_B4021_ = new_B4036_ | new_B4035_;
  assign new_B4020_ = new_B4031_ & new_B4030_;
  assign new_B4019_ = new_B4033_ & new_B4032_;
  assign new_B4018_ = new_B4028_ | new_B4027_;
  assign new_B4017_ = new_B4006_ | new_B4029_;
  assign B4016 = new_B4017_ | new_B4026_;
  assign B4015 = new_B4024_ & new_B4025_;
  assign B4014 = new_B4024_ & new_B4023_;
  assign B4013 = new_B4022_ | new_B4021_;
  assign B4012 = new_B4020_ | new_B4019_;
  assign B4011 = new_B4018_ & new_B4017_;
  assign new_B4010_ = new_C9692_;
  assign new_B4009_ = new_C9625_;
  assign new_B4008_ = new_C9558_;
  assign new_B4007_ = new_C9491_;
  assign new_B4006_ = new_C9424_;
  assign new_B4005_ = new_C9357_;
  assign new_B4004_ = ~new_B3943_ & new_B3957_;
  assign new_B4003_ = new_B3943_ & ~new_B3957_;
  assign new_B4002_ = new_B3943_ & ~new_B3957_;
  assign new_B4001_ = ~new_B3943_ & ~new_B3957_;
  assign new_B4000_ = new_B3943_ & new_B3957_;
  assign new_B3999_ = new_B4003_ | new_B4004_;
  assign new_B3998_ = ~new_B3943_ & new_B3957_;
  assign new_B3997_ = new_B4001_ | new_B4002_;
  assign new_B3996_ = ~new_B3972_ & ~new_B3992_;
  assign new_B3995_ = new_B3972_ & new_B3992_;
  assign new_B3994_ = ~new_B3939_ | ~new_B3964_;
  assign new_B3993_ = new_B3957_ & new_B3994_;
  assign new_B3992_ = new_B3940_ | new_B3941_;
  assign new_B3991_ = new_B3940_ | new_B3957_;
  assign new_B3990_ = ~new_B3957_ & ~new_B3993_;
  assign new_B3989_ = new_B3957_ | new_B3994_;
  assign new_B3988_ = new_B3940_ & ~new_B3941_;
  assign new_B3987_ = ~new_B3940_ & new_B3941_;
  assign new_B3986_ = new_B3950_ | new_B3983_;
  assign new_B3985_ = ~new_B3950_ & ~new_B3984_;
  assign new_B3984_ = new_B3950_ & new_B3983_;
  assign new_B3983_ = ~new_B3939_ | ~new_B3964_;
  assign new_B3982_ = ~new_B3940_ & new_B3950_;
  assign new_B3981_ = new_B3940_ & ~new_B3950_;
  assign new_B3980_ = new_B3942_ & new_B3979_;
  assign new_B3979_ = new_B3998_ | new_B3997_;
  assign new_B3978_ = ~new_B3942_ & new_B3977_;
  assign new_B3977_ = new_B4000_ | new_B3999_;
  assign new_B3976_ = new_B3942_ | new_B3975_;
  assign new_B3975_ = new_B3996_ | new_B3995_;
  assign new_B3974_ = ~new_B3954_ & ~new_B3964_;
  assign new_B3973_ = new_B3954_ & new_B3964_;
  assign new_B3972_ = ~new_B3954_ | new_B3964_;
  assign new_B3971_ = new_B3938_ & ~new_B3939_;
  assign new_B3970_ = ~new_B3938_ & new_B3939_;
  assign new_B3969_ = new_B3991_ & ~new_B3992_;
  assign new_B3968_ = ~new_B3991_ & new_B3992_;
  assign new_B3967_ = ~new_B3990_ | ~new_B3989_;
  assign new_B3966_ = new_B3982_ | new_B3981_;
  assign new_B3965_ = new_B3988_ | new_B3987_;
  assign new_B3964_ = new_B3978_ | new_B3980_;
  assign new_B3963_ = ~new_B3985_ | ~new_B3986_;
  assign new_B3962_ = new_B3938_ & ~new_B3939_;
  assign new_B3961_ = new_B3952_ & ~new_B3964_;
  assign new_B3960_ = ~new_B3952_ & new_B3964_;
  assign new_B3959_ = ~new_B3950_ & new_B3976_;
  assign new_B3958_ = new_B3974_ | new_B3973_;
  assign new_B3957_ = new_B3971_ | new_B3970_;
  assign new_B3956_ = new_B3939_ | new_B3972_;
  assign new_B3955_ = new_B3964_ & new_B3967_;
  assign new_B3954_ = new_B3969_ | new_B3968_;
  assign new_B3953_ = new_B3964_ & new_B3963_;
  assign new_B3952_ = new_B3966_ & new_B3965_;
  assign new_B3951_ = new_B3961_ | new_B3960_;
  assign new_B3950_ = new_B3939_ | new_B3962_;
  assign B3949 = new_B3950_ | new_B3959_;
  assign B3948 = new_B3957_ & new_B3958_;
  assign B3947 = new_B3957_ & new_B3956_;
  assign B3946 = new_B3955_ | new_B3954_;
  assign B3945 = new_B3953_ | new_B3952_;
  assign B3944 = new_B3951_ & new_B3950_;
  assign new_B3943_ = new_C9290_;
  assign new_B3942_ = new_C9223_;
  assign new_B3941_ = new_C9156_;
  assign new_B3940_ = new_C9089_;
  assign new_B3939_ = new_C9022_;
  assign new_B3938_ = new_C8955_;
  assign new_B3937_ = ~new_B3876_ & new_B3890_;
  assign new_B3936_ = new_B3876_ & ~new_B3890_;
  assign new_B3935_ = new_B3876_ & ~new_B3890_;
  assign new_B3934_ = ~new_B3876_ & ~new_B3890_;
  assign new_B3933_ = new_B3876_ & new_B3890_;
  assign new_B3932_ = new_B3936_ | new_B3937_;
  assign new_B3931_ = ~new_B3876_ & new_B3890_;
  assign new_B3930_ = new_B3934_ | new_B3935_;
  assign new_B3929_ = ~new_B3905_ & ~new_B3925_;
  assign new_B3928_ = new_B3905_ & new_B3925_;
  assign new_B3927_ = ~new_B3872_ | ~new_B3897_;
  assign new_B3926_ = new_B3890_ & new_B3927_;
  assign new_B3925_ = new_B3873_ | new_B3874_;
  assign new_B3924_ = new_B3873_ | new_B3890_;
  assign new_B3923_ = ~new_B3890_ & ~new_B3926_;
  assign new_B3922_ = new_B3890_ | new_B3927_;
  assign new_B3921_ = new_B3873_ & ~new_B3874_;
  assign new_B3920_ = ~new_B3873_ & new_B3874_;
  assign new_B3919_ = new_B3883_ | new_B3916_;
  assign new_B3918_ = ~new_B3883_ & ~new_B3917_;
  assign new_B3917_ = new_B3883_ & new_B3916_;
  assign new_B3916_ = ~new_B3872_ | ~new_B3897_;
  assign new_B3915_ = ~new_B3873_ & new_B3883_;
  assign new_B3914_ = new_B3873_ & ~new_B3883_;
  assign new_B3913_ = new_B3875_ & new_B3912_;
  assign new_B3912_ = new_B3931_ | new_B3930_;
  assign new_B3911_ = ~new_B3875_ & new_B3910_;
  assign new_B3910_ = new_B3933_ | new_B3932_;
  assign new_B3909_ = new_B3875_ | new_B3908_;
  assign new_B3908_ = new_B3929_ | new_B3928_;
  assign new_B3907_ = ~new_B3887_ & ~new_B3897_;
  assign new_B3906_ = new_B3887_ & new_B3897_;
  assign new_B3905_ = ~new_B3887_ | new_B3897_;
  assign new_B3904_ = new_B3871_ & ~new_B3872_;
  assign new_B3903_ = ~new_B3871_ & new_B3872_;
  assign new_B3902_ = new_B3924_ & ~new_B3925_;
  assign new_B3901_ = ~new_B3924_ & new_B3925_;
  assign new_B3900_ = ~new_B3923_ | ~new_B3922_;
  assign new_B3899_ = new_B3915_ | new_B3914_;
  assign new_B3898_ = new_B3921_ | new_B3920_;
  assign new_B3897_ = new_B3911_ | new_B3913_;
  assign new_B3896_ = ~new_B3918_ | ~new_B3919_;
  assign new_B3895_ = new_B3871_ & ~new_B3872_;
  assign new_B3894_ = new_B3885_ & ~new_B3897_;
  assign new_B3893_ = ~new_B3885_ & new_B3897_;
  assign new_B3892_ = ~new_B3883_ & new_B3909_;
  assign new_B3891_ = new_B3907_ | new_B3906_;
  assign new_B3890_ = new_B3904_ | new_B3903_;
  assign new_B3889_ = new_B3872_ | new_B3905_;
  assign new_B3888_ = new_B3897_ & new_B3900_;
  assign new_B3887_ = new_B3902_ | new_B3901_;
  assign new_B3886_ = new_B3897_ & new_B3896_;
  assign new_B3885_ = new_B3899_ & new_B3898_;
  assign new_B3884_ = new_B3894_ | new_B3893_;
  assign new_B3883_ = new_B3872_ | new_B3895_;
  assign B3882 = new_B3883_ | new_B3892_;
  assign B3881 = new_B3890_ & new_B3891_;
  assign B3880 = new_B3890_ & new_B3889_;
  assign B3879 = new_B3888_ | new_B3887_;
  assign B3878 = new_B3886_ | new_B3885_;
  assign B3877 = new_B3884_ & new_B3883_;
  assign new_B3876_ = new_C8888_;
  assign new_B3875_ = new_C8821_;
  assign new_B3874_ = new_C8754_;
  assign new_B3873_ = new_C8687_;
  assign new_B3872_ = new_C8620_;
  assign new_B3871_ = new_C8553_;
  assign new_B3870_ = ~new_B3809_ & new_B3823_;
  assign new_B3869_ = new_B3809_ & ~new_B3823_;
  assign new_B3868_ = new_B3809_ & ~new_B3823_;
  assign new_B3867_ = ~new_B3809_ & ~new_B3823_;
  assign new_B3866_ = new_B3809_ & new_B3823_;
  assign new_B3865_ = new_B3869_ | new_B3870_;
  assign new_B3864_ = ~new_B3809_ & new_B3823_;
  assign new_B3863_ = new_B3867_ | new_B3868_;
  assign new_B3862_ = ~new_B3838_ & ~new_B3858_;
  assign new_B3861_ = new_B3838_ & new_B3858_;
  assign new_B3860_ = ~new_B3805_ | ~new_B3830_;
  assign new_B3859_ = new_B3823_ & new_B3860_;
  assign new_B3858_ = new_B3806_ | new_B3807_;
  assign new_B3857_ = new_B3806_ | new_B3823_;
  assign new_B3856_ = ~new_B3823_ & ~new_B3859_;
  assign new_B3855_ = new_B3823_ | new_B3860_;
  assign new_B3854_ = new_B3806_ & ~new_B3807_;
  assign new_B3853_ = ~new_B3806_ & new_B3807_;
  assign new_B3852_ = new_B3816_ | new_B3849_;
  assign new_B3851_ = ~new_B3816_ & ~new_B3850_;
  assign new_B3850_ = new_B3816_ & new_B3849_;
  assign new_B3849_ = ~new_B3805_ | ~new_B3830_;
  assign new_B3848_ = ~new_B3806_ & new_B3816_;
  assign new_B3847_ = new_B3806_ & ~new_B3816_;
  assign new_B3846_ = new_B3808_ & new_B3845_;
  assign new_B3845_ = new_B3864_ | new_B3863_;
  assign new_B3844_ = ~new_B3808_ & new_B3843_;
  assign new_B3843_ = new_B3866_ | new_B3865_;
  assign new_B3842_ = new_B3808_ | new_B3841_;
  assign new_B3841_ = new_B3862_ | new_B3861_;
  assign new_B3840_ = ~new_B3820_ & ~new_B3830_;
  assign new_B3839_ = new_B3820_ & new_B3830_;
  assign new_B3838_ = ~new_B3820_ | new_B3830_;
  assign new_B3837_ = new_B3804_ & ~new_B3805_;
  assign new_B3836_ = ~new_B3804_ & new_B3805_;
  assign new_B3835_ = new_B3857_ & ~new_B3858_;
  assign new_B3834_ = ~new_B3857_ & new_B3858_;
  assign new_B3833_ = ~new_B3856_ | ~new_B3855_;
  assign new_B3832_ = new_B3848_ | new_B3847_;
  assign new_B3831_ = new_B3854_ | new_B3853_;
  assign new_B3830_ = new_B3844_ | new_B3846_;
  assign new_B3829_ = ~new_B3851_ | ~new_B3852_;
  assign new_B3828_ = new_B3804_ & ~new_B3805_;
  assign new_B3827_ = new_B3818_ & ~new_B3830_;
  assign new_B3826_ = ~new_B3818_ & new_B3830_;
  assign new_B3825_ = ~new_B3816_ & new_B3842_;
  assign new_B3824_ = new_B3840_ | new_B3839_;
  assign new_B3823_ = new_B3837_ | new_B3836_;
  assign new_B3822_ = new_B3805_ | new_B3838_;
  assign new_B3821_ = new_B3830_ & new_B3833_;
  assign new_B3820_ = new_B3835_ | new_B3834_;
  assign new_B3819_ = new_B3830_ & new_B3829_;
  assign new_B3818_ = new_B3832_ & new_B3831_;
  assign new_B3817_ = new_B3827_ | new_B3826_;
  assign new_B3816_ = new_B3805_ | new_B3828_;
  assign B3815 = new_B3816_ | new_B3825_;
  assign B3814 = new_B3823_ & new_B3824_;
  assign B3813 = new_B3823_ & new_B3822_;
  assign B3812 = new_B3821_ | new_B3820_;
  assign B3811 = new_B3819_ | new_B3818_;
  assign B3810 = new_B3817_ & new_B3816_;
  assign new_B3809_ = new_C8486_;
  assign new_B3808_ = new_C8419_;
  assign new_B3807_ = new_C8352_;
  assign new_B3806_ = new_C8285_;
  assign new_B3805_ = new_C8218_;
  assign new_B3804_ = new_C8151_;
  assign new_B3803_ = ~new_B3742_ & new_B3756_;
  assign new_B3802_ = new_B3742_ & ~new_B3756_;
  assign new_B3801_ = new_B3742_ & ~new_B3756_;
  assign new_B3800_ = ~new_B3742_ & ~new_B3756_;
  assign new_B3799_ = new_B3742_ & new_B3756_;
  assign new_B3798_ = new_B3802_ | new_B3803_;
  assign new_B3797_ = ~new_B3742_ & new_B3756_;
  assign new_B3796_ = new_B3800_ | new_B3801_;
  assign new_B3795_ = ~new_B3771_ & ~new_B3791_;
  assign new_B3794_ = new_B3771_ & new_B3791_;
  assign new_B3793_ = ~new_B3738_ | ~new_B3763_;
  assign new_B3792_ = new_B3756_ & new_B3793_;
  assign new_B3791_ = new_B3739_ | new_B3740_;
  assign new_B3790_ = new_B3739_ | new_B3756_;
  assign new_B3789_ = ~new_B3756_ & ~new_B3792_;
  assign new_B3788_ = new_B3756_ | new_B3793_;
  assign new_B3787_ = new_B3739_ & ~new_B3740_;
  assign new_B3786_ = ~new_B3739_ & new_B3740_;
  assign new_B3785_ = new_B3749_ | new_B3782_;
  assign new_B3784_ = ~new_B3749_ & ~new_B3783_;
  assign new_B3783_ = new_B3749_ & new_B3782_;
  assign new_B3782_ = ~new_B3738_ | ~new_B3763_;
  assign new_B3781_ = ~new_B3739_ & new_B3749_;
  assign new_B3780_ = new_B3739_ & ~new_B3749_;
  assign new_B3779_ = new_B3741_ & new_B3778_;
  assign new_B3778_ = new_B3797_ | new_B3796_;
  assign new_B3777_ = ~new_B3741_ & new_B3776_;
  assign new_B3776_ = new_B3799_ | new_B3798_;
  assign new_B3775_ = new_B3741_ | new_B3774_;
  assign new_B3774_ = new_B3795_ | new_B3794_;
  assign new_B3773_ = ~new_B3753_ & ~new_B3763_;
  assign new_B3772_ = new_B3753_ & new_B3763_;
  assign new_B3771_ = ~new_B3753_ | new_B3763_;
  assign new_B3770_ = new_B3737_ & ~new_B3738_;
  assign new_B3769_ = ~new_B3737_ & new_B3738_;
  assign new_B3768_ = new_B3790_ & ~new_B3791_;
  assign new_B3767_ = ~new_B3790_ & new_B3791_;
  assign new_B3766_ = ~new_B3789_ | ~new_B3788_;
  assign new_B3765_ = new_B3781_ | new_B3780_;
  assign new_B3764_ = new_B3787_ | new_B3786_;
  assign new_B3763_ = new_B3777_ | new_B3779_;
  assign new_B3762_ = ~new_B3784_ | ~new_B3785_;
  assign new_B3761_ = new_B3737_ & ~new_B3738_;
  assign new_B3760_ = new_B3751_ & ~new_B3763_;
  assign new_B3759_ = ~new_B3751_ & new_B3763_;
  assign new_B3758_ = ~new_B3749_ & new_B3775_;
  assign new_B3757_ = new_B3773_ | new_B3772_;
  assign new_B3756_ = new_B3770_ | new_B3769_;
  assign new_B3755_ = new_B3738_ | new_B3771_;
  assign new_B3754_ = new_B3763_ & new_B3766_;
  assign new_B3753_ = new_B3768_ | new_B3767_;
  assign new_B3752_ = new_B3763_ & new_B3762_;
  assign new_B3751_ = new_B3765_ & new_B3764_;
  assign new_B3750_ = new_B3760_ | new_B3759_;
  assign new_B3749_ = new_B3738_ | new_B3761_;
  assign B3748 = new_B3749_ | new_B3758_;
  assign B3747 = new_B3756_ & new_B3757_;
  assign B3746 = new_B3756_ & new_B3755_;
  assign B3745 = new_B3754_ | new_B3753_;
  assign B3744 = new_B3752_ | new_B3751_;
  assign B3743 = new_B3750_ & new_B3749_;
  assign new_B3742_ = new_C8084_;
  assign new_B3741_ = new_C8017_;
  assign new_B3740_ = new_C7950_;
  assign new_B3739_ = new_C7883_;
  assign new_B3738_ = new_C7816_;
  assign new_B3737_ = new_C7749_;
  assign new_B3736_ = ~new_B3675_ & new_B3689_;
  assign new_B3735_ = new_B3675_ & ~new_B3689_;
  assign new_B3734_ = new_B3675_ & ~new_B3689_;
  assign new_B3733_ = ~new_B3675_ & ~new_B3689_;
  assign new_B3732_ = new_B3675_ & new_B3689_;
  assign new_B3731_ = new_B3735_ | new_B3736_;
  assign new_B3730_ = ~new_B3675_ & new_B3689_;
  assign new_B3729_ = new_B3733_ | new_B3734_;
  assign new_B3728_ = ~new_B3704_ & ~new_B3724_;
  assign new_B3727_ = new_B3704_ & new_B3724_;
  assign new_B3726_ = ~new_B3671_ | ~new_B3696_;
  assign new_B3725_ = new_B3689_ & new_B3726_;
  assign new_B3724_ = new_B3672_ | new_B3673_;
  assign new_B3723_ = new_B3672_ | new_B3689_;
  assign new_B3722_ = ~new_B3689_ & ~new_B3725_;
  assign new_B3721_ = new_B3689_ | new_B3726_;
  assign new_B3720_ = new_B3672_ & ~new_B3673_;
  assign new_B3719_ = ~new_B3672_ & new_B3673_;
  assign new_B3718_ = new_B3682_ | new_B3715_;
  assign new_B3717_ = ~new_B3682_ & ~new_B3716_;
  assign new_B3716_ = new_B3682_ & new_B3715_;
  assign new_B3715_ = ~new_B3671_ | ~new_B3696_;
  assign new_B3714_ = ~new_B3672_ & new_B3682_;
  assign new_B3713_ = new_B3672_ & ~new_B3682_;
  assign new_B3712_ = new_B3674_ & new_B3711_;
  assign new_B3711_ = new_B3730_ | new_B3729_;
  assign new_B3710_ = ~new_B3674_ & new_B3709_;
  assign new_B3709_ = new_B3732_ | new_B3731_;
  assign new_B3708_ = new_B3674_ | new_B3707_;
  assign new_B3707_ = new_B3728_ | new_B3727_;
  assign new_B3706_ = ~new_B3686_ & ~new_B3696_;
  assign new_B3705_ = new_B3686_ & new_B3696_;
  assign new_B3704_ = ~new_B3686_ | new_B3696_;
  assign new_B3703_ = new_B3670_ & ~new_B3671_;
  assign new_B3702_ = ~new_B3670_ & new_B3671_;
  assign new_B3701_ = new_B3723_ & ~new_B3724_;
  assign new_B3700_ = ~new_B3723_ & new_B3724_;
  assign new_B3699_ = ~new_B3722_ | ~new_B3721_;
  assign new_B3698_ = new_B3714_ | new_B3713_;
  assign new_B3697_ = new_B3720_ | new_B3719_;
  assign new_B3696_ = new_B3710_ | new_B3712_;
  assign new_B3695_ = ~new_B3717_ | ~new_B3718_;
  assign new_B3694_ = new_B3670_ & ~new_B3671_;
  assign new_B3693_ = new_B3684_ & ~new_B3696_;
  assign new_B3692_ = ~new_B3684_ & new_B3696_;
  assign new_B3691_ = ~new_B3682_ & new_B3708_;
  assign new_B3690_ = new_B3706_ | new_B3705_;
  assign new_B3689_ = new_B3703_ | new_B3702_;
  assign new_B3688_ = new_B3671_ | new_B3704_;
  assign new_B3687_ = new_B3696_ & new_B3699_;
  assign new_B3686_ = new_B3701_ | new_B3700_;
  assign new_B3685_ = new_B3696_ & new_B3695_;
  assign new_B3684_ = new_B3698_ & new_B3697_;
  assign new_B3683_ = new_B3693_ | new_B3692_;
  assign new_B3682_ = new_B3671_ | new_B3694_;
  assign B3681 = new_B3682_ | new_B3691_;
  assign B3680 = new_B3689_ & new_B3690_;
  assign B3679 = new_B3689_ & new_B3688_;
  assign B3678 = new_B3687_ | new_B3686_;
  assign B3677 = new_B3685_ | new_B3684_;
  assign B3676 = new_B3683_ & new_B3682_;
  assign new_B3675_ = new_C7682_;
  assign new_B3674_ = new_C7615_;
  assign new_B3673_ = new_C7548_;
  assign new_B3672_ = new_C7481_;
  assign new_B3671_ = new_C7414_;
  assign new_B3670_ = new_C7347_;
  assign new_B3669_ = ~new_B3608_ & new_B3622_;
  assign new_B3668_ = new_B3608_ & ~new_B3622_;
  assign new_B3667_ = new_B3608_ & ~new_B3622_;
  assign new_B3666_ = ~new_B3608_ & ~new_B3622_;
  assign new_B3665_ = new_B3608_ & new_B3622_;
  assign new_B3664_ = new_B3668_ | new_B3669_;
  assign new_B3663_ = ~new_B3608_ & new_B3622_;
  assign new_B3662_ = new_B3666_ | new_B3667_;
  assign new_B3661_ = ~new_B3637_ & ~new_B3657_;
  assign new_B3660_ = new_B3637_ & new_B3657_;
  assign new_B3659_ = ~new_B3604_ | ~new_B3629_;
  assign new_B3658_ = new_B3622_ & new_B3659_;
  assign new_B3657_ = new_B3605_ | new_B3606_;
  assign new_B3656_ = new_B3605_ | new_B3622_;
  assign new_B3655_ = ~new_B3622_ & ~new_B3658_;
  assign new_B3654_ = new_B3622_ | new_B3659_;
  assign new_B3653_ = new_B3605_ & ~new_B3606_;
  assign new_B3652_ = ~new_B3605_ & new_B3606_;
  assign new_B3651_ = new_B3615_ | new_B3648_;
  assign new_B3650_ = ~new_B3615_ & ~new_B3649_;
  assign new_B3649_ = new_B3615_ & new_B3648_;
  assign new_B3648_ = ~new_B3604_ | ~new_B3629_;
  assign new_B3647_ = ~new_B3605_ & new_B3615_;
  assign new_B3646_ = new_B3605_ & ~new_B3615_;
  assign new_B3645_ = new_B3607_ & new_B3644_;
  assign new_B3644_ = new_B3663_ | new_B3662_;
  assign new_B3643_ = ~new_B3607_ & new_B3642_;
  assign new_B3642_ = new_B3665_ | new_B3664_;
  assign new_B3641_ = new_B3607_ | new_B3640_;
  assign new_B3640_ = new_B3661_ | new_B3660_;
  assign new_B3639_ = ~new_B3619_ & ~new_B3629_;
  assign new_B3638_ = new_B3619_ & new_B3629_;
  assign new_B3637_ = ~new_B3619_ | new_B3629_;
  assign new_B3636_ = new_B3603_ & ~new_B3604_;
  assign new_B3635_ = ~new_B3603_ & new_B3604_;
  assign new_B3634_ = new_B3656_ & ~new_B3657_;
  assign new_B3633_ = ~new_B3656_ & new_B3657_;
  assign new_B3632_ = ~new_B3655_ | ~new_B3654_;
  assign new_B3631_ = new_B3647_ | new_B3646_;
  assign new_B3630_ = new_B3653_ | new_B3652_;
  assign new_B3629_ = new_B3643_ | new_B3645_;
  assign new_B3628_ = ~new_B3650_ | ~new_B3651_;
  assign new_B3627_ = new_B3603_ & ~new_B3604_;
  assign new_B3626_ = new_B3617_ & ~new_B3629_;
  assign new_B3625_ = ~new_B3617_ & new_B3629_;
  assign new_B3624_ = ~new_B3615_ & new_B3641_;
  assign new_B3623_ = new_B3639_ | new_B3638_;
  assign new_B3622_ = new_B3636_ | new_B3635_;
  assign new_B3621_ = new_B3604_ | new_B3637_;
  assign new_B3620_ = new_B3629_ & new_B3632_;
  assign new_B3619_ = new_B3634_ | new_B3633_;
  assign new_B3618_ = new_B3629_ & new_B3628_;
  assign new_B3617_ = new_B3631_ & new_B3630_;
  assign new_B3616_ = new_B3626_ | new_B3625_;
  assign new_B3615_ = new_B3604_ | new_B3627_;
  assign B3614 = new_B3615_ | new_B3624_;
  assign B3613 = new_B3622_ & new_B3623_;
  assign B3612 = new_B3622_ & new_B3621_;
  assign B3611 = new_B3620_ | new_B3619_;
  assign B3610 = new_B3618_ | new_B3617_;
  assign B3609 = new_B3616_ & new_B3615_;
  assign new_B3608_ = new_C7280_;
  assign new_B3607_ = new_C7213_;
  assign new_B3606_ = new_C7146_;
  assign new_B3605_ = new_C7079_;
  assign new_B3604_ = new_C7012_;
  assign new_B3603_ = new_C6945_;
  assign new_B3602_ = ~new_B3541_ & new_B3555_;
  assign new_B3601_ = new_B3541_ & ~new_B3555_;
  assign new_B3600_ = new_B3541_ & ~new_B3555_;
  assign new_B3599_ = ~new_B3541_ & ~new_B3555_;
  assign new_B3598_ = new_B3541_ & new_B3555_;
  assign new_B3597_ = new_B3601_ | new_B3602_;
  assign new_B3596_ = ~new_B3541_ & new_B3555_;
  assign new_B3595_ = new_B3599_ | new_B3600_;
  assign new_B3594_ = ~new_B3570_ & ~new_B3590_;
  assign new_B3593_ = new_B3570_ & new_B3590_;
  assign new_B3592_ = ~new_B3537_ | ~new_B3562_;
  assign new_B3591_ = new_B3555_ & new_B3592_;
  assign new_B3590_ = new_B3538_ | new_B3539_;
  assign new_B3589_ = new_B3538_ | new_B3555_;
  assign new_B3588_ = ~new_B3555_ & ~new_B3591_;
  assign new_B3587_ = new_B3555_ | new_B3592_;
  assign new_B3586_ = new_B3538_ & ~new_B3539_;
  assign new_B3585_ = ~new_B3538_ & new_B3539_;
  assign new_B3584_ = new_B3548_ | new_B3581_;
  assign new_B3583_ = ~new_B3548_ & ~new_B3582_;
  assign new_B3582_ = new_B3548_ & new_B3581_;
  assign new_B3581_ = ~new_B3537_ | ~new_B3562_;
  assign new_B3580_ = ~new_B3538_ & new_B3548_;
  assign new_B3579_ = new_B3538_ & ~new_B3548_;
  assign new_B3578_ = new_B3540_ & new_B3577_;
  assign new_B3577_ = new_B3596_ | new_B3595_;
  assign new_B3576_ = ~new_B3540_ & new_B3575_;
  assign new_B3575_ = new_B3598_ | new_B3597_;
  assign new_B3574_ = new_B3540_ | new_B3573_;
  assign new_B3573_ = new_B3594_ | new_B3593_;
  assign new_B3572_ = ~new_B3552_ & ~new_B3562_;
  assign new_B3571_ = new_B3552_ & new_B3562_;
  assign new_B3570_ = ~new_B3552_ | new_B3562_;
  assign new_B3569_ = new_B3536_ & ~new_B3537_;
  assign new_B3568_ = ~new_B3536_ & new_B3537_;
  assign new_B3567_ = new_B3589_ & ~new_B3590_;
  assign new_B3566_ = ~new_B3589_ & new_B3590_;
  assign new_B3565_ = ~new_B3588_ | ~new_B3587_;
  assign new_B3564_ = new_B3580_ | new_B3579_;
  assign new_B3563_ = new_B3586_ | new_B3585_;
  assign new_B3562_ = new_B3576_ | new_B3578_;
  assign new_B3561_ = ~new_B3583_ | ~new_B3584_;
  assign new_B3560_ = new_B3536_ & ~new_B3537_;
  assign new_B3559_ = new_B3550_ & ~new_B3562_;
  assign new_B3558_ = ~new_B3550_ & new_B3562_;
  assign new_B3557_ = ~new_B3548_ & new_B3574_;
  assign new_B3556_ = new_B3572_ | new_B3571_;
  assign new_B3555_ = new_B3569_ | new_B3568_;
  assign new_B3554_ = new_B3537_ | new_B3570_;
  assign new_B3553_ = new_B3562_ & new_B3565_;
  assign new_B3552_ = new_B3567_ | new_B3566_;
  assign new_B3551_ = new_B3562_ & new_B3561_;
  assign new_B3550_ = new_B3564_ & new_B3563_;
  assign new_B3549_ = new_B3559_ | new_B3558_;
  assign new_B3548_ = new_B3537_ | new_B3560_;
  assign B3547 = new_B3548_ | new_B3557_;
  assign B3546 = new_B3555_ & new_B3556_;
  assign B3545 = new_B3555_ & new_B3554_;
  assign B3544 = new_B3553_ | new_B3552_;
  assign B3543 = new_B3551_ | new_B3550_;
  assign B3542 = new_B3549_ & new_B3548_;
  assign new_B3541_ = new_C6878_;
  assign new_B3540_ = new_C6811_;
  assign new_B3539_ = new_C6744_;
  assign new_B3538_ = new_C6677_;
  assign new_B3537_ = new_C6610_;
  assign new_B3536_ = new_C6543_;
  assign new_B3535_ = ~new_B3474_ & new_B3488_;
  assign new_B3534_ = new_B3474_ & ~new_B3488_;
  assign new_B3533_ = new_B3474_ & ~new_B3488_;
  assign new_B3532_ = ~new_B3474_ & ~new_B3488_;
  assign new_B3531_ = new_B3474_ & new_B3488_;
  assign new_B3530_ = new_B3534_ | new_B3535_;
  assign new_B3529_ = ~new_B3474_ & new_B3488_;
  assign new_B3528_ = new_B3532_ | new_B3533_;
  assign new_B3527_ = ~new_B3503_ & ~new_B3523_;
  assign new_B3526_ = new_B3503_ & new_B3523_;
  assign new_B3525_ = ~new_B3470_ | ~new_B3495_;
  assign new_B3524_ = new_B3488_ & new_B3525_;
  assign new_B3523_ = new_B3471_ | new_B3472_;
  assign new_B3522_ = new_B3471_ | new_B3488_;
  assign new_B3521_ = ~new_B3488_ & ~new_B3524_;
  assign new_B3520_ = new_B3488_ | new_B3525_;
  assign new_B3519_ = new_B3471_ & ~new_B3472_;
  assign new_B3518_ = ~new_B3471_ & new_B3472_;
  assign new_B3517_ = new_B3481_ | new_B3514_;
  assign new_B3516_ = ~new_B3481_ & ~new_B3515_;
  assign new_B3515_ = new_B3481_ & new_B3514_;
  assign new_B3514_ = ~new_B3470_ | ~new_B3495_;
  assign new_B3513_ = ~new_B3471_ & new_B3481_;
  assign new_B3512_ = new_B3471_ & ~new_B3481_;
  assign new_B3511_ = new_B3473_ & new_B3510_;
  assign new_B3510_ = new_B3529_ | new_B3528_;
  assign new_B3509_ = ~new_B3473_ & new_B3508_;
  assign new_B3508_ = new_B3531_ | new_B3530_;
  assign new_B3507_ = new_B3473_ | new_B3506_;
  assign new_B3506_ = new_B3527_ | new_B3526_;
  assign new_B3505_ = ~new_B3485_ & ~new_B3495_;
  assign new_B3504_ = new_B3485_ & new_B3495_;
  assign new_B3503_ = ~new_B3485_ | new_B3495_;
  assign new_B3502_ = new_B3469_ & ~new_B3470_;
  assign new_B3501_ = ~new_B3469_ & new_B3470_;
  assign new_B3500_ = new_B3522_ & ~new_B3523_;
  assign new_B3499_ = ~new_B3522_ & new_B3523_;
  assign new_B3498_ = ~new_B3521_ | ~new_B3520_;
  assign new_B3497_ = new_B3513_ | new_B3512_;
  assign new_B3496_ = new_B3519_ | new_B3518_;
  assign new_B3495_ = new_B3509_ | new_B3511_;
  assign new_B3494_ = ~new_B3516_ | ~new_B3517_;
  assign new_B3493_ = new_B3469_ & ~new_B3470_;
  assign new_B3492_ = new_B3483_ & ~new_B3495_;
  assign new_B3491_ = ~new_B3483_ & new_B3495_;
  assign new_B3490_ = ~new_B3481_ & new_B3507_;
  assign new_B3489_ = new_B3505_ | new_B3504_;
  assign new_B3488_ = new_B3502_ | new_B3501_;
  assign new_B3487_ = new_B3470_ | new_B3503_;
  assign new_B3486_ = new_B3495_ & new_B3498_;
  assign new_B3485_ = new_B3500_ | new_B3499_;
  assign new_B3484_ = new_B3495_ & new_B3494_;
  assign new_B3483_ = new_B3497_ & new_B3496_;
  assign new_B3482_ = new_B3492_ | new_B3491_;
  assign new_B3481_ = new_B3470_ | new_B3493_;
  assign B3480 = new_B3481_ | new_B3490_;
  assign B3479 = new_B3488_ & new_B3489_;
  assign B3478 = new_B3488_ & new_B3487_;
  assign B3477 = new_B3486_ | new_B3485_;
  assign B3476 = new_B3484_ | new_B3483_;
  assign B3475 = new_B3482_ & new_B3481_;
  assign new_B3474_ = new_C6476_;
  assign new_B3473_ = new_C6409_;
  assign new_B3472_ = new_C6342_;
  assign new_B3471_ = new_C6275_;
  assign new_B3470_ = new_C6208_;
  assign new_B3469_ = new_C6141_;
  assign new_B3468_ = ~new_B3407_ & new_B3421_;
  assign new_B3467_ = new_B3407_ & ~new_B3421_;
  assign new_B3466_ = new_B3407_ & ~new_B3421_;
  assign new_B3465_ = ~new_B3407_ & ~new_B3421_;
  assign new_B3464_ = new_B3407_ & new_B3421_;
  assign new_B3463_ = new_B3467_ | new_B3468_;
  assign new_B3462_ = ~new_B3407_ & new_B3421_;
  assign new_B3461_ = new_B3465_ | new_B3466_;
  assign new_B3460_ = ~new_B3436_ & ~new_B3456_;
  assign new_B3459_ = new_B3436_ & new_B3456_;
  assign new_B3458_ = ~new_B3403_ | ~new_B3428_;
  assign new_B3457_ = new_B3421_ & new_B3458_;
  assign new_B3456_ = new_B3404_ | new_B3405_;
  assign new_B3455_ = new_B3404_ | new_B3421_;
  assign new_B3454_ = ~new_B3421_ & ~new_B3457_;
  assign new_B3453_ = new_B3421_ | new_B3458_;
  assign new_B3452_ = new_B3404_ & ~new_B3405_;
  assign new_B3451_ = ~new_B3404_ & new_B3405_;
  assign new_B3450_ = new_B3414_ | new_B3447_;
  assign new_B3449_ = ~new_B3414_ & ~new_B3448_;
  assign new_B3448_ = new_B3414_ & new_B3447_;
  assign new_B3447_ = ~new_B3403_ | ~new_B3428_;
  assign new_B3446_ = ~new_B3404_ & new_B3414_;
  assign new_B3445_ = new_B3404_ & ~new_B3414_;
  assign new_B3444_ = new_B3406_ & new_B3443_;
  assign new_B3443_ = new_B3462_ | new_B3461_;
  assign new_B3442_ = ~new_B3406_ & new_B3441_;
  assign new_B3441_ = new_B3464_ | new_B3463_;
  assign new_B3440_ = new_B3406_ | new_B3439_;
  assign new_B3439_ = new_B3460_ | new_B3459_;
  assign new_B3438_ = ~new_B3418_ & ~new_B3428_;
  assign new_B3437_ = new_B3418_ & new_B3428_;
  assign new_B3436_ = ~new_B3418_ | new_B3428_;
  assign new_B3435_ = new_B3402_ & ~new_B3403_;
  assign new_B3434_ = ~new_B3402_ & new_B3403_;
  assign new_B3433_ = new_B3455_ & ~new_B3456_;
  assign new_B3432_ = ~new_B3455_ & new_B3456_;
  assign new_B3431_ = ~new_B3454_ | ~new_B3453_;
  assign new_B3430_ = new_B3446_ | new_B3445_;
  assign new_B3429_ = new_B3452_ | new_B3451_;
  assign new_B3428_ = new_B3442_ | new_B3444_;
  assign new_B3427_ = ~new_B3449_ | ~new_B3450_;
  assign new_B3426_ = new_B3402_ & ~new_B3403_;
  assign new_B3425_ = new_B3416_ & ~new_B3428_;
  assign new_B3424_ = ~new_B3416_ & new_B3428_;
  assign new_B3423_ = ~new_B3414_ & new_B3440_;
  assign new_B3422_ = new_B3438_ | new_B3437_;
  assign new_B3421_ = new_B3435_ | new_B3434_;
  assign new_B3420_ = new_B3403_ | new_B3436_;
  assign new_B3419_ = new_B3428_ & new_B3431_;
  assign new_B3418_ = new_B3433_ | new_B3432_;
  assign new_B3417_ = new_B3428_ & new_B3427_;
  assign new_B3416_ = new_B3430_ & new_B3429_;
  assign new_B3415_ = new_B3425_ | new_B3424_;
  assign new_B3414_ = new_B3403_ | new_B3426_;
  assign B3413 = new_B3414_ | new_B3423_;
  assign B3412 = new_B3421_ & new_B3422_;
  assign B3411 = new_B3421_ & new_B3420_;
  assign B3410 = new_B3419_ | new_B3418_;
  assign B3409 = new_B3417_ | new_B3416_;
  assign B3408 = new_B3415_ & new_B3414_;
  assign new_B3407_ = new_C6074_;
  assign new_B3406_ = new_C6007_;
  assign new_B3405_ = new_C5940_;
  assign new_B3404_ = new_C5873_;
  assign new_B3403_ = new_C5806_;
  assign new_B3402_ = new_C5739_;
  assign new_B3401_ = ~new_B3340_ & new_B3354_;
  assign new_B3400_ = new_B3340_ & ~new_B3354_;
  assign new_B3399_ = new_B3340_ & ~new_B3354_;
  assign new_B3398_ = ~new_B3340_ & ~new_B3354_;
  assign new_B3397_ = new_B3340_ & new_B3354_;
  assign new_B3396_ = new_B3400_ | new_B3401_;
  assign new_B3395_ = ~new_B3340_ & new_B3354_;
  assign new_B3394_ = new_B3398_ | new_B3399_;
  assign new_B3393_ = ~new_B3369_ & ~new_B3389_;
  assign new_B3392_ = new_B3369_ & new_B3389_;
  assign new_B3391_ = ~new_B3336_ | ~new_B3361_;
  assign new_B3390_ = new_B3354_ & new_B3391_;
  assign new_B3389_ = new_B3337_ | new_B3338_;
  assign new_B3388_ = new_B3337_ | new_B3354_;
  assign new_B3387_ = ~new_B3354_ & ~new_B3390_;
  assign new_B3386_ = new_B3354_ | new_B3391_;
  assign new_B3385_ = new_B3337_ & ~new_B3338_;
  assign new_B3384_ = ~new_B3337_ & new_B3338_;
  assign new_B3383_ = new_B3347_ | new_B3380_;
  assign new_B3382_ = ~new_B3347_ & ~new_B3381_;
  assign new_B3381_ = new_B3347_ & new_B3380_;
  assign new_B3380_ = ~new_B3336_ | ~new_B3361_;
  assign new_B3379_ = ~new_B3337_ & new_B3347_;
  assign new_B3378_ = new_B3337_ & ~new_B3347_;
  assign new_B3377_ = new_B3339_ & new_B3376_;
  assign new_B3376_ = new_B3395_ | new_B3394_;
  assign new_B3375_ = ~new_B3339_ & new_B3374_;
  assign new_B3374_ = new_B3397_ | new_B3396_;
  assign new_B3373_ = new_B3339_ | new_B3372_;
  assign new_B3372_ = new_B3393_ | new_B3392_;
  assign new_B3371_ = ~new_B3351_ & ~new_B3361_;
  assign new_B3370_ = new_B3351_ & new_B3361_;
  assign new_B3369_ = ~new_B3351_ | new_B3361_;
  assign new_B3368_ = new_B3335_ & ~new_B3336_;
  assign new_B3367_ = ~new_B3335_ & new_B3336_;
  assign new_B3366_ = new_B3388_ & ~new_B3389_;
  assign new_B3365_ = ~new_B3388_ & new_B3389_;
  assign new_B3364_ = ~new_B3387_ | ~new_B3386_;
  assign new_B3363_ = new_B3379_ | new_B3378_;
  assign new_B3362_ = new_B3385_ | new_B3384_;
  assign new_B3361_ = new_B3375_ | new_B3377_;
  assign new_B3360_ = ~new_B3382_ | ~new_B3383_;
  assign new_B3359_ = new_B3335_ & ~new_B3336_;
  assign new_B3358_ = new_B3349_ & ~new_B3361_;
  assign new_B3357_ = ~new_B3349_ & new_B3361_;
  assign new_B3356_ = ~new_B3347_ & new_B3373_;
  assign new_B3355_ = new_B3371_ | new_B3370_;
  assign new_B3354_ = new_B3368_ | new_B3367_;
  assign new_B3353_ = new_B3336_ | new_B3369_;
  assign new_B3352_ = new_B3361_ & new_B3364_;
  assign new_B3351_ = new_B3366_ | new_B3365_;
  assign new_B3350_ = new_B3361_ & new_B3360_;
  assign new_B3349_ = new_B3363_ & new_B3362_;
  assign new_B3348_ = new_B3358_ | new_B3357_;
  assign new_B3347_ = new_B3336_ | new_B3359_;
  assign B3346 = new_B3347_ | new_B3356_;
  assign B3345 = new_B3354_ & new_B3355_;
  assign B3344 = new_B3354_ & new_B3353_;
  assign B3343 = new_B3352_ | new_B3351_;
  assign B3342 = new_B3350_ | new_B3349_;
  assign B3341 = new_B3348_ & new_B3347_;
  assign new_B3340_ = new_C5672_;
  assign new_B3339_ = new_C5605_;
  assign new_B3338_ = new_C5538_;
  assign new_B3337_ = new_C5471_;
  assign new_B3336_ = new_C5404_;
  assign new_B3335_ = new_C5337_;
  assign new_B3334_ = ~new_B3273_ & new_B3287_;
  assign new_B3333_ = new_B3273_ & ~new_B3287_;
  assign new_B3332_ = new_B3273_ & ~new_B3287_;
  assign new_B3331_ = ~new_B3273_ & ~new_B3287_;
  assign new_B3330_ = new_B3273_ & new_B3287_;
  assign new_B3329_ = new_B3333_ | new_B3334_;
  assign new_B3328_ = ~new_B3273_ & new_B3287_;
  assign new_B3327_ = new_B3331_ | new_B3332_;
  assign new_B3326_ = ~new_B3302_ & ~new_B3322_;
  assign new_B3325_ = new_B3302_ & new_B3322_;
  assign new_B3324_ = ~new_B3269_ | ~new_B3294_;
  assign new_B3323_ = new_B3287_ & new_B3324_;
  assign new_B3322_ = new_B3270_ | new_B3271_;
  assign new_B3321_ = new_B3270_ | new_B3287_;
  assign new_B3320_ = ~new_B3287_ & ~new_B3323_;
  assign new_B3319_ = new_B3287_ | new_B3324_;
  assign new_B3318_ = new_B3270_ & ~new_B3271_;
  assign new_B3317_ = ~new_B3270_ & new_B3271_;
  assign new_B3316_ = new_B3280_ | new_B3313_;
  assign new_B3315_ = ~new_B3280_ & ~new_B3314_;
  assign new_B3314_ = new_B3280_ & new_B3313_;
  assign new_B3313_ = ~new_B3269_ | ~new_B3294_;
  assign new_B3312_ = ~new_B3270_ & new_B3280_;
  assign new_B3311_ = new_B3270_ & ~new_B3280_;
  assign new_B3310_ = new_B3272_ & new_B3309_;
  assign new_B3309_ = new_B3328_ | new_B3327_;
  assign new_B3308_ = ~new_B3272_ & new_B3307_;
  assign new_B3307_ = new_B3330_ | new_B3329_;
  assign new_B3306_ = new_B3272_ | new_B3305_;
  assign new_B3305_ = new_B3326_ | new_B3325_;
  assign new_B3304_ = ~new_B3284_ & ~new_B3294_;
  assign new_B3303_ = new_B3284_ & new_B3294_;
  assign new_B3302_ = ~new_B3284_ | new_B3294_;
  assign new_B3301_ = new_B3268_ & ~new_B3269_;
  assign new_B3300_ = ~new_B3268_ & new_B3269_;
  assign new_B3299_ = new_B3321_ & ~new_B3322_;
  assign new_B3298_ = ~new_B3321_ & new_B3322_;
  assign new_B3297_ = ~new_B3320_ | ~new_B3319_;
  assign new_B3296_ = new_B3312_ | new_B3311_;
  assign new_B3295_ = new_B3318_ | new_B3317_;
  assign new_B3294_ = new_B3308_ | new_B3310_;
  assign new_B3293_ = ~new_B3315_ | ~new_B3316_;
  assign new_B3292_ = new_B3268_ & ~new_B3269_;
  assign new_B3291_ = new_B3282_ & ~new_B3294_;
  assign new_B3290_ = ~new_B3282_ & new_B3294_;
  assign new_B3289_ = ~new_B3280_ & new_B3306_;
  assign new_B3288_ = new_B3304_ | new_B3303_;
  assign new_B3287_ = new_B3301_ | new_B3300_;
  assign new_B3286_ = new_B3269_ | new_B3302_;
  assign new_B3285_ = new_B3294_ & new_B3297_;
  assign new_B3284_ = new_B3299_ | new_B3298_;
  assign new_B3283_ = new_B3294_ & new_B3293_;
  assign new_B3282_ = new_B3296_ & new_B3295_;
  assign new_B3281_ = new_B3291_ | new_B3290_;
  assign new_B3280_ = new_B3269_ | new_B3292_;
  assign B3279 = new_B3280_ | new_B3289_;
  assign B3278 = new_B3287_ & new_B3288_;
  assign B3277 = new_B3287_ & new_B3286_;
  assign B3276 = new_B3285_ | new_B3284_;
  assign B3275 = new_B3283_ | new_B3282_;
  assign B3274 = new_B3281_ & new_B3280_;
  assign new_B3273_ = new_C5270_;
  assign new_B3272_ = new_C5203_;
  assign new_B3271_ = new_C5136_;
  assign new_B3270_ = new_C5069_;
  assign new_B3269_ = new_C5002_;
  assign new_B3268_ = new_C4935_;
  assign new_B3267_ = ~new_B3206_ & new_B3220_;
  assign new_B3266_ = new_B3206_ & ~new_B3220_;
  assign new_B3265_ = new_B3206_ & ~new_B3220_;
  assign new_B3264_ = ~new_B3206_ & ~new_B3220_;
  assign new_B3263_ = new_B3206_ & new_B3220_;
  assign new_B3262_ = new_B3266_ | new_B3267_;
  assign new_B3261_ = ~new_B3206_ & new_B3220_;
  assign new_B3260_ = new_B3264_ | new_B3265_;
  assign new_B3259_ = ~new_B3235_ & ~new_B3255_;
  assign new_B3258_ = new_B3235_ & new_B3255_;
  assign new_B3257_ = ~new_B3202_ | ~new_B3227_;
  assign new_B3256_ = new_B3220_ & new_B3257_;
  assign new_B3255_ = new_B3203_ | new_B3204_;
  assign new_B3254_ = new_B3203_ | new_B3220_;
  assign new_B3253_ = ~new_B3220_ & ~new_B3256_;
  assign new_B3252_ = new_B3220_ | new_B3257_;
  assign new_B3251_ = new_B3203_ & ~new_B3204_;
  assign new_B3250_ = ~new_B3203_ & new_B3204_;
  assign new_B3249_ = new_B3213_ | new_B3246_;
  assign new_B3248_ = ~new_B3213_ & ~new_B3247_;
  assign new_B3247_ = new_B3213_ & new_B3246_;
  assign new_B3246_ = ~new_B3202_ | ~new_B3227_;
  assign new_B3245_ = ~new_B3203_ & new_B3213_;
  assign new_B3244_ = new_B3203_ & ~new_B3213_;
  assign new_B3243_ = new_B3205_ & new_B3242_;
  assign new_B3242_ = new_B3261_ | new_B3260_;
  assign new_B3241_ = ~new_B3205_ & new_B3240_;
  assign new_B3240_ = new_B3263_ | new_B3262_;
  assign new_B3239_ = new_B3205_ | new_B3238_;
  assign new_B3238_ = new_B3259_ | new_B3258_;
  assign new_B3237_ = ~new_B3217_ & ~new_B3227_;
  assign new_B3236_ = new_B3217_ & new_B3227_;
  assign new_B3235_ = ~new_B3217_ | new_B3227_;
  assign new_B3234_ = new_B3201_ & ~new_B3202_;
  assign new_B3233_ = ~new_B3201_ & new_B3202_;
  assign new_B3232_ = new_B3254_ & ~new_B3255_;
  assign new_B3231_ = ~new_B3254_ & new_B3255_;
  assign new_B3230_ = ~new_B3253_ | ~new_B3252_;
  assign new_B3229_ = new_B3245_ | new_B3244_;
  assign new_B3228_ = new_B3251_ | new_B3250_;
  assign new_B3227_ = new_B3241_ | new_B3243_;
  assign new_B3226_ = ~new_B3248_ | ~new_B3249_;
  assign new_B3225_ = new_B3201_ & ~new_B3202_;
  assign new_B3224_ = new_B3215_ & ~new_B3227_;
  assign new_B3223_ = ~new_B3215_ & new_B3227_;
  assign new_B3222_ = ~new_B3213_ & new_B3239_;
  assign new_B3221_ = new_B3237_ | new_B3236_;
  assign new_B3220_ = new_B3234_ | new_B3233_;
  assign new_B3219_ = new_B3202_ | new_B3235_;
  assign new_B3218_ = new_B3227_ & new_B3230_;
  assign new_B3217_ = new_B3232_ | new_B3231_;
  assign new_B3216_ = new_B3227_ & new_B3226_;
  assign new_B3215_ = new_B3229_ & new_B3228_;
  assign new_B3214_ = new_B3224_ | new_B3223_;
  assign new_B3213_ = new_B3202_ | new_B3225_;
  assign B3212 = new_B3213_ | new_B3222_;
  assign B3211 = new_B3220_ & new_B3221_;
  assign B3210 = new_B3220_ & new_B3219_;
  assign B3209 = new_B3218_ | new_B3217_;
  assign B3208 = new_B3216_ | new_B3215_;
  assign B3207 = new_B3214_ & new_B3213_;
  assign new_B3206_ = new_C4868_;
  assign new_B3205_ = new_C4801_;
  assign new_B3204_ = new_C4734_;
  assign new_B3203_ = new_C4667_;
  assign new_B3202_ = new_C4600_;
  assign new_B3201_ = new_C4533_;
  assign new_B3200_ = ~new_B3139_ & new_B3153_;
  assign new_B3199_ = new_B3139_ & ~new_B3153_;
  assign new_B3198_ = new_B3139_ & ~new_B3153_;
  assign new_B3197_ = ~new_B3139_ & ~new_B3153_;
  assign new_B3196_ = new_B3139_ & new_B3153_;
  assign new_B3195_ = new_B3199_ | new_B3200_;
  assign new_B3194_ = ~new_B3139_ & new_B3153_;
  assign new_B3193_ = new_B3197_ | new_B3198_;
  assign new_B3192_ = ~new_B3168_ & ~new_B3188_;
  assign new_B3191_ = new_B3168_ & new_B3188_;
  assign new_B3190_ = ~new_B3135_ | ~new_B3160_;
  assign new_B3189_ = new_B3153_ & new_B3190_;
  assign new_B3188_ = new_B3136_ | new_B3137_;
  assign new_B3187_ = new_B3136_ | new_B3153_;
  assign new_B3186_ = ~new_B3153_ & ~new_B3189_;
  assign new_B3185_ = new_B3153_ | new_B3190_;
  assign new_B3184_ = new_B3136_ & ~new_B3137_;
  assign new_B3183_ = ~new_B3136_ & new_B3137_;
  assign new_B3182_ = new_B3146_ | new_B3179_;
  assign new_B3181_ = ~new_B3146_ & ~new_B3180_;
  assign new_B3180_ = new_B3146_ & new_B3179_;
  assign new_B3179_ = ~new_B3135_ | ~new_B3160_;
  assign new_B3178_ = ~new_B3136_ & new_B3146_;
  assign new_B3177_ = new_B3136_ & ~new_B3146_;
  assign new_B3176_ = new_B3138_ & new_B3175_;
  assign new_B3175_ = new_B3194_ | new_B3193_;
  assign new_B3174_ = ~new_B3138_ & new_B3173_;
  assign new_B3173_ = new_B3196_ | new_B3195_;
  assign new_B3172_ = new_B3138_ | new_B3171_;
  assign new_B3171_ = new_B3192_ | new_B3191_;
  assign new_B3170_ = ~new_B3150_ & ~new_B3160_;
  assign new_B3169_ = new_B3150_ & new_B3160_;
  assign new_B3168_ = ~new_B3150_ | new_B3160_;
  assign new_B3167_ = new_B3134_ & ~new_B3135_;
  assign new_B3166_ = ~new_B3134_ & new_B3135_;
  assign new_B3165_ = new_B3187_ & ~new_B3188_;
  assign new_B3164_ = ~new_B3187_ & new_B3188_;
  assign new_B3163_ = ~new_B3186_ | ~new_B3185_;
  assign new_B3162_ = new_B3178_ | new_B3177_;
  assign new_B3161_ = new_B3184_ | new_B3183_;
  assign new_B3160_ = new_B3174_ | new_B3176_;
  assign new_B3159_ = ~new_B3181_ | ~new_B3182_;
  assign new_B3158_ = new_B3134_ & ~new_B3135_;
  assign new_B3157_ = new_B3148_ & ~new_B3160_;
  assign new_B3156_ = ~new_B3148_ & new_B3160_;
  assign new_B3155_ = ~new_B3146_ & new_B3172_;
  assign new_B3154_ = new_B3170_ | new_B3169_;
  assign new_B3153_ = new_B3167_ | new_B3166_;
  assign new_B3152_ = new_B3135_ | new_B3168_;
  assign new_B3151_ = new_B3160_ & new_B3163_;
  assign new_B3150_ = new_B3165_ | new_B3164_;
  assign new_B3149_ = new_B3160_ & new_B3159_;
  assign new_B3148_ = new_B3162_ & new_B3161_;
  assign new_B3147_ = new_B3157_ | new_B3156_;
  assign new_B3146_ = new_B3135_ | new_B3158_;
  assign B3145 = new_B3146_ | new_B3155_;
  assign B3144 = new_B3153_ & new_B3154_;
  assign B3143 = new_B3153_ & new_B3152_;
  assign B3142 = new_B3151_ | new_B3150_;
  assign B3141 = new_B3149_ | new_B3148_;
  assign B3140 = new_B3147_ & new_B3146_;
  assign new_B3139_ = new_C4466_;
  assign new_B3138_ = new_C4399_;
  assign new_B3137_ = new_C4332_;
  assign new_B3136_ = new_C4265_;
  assign new_B3135_ = new_C4198_;
  assign new_B3134_ = new_C4131_;
  assign new_B3133_ = ~new_B3072_ & new_B3086_;
  assign new_B3132_ = new_B3072_ & ~new_B3086_;
  assign new_B3131_ = new_B3072_ & ~new_B3086_;
  assign new_B3130_ = ~new_B3072_ & ~new_B3086_;
  assign new_B3129_ = new_B3072_ & new_B3086_;
  assign new_B3128_ = new_B3132_ | new_B3133_;
  assign new_B3127_ = ~new_B3072_ & new_B3086_;
  assign new_B3126_ = new_B3130_ | new_B3131_;
  assign new_B3125_ = ~new_B3101_ & ~new_B3121_;
  assign new_B3124_ = new_B3101_ & new_B3121_;
  assign new_B3123_ = ~new_B3068_ | ~new_B3093_;
  assign new_B3122_ = new_B3086_ & new_B3123_;
  assign new_B3121_ = new_B3069_ | new_B3070_;
  assign new_B3120_ = new_B3069_ | new_B3086_;
  assign new_B3119_ = ~new_B3086_ & ~new_B3122_;
  assign new_B3118_ = new_B3086_ | new_B3123_;
  assign new_B3117_ = new_B3069_ & ~new_B3070_;
  assign new_B3116_ = ~new_B3069_ & new_B3070_;
  assign new_B3115_ = new_B3079_ | new_B3112_;
  assign new_B3114_ = ~new_B3079_ & ~new_B3113_;
  assign new_B3113_ = new_B3079_ & new_B3112_;
  assign new_B3112_ = ~new_B3068_ | ~new_B3093_;
  assign new_B3111_ = ~new_B3069_ & new_B3079_;
  assign new_B3110_ = new_B3069_ & ~new_B3079_;
  assign new_B3109_ = new_B3071_ & new_B3108_;
  assign new_B3108_ = new_B3127_ | new_B3126_;
  assign new_B3107_ = ~new_B3071_ & new_B3106_;
  assign new_B3106_ = new_B3129_ | new_B3128_;
  assign new_B3105_ = new_B3071_ | new_B3104_;
  assign new_B3104_ = new_B3125_ | new_B3124_;
  assign new_B3103_ = ~new_B3083_ & ~new_B3093_;
  assign new_B3102_ = new_B3083_ & new_B3093_;
  assign new_B3101_ = ~new_B3083_ | new_B3093_;
  assign new_B3100_ = new_B3067_ & ~new_B3068_;
  assign new_B3099_ = ~new_B3067_ & new_B3068_;
  assign new_B3098_ = new_B3120_ & ~new_B3121_;
  assign new_B3097_ = ~new_B3120_ & new_B3121_;
  assign new_B3096_ = ~new_B3119_ | ~new_B3118_;
  assign new_B3095_ = new_B3111_ | new_B3110_;
  assign new_B3094_ = new_B3117_ | new_B3116_;
  assign new_B3093_ = new_B3107_ | new_B3109_;
  assign new_B3092_ = ~new_B3114_ | ~new_B3115_;
  assign new_B3091_ = new_B3067_ & ~new_B3068_;
  assign new_B3090_ = new_B3081_ & ~new_B3093_;
  assign new_B3089_ = ~new_B3081_ & new_B3093_;
  assign new_B3088_ = ~new_B3079_ & new_B3105_;
  assign new_B3087_ = new_B3103_ | new_B3102_;
  assign new_B3086_ = new_B3100_ | new_B3099_;
  assign new_B3085_ = new_B3068_ | new_B3101_;
  assign new_B3084_ = new_B3093_ & new_B3096_;
  assign new_B3083_ = new_B3098_ | new_B3097_;
  assign new_B3082_ = new_B3093_ & new_B3092_;
  assign new_B3081_ = new_B3095_ & new_B3094_;
  assign new_B3080_ = new_B3090_ | new_B3089_;
  assign new_B3079_ = new_B3068_ | new_B3091_;
  assign B3078 = new_B3079_ | new_B3088_;
  assign B3077 = new_B3086_ & new_B3087_;
  assign B3076 = new_B3086_ & new_B3085_;
  assign B3075 = new_B3084_ | new_B3083_;
  assign B3074 = new_B3082_ | new_B3081_;
  assign B3073 = new_B3080_ & new_B3079_;
  assign new_B3072_ = new_C4064_;
  assign new_B3071_ = new_C3997_;
  assign new_B3070_ = new_C3930_;
  assign new_B3069_ = new_C3863_;
  assign new_B3068_ = new_C3796_;
  assign new_B3067_ = new_C3729_;
  assign new_B3066_ = ~new_B3005_ & new_B3019_;
  assign new_B3065_ = new_B3005_ & ~new_B3019_;
  assign new_B3064_ = new_B3005_ & ~new_B3019_;
  assign new_B3063_ = ~new_B3005_ & ~new_B3019_;
  assign new_B3062_ = new_B3005_ & new_B3019_;
  assign new_B3061_ = new_B3065_ | new_B3066_;
  assign new_B3060_ = ~new_B3005_ & new_B3019_;
  assign new_B3059_ = new_B3063_ | new_B3064_;
  assign new_B3058_ = ~new_B3034_ & ~new_B3054_;
  assign new_B3057_ = new_B3034_ & new_B3054_;
  assign new_B3056_ = ~new_B3001_ | ~new_B3026_;
  assign new_B3055_ = new_B3019_ & new_B3056_;
  assign new_B3054_ = new_B3002_ | new_B3003_;
  assign new_B3053_ = new_B3002_ | new_B3019_;
  assign new_B3052_ = ~new_B3019_ & ~new_B3055_;
  assign new_B3051_ = new_B3019_ | new_B3056_;
  assign new_B3050_ = new_B3002_ & ~new_B3003_;
  assign new_B3049_ = ~new_B3002_ & new_B3003_;
  assign new_B3048_ = new_B3012_ | new_B3045_;
  assign new_B3047_ = ~new_B3012_ & ~new_B3046_;
  assign new_B3046_ = new_B3012_ & new_B3045_;
  assign new_B3045_ = ~new_B3001_ | ~new_B3026_;
  assign new_B3044_ = ~new_B3002_ & new_B3012_;
  assign new_B3043_ = new_B3002_ & ~new_B3012_;
  assign new_B3042_ = new_B3004_ & new_B3041_;
  assign new_B3041_ = new_B3060_ | new_B3059_;
  assign new_B3040_ = ~new_B3004_ & new_B3039_;
  assign new_B3039_ = new_B3062_ | new_B3061_;
  assign new_B3038_ = new_B3004_ | new_B3037_;
  assign new_B3037_ = new_B3058_ | new_B3057_;
  assign new_B3036_ = ~new_B3016_ & ~new_B3026_;
  assign new_B3035_ = new_B3016_ & new_B3026_;
  assign new_B3034_ = ~new_B3016_ | new_B3026_;
  assign new_B3033_ = new_B3000_ & ~new_B3001_;
  assign new_B3032_ = ~new_B3000_ & new_B3001_;
  assign new_B3031_ = new_B3053_ & ~new_B3054_;
  assign new_B3030_ = ~new_B3053_ & new_B3054_;
  assign new_B3029_ = ~new_B3052_ | ~new_B3051_;
  assign new_B3028_ = new_B3044_ | new_B3043_;
  assign new_B3027_ = new_B3050_ | new_B3049_;
  assign new_B3026_ = new_B3040_ | new_B3042_;
  assign new_B3025_ = ~new_B3047_ | ~new_B3048_;
  assign new_B3024_ = new_B3000_ & ~new_B3001_;
  assign new_B3023_ = new_B3014_ & ~new_B3026_;
  assign new_B3022_ = ~new_B3014_ & new_B3026_;
  assign new_B3021_ = ~new_B3012_ & new_B3038_;
  assign new_B3020_ = new_B3036_ | new_B3035_;
  assign new_B3019_ = new_B3033_ | new_B3032_;
  assign new_B3018_ = new_B3001_ | new_B3034_;
  assign new_B3017_ = new_B3026_ & new_B3029_;
  assign new_B3016_ = new_B3031_ | new_B3030_;
  assign new_B3015_ = new_B3026_ & new_B3025_;
  assign new_B3014_ = new_B3028_ & new_B3027_;
  assign new_B3013_ = new_B3023_ | new_B3022_;
  assign new_B3012_ = new_B3001_ | new_B3024_;
  assign B3011 = new_B3012_ | new_B3021_;
  assign B3010 = new_B3019_ & new_B3020_;
  assign B3009 = new_B3019_ & new_B3018_;
  assign B3008 = new_B3017_ | new_B3016_;
  assign B3007 = new_B3015_ | new_B3014_;
  assign B3006 = new_B3013_ & new_B3012_;
  assign new_B3005_ = new_C3662_;
  assign new_B3004_ = new_C3595_;
  assign new_B3003_ = new_C3528_;
  assign new_B3002_ = new_C3461_;
  assign new_B3001_ = new_C3394_;
  assign new_B3000_ = new_C3327_;
  assign new_B2999_ = ~new_B2938_ & new_B2952_;
  assign new_B2998_ = new_B2938_ & ~new_B2952_;
  assign new_B2997_ = new_B2938_ & ~new_B2952_;
  assign new_B2996_ = ~new_B2938_ & ~new_B2952_;
  assign new_B2995_ = new_B2938_ & new_B2952_;
  assign new_B2994_ = new_B2998_ | new_B2999_;
  assign new_B2993_ = ~new_B2938_ & new_B2952_;
  assign new_B2992_ = new_B2996_ | new_B2997_;
  assign new_B2991_ = ~new_B2967_ & ~new_B2987_;
  assign new_B2990_ = new_B2967_ & new_B2987_;
  assign new_B2989_ = ~new_B2934_ | ~new_B2959_;
  assign new_B2988_ = new_B2952_ & new_B2989_;
  assign new_B2987_ = new_B2935_ | new_B2936_;
  assign new_B2986_ = new_B2935_ | new_B2952_;
  assign new_B2985_ = ~new_B2952_ & ~new_B2988_;
  assign new_B2984_ = new_B2952_ | new_B2989_;
  assign new_B2983_ = new_B2935_ & ~new_B2936_;
  assign new_B2982_ = ~new_B2935_ & new_B2936_;
  assign new_B2981_ = new_B2945_ | new_B2978_;
  assign new_B2980_ = ~new_B2945_ & ~new_B2979_;
  assign new_B2979_ = new_B2945_ & new_B2978_;
  assign new_B2978_ = ~new_B2934_ | ~new_B2959_;
  assign new_B2977_ = ~new_B2935_ & new_B2945_;
  assign new_B2976_ = new_B2935_ & ~new_B2945_;
  assign new_B2975_ = new_B2937_ & new_B2974_;
  assign new_B2974_ = new_B2993_ | new_B2992_;
  assign new_B2973_ = ~new_B2937_ & new_B2972_;
  assign new_B2972_ = new_B2995_ | new_B2994_;
  assign new_B2971_ = new_B2937_ | new_B2970_;
  assign new_B2970_ = new_B2991_ | new_B2990_;
  assign new_B2969_ = ~new_B2949_ & ~new_B2959_;
  assign new_B2968_ = new_B2949_ & new_B2959_;
  assign new_B2967_ = ~new_B2949_ | new_B2959_;
  assign new_B2966_ = new_B2933_ & ~new_B2934_;
  assign new_B2965_ = ~new_B2933_ & new_B2934_;
  assign new_B2964_ = new_B2986_ & ~new_B2987_;
  assign new_B2963_ = ~new_B2986_ & new_B2987_;
  assign new_B2962_ = ~new_B2985_ | ~new_B2984_;
  assign new_B2961_ = new_B2977_ | new_B2976_;
  assign new_B2960_ = new_B2983_ | new_B2982_;
  assign new_B2959_ = new_B2973_ | new_B2975_;
  assign new_B2958_ = ~new_B2980_ | ~new_B2981_;
  assign new_B2957_ = new_B2933_ & ~new_B2934_;
  assign new_B2956_ = new_B2947_ & ~new_B2959_;
  assign new_B2955_ = ~new_B2947_ & new_B2959_;
  assign new_B2954_ = ~new_B2945_ & new_B2971_;
  assign new_B2953_ = new_B2969_ | new_B2968_;
  assign new_B2952_ = new_B2966_ | new_B2965_;
  assign new_B2951_ = new_B2934_ | new_B2967_;
  assign new_B2950_ = new_B2959_ & new_B2962_;
  assign new_B2949_ = new_B2964_ | new_B2963_;
  assign new_B2948_ = new_B2959_ & new_B2958_;
  assign new_B2947_ = new_B2961_ & new_B2960_;
  assign new_B2946_ = new_B2956_ | new_B2955_;
  assign new_B2945_ = new_B2934_ | new_B2957_;
  assign B2944 = new_B2945_ | new_B2954_;
  assign B2943 = new_B2952_ & new_B2953_;
  assign B2942 = new_B2952_ & new_B2951_;
  assign B2941 = new_B2950_ | new_B2949_;
  assign B2940 = new_B2948_ | new_B2947_;
  assign B2939 = new_B2946_ & new_B2945_;
  assign new_B2938_ = new_C3260_;
  assign new_B2937_ = new_C3193_;
  assign new_B2936_ = new_C3126_;
  assign new_B2935_ = new_C3059_;
  assign new_B2934_ = new_C2992_;
  assign new_B2933_ = new_C2925_;
  assign new_B2932_ = ~new_B2871_ & new_B2885_;
  assign new_B2931_ = new_B2871_ & ~new_B2885_;
  assign new_B2930_ = new_B2871_ & ~new_B2885_;
  assign new_B2929_ = ~new_B2871_ & ~new_B2885_;
  assign new_B2928_ = new_B2871_ & new_B2885_;
  assign new_B2927_ = new_B2931_ | new_B2932_;
  assign new_B2926_ = ~new_B2871_ & new_B2885_;
  assign new_B2925_ = new_B2929_ | new_B2930_;
  assign new_B2924_ = ~new_B2900_ & ~new_B2920_;
  assign new_B2923_ = new_B2900_ & new_B2920_;
  assign new_B2922_ = ~new_B2867_ | ~new_B2892_;
  assign new_B2921_ = new_B2885_ & new_B2922_;
  assign new_B2920_ = new_B2868_ | new_B2869_;
  assign new_B2919_ = new_B2868_ | new_B2885_;
  assign new_B2918_ = ~new_B2885_ & ~new_B2921_;
  assign new_B2917_ = new_B2885_ | new_B2922_;
  assign new_B2916_ = new_B2868_ & ~new_B2869_;
  assign new_B2915_ = ~new_B2868_ & new_B2869_;
  assign new_B2914_ = new_B2878_ | new_B2911_;
  assign new_B2913_ = ~new_B2878_ & ~new_B2912_;
  assign new_B2912_ = new_B2878_ & new_B2911_;
  assign new_B2911_ = ~new_B2867_ | ~new_B2892_;
  assign new_B2910_ = ~new_B2868_ & new_B2878_;
  assign new_B2909_ = new_B2868_ & ~new_B2878_;
  assign new_B2908_ = new_B2870_ & new_B2907_;
  assign new_B2907_ = new_B2926_ | new_B2925_;
  assign new_B2906_ = ~new_B2870_ & new_B2905_;
  assign new_B2905_ = new_B2928_ | new_B2927_;
  assign new_B2904_ = new_B2870_ | new_B2903_;
  assign new_B2903_ = new_B2924_ | new_B2923_;
  assign new_B2902_ = ~new_B2882_ & ~new_B2892_;
  assign new_B2901_ = new_B2882_ & new_B2892_;
  assign new_B2900_ = ~new_B2882_ | new_B2892_;
  assign new_B2899_ = new_B2866_ & ~new_B2867_;
  assign new_B2898_ = ~new_B2866_ & new_B2867_;
  assign new_B2897_ = new_B2919_ & ~new_B2920_;
  assign new_B2896_ = ~new_B2919_ & new_B2920_;
  assign new_B2895_ = ~new_B2918_ | ~new_B2917_;
  assign new_B2894_ = new_B2910_ | new_B2909_;
  assign new_B2893_ = new_B2916_ | new_B2915_;
  assign new_B2892_ = new_B2906_ | new_B2908_;
  assign new_B2891_ = ~new_B2913_ | ~new_B2914_;
  assign new_B2890_ = new_B2866_ & ~new_B2867_;
  assign new_B2889_ = new_B2880_ & ~new_B2892_;
  assign new_B2888_ = ~new_B2880_ & new_B2892_;
  assign new_B2887_ = ~new_B2878_ & new_B2904_;
  assign new_B2886_ = new_B2902_ | new_B2901_;
  assign new_B2885_ = new_B2899_ | new_B2898_;
  assign new_B2884_ = new_B2867_ | new_B2900_;
  assign new_B2883_ = new_B2892_ & new_B2895_;
  assign new_B2882_ = new_B2897_ | new_B2896_;
  assign new_B2881_ = new_B2892_ & new_B2891_;
  assign new_B2880_ = new_B2894_ & new_B2893_;
  assign new_B2879_ = new_B2889_ | new_B2888_;
  assign new_B2878_ = new_B2867_ | new_B2890_;
  assign B2877 = new_B2878_ | new_B2887_;
  assign B2876 = new_B2885_ & new_B2886_;
  assign B2875 = new_B2885_ & new_B2884_;
  assign B2874 = new_B2883_ | new_B2882_;
  assign B2873 = new_B2881_ | new_B2880_;
  assign B2872 = new_B2879_ & new_B2878_;
  assign new_B2871_ = new_C2858_;
  assign new_B2870_ = new_C2791_;
  assign new_B2869_ = new_C2724_;
  assign new_B2868_ = new_C2657_;
  assign new_B2867_ = new_C2590_;
  assign new_B2866_ = new_C2524_;
  assign new_B2865_ = ~new_B2804_ & new_B2818_;
  assign new_B2864_ = new_B2804_ & ~new_B2818_;
  assign new_B2863_ = new_B2804_ & ~new_B2818_;
  assign new_B2862_ = ~new_B2804_ & ~new_B2818_;
  assign new_B2861_ = new_B2804_ & new_B2818_;
  assign new_B2860_ = new_B2864_ | new_B2865_;
  assign new_B2859_ = ~new_B2804_ & new_B2818_;
  assign new_B2858_ = new_B2862_ | new_B2863_;
  assign new_B2857_ = ~new_B2833_ & ~new_B2853_;
  assign new_B2856_ = new_B2833_ & new_B2853_;
  assign new_B2855_ = ~new_B2800_ | ~new_B2825_;
  assign new_B2854_ = new_B2818_ & new_B2855_;
  assign new_B2853_ = new_B2801_ | new_B2802_;
  assign new_B2852_ = new_B2801_ | new_B2818_;
  assign new_B2851_ = ~new_B2818_ & ~new_B2854_;
  assign new_B2850_ = new_B2818_ | new_B2855_;
  assign new_B2849_ = new_B2801_ & ~new_B2802_;
  assign new_B2848_ = ~new_B2801_ & new_B2802_;
  assign new_B2847_ = new_B2811_ | new_B2844_;
  assign new_B2846_ = ~new_B2811_ & ~new_B2845_;
  assign new_B2845_ = new_B2811_ & new_B2844_;
  assign new_B2844_ = ~new_B2800_ | ~new_B2825_;
  assign new_B2843_ = ~new_B2801_ & new_B2811_;
  assign new_B2842_ = new_B2801_ & ~new_B2811_;
  assign new_B2841_ = new_B2803_ & new_B2840_;
  assign new_B2840_ = new_B2859_ | new_B2858_;
  assign new_B2839_ = ~new_B2803_ & new_B2838_;
  assign new_B2838_ = new_B2861_ | new_B2860_;
  assign new_B2837_ = new_B2803_ | new_B2836_;
  assign new_B2836_ = new_B2857_ | new_B2856_;
  assign new_B2835_ = ~new_B2815_ & ~new_B2825_;
  assign new_B2834_ = new_B2815_ & new_B2825_;
  assign new_B2833_ = ~new_B2815_ | new_B2825_;
  assign new_B2832_ = new_B2799_ & ~new_B2800_;
  assign new_B2831_ = ~new_B2799_ & new_B2800_;
  assign new_B2830_ = new_B2852_ & ~new_B2853_;
  assign new_B2829_ = ~new_B2852_ & new_B2853_;
  assign new_B2828_ = ~new_B2851_ | ~new_B2850_;
  assign new_B2827_ = new_B2843_ | new_B2842_;
  assign new_B2826_ = new_B2849_ | new_B2848_;
  assign new_B2825_ = new_B2839_ | new_B2841_;
  assign new_B2824_ = ~new_B2846_ | ~new_B2847_;
  assign new_B2823_ = new_B2799_ & ~new_B2800_;
  assign new_B2822_ = new_B2813_ & ~new_B2825_;
  assign new_B2821_ = ~new_B2813_ & new_B2825_;
  assign new_B2820_ = ~new_B2811_ & new_B2837_;
  assign new_B2819_ = new_B2835_ | new_B2834_;
  assign new_B2818_ = new_B2832_ | new_B2831_;
  assign new_B2817_ = new_B2800_ | new_B2833_;
  assign new_B2816_ = new_B2825_ & new_B2828_;
  assign new_B2815_ = new_B2830_ | new_B2829_;
  assign new_B2814_ = new_B2825_ & new_B2824_;
  assign new_B2813_ = new_B2827_ & new_B2826_;
  assign new_B2812_ = new_B2822_ | new_B2821_;
  assign new_B2811_ = new_B2800_ | new_B2823_;
  assign B2810 = new_B2811_ | new_B2820_;
  assign B2809 = new_B2818_ & new_B2819_;
  assign B2808 = new_B2818_ & new_B2817_;
  assign B2807 = new_B2816_ | new_B2815_;
  assign B2806 = new_B2814_ | new_B2813_;
  assign B2805 = new_B2812_ & new_B2811_;
  assign new_B2804_ = new_D6928_;
  assign new_B2803_ = new_D6861_;
  assign new_B2802_ = new_D6794_;
  assign new_B2801_ = new_D6727_;
  assign new_B2800_ = new_D6660_;
  assign new_B2799_ = new_D6593_;
  assign new_B2798_ = ~new_B2737_ & new_B2751_;
  assign new_B2797_ = new_B2737_ & ~new_B2751_;
  assign new_B2796_ = new_B2737_ & ~new_B2751_;
  assign new_B2795_ = ~new_B2737_ & ~new_B2751_;
  assign new_B2794_ = new_B2737_ & new_B2751_;
  assign new_B2793_ = new_B2797_ | new_B2798_;
  assign new_B2792_ = ~new_B2737_ & new_B2751_;
  assign new_B2791_ = new_B2795_ | new_B2796_;
  assign new_B2790_ = ~new_B2766_ & ~new_B2786_;
  assign new_B2789_ = new_B2766_ & new_B2786_;
  assign new_B2788_ = ~new_B2733_ | ~new_B2758_;
  assign new_B2787_ = new_B2751_ & new_B2788_;
  assign new_B2786_ = new_B2734_ | new_B2735_;
  assign new_B2785_ = new_B2734_ | new_B2751_;
  assign new_B2784_ = ~new_B2751_ & ~new_B2787_;
  assign new_B2783_ = new_B2751_ | new_B2788_;
  assign new_B2782_ = new_B2734_ & ~new_B2735_;
  assign new_B2781_ = ~new_B2734_ & new_B2735_;
  assign new_B2780_ = new_B2744_ | new_B2777_;
  assign new_B2779_ = ~new_B2744_ & ~new_B2778_;
  assign new_B2778_ = new_B2744_ & new_B2777_;
  assign new_B2777_ = ~new_B2733_ | ~new_B2758_;
  assign new_B2776_ = ~new_B2734_ & new_B2744_;
  assign new_B2775_ = new_B2734_ & ~new_B2744_;
  assign new_B2774_ = new_B2736_ & new_B2773_;
  assign new_B2773_ = new_B2792_ | new_B2791_;
  assign new_B2772_ = ~new_B2736_ & new_B2771_;
  assign new_B2771_ = new_B2794_ | new_B2793_;
  assign new_B2770_ = new_B2736_ | new_B2769_;
  assign new_B2769_ = new_B2790_ | new_B2789_;
  assign new_B2768_ = ~new_B2748_ & ~new_B2758_;
  assign new_B2767_ = new_B2748_ & new_B2758_;
  assign new_B2766_ = ~new_B2748_ | new_B2758_;
  assign new_B2765_ = new_B2732_ & ~new_B2733_;
  assign new_B2764_ = ~new_B2732_ & new_B2733_;
  assign new_B2763_ = new_B2785_ & ~new_B2786_;
  assign new_B2762_ = ~new_B2785_ & new_B2786_;
  assign new_B2761_ = ~new_B2784_ | ~new_B2783_;
  assign new_B2760_ = new_B2776_ | new_B2775_;
  assign new_B2759_ = new_B2782_ | new_B2781_;
  assign new_B2758_ = new_B2772_ | new_B2774_;
  assign new_B2757_ = ~new_B2779_ | ~new_B2780_;
  assign new_B2756_ = new_B2732_ & ~new_B2733_;
  assign new_B2755_ = new_B2746_ & ~new_B2758_;
  assign new_B2754_ = ~new_B2746_ & new_B2758_;
  assign new_B2753_ = ~new_B2744_ & new_B2770_;
  assign new_B2752_ = new_B2768_ | new_B2767_;
  assign new_B2751_ = new_B2765_ | new_B2764_;
  assign new_B2750_ = new_B2733_ | new_B2766_;
  assign new_B2749_ = new_B2758_ & new_B2761_;
  assign new_B2748_ = new_B2763_ | new_B2762_;
  assign new_B2747_ = new_B2758_ & new_B2757_;
  assign new_B2746_ = new_B2760_ & new_B2759_;
  assign new_B2745_ = new_B2755_ | new_B2754_;
  assign new_B2744_ = new_B2733_ | new_B2756_;
  assign B2743 = new_B2744_ | new_B2753_;
  assign B2742 = new_B2751_ & new_B2752_;
  assign B2741 = new_B2751_ & new_B2750_;
  assign B2740 = new_B2749_ | new_B2748_;
  assign B2739 = new_B2747_ | new_B2746_;
  assign B2738 = new_B2745_ & new_B2744_;
  assign new_B2737_ = new_D6526_;
  assign new_B2736_ = new_D6459_;
  assign new_B2735_ = new_D6392_;
  assign new_B2734_ = new_D6325_;
  assign new_B2733_ = new_D6258_;
  assign new_B2732_ = new_D6191_;
  assign new_B2731_ = ~new_B2670_ & new_B2684_;
  assign new_B2730_ = new_B2670_ & ~new_B2684_;
  assign new_B2729_ = new_B2670_ & ~new_B2684_;
  assign new_B2728_ = ~new_B2670_ & ~new_B2684_;
  assign new_B2727_ = new_B2670_ & new_B2684_;
  assign new_B2726_ = new_B2730_ | new_B2731_;
  assign new_B2725_ = ~new_B2670_ & new_B2684_;
  assign new_B2724_ = new_B2728_ | new_B2729_;
  assign new_B2723_ = ~new_B2699_ & ~new_B2719_;
  assign new_B2722_ = new_B2699_ & new_B2719_;
  assign new_B2721_ = ~new_B2666_ | ~new_B2691_;
  assign new_B2720_ = new_B2684_ & new_B2721_;
  assign new_B2719_ = new_B2667_ | new_B2668_;
  assign new_B2718_ = new_B2667_ | new_B2684_;
  assign new_B2717_ = ~new_B2684_ & ~new_B2720_;
  assign new_B2716_ = new_B2684_ | new_B2721_;
  assign new_B2715_ = new_B2667_ & ~new_B2668_;
  assign new_B2714_ = ~new_B2667_ & new_B2668_;
  assign new_B2713_ = new_B2677_ | new_B2710_;
  assign new_B2712_ = ~new_B2677_ & ~new_B2711_;
  assign new_B2711_ = new_B2677_ & new_B2710_;
  assign new_B2710_ = ~new_B2666_ | ~new_B2691_;
  assign new_B2709_ = ~new_B2667_ & new_B2677_;
  assign new_B2708_ = new_B2667_ & ~new_B2677_;
  assign new_B2707_ = new_B2669_ & new_B2706_;
  assign new_B2706_ = new_B2725_ | new_B2724_;
  assign new_B2705_ = ~new_B2669_ & new_B2704_;
  assign new_B2704_ = new_B2727_ | new_B2726_;
  assign new_B2703_ = new_B2669_ | new_B2702_;
  assign new_B2702_ = new_B2723_ | new_B2722_;
  assign new_B2701_ = ~new_B2681_ & ~new_B2691_;
  assign new_B2700_ = new_B2681_ & new_B2691_;
  assign new_B2699_ = ~new_B2681_ | new_B2691_;
  assign new_B2698_ = new_B2665_ & ~new_B2666_;
  assign new_B2697_ = ~new_B2665_ & new_B2666_;
  assign new_B2696_ = new_B2718_ & ~new_B2719_;
  assign new_B2695_ = ~new_B2718_ & new_B2719_;
  assign new_B2694_ = ~new_B2717_ | ~new_B2716_;
  assign new_B2693_ = new_B2709_ | new_B2708_;
  assign new_B2692_ = new_B2715_ | new_B2714_;
  assign new_B2691_ = new_B2705_ | new_B2707_;
  assign new_B2690_ = ~new_B2712_ | ~new_B2713_;
  assign new_B2689_ = new_B2665_ & ~new_B2666_;
  assign new_B2688_ = new_B2679_ & ~new_B2691_;
  assign new_B2687_ = ~new_B2679_ & new_B2691_;
  assign new_B2686_ = ~new_B2677_ & new_B2703_;
  assign new_B2685_ = new_B2701_ | new_B2700_;
  assign new_B2684_ = new_B2698_ | new_B2697_;
  assign new_B2683_ = new_B2666_ | new_B2699_;
  assign new_B2682_ = new_B2691_ & new_B2694_;
  assign new_B2681_ = new_B2696_ | new_B2695_;
  assign new_B2680_ = new_B2691_ & new_B2690_;
  assign new_B2679_ = new_B2693_ & new_B2692_;
  assign new_B2678_ = new_B2688_ | new_B2687_;
  assign new_B2677_ = new_B2666_ | new_B2689_;
  assign B2676 = new_B2677_ | new_B2686_;
  assign B2675 = new_B2684_ & new_B2685_;
  assign B2674 = new_B2684_ & new_B2683_;
  assign B2673 = new_B2682_ | new_B2681_;
  assign B2672 = new_B2680_ | new_B2679_;
  assign B2671 = new_B2678_ & new_B2677_;
  assign new_B2670_ = new_D6124_;
  assign new_B2669_ = new_D6057_;
  assign new_B2668_ = new_D5990_;
  assign new_B2667_ = new_D5923_;
  assign new_B2666_ = new_D5856_;
  assign new_B2665_ = new_D5789_;
  assign new_B2664_ = ~new_B2603_ & new_B2617_;
  assign new_B2663_ = new_B2603_ & ~new_B2617_;
  assign new_B2662_ = new_B2603_ & ~new_B2617_;
  assign new_B2661_ = ~new_B2603_ & ~new_B2617_;
  assign new_B2660_ = new_B2603_ & new_B2617_;
  assign new_B2659_ = new_B2663_ | new_B2664_;
  assign new_B2658_ = ~new_B2603_ & new_B2617_;
  assign new_B2657_ = new_B2661_ | new_B2662_;
  assign new_B2656_ = ~new_B2632_ & ~new_B2652_;
  assign new_B2655_ = new_B2632_ & new_B2652_;
  assign new_B2654_ = ~new_B2599_ | ~new_B2624_;
  assign new_B2653_ = new_B2617_ & new_B2654_;
  assign new_B2652_ = new_B2600_ | new_B2601_;
  assign new_B2651_ = new_B2600_ | new_B2617_;
  assign new_B2650_ = ~new_B2617_ & ~new_B2653_;
  assign new_B2649_ = new_B2617_ | new_B2654_;
  assign new_B2648_ = new_B2600_ & ~new_B2601_;
  assign new_B2647_ = ~new_B2600_ & new_B2601_;
  assign new_B2646_ = new_B2610_ | new_B2643_;
  assign new_B2645_ = ~new_B2610_ & ~new_B2644_;
  assign new_B2644_ = new_B2610_ & new_B2643_;
  assign new_B2643_ = ~new_B2599_ | ~new_B2624_;
  assign new_B2642_ = ~new_B2600_ & new_B2610_;
  assign new_B2641_ = new_B2600_ & ~new_B2610_;
  assign new_B2640_ = new_B2602_ & new_B2639_;
  assign new_B2639_ = new_B2658_ | new_B2657_;
  assign new_B2638_ = ~new_B2602_ & new_B2637_;
  assign new_B2637_ = new_B2660_ | new_B2659_;
  assign new_B2636_ = new_B2602_ | new_B2635_;
  assign new_B2635_ = new_B2656_ | new_B2655_;
  assign new_B2634_ = ~new_B2614_ & ~new_B2624_;
  assign new_B2633_ = new_B2614_ & new_B2624_;
  assign new_B2632_ = ~new_B2614_ | new_B2624_;
  assign new_B2631_ = new_B2598_ & ~new_B2599_;
  assign new_B2630_ = ~new_B2598_ & new_B2599_;
  assign new_B2629_ = new_B2651_ & ~new_B2652_;
  assign new_B2628_ = ~new_B2651_ & new_B2652_;
  assign new_B2627_ = ~new_B2650_ | ~new_B2649_;
  assign new_B2626_ = new_B2642_ | new_B2641_;
  assign new_B2625_ = new_B2648_ | new_B2647_;
  assign new_B2624_ = new_B2638_ | new_B2640_;
  assign new_B2623_ = ~new_B2645_ | ~new_B2646_;
  assign new_B2622_ = new_B2598_ & ~new_B2599_;
  assign new_B2621_ = new_B2612_ & ~new_B2624_;
  assign new_B2620_ = ~new_B2612_ & new_B2624_;
  assign new_B2619_ = ~new_B2610_ & new_B2636_;
  assign new_B2618_ = new_B2634_ | new_B2633_;
  assign new_B2617_ = new_B2631_ | new_B2630_;
  assign new_B2616_ = new_B2599_ | new_B2632_;
  assign new_B2615_ = new_B2624_ & new_B2627_;
  assign new_B2614_ = new_B2629_ | new_B2628_;
  assign new_B2613_ = new_B2624_ & new_B2623_;
  assign new_B2612_ = new_B2626_ & new_B2625_;
  assign new_B2611_ = new_B2621_ | new_B2620_;
  assign new_B2610_ = new_B2599_ | new_B2622_;
  assign B2609 = new_B2610_ | new_B2619_;
  assign B2608 = new_B2617_ & new_B2618_;
  assign B2607 = new_B2617_ & new_B2616_;
  assign B2606 = new_B2615_ | new_B2614_;
  assign B2605 = new_B2613_ | new_B2612_;
  assign B2604 = new_B2611_ & new_B2610_;
  assign new_B2603_ = new_D5722_;
  assign new_B2602_ = new_D5655_;
  assign new_B2601_ = new_D5588_;
  assign new_B2600_ = new_D5521_;
  assign new_B2599_ = new_D5454_;
  assign new_B2598_ = new_D5387_;
  assign new_B2597_ = ~new_B2536_ & new_B2550_;
  assign new_B2596_ = new_B2536_ & ~new_B2550_;
  assign new_B2595_ = new_B2536_ & ~new_B2550_;
  assign new_B2594_ = ~new_B2536_ & ~new_B2550_;
  assign new_B2593_ = new_B2536_ & new_B2550_;
  assign new_B2592_ = new_B2596_ | new_B2597_;
  assign new_B2591_ = ~new_B2536_ & new_B2550_;
  assign new_B2590_ = new_B2594_ | new_B2595_;
  assign new_B2589_ = ~new_B2565_ & ~new_B2585_;
  assign new_B2588_ = new_B2565_ & new_B2585_;
  assign new_B2587_ = ~new_B2532_ | ~new_B2557_;
  assign new_B2586_ = new_B2550_ & new_B2587_;
  assign new_B2585_ = new_B2533_ | new_B2534_;
  assign new_B2584_ = new_B2533_ | new_B2550_;
  assign new_B2583_ = ~new_B2550_ & ~new_B2586_;
  assign new_B2582_ = new_B2550_ | new_B2587_;
  assign new_B2581_ = new_B2533_ & ~new_B2534_;
  assign new_B2580_ = ~new_B2533_ & new_B2534_;
  assign new_B2579_ = new_B2543_ | new_B2576_;
  assign new_B2578_ = ~new_B2543_ & ~new_B2577_;
  assign new_B2577_ = new_B2543_ & new_B2576_;
  assign new_B2576_ = ~new_B2532_ | ~new_B2557_;
  assign new_B2575_ = ~new_B2533_ & new_B2543_;
  assign new_B2574_ = new_B2533_ & ~new_B2543_;
  assign new_B2573_ = new_B2535_ & new_B2572_;
  assign new_B2572_ = new_B2591_ | new_B2590_;
  assign new_B2571_ = ~new_B2535_ & new_B2570_;
  assign new_B2570_ = new_B2593_ | new_B2592_;
  assign new_B2569_ = new_B2535_ | new_B2568_;
  assign new_B2568_ = new_B2589_ | new_B2588_;
  assign new_B2567_ = ~new_B2547_ & ~new_B2557_;
  assign new_B2566_ = new_B2547_ & new_B2557_;
  assign new_B2565_ = ~new_B2547_ | new_B2557_;
  assign new_B2564_ = new_B2531_ & ~new_B2532_;
  assign new_B2563_ = ~new_B2531_ & new_B2532_;
  assign new_B2562_ = new_B2584_ & ~new_B2585_;
  assign new_B2561_ = ~new_B2584_ & new_B2585_;
  assign new_B2560_ = ~new_B2583_ | ~new_B2582_;
  assign new_B2559_ = new_B2575_ | new_B2574_;
  assign new_B2558_ = new_B2581_ | new_B2580_;
  assign new_B2557_ = new_B2571_ | new_B2573_;
  assign new_B2556_ = ~new_B2578_ | ~new_B2579_;
  assign new_B2555_ = new_B2531_ & ~new_B2532_;
  assign new_B2554_ = new_B2545_ & ~new_B2557_;
  assign new_B2553_ = ~new_B2545_ & new_B2557_;
  assign new_B2552_ = ~new_B2543_ & new_B2569_;
  assign new_B2551_ = new_B2567_ | new_B2566_;
  assign new_B2550_ = new_B2564_ | new_B2563_;
  assign new_B2549_ = new_B2532_ | new_B2565_;
  assign new_B2548_ = new_B2557_ & new_B2560_;
  assign new_B2547_ = new_B2562_ | new_B2561_;
  assign new_B2546_ = new_B2557_ & new_B2556_;
  assign new_B2545_ = new_B2559_ & new_B2558_;
  assign new_B2544_ = new_B2554_ | new_B2553_;
  assign new_B2543_ = new_B2532_ | new_B2555_;
  assign B2542 = new_B2543_ | new_B2552_;
  assign B2541 = new_B2550_ & new_B2551_;
  assign B2540 = new_B2550_ & new_B2549_;
  assign B2539 = new_B2548_ | new_B2547_;
  assign B2538 = new_B2546_ | new_B2545_;
  assign B2537 = new_B2544_ & new_B2543_;
  assign new_B2536_ = new_D5320_;
  assign new_B2535_ = new_D5253_;
  assign new_B2534_ = new_D5186_;
  assign new_B2533_ = new_D5119_;
  assign new_B2532_ = new_D5052_;
  assign new_B2531_ = new_D4985_;
  assign new_B2530_ = ~new_B2469_ & new_B2483_;
  assign new_B2529_ = new_B2469_ & ~new_B2483_;
  assign new_B2528_ = new_B2469_ & ~new_B2483_;
  assign new_B2527_ = ~new_B2469_ & ~new_B2483_;
  assign new_B2526_ = new_B2469_ & new_B2483_;
  assign new_B2525_ = new_B2529_ | new_B2530_;
  assign new_B2524_ = ~new_B2469_ & new_B2483_;
  assign new_B2523_ = new_B2527_ | new_B2528_;
  assign new_B2522_ = ~new_B2498_ & ~new_B2518_;
  assign new_B2521_ = new_B2498_ & new_B2518_;
  assign new_B2520_ = ~new_B2465_ | ~new_B2490_;
  assign new_B2519_ = new_B2483_ & new_B2520_;
  assign new_B2518_ = new_B2466_ | new_B2467_;
  assign new_B2517_ = new_B2466_ | new_B2483_;
  assign new_B2516_ = ~new_B2483_ & ~new_B2519_;
  assign new_B2515_ = new_B2483_ | new_B2520_;
  assign new_B2514_ = new_B2466_ & ~new_B2467_;
  assign new_B2513_ = ~new_B2466_ & new_B2467_;
  assign new_B2512_ = new_B2476_ | new_B2509_;
  assign new_B2511_ = ~new_B2476_ & ~new_B2510_;
  assign new_B2510_ = new_B2476_ & new_B2509_;
  assign new_B2509_ = ~new_B2465_ | ~new_B2490_;
  assign new_B2508_ = ~new_B2466_ & new_B2476_;
  assign new_B2507_ = new_B2466_ & ~new_B2476_;
  assign new_B2506_ = new_B2468_ & new_B2505_;
  assign new_B2505_ = new_B2524_ | new_B2523_;
  assign new_B2504_ = ~new_B2468_ & new_B2503_;
  assign new_B2503_ = new_B2526_ | new_B2525_;
  assign new_B2502_ = new_B2468_ | new_B2501_;
  assign new_B2501_ = new_B2522_ | new_B2521_;
  assign new_B2500_ = ~new_B2480_ & ~new_B2490_;
  assign new_B2499_ = new_B2480_ & new_B2490_;
  assign new_B2498_ = ~new_B2480_ | new_B2490_;
  assign new_B2497_ = new_B2464_ & ~new_B2465_;
  assign new_B2496_ = ~new_B2464_ & new_B2465_;
  assign new_B2495_ = new_B2517_ & ~new_B2518_;
  assign new_B2494_ = ~new_B2517_ & new_B2518_;
  assign new_B2493_ = ~new_B2516_ | ~new_B2515_;
  assign new_B2492_ = new_B2508_ | new_B2507_;
  assign new_B2491_ = new_B2514_ | new_B2513_;
  assign new_B2490_ = new_B2504_ | new_B2506_;
  assign new_B2489_ = ~new_B2511_ | ~new_B2512_;
  assign new_B2488_ = new_B2464_ & ~new_B2465_;
  assign new_B2487_ = new_B2478_ & ~new_B2490_;
  assign new_B2486_ = ~new_B2478_ & new_B2490_;
  assign new_B2485_ = ~new_B2476_ & new_B2502_;
  assign new_B2484_ = new_B2500_ | new_B2499_;
  assign new_B2483_ = new_B2497_ | new_B2496_;
  assign new_B2482_ = new_B2465_ | new_B2498_;
  assign new_B2481_ = new_B2490_ & new_B2493_;
  assign new_B2480_ = new_B2495_ | new_B2494_;
  assign new_B2479_ = new_B2490_ & new_B2489_;
  assign new_B2478_ = new_B2492_ & new_B2491_;
  assign new_B2477_ = new_B2487_ | new_B2486_;
  assign new_B2476_ = new_B2465_ | new_B2488_;
  assign B2475 = new_B2476_ | new_B2485_;
  assign B2474 = new_B2483_ & new_B2484_;
  assign B2473 = new_B2483_ & new_B2482_;
  assign B2472 = new_B2481_ | new_B2480_;
  assign B2471 = new_B2479_ | new_B2478_;
  assign B2470 = new_B2477_ & new_B2476_;
  assign new_B2469_ = new_D4918_;
  assign new_B2468_ = new_D4851_;
  assign new_B2467_ = new_D4784_;
  assign new_B2466_ = new_D4717_;
  assign new_B2465_ = new_D4650_;
  assign new_B2464_ = new_D4583_;
  assign new_B2463_ = ~new_B2402_ & new_B2416_;
  assign new_B2462_ = new_B2402_ & ~new_B2416_;
  assign new_B2461_ = new_B2402_ & ~new_B2416_;
  assign new_B2460_ = ~new_B2402_ & ~new_B2416_;
  assign new_B2459_ = new_B2402_ & new_B2416_;
  assign new_B2458_ = new_B2462_ | new_B2463_;
  assign new_B2457_ = ~new_B2402_ & new_B2416_;
  assign new_B2456_ = new_B2460_ | new_B2461_;
  assign new_B2455_ = ~new_B2431_ & ~new_B2451_;
  assign new_B2454_ = new_B2431_ & new_B2451_;
  assign new_B2453_ = ~new_B2398_ | ~new_B2423_;
  assign new_B2452_ = new_B2416_ & new_B2453_;
  assign new_B2451_ = new_B2399_ | new_B2400_;
  assign new_B2450_ = new_B2399_ | new_B2416_;
  assign new_B2449_ = ~new_B2416_ & ~new_B2452_;
  assign new_B2448_ = new_B2416_ | new_B2453_;
  assign new_B2447_ = new_B2399_ & ~new_B2400_;
  assign new_B2446_ = ~new_B2399_ & new_B2400_;
  assign new_B2445_ = new_B2409_ | new_B2442_;
  assign new_B2444_ = ~new_B2409_ & ~new_B2443_;
  assign new_B2443_ = new_B2409_ & new_B2442_;
  assign new_B2442_ = ~new_B2398_ | ~new_B2423_;
  assign new_B2441_ = ~new_B2399_ & new_B2409_;
  assign new_B2440_ = new_B2399_ & ~new_B2409_;
  assign new_B2439_ = new_B2401_ & new_B2438_;
  assign new_B2438_ = new_B2457_ | new_B2456_;
  assign new_B2437_ = ~new_B2401_ & new_B2436_;
  assign new_B2436_ = new_B2459_ | new_B2458_;
  assign new_B2435_ = new_B2401_ | new_B2434_;
  assign new_B2434_ = new_B2455_ | new_B2454_;
  assign new_B2433_ = ~new_B2413_ & ~new_B2423_;
  assign new_B2432_ = new_B2413_ & new_B2423_;
  assign new_B2431_ = ~new_B2413_ | new_B2423_;
  assign new_B2430_ = new_B2397_ & ~new_B2398_;
  assign new_B2429_ = ~new_B2397_ & new_B2398_;
  assign new_B2428_ = new_B2450_ & ~new_B2451_;
  assign new_B2427_ = ~new_B2450_ & new_B2451_;
  assign new_B2426_ = ~new_B2449_ | ~new_B2448_;
  assign new_B2425_ = new_B2441_ | new_B2440_;
  assign new_B2424_ = new_B2447_ | new_B2446_;
  assign new_B2423_ = new_B2437_ | new_B2439_;
  assign new_B2422_ = ~new_B2444_ | ~new_B2445_;
  assign new_B2421_ = new_B2397_ & ~new_B2398_;
  assign new_B2420_ = new_B2411_ & ~new_B2423_;
  assign new_B2419_ = ~new_B2411_ & new_B2423_;
  assign new_B2418_ = ~new_B2409_ & new_B2435_;
  assign new_B2417_ = new_B2433_ | new_B2432_;
  assign new_B2416_ = new_B2430_ | new_B2429_;
  assign new_B2415_ = new_B2398_ | new_B2431_;
  assign new_B2414_ = new_B2423_ & new_B2426_;
  assign new_B2413_ = new_B2428_ | new_B2427_;
  assign new_B2412_ = new_B2423_ & new_B2422_;
  assign new_B2411_ = new_B2425_ & new_B2424_;
  assign new_B2410_ = new_B2420_ | new_B2419_;
  assign new_B2409_ = new_B2398_ | new_B2421_;
  assign B2408 = new_B2409_ | new_B2418_;
  assign B2407 = new_B2416_ & new_B2417_;
  assign B2406 = new_B2416_ & new_B2415_;
  assign B2405 = new_B2414_ | new_B2413_;
  assign B2404 = new_B2412_ | new_B2411_;
  assign B2403 = new_B2410_ & new_B2409_;
  assign new_B2402_ = new_D4516_;
  assign new_B2401_ = new_D4449_;
  assign new_B2400_ = new_D4382_;
  assign new_B2399_ = new_D4315_;
  assign new_B2398_ = new_D4248_;
  assign new_B2397_ = new_D4181_;
  assign new_B2396_ = ~new_B2335_ & new_B2349_;
  assign new_B2395_ = new_B2335_ & ~new_B2349_;
  assign new_B2394_ = new_B2335_ & ~new_B2349_;
  assign new_B2393_ = ~new_B2335_ & ~new_B2349_;
  assign new_B2392_ = new_B2335_ & new_B2349_;
  assign new_B2391_ = new_B2395_ | new_B2396_;
  assign new_B2390_ = ~new_B2335_ & new_B2349_;
  assign new_B2389_ = new_B2393_ | new_B2394_;
  assign new_B2388_ = ~new_B2364_ & ~new_B2384_;
  assign new_B2387_ = new_B2364_ & new_B2384_;
  assign new_B2386_ = ~new_B2331_ | ~new_B2356_;
  assign new_B2385_ = new_B2349_ & new_B2386_;
  assign new_B2384_ = new_B2332_ | new_B2333_;
  assign new_B2383_ = new_B2332_ | new_B2349_;
  assign new_B2382_ = ~new_B2349_ & ~new_B2385_;
  assign new_B2381_ = new_B2349_ | new_B2386_;
  assign new_B2380_ = new_B2332_ & ~new_B2333_;
  assign new_B2379_ = ~new_B2332_ & new_B2333_;
  assign new_B2378_ = new_B2342_ | new_B2375_;
  assign new_B2377_ = ~new_B2342_ & ~new_B2376_;
  assign new_B2376_ = new_B2342_ & new_B2375_;
  assign new_B2375_ = ~new_B2331_ | ~new_B2356_;
  assign new_B2374_ = ~new_B2332_ & new_B2342_;
  assign new_B2373_ = new_B2332_ & ~new_B2342_;
  assign new_B2372_ = new_B2334_ & new_B2371_;
  assign new_B2371_ = new_B2390_ | new_B2389_;
  assign new_B2370_ = ~new_B2334_ & new_B2369_;
  assign new_B2369_ = new_B2392_ | new_B2391_;
  assign new_B2368_ = new_B2334_ | new_B2367_;
  assign new_B2367_ = new_B2388_ | new_B2387_;
  assign new_B2366_ = ~new_B2346_ & ~new_B2356_;
  assign new_B2365_ = new_B2346_ & new_B2356_;
  assign new_B2364_ = ~new_B2346_ | new_B2356_;
  assign new_B2363_ = new_B2330_ & ~new_B2331_;
  assign new_B2362_ = ~new_B2330_ & new_B2331_;
  assign new_B2361_ = new_B2383_ & ~new_B2384_;
  assign new_B2360_ = ~new_B2383_ & new_B2384_;
  assign new_B2359_ = ~new_B2382_ | ~new_B2381_;
  assign new_B2358_ = new_B2374_ | new_B2373_;
  assign new_B2357_ = new_B2380_ | new_B2379_;
  assign new_B2356_ = new_B2370_ | new_B2372_;
  assign new_B2355_ = ~new_B2377_ | ~new_B2378_;
  assign new_B2354_ = new_B2330_ & ~new_B2331_;
  assign new_B2353_ = new_B2344_ & ~new_B2356_;
  assign new_B2352_ = ~new_B2344_ & new_B2356_;
  assign new_B2351_ = ~new_B2342_ & new_B2368_;
  assign new_B2350_ = new_B2366_ | new_B2365_;
  assign new_B2349_ = new_B2363_ | new_B2362_;
  assign new_B2348_ = new_B2331_ | new_B2364_;
  assign new_B2347_ = new_B2356_ & new_B2359_;
  assign new_B2346_ = new_B2361_ | new_B2360_;
  assign new_B2345_ = new_B2356_ & new_B2355_;
  assign new_B2344_ = new_B2358_ & new_B2357_;
  assign new_B2343_ = new_B2353_ | new_B2352_;
  assign new_B2342_ = new_B2331_ | new_B2354_;
  assign B2341 = new_B2342_ | new_B2351_;
  assign B2340 = new_B2349_ & new_B2350_;
  assign B2339 = new_B2349_ & new_B2348_;
  assign B2338 = new_B2347_ | new_B2346_;
  assign B2337 = new_B2345_ | new_B2344_;
  assign B2336 = new_B2343_ & new_B2342_;
  assign new_B2335_ = new_D4114_;
  assign new_B2334_ = new_D4047_;
  assign new_B2333_ = new_D3980_;
  assign new_B2332_ = new_D3913_;
  assign new_B2331_ = new_D3846_;
  assign new_B2330_ = new_D3779_;
  assign new_B2329_ = ~new_B2268_ & new_B2282_;
  assign new_B2328_ = new_B2268_ & ~new_B2282_;
  assign new_B2327_ = new_B2268_ & ~new_B2282_;
  assign new_B2326_ = ~new_B2268_ & ~new_B2282_;
  assign new_B2325_ = new_B2268_ & new_B2282_;
  assign new_B2324_ = new_B2328_ | new_B2329_;
  assign new_B2323_ = ~new_B2268_ & new_B2282_;
  assign new_B2322_ = new_B2326_ | new_B2327_;
  assign new_B2321_ = ~new_B2297_ & ~new_B2317_;
  assign new_B2320_ = new_B2297_ & new_B2317_;
  assign new_B2319_ = ~new_B2264_ | ~new_B2289_;
  assign new_B2318_ = new_B2282_ & new_B2319_;
  assign new_B2317_ = new_B2265_ | new_B2266_;
  assign new_B2316_ = new_B2265_ | new_B2282_;
  assign new_B2315_ = ~new_B2282_ & ~new_B2318_;
  assign new_B2314_ = new_B2282_ | new_B2319_;
  assign new_B2313_ = new_B2265_ & ~new_B2266_;
  assign new_B2312_ = ~new_B2265_ & new_B2266_;
  assign new_B2311_ = new_B2275_ | new_B2308_;
  assign new_B2310_ = ~new_B2275_ & ~new_B2309_;
  assign new_B2309_ = new_B2275_ & new_B2308_;
  assign new_B2308_ = ~new_B2264_ | ~new_B2289_;
  assign new_B2307_ = ~new_B2265_ & new_B2275_;
  assign new_B2306_ = new_B2265_ & ~new_B2275_;
  assign new_B2305_ = new_B2267_ & new_B2304_;
  assign new_B2304_ = new_B2323_ | new_B2322_;
  assign new_B2303_ = ~new_B2267_ & new_B2302_;
  assign new_B2302_ = new_B2325_ | new_B2324_;
  assign new_B2301_ = new_B2267_ | new_B2300_;
  assign new_B2300_ = new_B2321_ | new_B2320_;
  assign new_B2299_ = ~new_B2279_ & ~new_B2289_;
  assign new_B2298_ = new_B2279_ & new_B2289_;
  assign new_B2297_ = ~new_B2279_ | new_B2289_;
  assign new_B2296_ = new_B2263_ & ~new_B2264_;
  assign new_B2295_ = ~new_B2263_ & new_B2264_;
  assign new_B2294_ = new_B2316_ & ~new_B2317_;
  assign new_B2293_ = ~new_B2316_ & new_B2317_;
  assign new_B2292_ = ~new_B2315_ | ~new_B2314_;
  assign new_B2291_ = new_B2307_ | new_B2306_;
  assign new_B2290_ = new_B2313_ | new_B2312_;
  assign new_B2289_ = new_B2303_ | new_B2305_;
  assign new_B2288_ = ~new_B2310_ | ~new_B2311_;
  assign new_B2287_ = new_B2263_ & ~new_B2264_;
  assign new_B2286_ = new_B2277_ & ~new_B2289_;
  assign new_B2285_ = ~new_B2277_ & new_B2289_;
  assign new_B2284_ = ~new_B2275_ & new_B2301_;
  assign new_B2283_ = new_B2299_ | new_B2298_;
  assign new_B2282_ = new_B2296_ | new_B2295_;
  assign new_B2281_ = new_B2264_ | new_B2297_;
  assign new_B2280_ = new_B2289_ & new_B2292_;
  assign new_B2279_ = new_B2294_ | new_B2293_;
  assign new_B2278_ = new_B2289_ & new_B2288_;
  assign new_B2277_ = new_B2291_ & new_B2290_;
  assign new_B2276_ = new_B2286_ | new_B2285_;
  assign new_B2275_ = new_B2264_ | new_B2287_;
  assign B2274 = new_B2275_ | new_B2284_;
  assign B2273 = new_B2282_ & new_B2283_;
  assign B2272 = new_B2282_ & new_B2281_;
  assign B2271 = new_B2280_ | new_B2279_;
  assign B2270 = new_B2278_ | new_B2277_;
  assign B2269 = new_B2276_ & new_B2275_;
  assign new_B2268_ = new_D3712_;
  assign new_B2267_ = new_D3645_;
  assign new_B2266_ = new_D3578_;
  assign new_B2265_ = new_D3511_;
  assign new_B2264_ = new_D3444_;
  assign new_B2263_ = new_D3377_;
  assign new_B2262_ = ~new_B2201_ & new_B2215_;
  assign new_B2261_ = new_B2201_ & ~new_B2215_;
  assign new_B2260_ = new_B2201_ & ~new_B2215_;
  assign new_B2259_ = ~new_B2201_ & ~new_B2215_;
  assign new_B2258_ = new_B2201_ & new_B2215_;
  assign new_B2257_ = new_B2261_ | new_B2262_;
  assign new_B2256_ = ~new_B2201_ & new_B2215_;
  assign new_B2255_ = new_B2259_ | new_B2260_;
  assign new_B2254_ = ~new_B2230_ & ~new_B2250_;
  assign new_B2253_ = new_B2230_ & new_B2250_;
  assign new_B2252_ = ~new_B2197_ | ~new_B2222_;
  assign new_B2251_ = new_B2215_ & new_B2252_;
  assign new_B2250_ = new_B2198_ | new_B2199_;
  assign new_B2249_ = new_B2198_ | new_B2215_;
  assign new_B2248_ = ~new_B2215_ & ~new_B2251_;
  assign new_B2247_ = new_B2215_ | new_B2252_;
  assign new_B2246_ = new_B2198_ & ~new_B2199_;
  assign new_B2245_ = ~new_B2198_ & new_B2199_;
  assign new_B2244_ = new_B2208_ | new_B2241_;
  assign new_B2243_ = ~new_B2208_ & ~new_B2242_;
  assign new_B2242_ = new_B2208_ & new_B2241_;
  assign new_B2241_ = ~new_B2197_ | ~new_B2222_;
  assign new_B2240_ = ~new_B2198_ & new_B2208_;
  assign new_B2239_ = new_B2198_ & ~new_B2208_;
  assign new_B2238_ = new_B2200_ & new_B2237_;
  assign new_B2237_ = new_B2256_ | new_B2255_;
  assign new_B2236_ = ~new_B2200_ & new_B2235_;
  assign new_B2235_ = new_B2258_ | new_B2257_;
  assign new_B2234_ = new_B2200_ | new_B2233_;
  assign new_B2233_ = new_B2254_ | new_B2253_;
  assign new_B2232_ = ~new_B2212_ & ~new_B2222_;
  assign new_B2231_ = new_B2212_ & new_B2222_;
  assign new_B2230_ = ~new_B2212_ | new_B2222_;
  assign new_B2229_ = new_B2196_ & ~new_B2197_;
  assign new_B2228_ = ~new_B2196_ & new_B2197_;
  assign new_B2227_ = new_B2249_ & ~new_B2250_;
  assign new_B2226_ = ~new_B2249_ & new_B2250_;
  assign new_B2225_ = ~new_B2248_ | ~new_B2247_;
  assign new_B2224_ = new_B2240_ | new_B2239_;
  assign new_B2223_ = new_B2246_ | new_B2245_;
  assign new_B2222_ = new_B2236_ | new_B2238_;
  assign new_B2221_ = ~new_B2243_ | ~new_B2244_;
  assign new_B2220_ = new_B2196_ & ~new_B2197_;
  assign new_B2219_ = new_B2210_ & ~new_B2222_;
  assign new_B2218_ = ~new_B2210_ & new_B2222_;
  assign new_B2217_ = ~new_B2208_ & new_B2234_;
  assign new_B2216_ = new_B2232_ | new_B2231_;
  assign new_B2215_ = new_B2229_ | new_B2228_;
  assign new_B2214_ = new_B2197_ | new_B2230_;
  assign new_B2213_ = new_B2222_ & new_B2225_;
  assign new_B2212_ = new_B2227_ | new_B2226_;
  assign new_B2211_ = new_B2222_ & new_B2221_;
  assign new_B2210_ = new_B2224_ & new_B2223_;
  assign new_B2209_ = new_B2219_ | new_B2218_;
  assign new_B2208_ = new_B2197_ | new_B2220_;
  assign B2207 = new_B2208_ | new_B2217_;
  assign B2206 = new_B2215_ & new_B2216_;
  assign B2205 = new_B2215_ & new_B2214_;
  assign B2204 = new_B2213_ | new_B2212_;
  assign B2203 = new_B2211_ | new_B2210_;
  assign B2202 = new_B2209_ & new_B2208_;
  assign new_B2201_ = new_D3310_;
  assign new_B2200_ = new_D3243_;
  assign new_B2199_ = new_D3176_;
  assign new_B2198_ = new_D3109_;
  assign new_B2197_ = new_D3042_;
  assign new_B2196_ = new_D2975_;
  assign new_B2195_ = ~new_B2134_ & new_B2148_;
  assign new_B2194_ = new_B2134_ & ~new_B2148_;
  assign new_B2193_ = new_B2134_ & ~new_B2148_;
  assign new_B2192_ = ~new_B2134_ & ~new_B2148_;
  assign new_B2191_ = new_B2134_ & new_B2148_;
  assign new_B2190_ = new_B2194_ | new_B2195_;
  assign new_B2189_ = ~new_B2134_ & new_B2148_;
  assign new_B2188_ = new_B2192_ | new_B2193_;
  assign new_B2187_ = ~new_B2163_ & ~new_B2183_;
  assign new_B2186_ = new_B2163_ & new_B2183_;
  assign new_B2185_ = ~new_B2130_ | ~new_B2155_;
  assign new_B2184_ = new_B2148_ & new_B2185_;
  assign new_B2183_ = new_B2131_ | new_B2132_;
  assign new_B2182_ = new_B2131_ | new_B2148_;
  assign new_B2181_ = ~new_B2148_ & ~new_B2184_;
  assign new_B2180_ = new_B2148_ | new_B2185_;
  assign new_B2179_ = new_B2131_ & ~new_B2132_;
  assign new_B2178_ = ~new_B2131_ & new_B2132_;
  assign new_B2177_ = new_B2141_ | new_B2174_;
  assign new_B2176_ = ~new_B2141_ & ~new_B2175_;
  assign new_B2175_ = new_B2141_ & new_B2174_;
  assign new_B2174_ = ~new_B2130_ | ~new_B2155_;
  assign new_B2173_ = ~new_B2131_ & new_B2141_;
  assign new_B2172_ = new_B2131_ & ~new_B2141_;
  assign new_B2171_ = new_B2133_ & new_B2170_;
  assign new_B2170_ = new_B2189_ | new_B2188_;
  assign new_B2169_ = ~new_B2133_ & new_B2168_;
  assign new_B2168_ = new_B2191_ | new_B2190_;
  assign new_B2167_ = new_B2133_ | new_B2166_;
  assign new_B2166_ = new_B2187_ | new_B2186_;
  assign new_B2165_ = ~new_B2145_ & ~new_B2155_;
  assign new_B2164_ = new_B2145_ & new_B2155_;
  assign new_B2163_ = ~new_B2145_ | new_B2155_;
  assign new_B2162_ = new_B2129_ & ~new_B2130_;
  assign new_B2161_ = ~new_B2129_ & new_B2130_;
  assign new_B2160_ = new_B2182_ & ~new_B2183_;
  assign new_B2159_ = ~new_B2182_ & new_B2183_;
  assign new_B2158_ = ~new_B2181_ | ~new_B2180_;
  assign new_B2157_ = new_B2173_ | new_B2172_;
  assign new_B2156_ = new_B2179_ | new_B2178_;
  assign new_B2155_ = new_B2169_ | new_B2171_;
  assign new_B2154_ = ~new_B2176_ | ~new_B2177_;
  assign new_B2153_ = new_B2129_ & ~new_B2130_;
  assign new_B2152_ = new_B2143_ & ~new_B2155_;
  assign new_B2151_ = ~new_B2143_ & new_B2155_;
  assign new_B2150_ = ~new_B2141_ & new_B2167_;
  assign new_B2149_ = new_B2165_ | new_B2164_;
  assign new_B2148_ = new_B2162_ | new_B2161_;
  assign new_B2147_ = new_B2130_ | new_B2163_;
  assign new_B2146_ = new_B2155_ & new_B2158_;
  assign new_B2145_ = new_B2160_ | new_B2159_;
  assign new_B2144_ = new_B2155_ & new_B2154_;
  assign new_B2143_ = new_B2157_ & new_B2156_;
  assign new_B2142_ = new_B2152_ | new_B2151_;
  assign new_B2141_ = new_B2130_ | new_B2153_;
  assign B2140 = new_B2141_ | new_B2150_;
  assign B2139 = new_B2148_ & new_B2149_;
  assign B2138 = new_B2148_ & new_B2147_;
  assign B2137 = new_B2146_ | new_B2145_;
  assign B2136 = new_B2144_ | new_B2143_;
  assign B2135 = new_B2142_ & new_B2141_;
  assign new_B2134_ = new_D2908_;
  assign new_B2133_ = new_D2841_;
  assign new_B2132_ = new_D2774_;
  assign new_B2131_ = new_D2707_;
  assign new_B2130_ = new_D2640_;
  assign new_B2129_ = new_D2573_;
  assign new_B2128_ = ~new_B2067_ & new_B2081_;
  assign new_B2127_ = new_B2067_ & ~new_B2081_;
  assign new_B2126_ = new_B2067_ & ~new_B2081_;
  assign new_B2125_ = ~new_B2067_ & ~new_B2081_;
  assign new_B2124_ = new_B2067_ & new_B2081_;
  assign new_B2123_ = new_B2127_ | new_B2128_;
  assign new_B2122_ = ~new_B2067_ & new_B2081_;
  assign new_B2121_ = new_B2125_ | new_B2126_;
  assign new_B2120_ = ~new_B2096_ & ~new_B2116_;
  assign new_B2119_ = new_B2096_ & new_B2116_;
  assign new_B2118_ = ~new_B2063_ | ~new_B2088_;
  assign new_B2117_ = new_B2081_ & new_B2118_;
  assign new_B2116_ = new_B2064_ | new_B2065_;
  assign new_B2115_ = new_B2064_ | new_B2081_;
  assign new_B2114_ = ~new_B2081_ & ~new_B2117_;
  assign new_B2113_ = new_B2081_ | new_B2118_;
  assign new_B2112_ = new_B2064_ & ~new_B2065_;
  assign new_B2111_ = ~new_B2064_ & new_B2065_;
  assign new_B2110_ = new_B2074_ | new_B2107_;
  assign new_B2109_ = ~new_B2074_ & ~new_B2108_;
  assign new_B2108_ = new_B2074_ & new_B2107_;
  assign new_B2107_ = ~new_B2063_ | ~new_B2088_;
  assign new_B2106_ = ~new_B2064_ & new_B2074_;
  assign new_B2105_ = new_B2064_ & ~new_B2074_;
  assign new_B2104_ = new_B2066_ & new_B2103_;
  assign new_B2103_ = new_B2122_ | new_B2121_;
  assign new_B2102_ = ~new_B2066_ & new_B2101_;
  assign new_B2101_ = new_B2124_ | new_B2123_;
  assign new_B2100_ = new_B2066_ | new_B2099_;
  assign new_B2099_ = new_B2120_ | new_B2119_;
  assign new_B2098_ = ~new_B2078_ & ~new_B2088_;
  assign new_B2097_ = new_B2078_ & new_B2088_;
  assign new_B2096_ = ~new_B2078_ | new_B2088_;
  assign new_B2095_ = new_B2062_ & ~new_B2063_;
  assign new_B2094_ = ~new_B2062_ & new_B2063_;
  assign new_B2093_ = new_B2115_ & ~new_B2116_;
  assign new_B2092_ = ~new_B2115_ & new_B2116_;
  assign new_B2091_ = ~new_B2114_ | ~new_B2113_;
  assign new_B2090_ = new_B2106_ | new_B2105_;
  assign new_B2089_ = new_B2112_ | new_B2111_;
  assign new_B2088_ = new_B2102_ | new_B2104_;
  assign new_B2087_ = ~new_B2109_ | ~new_B2110_;
  assign new_B2086_ = new_B2062_ & ~new_B2063_;
  assign new_B2085_ = new_B2076_ & ~new_B2088_;
  assign new_B2084_ = ~new_B2076_ & new_B2088_;
  assign new_B2083_ = ~new_B2074_ & new_B2100_;
  assign new_B2082_ = new_B2098_ | new_B2097_;
  assign new_B2081_ = new_B2095_ | new_B2094_;
  assign new_B2080_ = new_B2063_ | new_B2096_;
  assign new_B2079_ = new_B2088_ & new_B2091_;
  assign new_B2078_ = new_B2093_ | new_B2092_;
  assign new_B2077_ = new_B2088_ & new_B2087_;
  assign new_B2076_ = new_B2090_ & new_B2089_;
  assign new_B2075_ = new_B2085_ | new_B2084_;
  assign new_B2074_ = new_B2063_ | new_B2086_;
  assign B2073 = new_B2074_ | new_B2083_;
  assign B2072 = new_B2081_ & new_B2082_;
  assign B2071 = new_B2081_ & new_B2080_;
  assign B2070 = new_B2079_ | new_B2078_;
  assign B2069 = new_B2077_ | new_B2076_;
  assign B2068 = new_B2075_ & new_B2074_;
  assign new_B2067_ = new_D2506_;
  assign new_B2066_ = new_D2439_;
  assign new_B2065_ = new_D2372_;
  assign new_B2064_ = new_D2305_;
  assign new_B2063_ = new_D2238_;
  assign new_B2062_ = new_D2171_;
  assign new_B2061_ = ~new_B2000_ & new_B2014_;
  assign new_B2060_ = new_B2000_ & ~new_B2014_;
  assign new_B2059_ = new_B2000_ & ~new_B2014_;
  assign new_B2058_ = ~new_B2000_ & ~new_B2014_;
  assign new_B2057_ = new_B2000_ & new_B2014_;
  assign new_B2056_ = new_B2060_ | new_B2061_;
  assign new_B2055_ = ~new_B2000_ & new_B2014_;
  assign new_B2054_ = new_B2058_ | new_B2059_;
  assign new_B2053_ = ~new_B2029_ & ~new_B2049_;
  assign new_B2052_ = new_B2029_ & new_B2049_;
  assign new_B2051_ = ~new_B1996_ | ~new_B2021_;
  assign new_B2050_ = new_B2014_ & new_B2051_;
  assign new_B2049_ = new_B1997_ | new_B1998_;
  assign new_B2048_ = new_B1997_ | new_B2014_;
  assign new_B2047_ = ~new_B2014_ & ~new_B2050_;
  assign new_B2046_ = new_B2014_ | new_B2051_;
  assign new_B2045_ = new_B1997_ & ~new_B1998_;
  assign new_B2044_ = ~new_B1997_ & new_B1998_;
  assign new_B2043_ = new_B2007_ | new_B2040_;
  assign new_B2042_ = ~new_B2007_ & ~new_B2041_;
  assign new_B2041_ = new_B2007_ & new_B2040_;
  assign new_B2040_ = ~new_B1996_ | ~new_B2021_;
  assign new_B2039_ = ~new_B1997_ & new_B2007_;
  assign new_B2038_ = new_B1997_ & ~new_B2007_;
  assign new_B2037_ = new_B1999_ & new_B2036_;
  assign new_B2036_ = new_B2055_ | new_B2054_;
  assign new_B2035_ = ~new_B1999_ & new_B2034_;
  assign new_B2034_ = new_B2057_ | new_B2056_;
  assign new_B2033_ = new_B1999_ | new_B2032_;
  assign new_B2032_ = new_B2053_ | new_B2052_;
  assign new_B2031_ = ~new_B2011_ & ~new_B2021_;
  assign new_B2030_ = new_B2011_ & new_B2021_;
  assign new_B2029_ = ~new_B2011_ | new_B2021_;
  assign new_B2028_ = new_B1995_ & ~new_B1996_;
  assign new_B2027_ = ~new_B1995_ & new_B1996_;
  assign new_B2026_ = new_B2048_ & ~new_B2049_;
  assign new_B2025_ = ~new_B2048_ & new_B2049_;
  assign new_B2024_ = ~new_B2047_ | ~new_B2046_;
  assign new_B2023_ = new_B2039_ | new_B2038_;
  assign new_B2022_ = new_B2045_ | new_B2044_;
  assign new_B2021_ = new_B2035_ | new_B2037_;
  assign new_B2020_ = ~new_B2042_ | ~new_B2043_;
  assign new_B2019_ = new_B1995_ & ~new_B1996_;
  assign new_B2018_ = new_B2009_ & ~new_B2021_;
  assign new_B2017_ = ~new_B2009_ & new_B2021_;
  assign new_B2016_ = ~new_B2007_ & new_B2033_;
  assign new_B2015_ = new_B2031_ | new_B2030_;
  assign new_B2014_ = new_B2028_ | new_B2027_;
  assign new_B2013_ = new_B1996_ | new_B2029_;
  assign new_B2012_ = new_B2021_ & new_B2024_;
  assign new_B2011_ = new_B2026_ | new_B2025_;
  assign new_B2010_ = new_B2021_ & new_B2020_;
  assign new_B2009_ = new_B2023_ & new_B2022_;
  assign new_B2008_ = new_B2018_ | new_B2017_;
  assign new_B2007_ = new_B1996_ | new_B2019_;
  assign B2006 = new_B2007_ | new_B2016_;
  assign B2005 = new_B2014_ & new_B2015_;
  assign B2004 = new_B2014_ & new_B2013_;
  assign B2003 = new_B2012_ | new_B2011_;
  assign B2002 = new_B2010_ | new_B2009_;
  assign B2001 = new_B2008_ & new_B2007_;
  assign new_B2000_ = new_D2104_;
  assign new_B1999_ = new_D2037_;
  assign new_B1998_ = new_D1970_;
  assign new_B1997_ = new_D1903_;
  assign new_B1996_ = new_D1836_;
  assign new_B1995_ = new_D1769_;
  assign new_B1994_ = ~new_B1933_ & new_B1947_;
  assign new_B1993_ = new_B1933_ & ~new_B1947_;
  assign new_B1992_ = new_B1933_ & ~new_B1947_;
  assign new_B1991_ = ~new_B1933_ & ~new_B1947_;
  assign new_B1990_ = new_B1933_ & new_B1947_;
  assign new_B1989_ = new_B1993_ | new_B1994_;
  assign new_B1988_ = ~new_B1933_ & new_B1947_;
  assign new_B1987_ = new_B1991_ | new_B1992_;
  assign new_B1986_ = ~new_B1962_ & ~new_B1982_;
  assign new_B1985_ = new_B1962_ & new_B1982_;
  assign new_B1984_ = ~new_B1929_ | ~new_B1954_;
  assign new_B1983_ = new_B1947_ & new_B1984_;
  assign new_B1982_ = new_B1930_ | new_B1931_;
  assign new_B1981_ = new_B1930_ | new_B1947_;
  assign new_B1980_ = ~new_B1947_ & ~new_B1983_;
  assign new_B1979_ = new_B1947_ | new_B1984_;
  assign new_B1978_ = new_B1930_ & ~new_B1931_;
  assign new_B1977_ = ~new_B1930_ & new_B1931_;
  assign new_B1976_ = new_B1940_ | new_B1973_;
  assign new_B1975_ = ~new_B1940_ & ~new_B1974_;
  assign new_B1974_ = new_B1940_ & new_B1973_;
  assign new_B1973_ = ~new_B1929_ | ~new_B1954_;
  assign new_B1972_ = ~new_B1930_ & new_B1940_;
  assign new_B1971_ = new_B1930_ & ~new_B1940_;
  assign new_B1970_ = new_B1932_ & new_B1969_;
  assign new_B1969_ = new_B1988_ | new_B1987_;
  assign new_B1968_ = ~new_B1932_ & new_B1967_;
  assign new_B1967_ = new_B1990_ | new_B1989_;
  assign new_B1966_ = new_B1932_ | new_B1965_;
  assign new_B1965_ = new_B1986_ | new_B1985_;
  assign new_B1964_ = ~new_B1944_ & ~new_B1954_;
  assign new_B1963_ = new_B1944_ & new_B1954_;
  assign new_B1962_ = ~new_B1944_ | new_B1954_;
  assign new_B1961_ = new_B1928_ & ~new_B1929_;
  assign new_B1960_ = ~new_B1928_ & new_B1929_;
  assign new_B1959_ = new_B1981_ & ~new_B1982_;
  assign new_B1958_ = ~new_B1981_ & new_B1982_;
  assign new_B1957_ = ~new_B1980_ | ~new_B1979_;
  assign new_B1956_ = new_B1972_ | new_B1971_;
  assign new_B1955_ = new_B1978_ | new_B1977_;
  assign new_B1954_ = new_B1968_ | new_B1970_;
  assign new_B1953_ = ~new_B1975_ | ~new_B1976_;
  assign new_B1952_ = new_B1928_ & ~new_B1929_;
  assign new_B1951_ = new_B1942_ & ~new_B1954_;
  assign new_B1950_ = ~new_B1942_ & new_B1954_;
  assign new_B1949_ = ~new_B1940_ & new_B1966_;
  assign new_B1948_ = new_B1964_ | new_B1963_;
  assign new_B1947_ = new_B1961_ | new_B1960_;
  assign new_B1946_ = new_B1929_ | new_B1962_;
  assign new_B1945_ = new_B1954_ & new_B1957_;
  assign new_B1944_ = new_B1959_ | new_B1958_;
  assign new_B1943_ = new_B1954_ & new_B1953_;
  assign new_B1942_ = new_B1956_ & new_B1955_;
  assign new_B1941_ = new_B1951_ | new_B1950_;
  assign new_B1940_ = new_B1929_ | new_B1952_;
  assign B1939 = new_B1940_ | new_B1949_;
  assign B1938 = new_B1947_ & new_B1948_;
  assign B1937 = new_B1947_ & new_B1946_;
  assign B1936 = new_B1945_ | new_B1944_;
  assign B1935 = new_B1943_ | new_B1942_;
  assign B1934 = new_B1941_ & new_B1940_;
  assign new_B1933_ = new_D1702_;
  assign new_B1932_ = new_D1635_;
  assign new_B1931_ = new_D1568_;
  assign new_B1930_ = new_D1501_;
  assign new_B1929_ = new_D1434_;
  assign new_B1928_ = new_D1367_;
  assign new_B1927_ = ~new_B1866_ & new_B1880_;
  assign new_B1926_ = new_B1866_ & ~new_B1880_;
  assign new_B1925_ = new_B1866_ & ~new_B1880_;
  assign new_B1924_ = ~new_B1866_ & ~new_B1880_;
  assign new_B1923_ = new_B1866_ & new_B1880_;
  assign new_B1922_ = new_B1926_ | new_B1927_;
  assign new_B1921_ = ~new_B1866_ & new_B1880_;
  assign new_B1920_ = new_B1924_ | new_B1925_;
  assign new_B1919_ = ~new_B1895_ & ~new_B1915_;
  assign new_B1918_ = new_B1895_ & new_B1915_;
  assign new_B1917_ = ~new_B1862_ | ~new_B1887_;
  assign new_B1916_ = new_B1880_ & new_B1917_;
  assign new_B1915_ = new_B1863_ | new_B1864_;
  assign new_B1914_ = new_B1863_ | new_B1880_;
  assign new_B1913_ = ~new_B1880_ & ~new_B1916_;
  assign new_B1912_ = new_B1880_ | new_B1917_;
  assign new_B1911_ = new_B1863_ & ~new_B1864_;
  assign new_B1910_ = ~new_B1863_ & new_B1864_;
  assign new_B1909_ = new_B1873_ | new_B1906_;
  assign new_B1908_ = ~new_B1873_ & ~new_B1907_;
  assign new_B1907_ = new_B1873_ & new_B1906_;
  assign new_B1906_ = ~new_B1862_ | ~new_B1887_;
  assign new_B1905_ = ~new_B1863_ & new_B1873_;
  assign new_B1904_ = new_B1863_ & ~new_B1873_;
  assign new_B1903_ = new_B1865_ & new_B1902_;
  assign new_B1902_ = new_B1921_ | new_B1920_;
  assign new_B1901_ = ~new_B1865_ & new_B1900_;
  assign new_B1900_ = new_B1923_ | new_B1922_;
  assign new_B1899_ = new_B1865_ | new_B1898_;
  assign new_B1898_ = new_B1919_ | new_B1918_;
  assign new_B1897_ = ~new_B1877_ & ~new_B1887_;
  assign new_B1896_ = new_B1877_ & new_B1887_;
  assign new_B1895_ = ~new_B1877_ | new_B1887_;
  assign new_B1894_ = new_B1861_ & ~new_B1862_;
  assign new_B1893_ = ~new_B1861_ & new_B1862_;
  assign new_B1892_ = new_B1914_ & ~new_B1915_;
  assign new_B1891_ = ~new_B1914_ & new_B1915_;
  assign new_B1890_ = ~new_B1913_ | ~new_B1912_;
  assign new_B1889_ = new_B1905_ | new_B1904_;
  assign new_B1888_ = new_B1911_ | new_B1910_;
  assign new_B1887_ = new_B1901_ | new_B1903_;
  assign new_B1886_ = ~new_B1908_ | ~new_B1909_;
  assign new_B1885_ = new_B1861_ & ~new_B1862_;
  assign new_B1884_ = new_B1875_ & ~new_B1887_;
  assign new_B1883_ = ~new_B1875_ & new_B1887_;
  assign new_B1882_ = ~new_B1873_ & new_B1899_;
  assign new_B1881_ = new_B1897_ | new_B1896_;
  assign new_B1880_ = new_B1894_ | new_B1893_;
  assign new_B1879_ = new_B1862_ | new_B1895_;
  assign new_B1878_ = new_B1887_ & new_B1890_;
  assign new_B1877_ = new_B1892_ | new_B1891_;
  assign new_B1876_ = new_B1887_ & new_B1886_;
  assign new_B1875_ = new_B1889_ & new_B1888_;
  assign new_B1874_ = new_B1884_ | new_B1883_;
  assign new_B1873_ = new_B1862_ | new_B1885_;
  assign B1872 = new_B1873_ | new_B1882_;
  assign B1871 = new_B1880_ & new_B1881_;
  assign B1870 = new_B1880_ & new_B1879_;
  assign B1869 = new_B1878_ | new_B1877_;
  assign B1868 = new_B1876_ | new_B1875_;
  assign B1867 = new_B1874_ & new_B1873_;
  assign new_B1866_ = new_D1300_;
  assign new_B1865_ = new_D1233_;
  assign new_B1864_ = new_D1166_;
  assign new_B1863_ = new_D1099_;
  assign new_B1862_ = new_D1032_;
  assign new_B1861_ = new_D965_;
  assign new_B1860_ = ~new_B1799_ & new_B1813_;
  assign new_B1859_ = new_B1799_ & ~new_B1813_;
  assign new_B1858_ = new_B1799_ & ~new_B1813_;
  assign new_B1857_ = ~new_B1799_ & ~new_B1813_;
  assign new_B1856_ = new_B1799_ & new_B1813_;
  assign new_B1855_ = new_B1859_ | new_B1860_;
  assign new_B1854_ = ~new_B1799_ & new_B1813_;
  assign new_B1853_ = new_B1857_ | new_B1858_;
  assign new_B1852_ = ~new_B1828_ & ~new_B1848_;
  assign new_B1851_ = new_B1828_ & new_B1848_;
  assign new_B1850_ = ~new_B1795_ | ~new_B1820_;
  assign new_B1849_ = new_B1813_ & new_B1850_;
  assign new_B1848_ = new_B1796_ | new_B1797_;
  assign new_B1847_ = new_B1796_ | new_B1813_;
  assign new_B1846_ = ~new_B1813_ & ~new_B1849_;
  assign new_B1845_ = new_B1813_ | new_B1850_;
  assign new_B1844_ = new_B1796_ & ~new_B1797_;
  assign new_B1843_ = ~new_B1796_ & new_B1797_;
  assign new_B1842_ = new_B1806_ | new_B1839_;
  assign new_B1841_ = ~new_B1806_ & ~new_B1840_;
  assign new_B1840_ = new_B1806_ & new_B1839_;
  assign new_B1839_ = ~new_B1795_ | ~new_B1820_;
  assign new_B1838_ = ~new_B1796_ & new_B1806_;
  assign new_B1837_ = new_B1796_ & ~new_B1806_;
  assign new_B1836_ = new_B1798_ & new_B1835_;
  assign new_B1835_ = new_B1854_ | new_B1853_;
  assign new_B1834_ = ~new_B1798_ & new_B1833_;
  assign new_B1833_ = new_B1856_ | new_B1855_;
  assign new_B1832_ = new_B1798_ | new_B1831_;
  assign new_B1831_ = new_B1852_ | new_B1851_;
  assign new_B1830_ = ~new_B1810_ & ~new_B1820_;
  assign new_B1829_ = new_B1810_ & new_B1820_;
  assign new_B1828_ = ~new_B1810_ | new_B1820_;
  assign new_B1827_ = new_B1794_ & ~new_B1795_;
  assign new_B1826_ = ~new_B1794_ & new_B1795_;
  assign new_B1825_ = new_B1847_ & ~new_B1848_;
  assign new_B1824_ = ~new_B1847_ & new_B1848_;
  assign new_B1823_ = ~new_B1846_ | ~new_B1845_;
  assign new_B1822_ = new_B1838_ | new_B1837_;
  assign new_B1821_ = new_B1844_ | new_B1843_;
  assign new_B1820_ = new_B1834_ | new_B1836_;
  assign new_B1819_ = ~new_B1841_ | ~new_B1842_;
  assign new_B1818_ = new_B1794_ & ~new_B1795_;
  assign new_B1817_ = new_B1808_ & ~new_B1820_;
  assign new_B1816_ = ~new_B1808_ & new_B1820_;
  assign new_B1815_ = ~new_B1806_ & new_B1832_;
  assign new_B1814_ = new_B1830_ | new_B1829_;
  assign new_B1813_ = new_B1827_ | new_B1826_;
  assign new_B1812_ = new_B1795_ | new_B1828_;
  assign new_B1811_ = new_B1820_ & new_B1823_;
  assign new_B1810_ = new_B1825_ | new_B1824_;
  assign new_B1809_ = new_B1820_ & new_B1819_;
  assign new_B1808_ = new_B1822_ & new_B1821_;
  assign new_B1807_ = new_B1817_ | new_B1816_;
  assign new_B1806_ = new_B1795_ | new_B1818_;
  assign B1805 = new_B1806_ | new_B1815_;
  assign B1804 = new_B1813_ & new_B1814_;
  assign B1803 = new_B1813_ & new_B1812_;
  assign B1802 = new_B1811_ | new_B1810_;
  assign B1801 = new_B1809_ | new_B1808_;
  assign B1800 = new_B1807_ & new_B1806_;
  assign new_B1799_ = new_D898_;
  assign new_B1798_ = new_D831_;
  assign new_B1797_ = new_D764_;
  assign new_B1796_ = new_D697_;
  assign new_B1795_ = new_D630_;
  assign new_B1794_ = new_D563_;
  assign new_B1793_ = ~new_B1732_ & new_B1746_;
  assign new_B1792_ = new_B1732_ & ~new_B1746_;
  assign new_B1791_ = new_B1732_ & ~new_B1746_;
  assign new_B1790_ = ~new_B1732_ & ~new_B1746_;
  assign new_B1789_ = new_B1732_ & new_B1746_;
  assign new_B1788_ = new_B1792_ | new_B1793_;
  assign new_B1787_ = ~new_B1732_ & new_B1746_;
  assign new_B1786_ = new_B1790_ | new_B1791_;
  assign new_B1785_ = ~new_B1761_ & ~new_B1781_;
  assign new_B1784_ = new_B1761_ & new_B1781_;
  assign new_B1783_ = ~new_B1728_ | ~new_B1753_;
  assign new_B1782_ = new_B1746_ & new_B1783_;
  assign new_B1781_ = new_B1729_ | new_B1730_;
  assign new_B1780_ = new_B1729_ | new_B1746_;
  assign new_B1779_ = ~new_B1746_ & ~new_B1782_;
  assign new_B1778_ = new_B1746_ | new_B1783_;
  assign new_B1777_ = new_B1729_ & ~new_B1730_;
  assign new_B1776_ = ~new_B1729_ & new_B1730_;
  assign new_B1775_ = new_B1739_ | new_B1772_;
  assign new_B1774_ = ~new_B1739_ & ~new_B1773_;
  assign new_B1773_ = new_B1739_ & new_B1772_;
  assign new_B1772_ = ~new_B1728_ | ~new_B1753_;
  assign new_B1771_ = ~new_B1729_ & new_B1739_;
  assign new_B1770_ = new_B1729_ & ~new_B1739_;
  assign new_B1769_ = new_B1731_ & new_B1768_;
  assign new_B1768_ = new_B1787_ | new_B1786_;
  assign new_B1767_ = ~new_B1731_ & new_B1766_;
  assign new_B1766_ = new_B1789_ | new_B1788_;
  assign new_B1765_ = new_B1731_ | new_B1764_;
  assign new_B1764_ = new_B1785_ | new_B1784_;
  assign new_B1763_ = ~new_B1743_ & ~new_B1753_;
  assign new_B1762_ = new_B1743_ & new_B1753_;
  assign new_B1761_ = ~new_B1743_ | new_B1753_;
  assign new_B1760_ = new_B1727_ & ~new_B1728_;
  assign new_B1759_ = ~new_B1727_ & new_B1728_;
  assign new_B1758_ = new_B1780_ & ~new_B1781_;
  assign new_B1757_ = ~new_B1780_ & new_B1781_;
  assign new_B1756_ = ~new_B1779_ | ~new_B1778_;
  assign new_B1755_ = new_B1771_ | new_B1770_;
  assign new_B1754_ = new_B1777_ | new_B1776_;
  assign new_B1753_ = new_B1767_ | new_B1769_;
  assign new_B1752_ = ~new_B1774_ | ~new_B1775_;
  assign new_B1751_ = new_B1727_ & ~new_B1728_;
  assign new_B1750_ = new_B1741_ & ~new_B1753_;
  assign new_B1749_ = ~new_B1741_ & new_B1753_;
  assign new_B1748_ = ~new_B1739_ & new_B1765_;
  assign new_B1747_ = new_B1763_ | new_B1762_;
  assign new_B1746_ = new_B1760_ | new_B1759_;
  assign new_B1745_ = new_B1728_ | new_B1761_;
  assign new_B1744_ = new_B1753_ & new_B1756_;
  assign new_B1743_ = new_B1758_ | new_B1757_;
  assign new_B1742_ = new_B1753_ & new_B1752_;
  assign new_B1741_ = new_B1755_ & new_B1754_;
  assign new_B1740_ = new_B1750_ | new_B1749_;
  assign new_B1739_ = new_B1728_ | new_B1751_;
  assign B1738 = new_B1739_ | new_B1748_;
  assign B1737 = new_B1746_ & new_B1747_;
  assign B1736 = new_B1746_ & new_B1745_;
  assign B1735 = new_B1744_ | new_B1743_;
  assign B1734 = new_B1742_ | new_B1741_;
  assign B1733 = new_B1740_ & new_B1739_;
  assign new_B1732_ = new_D496_;
  assign new_B1731_ = new_D429_;
  assign new_B1730_ = new_D362_;
  assign new_B1729_ = new_D295_;
  assign new_B1728_ = new_D228_;
  assign new_B1727_ = new_D161_;
  assign new_B1726_ = ~new_B1665_ & new_B1679_;
  assign new_B1725_ = new_B1665_ & ~new_B1679_;
  assign new_B1724_ = new_B1665_ & ~new_B1679_;
  assign new_B1723_ = ~new_B1665_ & ~new_B1679_;
  assign new_B1722_ = new_B1665_ & new_B1679_;
  assign new_B1721_ = new_B1725_ | new_B1726_;
  assign new_B1720_ = ~new_B1665_ & new_B1679_;
  assign new_B1719_ = new_B1723_ | new_B1724_;
  assign new_B1718_ = ~new_B1694_ & ~new_B1714_;
  assign new_B1717_ = new_B1694_ & new_B1714_;
  assign new_B1716_ = ~new_B1661_ | ~new_B1686_;
  assign new_B1715_ = new_B1679_ & new_B1716_;
  assign new_B1714_ = new_B1662_ | new_B1663_;
  assign new_B1713_ = new_B1662_ | new_B1679_;
  assign new_B1712_ = ~new_B1679_ & ~new_B1715_;
  assign new_B1711_ = new_B1679_ | new_B1716_;
  assign new_B1710_ = new_B1662_ & ~new_B1663_;
  assign new_B1709_ = ~new_B1662_ & new_B1663_;
  assign new_B1708_ = new_B1672_ | new_B1705_;
  assign new_B1707_ = ~new_B1672_ & ~new_B1706_;
  assign new_B1706_ = new_B1672_ & new_B1705_;
  assign new_B1705_ = ~new_B1661_ | ~new_B1686_;
  assign new_B1704_ = ~new_B1662_ & new_B1672_;
  assign new_B1703_ = new_B1662_ & ~new_B1672_;
  assign new_B1702_ = new_B1664_ & new_B1701_;
  assign new_B1701_ = new_B1720_ | new_B1719_;
  assign new_B1700_ = ~new_B1664_ & new_B1699_;
  assign new_B1699_ = new_B1722_ | new_B1721_;
  assign new_B1698_ = new_B1664_ | new_B1697_;
  assign new_B1697_ = new_B1718_ | new_B1717_;
  assign new_B1696_ = ~new_B1676_ & ~new_B1686_;
  assign new_B1695_ = new_B1676_ & new_B1686_;
  assign new_B1694_ = ~new_B1676_ | new_B1686_;
  assign new_B1693_ = new_B1660_ & ~new_B1661_;
  assign new_B1692_ = ~new_B1660_ & new_B1661_;
  assign new_B1691_ = new_B1713_ & ~new_B1714_;
  assign new_B1690_ = ~new_B1713_ & new_B1714_;
  assign new_B1689_ = ~new_B1712_ | ~new_B1711_;
  assign new_B1688_ = new_B1704_ | new_B1703_;
  assign new_B1687_ = new_B1710_ | new_B1709_;
  assign new_B1686_ = new_B1700_ | new_B1702_;
  assign new_B1685_ = ~new_B1707_ | ~new_B1708_;
  assign new_B1684_ = new_B1660_ & ~new_B1661_;
  assign new_B1683_ = new_B1674_ & ~new_B1686_;
  assign new_B1682_ = ~new_B1674_ & new_B1686_;
  assign new_B1681_ = ~new_B1672_ & new_B1698_;
  assign new_B1680_ = new_B1696_ | new_B1695_;
  assign new_B1679_ = new_B1693_ | new_B1692_;
  assign new_B1678_ = new_B1661_ | new_B1694_;
  assign new_B1677_ = new_B1686_ & new_B1689_;
  assign new_B1676_ = new_B1691_ | new_B1690_;
  assign new_B1675_ = new_B1686_ & new_B1685_;
  assign new_B1674_ = new_B1688_ & new_B1687_;
  assign new_B1673_ = new_B1683_ | new_B1682_;
  assign new_B1672_ = new_B1661_ | new_B1684_;
  assign B1671 = new_B1672_ | new_B1681_;
  assign B1670 = new_B1679_ & new_B1680_;
  assign B1669 = new_B1679_ & new_B1678_;
  assign B1668 = new_B1677_ | new_B1676_;
  assign B1667 = new_B1675_ | new_B1674_;
  assign B1666 = new_B1673_ & new_B1672_;
  assign new_B1665_ = new_D94_;
  assign new_B1664_ = new_D27_;
  assign new_B1663_ = new_C9959_;
  assign new_B1662_ = new_C9892_;
  assign new_B1661_ = new_C9825_;
  assign new_B1660_ = new_C9758_;
  assign new_B1659_ = ~new_B1598_ & new_B1612_;
  assign new_B1658_ = new_B1598_ & ~new_B1612_;
  assign new_B1657_ = new_B1598_ & ~new_B1612_;
  assign new_B1656_ = ~new_B1598_ & ~new_B1612_;
  assign new_B1655_ = new_B1598_ & new_B1612_;
  assign new_B1654_ = new_B1658_ | new_B1659_;
  assign new_B1653_ = ~new_B1598_ & new_B1612_;
  assign new_B1652_ = new_B1656_ | new_B1657_;
  assign new_B1651_ = ~new_B1627_ & ~new_B1647_;
  assign new_B1650_ = new_B1627_ & new_B1647_;
  assign new_B1649_ = ~new_B1594_ | ~new_B1619_;
  assign new_B1648_ = new_B1612_ & new_B1649_;
  assign new_B1647_ = new_B1595_ | new_B1596_;
  assign new_B1646_ = new_B1595_ | new_B1612_;
  assign new_B1645_ = ~new_B1612_ & ~new_B1648_;
  assign new_B1644_ = new_B1612_ | new_B1649_;
  assign new_B1643_ = new_B1595_ & ~new_B1596_;
  assign new_B1642_ = ~new_B1595_ & new_B1596_;
  assign new_B1641_ = new_B1605_ | new_B1638_;
  assign new_B1640_ = ~new_B1605_ & ~new_B1639_;
  assign new_B1639_ = new_B1605_ & new_B1638_;
  assign new_B1638_ = ~new_B1594_ | ~new_B1619_;
  assign new_B1637_ = ~new_B1595_ & new_B1605_;
  assign new_B1636_ = new_B1595_ & ~new_B1605_;
  assign new_B1635_ = new_B1597_ & new_B1634_;
  assign new_B1634_ = new_B1653_ | new_B1652_;
  assign new_B1633_ = ~new_B1597_ & new_B1632_;
  assign new_B1632_ = new_B1655_ | new_B1654_;
  assign new_B1631_ = new_B1597_ | new_B1630_;
  assign new_B1630_ = new_B1651_ | new_B1650_;
  assign new_B1629_ = ~new_B1609_ & ~new_B1619_;
  assign new_B1628_ = new_B1609_ & new_B1619_;
  assign new_B1627_ = ~new_B1609_ | new_B1619_;
  assign new_B1626_ = new_B1593_ & ~new_B1594_;
  assign new_B1625_ = ~new_B1593_ & new_B1594_;
  assign new_B1624_ = new_B1646_ & ~new_B1647_;
  assign new_B1623_ = ~new_B1646_ & new_B1647_;
  assign new_B1622_ = ~new_B1645_ | ~new_B1644_;
  assign new_B1621_ = new_B1637_ | new_B1636_;
  assign new_B1620_ = new_B1643_ | new_B1642_;
  assign new_B1619_ = new_B1633_ | new_B1635_;
  assign new_B1618_ = ~new_B1640_ | ~new_B1641_;
  assign new_B1617_ = new_B1593_ & ~new_B1594_;
  assign new_B1616_ = new_B1607_ & ~new_B1619_;
  assign new_B1615_ = ~new_B1607_ & new_B1619_;
  assign new_B1614_ = ~new_B1605_ & new_B1631_;
  assign new_B1613_ = new_B1629_ | new_B1628_;
  assign new_B1612_ = new_B1626_ | new_B1625_;
  assign new_B1611_ = new_B1594_ | new_B1627_;
  assign new_B1610_ = new_B1619_ & new_B1622_;
  assign new_B1609_ = new_B1624_ | new_B1623_;
  assign new_B1608_ = new_B1619_ & new_B1618_;
  assign new_B1607_ = new_B1621_ & new_B1620_;
  assign new_B1606_ = new_B1616_ | new_B1615_;
  assign new_B1605_ = new_B1594_ | new_B1617_;
  assign B1604 = new_B1605_ | new_B1614_;
  assign B1603 = new_B1612_ & new_B1613_;
  assign B1602 = new_B1612_ & new_B1611_;
  assign B1601 = new_B1610_ | new_B1609_;
  assign B1600 = new_B1608_ | new_B1607_;
  assign B1599 = new_B1606_ & new_B1605_;
  assign new_B1598_ = new_C9691_;
  assign new_B1597_ = new_C9624_;
  assign new_B1596_ = new_C9557_;
  assign new_B1595_ = new_C9490_;
  assign new_B1594_ = new_C9423_;
  assign new_B1593_ = new_C9356_;
  assign new_B1592_ = ~new_B1531_ & new_B1545_;
  assign new_B1591_ = new_B1531_ & ~new_B1545_;
  assign new_B1590_ = new_B1531_ & ~new_B1545_;
  assign new_B1589_ = ~new_B1531_ & ~new_B1545_;
  assign new_B1588_ = new_B1531_ & new_B1545_;
  assign new_B1587_ = new_B1591_ | new_B1592_;
  assign new_B1586_ = ~new_B1531_ & new_B1545_;
  assign new_B1585_ = new_B1589_ | new_B1590_;
  assign new_B1584_ = ~new_B1560_ & ~new_B1580_;
  assign new_B1583_ = new_B1560_ & new_B1580_;
  assign new_B1582_ = ~new_B1527_ | ~new_B1552_;
  assign new_B1581_ = new_B1545_ & new_B1582_;
  assign new_B1580_ = new_B1528_ | new_B1529_;
  assign new_B1579_ = new_B1528_ | new_B1545_;
  assign new_B1578_ = ~new_B1545_ & ~new_B1581_;
  assign new_B1577_ = new_B1545_ | new_B1582_;
  assign new_B1576_ = new_B1528_ & ~new_B1529_;
  assign new_B1575_ = ~new_B1528_ & new_B1529_;
  assign new_B1574_ = new_B1538_ | new_B1571_;
  assign new_B1573_ = ~new_B1538_ & ~new_B1572_;
  assign new_B1572_ = new_B1538_ & new_B1571_;
  assign new_B1571_ = ~new_B1527_ | ~new_B1552_;
  assign new_B1570_ = ~new_B1528_ & new_B1538_;
  assign new_B1569_ = new_B1528_ & ~new_B1538_;
  assign new_B1568_ = new_B1530_ & new_B1567_;
  assign new_B1567_ = new_B1586_ | new_B1585_;
  assign new_B1566_ = ~new_B1530_ & new_B1565_;
  assign new_B1565_ = new_B1588_ | new_B1587_;
  assign new_B1564_ = new_B1530_ | new_B1563_;
  assign new_B1563_ = new_B1584_ | new_B1583_;
  assign new_B1562_ = ~new_B1542_ & ~new_B1552_;
  assign new_B1561_ = new_B1542_ & new_B1552_;
  assign new_B1560_ = ~new_B1542_ | new_B1552_;
  assign new_B1559_ = new_B1526_ & ~new_B1527_;
  assign new_B1558_ = ~new_B1526_ & new_B1527_;
  assign new_B1557_ = new_B1579_ & ~new_B1580_;
  assign new_B1556_ = ~new_B1579_ & new_B1580_;
  assign new_B1555_ = ~new_B1578_ | ~new_B1577_;
  assign new_B1554_ = new_B1570_ | new_B1569_;
  assign new_B1553_ = new_B1576_ | new_B1575_;
  assign new_B1552_ = new_B1566_ | new_B1568_;
  assign new_B1551_ = ~new_B1573_ | ~new_B1574_;
  assign new_B1550_ = new_B1526_ & ~new_B1527_;
  assign new_B1549_ = new_B1540_ & ~new_B1552_;
  assign new_B1548_ = ~new_B1540_ & new_B1552_;
  assign new_B1547_ = ~new_B1538_ & new_B1564_;
  assign new_B1546_ = new_B1562_ | new_B1561_;
  assign new_B1545_ = new_B1559_ | new_B1558_;
  assign new_B1544_ = new_B1527_ | new_B1560_;
  assign new_B1543_ = new_B1552_ & new_B1555_;
  assign new_B1542_ = new_B1557_ | new_B1556_;
  assign new_B1541_ = new_B1552_ & new_B1551_;
  assign new_B1540_ = new_B1554_ & new_B1553_;
  assign new_B1539_ = new_B1549_ | new_B1548_;
  assign new_B1538_ = new_B1527_ | new_B1550_;
  assign B1537 = new_B1538_ | new_B1547_;
  assign B1536 = new_B1545_ & new_B1546_;
  assign B1535 = new_B1545_ & new_B1544_;
  assign B1534 = new_B1543_ | new_B1542_;
  assign B1533 = new_B1541_ | new_B1540_;
  assign B1532 = new_B1539_ & new_B1538_;
  assign new_B1531_ = new_C9289_;
  assign new_B1530_ = new_C9222_;
  assign new_B1529_ = new_C9155_;
  assign new_B1528_ = new_C9088_;
  assign new_B1527_ = new_C9021_;
  assign new_B1526_ = new_C8954_;
  assign new_B1525_ = ~new_B1464_ & new_B1478_;
  assign new_B1524_ = new_B1464_ & ~new_B1478_;
  assign new_B1523_ = new_B1464_ & ~new_B1478_;
  assign new_B1522_ = ~new_B1464_ & ~new_B1478_;
  assign new_B1521_ = new_B1464_ & new_B1478_;
  assign new_B1520_ = new_B1524_ | new_B1525_;
  assign new_B1519_ = ~new_B1464_ & new_B1478_;
  assign new_B1518_ = new_B1522_ | new_B1523_;
  assign new_B1517_ = ~new_B1493_ & ~new_B1513_;
  assign new_B1516_ = new_B1493_ & new_B1513_;
  assign new_B1515_ = ~new_B1460_ | ~new_B1485_;
  assign new_B1514_ = new_B1478_ & new_B1515_;
  assign new_B1513_ = new_B1461_ | new_B1462_;
  assign new_B1512_ = new_B1461_ | new_B1478_;
  assign new_B1511_ = ~new_B1478_ & ~new_B1514_;
  assign new_B1510_ = new_B1478_ | new_B1515_;
  assign new_B1509_ = new_B1461_ & ~new_B1462_;
  assign new_B1508_ = ~new_B1461_ & new_B1462_;
  assign new_B1507_ = new_B1471_ | new_B1504_;
  assign new_B1506_ = ~new_B1471_ & ~new_B1505_;
  assign new_B1505_ = new_B1471_ & new_B1504_;
  assign new_B1504_ = ~new_B1460_ | ~new_B1485_;
  assign new_B1503_ = ~new_B1461_ & new_B1471_;
  assign new_B1502_ = new_B1461_ & ~new_B1471_;
  assign new_B1501_ = new_B1463_ & new_B1500_;
  assign new_B1500_ = new_B1519_ | new_B1518_;
  assign new_B1499_ = ~new_B1463_ & new_B1498_;
  assign new_B1498_ = new_B1521_ | new_B1520_;
  assign new_B1497_ = new_B1463_ | new_B1496_;
  assign new_B1496_ = new_B1517_ | new_B1516_;
  assign new_B1495_ = ~new_B1475_ & ~new_B1485_;
  assign new_B1494_ = new_B1475_ & new_B1485_;
  assign new_B1493_ = ~new_B1475_ | new_B1485_;
  assign new_B1492_ = new_B1459_ & ~new_B1460_;
  assign new_B1491_ = ~new_B1459_ & new_B1460_;
  assign new_B1490_ = new_B1512_ & ~new_B1513_;
  assign new_B1489_ = ~new_B1512_ & new_B1513_;
  assign new_B1488_ = ~new_B1511_ | ~new_B1510_;
  assign new_B1487_ = new_B1503_ | new_B1502_;
  assign new_B1486_ = new_B1509_ | new_B1508_;
  assign new_B1485_ = new_B1499_ | new_B1501_;
  assign new_B1484_ = ~new_B1506_ | ~new_B1507_;
  assign new_B1483_ = new_B1459_ & ~new_B1460_;
  assign new_B1482_ = new_B1473_ & ~new_B1485_;
  assign new_B1481_ = ~new_B1473_ & new_B1485_;
  assign new_B1480_ = ~new_B1471_ & new_B1497_;
  assign new_B1479_ = new_B1495_ | new_B1494_;
  assign new_B1478_ = new_B1492_ | new_B1491_;
  assign new_B1477_ = new_B1460_ | new_B1493_;
  assign new_B1476_ = new_B1485_ & new_B1488_;
  assign new_B1475_ = new_B1490_ | new_B1489_;
  assign new_B1474_ = new_B1485_ & new_B1484_;
  assign new_B1473_ = new_B1487_ & new_B1486_;
  assign new_B1472_ = new_B1482_ | new_B1481_;
  assign new_B1471_ = new_B1460_ | new_B1483_;
  assign B1470 = new_B1471_ | new_B1480_;
  assign B1469 = new_B1478_ & new_B1479_;
  assign B1468 = new_B1478_ & new_B1477_;
  assign B1467 = new_B1476_ | new_B1475_;
  assign B1466 = new_B1474_ | new_B1473_;
  assign B1465 = new_B1472_ & new_B1471_;
  assign new_B1464_ = new_C8887_;
  assign new_B1463_ = new_C8820_;
  assign new_B1462_ = new_C8753_;
  assign new_B1461_ = new_C8686_;
  assign new_B1460_ = new_C8619_;
  assign new_B1459_ = new_C8552_;
  assign new_B1458_ = ~new_B1397_ & new_B1411_;
  assign new_B1457_ = new_B1397_ & ~new_B1411_;
  assign new_B1456_ = new_B1397_ & ~new_B1411_;
  assign new_B1455_ = ~new_B1397_ & ~new_B1411_;
  assign new_B1454_ = new_B1397_ & new_B1411_;
  assign new_B1453_ = new_B1457_ | new_B1458_;
  assign new_B1452_ = ~new_B1397_ & new_B1411_;
  assign new_B1451_ = new_B1455_ | new_B1456_;
  assign new_B1450_ = ~new_B1426_ & ~new_B1446_;
  assign new_B1449_ = new_B1426_ & new_B1446_;
  assign new_B1448_ = ~new_B1393_ | ~new_B1418_;
  assign new_B1447_ = new_B1411_ & new_B1448_;
  assign new_B1446_ = new_B1394_ | new_B1395_;
  assign new_B1445_ = new_B1394_ | new_B1411_;
  assign new_B1444_ = ~new_B1411_ & ~new_B1447_;
  assign new_B1443_ = new_B1411_ | new_B1448_;
  assign new_B1442_ = new_B1394_ & ~new_B1395_;
  assign new_B1441_ = ~new_B1394_ & new_B1395_;
  assign new_B1440_ = new_B1404_ | new_B1437_;
  assign new_B1439_ = ~new_B1404_ & ~new_B1438_;
  assign new_B1438_ = new_B1404_ & new_B1437_;
  assign new_B1437_ = ~new_B1393_ | ~new_B1418_;
  assign new_B1436_ = ~new_B1394_ & new_B1404_;
  assign new_B1435_ = new_B1394_ & ~new_B1404_;
  assign new_B1434_ = new_B1396_ & new_B1433_;
  assign new_B1433_ = new_B1452_ | new_B1451_;
  assign new_B1432_ = ~new_B1396_ & new_B1431_;
  assign new_B1431_ = new_B1454_ | new_B1453_;
  assign new_B1430_ = new_B1396_ | new_B1429_;
  assign new_B1429_ = new_B1450_ | new_B1449_;
  assign new_B1428_ = ~new_B1408_ & ~new_B1418_;
  assign new_B1427_ = new_B1408_ & new_B1418_;
  assign new_B1426_ = ~new_B1408_ | new_B1418_;
  assign new_B1425_ = new_B1392_ & ~new_B1393_;
  assign new_B1424_ = ~new_B1392_ & new_B1393_;
  assign new_B1423_ = new_B1445_ & ~new_B1446_;
  assign new_B1422_ = ~new_B1445_ & new_B1446_;
  assign new_B1421_ = ~new_B1444_ | ~new_B1443_;
  assign new_B1420_ = new_B1436_ | new_B1435_;
  assign new_B1419_ = new_B1442_ | new_B1441_;
  assign new_B1418_ = new_B1432_ | new_B1434_;
  assign new_B1417_ = ~new_B1439_ | ~new_B1440_;
  assign new_B1416_ = new_B1392_ & ~new_B1393_;
  assign new_B1415_ = new_B1406_ & ~new_B1418_;
  assign new_B1414_ = ~new_B1406_ & new_B1418_;
  assign new_B1413_ = ~new_B1404_ & new_B1430_;
  assign new_B1412_ = new_B1428_ | new_B1427_;
  assign new_B1411_ = new_B1425_ | new_B1424_;
  assign new_B1410_ = new_B1393_ | new_B1426_;
  assign new_B1409_ = new_B1418_ & new_B1421_;
  assign new_B1408_ = new_B1423_ | new_B1422_;
  assign new_B1407_ = new_B1418_ & new_B1417_;
  assign new_B1406_ = new_B1420_ & new_B1419_;
  assign new_B1405_ = new_B1415_ | new_B1414_;
  assign new_B1404_ = new_B1393_ | new_B1416_;
  assign B1403 = new_B1404_ | new_B1413_;
  assign B1402 = new_B1411_ & new_B1412_;
  assign B1401 = new_B1411_ & new_B1410_;
  assign B1400 = new_B1409_ | new_B1408_;
  assign B1399 = new_B1407_ | new_B1406_;
  assign B1398 = new_B1405_ & new_B1404_;
  assign new_B1397_ = new_C8485_;
  assign new_B1396_ = new_C8418_;
  assign new_B1395_ = new_C8351_;
  assign new_B1394_ = new_C8284_;
  assign new_B1393_ = new_C8217_;
  assign new_B1392_ = new_C8150_;
  assign new_B1391_ = ~new_B1330_ & new_B1344_;
  assign new_B1390_ = new_B1330_ & ~new_B1344_;
  assign new_B1389_ = new_B1330_ & ~new_B1344_;
  assign new_B1388_ = ~new_B1330_ & ~new_B1344_;
  assign new_B1387_ = new_B1330_ & new_B1344_;
  assign new_B1386_ = new_B1390_ | new_B1391_;
  assign new_B1385_ = ~new_B1330_ & new_B1344_;
  assign new_B1384_ = new_B1388_ | new_B1389_;
  assign new_B1383_ = ~new_B1359_ & ~new_B1379_;
  assign new_B1382_ = new_B1359_ & new_B1379_;
  assign new_B1381_ = ~new_B1326_ | ~new_B1351_;
  assign new_B1380_ = new_B1344_ & new_B1381_;
  assign new_B1379_ = new_B1327_ | new_B1328_;
  assign new_B1378_ = new_B1327_ | new_B1344_;
  assign new_B1377_ = ~new_B1344_ & ~new_B1380_;
  assign new_B1376_ = new_B1344_ | new_B1381_;
  assign new_B1375_ = new_B1327_ & ~new_B1328_;
  assign new_B1374_ = ~new_B1327_ & new_B1328_;
  assign new_B1373_ = new_B1337_ | new_B1370_;
  assign new_B1372_ = ~new_B1337_ & ~new_B1371_;
  assign new_B1371_ = new_B1337_ & new_B1370_;
  assign new_B1370_ = ~new_B1326_ | ~new_B1351_;
  assign new_B1369_ = ~new_B1327_ & new_B1337_;
  assign new_B1368_ = new_B1327_ & ~new_B1337_;
  assign new_B1367_ = new_B1329_ & new_B1366_;
  assign new_B1366_ = new_B1385_ | new_B1384_;
  assign new_B1365_ = ~new_B1329_ & new_B1364_;
  assign new_B1364_ = new_B1387_ | new_B1386_;
  assign new_B1363_ = new_B1329_ | new_B1362_;
  assign new_B1362_ = new_B1383_ | new_B1382_;
  assign new_B1361_ = ~new_B1341_ & ~new_B1351_;
  assign new_B1360_ = new_B1341_ & new_B1351_;
  assign new_B1359_ = ~new_B1341_ | new_B1351_;
  assign new_B1358_ = new_B1325_ & ~new_B1326_;
  assign new_B1357_ = ~new_B1325_ & new_B1326_;
  assign new_B1356_ = new_B1378_ & ~new_B1379_;
  assign new_B1355_ = ~new_B1378_ & new_B1379_;
  assign new_B1354_ = ~new_B1377_ | ~new_B1376_;
  assign new_B1353_ = new_B1369_ | new_B1368_;
  assign new_B1352_ = new_B1375_ | new_B1374_;
  assign new_B1351_ = new_B1365_ | new_B1367_;
  assign new_B1350_ = ~new_B1372_ | ~new_B1373_;
  assign new_B1349_ = new_B1325_ & ~new_B1326_;
  assign new_B1348_ = new_B1339_ & ~new_B1351_;
  assign new_B1347_ = ~new_B1339_ & new_B1351_;
  assign new_B1346_ = ~new_B1337_ & new_B1363_;
  assign new_B1345_ = new_B1361_ | new_B1360_;
  assign new_B1344_ = new_B1358_ | new_B1357_;
  assign new_B1343_ = new_B1326_ | new_B1359_;
  assign new_B1342_ = new_B1351_ & new_B1354_;
  assign new_B1341_ = new_B1356_ | new_B1355_;
  assign new_B1340_ = new_B1351_ & new_B1350_;
  assign new_B1339_ = new_B1353_ & new_B1352_;
  assign new_B1338_ = new_B1348_ | new_B1347_;
  assign new_B1337_ = new_B1326_ | new_B1349_;
  assign B1336 = new_B1337_ | new_B1346_;
  assign B1335 = new_B1344_ & new_B1345_;
  assign B1334 = new_B1344_ & new_B1343_;
  assign B1333 = new_B1342_ | new_B1341_;
  assign B1332 = new_B1340_ | new_B1339_;
  assign B1331 = new_B1338_ & new_B1337_;
  assign new_B1330_ = new_C8083_;
  assign new_B1329_ = new_C8016_;
  assign new_B1328_ = new_C7949_;
  assign new_B1327_ = new_C7882_;
  assign new_B1326_ = new_C7815_;
  assign new_B1325_ = new_C7748_;
  assign new_B1324_ = ~new_B1263_ & new_B1277_;
  assign new_B1323_ = new_B1263_ & ~new_B1277_;
  assign new_B1322_ = new_B1263_ & ~new_B1277_;
  assign new_B1321_ = ~new_B1263_ & ~new_B1277_;
  assign new_B1320_ = new_B1263_ & new_B1277_;
  assign new_B1319_ = new_B1323_ | new_B1324_;
  assign new_B1318_ = ~new_B1263_ & new_B1277_;
  assign new_B1317_ = new_B1321_ | new_B1322_;
  assign new_B1316_ = ~new_B1292_ & ~new_B1312_;
  assign new_B1315_ = new_B1292_ & new_B1312_;
  assign new_B1314_ = ~new_B1259_ | ~new_B1284_;
  assign new_B1313_ = new_B1277_ & new_B1314_;
  assign new_B1312_ = new_B1260_ | new_B1261_;
  assign new_B1311_ = new_B1260_ | new_B1277_;
  assign new_B1310_ = ~new_B1277_ & ~new_B1313_;
  assign new_B1309_ = new_B1277_ | new_B1314_;
  assign new_B1308_ = new_B1260_ & ~new_B1261_;
  assign new_B1307_ = ~new_B1260_ & new_B1261_;
  assign new_B1306_ = new_B1270_ | new_B1303_;
  assign new_B1305_ = ~new_B1270_ & ~new_B1304_;
  assign new_B1304_ = new_B1270_ & new_B1303_;
  assign new_B1303_ = ~new_B1259_ | ~new_B1284_;
  assign new_B1302_ = ~new_B1260_ & new_B1270_;
  assign new_B1301_ = new_B1260_ & ~new_B1270_;
  assign new_B1300_ = new_B1262_ & new_B1299_;
  assign new_B1299_ = new_B1318_ | new_B1317_;
  assign new_B1298_ = ~new_B1262_ & new_B1297_;
  assign new_B1297_ = new_B1320_ | new_B1319_;
  assign new_B1296_ = new_B1262_ | new_B1295_;
  assign new_B1295_ = new_B1316_ | new_B1315_;
  assign new_B1294_ = ~new_B1274_ & ~new_B1284_;
  assign new_B1293_ = new_B1274_ & new_B1284_;
  assign new_B1292_ = ~new_B1274_ | new_B1284_;
  assign new_B1291_ = new_B1258_ & ~new_B1259_;
  assign new_B1290_ = ~new_B1258_ & new_B1259_;
  assign new_B1289_ = new_B1311_ & ~new_B1312_;
  assign new_B1288_ = ~new_B1311_ & new_B1312_;
  assign new_B1287_ = ~new_B1310_ | ~new_B1309_;
  assign new_B1286_ = new_B1302_ | new_B1301_;
  assign new_B1285_ = new_B1308_ | new_B1307_;
  assign new_B1284_ = new_B1298_ | new_B1300_;
  assign new_B1283_ = ~new_B1305_ | ~new_B1306_;
  assign new_B1282_ = new_B1258_ & ~new_B1259_;
  assign new_B1281_ = new_B1272_ & ~new_B1284_;
  assign new_B1280_ = ~new_B1272_ & new_B1284_;
  assign new_B1279_ = ~new_B1270_ & new_B1296_;
  assign new_B1278_ = new_B1294_ | new_B1293_;
  assign new_B1277_ = new_B1291_ | new_B1290_;
  assign new_B1276_ = new_B1259_ | new_B1292_;
  assign new_B1275_ = new_B1284_ & new_B1287_;
  assign new_B1274_ = new_B1289_ | new_B1288_;
  assign new_B1273_ = new_B1284_ & new_B1283_;
  assign new_B1272_ = new_B1286_ & new_B1285_;
  assign new_B1271_ = new_B1281_ | new_B1280_;
  assign new_B1270_ = new_B1259_ | new_B1282_;
  assign B1269 = new_B1270_ | new_B1279_;
  assign B1268 = new_B1277_ & new_B1278_;
  assign B1267 = new_B1277_ & new_B1276_;
  assign B1266 = new_B1275_ | new_B1274_;
  assign B1265 = new_B1273_ | new_B1272_;
  assign B1264 = new_B1271_ & new_B1270_;
  assign new_B1263_ = new_C7681_;
  assign new_B1262_ = new_C7614_;
  assign new_B1261_ = new_C7547_;
  assign new_B1260_ = new_C7480_;
  assign new_B1259_ = new_C7413_;
  assign new_B1258_ = new_C7346_;
  assign new_B1257_ = ~new_B1196_ & new_B1210_;
  assign new_B1256_ = new_B1196_ & ~new_B1210_;
  assign new_B1255_ = new_B1196_ & ~new_B1210_;
  assign new_B1254_ = ~new_B1196_ & ~new_B1210_;
  assign new_B1253_ = new_B1196_ & new_B1210_;
  assign new_B1252_ = new_B1256_ | new_B1257_;
  assign new_B1251_ = ~new_B1196_ & new_B1210_;
  assign new_B1250_ = new_B1254_ | new_B1255_;
  assign new_B1249_ = ~new_B1225_ & ~new_B1245_;
  assign new_B1248_ = new_B1225_ & new_B1245_;
  assign new_B1247_ = ~new_B1192_ | ~new_B1217_;
  assign new_B1246_ = new_B1210_ & new_B1247_;
  assign new_B1245_ = new_B1193_ | new_B1194_;
  assign new_B1244_ = new_B1193_ | new_B1210_;
  assign new_B1243_ = ~new_B1210_ & ~new_B1246_;
  assign new_B1242_ = new_B1210_ | new_B1247_;
  assign new_B1241_ = new_B1193_ & ~new_B1194_;
  assign new_B1240_ = ~new_B1193_ & new_B1194_;
  assign new_B1239_ = new_B1203_ | new_B1236_;
  assign new_B1238_ = ~new_B1203_ & ~new_B1237_;
  assign new_B1237_ = new_B1203_ & new_B1236_;
  assign new_B1236_ = ~new_B1192_ | ~new_B1217_;
  assign new_B1235_ = ~new_B1193_ & new_B1203_;
  assign new_B1234_ = new_B1193_ & ~new_B1203_;
  assign new_B1233_ = new_B1195_ & new_B1232_;
  assign new_B1232_ = new_B1251_ | new_B1250_;
  assign new_B1231_ = ~new_B1195_ & new_B1230_;
  assign new_B1230_ = new_B1253_ | new_B1252_;
  assign new_B1229_ = new_B1195_ | new_B1228_;
  assign new_B1228_ = new_B1249_ | new_B1248_;
  assign new_B1227_ = ~new_B1207_ & ~new_B1217_;
  assign new_B1226_ = new_B1207_ & new_B1217_;
  assign new_B1225_ = ~new_B1207_ | new_B1217_;
  assign new_B1224_ = new_B1191_ & ~new_B1192_;
  assign new_B1223_ = ~new_B1191_ & new_B1192_;
  assign new_B1222_ = new_B1244_ & ~new_B1245_;
  assign new_B1221_ = ~new_B1244_ & new_B1245_;
  assign new_B1220_ = ~new_B1243_ | ~new_B1242_;
  assign new_B1219_ = new_B1235_ | new_B1234_;
  assign new_B1218_ = new_B1241_ | new_B1240_;
  assign new_B1217_ = new_B1231_ | new_B1233_;
  assign new_B1216_ = ~new_B1238_ | ~new_B1239_;
  assign new_B1215_ = new_B1191_ & ~new_B1192_;
  assign new_B1214_ = new_B1205_ & ~new_B1217_;
  assign new_B1213_ = ~new_B1205_ & new_B1217_;
  assign new_B1212_ = ~new_B1203_ & new_B1229_;
  assign new_B1211_ = new_B1227_ | new_B1226_;
  assign new_B1210_ = new_B1224_ | new_B1223_;
  assign new_B1209_ = new_B1192_ | new_B1225_;
  assign new_B1208_ = new_B1217_ & new_B1220_;
  assign new_B1207_ = new_B1222_ | new_B1221_;
  assign new_B1206_ = new_B1217_ & new_B1216_;
  assign new_B1205_ = new_B1219_ & new_B1218_;
  assign new_B1204_ = new_B1214_ | new_B1213_;
  assign new_B1203_ = new_B1192_ | new_B1215_;
  assign B1202 = new_B1203_ | new_B1212_;
  assign B1201 = new_B1210_ & new_B1211_;
  assign B1200 = new_B1210_ & new_B1209_;
  assign B1199 = new_B1208_ | new_B1207_;
  assign B1198 = new_B1206_ | new_B1205_;
  assign B1197 = new_B1204_ & new_B1203_;
  assign new_B1196_ = new_C7279_;
  assign new_B1195_ = new_C7212_;
  assign new_B1194_ = new_C7145_;
  assign new_B1193_ = new_C7078_;
  assign new_B1192_ = new_C7011_;
  assign new_B1191_ = new_C6944_;
  assign new_B1190_ = ~new_B1129_ & new_B1143_;
  assign new_B1189_ = new_B1129_ & ~new_B1143_;
  assign new_B1188_ = new_B1129_ & ~new_B1143_;
  assign new_B1187_ = ~new_B1129_ & ~new_B1143_;
  assign new_B1186_ = new_B1129_ & new_B1143_;
  assign new_B1185_ = new_B1189_ | new_B1190_;
  assign new_B1184_ = ~new_B1129_ & new_B1143_;
  assign new_B1183_ = new_B1187_ | new_B1188_;
  assign new_B1182_ = ~new_B1158_ & ~new_B1178_;
  assign new_B1181_ = new_B1158_ & new_B1178_;
  assign new_B1180_ = ~new_B1125_ | ~new_B1150_;
  assign new_B1179_ = new_B1143_ & new_B1180_;
  assign new_B1178_ = new_B1126_ | new_B1127_;
  assign new_B1177_ = new_B1126_ | new_B1143_;
  assign new_B1176_ = ~new_B1143_ & ~new_B1179_;
  assign new_B1175_ = new_B1143_ | new_B1180_;
  assign new_B1174_ = new_B1126_ & ~new_B1127_;
  assign new_B1173_ = ~new_B1126_ & new_B1127_;
  assign new_B1172_ = new_B1136_ | new_B1169_;
  assign new_B1171_ = ~new_B1136_ & ~new_B1170_;
  assign new_B1170_ = new_B1136_ & new_B1169_;
  assign new_B1169_ = ~new_B1125_ | ~new_B1150_;
  assign new_B1168_ = ~new_B1126_ & new_B1136_;
  assign new_B1167_ = new_B1126_ & ~new_B1136_;
  assign new_B1166_ = new_B1128_ & new_B1165_;
  assign new_B1165_ = new_B1184_ | new_B1183_;
  assign new_B1164_ = ~new_B1128_ & new_B1163_;
  assign new_B1163_ = new_B1186_ | new_B1185_;
  assign new_B1162_ = new_B1128_ | new_B1161_;
  assign new_B1161_ = new_B1182_ | new_B1181_;
  assign new_B1160_ = ~new_B1140_ & ~new_B1150_;
  assign new_B1159_ = new_B1140_ & new_B1150_;
  assign new_B1158_ = ~new_B1140_ | new_B1150_;
  assign new_B1157_ = new_B1124_ & ~new_B1125_;
  assign new_B1156_ = ~new_B1124_ & new_B1125_;
  assign new_B1155_ = new_B1177_ & ~new_B1178_;
  assign new_B1154_ = ~new_B1177_ & new_B1178_;
  assign new_B1153_ = ~new_B1176_ | ~new_B1175_;
  assign new_B1152_ = new_B1168_ | new_B1167_;
  assign new_B1151_ = new_B1174_ | new_B1173_;
  assign new_B1150_ = new_B1164_ | new_B1166_;
  assign new_B1149_ = ~new_B1171_ | ~new_B1172_;
  assign new_B1148_ = new_B1124_ & ~new_B1125_;
  assign new_B1147_ = new_B1138_ & ~new_B1150_;
  assign new_B1146_ = ~new_B1138_ & new_B1150_;
  assign new_B1145_ = ~new_B1136_ & new_B1162_;
  assign new_B1144_ = new_B1160_ | new_B1159_;
  assign new_B1143_ = new_B1157_ | new_B1156_;
  assign new_B1142_ = new_B1125_ | new_B1158_;
  assign new_B1141_ = new_B1150_ & new_B1153_;
  assign new_B1140_ = new_B1155_ | new_B1154_;
  assign new_B1139_ = new_B1150_ & new_B1149_;
  assign new_B1138_ = new_B1152_ & new_B1151_;
  assign new_B1137_ = new_B1147_ | new_B1146_;
  assign new_B1136_ = new_B1125_ | new_B1148_;
  assign B1135 = new_B1136_ | new_B1145_;
  assign B1134 = new_B1143_ & new_B1144_;
  assign B1133 = new_B1143_ & new_B1142_;
  assign B1132 = new_B1141_ | new_B1140_;
  assign B1131 = new_B1139_ | new_B1138_;
  assign B1130 = new_B1137_ & new_B1136_;
  assign new_B1129_ = new_C6877_;
  assign new_B1128_ = new_C6810_;
  assign new_B1127_ = new_C6743_;
  assign new_B1126_ = new_C6676_;
  assign new_B1125_ = new_C6609_;
  assign new_B1124_ = new_C6542_;
  assign new_B1123_ = ~new_B1062_ & new_B1076_;
  assign new_B1122_ = new_B1062_ & ~new_B1076_;
  assign new_B1121_ = new_B1062_ & ~new_B1076_;
  assign new_B1120_ = ~new_B1062_ & ~new_B1076_;
  assign new_B1119_ = new_B1062_ & new_B1076_;
  assign new_B1118_ = new_B1122_ | new_B1123_;
  assign new_B1117_ = ~new_B1062_ & new_B1076_;
  assign new_B1116_ = new_B1120_ | new_B1121_;
  assign new_B1115_ = ~new_B1091_ & ~new_B1111_;
  assign new_B1114_ = new_B1091_ & new_B1111_;
  assign new_B1113_ = ~new_B1058_ | ~new_B1083_;
  assign new_B1112_ = new_B1076_ & new_B1113_;
  assign new_B1111_ = new_B1059_ | new_B1060_;
  assign new_B1110_ = new_B1059_ | new_B1076_;
  assign new_B1109_ = ~new_B1076_ & ~new_B1112_;
  assign new_B1108_ = new_B1076_ | new_B1113_;
  assign new_B1107_ = new_B1059_ & ~new_B1060_;
  assign new_B1106_ = ~new_B1059_ & new_B1060_;
  assign new_B1105_ = new_B1069_ | new_B1102_;
  assign new_B1104_ = ~new_B1069_ & ~new_B1103_;
  assign new_B1103_ = new_B1069_ & new_B1102_;
  assign new_B1102_ = ~new_B1058_ | ~new_B1083_;
  assign new_B1101_ = ~new_B1059_ & new_B1069_;
  assign new_B1100_ = new_B1059_ & ~new_B1069_;
  assign new_B1099_ = new_B1061_ & new_B1098_;
  assign new_B1098_ = new_B1117_ | new_B1116_;
  assign new_B1097_ = ~new_B1061_ & new_B1096_;
  assign new_B1096_ = new_B1119_ | new_B1118_;
  assign new_B1095_ = new_B1061_ | new_B1094_;
  assign new_B1094_ = new_B1115_ | new_B1114_;
  assign new_B1093_ = ~new_B1073_ & ~new_B1083_;
  assign new_B1092_ = new_B1073_ & new_B1083_;
  assign new_B1091_ = ~new_B1073_ | new_B1083_;
  assign new_B1090_ = new_B1057_ & ~new_B1058_;
  assign new_B1089_ = ~new_B1057_ & new_B1058_;
  assign new_B1088_ = new_B1110_ & ~new_B1111_;
  assign new_B1087_ = ~new_B1110_ & new_B1111_;
  assign new_B1086_ = ~new_B1109_ | ~new_B1108_;
  assign new_B1085_ = new_B1101_ | new_B1100_;
  assign new_B1084_ = new_B1107_ | new_B1106_;
  assign new_B1083_ = new_B1097_ | new_B1099_;
  assign new_B1082_ = ~new_B1104_ | ~new_B1105_;
  assign new_B1081_ = new_B1057_ & ~new_B1058_;
  assign new_B1080_ = new_B1071_ & ~new_B1083_;
  assign new_B1079_ = ~new_B1071_ & new_B1083_;
  assign new_B1078_ = ~new_B1069_ & new_B1095_;
  assign new_B1077_ = new_B1093_ | new_B1092_;
  assign new_B1076_ = new_B1090_ | new_B1089_;
  assign new_B1075_ = new_B1058_ | new_B1091_;
  assign new_B1074_ = new_B1083_ & new_B1086_;
  assign new_B1073_ = new_B1088_ | new_B1087_;
  assign new_B1072_ = new_B1083_ & new_B1082_;
  assign new_B1071_ = new_B1085_ & new_B1084_;
  assign new_B1070_ = new_B1080_ | new_B1079_;
  assign new_B1069_ = new_B1058_ | new_B1081_;
  assign B1068 = new_B1069_ | new_B1078_;
  assign B1067 = new_B1076_ & new_B1077_;
  assign B1066 = new_B1076_ & new_B1075_;
  assign B1065 = new_B1074_ | new_B1073_;
  assign B1064 = new_B1072_ | new_B1071_;
  assign B1063 = new_B1070_ & new_B1069_;
  assign new_B1062_ = new_C6475_;
  assign new_B1061_ = new_C6408_;
  assign new_B1060_ = new_C6341_;
  assign new_B1059_ = new_C6274_;
  assign new_B1058_ = new_C6207_;
  assign new_B1057_ = new_C6140_;
  assign new_B1056_ = ~new_B995_ & new_B1009_;
  assign new_B1055_ = new_B995_ & ~new_B1009_;
  assign new_B1054_ = new_B995_ & ~new_B1009_;
  assign new_B1053_ = ~new_B995_ & ~new_B1009_;
  assign new_B1052_ = new_B995_ & new_B1009_;
  assign new_B1051_ = new_B1055_ | new_B1056_;
  assign new_B1050_ = ~new_B995_ & new_B1009_;
  assign new_B1049_ = new_B1053_ | new_B1054_;
  assign new_B1048_ = ~new_B1024_ & ~new_B1044_;
  assign new_B1047_ = new_B1024_ & new_B1044_;
  assign new_B1046_ = ~new_B991_ | ~new_B1016_;
  assign new_B1045_ = new_B1009_ & new_B1046_;
  assign new_B1044_ = new_B992_ | new_B993_;
  assign new_B1043_ = new_B992_ | new_B1009_;
  assign new_B1042_ = ~new_B1009_ & ~new_B1045_;
  assign new_B1041_ = new_B1009_ | new_B1046_;
  assign new_B1040_ = new_B992_ & ~new_B993_;
  assign new_B1039_ = ~new_B992_ & new_B993_;
  assign new_B1038_ = new_B1002_ | new_B1035_;
  assign new_B1037_ = ~new_B1002_ & ~new_B1036_;
  assign new_B1036_ = new_B1002_ & new_B1035_;
  assign new_B1035_ = ~new_B991_ | ~new_B1016_;
  assign new_B1034_ = ~new_B992_ & new_B1002_;
  assign new_B1033_ = new_B992_ & ~new_B1002_;
  assign new_B1032_ = new_B994_ & new_B1031_;
  assign new_B1031_ = new_B1050_ | new_B1049_;
  assign new_B1030_ = ~new_B994_ & new_B1029_;
  assign new_B1029_ = new_B1052_ | new_B1051_;
  assign new_B1028_ = new_B994_ | new_B1027_;
  assign new_B1027_ = new_B1048_ | new_B1047_;
  assign new_B1026_ = ~new_B1006_ & ~new_B1016_;
  assign new_B1025_ = new_B1006_ & new_B1016_;
  assign new_B1024_ = ~new_B1006_ | new_B1016_;
  assign new_B1023_ = new_B990_ & ~new_B991_;
  assign new_B1022_ = ~new_B990_ & new_B991_;
  assign new_B1021_ = new_B1043_ & ~new_B1044_;
  assign new_B1020_ = ~new_B1043_ & new_B1044_;
  assign new_B1019_ = ~new_B1042_ | ~new_B1041_;
  assign new_B1018_ = new_B1034_ | new_B1033_;
  assign new_B1017_ = new_B1040_ | new_B1039_;
  assign new_B1016_ = new_B1030_ | new_B1032_;
  assign new_B1015_ = ~new_B1037_ | ~new_B1038_;
  assign new_B1014_ = new_B990_ & ~new_B991_;
  assign new_B1013_ = new_B1004_ & ~new_B1016_;
  assign new_B1012_ = ~new_B1004_ & new_B1016_;
  assign new_B1011_ = ~new_B1002_ & new_B1028_;
  assign new_B1010_ = new_B1026_ | new_B1025_;
  assign new_B1009_ = new_B1023_ | new_B1022_;
  assign new_B1008_ = new_B991_ | new_B1024_;
  assign new_B1007_ = new_B1016_ & new_B1019_;
  assign new_B1006_ = new_B1021_ | new_B1020_;
  assign new_B1005_ = new_B1016_ & new_B1015_;
  assign new_B1004_ = new_B1018_ & new_B1017_;
  assign new_B1003_ = new_B1013_ | new_B1012_;
  assign new_B1002_ = new_B991_ | new_B1014_;
  assign B1001 = new_B1002_ | new_B1011_;
  assign B1000 = new_B1009_ & new_B1010_;
  assign B999 = new_B1009_ & new_B1008_;
  assign B998 = new_B1007_ | new_B1006_;
  assign B997 = new_B1005_ | new_B1004_;
  assign B996 = new_B1003_ & new_B1002_;
  assign new_B995_ = new_C6073_;
  assign new_B994_ = new_C6006_;
  assign new_B993_ = new_C5939_;
  assign new_B992_ = new_C5872_;
  assign new_B991_ = new_C5805_;
  assign new_B990_ = new_C5738_;
  assign new_B989_ = ~new_B928_ & new_B942_;
  assign new_B988_ = new_B928_ & ~new_B942_;
  assign new_B987_ = new_B928_ & ~new_B942_;
  assign new_B986_ = ~new_B928_ & ~new_B942_;
  assign new_B985_ = new_B928_ & new_B942_;
  assign new_B984_ = new_B988_ | new_B989_;
  assign new_B983_ = ~new_B928_ & new_B942_;
  assign new_B982_ = new_B986_ | new_B987_;
  assign new_B981_ = ~new_B957_ & ~new_B977_;
  assign new_B980_ = new_B957_ & new_B977_;
  assign new_B979_ = ~new_B924_ | ~new_B949_;
  assign new_B978_ = new_B942_ & new_B979_;
  assign new_B977_ = new_B925_ | new_B926_;
  assign new_B976_ = new_B925_ | new_B942_;
  assign new_B975_ = ~new_B942_ & ~new_B978_;
  assign new_B974_ = new_B942_ | new_B979_;
  assign new_B973_ = new_B925_ & ~new_B926_;
  assign new_B972_ = ~new_B925_ & new_B926_;
  assign new_B971_ = new_B935_ | new_B968_;
  assign new_B970_ = ~new_B935_ & ~new_B969_;
  assign new_B969_ = new_B935_ & new_B968_;
  assign new_B968_ = ~new_B924_ | ~new_B949_;
  assign new_B967_ = ~new_B925_ & new_B935_;
  assign new_B966_ = new_B925_ & ~new_B935_;
  assign new_B965_ = new_B927_ & new_B964_;
  assign new_B964_ = new_B983_ | new_B982_;
  assign new_B963_ = ~new_B927_ & new_B962_;
  assign new_B962_ = new_B985_ | new_B984_;
  assign new_B961_ = new_B927_ | new_B960_;
  assign new_B960_ = new_B981_ | new_B980_;
  assign new_B959_ = ~new_B939_ & ~new_B949_;
  assign new_B958_ = new_B939_ & new_B949_;
  assign new_B957_ = ~new_B939_ | new_B949_;
  assign new_B956_ = new_B923_ & ~new_B924_;
  assign new_B955_ = ~new_B923_ & new_B924_;
  assign new_B954_ = new_B976_ & ~new_B977_;
  assign new_B953_ = ~new_B976_ & new_B977_;
  assign new_B952_ = ~new_B975_ | ~new_B974_;
  assign new_B951_ = new_B967_ | new_B966_;
  assign new_B950_ = new_B973_ | new_B972_;
  assign new_B949_ = new_B963_ | new_B965_;
  assign new_B948_ = ~new_B970_ | ~new_B971_;
  assign new_B947_ = new_B923_ & ~new_B924_;
  assign new_B946_ = new_B937_ & ~new_B949_;
  assign new_B945_ = ~new_B937_ & new_B949_;
  assign new_B944_ = ~new_B935_ & new_B961_;
  assign new_B943_ = new_B959_ | new_B958_;
  assign new_B942_ = new_B956_ | new_B955_;
  assign new_B941_ = new_B924_ | new_B957_;
  assign new_B940_ = new_B949_ & new_B952_;
  assign new_B939_ = new_B954_ | new_B953_;
  assign new_B938_ = new_B949_ & new_B948_;
  assign new_B937_ = new_B951_ & new_B950_;
  assign new_B936_ = new_B946_ | new_B945_;
  assign new_B935_ = new_B924_ | new_B947_;
  assign B934 = new_B935_ | new_B944_;
  assign B933 = new_B942_ & new_B943_;
  assign B932 = new_B942_ & new_B941_;
  assign B931 = new_B940_ | new_B939_;
  assign B930 = new_B938_ | new_B937_;
  assign B929 = new_B936_ & new_B935_;
  assign new_B928_ = new_C5671_;
  assign new_B927_ = new_C5604_;
  assign new_B926_ = new_C5537_;
  assign new_B925_ = new_C5470_;
  assign new_B924_ = new_C5403_;
  assign new_B923_ = new_C5336_;
  assign new_B922_ = ~new_B861_ & new_B875_;
  assign new_B921_ = new_B861_ & ~new_B875_;
  assign new_B920_ = new_B861_ & ~new_B875_;
  assign new_B919_ = ~new_B861_ & ~new_B875_;
  assign new_B918_ = new_B861_ & new_B875_;
  assign new_B917_ = new_B921_ | new_B922_;
  assign new_B916_ = ~new_B861_ & new_B875_;
  assign new_B915_ = new_B919_ | new_B920_;
  assign new_B914_ = ~new_B890_ & ~new_B910_;
  assign new_B913_ = new_B890_ & new_B910_;
  assign new_B912_ = ~new_B857_ | ~new_B882_;
  assign new_B911_ = new_B875_ & new_B912_;
  assign new_B910_ = new_B858_ | new_B859_;
  assign new_B909_ = new_B858_ | new_B875_;
  assign new_B908_ = ~new_B875_ & ~new_B911_;
  assign new_B907_ = new_B875_ | new_B912_;
  assign new_B906_ = new_B858_ & ~new_B859_;
  assign new_B905_ = ~new_B858_ & new_B859_;
  assign new_B904_ = new_B868_ | new_B901_;
  assign new_B903_ = ~new_B868_ & ~new_B902_;
  assign new_B902_ = new_B868_ & new_B901_;
  assign new_B901_ = ~new_B857_ | ~new_B882_;
  assign new_B900_ = ~new_B858_ & new_B868_;
  assign new_B899_ = new_B858_ & ~new_B868_;
  assign new_B898_ = new_B860_ & new_B897_;
  assign new_B897_ = new_B916_ | new_B915_;
  assign new_B896_ = ~new_B860_ & new_B895_;
  assign new_B895_ = new_B918_ | new_B917_;
  assign new_B894_ = new_B860_ | new_B893_;
  assign new_B893_ = new_B914_ | new_B913_;
  assign new_B892_ = ~new_B872_ & ~new_B882_;
  assign new_B891_ = new_B872_ & new_B882_;
  assign new_B890_ = ~new_B872_ | new_B882_;
  assign new_B889_ = new_B856_ & ~new_B857_;
  assign new_B888_ = ~new_B856_ & new_B857_;
  assign new_B887_ = new_B909_ & ~new_B910_;
  assign new_B886_ = ~new_B909_ & new_B910_;
  assign new_B885_ = ~new_B908_ | ~new_B907_;
  assign new_B884_ = new_B900_ | new_B899_;
  assign new_B883_ = new_B906_ | new_B905_;
  assign new_B882_ = new_B896_ | new_B898_;
  assign new_B881_ = ~new_B903_ | ~new_B904_;
  assign new_B880_ = new_B856_ & ~new_B857_;
  assign new_B879_ = new_B870_ & ~new_B882_;
  assign new_B878_ = ~new_B870_ & new_B882_;
  assign new_B877_ = ~new_B868_ & new_B894_;
  assign new_B876_ = new_B892_ | new_B891_;
  assign new_B875_ = new_B889_ | new_B888_;
  assign new_B874_ = new_B857_ | new_B890_;
  assign new_B873_ = new_B882_ & new_B885_;
  assign new_B872_ = new_B887_ | new_B886_;
  assign new_B871_ = new_B882_ & new_B881_;
  assign new_B870_ = new_B884_ & new_B883_;
  assign new_B869_ = new_B879_ | new_B878_;
  assign new_B868_ = new_B857_ | new_B880_;
  assign B867 = new_B868_ | new_B877_;
  assign B866 = new_B875_ & new_B876_;
  assign B865 = new_B875_ & new_B874_;
  assign B864 = new_B873_ | new_B872_;
  assign B863 = new_B871_ | new_B870_;
  assign B862 = new_B869_ & new_B868_;
  assign new_B861_ = new_C5269_;
  assign new_B860_ = new_C5202_;
  assign new_B859_ = new_C5135_;
  assign new_B858_ = new_C5068_;
  assign new_B857_ = new_C5001_;
  assign new_B856_ = new_C4934_;
  assign new_B855_ = ~new_B794_ & new_B808_;
  assign new_B854_ = new_B794_ & ~new_B808_;
  assign new_B853_ = new_B794_ & ~new_B808_;
  assign new_B852_ = ~new_B794_ & ~new_B808_;
  assign new_B851_ = new_B794_ & new_B808_;
  assign new_B850_ = new_B854_ | new_B855_;
  assign new_B849_ = ~new_B794_ & new_B808_;
  assign new_B848_ = new_B852_ | new_B853_;
  assign new_B847_ = ~new_B823_ & ~new_B843_;
  assign new_B846_ = new_B823_ & new_B843_;
  assign new_B845_ = ~new_B790_ | ~new_B815_;
  assign new_B844_ = new_B808_ & new_B845_;
  assign new_B843_ = new_B791_ | new_B792_;
  assign new_B842_ = new_B791_ | new_B808_;
  assign new_B841_ = ~new_B808_ & ~new_B844_;
  assign new_B840_ = new_B808_ | new_B845_;
  assign new_B839_ = new_B791_ & ~new_B792_;
  assign new_B838_ = ~new_B791_ & new_B792_;
  assign new_B837_ = new_B801_ | new_B834_;
  assign new_B836_ = ~new_B801_ & ~new_B835_;
  assign new_B835_ = new_B801_ & new_B834_;
  assign new_B834_ = ~new_B790_ | ~new_B815_;
  assign new_B833_ = ~new_B791_ & new_B801_;
  assign new_B832_ = new_B791_ & ~new_B801_;
  assign new_B831_ = new_B793_ & new_B830_;
  assign new_B830_ = new_B849_ | new_B848_;
  assign new_B829_ = ~new_B793_ & new_B828_;
  assign new_B828_ = new_B851_ | new_B850_;
  assign new_B827_ = new_B793_ | new_B826_;
  assign new_B826_ = new_B847_ | new_B846_;
  assign new_B825_ = ~new_B805_ & ~new_B815_;
  assign new_B824_ = new_B805_ & new_B815_;
  assign new_B823_ = ~new_B805_ | new_B815_;
  assign new_B822_ = new_B789_ & ~new_B790_;
  assign new_B821_ = ~new_B789_ & new_B790_;
  assign new_B820_ = new_B842_ & ~new_B843_;
  assign new_B819_ = ~new_B842_ & new_B843_;
  assign new_B818_ = ~new_B841_ | ~new_B840_;
  assign new_B817_ = new_B833_ | new_B832_;
  assign new_B816_ = new_B839_ | new_B838_;
  assign new_B815_ = new_B829_ | new_B831_;
  assign new_B814_ = ~new_B836_ | ~new_B837_;
  assign new_B813_ = new_B789_ & ~new_B790_;
  assign new_B812_ = new_B803_ & ~new_B815_;
  assign new_B811_ = ~new_B803_ & new_B815_;
  assign new_B810_ = ~new_B801_ & new_B827_;
  assign new_B809_ = new_B825_ | new_B824_;
  assign new_B808_ = new_B822_ | new_B821_;
  assign new_B807_ = new_B790_ | new_B823_;
  assign new_B806_ = new_B815_ & new_B818_;
  assign new_B805_ = new_B820_ | new_B819_;
  assign new_B804_ = new_B815_ & new_B814_;
  assign new_B803_ = new_B817_ & new_B816_;
  assign new_B802_ = new_B812_ | new_B811_;
  assign new_B801_ = new_B790_ | new_B813_;
  assign B800 = new_B801_ | new_B810_;
  assign B799 = new_B808_ & new_B809_;
  assign B798 = new_B808_ & new_B807_;
  assign B797 = new_B806_ | new_B805_;
  assign B796 = new_B804_ | new_B803_;
  assign B795 = new_B802_ & new_B801_;
  assign new_B794_ = new_C4867_;
  assign new_B793_ = new_C4800_;
  assign new_B792_ = new_C4733_;
  assign new_B791_ = new_C4666_;
  assign new_B790_ = new_C4599_;
  assign new_B789_ = new_C4532_;
  assign new_B788_ = ~new_B727_ & new_B741_;
  assign new_B787_ = new_B727_ & ~new_B741_;
  assign new_B786_ = new_B727_ & ~new_B741_;
  assign new_B785_ = ~new_B727_ & ~new_B741_;
  assign new_B784_ = new_B727_ & new_B741_;
  assign new_B783_ = new_B787_ | new_B788_;
  assign new_B782_ = ~new_B727_ & new_B741_;
  assign new_B781_ = new_B785_ | new_B786_;
  assign new_B780_ = ~new_B756_ & ~new_B776_;
  assign new_B779_ = new_B756_ & new_B776_;
  assign new_B778_ = ~new_B723_ | ~new_B748_;
  assign new_B777_ = new_B741_ & new_B778_;
  assign new_B776_ = new_B724_ | new_B725_;
  assign new_B775_ = new_B724_ | new_B741_;
  assign new_B774_ = ~new_B741_ & ~new_B777_;
  assign new_B773_ = new_B741_ | new_B778_;
  assign new_B772_ = new_B724_ & ~new_B725_;
  assign new_B771_ = ~new_B724_ & new_B725_;
  assign new_B770_ = new_B734_ | new_B767_;
  assign new_B769_ = ~new_B734_ & ~new_B768_;
  assign new_B768_ = new_B734_ & new_B767_;
  assign new_B767_ = ~new_B723_ | ~new_B748_;
  assign new_B766_ = ~new_B724_ & new_B734_;
  assign new_B765_ = new_B724_ & ~new_B734_;
  assign new_B764_ = new_B726_ & new_B763_;
  assign new_B763_ = new_B782_ | new_B781_;
  assign new_B762_ = ~new_B726_ & new_B761_;
  assign new_B761_ = new_B784_ | new_B783_;
  assign new_B760_ = new_B726_ | new_B759_;
  assign new_B759_ = new_B780_ | new_B779_;
  assign new_B758_ = ~new_B738_ & ~new_B748_;
  assign new_B757_ = new_B738_ & new_B748_;
  assign new_B756_ = ~new_B738_ | new_B748_;
  assign new_B755_ = new_B722_ & ~new_B723_;
  assign new_B754_ = ~new_B722_ & new_B723_;
  assign new_B753_ = new_B775_ & ~new_B776_;
  assign new_B752_ = ~new_B775_ & new_B776_;
  assign new_B751_ = ~new_B774_ | ~new_B773_;
  assign new_B750_ = new_B766_ | new_B765_;
  assign new_B749_ = new_B772_ | new_B771_;
  assign new_B748_ = new_B762_ | new_B764_;
  assign new_B747_ = ~new_B769_ | ~new_B770_;
  assign new_B746_ = new_B722_ & ~new_B723_;
  assign new_B745_ = new_B736_ & ~new_B748_;
  assign new_B744_ = ~new_B736_ & new_B748_;
  assign new_B743_ = ~new_B734_ & new_B760_;
  assign new_B742_ = new_B758_ | new_B757_;
  assign new_B741_ = new_B755_ | new_B754_;
  assign new_B740_ = new_B723_ | new_B756_;
  assign new_B739_ = new_B748_ & new_B751_;
  assign new_B738_ = new_B753_ | new_B752_;
  assign new_B737_ = new_B748_ & new_B747_;
  assign new_B736_ = new_B750_ & new_B749_;
  assign new_B735_ = new_B745_ | new_B744_;
  assign new_B734_ = new_B723_ | new_B746_;
  assign B733 = new_B734_ | new_B743_;
  assign B732 = new_B741_ & new_B742_;
  assign B731 = new_B741_ & new_B740_;
  assign B730 = new_B739_ | new_B738_;
  assign B729 = new_B737_ | new_B736_;
  assign B728 = new_B735_ & new_B734_;
  assign new_B727_ = new_C4465_;
  assign new_B726_ = new_C4398_;
  assign new_B725_ = new_C4331_;
  assign new_B724_ = new_C4264_;
  assign new_B723_ = new_C4197_;
  assign new_B722_ = new_C4130_;
  assign new_B721_ = ~new_B660_ & new_B674_;
  assign new_B720_ = new_B660_ & ~new_B674_;
  assign new_B719_ = new_B660_ & ~new_B674_;
  assign new_B718_ = ~new_B660_ & ~new_B674_;
  assign new_B717_ = new_B660_ & new_B674_;
  assign new_B716_ = new_B720_ | new_B721_;
  assign new_B715_ = ~new_B660_ & new_B674_;
  assign new_B714_ = new_B718_ | new_B719_;
  assign new_B713_ = ~new_B689_ & ~new_B709_;
  assign new_B712_ = new_B689_ & new_B709_;
  assign new_B711_ = ~new_B656_ | ~new_B681_;
  assign new_B710_ = new_B674_ & new_B711_;
  assign new_B709_ = new_B657_ | new_B658_;
  assign new_B708_ = new_B657_ | new_B674_;
  assign new_B707_ = ~new_B674_ & ~new_B710_;
  assign new_B706_ = new_B674_ | new_B711_;
  assign new_B705_ = new_B657_ & ~new_B658_;
  assign new_B704_ = ~new_B657_ & new_B658_;
  assign new_B703_ = new_B667_ | new_B700_;
  assign new_B702_ = ~new_B667_ & ~new_B701_;
  assign new_B701_ = new_B667_ & new_B700_;
  assign new_B700_ = ~new_B656_ | ~new_B681_;
  assign new_B699_ = ~new_B657_ & new_B667_;
  assign new_B698_ = new_B657_ & ~new_B667_;
  assign new_B697_ = new_B659_ & new_B696_;
  assign new_B696_ = new_B715_ | new_B714_;
  assign new_B695_ = ~new_B659_ & new_B694_;
  assign new_B694_ = new_B717_ | new_B716_;
  assign new_B693_ = new_B659_ | new_B692_;
  assign new_B692_ = new_B713_ | new_B712_;
  assign new_B691_ = ~new_B671_ & ~new_B681_;
  assign new_B690_ = new_B671_ & new_B681_;
  assign new_B689_ = ~new_B671_ | new_B681_;
  assign new_B688_ = new_B655_ & ~new_B656_;
  assign new_B687_ = ~new_B655_ & new_B656_;
  assign new_B686_ = new_B708_ & ~new_B709_;
  assign new_B685_ = ~new_B708_ & new_B709_;
  assign new_B684_ = ~new_B707_ | ~new_B706_;
  assign new_B683_ = new_B699_ | new_B698_;
  assign new_B682_ = new_B705_ | new_B704_;
  assign new_B681_ = new_B695_ | new_B697_;
  assign new_B680_ = ~new_B702_ | ~new_B703_;
  assign new_B679_ = new_B655_ & ~new_B656_;
  assign new_B678_ = new_B669_ & ~new_B681_;
  assign new_B677_ = ~new_B669_ & new_B681_;
  assign new_B676_ = ~new_B667_ & new_B693_;
  assign new_B675_ = new_B691_ | new_B690_;
  assign new_B674_ = new_B688_ | new_B687_;
  assign new_B673_ = new_B656_ | new_B689_;
  assign new_B672_ = new_B681_ & new_B684_;
  assign new_B671_ = new_B686_ | new_B685_;
  assign new_B670_ = new_B681_ & new_B680_;
  assign new_B669_ = new_B683_ & new_B682_;
  assign new_B668_ = new_B678_ | new_B677_;
  assign new_B667_ = new_B656_ | new_B679_;
  assign B666 = new_B667_ | new_B676_;
  assign B665 = new_B674_ & new_B675_;
  assign B664 = new_B674_ & new_B673_;
  assign B663 = new_B672_ | new_B671_;
  assign B662 = new_B670_ | new_B669_;
  assign B661 = new_B668_ & new_B667_;
  assign new_B660_ = new_C4063_;
  assign new_B659_ = new_C3996_;
  assign new_B658_ = new_C3929_;
  assign new_B657_ = new_C3862_;
  assign new_B656_ = new_C3795_;
  assign new_B655_ = new_C3728_;
  assign new_B654_ = ~new_B593_ & new_B607_;
  assign new_B653_ = new_B593_ & ~new_B607_;
  assign new_B652_ = new_B593_ & ~new_B607_;
  assign new_B651_ = ~new_B593_ & ~new_B607_;
  assign new_B650_ = new_B593_ & new_B607_;
  assign new_B649_ = new_B653_ | new_B654_;
  assign new_B648_ = ~new_B593_ & new_B607_;
  assign new_B647_ = new_B651_ | new_B652_;
  assign new_B646_ = ~new_B622_ & ~new_B642_;
  assign new_B645_ = new_B622_ & new_B642_;
  assign new_B644_ = ~new_B589_ | ~new_B614_;
  assign new_B643_ = new_B607_ & new_B644_;
  assign new_B642_ = new_B590_ | new_B591_;
  assign new_B641_ = new_B590_ | new_B607_;
  assign new_B640_ = ~new_B607_ & ~new_B643_;
  assign new_B639_ = new_B607_ | new_B644_;
  assign new_B638_ = new_B590_ & ~new_B591_;
  assign new_B637_ = ~new_B590_ & new_B591_;
  assign new_B636_ = new_B600_ | new_B633_;
  assign new_B635_ = ~new_B600_ & ~new_B634_;
  assign new_B634_ = new_B600_ & new_B633_;
  assign new_B633_ = ~new_B589_ | ~new_B614_;
  assign new_B632_ = ~new_B590_ & new_B600_;
  assign new_B631_ = new_B590_ & ~new_B600_;
  assign new_B630_ = new_B592_ & new_B629_;
  assign new_B629_ = new_B648_ | new_B647_;
  assign new_B628_ = ~new_B592_ & new_B627_;
  assign new_B627_ = new_B650_ | new_B649_;
  assign new_B626_ = new_B592_ | new_B625_;
  assign new_B625_ = new_B646_ | new_B645_;
  assign new_B624_ = ~new_B604_ & ~new_B614_;
  assign new_B623_ = new_B604_ & new_B614_;
  assign new_B622_ = ~new_B604_ | new_B614_;
  assign new_B621_ = new_B588_ & ~new_B589_;
  assign new_B620_ = ~new_B588_ & new_B589_;
  assign new_B619_ = new_B641_ & ~new_B642_;
  assign new_B618_ = ~new_B641_ & new_B642_;
  assign new_B617_ = ~new_B640_ | ~new_B639_;
  assign new_B616_ = new_B632_ | new_B631_;
  assign new_B615_ = new_B638_ | new_B637_;
  assign new_B614_ = new_B628_ | new_B630_;
  assign new_B613_ = ~new_B635_ | ~new_B636_;
  assign new_B612_ = new_B588_ & ~new_B589_;
  assign new_B611_ = new_B602_ & ~new_B614_;
  assign new_B610_ = ~new_B602_ & new_B614_;
  assign new_B609_ = ~new_B600_ & new_B626_;
  assign new_B608_ = new_B624_ | new_B623_;
  assign new_B607_ = new_B621_ | new_B620_;
  assign new_B606_ = new_B589_ | new_B622_;
  assign new_B605_ = new_B614_ & new_B617_;
  assign new_B604_ = new_B619_ | new_B618_;
  assign new_B603_ = new_B614_ & new_B613_;
  assign new_B602_ = new_B616_ & new_B615_;
  assign new_B601_ = new_B611_ | new_B610_;
  assign new_B600_ = new_B589_ | new_B612_;
  assign B599 = new_B600_ | new_B609_;
  assign B598 = new_B607_ & new_B608_;
  assign B597 = new_B607_ & new_B606_;
  assign B596 = new_B605_ | new_B604_;
  assign B595 = new_B603_ | new_B602_;
  assign B594 = new_B601_ & new_B600_;
  assign new_B593_ = new_C3661_;
  assign new_B592_ = new_C3594_;
  assign new_B591_ = new_C3527_;
  assign new_B590_ = new_C3460_;
  assign new_B589_ = new_C3393_;
  assign new_B588_ = new_C3326_;
  assign new_B587_ = ~new_B526_ & new_B540_;
  assign new_B586_ = new_B526_ & ~new_B540_;
  assign new_B585_ = new_B526_ & ~new_B540_;
  assign new_B584_ = ~new_B526_ & ~new_B540_;
  assign new_B583_ = new_B526_ & new_B540_;
  assign new_B582_ = new_B586_ | new_B587_;
  assign new_B581_ = ~new_B526_ & new_B540_;
  assign new_B580_ = new_B584_ | new_B585_;
  assign new_B579_ = ~new_B555_ & ~new_B575_;
  assign new_B578_ = new_B555_ & new_B575_;
  assign new_B577_ = ~new_B522_ | ~new_B547_;
  assign new_B576_ = new_B540_ & new_B577_;
  assign new_B575_ = new_B523_ | new_B524_;
  assign new_B574_ = new_B523_ | new_B540_;
  assign new_B573_ = ~new_B540_ & ~new_B576_;
  assign new_B572_ = new_B540_ | new_B577_;
  assign new_B571_ = new_B523_ & ~new_B524_;
  assign new_B570_ = ~new_B523_ & new_B524_;
  assign new_B569_ = new_B533_ | new_B566_;
  assign new_B568_ = ~new_B533_ & ~new_B567_;
  assign new_B567_ = new_B533_ & new_B566_;
  assign new_B566_ = ~new_B522_ | ~new_B547_;
  assign new_B565_ = ~new_B523_ & new_B533_;
  assign new_B564_ = new_B523_ & ~new_B533_;
  assign new_B563_ = new_B525_ & new_B562_;
  assign new_B562_ = new_B581_ | new_B580_;
  assign new_B561_ = ~new_B525_ & new_B560_;
  assign new_B560_ = new_B583_ | new_B582_;
  assign new_B559_ = new_B525_ | new_B558_;
  assign new_B558_ = new_B579_ | new_B578_;
  assign new_B557_ = ~new_B537_ & ~new_B547_;
  assign new_B556_ = new_B537_ & new_B547_;
  assign new_B555_ = ~new_B537_ | new_B547_;
  assign new_B554_ = new_B521_ & ~new_B522_;
  assign new_B553_ = ~new_B521_ & new_B522_;
  assign new_B552_ = new_B574_ & ~new_B575_;
  assign new_B551_ = ~new_B574_ & new_B575_;
  assign new_B550_ = ~new_B573_ | ~new_B572_;
  assign new_B549_ = new_B565_ | new_B564_;
  assign new_B548_ = new_B571_ | new_B570_;
  assign new_B547_ = new_B561_ | new_B563_;
  assign new_B546_ = ~new_B568_ | ~new_B569_;
  assign new_B545_ = new_B521_ & ~new_B522_;
  assign new_B544_ = new_B535_ & ~new_B547_;
  assign new_B543_ = ~new_B535_ & new_B547_;
  assign new_B542_ = ~new_B533_ & new_B559_;
  assign new_B541_ = new_B557_ | new_B556_;
  assign new_B540_ = new_B554_ | new_B553_;
  assign new_B539_ = new_B522_ | new_B555_;
  assign new_B538_ = new_B547_ & new_B550_;
  assign new_B537_ = new_B552_ | new_B551_;
  assign new_B536_ = new_B547_ & new_B546_;
  assign new_B535_ = new_B549_ & new_B548_;
  assign new_B534_ = new_B544_ | new_B543_;
  assign new_B533_ = new_B522_ | new_B545_;
  assign B532 = new_B533_ | new_B542_;
  assign B531 = new_B540_ & new_B541_;
  assign B530 = new_B540_ & new_B539_;
  assign B529 = new_B538_ | new_B537_;
  assign B528 = new_B536_ | new_B535_;
  assign B527 = new_B534_ & new_B533_;
  assign new_B526_ = new_C3259_;
  assign new_B525_ = new_C3192_;
  assign new_B524_ = new_C3125_;
  assign new_B523_ = new_C3058_;
  assign new_B522_ = new_C2991_;
  assign new_B521_ = new_C2924_;
  assign new_B520_ = ~new_B459_ & new_B473_;
  assign new_B519_ = new_B459_ & ~new_B473_;
  assign new_B518_ = new_B459_ & ~new_B473_;
  assign new_B517_ = ~new_B459_ & ~new_B473_;
  assign new_B516_ = new_B459_ & new_B473_;
  assign new_B515_ = new_B519_ | new_B520_;
  assign new_B514_ = ~new_B459_ & new_B473_;
  assign new_B513_ = new_B517_ | new_B518_;
  assign new_B512_ = ~new_B488_ & ~new_B508_;
  assign new_B511_ = new_B488_ & new_B508_;
  assign new_B510_ = ~new_B455_ | ~new_B480_;
  assign new_B509_ = new_B473_ & new_B510_;
  assign new_B508_ = new_B456_ | new_B457_;
  assign new_B507_ = new_B456_ | new_B473_;
  assign new_B506_ = ~new_B473_ & ~new_B509_;
  assign new_B505_ = new_B473_ | new_B510_;
  assign new_B504_ = new_B456_ & ~new_B457_;
  assign new_B503_ = ~new_B456_ & new_B457_;
  assign new_B502_ = new_B466_ | new_B499_;
  assign new_B501_ = ~new_B466_ & ~new_B500_;
  assign new_B500_ = new_B466_ & new_B499_;
  assign new_B499_ = ~new_B455_ | ~new_B480_;
  assign new_B498_ = ~new_B456_ & new_B466_;
  assign new_B497_ = new_B456_ & ~new_B466_;
  assign new_B496_ = new_B458_ & new_B495_;
  assign new_B495_ = new_B514_ | new_B513_;
  assign new_B494_ = ~new_B458_ & new_B493_;
  assign new_B493_ = new_B516_ | new_B515_;
  assign new_B492_ = new_B458_ | new_B491_;
  assign new_B491_ = new_B512_ | new_B511_;
  assign new_B490_ = ~new_B470_ & ~new_B480_;
  assign new_B489_ = new_B470_ & new_B480_;
  assign new_B488_ = ~new_B470_ | new_B480_;
  assign new_B487_ = new_B454_ & ~new_B455_;
  assign new_B486_ = ~new_B454_ & new_B455_;
  assign new_B485_ = new_B507_ & ~new_B508_;
  assign new_B484_ = ~new_B507_ & new_B508_;
  assign new_B483_ = ~new_B506_ | ~new_B505_;
  assign new_B482_ = new_B498_ | new_B497_;
  assign new_B481_ = new_B504_ | new_B503_;
  assign new_B480_ = new_B494_ | new_B496_;
  assign new_B479_ = ~new_B501_ | ~new_B502_;
  assign new_B478_ = new_B454_ & ~new_B455_;
  assign new_B477_ = new_B468_ & ~new_B480_;
  assign new_B476_ = ~new_B468_ & new_B480_;
  assign new_B475_ = ~new_B466_ & new_B492_;
  assign new_B474_ = new_B490_ | new_B489_;
  assign new_B473_ = new_B487_ | new_B486_;
  assign new_B472_ = new_B455_ | new_B488_;
  assign new_B471_ = new_B480_ & new_B483_;
  assign new_B470_ = new_B485_ | new_B484_;
  assign new_B469_ = new_B480_ & new_B479_;
  assign new_B468_ = new_B482_ & new_B481_;
  assign new_B467_ = new_B477_ | new_B476_;
  assign new_B466_ = new_B455_ | new_B478_;
  assign B465 = new_B466_ | new_B475_;
  assign B464 = new_B473_ & new_B474_;
  assign B463 = new_B473_ & new_B472_;
  assign B462 = new_B471_ | new_B470_;
  assign B461 = new_B469_ | new_B468_;
  assign B460 = new_B467_ & new_B466_;
  assign new_B459_ = new_C2857_;
  assign new_B458_ = new_C2790_;
  assign new_B457_ = new_C2723_;
  assign new_B456_ = new_C2656_;
  assign new_B455_ = new_C2589_;
  assign new_B454_ = new_C2525_;
  assign new_B453_ = ~new_B392_ & new_B406_;
  assign new_B452_ = new_B392_ & ~new_B406_;
  assign new_B451_ = new_B392_ & ~new_B406_;
  assign new_B450_ = ~new_B392_ & ~new_B406_;
  assign new_B449_ = new_B392_ & new_B406_;
  assign new_B448_ = new_B452_ | new_B453_;
  assign new_B447_ = ~new_B392_ & new_B406_;
  assign new_B446_ = new_B450_ | new_B451_;
  assign new_B445_ = ~new_B421_ & ~new_B441_;
  assign new_B444_ = new_B421_ & new_B441_;
  assign new_B443_ = ~new_B388_ | ~new_B413_;
  assign new_B442_ = new_B406_ & new_B443_;
  assign new_B441_ = new_B389_ | new_B390_;
  assign new_B440_ = new_B389_ | new_B406_;
  assign new_B439_ = ~new_B406_ & ~new_B442_;
  assign new_B438_ = new_B406_ | new_B443_;
  assign new_B437_ = new_B389_ & ~new_B390_;
  assign new_B436_ = ~new_B389_ & new_B390_;
  assign new_B435_ = new_B399_ | new_B432_;
  assign new_B434_ = ~new_B399_ & ~new_B433_;
  assign new_B433_ = new_B399_ & new_B432_;
  assign new_B432_ = ~new_B388_ | ~new_B413_;
  assign new_B431_ = ~new_B389_ & new_B399_;
  assign new_B430_ = new_B389_ & ~new_B399_;
  assign new_B429_ = new_B391_ & new_B428_;
  assign new_B428_ = new_B447_ | new_B446_;
  assign new_B427_ = ~new_B391_ & new_B426_;
  assign new_B426_ = new_B449_ | new_B448_;
  assign new_B425_ = new_B391_ | new_B424_;
  assign new_B424_ = new_B445_ | new_B444_;
  assign new_B423_ = ~new_B403_ & ~new_B413_;
  assign new_B422_ = new_B403_ & new_B413_;
  assign new_B421_ = ~new_B403_ | new_B413_;
  assign new_B420_ = new_B387_ & ~new_B388_;
  assign new_B419_ = ~new_B387_ & new_B388_;
  assign new_B418_ = new_B440_ & ~new_B441_;
  assign new_B417_ = ~new_B440_ & new_B441_;
  assign new_B416_ = ~new_B439_ | ~new_B438_;
  assign new_B415_ = new_B431_ | new_B430_;
  assign new_B414_ = new_B437_ | new_B436_;
  assign new_B413_ = new_B427_ | new_B429_;
  assign new_B412_ = ~new_B434_ | ~new_B435_;
  assign new_B411_ = new_B387_ & ~new_B388_;
  assign new_B410_ = new_B401_ & ~new_B413_;
  assign new_B409_ = ~new_B401_ & new_B413_;
  assign new_B408_ = ~new_B399_ & new_B425_;
  assign new_B407_ = new_B423_ | new_B422_;
  assign new_B406_ = new_B420_ | new_B419_;
  assign new_B405_ = new_B388_ | new_B421_;
  assign new_B404_ = new_B413_ & new_B416_;
  assign new_B403_ = new_B418_ | new_B417_;
  assign new_B402_ = new_B413_ & new_B412_;
  assign new_B401_ = new_B415_ & new_B414_;
  assign new_B400_ = new_B410_ | new_B409_;
  assign new_B399_ = new_B388_ | new_B411_;
  assign B398 = new_B399_ | new_B408_;
  assign B397 = new_B406_ & new_B407_;
  assign B396 = new_B406_ & new_B405_;
  assign B395 = new_B404_ | new_B403_;
  assign B394 = new_B402_ | new_B401_;
  assign B393 = new_B400_ & new_B399_;
  assign new_B392_ = new_D6927_;
  assign new_B391_ = new_D6860_;
  assign new_B390_ = new_D6793_;
  assign new_B389_ = new_D6726_;
  assign new_B388_ = new_D6659_;
  assign new_B387_ = new_D6592_;
  assign new_B386_ = ~new_B325_ & new_B339_;
  assign new_B385_ = new_B325_ & ~new_B339_;
  assign new_B384_ = new_B325_ & ~new_B339_;
  assign new_B383_ = ~new_B325_ & ~new_B339_;
  assign new_B382_ = new_B325_ & new_B339_;
  assign new_B381_ = new_B385_ | new_B386_;
  assign new_B380_ = ~new_B325_ & new_B339_;
  assign new_B379_ = new_B383_ | new_B384_;
  assign new_B378_ = ~new_B354_ & ~new_B374_;
  assign new_B377_ = new_B354_ & new_B374_;
  assign new_B376_ = ~new_B321_ | ~new_B346_;
  assign new_B375_ = new_B339_ & new_B376_;
  assign new_B374_ = new_B322_ | new_B323_;
  assign new_B373_ = new_B322_ | new_B339_;
  assign new_B372_ = ~new_B339_ & ~new_B375_;
  assign new_B371_ = new_B339_ | new_B376_;
  assign new_B370_ = new_B322_ & ~new_B323_;
  assign new_B369_ = ~new_B322_ & new_B323_;
  assign new_B368_ = new_B332_ | new_B365_;
  assign new_B367_ = ~new_B332_ & ~new_B366_;
  assign new_B366_ = new_B332_ & new_B365_;
  assign new_B365_ = ~new_B321_ | ~new_B346_;
  assign new_B364_ = ~new_B322_ & new_B332_;
  assign new_B363_ = new_B322_ & ~new_B332_;
  assign new_B362_ = new_B324_ & new_B361_;
  assign new_B361_ = new_B380_ | new_B379_;
  assign new_B360_ = ~new_B324_ & new_B359_;
  assign new_B359_ = new_B382_ | new_B381_;
  assign new_B358_ = new_B324_ | new_B357_;
  assign new_B357_ = new_B378_ | new_B377_;
  assign new_B356_ = ~new_B336_ & ~new_B346_;
  assign new_B355_ = new_B336_ & new_B346_;
  assign new_B354_ = ~new_B336_ | new_B346_;
  assign new_B353_ = new_B320_ & ~new_B321_;
  assign new_B352_ = ~new_B320_ & new_B321_;
  assign new_B351_ = new_B373_ & ~new_B374_;
  assign new_B350_ = ~new_B373_ & new_B374_;
  assign new_B349_ = ~new_B372_ | ~new_B371_;
  assign new_B348_ = new_B364_ | new_B363_;
  assign new_B347_ = new_B370_ | new_B369_;
  assign new_B346_ = new_B360_ | new_B362_;
  assign new_B345_ = ~new_B367_ | ~new_B368_;
  assign new_B344_ = new_B320_ & ~new_B321_;
  assign new_B343_ = new_B334_ & ~new_B346_;
  assign new_B342_ = ~new_B334_ & new_B346_;
  assign new_B341_ = ~new_B332_ & new_B358_;
  assign new_B340_ = new_B356_ | new_B355_;
  assign new_B339_ = new_B353_ | new_B352_;
  assign new_B338_ = new_B321_ | new_B354_;
  assign new_B337_ = new_B346_ & new_B349_;
  assign new_B336_ = new_B351_ | new_B350_;
  assign new_B335_ = new_B346_ & new_B345_;
  assign new_B334_ = new_B348_ & new_B347_;
  assign new_B333_ = new_B343_ | new_B342_;
  assign new_B332_ = new_B321_ | new_B344_;
  assign B331 = new_B332_ | new_B341_;
  assign B330 = new_B339_ & new_B340_;
  assign B329 = new_B339_ & new_B338_;
  assign B328 = new_B337_ | new_B336_;
  assign B327 = new_B335_ | new_B334_;
  assign B326 = new_B333_ & new_B332_;
  assign new_B325_ = new_D6525_;
  assign new_B324_ = new_D6458_;
  assign new_B323_ = new_D6391_;
  assign new_B322_ = new_D6324_;
  assign new_B321_ = new_D6257_;
  assign new_B320_ = new_D6190_;
  assign new_B319_ = ~new_B258_ & new_B272_;
  assign new_B318_ = new_B258_ & ~new_B272_;
  assign new_B317_ = new_B258_ & ~new_B272_;
  assign new_B316_ = ~new_B258_ & ~new_B272_;
  assign new_B315_ = new_B258_ & new_B272_;
  assign new_B314_ = new_B318_ | new_B319_;
  assign new_B313_ = ~new_B258_ & new_B272_;
  assign new_B312_ = new_B316_ | new_B317_;
  assign new_B311_ = ~new_B287_ & ~new_B307_;
  assign new_B310_ = new_B287_ & new_B307_;
  assign new_B309_ = ~new_B254_ | ~new_B279_;
  assign new_B308_ = new_B272_ & new_B309_;
  assign new_B307_ = new_B255_ | new_B256_;
  assign new_B306_ = new_B255_ | new_B272_;
  assign new_B305_ = ~new_B272_ & ~new_B308_;
  assign new_B304_ = new_B272_ | new_B309_;
  assign new_B303_ = new_B255_ & ~new_B256_;
  assign new_B302_ = ~new_B255_ & new_B256_;
  assign new_B301_ = new_B265_ | new_B298_;
  assign new_B300_ = ~new_B265_ & ~new_B299_;
  assign new_B299_ = new_B265_ & new_B298_;
  assign new_B298_ = ~new_B254_ | ~new_B279_;
  assign new_B297_ = ~new_B255_ & new_B265_;
  assign new_B296_ = new_B255_ & ~new_B265_;
  assign new_B295_ = new_B257_ & new_B294_;
  assign new_B294_ = new_B313_ | new_B312_;
  assign new_B293_ = ~new_B257_ & new_B292_;
  assign new_B292_ = new_B315_ | new_B314_;
  assign new_B291_ = new_B257_ | new_B290_;
  assign new_B290_ = new_B311_ | new_B310_;
  assign new_B289_ = ~new_B269_ & ~new_B279_;
  assign new_B288_ = new_B269_ & new_B279_;
  assign new_B287_ = ~new_B269_ | new_B279_;
  assign new_B286_ = new_B253_ & ~new_B254_;
  assign new_B285_ = ~new_B253_ & new_B254_;
  assign new_B284_ = new_B306_ & ~new_B307_;
  assign new_B283_ = ~new_B306_ & new_B307_;
  assign new_B282_ = ~new_B305_ | ~new_B304_;
  assign new_B281_ = new_B297_ | new_B296_;
  assign new_B280_ = new_B303_ | new_B302_;
  assign new_B279_ = new_B293_ | new_B295_;
  assign new_B278_ = ~new_B300_ | ~new_B301_;
  assign new_B277_ = new_B253_ & ~new_B254_;
  assign new_B276_ = new_B267_ & ~new_B279_;
  assign new_B275_ = ~new_B267_ & new_B279_;
  assign new_B274_ = ~new_B265_ & new_B291_;
  assign new_B273_ = new_B289_ | new_B288_;
  assign new_B272_ = new_B286_ | new_B285_;
  assign new_B271_ = new_B254_ | new_B287_;
  assign new_B270_ = new_B279_ & new_B282_;
  assign new_B269_ = new_B284_ | new_B283_;
  assign new_B268_ = new_B279_ & new_B278_;
  assign new_B267_ = new_B281_ & new_B280_;
  assign new_B266_ = new_B276_ | new_B275_;
  assign new_B265_ = new_B254_ | new_B277_;
  assign B264 = new_B265_ | new_B274_;
  assign B263 = new_B272_ & new_B273_;
  assign B262 = new_B272_ & new_B271_;
  assign B261 = new_B270_ | new_B269_;
  assign B260 = new_B268_ | new_B267_;
  assign B259 = new_B266_ & new_B265_;
  assign new_B258_ = new_D6123_;
  assign new_B257_ = new_D6056_;
  assign new_B256_ = new_D5989_;
  assign new_B255_ = new_D5922_;
  assign new_B254_ = new_D5855_;
  assign new_B253_ = new_D5788_;
  assign new_B252_ = ~new_B191_ & new_B205_;
  assign new_B251_ = new_B191_ & ~new_B205_;
  assign new_B250_ = new_B191_ & ~new_B205_;
  assign new_B249_ = ~new_B191_ & ~new_B205_;
  assign new_B248_ = new_B191_ & new_B205_;
  assign new_B247_ = new_B251_ | new_B252_;
  assign new_B246_ = ~new_B191_ & new_B205_;
  assign new_B245_ = new_B249_ | new_B250_;
  assign new_B244_ = ~new_B220_ & ~new_B240_;
  assign new_B243_ = new_B220_ & new_B240_;
  assign new_B242_ = ~new_B187_ | ~new_B212_;
  assign new_B241_ = new_B205_ & new_B242_;
  assign new_B240_ = new_B188_ | new_B189_;
  assign new_B239_ = new_B188_ | new_B205_;
  assign new_B238_ = ~new_B205_ & ~new_B241_;
  assign new_B237_ = new_B205_ | new_B242_;
  assign new_B236_ = new_B188_ & ~new_B189_;
  assign new_B235_ = ~new_B188_ & new_B189_;
  assign new_B234_ = new_B198_ | new_B231_;
  assign new_B233_ = ~new_B198_ & ~new_B232_;
  assign new_B232_ = new_B198_ & new_B231_;
  assign new_B231_ = ~new_B187_ | ~new_B212_;
  assign new_B230_ = ~new_B188_ & new_B198_;
  assign new_B229_ = new_B188_ & ~new_B198_;
  assign new_B228_ = new_B190_ & new_B227_;
  assign new_B227_ = new_B246_ | new_B245_;
  assign new_B226_ = ~new_B190_ & new_B225_;
  assign new_B225_ = new_B248_ | new_B247_;
  assign new_B224_ = new_B190_ | new_B223_;
  assign new_B223_ = new_B244_ | new_B243_;
  assign new_B222_ = ~new_B202_ & ~new_B212_;
  assign new_B221_ = new_B202_ & new_B212_;
  assign new_B220_ = ~new_B202_ | new_B212_;
  assign new_B219_ = new_B186_ & ~new_B187_;
  assign new_B218_ = ~new_B186_ & new_B187_;
  assign new_B217_ = new_B239_ & ~new_B240_;
  assign new_B216_ = ~new_B239_ & new_B240_;
  assign new_B215_ = ~new_B238_ | ~new_B237_;
  assign new_B214_ = new_B230_ | new_B229_;
  assign new_B213_ = new_B236_ | new_B235_;
  assign new_B212_ = new_B226_ | new_B228_;
  assign new_B211_ = ~new_B233_ | ~new_B234_;
  assign new_B210_ = new_B186_ & ~new_B187_;
  assign new_B209_ = new_B200_ & ~new_B212_;
  assign new_B208_ = ~new_B200_ & new_B212_;
  assign new_B207_ = ~new_B198_ & new_B224_;
  assign new_B206_ = new_B222_ | new_B221_;
  assign new_B205_ = new_B219_ | new_B218_;
  assign new_B204_ = new_B187_ | new_B220_;
  assign new_B203_ = new_B212_ & new_B215_;
  assign new_B202_ = new_B217_ | new_B216_;
  assign new_B201_ = new_B212_ & new_B211_;
  assign new_B200_ = new_B214_ & new_B213_;
  assign new_B199_ = new_B209_ | new_B208_;
  assign new_B198_ = new_B187_ | new_B210_;
  assign B197 = new_B198_ | new_B207_;
  assign B196 = new_B205_ & new_B206_;
  assign B195 = new_B205_ & new_B204_;
  assign B194 = new_B203_ | new_B202_;
  assign B193 = new_B201_ | new_B200_;
  assign B192 = new_B199_ & new_B198_;
  assign new_B191_ = new_D5721_;
  assign new_B190_ = new_D5654_;
  assign new_B189_ = new_D5587_;
  assign new_B188_ = new_D5520_;
  assign new_B187_ = new_D5453_;
  assign new_B186_ = new_D5386_;
  assign new_B185_ = ~new_B124_ & new_B138_;
  assign new_B184_ = new_B124_ & ~new_B138_;
  assign new_B183_ = new_B124_ & ~new_B138_;
  assign new_B182_ = ~new_B124_ & ~new_B138_;
  assign new_B181_ = new_B124_ & new_B138_;
  assign new_B180_ = new_B184_ | new_B185_;
  assign new_B179_ = ~new_B124_ & new_B138_;
  assign new_B178_ = new_B182_ | new_B183_;
  assign new_B177_ = ~new_B153_ & ~new_B173_;
  assign new_B176_ = new_B153_ & new_B173_;
  assign new_B175_ = ~new_B120_ | ~new_B145_;
  assign new_B174_ = new_B138_ & new_B175_;
  assign new_B173_ = new_B121_ | new_B122_;
  assign new_B172_ = new_B121_ | new_B138_;
  assign new_B171_ = ~new_B138_ & ~new_B174_;
  assign new_B170_ = new_B138_ | new_B175_;
  assign new_B169_ = new_B121_ & ~new_B122_;
  assign new_B168_ = ~new_B121_ & new_B122_;
  assign new_B167_ = new_B131_ | new_B164_;
  assign new_B166_ = ~new_B131_ & ~new_B165_;
  assign new_B165_ = new_B131_ & new_B164_;
  assign new_B164_ = ~new_B120_ | ~new_B145_;
  assign new_B163_ = ~new_B121_ & new_B131_;
  assign new_B162_ = new_B121_ & ~new_B131_;
  assign new_B161_ = new_B123_ & new_B160_;
  assign new_B160_ = new_B179_ | new_B178_;
  assign new_B159_ = ~new_B123_ & new_B158_;
  assign new_B158_ = new_B181_ | new_B180_;
  assign new_B157_ = new_B123_ | new_B156_;
  assign new_B156_ = new_B177_ | new_B176_;
  assign new_B155_ = ~new_B135_ & ~new_B145_;
  assign new_B154_ = new_B135_ & new_B145_;
  assign new_B153_ = ~new_B135_ | new_B145_;
  assign new_B152_ = new_B119_ & ~new_B120_;
  assign new_B151_ = ~new_B119_ & new_B120_;
  assign new_B150_ = new_B172_ & ~new_B173_;
  assign new_B149_ = ~new_B172_ & new_B173_;
  assign new_B148_ = ~new_B171_ | ~new_B170_;
  assign new_B147_ = new_B163_ | new_B162_;
  assign new_B146_ = new_B169_ | new_B168_;
  assign new_B145_ = new_B159_ | new_B161_;
  assign new_B144_ = ~new_B166_ | ~new_B167_;
  assign new_B143_ = new_B119_ & ~new_B120_;
  assign new_B142_ = new_B133_ & ~new_B145_;
  assign new_B141_ = ~new_B133_ & new_B145_;
  assign new_B140_ = ~new_B131_ & new_B157_;
  assign new_B139_ = new_B155_ | new_B154_;
  assign new_B138_ = new_B152_ | new_B151_;
  assign new_B137_ = new_B120_ | new_B153_;
  assign new_B136_ = new_B145_ & new_B148_;
  assign new_B135_ = new_B150_ | new_B149_;
  assign new_B134_ = new_B145_ & new_B144_;
  assign new_B133_ = new_B147_ & new_B146_;
  assign new_B132_ = new_B142_ | new_B141_;
  assign new_B131_ = new_B120_ | new_B143_;
  assign B130 = new_B131_ | new_B140_;
  assign B129 = new_B138_ & new_B139_;
  assign B128 = new_B138_ & new_B137_;
  assign B127 = new_B136_ | new_B135_;
  assign B126 = new_B134_ | new_B133_;
  assign B125 = new_B132_ & new_B131_;
  assign new_B124_ = new_D5319_;
  assign new_B123_ = new_D5252_;
  assign new_B122_ = new_D5185_;
  assign new_B121_ = new_D5118_;
  assign new_B120_ = new_D5051_;
  assign new_B119_ = new_D4984_;
  assign new_B118_ = ~new_B57_ & new_B71_;
  assign new_B117_ = new_B57_ & ~new_B71_;
  assign new_B116_ = new_B57_ & ~new_B71_;
  assign new_B115_ = ~new_B57_ & ~new_B71_;
  assign new_B114_ = new_B57_ & new_B71_;
  assign new_B113_ = new_B117_ | new_B118_;
  assign new_B112_ = ~new_B57_ & new_B71_;
  assign new_B111_ = new_B115_ | new_B116_;
  assign new_B110_ = ~new_B86_ & ~new_B106_;
  assign new_B109_ = new_B86_ & new_B106_;
  assign new_B108_ = ~new_B53_ | ~new_B78_;
  assign new_B107_ = new_B71_ & new_B108_;
  assign new_B106_ = new_B54_ | new_B55_;
  assign new_B105_ = new_B54_ | new_B71_;
  assign new_B104_ = ~new_B71_ & ~new_B107_;
  assign new_B103_ = new_B71_ | new_B108_;
  assign new_B102_ = new_B54_ & ~new_B55_;
  assign new_B101_ = ~new_B54_ & new_B55_;
  assign new_B100_ = new_B64_ | new_B97_;
  assign new_B99_ = ~new_B64_ & ~new_B98_;
  assign new_B98_ = new_B64_ & new_B97_;
  assign new_B97_ = ~new_B53_ | ~new_B78_;
  assign new_B96_ = ~new_B54_ & new_B64_;
  assign new_B95_ = new_B54_ & ~new_B64_;
  assign new_B94_ = new_B56_ & new_B93_;
  assign new_B93_ = new_B112_ | new_B111_;
  assign new_B92_ = ~new_B56_ & new_B91_;
  assign new_B91_ = new_B114_ | new_B113_;
  assign new_B90_ = new_B56_ | new_B89_;
  assign new_B89_ = new_B110_ | new_B109_;
  assign new_B88_ = ~new_B68_ & ~new_B78_;
  assign new_B87_ = new_B68_ & new_B78_;
  assign new_B86_ = ~new_B68_ | new_B78_;
  assign new_B85_ = new_B52_ & ~new_B53_;
  assign new_B84_ = ~new_B52_ & new_B53_;
  assign new_B83_ = new_B105_ & ~new_B106_;
  assign new_B82_ = ~new_B105_ & new_B106_;
  assign new_B81_ = ~new_B104_ | ~new_B103_;
  assign new_B80_ = new_B96_ | new_B95_;
  assign new_B79_ = new_B102_ | new_B101_;
  assign new_B78_ = new_B92_ | new_B94_;
  assign new_B77_ = ~new_B99_ | ~new_B100_;
  assign new_B76_ = new_B52_ & ~new_B53_;
  assign new_B75_ = new_B66_ & ~new_B78_;
  assign new_B74_ = ~new_B66_ & new_B78_;
  assign new_B73_ = ~new_B64_ & new_B90_;
  assign new_B72_ = new_B88_ | new_B87_;
  assign new_B71_ = new_B85_ | new_B84_;
  assign new_B70_ = new_B53_ | new_B86_;
  assign new_B69_ = new_B78_ & new_B81_;
  assign new_B68_ = new_B83_ | new_B82_;
  assign new_B67_ = new_B78_ & new_B77_;
  assign new_B66_ = new_B80_ & new_B79_;
  assign new_B65_ = new_B75_ | new_B74_;
  assign new_B64_ = new_B53_ | new_B76_;
  assign B63 = new_B64_ | new_B73_;
  assign B62 = new_B71_ & new_B72_;
  assign B61 = new_B71_ & new_B70_;
  assign B60 = new_B69_ | new_B68_;
  assign B59 = new_B67_ | new_B66_;
  assign B58 = new_B65_ & new_B64_;
  assign new_B57_ = new_D4917_;
  assign new_B56_ = new_D4850_;
  assign new_B55_ = new_D4783_;
  assign new_B54_ = new_D4716_;
  assign new_B53_ = new_D4649_;
  assign new_B52_ = new_D4582_;
  assign new_B51_ = ~new_A9989_ & new_B4_;
  assign new_B50_ = new_A9989_ & ~new_B4_;
  assign new_B49_ = new_A9989_ & ~new_B4_;
  assign new_B48_ = ~new_A9989_ & ~new_B4_;
  assign new_B47_ = new_A9989_ & new_B4_;
  assign new_B46_ = new_B50_ | new_B51_;
  assign new_B45_ = ~new_A9989_ & new_B4_;
  assign new_B44_ = new_B48_ | new_B49_;
  assign new_B43_ = ~new_B19_ & ~new_B39_;
  assign new_B42_ = new_B19_ & new_B39_;
  assign new_B41_ = ~new_A9985_ | ~new_B11_;
  assign new_B40_ = new_B4_ & new_B41_;
  assign new_B39_ = new_A9986_ | new_A9987_;
  assign new_B38_ = new_A9986_ | new_B4_;
  assign new_B37_ = ~new_B4_ & ~new_B40_;
  assign new_B36_ = new_B4_ | new_B41_;
  assign new_B35_ = new_A9986_ & ~new_A9987_;
  assign new_B34_ = ~new_A9986_ & new_A9987_;
  assign new_B33_ = new_A9996_ | new_B30_;
  assign new_B32_ = ~new_A9996_ & ~new_B31_;
  assign new_B31_ = new_A9996_ & new_B30_;
  assign new_B30_ = ~new_A9985_ | ~new_B11_;
  assign new_B29_ = ~new_A9986_ & new_A9996_;
  assign new_B28_ = new_A9986_ & ~new_A9996_;
  assign new_B27_ = new_A9988_ & new_B26_;
  assign new_B26_ = new_B45_ | new_B44_;
  assign new_B25_ = ~new_A9988_ & new_B24_;
  assign new_B24_ = new_B47_ | new_B46_;
  assign new_B23_ = new_A9988_ | new_B22_;
  assign new_B22_ = new_B43_ | new_B42_;
  assign new_B21_ = ~new_B1_ & ~new_B11_;
  assign new_B20_ = new_B1_ & new_B11_;
  assign new_B19_ = ~new_B1_ | new_B11_;
  assign new_B18_ = new_A9984_ & ~new_A9985_;
  assign new_B17_ = ~new_A9984_ & new_A9985_;
  assign new_B16_ = new_B38_ & ~new_B39_;
  assign new_B15_ = ~new_B38_ & new_B39_;
  assign new_B14_ = ~new_B37_ | ~new_B36_;
  assign new_B13_ = new_B29_ | new_B28_;
  assign new_B12_ = new_B35_ | new_B34_;
  assign new_B11_ = new_B25_ | new_B27_;
  assign new_B10_ = ~new_B32_ | ~new_B33_;
  assign new_B9_ = new_A9984_ & ~new_A9985_;
  assign new_B8_ = new_A9998_ & ~new_B11_;
  assign new_B7_ = ~new_A9998_ & new_B11_;
  assign new_B6_ = ~new_A9996_ & new_B23_;
  assign new_B5_ = new_B21_ | new_B20_;
  assign new_B4_ = new_B18_ | new_B17_;
  assign new_B3_ = new_A9985_ | new_B19_;
  assign new_B2_ = new_B11_ & new_B14_;
  assign new_B1_ = new_B16_ | new_B15_;
  assign new_A9999_ = new_B11_ & new_B10_;
  assign new_A9998_ = new_B13_ & new_B12_;
  assign new_A9997_ = new_B8_ | new_B7_;
  assign new_A9996_ = new_A9985_ | new_B9_;
  assign A9995 = new_A9996_ | new_B6_;
  assign A9994 = new_B4_ & new_B5_;
  assign A9993 = new_B4_ & new_B3_;
  assign A9992 = new_B2_ | new_B1_;
  assign A9991 = new_A9999_ | new_A9998_;
  assign A9990 = new_A9997_ & new_A9996_;
  assign new_A9989_ = new_D4515_;
  assign new_A9988_ = new_D4448_;
  assign new_A9987_ = new_D4381_;
  assign new_A9986_ = new_D4314_;
  assign new_A9985_ = new_D4247_;
  assign new_A9984_ = new_D4180_;
  assign new_A9983_ = ~new_A9922_ & new_A9936_;
  assign new_A9982_ = new_A9922_ & ~new_A9936_;
  assign new_A9981_ = new_A9922_ & ~new_A9936_;
  assign new_A9980_ = ~new_A9922_ & ~new_A9936_;
  assign new_A9979_ = new_A9922_ & new_A9936_;
  assign new_A9978_ = new_A9982_ | new_A9983_;
  assign new_A9977_ = ~new_A9922_ & new_A9936_;
  assign new_A9976_ = new_A9980_ | new_A9981_;
  assign new_A9975_ = ~new_A9951_ & ~new_A9971_;
  assign new_A9974_ = new_A9951_ & new_A9971_;
  assign new_A9973_ = ~new_A9918_ | ~new_A9943_;
  assign new_A9972_ = new_A9936_ & new_A9973_;
  assign new_A9971_ = new_A9919_ | new_A9920_;
  assign new_A9970_ = new_A9919_ | new_A9936_;
  assign new_A9969_ = ~new_A9936_ & ~new_A9972_;
  assign new_A9968_ = new_A9936_ | new_A9973_;
  assign new_A9967_ = new_A9919_ & ~new_A9920_;
  assign new_A9966_ = ~new_A9919_ & new_A9920_;
  assign new_A9965_ = new_A9929_ | new_A9962_;
  assign new_A9964_ = ~new_A9929_ & ~new_A9963_;
  assign new_A9963_ = new_A9929_ & new_A9962_;
  assign new_A9962_ = ~new_A9918_ | ~new_A9943_;
  assign new_A9961_ = ~new_A9919_ & new_A9929_;
  assign new_A9960_ = new_A9919_ & ~new_A9929_;
  assign new_A9959_ = new_A9921_ & new_A9958_;
  assign new_A9958_ = new_A9977_ | new_A9976_;
  assign new_A9957_ = ~new_A9921_ & new_A9956_;
  assign new_A9956_ = new_A9979_ | new_A9978_;
  assign new_A9955_ = new_A9921_ | new_A9954_;
  assign new_A9954_ = new_A9975_ | new_A9974_;
  assign new_A9953_ = ~new_A9933_ & ~new_A9943_;
  assign new_A9952_ = new_A9933_ & new_A9943_;
  assign new_A9951_ = ~new_A9933_ | new_A9943_;
  assign new_A9950_ = new_A9917_ & ~new_A9918_;
  assign new_A9949_ = ~new_A9917_ & new_A9918_;
  assign new_A9948_ = new_A9970_ & ~new_A9971_;
  assign new_A9947_ = ~new_A9970_ & new_A9971_;
  assign new_A9946_ = ~new_A9969_ | ~new_A9968_;
  assign new_A9945_ = new_A9961_ | new_A9960_;
  assign new_A9944_ = new_A9967_ | new_A9966_;
  assign new_A9943_ = new_A9957_ | new_A9959_;
  assign new_A9942_ = ~new_A9964_ | ~new_A9965_;
  assign new_A9941_ = new_A9917_ & ~new_A9918_;
  assign new_A9940_ = new_A9931_ & ~new_A9943_;
  assign new_A9939_ = ~new_A9931_ & new_A9943_;
  assign new_A9938_ = ~new_A9929_ & new_A9955_;
  assign new_A9937_ = new_A9953_ | new_A9952_;
  assign new_A9936_ = new_A9950_ | new_A9949_;
  assign new_A9935_ = new_A9918_ | new_A9951_;
  assign new_A9934_ = new_A9943_ & new_A9946_;
  assign new_A9933_ = new_A9948_ | new_A9947_;
  assign new_A9932_ = new_A9943_ & new_A9942_;
  assign new_A9931_ = new_A9945_ & new_A9944_;
  assign new_A9930_ = new_A9940_ | new_A9939_;
  assign new_A9929_ = new_A9918_ | new_A9941_;
  assign A9928 = new_A9929_ | new_A9938_;
  assign A9927 = new_A9936_ & new_A9937_;
  assign A9926 = new_A9936_ & new_A9935_;
  assign A9925 = new_A9934_ | new_A9933_;
  assign A9924 = new_A9932_ | new_A9931_;
  assign A9923 = new_A9930_ & new_A9929_;
  assign new_A9922_ = new_D4113_;
  assign new_A9921_ = new_D4046_;
  assign new_A9920_ = new_D3979_;
  assign new_A9919_ = new_D3912_;
  assign new_A9918_ = new_D3845_;
  assign new_A9917_ = new_D3778_;
  assign new_A9916_ = ~new_A9855_ & new_A9869_;
  assign new_A9915_ = new_A9855_ & ~new_A9869_;
  assign new_A9914_ = new_A9855_ & ~new_A9869_;
  assign new_A9913_ = ~new_A9855_ & ~new_A9869_;
  assign new_A9912_ = new_A9855_ & new_A9869_;
  assign new_A9911_ = new_A9915_ | new_A9916_;
  assign new_A9910_ = ~new_A9855_ & new_A9869_;
  assign new_A9909_ = new_A9913_ | new_A9914_;
  assign new_A9908_ = ~new_A9884_ & ~new_A9904_;
  assign new_A9907_ = new_A9884_ & new_A9904_;
  assign new_A9906_ = ~new_A9851_ | ~new_A9876_;
  assign new_A9905_ = new_A9869_ & new_A9906_;
  assign new_A9904_ = new_A9852_ | new_A9853_;
  assign new_A9903_ = new_A9852_ | new_A9869_;
  assign new_A9902_ = ~new_A9869_ & ~new_A9905_;
  assign new_A9901_ = new_A9869_ | new_A9906_;
  assign new_A9900_ = new_A9852_ & ~new_A9853_;
  assign new_A9899_ = ~new_A9852_ & new_A9853_;
  assign new_A9898_ = new_A9862_ | new_A9895_;
  assign new_A9897_ = ~new_A9862_ & ~new_A9896_;
  assign new_A9896_ = new_A9862_ & new_A9895_;
  assign new_A9895_ = ~new_A9851_ | ~new_A9876_;
  assign new_A9894_ = ~new_A9852_ & new_A9862_;
  assign new_A9893_ = new_A9852_ & ~new_A9862_;
  assign new_A9892_ = new_A9854_ & new_A9891_;
  assign new_A9891_ = new_A9910_ | new_A9909_;
  assign new_A9890_ = ~new_A9854_ & new_A9889_;
  assign new_A9889_ = new_A9912_ | new_A9911_;
  assign new_A9888_ = new_A9854_ | new_A9887_;
  assign new_A9887_ = new_A9908_ | new_A9907_;
  assign new_A9886_ = ~new_A9866_ & ~new_A9876_;
  assign new_A9885_ = new_A9866_ & new_A9876_;
  assign new_A9884_ = ~new_A9866_ | new_A9876_;
  assign new_A9883_ = new_A9850_ & ~new_A9851_;
  assign new_A9882_ = ~new_A9850_ & new_A9851_;
  assign new_A9881_ = new_A9903_ & ~new_A9904_;
  assign new_A9880_ = ~new_A9903_ & new_A9904_;
  assign new_A9879_ = ~new_A9902_ | ~new_A9901_;
  assign new_A9878_ = new_A9894_ | new_A9893_;
  assign new_A9877_ = new_A9900_ | new_A9899_;
  assign new_A9876_ = new_A9890_ | new_A9892_;
  assign new_A9875_ = ~new_A9897_ | ~new_A9898_;
  assign new_A9874_ = new_A9850_ & ~new_A9851_;
  assign new_A9873_ = new_A9864_ & ~new_A9876_;
  assign new_A9872_ = ~new_A9864_ & new_A9876_;
  assign new_A9871_ = ~new_A9862_ & new_A9888_;
  assign new_A9870_ = new_A9886_ | new_A9885_;
  assign new_A9869_ = new_A9883_ | new_A9882_;
  assign new_A9868_ = new_A9851_ | new_A9884_;
  assign new_A9867_ = new_A9876_ & new_A9879_;
  assign new_A9866_ = new_A9881_ | new_A9880_;
  assign new_A9865_ = new_A9876_ & new_A9875_;
  assign new_A9864_ = new_A9878_ & new_A9877_;
  assign new_A9863_ = new_A9873_ | new_A9872_;
  assign new_A9862_ = new_A9851_ | new_A9874_;
  assign A9861 = new_A9862_ | new_A9871_;
  assign A9860 = new_A9869_ & new_A9870_;
  assign A9859 = new_A9869_ & new_A9868_;
  assign A9858 = new_A9867_ | new_A9866_;
  assign A9857 = new_A9865_ | new_A9864_;
  assign A9856 = new_A9863_ & new_A9862_;
  assign new_A9855_ = new_D3711_;
  assign new_A9854_ = new_D3644_;
  assign new_A9853_ = new_D3577_;
  assign new_A9852_ = new_D3510_;
  assign new_A9851_ = new_D3443_;
  assign new_A9850_ = new_D3376_;
  assign new_A9849_ = ~new_A9788_ & new_A9802_;
  assign new_A9848_ = new_A9788_ & ~new_A9802_;
  assign new_A9847_ = new_A9788_ & ~new_A9802_;
  assign new_A9846_ = ~new_A9788_ & ~new_A9802_;
  assign new_A9845_ = new_A9788_ & new_A9802_;
  assign new_A9844_ = new_A9848_ | new_A9849_;
  assign new_A9843_ = ~new_A9788_ & new_A9802_;
  assign new_A9842_ = new_A9846_ | new_A9847_;
  assign new_A9841_ = ~new_A9817_ & ~new_A9837_;
  assign new_A9840_ = new_A9817_ & new_A9837_;
  assign new_A9839_ = ~new_A9784_ | ~new_A9809_;
  assign new_A9838_ = new_A9802_ & new_A9839_;
  assign new_A9837_ = new_A9785_ | new_A9786_;
  assign new_A9836_ = new_A9785_ | new_A9802_;
  assign new_A9835_ = ~new_A9802_ & ~new_A9838_;
  assign new_A9834_ = new_A9802_ | new_A9839_;
  assign new_A9833_ = new_A9785_ & ~new_A9786_;
  assign new_A9832_ = ~new_A9785_ & new_A9786_;
  assign new_A9831_ = new_A9795_ | new_A9828_;
  assign new_A9830_ = ~new_A9795_ & ~new_A9829_;
  assign new_A9829_ = new_A9795_ & new_A9828_;
  assign new_A9828_ = ~new_A9784_ | ~new_A9809_;
  assign new_A9827_ = ~new_A9785_ & new_A9795_;
  assign new_A9826_ = new_A9785_ & ~new_A9795_;
  assign new_A9825_ = new_A9787_ & new_A9824_;
  assign new_A9824_ = new_A9843_ | new_A9842_;
  assign new_A9823_ = ~new_A9787_ & new_A9822_;
  assign new_A9822_ = new_A9845_ | new_A9844_;
  assign new_A9821_ = new_A9787_ | new_A9820_;
  assign new_A9820_ = new_A9841_ | new_A9840_;
  assign new_A9819_ = ~new_A9799_ & ~new_A9809_;
  assign new_A9818_ = new_A9799_ & new_A9809_;
  assign new_A9817_ = ~new_A9799_ | new_A9809_;
  assign new_A9816_ = new_A9783_ & ~new_A9784_;
  assign new_A9815_ = ~new_A9783_ & new_A9784_;
  assign new_A9814_ = new_A9836_ & ~new_A9837_;
  assign new_A9813_ = ~new_A9836_ & new_A9837_;
  assign new_A9812_ = ~new_A9835_ | ~new_A9834_;
  assign new_A9811_ = new_A9827_ | new_A9826_;
  assign new_A9810_ = new_A9833_ | new_A9832_;
  assign new_A9809_ = new_A9823_ | new_A9825_;
  assign new_A9808_ = ~new_A9830_ | ~new_A9831_;
  assign new_A9807_ = new_A9783_ & ~new_A9784_;
  assign new_A9806_ = new_A9797_ & ~new_A9809_;
  assign new_A9805_ = ~new_A9797_ & new_A9809_;
  assign new_A9804_ = ~new_A9795_ & new_A9821_;
  assign new_A9803_ = new_A9819_ | new_A9818_;
  assign new_A9802_ = new_A9816_ | new_A9815_;
  assign new_A9801_ = new_A9784_ | new_A9817_;
  assign new_A9800_ = new_A9809_ & new_A9812_;
  assign new_A9799_ = new_A9814_ | new_A9813_;
  assign new_A9798_ = new_A9809_ & new_A9808_;
  assign new_A9797_ = new_A9811_ & new_A9810_;
  assign new_A9796_ = new_A9806_ | new_A9805_;
  assign new_A9795_ = new_A9784_ | new_A9807_;
  assign A9794 = new_A9795_ | new_A9804_;
  assign A9793 = new_A9802_ & new_A9803_;
  assign A9792 = new_A9802_ & new_A9801_;
  assign A9791 = new_A9800_ | new_A9799_;
  assign A9790 = new_A9798_ | new_A9797_;
  assign A9789 = new_A9796_ & new_A9795_;
  assign new_A9788_ = new_D3309_;
  assign new_A9787_ = new_D3242_;
  assign new_A9786_ = new_D3175_;
  assign new_A9785_ = new_D3108_;
  assign new_A9784_ = new_D3041_;
  assign new_A9783_ = new_D2974_;
  assign new_A9782_ = ~new_A9721_ & new_A9735_;
  assign new_A9781_ = new_A9721_ & ~new_A9735_;
  assign new_A9780_ = new_A9721_ & ~new_A9735_;
  assign new_A9779_ = ~new_A9721_ & ~new_A9735_;
  assign new_A9778_ = new_A9721_ & new_A9735_;
  assign new_A9777_ = new_A9781_ | new_A9782_;
  assign new_A9776_ = ~new_A9721_ & new_A9735_;
  assign new_A9775_ = new_A9779_ | new_A9780_;
  assign new_A9774_ = ~new_A9750_ & ~new_A9770_;
  assign new_A9773_ = new_A9750_ & new_A9770_;
  assign new_A9772_ = ~new_A9717_ | ~new_A9742_;
  assign new_A9771_ = new_A9735_ & new_A9772_;
  assign new_A9770_ = new_A9718_ | new_A9719_;
  assign new_A9769_ = new_A9718_ | new_A9735_;
  assign new_A9768_ = ~new_A9735_ & ~new_A9771_;
  assign new_A9767_ = new_A9735_ | new_A9772_;
  assign new_A9766_ = new_A9718_ & ~new_A9719_;
  assign new_A9765_ = ~new_A9718_ & new_A9719_;
  assign new_A9764_ = new_A9728_ | new_A9761_;
  assign new_A9763_ = ~new_A9728_ & ~new_A9762_;
  assign new_A9762_ = new_A9728_ & new_A9761_;
  assign new_A9761_ = ~new_A9717_ | ~new_A9742_;
  assign new_A9760_ = ~new_A9718_ & new_A9728_;
  assign new_A9759_ = new_A9718_ & ~new_A9728_;
  assign new_A9758_ = new_A9720_ & new_A9757_;
  assign new_A9757_ = new_A9776_ | new_A9775_;
  assign new_A9756_ = ~new_A9720_ & new_A9755_;
  assign new_A9755_ = new_A9778_ | new_A9777_;
  assign new_A9754_ = new_A9720_ | new_A9753_;
  assign new_A9753_ = new_A9774_ | new_A9773_;
  assign new_A9752_ = ~new_A9732_ & ~new_A9742_;
  assign new_A9751_ = new_A9732_ & new_A9742_;
  assign new_A9750_ = ~new_A9732_ | new_A9742_;
  assign new_A9749_ = new_A9716_ & ~new_A9717_;
  assign new_A9748_ = ~new_A9716_ & new_A9717_;
  assign new_A9747_ = new_A9769_ & ~new_A9770_;
  assign new_A9746_ = ~new_A9769_ & new_A9770_;
  assign new_A9745_ = ~new_A9768_ | ~new_A9767_;
  assign new_A9744_ = new_A9760_ | new_A9759_;
  assign new_A9743_ = new_A9766_ | new_A9765_;
  assign new_A9742_ = new_A9756_ | new_A9758_;
  assign new_A9741_ = ~new_A9763_ | ~new_A9764_;
  assign new_A9740_ = new_A9716_ & ~new_A9717_;
  assign new_A9739_ = new_A9730_ & ~new_A9742_;
  assign new_A9738_ = ~new_A9730_ & new_A9742_;
  assign new_A9737_ = ~new_A9728_ & new_A9754_;
  assign new_A9736_ = new_A9752_ | new_A9751_;
  assign new_A9735_ = new_A9749_ | new_A9748_;
  assign new_A9734_ = new_A9717_ | new_A9750_;
  assign new_A9733_ = new_A9742_ & new_A9745_;
  assign new_A9732_ = new_A9747_ | new_A9746_;
  assign new_A9731_ = new_A9742_ & new_A9741_;
  assign new_A9730_ = new_A9744_ & new_A9743_;
  assign new_A9729_ = new_A9739_ | new_A9738_;
  assign new_A9728_ = new_A9717_ | new_A9740_;
  assign A9727 = new_A9728_ | new_A9737_;
  assign A9726 = new_A9735_ & new_A9736_;
  assign A9725 = new_A9735_ & new_A9734_;
  assign A9724 = new_A9733_ | new_A9732_;
  assign A9723 = new_A9731_ | new_A9730_;
  assign A9722 = new_A9729_ & new_A9728_;
  assign new_A9721_ = new_D2907_;
  assign new_A9720_ = new_D2840_;
  assign new_A9719_ = new_D2773_;
  assign new_A9718_ = new_D2706_;
  assign new_A9717_ = new_D2639_;
  assign new_A9716_ = new_D2572_;
  assign new_A9715_ = ~new_A9654_ & new_A9668_;
  assign new_A9714_ = new_A9654_ & ~new_A9668_;
  assign new_A9713_ = new_A9654_ & ~new_A9668_;
  assign new_A9712_ = ~new_A9654_ & ~new_A9668_;
  assign new_A9711_ = new_A9654_ & new_A9668_;
  assign new_A9710_ = new_A9714_ | new_A9715_;
  assign new_A9709_ = ~new_A9654_ & new_A9668_;
  assign new_A9708_ = new_A9712_ | new_A9713_;
  assign new_A9707_ = ~new_A9683_ & ~new_A9703_;
  assign new_A9706_ = new_A9683_ & new_A9703_;
  assign new_A9705_ = ~new_A9650_ | ~new_A9675_;
  assign new_A9704_ = new_A9668_ & new_A9705_;
  assign new_A9703_ = new_A9651_ | new_A9652_;
  assign new_A9702_ = new_A9651_ | new_A9668_;
  assign new_A9701_ = ~new_A9668_ & ~new_A9704_;
  assign new_A9700_ = new_A9668_ | new_A9705_;
  assign new_A9699_ = new_A9651_ & ~new_A9652_;
  assign new_A9698_ = ~new_A9651_ & new_A9652_;
  assign new_A9697_ = new_A9661_ | new_A9694_;
  assign new_A9696_ = ~new_A9661_ & ~new_A9695_;
  assign new_A9695_ = new_A9661_ & new_A9694_;
  assign new_A9694_ = ~new_A9650_ | ~new_A9675_;
  assign new_A9693_ = ~new_A9651_ & new_A9661_;
  assign new_A9692_ = new_A9651_ & ~new_A9661_;
  assign new_A9691_ = new_A9653_ & new_A9690_;
  assign new_A9690_ = new_A9709_ | new_A9708_;
  assign new_A9689_ = ~new_A9653_ & new_A9688_;
  assign new_A9688_ = new_A9711_ | new_A9710_;
  assign new_A9687_ = new_A9653_ | new_A9686_;
  assign new_A9686_ = new_A9707_ | new_A9706_;
  assign new_A9685_ = ~new_A9665_ & ~new_A9675_;
  assign new_A9684_ = new_A9665_ & new_A9675_;
  assign new_A9683_ = ~new_A9665_ | new_A9675_;
  assign new_A9682_ = new_A9649_ & ~new_A9650_;
  assign new_A9681_ = ~new_A9649_ & new_A9650_;
  assign new_A9680_ = new_A9702_ & ~new_A9703_;
  assign new_A9679_ = ~new_A9702_ & new_A9703_;
  assign new_A9678_ = ~new_A9701_ | ~new_A9700_;
  assign new_A9677_ = new_A9693_ | new_A9692_;
  assign new_A9676_ = new_A9699_ | new_A9698_;
  assign new_A9675_ = new_A9689_ | new_A9691_;
  assign new_A9674_ = ~new_A9696_ | ~new_A9697_;
  assign new_A9673_ = new_A9649_ & ~new_A9650_;
  assign new_A9672_ = new_A9663_ & ~new_A9675_;
  assign new_A9671_ = ~new_A9663_ & new_A9675_;
  assign new_A9670_ = ~new_A9661_ & new_A9687_;
  assign new_A9669_ = new_A9685_ | new_A9684_;
  assign new_A9668_ = new_A9682_ | new_A9681_;
  assign new_A9667_ = new_A9650_ | new_A9683_;
  assign new_A9666_ = new_A9675_ & new_A9678_;
  assign new_A9665_ = new_A9680_ | new_A9679_;
  assign new_A9664_ = new_A9675_ & new_A9674_;
  assign new_A9663_ = new_A9677_ & new_A9676_;
  assign new_A9662_ = new_A9672_ | new_A9671_;
  assign new_A9661_ = new_A9650_ | new_A9673_;
  assign A9660 = new_A9661_ | new_A9670_;
  assign A9659 = new_A9668_ & new_A9669_;
  assign A9658 = new_A9668_ & new_A9667_;
  assign A9657 = new_A9666_ | new_A9665_;
  assign A9656 = new_A9664_ | new_A9663_;
  assign A9655 = new_A9662_ & new_A9661_;
  assign new_A9654_ = new_D2505_;
  assign new_A9653_ = new_D2438_;
  assign new_A9652_ = new_D2371_;
  assign new_A9651_ = new_D2304_;
  assign new_A9650_ = new_D2237_;
  assign new_A9649_ = new_D2170_;
  assign new_A9648_ = ~new_A9587_ & new_A9601_;
  assign new_A9647_ = new_A9587_ & ~new_A9601_;
  assign new_A9646_ = new_A9587_ & ~new_A9601_;
  assign new_A9645_ = ~new_A9587_ & ~new_A9601_;
  assign new_A9644_ = new_A9587_ & new_A9601_;
  assign new_A9643_ = new_A9647_ | new_A9648_;
  assign new_A9642_ = ~new_A9587_ & new_A9601_;
  assign new_A9641_ = new_A9645_ | new_A9646_;
  assign new_A9640_ = ~new_A9616_ & ~new_A9636_;
  assign new_A9639_ = new_A9616_ & new_A9636_;
  assign new_A9638_ = ~new_A9583_ | ~new_A9608_;
  assign new_A9637_ = new_A9601_ & new_A9638_;
  assign new_A9636_ = new_A9584_ | new_A9585_;
  assign new_A9635_ = new_A9584_ | new_A9601_;
  assign new_A9634_ = ~new_A9601_ & ~new_A9637_;
  assign new_A9633_ = new_A9601_ | new_A9638_;
  assign new_A9632_ = new_A9584_ & ~new_A9585_;
  assign new_A9631_ = ~new_A9584_ & new_A9585_;
  assign new_A9630_ = new_A9594_ | new_A9627_;
  assign new_A9629_ = ~new_A9594_ & ~new_A9628_;
  assign new_A9628_ = new_A9594_ & new_A9627_;
  assign new_A9627_ = ~new_A9583_ | ~new_A9608_;
  assign new_A9626_ = ~new_A9584_ & new_A9594_;
  assign new_A9625_ = new_A9584_ & ~new_A9594_;
  assign new_A9624_ = new_A9586_ & new_A9623_;
  assign new_A9623_ = new_A9642_ | new_A9641_;
  assign new_A9622_ = ~new_A9586_ & new_A9621_;
  assign new_A9621_ = new_A9644_ | new_A9643_;
  assign new_A9620_ = new_A9586_ | new_A9619_;
  assign new_A9619_ = new_A9640_ | new_A9639_;
  assign new_A9618_ = ~new_A9598_ & ~new_A9608_;
  assign new_A9617_ = new_A9598_ & new_A9608_;
  assign new_A9616_ = ~new_A9598_ | new_A9608_;
  assign new_A9615_ = new_A9582_ & ~new_A9583_;
  assign new_A9614_ = ~new_A9582_ & new_A9583_;
  assign new_A9613_ = new_A9635_ & ~new_A9636_;
  assign new_A9612_ = ~new_A9635_ & new_A9636_;
  assign new_A9611_ = ~new_A9634_ | ~new_A9633_;
  assign new_A9610_ = new_A9626_ | new_A9625_;
  assign new_A9609_ = new_A9632_ | new_A9631_;
  assign new_A9608_ = new_A9622_ | new_A9624_;
  assign new_A9607_ = ~new_A9629_ | ~new_A9630_;
  assign new_A9606_ = new_A9582_ & ~new_A9583_;
  assign new_A9605_ = new_A9596_ & ~new_A9608_;
  assign new_A9604_ = ~new_A9596_ & new_A9608_;
  assign new_A9603_ = ~new_A9594_ & new_A9620_;
  assign new_A9602_ = new_A9618_ | new_A9617_;
  assign new_A9601_ = new_A9615_ | new_A9614_;
  assign new_A9600_ = new_A9583_ | new_A9616_;
  assign new_A9599_ = new_A9608_ & new_A9611_;
  assign new_A9598_ = new_A9613_ | new_A9612_;
  assign new_A9597_ = new_A9608_ & new_A9607_;
  assign new_A9596_ = new_A9610_ & new_A9609_;
  assign new_A9595_ = new_A9605_ | new_A9604_;
  assign new_A9594_ = new_A9583_ | new_A9606_;
  assign A9593 = new_A9594_ | new_A9603_;
  assign A9592 = new_A9601_ & new_A9602_;
  assign A9591 = new_A9601_ & new_A9600_;
  assign A9590 = new_A9599_ | new_A9598_;
  assign A9589 = new_A9597_ | new_A9596_;
  assign A9588 = new_A9595_ & new_A9594_;
  assign new_A9587_ = new_D2103_;
  assign new_A9586_ = new_D2036_;
  assign new_A9585_ = new_D1969_;
  assign new_A9584_ = new_D1902_;
  assign new_A9583_ = new_D1835_;
  assign new_A9582_ = new_D1768_;
  assign new_A9581_ = ~new_A9520_ & new_A9534_;
  assign new_A9580_ = new_A9520_ & ~new_A9534_;
  assign new_A9579_ = new_A9520_ & ~new_A9534_;
  assign new_A9578_ = ~new_A9520_ & ~new_A9534_;
  assign new_A9577_ = new_A9520_ & new_A9534_;
  assign new_A9576_ = new_A9580_ | new_A9581_;
  assign new_A9575_ = ~new_A9520_ & new_A9534_;
  assign new_A9574_ = new_A9578_ | new_A9579_;
  assign new_A9573_ = ~new_A9549_ & ~new_A9569_;
  assign new_A9572_ = new_A9549_ & new_A9569_;
  assign new_A9571_ = ~new_A9516_ | ~new_A9541_;
  assign new_A9570_ = new_A9534_ & new_A9571_;
  assign new_A9569_ = new_A9517_ | new_A9518_;
  assign new_A9568_ = new_A9517_ | new_A9534_;
  assign new_A9567_ = ~new_A9534_ & ~new_A9570_;
  assign new_A9566_ = new_A9534_ | new_A9571_;
  assign new_A9565_ = new_A9517_ & ~new_A9518_;
  assign new_A9564_ = ~new_A9517_ & new_A9518_;
  assign new_A9563_ = new_A9527_ | new_A9560_;
  assign new_A9562_ = ~new_A9527_ & ~new_A9561_;
  assign new_A9561_ = new_A9527_ & new_A9560_;
  assign new_A9560_ = ~new_A9516_ | ~new_A9541_;
  assign new_A9559_ = ~new_A9517_ & new_A9527_;
  assign new_A9558_ = new_A9517_ & ~new_A9527_;
  assign new_A9557_ = new_A9519_ & new_A9556_;
  assign new_A9556_ = new_A9575_ | new_A9574_;
  assign new_A9555_ = ~new_A9519_ & new_A9554_;
  assign new_A9554_ = new_A9577_ | new_A9576_;
  assign new_A9553_ = new_A9519_ | new_A9552_;
  assign new_A9552_ = new_A9573_ | new_A9572_;
  assign new_A9551_ = ~new_A9531_ & ~new_A9541_;
  assign new_A9550_ = new_A9531_ & new_A9541_;
  assign new_A9549_ = ~new_A9531_ | new_A9541_;
  assign new_A9548_ = new_A9515_ & ~new_A9516_;
  assign new_A9547_ = ~new_A9515_ & new_A9516_;
  assign new_A9546_ = new_A9568_ & ~new_A9569_;
  assign new_A9545_ = ~new_A9568_ & new_A9569_;
  assign new_A9544_ = ~new_A9567_ | ~new_A9566_;
  assign new_A9543_ = new_A9559_ | new_A9558_;
  assign new_A9542_ = new_A9565_ | new_A9564_;
  assign new_A9541_ = new_A9555_ | new_A9557_;
  assign new_A9540_ = ~new_A9562_ | ~new_A9563_;
  assign new_A9539_ = new_A9515_ & ~new_A9516_;
  assign new_A9538_ = new_A9529_ & ~new_A9541_;
  assign new_A9537_ = ~new_A9529_ & new_A9541_;
  assign new_A9536_ = ~new_A9527_ & new_A9553_;
  assign new_A9535_ = new_A9551_ | new_A9550_;
  assign new_A9534_ = new_A9548_ | new_A9547_;
  assign new_A9533_ = new_A9516_ | new_A9549_;
  assign new_A9532_ = new_A9541_ & new_A9544_;
  assign new_A9531_ = new_A9546_ | new_A9545_;
  assign new_A9530_ = new_A9541_ & new_A9540_;
  assign new_A9529_ = new_A9543_ & new_A9542_;
  assign new_A9528_ = new_A9538_ | new_A9537_;
  assign new_A9527_ = new_A9516_ | new_A9539_;
  assign A9526 = new_A9527_ | new_A9536_;
  assign A9525 = new_A9534_ & new_A9535_;
  assign A9524 = new_A9534_ & new_A9533_;
  assign A9523 = new_A9532_ | new_A9531_;
  assign A9522 = new_A9530_ | new_A9529_;
  assign A9521 = new_A9528_ & new_A9527_;
  assign new_A9520_ = new_D1701_;
  assign new_A9519_ = new_D1634_;
  assign new_A9518_ = new_D1567_;
  assign new_A9517_ = new_D1500_;
  assign new_A9516_ = new_D1433_;
  assign new_A9515_ = new_D1366_;
  assign new_A9514_ = ~new_A9453_ & new_A9467_;
  assign new_A9513_ = new_A9453_ & ~new_A9467_;
  assign new_A9512_ = new_A9453_ & ~new_A9467_;
  assign new_A9511_ = ~new_A9453_ & ~new_A9467_;
  assign new_A9510_ = new_A9453_ & new_A9467_;
  assign new_A9509_ = new_A9513_ | new_A9514_;
  assign new_A9508_ = ~new_A9453_ & new_A9467_;
  assign new_A9507_ = new_A9511_ | new_A9512_;
  assign new_A9506_ = ~new_A9482_ & ~new_A9502_;
  assign new_A9505_ = new_A9482_ & new_A9502_;
  assign new_A9504_ = ~new_A9449_ | ~new_A9474_;
  assign new_A9503_ = new_A9467_ & new_A9504_;
  assign new_A9502_ = new_A9450_ | new_A9451_;
  assign new_A9501_ = new_A9450_ | new_A9467_;
  assign new_A9500_ = ~new_A9467_ & ~new_A9503_;
  assign new_A9499_ = new_A9467_ | new_A9504_;
  assign new_A9498_ = new_A9450_ & ~new_A9451_;
  assign new_A9497_ = ~new_A9450_ & new_A9451_;
  assign new_A9496_ = new_A9460_ | new_A9493_;
  assign new_A9495_ = ~new_A9460_ & ~new_A9494_;
  assign new_A9494_ = new_A9460_ & new_A9493_;
  assign new_A9493_ = ~new_A9449_ | ~new_A9474_;
  assign new_A9492_ = ~new_A9450_ & new_A9460_;
  assign new_A9491_ = new_A9450_ & ~new_A9460_;
  assign new_A9490_ = new_A9452_ & new_A9489_;
  assign new_A9489_ = new_A9508_ | new_A9507_;
  assign new_A9488_ = ~new_A9452_ & new_A9487_;
  assign new_A9487_ = new_A9510_ | new_A9509_;
  assign new_A9486_ = new_A9452_ | new_A9485_;
  assign new_A9485_ = new_A9506_ | new_A9505_;
  assign new_A9484_ = ~new_A9464_ & ~new_A9474_;
  assign new_A9483_ = new_A9464_ & new_A9474_;
  assign new_A9482_ = ~new_A9464_ | new_A9474_;
  assign new_A9481_ = new_A9448_ & ~new_A9449_;
  assign new_A9480_ = ~new_A9448_ & new_A9449_;
  assign new_A9479_ = new_A9501_ & ~new_A9502_;
  assign new_A9478_ = ~new_A9501_ & new_A9502_;
  assign new_A9477_ = ~new_A9500_ | ~new_A9499_;
  assign new_A9476_ = new_A9492_ | new_A9491_;
  assign new_A9475_ = new_A9498_ | new_A9497_;
  assign new_A9474_ = new_A9488_ | new_A9490_;
  assign new_A9473_ = ~new_A9495_ | ~new_A9496_;
  assign new_A9472_ = new_A9448_ & ~new_A9449_;
  assign new_A9471_ = new_A9462_ & ~new_A9474_;
  assign new_A9470_ = ~new_A9462_ & new_A9474_;
  assign new_A9469_ = ~new_A9460_ & new_A9486_;
  assign new_A9468_ = new_A9484_ | new_A9483_;
  assign new_A9467_ = new_A9481_ | new_A9480_;
  assign new_A9466_ = new_A9449_ | new_A9482_;
  assign new_A9465_ = new_A9474_ & new_A9477_;
  assign new_A9464_ = new_A9479_ | new_A9478_;
  assign new_A9463_ = new_A9474_ & new_A9473_;
  assign new_A9462_ = new_A9476_ & new_A9475_;
  assign new_A9461_ = new_A9471_ | new_A9470_;
  assign new_A9460_ = new_A9449_ | new_A9472_;
  assign A9459 = new_A9460_ | new_A9469_;
  assign A9458 = new_A9467_ & new_A9468_;
  assign A9457 = new_A9467_ & new_A9466_;
  assign A9456 = new_A9465_ | new_A9464_;
  assign A9455 = new_A9463_ | new_A9462_;
  assign A9454 = new_A9461_ & new_A9460_;
  assign new_A9453_ = new_D1299_;
  assign new_A9452_ = new_D1232_;
  assign new_A9451_ = new_D1165_;
  assign new_A9450_ = new_D1098_;
  assign new_A9449_ = new_D1031_;
  assign new_A9448_ = new_D964_;
  assign new_A9447_ = ~new_A9386_ & new_A9400_;
  assign new_A9446_ = new_A9386_ & ~new_A9400_;
  assign new_A9445_ = new_A9386_ & ~new_A9400_;
  assign new_A9444_ = ~new_A9386_ & ~new_A9400_;
  assign new_A9443_ = new_A9386_ & new_A9400_;
  assign new_A9442_ = new_A9446_ | new_A9447_;
  assign new_A9441_ = ~new_A9386_ & new_A9400_;
  assign new_A9440_ = new_A9444_ | new_A9445_;
  assign new_A9439_ = ~new_A9415_ & ~new_A9435_;
  assign new_A9438_ = new_A9415_ & new_A9435_;
  assign new_A9437_ = ~new_A9382_ | ~new_A9407_;
  assign new_A9436_ = new_A9400_ & new_A9437_;
  assign new_A9435_ = new_A9383_ | new_A9384_;
  assign new_A9434_ = new_A9383_ | new_A9400_;
  assign new_A9433_ = ~new_A9400_ & ~new_A9436_;
  assign new_A9432_ = new_A9400_ | new_A9437_;
  assign new_A9431_ = new_A9383_ & ~new_A9384_;
  assign new_A9430_ = ~new_A9383_ & new_A9384_;
  assign new_A9429_ = new_A9393_ | new_A9426_;
  assign new_A9428_ = ~new_A9393_ & ~new_A9427_;
  assign new_A9427_ = new_A9393_ & new_A9426_;
  assign new_A9426_ = ~new_A9382_ | ~new_A9407_;
  assign new_A9425_ = ~new_A9383_ & new_A9393_;
  assign new_A9424_ = new_A9383_ & ~new_A9393_;
  assign new_A9423_ = new_A9385_ & new_A9422_;
  assign new_A9422_ = new_A9441_ | new_A9440_;
  assign new_A9421_ = ~new_A9385_ & new_A9420_;
  assign new_A9420_ = new_A9443_ | new_A9442_;
  assign new_A9419_ = new_A9385_ | new_A9418_;
  assign new_A9418_ = new_A9439_ | new_A9438_;
  assign new_A9417_ = ~new_A9397_ & ~new_A9407_;
  assign new_A9416_ = new_A9397_ & new_A9407_;
  assign new_A9415_ = ~new_A9397_ | new_A9407_;
  assign new_A9414_ = new_A9381_ & ~new_A9382_;
  assign new_A9413_ = ~new_A9381_ & new_A9382_;
  assign new_A9412_ = new_A9434_ & ~new_A9435_;
  assign new_A9411_ = ~new_A9434_ & new_A9435_;
  assign new_A9410_ = ~new_A9433_ | ~new_A9432_;
  assign new_A9409_ = new_A9425_ | new_A9424_;
  assign new_A9408_ = new_A9431_ | new_A9430_;
  assign new_A9407_ = new_A9421_ | new_A9423_;
  assign new_A9406_ = ~new_A9428_ | ~new_A9429_;
  assign new_A9405_ = new_A9381_ & ~new_A9382_;
  assign new_A9404_ = new_A9395_ & ~new_A9407_;
  assign new_A9403_ = ~new_A9395_ & new_A9407_;
  assign new_A9402_ = ~new_A9393_ & new_A9419_;
  assign new_A9401_ = new_A9417_ | new_A9416_;
  assign new_A9400_ = new_A9414_ | new_A9413_;
  assign new_A9399_ = new_A9382_ | new_A9415_;
  assign new_A9398_ = new_A9407_ & new_A9410_;
  assign new_A9397_ = new_A9412_ | new_A9411_;
  assign new_A9396_ = new_A9407_ & new_A9406_;
  assign new_A9395_ = new_A9409_ & new_A9408_;
  assign new_A9394_ = new_A9404_ | new_A9403_;
  assign new_A9393_ = new_A9382_ | new_A9405_;
  assign A9392 = new_A9393_ | new_A9402_;
  assign A9391 = new_A9400_ & new_A9401_;
  assign A9390 = new_A9400_ & new_A9399_;
  assign A9389 = new_A9398_ | new_A9397_;
  assign A9388 = new_A9396_ | new_A9395_;
  assign A9387 = new_A9394_ & new_A9393_;
  assign new_A9386_ = new_D897_;
  assign new_A9385_ = new_D830_;
  assign new_A9384_ = new_D763_;
  assign new_A9383_ = new_D696_;
  assign new_A9382_ = new_D629_;
  assign new_A9381_ = new_D562_;
  assign new_A9380_ = ~new_A9319_ & new_A9333_;
  assign new_A9379_ = new_A9319_ & ~new_A9333_;
  assign new_A9378_ = new_A9319_ & ~new_A9333_;
  assign new_A9377_ = ~new_A9319_ & ~new_A9333_;
  assign new_A9376_ = new_A9319_ & new_A9333_;
  assign new_A9375_ = new_A9379_ | new_A9380_;
  assign new_A9374_ = ~new_A9319_ & new_A9333_;
  assign new_A9373_ = new_A9377_ | new_A9378_;
  assign new_A9372_ = ~new_A9348_ & ~new_A9368_;
  assign new_A9371_ = new_A9348_ & new_A9368_;
  assign new_A9370_ = ~new_A9315_ | ~new_A9340_;
  assign new_A9369_ = new_A9333_ & new_A9370_;
  assign new_A9368_ = new_A9316_ | new_A9317_;
  assign new_A9367_ = new_A9316_ | new_A9333_;
  assign new_A9366_ = ~new_A9333_ & ~new_A9369_;
  assign new_A9365_ = new_A9333_ | new_A9370_;
  assign new_A9364_ = new_A9316_ & ~new_A9317_;
  assign new_A9363_ = ~new_A9316_ & new_A9317_;
  assign new_A9362_ = new_A9326_ | new_A9359_;
  assign new_A9361_ = ~new_A9326_ & ~new_A9360_;
  assign new_A9360_ = new_A9326_ & new_A9359_;
  assign new_A9359_ = ~new_A9315_ | ~new_A9340_;
  assign new_A9358_ = ~new_A9316_ & new_A9326_;
  assign new_A9357_ = new_A9316_ & ~new_A9326_;
  assign new_A9356_ = new_A9318_ & new_A9355_;
  assign new_A9355_ = new_A9374_ | new_A9373_;
  assign new_A9354_ = ~new_A9318_ & new_A9353_;
  assign new_A9353_ = new_A9376_ | new_A9375_;
  assign new_A9352_ = new_A9318_ | new_A9351_;
  assign new_A9351_ = new_A9372_ | new_A9371_;
  assign new_A9350_ = ~new_A9330_ & ~new_A9340_;
  assign new_A9349_ = new_A9330_ & new_A9340_;
  assign new_A9348_ = ~new_A9330_ | new_A9340_;
  assign new_A9347_ = new_A9314_ & ~new_A9315_;
  assign new_A9346_ = ~new_A9314_ & new_A9315_;
  assign new_A9345_ = new_A9367_ & ~new_A9368_;
  assign new_A9344_ = ~new_A9367_ & new_A9368_;
  assign new_A9343_ = ~new_A9366_ | ~new_A9365_;
  assign new_A9342_ = new_A9358_ | new_A9357_;
  assign new_A9341_ = new_A9364_ | new_A9363_;
  assign new_A9340_ = new_A9354_ | new_A9356_;
  assign new_A9339_ = ~new_A9361_ | ~new_A9362_;
  assign new_A9338_ = new_A9314_ & ~new_A9315_;
  assign new_A9337_ = new_A9328_ & ~new_A9340_;
  assign new_A9336_ = ~new_A9328_ & new_A9340_;
  assign new_A9335_ = ~new_A9326_ & new_A9352_;
  assign new_A9334_ = new_A9350_ | new_A9349_;
  assign new_A9333_ = new_A9347_ | new_A9346_;
  assign new_A9332_ = new_A9315_ | new_A9348_;
  assign new_A9331_ = new_A9340_ & new_A9343_;
  assign new_A9330_ = new_A9345_ | new_A9344_;
  assign new_A9329_ = new_A9340_ & new_A9339_;
  assign new_A9328_ = new_A9342_ & new_A9341_;
  assign new_A9327_ = new_A9337_ | new_A9336_;
  assign new_A9326_ = new_A9315_ | new_A9338_;
  assign A9325 = new_A9326_ | new_A9335_;
  assign A9324 = new_A9333_ & new_A9334_;
  assign A9323 = new_A9333_ & new_A9332_;
  assign A9322 = new_A9331_ | new_A9330_;
  assign A9321 = new_A9329_ | new_A9328_;
  assign A9320 = new_A9327_ & new_A9326_;
  assign new_A9319_ = new_D495_;
  assign new_A9318_ = new_D428_;
  assign new_A9317_ = new_D361_;
  assign new_A9316_ = new_D294_;
  assign new_A9315_ = new_D227_;
  assign new_A9314_ = new_D160_;
  assign new_A9313_ = ~new_A9252_ & new_A9266_;
  assign new_A9312_ = new_A9252_ & ~new_A9266_;
  assign new_A9311_ = new_A9252_ & ~new_A9266_;
  assign new_A9310_ = ~new_A9252_ & ~new_A9266_;
  assign new_A9309_ = new_A9252_ & new_A9266_;
  assign new_A9308_ = new_A9312_ | new_A9313_;
  assign new_A9307_ = ~new_A9252_ & new_A9266_;
  assign new_A9306_ = new_A9310_ | new_A9311_;
  assign new_A9305_ = ~new_A9281_ & ~new_A9301_;
  assign new_A9304_ = new_A9281_ & new_A9301_;
  assign new_A9303_ = ~new_A9248_ | ~new_A9273_;
  assign new_A9302_ = new_A9266_ & new_A9303_;
  assign new_A9301_ = new_A9249_ | new_A9250_;
  assign new_A9300_ = new_A9249_ | new_A9266_;
  assign new_A9299_ = ~new_A9266_ & ~new_A9302_;
  assign new_A9298_ = new_A9266_ | new_A9303_;
  assign new_A9297_ = new_A9249_ & ~new_A9250_;
  assign new_A9296_ = ~new_A9249_ & new_A9250_;
  assign new_A9295_ = new_A9259_ | new_A9292_;
  assign new_A9294_ = ~new_A9259_ & ~new_A9293_;
  assign new_A9293_ = new_A9259_ & new_A9292_;
  assign new_A9292_ = ~new_A9248_ | ~new_A9273_;
  assign new_A9291_ = ~new_A9249_ & new_A9259_;
  assign new_A9290_ = new_A9249_ & ~new_A9259_;
  assign new_A9289_ = new_A9251_ & new_A9288_;
  assign new_A9288_ = new_A9307_ | new_A9306_;
  assign new_A9287_ = ~new_A9251_ & new_A9286_;
  assign new_A9286_ = new_A9309_ | new_A9308_;
  assign new_A9285_ = new_A9251_ | new_A9284_;
  assign new_A9284_ = new_A9305_ | new_A9304_;
  assign new_A9283_ = ~new_A9263_ & ~new_A9273_;
  assign new_A9282_ = new_A9263_ & new_A9273_;
  assign new_A9281_ = ~new_A9263_ | new_A9273_;
  assign new_A9280_ = new_A9247_ & ~new_A9248_;
  assign new_A9279_ = ~new_A9247_ & new_A9248_;
  assign new_A9278_ = new_A9300_ & ~new_A9301_;
  assign new_A9277_ = ~new_A9300_ & new_A9301_;
  assign new_A9276_ = ~new_A9299_ | ~new_A9298_;
  assign new_A9275_ = new_A9291_ | new_A9290_;
  assign new_A9274_ = new_A9297_ | new_A9296_;
  assign new_A9273_ = new_A9287_ | new_A9289_;
  assign new_A9272_ = ~new_A9294_ | ~new_A9295_;
  assign new_A9271_ = new_A9247_ & ~new_A9248_;
  assign new_A9270_ = new_A9261_ & ~new_A9273_;
  assign new_A9269_ = ~new_A9261_ & new_A9273_;
  assign new_A9268_ = ~new_A9259_ & new_A9285_;
  assign new_A9267_ = new_A9283_ | new_A9282_;
  assign new_A9266_ = new_A9280_ | new_A9279_;
  assign new_A9265_ = new_A9248_ | new_A9281_;
  assign new_A9264_ = new_A9273_ & new_A9276_;
  assign new_A9263_ = new_A9278_ | new_A9277_;
  assign new_A9262_ = new_A9273_ & new_A9272_;
  assign new_A9261_ = new_A9275_ & new_A9274_;
  assign new_A9260_ = new_A9270_ | new_A9269_;
  assign new_A9259_ = new_A9248_ | new_A9271_;
  assign A9258 = new_A9259_ | new_A9268_;
  assign A9257 = new_A9266_ & new_A9267_;
  assign A9256 = new_A9266_ & new_A9265_;
  assign A9255 = new_A9264_ | new_A9263_;
  assign A9254 = new_A9262_ | new_A9261_;
  assign A9253 = new_A9260_ & new_A9259_;
  assign new_A9252_ = new_D93_;
  assign new_A9251_ = new_D26_;
  assign new_A9250_ = new_C9958_;
  assign new_A9249_ = new_C9891_;
  assign new_A9248_ = new_C9824_;
  assign new_A9247_ = new_C9757_;
  assign new_A9246_ = ~new_A9185_ & new_A9199_;
  assign new_A9245_ = new_A9185_ & ~new_A9199_;
  assign new_A9244_ = new_A9185_ & ~new_A9199_;
  assign new_A9243_ = ~new_A9185_ & ~new_A9199_;
  assign new_A9242_ = new_A9185_ & new_A9199_;
  assign new_A9241_ = new_A9245_ | new_A9246_;
  assign new_A9240_ = ~new_A9185_ & new_A9199_;
  assign new_A9239_ = new_A9243_ | new_A9244_;
  assign new_A9238_ = ~new_A9214_ & ~new_A9234_;
  assign new_A9237_ = new_A9214_ & new_A9234_;
  assign new_A9236_ = ~new_A9181_ | ~new_A9206_;
  assign new_A9235_ = new_A9199_ & new_A9236_;
  assign new_A9234_ = new_A9182_ | new_A9183_;
  assign new_A9233_ = new_A9182_ | new_A9199_;
  assign new_A9232_ = ~new_A9199_ & ~new_A9235_;
  assign new_A9231_ = new_A9199_ | new_A9236_;
  assign new_A9230_ = new_A9182_ & ~new_A9183_;
  assign new_A9229_ = ~new_A9182_ & new_A9183_;
  assign new_A9228_ = new_A9192_ | new_A9225_;
  assign new_A9227_ = ~new_A9192_ & ~new_A9226_;
  assign new_A9226_ = new_A9192_ & new_A9225_;
  assign new_A9225_ = ~new_A9181_ | ~new_A9206_;
  assign new_A9224_ = ~new_A9182_ & new_A9192_;
  assign new_A9223_ = new_A9182_ & ~new_A9192_;
  assign new_A9222_ = new_A9184_ & new_A9221_;
  assign new_A9221_ = new_A9240_ | new_A9239_;
  assign new_A9220_ = ~new_A9184_ & new_A9219_;
  assign new_A9219_ = new_A9242_ | new_A9241_;
  assign new_A9218_ = new_A9184_ | new_A9217_;
  assign new_A9217_ = new_A9238_ | new_A9237_;
  assign new_A9216_ = ~new_A9196_ & ~new_A9206_;
  assign new_A9215_ = new_A9196_ & new_A9206_;
  assign new_A9214_ = ~new_A9196_ | new_A9206_;
  assign new_A9213_ = new_A9180_ & ~new_A9181_;
  assign new_A9212_ = ~new_A9180_ & new_A9181_;
  assign new_A9211_ = new_A9233_ & ~new_A9234_;
  assign new_A9210_ = ~new_A9233_ & new_A9234_;
  assign new_A9209_ = ~new_A9232_ | ~new_A9231_;
  assign new_A9208_ = new_A9224_ | new_A9223_;
  assign new_A9207_ = new_A9230_ | new_A9229_;
  assign new_A9206_ = new_A9220_ | new_A9222_;
  assign new_A9205_ = ~new_A9227_ | ~new_A9228_;
  assign new_A9204_ = new_A9180_ & ~new_A9181_;
  assign new_A9203_ = new_A9194_ & ~new_A9206_;
  assign new_A9202_ = ~new_A9194_ & new_A9206_;
  assign new_A9201_ = ~new_A9192_ & new_A9218_;
  assign new_A9200_ = new_A9216_ | new_A9215_;
  assign new_A9199_ = new_A9213_ | new_A9212_;
  assign new_A9198_ = new_A9181_ | new_A9214_;
  assign new_A9197_ = new_A9206_ & new_A9209_;
  assign new_A9196_ = new_A9211_ | new_A9210_;
  assign new_A9195_ = new_A9206_ & new_A9205_;
  assign new_A9194_ = new_A9208_ & new_A9207_;
  assign new_A9193_ = new_A9203_ | new_A9202_;
  assign new_A9192_ = new_A9181_ | new_A9204_;
  assign A9191 = new_A9192_ | new_A9201_;
  assign A9190 = new_A9199_ & new_A9200_;
  assign A9189 = new_A9199_ & new_A9198_;
  assign A9188 = new_A9197_ | new_A9196_;
  assign A9187 = new_A9195_ | new_A9194_;
  assign A9186 = new_A9193_ & new_A9192_;
  assign new_A9185_ = new_C9690_;
  assign new_A9184_ = new_C9623_;
  assign new_A9183_ = new_C9556_;
  assign new_A9182_ = new_C9489_;
  assign new_A9181_ = new_C9422_;
  assign new_A9180_ = new_C9355_;
  assign new_A9179_ = ~new_A9118_ & new_A9132_;
  assign new_A9178_ = new_A9118_ & ~new_A9132_;
  assign new_A9177_ = new_A9118_ & ~new_A9132_;
  assign new_A9176_ = ~new_A9118_ & ~new_A9132_;
  assign new_A9175_ = new_A9118_ & new_A9132_;
  assign new_A9174_ = new_A9178_ | new_A9179_;
  assign new_A9173_ = ~new_A9118_ & new_A9132_;
  assign new_A9172_ = new_A9176_ | new_A9177_;
  assign new_A9171_ = ~new_A9147_ & ~new_A9167_;
  assign new_A9170_ = new_A9147_ & new_A9167_;
  assign new_A9169_ = ~new_A9114_ | ~new_A9139_;
  assign new_A9168_ = new_A9132_ & new_A9169_;
  assign new_A9167_ = new_A9115_ | new_A9116_;
  assign new_A9166_ = new_A9115_ | new_A9132_;
  assign new_A9165_ = ~new_A9132_ & ~new_A9168_;
  assign new_A9164_ = new_A9132_ | new_A9169_;
  assign new_A9163_ = new_A9115_ & ~new_A9116_;
  assign new_A9162_ = ~new_A9115_ & new_A9116_;
  assign new_A9161_ = new_A9125_ | new_A9158_;
  assign new_A9160_ = ~new_A9125_ & ~new_A9159_;
  assign new_A9159_ = new_A9125_ & new_A9158_;
  assign new_A9158_ = ~new_A9114_ | ~new_A9139_;
  assign new_A9157_ = ~new_A9115_ & new_A9125_;
  assign new_A9156_ = new_A9115_ & ~new_A9125_;
  assign new_A9155_ = new_A9117_ & new_A9154_;
  assign new_A9154_ = new_A9173_ | new_A9172_;
  assign new_A9153_ = ~new_A9117_ & new_A9152_;
  assign new_A9152_ = new_A9175_ | new_A9174_;
  assign new_A9151_ = new_A9117_ | new_A9150_;
  assign new_A9150_ = new_A9171_ | new_A9170_;
  assign new_A9149_ = ~new_A9129_ & ~new_A9139_;
  assign new_A9148_ = new_A9129_ & new_A9139_;
  assign new_A9147_ = ~new_A9129_ | new_A9139_;
  assign new_A9146_ = new_A9113_ & ~new_A9114_;
  assign new_A9145_ = ~new_A9113_ & new_A9114_;
  assign new_A9144_ = new_A9166_ & ~new_A9167_;
  assign new_A9143_ = ~new_A9166_ & new_A9167_;
  assign new_A9142_ = ~new_A9165_ | ~new_A9164_;
  assign new_A9141_ = new_A9157_ | new_A9156_;
  assign new_A9140_ = new_A9163_ | new_A9162_;
  assign new_A9139_ = new_A9153_ | new_A9155_;
  assign new_A9138_ = ~new_A9160_ | ~new_A9161_;
  assign new_A9137_ = new_A9113_ & ~new_A9114_;
  assign new_A9136_ = new_A9127_ & ~new_A9139_;
  assign new_A9135_ = ~new_A9127_ & new_A9139_;
  assign new_A9134_ = ~new_A9125_ & new_A9151_;
  assign new_A9133_ = new_A9149_ | new_A9148_;
  assign new_A9132_ = new_A9146_ | new_A9145_;
  assign new_A9131_ = new_A9114_ | new_A9147_;
  assign new_A9130_ = new_A9139_ & new_A9142_;
  assign new_A9129_ = new_A9144_ | new_A9143_;
  assign new_A9128_ = new_A9139_ & new_A9138_;
  assign new_A9127_ = new_A9141_ & new_A9140_;
  assign new_A9126_ = new_A9136_ | new_A9135_;
  assign new_A9125_ = new_A9114_ | new_A9137_;
  assign A9124 = new_A9125_ | new_A9134_;
  assign A9123 = new_A9132_ & new_A9133_;
  assign A9122 = new_A9132_ & new_A9131_;
  assign A9121 = new_A9130_ | new_A9129_;
  assign A9120 = new_A9128_ | new_A9127_;
  assign A9119 = new_A9126_ & new_A9125_;
  assign new_A9118_ = new_C9288_;
  assign new_A9117_ = new_C9221_;
  assign new_A9116_ = new_C9154_;
  assign new_A9115_ = new_C9087_;
  assign new_A9114_ = new_C9020_;
  assign new_A9113_ = new_C8953_;
  assign new_A9112_ = ~new_A9051_ & new_A9065_;
  assign new_A9111_ = new_A9051_ & ~new_A9065_;
  assign new_A9110_ = new_A9051_ & ~new_A9065_;
  assign new_A9109_ = ~new_A9051_ & ~new_A9065_;
  assign new_A9108_ = new_A9051_ & new_A9065_;
  assign new_A9107_ = new_A9111_ | new_A9112_;
  assign new_A9106_ = ~new_A9051_ & new_A9065_;
  assign new_A9105_ = new_A9109_ | new_A9110_;
  assign new_A9104_ = ~new_A9080_ & ~new_A9100_;
  assign new_A9103_ = new_A9080_ & new_A9100_;
  assign new_A9102_ = ~new_A9047_ | ~new_A9072_;
  assign new_A9101_ = new_A9065_ & new_A9102_;
  assign new_A9100_ = new_A9048_ | new_A9049_;
  assign new_A9099_ = new_A9048_ | new_A9065_;
  assign new_A9098_ = ~new_A9065_ & ~new_A9101_;
  assign new_A9097_ = new_A9065_ | new_A9102_;
  assign new_A9096_ = new_A9048_ & ~new_A9049_;
  assign new_A9095_ = ~new_A9048_ & new_A9049_;
  assign new_A9094_ = new_A9058_ | new_A9091_;
  assign new_A9093_ = ~new_A9058_ & ~new_A9092_;
  assign new_A9092_ = new_A9058_ & new_A9091_;
  assign new_A9091_ = ~new_A9047_ | ~new_A9072_;
  assign new_A9090_ = ~new_A9048_ & new_A9058_;
  assign new_A9089_ = new_A9048_ & ~new_A9058_;
  assign new_A9088_ = new_A9050_ & new_A9087_;
  assign new_A9087_ = new_A9106_ | new_A9105_;
  assign new_A9086_ = ~new_A9050_ & new_A9085_;
  assign new_A9085_ = new_A9108_ | new_A9107_;
  assign new_A9084_ = new_A9050_ | new_A9083_;
  assign new_A9083_ = new_A9104_ | new_A9103_;
  assign new_A9082_ = ~new_A9062_ & ~new_A9072_;
  assign new_A9081_ = new_A9062_ & new_A9072_;
  assign new_A9080_ = ~new_A9062_ | new_A9072_;
  assign new_A9079_ = new_A9046_ & ~new_A9047_;
  assign new_A9078_ = ~new_A9046_ & new_A9047_;
  assign new_A9077_ = new_A9099_ & ~new_A9100_;
  assign new_A9076_ = ~new_A9099_ & new_A9100_;
  assign new_A9075_ = ~new_A9098_ | ~new_A9097_;
  assign new_A9074_ = new_A9090_ | new_A9089_;
  assign new_A9073_ = new_A9096_ | new_A9095_;
  assign new_A9072_ = new_A9086_ | new_A9088_;
  assign new_A9071_ = ~new_A9093_ | ~new_A9094_;
  assign new_A9070_ = new_A9046_ & ~new_A9047_;
  assign new_A9069_ = new_A9060_ & ~new_A9072_;
  assign new_A9068_ = ~new_A9060_ & new_A9072_;
  assign new_A9067_ = ~new_A9058_ & new_A9084_;
  assign new_A9066_ = new_A9082_ | new_A9081_;
  assign new_A9065_ = new_A9079_ | new_A9078_;
  assign new_A9064_ = new_A9047_ | new_A9080_;
  assign new_A9063_ = new_A9072_ & new_A9075_;
  assign new_A9062_ = new_A9077_ | new_A9076_;
  assign new_A9061_ = new_A9072_ & new_A9071_;
  assign new_A9060_ = new_A9074_ & new_A9073_;
  assign new_A9059_ = new_A9069_ | new_A9068_;
  assign new_A9058_ = new_A9047_ | new_A9070_;
  assign A9057 = new_A9058_ | new_A9067_;
  assign A9056 = new_A9065_ & new_A9066_;
  assign A9055 = new_A9065_ & new_A9064_;
  assign A9054 = new_A9063_ | new_A9062_;
  assign A9053 = new_A9061_ | new_A9060_;
  assign A9052 = new_A9059_ & new_A9058_;
  assign new_A9051_ = new_C8886_;
  assign new_A9050_ = new_C8819_;
  assign new_A9049_ = new_C8752_;
  assign new_A9048_ = new_C8685_;
  assign new_A9047_ = new_C8618_;
  assign new_A9046_ = new_C8551_;
  assign new_A9045_ = ~new_A8984_ & new_A8998_;
  assign new_A9044_ = new_A8984_ & ~new_A8998_;
  assign new_A9043_ = new_A8984_ & ~new_A8998_;
  assign new_A9042_ = ~new_A8984_ & ~new_A8998_;
  assign new_A9041_ = new_A8984_ & new_A8998_;
  assign new_A9040_ = new_A9044_ | new_A9045_;
  assign new_A9039_ = ~new_A8984_ & new_A8998_;
  assign new_A9038_ = new_A9042_ | new_A9043_;
  assign new_A9037_ = ~new_A9013_ & ~new_A9033_;
  assign new_A9036_ = new_A9013_ & new_A9033_;
  assign new_A9035_ = ~new_A8980_ | ~new_A9005_;
  assign new_A9034_ = new_A8998_ & new_A9035_;
  assign new_A9033_ = new_A8981_ | new_A8982_;
  assign new_A9032_ = new_A8981_ | new_A8998_;
  assign new_A9031_ = ~new_A8998_ & ~new_A9034_;
  assign new_A9030_ = new_A8998_ | new_A9035_;
  assign new_A9029_ = new_A8981_ & ~new_A8982_;
  assign new_A9028_ = ~new_A8981_ & new_A8982_;
  assign new_A9027_ = new_A8991_ | new_A9024_;
  assign new_A9026_ = ~new_A8991_ & ~new_A9025_;
  assign new_A9025_ = new_A8991_ & new_A9024_;
  assign new_A9024_ = ~new_A8980_ | ~new_A9005_;
  assign new_A9023_ = ~new_A8981_ & new_A8991_;
  assign new_A9022_ = new_A8981_ & ~new_A8991_;
  assign new_A9021_ = new_A8983_ & new_A9020_;
  assign new_A9020_ = new_A9039_ | new_A9038_;
  assign new_A9019_ = ~new_A8983_ & new_A9018_;
  assign new_A9018_ = new_A9041_ | new_A9040_;
  assign new_A9017_ = new_A8983_ | new_A9016_;
  assign new_A9016_ = new_A9037_ | new_A9036_;
  assign new_A9015_ = ~new_A8995_ & ~new_A9005_;
  assign new_A9014_ = new_A8995_ & new_A9005_;
  assign new_A9013_ = ~new_A8995_ | new_A9005_;
  assign new_A9012_ = new_A8979_ & ~new_A8980_;
  assign new_A9011_ = ~new_A8979_ & new_A8980_;
  assign new_A9010_ = new_A9032_ & ~new_A9033_;
  assign new_A9009_ = ~new_A9032_ & new_A9033_;
  assign new_A9008_ = ~new_A9031_ | ~new_A9030_;
  assign new_A9007_ = new_A9023_ | new_A9022_;
  assign new_A9006_ = new_A9029_ | new_A9028_;
  assign new_A9005_ = new_A9019_ | new_A9021_;
  assign new_A9004_ = ~new_A9026_ | ~new_A9027_;
  assign new_A9003_ = new_A8979_ & ~new_A8980_;
  assign new_A9002_ = new_A8993_ & ~new_A9005_;
  assign new_A9001_ = ~new_A8993_ & new_A9005_;
  assign new_A9000_ = ~new_A8991_ & new_A9017_;
  assign new_A8999_ = new_A9015_ | new_A9014_;
  assign new_A8998_ = new_A9012_ | new_A9011_;
  assign new_A8997_ = new_A8980_ | new_A9013_;
  assign new_A8996_ = new_A9005_ & new_A9008_;
  assign new_A8995_ = new_A9010_ | new_A9009_;
  assign new_A8994_ = new_A9005_ & new_A9004_;
  assign new_A8993_ = new_A9007_ & new_A9006_;
  assign new_A8992_ = new_A9002_ | new_A9001_;
  assign new_A8991_ = new_A8980_ | new_A9003_;
  assign A8990 = new_A8991_ | new_A9000_;
  assign A8989 = new_A8998_ & new_A8999_;
  assign A8988 = new_A8998_ & new_A8997_;
  assign A8987 = new_A8996_ | new_A8995_;
  assign A8986 = new_A8994_ | new_A8993_;
  assign A8985 = new_A8992_ & new_A8991_;
  assign new_A8984_ = new_C8484_;
  assign new_A8983_ = new_C8417_;
  assign new_A8982_ = new_C8350_;
  assign new_A8981_ = new_C8283_;
  assign new_A8980_ = new_C8216_;
  assign new_A8979_ = new_C8149_;
  assign new_A8978_ = ~new_A8917_ & new_A8931_;
  assign new_A8977_ = new_A8917_ & ~new_A8931_;
  assign new_A8976_ = new_A8917_ & ~new_A8931_;
  assign new_A8975_ = ~new_A8917_ & ~new_A8931_;
  assign new_A8974_ = new_A8917_ & new_A8931_;
  assign new_A8973_ = new_A8977_ | new_A8978_;
  assign new_A8972_ = ~new_A8917_ & new_A8931_;
  assign new_A8971_ = new_A8975_ | new_A8976_;
  assign new_A8970_ = ~new_A8946_ & ~new_A8966_;
  assign new_A8969_ = new_A8946_ & new_A8966_;
  assign new_A8968_ = ~new_A8913_ | ~new_A8938_;
  assign new_A8967_ = new_A8931_ & new_A8968_;
  assign new_A8966_ = new_A8914_ | new_A8915_;
  assign new_A8965_ = new_A8914_ | new_A8931_;
  assign new_A8964_ = ~new_A8931_ & ~new_A8967_;
  assign new_A8963_ = new_A8931_ | new_A8968_;
  assign new_A8962_ = new_A8914_ & ~new_A8915_;
  assign new_A8961_ = ~new_A8914_ & new_A8915_;
  assign new_A8960_ = new_A8924_ | new_A8957_;
  assign new_A8959_ = ~new_A8924_ & ~new_A8958_;
  assign new_A8958_ = new_A8924_ & new_A8957_;
  assign new_A8957_ = ~new_A8913_ | ~new_A8938_;
  assign new_A8956_ = ~new_A8914_ & new_A8924_;
  assign new_A8955_ = new_A8914_ & ~new_A8924_;
  assign new_A8954_ = new_A8916_ & new_A8953_;
  assign new_A8953_ = new_A8972_ | new_A8971_;
  assign new_A8952_ = ~new_A8916_ & new_A8951_;
  assign new_A8951_ = new_A8974_ | new_A8973_;
  assign new_A8950_ = new_A8916_ | new_A8949_;
  assign new_A8949_ = new_A8970_ | new_A8969_;
  assign new_A8948_ = ~new_A8928_ & ~new_A8938_;
  assign new_A8947_ = new_A8928_ & new_A8938_;
  assign new_A8946_ = ~new_A8928_ | new_A8938_;
  assign new_A8945_ = new_A8912_ & ~new_A8913_;
  assign new_A8944_ = ~new_A8912_ & new_A8913_;
  assign new_A8943_ = new_A8965_ & ~new_A8966_;
  assign new_A8942_ = ~new_A8965_ & new_A8966_;
  assign new_A8941_ = ~new_A8964_ | ~new_A8963_;
  assign new_A8940_ = new_A8956_ | new_A8955_;
  assign new_A8939_ = new_A8962_ | new_A8961_;
  assign new_A8938_ = new_A8952_ | new_A8954_;
  assign new_A8937_ = ~new_A8959_ | ~new_A8960_;
  assign new_A8936_ = new_A8912_ & ~new_A8913_;
  assign new_A8935_ = new_A8926_ & ~new_A8938_;
  assign new_A8934_ = ~new_A8926_ & new_A8938_;
  assign new_A8933_ = ~new_A8924_ & new_A8950_;
  assign new_A8932_ = new_A8948_ | new_A8947_;
  assign new_A8931_ = new_A8945_ | new_A8944_;
  assign new_A8930_ = new_A8913_ | new_A8946_;
  assign new_A8929_ = new_A8938_ & new_A8941_;
  assign new_A8928_ = new_A8943_ | new_A8942_;
  assign new_A8927_ = new_A8938_ & new_A8937_;
  assign new_A8926_ = new_A8940_ & new_A8939_;
  assign new_A8925_ = new_A8935_ | new_A8934_;
  assign new_A8924_ = new_A8913_ | new_A8936_;
  assign A8923 = new_A8924_ | new_A8933_;
  assign A8922 = new_A8931_ & new_A8932_;
  assign A8921 = new_A8931_ & new_A8930_;
  assign A8920 = new_A8929_ | new_A8928_;
  assign A8919 = new_A8927_ | new_A8926_;
  assign A8918 = new_A8925_ & new_A8924_;
  assign new_A8917_ = new_C8082_;
  assign new_A8916_ = new_C8015_;
  assign new_A8915_ = new_C7948_;
  assign new_A8914_ = new_C7881_;
  assign new_A8913_ = new_C7814_;
  assign new_A8912_ = new_C7747_;
  assign new_A8911_ = ~new_A8850_ & new_A8864_;
  assign new_A8910_ = new_A8850_ & ~new_A8864_;
  assign new_A8909_ = new_A8850_ & ~new_A8864_;
  assign new_A8908_ = ~new_A8850_ & ~new_A8864_;
  assign new_A8907_ = new_A8850_ & new_A8864_;
  assign new_A8906_ = new_A8910_ | new_A8911_;
  assign new_A8905_ = ~new_A8850_ & new_A8864_;
  assign new_A8904_ = new_A8908_ | new_A8909_;
  assign new_A8903_ = ~new_A8879_ & ~new_A8899_;
  assign new_A8902_ = new_A8879_ & new_A8899_;
  assign new_A8901_ = ~new_A8846_ | ~new_A8871_;
  assign new_A8900_ = new_A8864_ & new_A8901_;
  assign new_A8899_ = new_A8847_ | new_A8848_;
  assign new_A8898_ = new_A8847_ | new_A8864_;
  assign new_A8897_ = ~new_A8864_ & ~new_A8900_;
  assign new_A8896_ = new_A8864_ | new_A8901_;
  assign new_A8895_ = new_A8847_ & ~new_A8848_;
  assign new_A8894_ = ~new_A8847_ & new_A8848_;
  assign new_A8893_ = new_A8857_ | new_A8890_;
  assign new_A8892_ = ~new_A8857_ & ~new_A8891_;
  assign new_A8891_ = new_A8857_ & new_A8890_;
  assign new_A8890_ = ~new_A8846_ | ~new_A8871_;
  assign new_A8889_ = ~new_A8847_ & new_A8857_;
  assign new_A8888_ = new_A8847_ & ~new_A8857_;
  assign new_A8887_ = new_A8849_ & new_A8886_;
  assign new_A8886_ = new_A8905_ | new_A8904_;
  assign new_A8885_ = ~new_A8849_ & new_A8884_;
  assign new_A8884_ = new_A8907_ | new_A8906_;
  assign new_A8883_ = new_A8849_ | new_A8882_;
  assign new_A8882_ = new_A8903_ | new_A8902_;
  assign new_A8881_ = ~new_A8861_ & ~new_A8871_;
  assign new_A8880_ = new_A8861_ & new_A8871_;
  assign new_A8879_ = ~new_A8861_ | new_A8871_;
  assign new_A8878_ = new_A8845_ & ~new_A8846_;
  assign new_A8877_ = ~new_A8845_ & new_A8846_;
  assign new_A8876_ = new_A8898_ & ~new_A8899_;
  assign new_A8875_ = ~new_A8898_ & new_A8899_;
  assign new_A8874_ = ~new_A8897_ | ~new_A8896_;
  assign new_A8873_ = new_A8889_ | new_A8888_;
  assign new_A8872_ = new_A8895_ | new_A8894_;
  assign new_A8871_ = new_A8885_ | new_A8887_;
  assign new_A8870_ = ~new_A8892_ | ~new_A8893_;
  assign new_A8869_ = new_A8845_ & ~new_A8846_;
  assign new_A8868_ = new_A8859_ & ~new_A8871_;
  assign new_A8867_ = ~new_A8859_ & new_A8871_;
  assign new_A8866_ = ~new_A8857_ & new_A8883_;
  assign new_A8865_ = new_A8881_ | new_A8880_;
  assign new_A8864_ = new_A8878_ | new_A8877_;
  assign new_A8863_ = new_A8846_ | new_A8879_;
  assign new_A8862_ = new_A8871_ & new_A8874_;
  assign new_A8861_ = new_A8876_ | new_A8875_;
  assign new_A8860_ = new_A8871_ & new_A8870_;
  assign new_A8859_ = new_A8873_ & new_A8872_;
  assign new_A8858_ = new_A8868_ | new_A8867_;
  assign new_A8857_ = new_A8846_ | new_A8869_;
  assign A8856 = new_A8857_ | new_A8866_;
  assign A8855 = new_A8864_ & new_A8865_;
  assign A8854 = new_A8864_ & new_A8863_;
  assign A8853 = new_A8862_ | new_A8861_;
  assign A8852 = new_A8860_ | new_A8859_;
  assign A8851 = new_A8858_ & new_A8857_;
  assign new_A8850_ = new_C7680_;
  assign new_A8849_ = new_C7613_;
  assign new_A8848_ = new_C7546_;
  assign new_A8847_ = new_C7479_;
  assign new_A8846_ = new_C7412_;
  assign new_A8845_ = new_C7345_;
  assign new_A8844_ = ~new_A8783_ & new_A8797_;
  assign new_A8843_ = new_A8783_ & ~new_A8797_;
  assign new_A8842_ = new_A8783_ & ~new_A8797_;
  assign new_A8841_ = ~new_A8783_ & ~new_A8797_;
  assign new_A8840_ = new_A8783_ & new_A8797_;
  assign new_A8839_ = new_A8843_ | new_A8844_;
  assign new_A8838_ = ~new_A8783_ & new_A8797_;
  assign new_A8837_ = new_A8841_ | new_A8842_;
  assign new_A8836_ = ~new_A8812_ & ~new_A8832_;
  assign new_A8835_ = new_A8812_ & new_A8832_;
  assign new_A8834_ = ~new_A8779_ | ~new_A8804_;
  assign new_A8833_ = new_A8797_ & new_A8834_;
  assign new_A8832_ = new_A8780_ | new_A8781_;
  assign new_A8831_ = new_A8780_ | new_A8797_;
  assign new_A8830_ = ~new_A8797_ & ~new_A8833_;
  assign new_A8829_ = new_A8797_ | new_A8834_;
  assign new_A8828_ = new_A8780_ & ~new_A8781_;
  assign new_A8827_ = ~new_A8780_ & new_A8781_;
  assign new_A8826_ = new_A8790_ | new_A8823_;
  assign new_A8825_ = ~new_A8790_ & ~new_A8824_;
  assign new_A8824_ = new_A8790_ & new_A8823_;
  assign new_A8823_ = ~new_A8779_ | ~new_A8804_;
  assign new_A8822_ = ~new_A8780_ & new_A8790_;
  assign new_A8821_ = new_A8780_ & ~new_A8790_;
  assign new_A8820_ = new_A8782_ & new_A8819_;
  assign new_A8819_ = new_A8838_ | new_A8837_;
  assign new_A8818_ = ~new_A8782_ & new_A8817_;
  assign new_A8817_ = new_A8840_ | new_A8839_;
  assign new_A8816_ = new_A8782_ | new_A8815_;
  assign new_A8815_ = new_A8836_ | new_A8835_;
  assign new_A8814_ = ~new_A8794_ & ~new_A8804_;
  assign new_A8813_ = new_A8794_ & new_A8804_;
  assign new_A8812_ = ~new_A8794_ | new_A8804_;
  assign new_A8811_ = new_A8778_ & ~new_A8779_;
  assign new_A8810_ = ~new_A8778_ & new_A8779_;
  assign new_A8809_ = new_A8831_ & ~new_A8832_;
  assign new_A8808_ = ~new_A8831_ & new_A8832_;
  assign new_A8807_ = ~new_A8830_ | ~new_A8829_;
  assign new_A8806_ = new_A8822_ | new_A8821_;
  assign new_A8805_ = new_A8828_ | new_A8827_;
  assign new_A8804_ = new_A8818_ | new_A8820_;
  assign new_A8803_ = ~new_A8825_ | ~new_A8826_;
  assign new_A8802_ = new_A8778_ & ~new_A8779_;
  assign new_A8801_ = new_A8792_ & ~new_A8804_;
  assign new_A8800_ = ~new_A8792_ & new_A8804_;
  assign new_A8799_ = ~new_A8790_ & new_A8816_;
  assign new_A8798_ = new_A8814_ | new_A8813_;
  assign new_A8797_ = new_A8811_ | new_A8810_;
  assign new_A8796_ = new_A8779_ | new_A8812_;
  assign new_A8795_ = new_A8804_ & new_A8807_;
  assign new_A8794_ = new_A8809_ | new_A8808_;
  assign new_A8793_ = new_A8804_ & new_A8803_;
  assign new_A8792_ = new_A8806_ & new_A8805_;
  assign new_A8791_ = new_A8801_ | new_A8800_;
  assign new_A8790_ = new_A8779_ | new_A8802_;
  assign A8789 = new_A8790_ | new_A8799_;
  assign A8788 = new_A8797_ & new_A8798_;
  assign A8787 = new_A8797_ & new_A8796_;
  assign A8786 = new_A8795_ | new_A8794_;
  assign A8785 = new_A8793_ | new_A8792_;
  assign A8784 = new_A8791_ & new_A8790_;
  assign new_A8783_ = new_C7278_;
  assign new_A8782_ = new_C7211_;
  assign new_A8781_ = new_C7144_;
  assign new_A8780_ = new_C7077_;
  assign new_A8779_ = new_C7010_;
  assign new_A8778_ = new_C6943_;
  assign new_A8777_ = ~new_A8716_ & new_A8730_;
  assign new_A8776_ = new_A8716_ & ~new_A8730_;
  assign new_A8775_ = new_A8716_ & ~new_A8730_;
  assign new_A8774_ = ~new_A8716_ & ~new_A8730_;
  assign new_A8773_ = new_A8716_ & new_A8730_;
  assign new_A8772_ = new_A8776_ | new_A8777_;
  assign new_A8771_ = ~new_A8716_ & new_A8730_;
  assign new_A8770_ = new_A8774_ | new_A8775_;
  assign new_A8769_ = ~new_A8745_ & ~new_A8765_;
  assign new_A8768_ = new_A8745_ & new_A8765_;
  assign new_A8767_ = ~new_A8712_ | ~new_A8737_;
  assign new_A8766_ = new_A8730_ & new_A8767_;
  assign new_A8765_ = new_A8713_ | new_A8714_;
  assign new_A8764_ = new_A8713_ | new_A8730_;
  assign new_A8763_ = ~new_A8730_ & ~new_A8766_;
  assign new_A8762_ = new_A8730_ | new_A8767_;
  assign new_A8761_ = new_A8713_ & ~new_A8714_;
  assign new_A8760_ = ~new_A8713_ & new_A8714_;
  assign new_A8759_ = new_A8723_ | new_A8756_;
  assign new_A8758_ = ~new_A8723_ & ~new_A8757_;
  assign new_A8757_ = new_A8723_ & new_A8756_;
  assign new_A8756_ = ~new_A8712_ | ~new_A8737_;
  assign new_A8755_ = ~new_A8713_ & new_A8723_;
  assign new_A8754_ = new_A8713_ & ~new_A8723_;
  assign new_A8753_ = new_A8715_ & new_A8752_;
  assign new_A8752_ = new_A8771_ | new_A8770_;
  assign new_A8751_ = ~new_A8715_ & new_A8750_;
  assign new_A8750_ = new_A8773_ | new_A8772_;
  assign new_A8749_ = new_A8715_ | new_A8748_;
  assign new_A8748_ = new_A8769_ | new_A8768_;
  assign new_A8747_ = ~new_A8727_ & ~new_A8737_;
  assign new_A8746_ = new_A8727_ & new_A8737_;
  assign new_A8745_ = ~new_A8727_ | new_A8737_;
  assign new_A8744_ = new_A8711_ & ~new_A8712_;
  assign new_A8743_ = ~new_A8711_ & new_A8712_;
  assign new_A8742_ = new_A8764_ & ~new_A8765_;
  assign new_A8741_ = ~new_A8764_ & new_A8765_;
  assign new_A8740_ = ~new_A8763_ | ~new_A8762_;
  assign new_A8739_ = new_A8755_ | new_A8754_;
  assign new_A8738_ = new_A8761_ | new_A8760_;
  assign new_A8737_ = new_A8751_ | new_A8753_;
  assign new_A8736_ = ~new_A8758_ | ~new_A8759_;
  assign new_A8735_ = new_A8711_ & ~new_A8712_;
  assign new_A8734_ = new_A8725_ & ~new_A8737_;
  assign new_A8733_ = ~new_A8725_ & new_A8737_;
  assign new_A8732_ = ~new_A8723_ & new_A8749_;
  assign new_A8731_ = new_A8747_ | new_A8746_;
  assign new_A8730_ = new_A8744_ | new_A8743_;
  assign new_A8729_ = new_A8712_ | new_A8745_;
  assign new_A8728_ = new_A8737_ & new_A8740_;
  assign new_A8727_ = new_A8742_ | new_A8741_;
  assign new_A8726_ = new_A8737_ & new_A8736_;
  assign new_A8725_ = new_A8739_ & new_A8738_;
  assign new_A8724_ = new_A8734_ | new_A8733_;
  assign new_A8723_ = new_A8712_ | new_A8735_;
  assign A8722 = new_A8723_ | new_A8732_;
  assign A8721 = new_A8730_ & new_A8731_;
  assign A8720 = new_A8730_ & new_A8729_;
  assign A8719 = new_A8728_ | new_A8727_;
  assign A8718 = new_A8726_ | new_A8725_;
  assign A8717 = new_A8724_ & new_A8723_;
  assign new_A8716_ = new_C6876_;
  assign new_A8715_ = new_C6809_;
  assign new_A8714_ = new_C6742_;
  assign new_A8713_ = new_C6675_;
  assign new_A8712_ = new_C6608_;
  assign new_A8711_ = new_C6541_;
  assign new_A8710_ = ~new_A8649_ & new_A8663_;
  assign new_A8709_ = new_A8649_ & ~new_A8663_;
  assign new_A8708_ = new_A8649_ & ~new_A8663_;
  assign new_A8707_ = ~new_A8649_ & ~new_A8663_;
  assign new_A8706_ = new_A8649_ & new_A8663_;
  assign new_A8705_ = new_A8709_ | new_A8710_;
  assign new_A8704_ = ~new_A8649_ & new_A8663_;
  assign new_A8703_ = new_A8707_ | new_A8708_;
  assign new_A8702_ = ~new_A8678_ & ~new_A8698_;
  assign new_A8701_ = new_A8678_ & new_A8698_;
  assign new_A8700_ = ~new_A8645_ | ~new_A8670_;
  assign new_A8699_ = new_A8663_ & new_A8700_;
  assign new_A8698_ = new_A8646_ | new_A8647_;
  assign new_A8697_ = new_A8646_ | new_A8663_;
  assign new_A8696_ = ~new_A8663_ & ~new_A8699_;
  assign new_A8695_ = new_A8663_ | new_A8700_;
  assign new_A8694_ = new_A8646_ & ~new_A8647_;
  assign new_A8693_ = ~new_A8646_ & new_A8647_;
  assign new_A8692_ = new_A8656_ | new_A8689_;
  assign new_A8691_ = ~new_A8656_ & ~new_A8690_;
  assign new_A8690_ = new_A8656_ & new_A8689_;
  assign new_A8689_ = ~new_A8645_ | ~new_A8670_;
  assign new_A8688_ = ~new_A8646_ & new_A8656_;
  assign new_A8687_ = new_A8646_ & ~new_A8656_;
  assign new_A8686_ = new_A8648_ & new_A8685_;
  assign new_A8685_ = new_A8704_ | new_A8703_;
  assign new_A8684_ = ~new_A8648_ & new_A8683_;
  assign new_A8683_ = new_A8706_ | new_A8705_;
  assign new_A8682_ = new_A8648_ | new_A8681_;
  assign new_A8681_ = new_A8702_ | new_A8701_;
  assign new_A8680_ = ~new_A8660_ & ~new_A8670_;
  assign new_A8679_ = new_A8660_ & new_A8670_;
  assign new_A8678_ = ~new_A8660_ | new_A8670_;
  assign new_A8677_ = new_A8644_ & ~new_A8645_;
  assign new_A8676_ = ~new_A8644_ & new_A8645_;
  assign new_A8675_ = new_A8697_ & ~new_A8698_;
  assign new_A8674_ = ~new_A8697_ & new_A8698_;
  assign new_A8673_ = ~new_A8696_ | ~new_A8695_;
  assign new_A8672_ = new_A8688_ | new_A8687_;
  assign new_A8671_ = new_A8694_ | new_A8693_;
  assign new_A8670_ = new_A8684_ | new_A8686_;
  assign new_A8669_ = ~new_A8691_ | ~new_A8692_;
  assign new_A8668_ = new_A8644_ & ~new_A8645_;
  assign new_A8667_ = new_A8658_ & ~new_A8670_;
  assign new_A8666_ = ~new_A8658_ & new_A8670_;
  assign new_A8665_ = ~new_A8656_ & new_A8682_;
  assign new_A8664_ = new_A8680_ | new_A8679_;
  assign new_A8663_ = new_A8677_ | new_A8676_;
  assign new_A8662_ = new_A8645_ | new_A8678_;
  assign new_A8661_ = new_A8670_ & new_A8673_;
  assign new_A8660_ = new_A8675_ | new_A8674_;
  assign new_A8659_ = new_A8670_ & new_A8669_;
  assign new_A8658_ = new_A8672_ & new_A8671_;
  assign new_A8657_ = new_A8667_ | new_A8666_;
  assign new_A8656_ = new_A8645_ | new_A8668_;
  assign A8655 = new_A8656_ | new_A8665_;
  assign A8654 = new_A8663_ & new_A8664_;
  assign A8653 = new_A8663_ & new_A8662_;
  assign A8652 = new_A8661_ | new_A8660_;
  assign A8651 = new_A8659_ | new_A8658_;
  assign A8650 = new_A8657_ & new_A8656_;
  assign new_A8649_ = new_C6474_;
  assign new_A8648_ = new_C6407_;
  assign new_A8647_ = new_C6340_;
  assign new_A8646_ = new_C6273_;
  assign new_A8645_ = new_C6206_;
  assign new_A8644_ = new_C6139_;
  assign new_A8643_ = ~new_A8582_ & new_A8596_;
  assign new_A8642_ = new_A8582_ & ~new_A8596_;
  assign new_A8641_ = new_A8582_ & ~new_A8596_;
  assign new_A8640_ = ~new_A8582_ & ~new_A8596_;
  assign new_A8639_ = new_A8582_ & new_A8596_;
  assign new_A8638_ = new_A8642_ | new_A8643_;
  assign new_A8637_ = ~new_A8582_ & new_A8596_;
  assign new_A8636_ = new_A8640_ | new_A8641_;
  assign new_A8635_ = ~new_A8611_ & ~new_A8631_;
  assign new_A8634_ = new_A8611_ & new_A8631_;
  assign new_A8633_ = ~new_A8578_ | ~new_A8603_;
  assign new_A8632_ = new_A8596_ & new_A8633_;
  assign new_A8631_ = new_A8579_ | new_A8580_;
  assign new_A8630_ = new_A8579_ | new_A8596_;
  assign new_A8629_ = ~new_A8596_ & ~new_A8632_;
  assign new_A8628_ = new_A8596_ | new_A8633_;
  assign new_A8627_ = new_A8579_ & ~new_A8580_;
  assign new_A8626_ = ~new_A8579_ & new_A8580_;
  assign new_A8625_ = new_A8589_ | new_A8622_;
  assign new_A8624_ = ~new_A8589_ & ~new_A8623_;
  assign new_A8623_ = new_A8589_ & new_A8622_;
  assign new_A8622_ = ~new_A8578_ | ~new_A8603_;
  assign new_A8621_ = ~new_A8579_ & new_A8589_;
  assign new_A8620_ = new_A8579_ & ~new_A8589_;
  assign new_A8619_ = new_A8581_ & new_A8618_;
  assign new_A8618_ = new_A8637_ | new_A8636_;
  assign new_A8617_ = ~new_A8581_ & new_A8616_;
  assign new_A8616_ = new_A8639_ | new_A8638_;
  assign new_A8615_ = new_A8581_ | new_A8614_;
  assign new_A8614_ = new_A8635_ | new_A8634_;
  assign new_A8613_ = ~new_A8593_ & ~new_A8603_;
  assign new_A8612_ = new_A8593_ & new_A8603_;
  assign new_A8611_ = ~new_A8593_ | new_A8603_;
  assign new_A8610_ = new_A8577_ & ~new_A8578_;
  assign new_A8609_ = ~new_A8577_ & new_A8578_;
  assign new_A8608_ = new_A8630_ & ~new_A8631_;
  assign new_A8607_ = ~new_A8630_ & new_A8631_;
  assign new_A8606_ = ~new_A8629_ | ~new_A8628_;
  assign new_A8605_ = new_A8621_ | new_A8620_;
  assign new_A8604_ = new_A8627_ | new_A8626_;
  assign new_A8603_ = new_A8617_ | new_A8619_;
  assign new_A8602_ = ~new_A8624_ | ~new_A8625_;
  assign new_A8601_ = new_A8577_ & ~new_A8578_;
  assign new_A8600_ = new_A8591_ & ~new_A8603_;
  assign new_A8599_ = ~new_A8591_ & new_A8603_;
  assign new_A8598_ = ~new_A8589_ & new_A8615_;
  assign new_A8597_ = new_A8613_ | new_A8612_;
  assign new_A8596_ = new_A8610_ | new_A8609_;
  assign new_A8595_ = new_A8578_ | new_A8611_;
  assign new_A8594_ = new_A8603_ & new_A8606_;
  assign new_A8593_ = new_A8608_ | new_A8607_;
  assign new_A8592_ = new_A8603_ & new_A8602_;
  assign new_A8591_ = new_A8605_ & new_A8604_;
  assign new_A8590_ = new_A8600_ | new_A8599_;
  assign new_A8589_ = new_A8578_ | new_A8601_;
  assign A8588 = new_A8589_ | new_A8598_;
  assign A8587 = new_A8596_ & new_A8597_;
  assign A8586 = new_A8596_ & new_A8595_;
  assign A8585 = new_A8594_ | new_A8593_;
  assign A8584 = new_A8592_ | new_A8591_;
  assign A8583 = new_A8590_ & new_A8589_;
  assign new_A8582_ = new_C6072_;
  assign new_A8581_ = new_C6005_;
  assign new_A8580_ = new_C5938_;
  assign new_A8579_ = new_C5871_;
  assign new_A8578_ = new_C5804_;
  assign new_A8577_ = new_C5737_;
  assign new_A8576_ = ~new_A8515_ & new_A8529_;
  assign new_A8575_ = new_A8515_ & ~new_A8529_;
  assign new_A8574_ = new_A8515_ & ~new_A8529_;
  assign new_A8573_ = ~new_A8515_ & ~new_A8529_;
  assign new_A8572_ = new_A8515_ & new_A8529_;
  assign new_A8571_ = new_A8575_ | new_A8576_;
  assign new_A8570_ = ~new_A8515_ & new_A8529_;
  assign new_A8569_ = new_A8573_ | new_A8574_;
  assign new_A8568_ = ~new_A8544_ & ~new_A8564_;
  assign new_A8567_ = new_A8544_ & new_A8564_;
  assign new_A8566_ = ~new_A8511_ | ~new_A8536_;
  assign new_A8565_ = new_A8529_ & new_A8566_;
  assign new_A8564_ = new_A8512_ | new_A8513_;
  assign new_A8563_ = new_A8512_ | new_A8529_;
  assign new_A8562_ = ~new_A8529_ & ~new_A8565_;
  assign new_A8561_ = new_A8529_ | new_A8566_;
  assign new_A8560_ = new_A8512_ & ~new_A8513_;
  assign new_A8559_ = ~new_A8512_ & new_A8513_;
  assign new_A8558_ = new_A8522_ | new_A8555_;
  assign new_A8557_ = ~new_A8522_ & ~new_A8556_;
  assign new_A8556_ = new_A8522_ & new_A8555_;
  assign new_A8555_ = ~new_A8511_ | ~new_A8536_;
  assign new_A8554_ = ~new_A8512_ & new_A8522_;
  assign new_A8553_ = new_A8512_ & ~new_A8522_;
  assign new_A8552_ = new_A8514_ & new_A8551_;
  assign new_A8551_ = new_A8570_ | new_A8569_;
  assign new_A8550_ = ~new_A8514_ & new_A8549_;
  assign new_A8549_ = new_A8572_ | new_A8571_;
  assign new_A8548_ = new_A8514_ | new_A8547_;
  assign new_A8547_ = new_A8568_ | new_A8567_;
  assign new_A8546_ = ~new_A8526_ & ~new_A8536_;
  assign new_A8545_ = new_A8526_ & new_A8536_;
  assign new_A8544_ = ~new_A8526_ | new_A8536_;
  assign new_A8543_ = new_A8510_ & ~new_A8511_;
  assign new_A8542_ = ~new_A8510_ & new_A8511_;
  assign new_A8541_ = new_A8563_ & ~new_A8564_;
  assign new_A8540_ = ~new_A8563_ & new_A8564_;
  assign new_A8539_ = ~new_A8562_ | ~new_A8561_;
  assign new_A8538_ = new_A8554_ | new_A8553_;
  assign new_A8537_ = new_A8560_ | new_A8559_;
  assign new_A8536_ = new_A8550_ | new_A8552_;
  assign new_A8535_ = ~new_A8557_ | ~new_A8558_;
  assign new_A8534_ = new_A8510_ & ~new_A8511_;
  assign new_A8533_ = new_A8524_ & ~new_A8536_;
  assign new_A8532_ = ~new_A8524_ & new_A8536_;
  assign new_A8531_ = ~new_A8522_ & new_A8548_;
  assign new_A8530_ = new_A8546_ | new_A8545_;
  assign new_A8529_ = new_A8543_ | new_A8542_;
  assign new_A8528_ = new_A8511_ | new_A8544_;
  assign new_A8527_ = new_A8536_ & new_A8539_;
  assign new_A8526_ = new_A8541_ | new_A8540_;
  assign new_A8525_ = new_A8536_ & new_A8535_;
  assign new_A8524_ = new_A8538_ & new_A8537_;
  assign new_A8523_ = new_A8533_ | new_A8532_;
  assign new_A8522_ = new_A8511_ | new_A8534_;
  assign A8521 = new_A8522_ | new_A8531_;
  assign A8520 = new_A8529_ & new_A8530_;
  assign A8519 = new_A8529_ & new_A8528_;
  assign A8518 = new_A8527_ | new_A8526_;
  assign A8517 = new_A8525_ | new_A8524_;
  assign A8516 = new_A8523_ & new_A8522_;
  assign new_A8515_ = new_C5670_;
  assign new_A8514_ = new_C5603_;
  assign new_A8513_ = new_C5536_;
  assign new_A8512_ = new_C5469_;
  assign new_A8511_ = new_C5402_;
  assign new_A8510_ = new_C5335_;
  assign new_A8509_ = ~new_A8448_ & new_A8462_;
  assign new_A8508_ = new_A8448_ & ~new_A8462_;
  assign new_A8507_ = new_A8448_ & ~new_A8462_;
  assign new_A8506_ = ~new_A8448_ & ~new_A8462_;
  assign new_A8505_ = new_A8448_ & new_A8462_;
  assign new_A8504_ = new_A8508_ | new_A8509_;
  assign new_A8503_ = ~new_A8448_ & new_A8462_;
  assign new_A8502_ = new_A8506_ | new_A8507_;
  assign new_A8501_ = ~new_A8477_ & ~new_A8497_;
  assign new_A8500_ = new_A8477_ & new_A8497_;
  assign new_A8499_ = ~new_A8444_ | ~new_A8469_;
  assign new_A8498_ = new_A8462_ & new_A8499_;
  assign new_A8497_ = new_A8445_ | new_A8446_;
  assign new_A8496_ = new_A8445_ | new_A8462_;
  assign new_A8495_ = ~new_A8462_ & ~new_A8498_;
  assign new_A8494_ = new_A8462_ | new_A8499_;
  assign new_A8493_ = new_A8445_ & ~new_A8446_;
  assign new_A8492_ = ~new_A8445_ & new_A8446_;
  assign new_A8491_ = new_A8455_ | new_A8488_;
  assign new_A8490_ = ~new_A8455_ & ~new_A8489_;
  assign new_A8489_ = new_A8455_ & new_A8488_;
  assign new_A8488_ = ~new_A8444_ | ~new_A8469_;
  assign new_A8487_ = ~new_A8445_ & new_A8455_;
  assign new_A8486_ = new_A8445_ & ~new_A8455_;
  assign new_A8485_ = new_A8447_ & new_A8484_;
  assign new_A8484_ = new_A8503_ | new_A8502_;
  assign new_A8483_ = ~new_A8447_ & new_A8482_;
  assign new_A8482_ = new_A8505_ | new_A8504_;
  assign new_A8481_ = new_A8447_ | new_A8480_;
  assign new_A8480_ = new_A8501_ | new_A8500_;
  assign new_A8479_ = ~new_A8459_ & ~new_A8469_;
  assign new_A8478_ = new_A8459_ & new_A8469_;
  assign new_A8477_ = ~new_A8459_ | new_A8469_;
  assign new_A8476_ = new_A8443_ & ~new_A8444_;
  assign new_A8475_ = ~new_A8443_ & new_A8444_;
  assign new_A8474_ = new_A8496_ & ~new_A8497_;
  assign new_A8473_ = ~new_A8496_ & new_A8497_;
  assign new_A8472_ = ~new_A8495_ | ~new_A8494_;
  assign new_A8471_ = new_A8487_ | new_A8486_;
  assign new_A8470_ = new_A8493_ | new_A8492_;
  assign new_A8469_ = new_A8483_ | new_A8485_;
  assign new_A8468_ = ~new_A8490_ | ~new_A8491_;
  assign new_A8467_ = new_A8443_ & ~new_A8444_;
  assign new_A8466_ = new_A8457_ & ~new_A8469_;
  assign new_A8465_ = ~new_A8457_ & new_A8469_;
  assign new_A8464_ = ~new_A8455_ & new_A8481_;
  assign new_A8463_ = new_A8479_ | new_A8478_;
  assign new_A8462_ = new_A8476_ | new_A8475_;
  assign new_A8461_ = new_A8444_ | new_A8477_;
  assign new_A8460_ = new_A8469_ & new_A8472_;
  assign new_A8459_ = new_A8474_ | new_A8473_;
  assign new_A8458_ = new_A8469_ & new_A8468_;
  assign new_A8457_ = new_A8471_ & new_A8470_;
  assign new_A8456_ = new_A8466_ | new_A8465_;
  assign new_A8455_ = new_A8444_ | new_A8467_;
  assign A8454 = new_A8455_ | new_A8464_;
  assign A8453 = new_A8462_ & new_A8463_;
  assign A8452 = new_A8462_ & new_A8461_;
  assign A8451 = new_A8460_ | new_A8459_;
  assign A8450 = new_A8458_ | new_A8457_;
  assign A8449 = new_A8456_ & new_A8455_;
  assign new_A8448_ = new_C5268_;
  assign new_A8447_ = new_C5201_;
  assign new_A8446_ = new_C5134_;
  assign new_A8445_ = new_C5067_;
  assign new_A8444_ = new_C5000_;
  assign new_A8443_ = new_C4933_;
  assign new_A8442_ = ~new_A8381_ & new_A8395_;
  assign new_A8441_ = new_A8381_ & ~new_A8395_;
  assign new_A8440_ = new_A8381_ & ~new_A8395_;
  assign new_A8439_ = ~new_A8381_ & ~new_A8395_;
  assign new_A8438_ = new_A8381_ & new_A8395_;
  assign new_A8437_ = new_A8441_ | new_A8442_;
  assign new_A8436_ = ~new_A8381_ & new_A8395_;
  assign new_A8435_ = new_A8439_ | new_A8440_;
  assign new_A8434_ = ~new_A8410_ & ~new_A8430_;
  assign new_A8433_ = new_A8410_ & new_A8430_;
  assign new_A8432_ = ~new_A8377_ | ~new_A8402_;
  assign new_A8431_ = new_A8395_ & new_A8432_;
  assign new_A8430_ = new_A8378_ | new_A8379_;
  assign new_A8429_ = new_A8378_ | new_A8395_;
  assign new_A8428_ = ~new_A8395_ & ~new_A8431_;
  assign new_A8427_ = new_A8395_ | new_A8432_;
  assign new_A8426_ = new_A8378_ & ~new_A8379_;
  assign new_A8425_ = ~new_A8378_ & new_A8379_;
  assign new_A8424_ = new_A8388_ | new_A8421_;
  assign new_A8423_ = ~new_A8388_ & ~new_A8422_;
  assign new_A8422_ = new_A8388_ & new_A8421_;
  assign new_A8421_ = ~new_A8377_ | ~new_A8402_;
  assign new_A8420_ = ~new_A8378_ & new_A8388_;
  assign new_A8419_ = new_A8378_ & ~new_A8388_;
  assign new_A8418_ = new_A8380_ & new_A8417_;
  assign new_A8417_ = new_A8436_ | new_A8435_;
  assign new_A8416_ = ~new_A8380_ & new_A8415_;
  assign new_A8415_ = new_A8438_ | new_A8437_;
  assign new_A8414_ = new_A8380_ | new_A8413_;
  assign new_A8413_ = new_A8434_ | new_A8433_;
  assign new_A8412_ = ~new_A8392_ & ~new_A8402_;
  assign new_A8411_ = new_A8392_ & new_A8402_;
  assign new_A8410_ = ~new_A8392_ | new_A8402_;
  assign new_A8409_ = new_A8376_ & ~new_A8377_;
  assign new_A8408_ = ~new_A8376_ & new_A8377_;
  assign new_A8407_ = new_A8429_ & ~new_A8430_;
  assign new_A8406_ = ~new_A8429_ & new_A8430_;
  assign new_A8405_ = ~new_A8428_ | ~new_A8427_;
  assign new_A8404_ = new_A8420_ | new_A8419_;
  assign new_A8403_ = new_A8426_ | new_A8425_;
  assign new_A8402_ = new_A8416_ | new_A8418_;
  assign new_A8401_ = ~new_A8423_ | ~new_A8424_;
  assign new_A8400_ = new_A8376_ & ~new_A8377_;
  assign new_A8399_ = new_A8390_ & ~new_A8402_;
  assign new_A8398_ = ~new_A8390_ & new_A8402_;
  assign new_A8397_ = ~new_A8388_ & new_A8414_;
  assign new_A8396_ = new_A8412_ | new_A8411_;
  assign new_A8395_ = new_A8409_ | new_A8408_;
  assign new_A8394_ = new_A8377_ | new_A8410_;
  assign new_A8393_ = new_A8402_ & new_A8405_;
  assign new_A8392_ = new_A8407_ | new_A8406_;
  assign new_A8391_ = new_A8402_ & new_A8401_;
  assign new_A8390_ = new_A8404_ & new_A8403_;
  assign new_A8389_ = new_A8399_ | new_A8398_;
  assign new_A8388_ = new_A8377_ | new_A8400_;
  assign A8387 = new_A8388_ | new_A8397_;
  assign A8386 = new_A8395_ & new_A8396_;
  assign A8385 = new_A8395_ & new_A8394_;
  assign A8384 = new_A8393_ | new_A8392_;
  assign A8383 = new_A8391_ | new_A8390_;
  assign A8382 = new_A8389_ & new_A8388_;
  assign new_A8381_ = new_C4866_;
  assign new_A8380_ = new_C4799_;
  assign new_A8379_ = new_C4732_;
  assign new_A8378_ = new_C4665_;
  assign new_A8377_ = new_C4598_;
  assign new_A8376_ = new_C4531_;
  assign new_A8375_ = ~new_A8314_ & new_A8328_;
  assign new_A8374_ = new_A8314_ & ~new_A8328_;
  assign new_A8373_ = new_A8314_ & ~new_A8328_;
  assign new_A8372_ = ~new_A8314_ & ~new_A8328_;
  assign new_A8371_ = new_A8314_ & new_A8328_;
  assign new_A8370_ = new_A8374_ | new_A8375_;
  assign new_A8369_ = ~new_A8314_ & new_A8328_;
  assign new_A8368_ = new_A8372_ | new_A8373_;
  assign new_A8367_ = ~new_A8343_ & ~new_A8363_;
  assign new_A8366_ = new_A8343_ & new_A8363_;
  assign new_A8365_ = ~new_A8310_ | ~new_A8335_;
  assign new_A8364_ = new_A8328_ & new_A8365_;
  assign new_A8363_ = new_A8311_ | new_A8312_;
  assign new_A8362_ = new_A8311_ | new_A8328_;
  assign new_A8361_ = ~new_A8328_ & ~new_A8364_;
  assign new_A8360_ = new_A8328_ | new_A8365_;
  assign new_A8359_ = new_A8311_ & ~new_A8312_;
  assign new_A8358_ = ~new_A8311_ & new_A8312_;
  assign new_A8357_ = new_A8321_ | new_A8354_;
  assign new_A8356_ = ~new_A8321_ & ~new_A8355_;
  assign new_A8355_ = new_A8321_ & new_A8354_;
  assign new_A8354_ = ~new_A8310_ | ~new_A8335_;
  assign new_A8353_ = ~new_A8311_ & new_A8321_;
  assign new_A8352_ = new_A8311_ & ~new_A8321_;
  assign new_A8351_ = new_A8313_ & new_A8350_;
  assign new_A8350_ = new_A8369_ | new_A8368_;
  assign new_A8349_ = ~new_A8313_ & new_A8348_;
  assign new_A8348_ = new_A8371_ | new_A8370_;
  assign new_A8347_ = new_A8313_ | new_A8346_;
  assign new_A8346_ = new_A8367_ | new_A8366_;
  assign new_A8345_ = ~new_A8325_ & ~new_A8335_;
  assign new_A8344_ = new_A8325_ & new_A8335_;
  assign new_A8343_ = ~new_A8325_ | new_A8335_;
  assign new_A8342_ = new_A8309_ & ~new_A8310_;
  assign new_A8341_ = ~new_A8309_ & new_A8310_;
  assign new_A8340_ = new_A8362_ & ~new_A8363_;
  assign new_A8339_ = ~new_A8362_ & new_A8363_;
  assign new_A8338_ = ~new_A8361_ | ~new_A8360_;
  assign new_A8337_ = new_A8353_ | new_A8352_;
  assign new_A8336_ = new_A8359_ | new_A8358_;
  assign new_A8335_ = new_A8349_ | new_A8351_;
  assign new_A8334_ = ~new_A8356_ | ~new_A8357_;
  assign new_A8333_ = new_A8309_ & ~new_A8310_;
  assign new_A8332_ = new_A8323_ & ~new_A8335_;
  assign new_A8331_ = ~new_A8323_ & new_A8335_;
  assign new_A8330_ = ~new_A8321_ & new_A8347_;
  assign new_A8329_ = new_A8345_ | new_A8344_;
  assign new_A8328_ = new_A8342_ | new_A8341_;
  assign new_A8327_ = new_A8310_ | new_A8343_;
  assign new_A8326_ = new_A8335_ & new_A8338_;
  assign new_A8325_ = new_A8340_ | new_A8339_;
  assign new_A8324_ = new_A8335_ & new_A8334_;
  assign new_A8323_ = new_A8337_ & new_A8336_;
  assign new_A8322_ = new_A8332_ | new_A8331_;
  assign new_A8321_ = new_A8310_ | new_A8333_;
  assign A8320 = new_A8321_ | new_A8330_;
  assign A8319 = new_A8328_ & new_A8329_;
  assign A8318 = new_A8328_ & new_A8327_;
  assign A8317 = new_A8326_ | new_A8325_;
  assign A8316 = new_A8324_ | new_A8323_;
  assign A8315 = new_A8322_ & new_A8321_;
  assign new_A8314_ = new_C4464_;
  assign new_A8313_ = new_C4397_;
  assign new_A8312_ = new_C4330_;
  assign new_A8311_ = new_C4263_;
  assign new_A8310_ = new_C4196_;
  assign new_A8309_ = new_C4129_;
  assign new_A8308_ = ~new_A8247_ & new_A8261_;
  assign new_A8307_ = new_A8247_ & ~new_A8261_;
  assign new_A8306_ = new_A8247_ & ~new_A8261_;
  assign new_A8305_ = ~new_A8247_ & ~new_A8261_;
  assign new_A8304_ = new_A8247_ & new_A8261_;
  assign new_A8303_ = new_A8307_ | new_A8308_;
  assign new_A8302_ = ~new_A8247_ & new_A8261_;
  assign new_A8301_ = new_A8305_ | new_A8306_;
  assign new_A8300_ = ~new_A8276_ & ~new_A8296_;
  assign new_A8299_ = new_A8276_ & new_A8296_;
  assign new_A8298_ = ~new_A8243_ | ~new_A8268_;
  assign new_A8297_ = new_A8261_ & new_A8298_;
  assign new_A8296_ = new_A8244_ | new_A8245_;
  assign new_A8295_ = new_A8244_ | new_A8261_;
  assign new_A8294_ = ~new_A8261_ & ~new_A8297_;
  assign new_A8293_ = new_A8261_ | new_A8298_;
  assign new_A8292_ = new_A8244_ & ~new_A8245_;
  assign new_A8291_ = ~new_A8244_ & new_A8245_;
  assign new_A8290_ = new_A8254_ | new_A8287_;
  assign new_A8289_ = ~new_A8254_ & ~new_A8288_;
  assign new_A8288_ = new_A8254_ & new_A8287_;
  assign new_A8287_ = ~new_A8243_ | ~new_A8268_;
  assign new_A8286_ = ~new_A8244_ & new_A8254_;
  assign new_A8285_ = new_A8244_ & ~new_A8254_;
  assign new_A8284_ = new_A8246_ & new_A8283_;
  assign new_A8283_ = new_A8302_ | new_A8301_;
  assign new_A8282_ = ~new_A8246_ & new_A8281_;
  assign new_A8281_ = new_A8304_ | new_A8303_;
  assign new_A8280_ = new_A8246_ | new_A8279_;
  assign new_A8279_ = new_A8300_ | new_A8299_;
  assign new_A8278_ = ~new_A8258_ & ~new_A8268_;
  assign new_A8277_ = new_A8258_ & new_A8268_;
  assign new_A8276_ = ~new_A8258_ | new_A8268_;
  assign new_A8275_ = new_A8242_ & ~new_A8243_;
  assign new_A8274_ = ~new_A8242_ & new_A8243_;
  assign new_A8273_ = new_A8295_ & ~new_A8296_;
  assign new_A8272_ = ~new_A8295_ & new_A8296_;
  assign new_A8271_ = ~new_A8294_ | ~new_A8293_;
  assign new_A8270_ = new_A8286_ | new_A8285_;
  assign new_A8269_ = new_A8292_ | new_A8291_;
  assign new_A8268_ = new_A8282_ | new_A8284_;
  assign new_A8267_ = ~new_A8289_ | ~new_A8290_;
  assign new_A8266_ = new_A8242_ & ~new_A8243_;
  assign new_A8265_ = new_A8256_ & ~new_A8268_;
  assign new_A8264_ = ~new_A8256_ & new_A8268_;
  assign new_A8263_ = ~new_A8254_ & new_A8280_;
  assign new_A8262_ = new_A8278_ | new_A8277_;
  assign new_A8261_ = new_A8275_ | new_A8274_;
  assign new_A8260_ = new_A8243_ | new_A8276_;
  assign new_A8259_ = new_A8268_ & new_A8271_;
  assign new_A8258_ = new_A8273_ | new_A8272_;
  assign new_A8257_ = new_A8268_ & new_A8267_;
  assign new_A8256_ = new_A8270_ & new_A8269_;
  assign new_A8255_ = new_A8265_ | new_A8264_;
  assign new_A8254_ = new_A8243_ | new_A8266_;
  assign A8253 = new_A8254_ | new_A8263_;
  assign A8252 = new_A8261_ & new_A8262_;
  assign A8251 = new_A8261_ & new_A8260_;
  assign A8250 = new_A8259_ | new_A8258_;
  assign A8249 = new_A8257_ | new_A8256_;
  assign A8248 = new_A8255_ & new_A8254_;
  assign new_A8247_ = new_C4062_;
  assign new_A8246_ = new_C3995_;
  assign new_A8245_ = new_C3928_;
  assign new_A8244_ = new_C3861_;
  assign new_A8243_ = new_C3794_;
  assign new_A8242_ = new_C3727_;
  assign new_A8241_ = ~new_A8180_ & new_A8194_;
  assign new_A8240_ = new_A8180_ & ~new_A8194_;
  assign new_A8239_ = new_A8180_ & ~new_A8194_;
  assign new_A8238_ = ~new_A8180_ & ~new_A8194_;
  assign new_A8237_ = new_A8180_ & new_A8194_;
  assign new_A8236_ = new_A8240_ | new_A8241_;
  assign new_A8235_ = ~new_A8180_ & new_A8194_;
  assign new_A8234_ = new_A8238_ | new_A8239_;
  assign new_A8233_ = ~new_A8209_ & ~new_A8229_;
  assign new_A8232_ = new_A8209_ & new_A8229_;
  assign new_A8231_ = ~new_A8176_ | ~new_A8201_;
  assign new_A8230_ = new_A8194_ & new_A8231_;
  assign new_A8229_ = new_A8177_ | new_A8178_;
  assign new_A8228_ = new_A8177_ | new_A8194_;
  assign new_A8227_ = ~new_A8194_ & ~new_A8230_;
  assign new_A8226_ = new_A8194_ | new_A8231_;
  assign new_A8225_ = new_A8177_ & ~new_A8178_;
  assign new_A8224_ = ~new_A8177_ & new_A8178_;
  assign new_A8223_ = new_A8187_ | new_A8220_;
  assign new_A8222_ = ~new_A8187_ & ~new_A8221_;
  assign new_A8221_ = new_A8187_ & new_A8220_;
  assign new_A8220_ = ~new_A8176_ | ~new_A8201_;
  assign new_A8219_ = ~new_A8177_ & new_A8187_;
  assign new_A8218_ = new_A8177_ & ~new_A8187_;
  assign new_A8217_ = new_A8179_ & new_A8216_;
  assign new_A8216_ = new_A8235_ | new_A8234_;
  assign new_A8215_ = ~new_A8179_ & new_A8214_;
  assign new_A8214_ = new_A8237_ | new_A8236_;
  assign new_A8213_ = new_A8179_ | new_A8212_;
  assign new_A8212_ = new_A8233_ | new_A8232_;
  assign new_A8211_ = ~new_A8191_ & ~new_A8201_;
  assign new_A8210_ = new_A8191_ & new_A8201_;
  assign new_A8209_ = ~new_A8191_ | new_A8201_;
  assign new_A8208_ = new_A8175_ & ~new_A8176_;
  assign new_A8207_ = ~new_A8175_ & new_A8176_;
  assign new_A8206_ = new_A8228_ & ~new_A8229_;
  assign new_A8205_ = ~new_A8228_ & new_A8229_;
  assign new_A8204_ = ~new_A8227_ | ~new_A8226_;
  assign new_A8203_ = new_A8219_ | new_A8218_;
  assign new_A8202_ = new_A8225_ | new_A8224_;
  assign new_A8201_ = new_A8215_ | new_A8217_;
  assign new_A8200_ = ~new_A8222_ | ~new_A8223_;
  assign new_A8199_ = new_A8175_ & ~new_A8176_;
  assign new_A8198_ = new_A8189_ & ~new_A8201_;
  assign new_A8197_ = ~new_A8189_ & new_A8201_;
  assign new_A8196_ = ~new_A8187_ & new_A8213_;
  assign new_A8195_ = new_A8211_ | new_A8210_;
  assign new_A8194_ = new_A8208_ | new_A8207_;
  assign new_A8193_ = new_A8176_ | new_A8209_;
  assign new_A8192_ = new_A8201_ & new_A8204_;
  assign new_A8191_ = new_A8206_ | new_A8205_;
  assign new_A8190_ = new_A8201_ & new_A8200_;
  assign new_A8189_ = new_A8203_ & new_A8202_;
  assign new_A8188_ = new_A8198_ | new_A8197_;
  assign new_A8187_ = new_A8176_ | new_A8199_;
  assign A8186 = new_A8187_ | new_A8196_;
  assign A8185 = new_A8194_ & new_A8195_;
  assign A8184 = new_A8194_ & new_A8193_;
  assign A8183 = new_A8192_ | new_A8191_;
  assign A8182 = new_A8190_ | new_A8189_;
  assign A8181 = new_A8188_ & new_A8187_;
  assign new_A8180_ = new_C3660_;
  assign new_A8179_ = new_C3593_;
  assign new_A8178_ = new_C3526_;
  assign new_A8177_ = new_C3459_;
  assign new_A8176_ = new_C3392_;
  assign new_A8175_ = new_C3325_;
  assign new_A8174_ = ~new_A8113_ & new_A8127_;
  assign new_A8173_ = new_A8113_ & ~new_A8127_;
  assign new_A8172_ = new_A8113_ & ~new_A8127_;
  assign new_A8171_ = ~new_A8113_ & ~new_A8127_;
  assign new_A8170_ = new_A8113_ & new_A8127_;
  assign new_A8169_ = new_A8173_ | new_A8174_;
  assign new_A8168_ = ~new_A8113_ & new_A8127_;
  assign new_A8167_ = new_A8171_ | new_A8172_;
  assign new_A8166_ = ~new_A8142_ & ~new_A8162_;
  assign new_A8165_ = new_A8142_ & new_A8162_;
  assign new_A8164_ = ~new_A8109_ | ~new_A8134_;
  assign new_A8163_ = new_A8127_ & new_A8164_;
  assign new_A8162_ = new_A8110_ | new_A8111_;
  assign new_A8161_ = new_A8110_ | new_A8127_;
  assign new_A8160_ = ~new_A8127_ & ~new_A8163_;
  assign new_A8159_ = new_A8127_ | new_A8164_;
  assign new_A8158_ = new_A8110_ & ~new_A8111_;
  assign new_A8157_ = ~new_A8110_ & new_A8111_;
  assign new_A8156_ = new_A8120_ | new_A8153_;
  assign new_A8155_ = ~new_A8120_ & ~new_A8154_;
  assign new_A8154_ = new_A8120_ & new_A8153_;
  assign new_A8153_ = ~new_A8109_ | ~new_A8134_;
  assign new_A8152_ = ~new_A8110_ & new_A8120_;
  assign new_A8151_ = new_A8110_ & ~new_A8120_;
  assign new_A8150_ = new_A8112_ & new_A8149_;
  assign new_A8149_ = new_A8168_ | new_A8167_;
  assign new_A8148_ = ~new_A8112_ & new_A8147_;
  assign new_A8147_ = new_A8170_ | new_A8169_;
  assign new_A8146_ = new_A8112_ | new_A8145_;
  assign new_A8145_ = new_A8166_ | new_A8165_;
  assign new_A8144_ = ~new_A8124_ & ~new_A8134_;
  assign new_A8143_ = new_A8124_ & new_A8134_;
  assign new_A8142_ = ~new_A8124_ | new_A8134_;
  assign new_A8141_ = new_A8108_ & ~new_A8109_;
  assign new_A8140_ = ~new_A8108_ & new_A8109_;
  assign new_A8139_ = new_A8161_ & ~new_A8162_;
  assign new_A8138_ = ~new_A8161_ & new_A8162_;
  assign new_A8137_ = ~new_A8160_ | ~new_A8159_;
  assign new_A8136_ = new_A8152_ | new_A8151_;
  assign new_A8135_ = new_A8158_ | new_A8157_;
  assign new_A8134_ = new_A8148_ | new_A8150_;
  assign new_A8133_ = ~new_A8155_ | ~new_A8156_;
  assign new_A8132_ = new_A8108_ & ~new_A8109_;
  assign new_A8131_ = new_A8122_ & ~new_A8134_;
  assign new_A8130_ = ~new_A8122_ & new_A8134_;
  assign new_A8129_ = ~new_A8120_ & new_A8146_;
  assign new_A8128_ = new_A8144_ | new_A8143_;
  assign new_A8127_ = new_A8141_ | new_A8140_;
  assign new_A8126_ = new_A8109_ | new_A8142_;
  assign new_A8125_ = new_A8134_ & new_A8137_;
  assign new_A8124_ = new_A8139_ | new_A8138_;
  assign new_A8123_ = new_A8134_ & new_A8133_;
  assign new_A8122_ = new_A8136_ & new_A8135_;
  assign new_A8121_ = new_A8131_ | new_A8130_;
  assign new_A8120_ = new_A8109_ | new_A8132_;
  assign A8119 = new_A8120_ | new_A8129_;
  assign A8118 = new_A8127_ & new_A8128_;
  assign A8117 = new_A8127_ & new_A8126_;
  assign A8116 = new_A8125_ | new_A8124_;
  assign A8115 = new_A8123_ | new_A8122_;
  assign A8114 = new_A8121_ & new_A8120_;
  assign new_A8113_ = new_C3258_;
  assign new_A8112_ = new_C3191_;
  assign new_A8111_ = new_C3124_;
  assign new_A8110_ = new_C3057_;
  assign new_A8109_ = new_C2990_;
  assign new_A8108_ = new_C2923_;
  assign new_A8041_ = new_C2856_;
  assign new_A8042_ = new_C2789_;
  assign new_A8043_ = new_C2722_;
  assign new_A8044_ = new_C2655_;
  assign new_A8045_ = new_C2588_;
  assign new_A8046_ = new_C2526_;
  assign A8047 = new_A8054_ & new_A8053_;
  assign A8048 = new_A8056_ | new_A8055_;
  assign A8049 = new_A8058_ | new_A8057_;
  assign A8050 = new_A8060_ & new_A8059_;
  assign A8051 = new_A8060_ & new_A8061_;
  assign A8052 = new_A8053_ | new_A8062_;
  assign new_A8053_ = new_A8042_ | new_A8065_;
  assign new_A8054_ = new_A8064_ | new_A8063_;
  assign new_A8055_ = new_A8069_ & new_A8068_;
  assign new_A8056_ = new_A8067_ & new_A8066_;
  assign new_A8057_ = new_A8072_ | new_A8071_;
  assign new_A8058_ = new_A8067_ & new_A8070_;
  assign new_A8059_ = new_A8042_ | new_A8075_;
  assign new_A8060_ = new_A8074_ | new_A8073_;
  assign new_A8061_ = new_A8077_ | new_A8076_;
  assign new_A8062_ = ~new_A8053_ & new_A8079_;
  assign new_A8063_ = ~new_A8055_ & new_A8067_;
  assign new_A8064_ = new_A8055_ & ~new_A8067_;
  assign new_A8065_ = new_A8041_ & ~new_A8042_;
  assign new_A8066_ = ~new_A8088_ | ~new_A8089_;
  assign new_A8067_ = new_A8081_ | new_A8083_;
  assign new_A8068_ = new_A8091_ | new_A8090_;
  assign new_A8069_ = new_A8085_ | new_A8084_;
  assign new_A8070_ = ~new_A8093_ | ~new_A8092_;
  assign new_A8071_ = ~new_A8094_ & new_A8095_;
  assign new_A8072_ = new_A8094_ & ~new_A8095_;
  assign new_A8073_ = ~new_A8041_ & new_A8042_;
  assign new_A8074_ = new_A8041_ & ~new_A8042_;
  assign new_A8075_ = ~new_A8057_ | new_A8067_;
  assign new_A8076_ = new_A8057_ & new_A8067_;
  assign new_A8077_ = ~new_A8057_ & ~new_A8067_;
  assign new_A8078_ = new_A8099_ | new_A8098_;
  assign new_A8079_ = new_A8045_ | new_A8078_;
  assign new_A8080_ = new_A8103_ | new_A8102_;
  assign new_A8081_ = ~new_A8045_ & new_A8080_;
  assign new_A8082_ = new_A8101_ | new_A8100_;
  assign new_A8083_ = new_A8045_ & new_A8082_;
  assign new_A8084_ = new_A8043_ & ~new_A8053_;
  assign new_A8085_ = ~new_A8043_ & new_A8053_;
  assign new_A8086_ = ~new_A8042_ | ~new_A8067_;
  assign new_A8087_ = new_A8053_ & new_A8086_;
  assign new_A8088_ = ~new_A8053_ & ~new_A8087_;
  assign new_A8089_ = new_A8053_ | new_A8086_;
  assign new_A8090_ = ~new_A8043_ & new_A8044_;
  assign new_A8091_ = new_A8043_ & ~new_A8044_;
  assign new_A8092_ = new_A8060_ | new_A8097_;
  assign new_A8093_ = ~new_A8060_ & ~new_A8096_;
  assign new_A8094_ = new_A8043_ | new_A8060_;
  assign new_A8095_ = new_A8043_ | new_A8044_;
  assign new_A8096_ = new_A8060_ & new_A8097_;
  assign new_A8097_ = ~new_A8042_ | ~new_A8067_;
  assign new_A8098_ = new_A8075_ & new_A8095_;
  assign new_A8099_ = ~new_A8075_ & ~new_A8095_;
  assign new_A8100_ = new_A8104_ | new_A8105_;
  assign new_A8101_ = ~new_A8046_ & new_A8060_;
  assign new_A8102_ = new_A8106_ | new_A8107_;
  assign new_A8103_ = new_A8046_ & new_A8060_;
  assign new_A8104_ = ~new_A8046_ & ~new_A8060_;
  assign new_A8105_ = new_A8046_ & ~new_A8060_;
  assign new_A8106_ = new_A8046_ & ~new_A8060_;
  assign new_A8107_ = ~new_A8046_ & new_A8060_;
endmodule


