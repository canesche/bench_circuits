// Benchmark "pci_bridge32" written by ABC on Thu Oct  8 22:04:25 2020

module pci_bridge32 ( clock, 
    wb_clk_i, wb_rst_i, wb_int_i, wbs_cyc_i, wbs_stb_i, wbs_we_i,
    wbm_ack_i, wbm_rty_i, wbm_err_i, pci_clk_i, pci_rst_i, pci_inta_i,
    pci_gnt_i, pci_frame_i, pci_irdy_i, pci_idsel_i, pci_devsel_i,
    pci_trdy_i, pci_stop_i, pci_par_i, pci_perr_i, \wbs_adr_i[0] ,
    \wbs_adr_i[1] , \wbs_adr_i[2] , \wbs_adr_i[3] , \wbs_adr_i[4] ,
    \wbs_adr_i[5] , \wbs_adr_i[6] , \wbs_adr_i[7] , \wbs_adr_i[8] ,
    \wbs_adr_i[9] , \wbs_adr_i[10] , \wbs_adr_i[11] , \wbs_adr_i[12] ,
    \wbs_adr_i[13] , \wbs_adr_i[14] , \wbs_adr_i[15] , \wbs_adr_i[16] ,
    \wbs_adr_i[17] , \wbs_adr_i[18] , \wbs_adr_i[19] , \wbs_adr_i[20] ,
    \wbs_adr_i[21] , \wbs_adr_i[22] , \wbs_adr_i[23] , \wbs_adr_i[24] ,
    \wbs_adr_i[25] , \wbs_adr_i[26] , \wbs_adr_i[27] , \wbs_adr_i[28] ,
    \wbs_adr_i[29] , \wbs_adr_i[30] , \wbs_adr_i[31] , \wbs_dat_i[0] ,
    \wbs_dat_i[1] , \wbs_dat_i[2] , \wbs_dat_i[3] , \wbs_dat_i[4] ,
    \wbs_dat_i[5] , \wbs_dat_i[6] , \wbs_dat_i[7] , \wbs_dat_i[8] ,
    \wbs_dat_i[9] , \wbs_dat_i[10] , \wbs_dat_i[11] , \wbs_dat_i[12] ,
    \wbs_dat_i[13] , \wbs_dat_i[14] , \wbs_dat_i[15] , \wbs_dat_i[16] ,
    \wbs_dat_i[17] , \wbs_dat_i[18] , \wbs_dat_i[19] , \wbs_dat_i[20] ,
    \wbs_dat_i[21] , \wbs_dat_i[22] , \wbs_dat_i[23] , \wbs_dat_i[24] ,
    \wbs_dat_i[25] , \wbs_dat_i[26] , \wbs_dat_i[27] , \wbs_dat_i[28] ,
    \wbs_dat_i[29] , \wbs_dat_i[30] , \wbs_dat_i[31] , \wbm_dat_i[0] ,
    \wbm_dat_i[1] , \wbm_dat_i[2] , \wbm_dat_i[3] , \wbm_dat_i[4] ,
    \wbm_dat_i[5] , \wbm_dat_i[6] , \wbm_dat_i[7] , \wbm_dat_i[8] ,
    \wbm_dat_i[9] , \wbm_dat_i[10] , \wbm_dat_i[11] , \wbm_dat_i[12] ,
    \wbm_dat_i[13] , \wbm_dat_i[14] , \wbm_dat_i[15] , \wbm_dat_i[16] ,
    \wbm_dat_i[17] , \wbm_dat_i[18] , \wbm_dat_i[19] , \wbm_dat_i[20] ,
    \wbm_dat_i[21] , \wbm_dat_i[22] , \wbm_dat_i[23] , \wbm_dat_i[24] ,
    \wbm_dat_i[25] , \wbm_dat_i[26] , \wbm_dat_i[27] , \wbm_dat_i[28] ,
    \wbm_dat_i[29] , \wbm_dat_i[30] , \wbm_dat_i[31] , \pci_ad_i[0] ,
    \pci_ad_i[1] , \pci_ad_i[2] , \pci_ad_i[3] , \pci_ad_i[4] ,
    \pci_ad_i[5] , \pci_ad_i[6] , \pci_ad_i[7] , \pci_ad_i[8] ,
    \pci_ad_i[9] , \pci_ad_i[10] , \pci_ad_i[11] , \pci_ad_i[12] ,
    \pci_ad_i[13] , \pci_ad_i[14] , \pci_ad_i[15] , \pci_ad_i[16] ,
    \pci_ad_i[17] , \pci_ad_i[18] , \pci_ad_i[19] , \pci_ad_i[20] ,
    \pci_ad_i[21] , \pci_ad_i[22] , \pci_ad_i[23] , \pci_ad_i[24] ,
    \pci_ad_i[25] , \pci_ad_i[26] , \pci_ad_i[27] , \pci_ad_i[28] ,
    \pci_ad_i[29] , \pci_ad_i[30] , \pci_ad_i[31] , \wbs_sel_i[0] ,
    \wbs_sel_i[1] , \wbs_sel_i[2] , \wbs_sel_i[3] , \pci_cbe_i[0] ,
    \pci_cbe_i[1] , \pci_cbe_i[2] , \pci_cbe_i[3] , \wbs_cti_i[0] ,
    \wbs_cti_i[1] , \wbs_cti_i[2] , \wbs_bte_i[0] , \wbs_bte_i[1] ,
    wb_rst_o, wb_int_o, wbs_ack_o, wbs_rty_o, wbs_err_o, wbm_cyc_o,
    wbm_stb_o, wbm_we_o, pci_rst_o, pci_inta_o, pci_rst_oe_o,
    pci_inta_oe_o, pci_req_o, pci_req_oe_o, pci_frame_o, pci_frame_oe_o,
    pci_irdy_oe_o, pci_devsel_oe_o, pci_trdy_oe_o, pci_stop_oe_o,
    pci_irdy_o, pci_devsel_o, pci_trdy_o, pci_stop_o, pci_par_o,
    pci_par_oe_o, pci_perr_o, pci_perr_oe_o, pci_serr_o, pci_serr_oe_o,
    \wbs_dat_o[0] , \wbs_dat_o[1] , \wbs_dat_o[2] , \wbs_dat_o[3] ,
    \wbs_dat_o[4] , \wbs_dat_o[5] , \wbs_dat_o[6] , \wbs_dat_o[7] ,
    \wbs_dat_o[8] , \wbs_dat_o[9] , \wbs_dat_o[10] , \wbs_dat_o[11] ,
    \wbs_dat_o[12] , \wbs_dat_o[13] , \wbs_dat_o[14] , \wbs_dat_o[15] ,
    \wbs_dat_o[16] , \wbs_dat_o[17] , \wbs_dat_o[18] , \wbs_dat_o[19] ,
    \wbs_dat_o[20] , \wbs_dat_o[21] , \wbs_dat_o[22] , \wbs_dat_o[23] ,
    \wbs_dat_o[24] , \wbs_dat_o[25] , \wbs_dat_o[26] , \wbs_dat_o[27] ,
    \wbs_dat_o[28] , \wbs_dat_o[29] , \wbs_dat_o[30] , \wbs_dat_o[31] ,
    \wbm_adr_o[0] , \wbm_adr_o[1] , \wbm_adr_o[2] , \wbm_adr_o[3] ,
    \wbm_adr_o[4] , \wbm_adr_o[5] , \wbm_adr_o[6] , \wbm_adr_o[7] ,
    \wbm_adr_o[8] , \wbm_adr_o[9] , \wbm_adr_o[10] , \wbm_adr_o[11] ,
    \wbm_adr_o[12] , \wbm_adr_o[13] , \wbm_adr_o[14] , \wbm_adr_o[15] ,
    \wbm_adr_o[16] , \wbm_adr_o[17] , \wbm_adr_o[18] , \wbm_adr_o[19] ,
    \wbm_adr_o[20] , \wbm_adr_o[21] , \wbm_adr_o[22] , \wbm_adr_o[23] ,
    \wbm_adr_o[24] , \wbm_adr_o[25] , \wbm_adr_o[26] , \wbm_adr_o[27] ,
    \wbm_adr_o[28] , \wbm_adr_o[29] , \wbm_adr_o[30] , \wbm_adr_o[31] ,
    \wbm_dat_o[0] , \wbm_dat_o[1] , \wbm_dat_o[2] , \wbm_dat_o[3] ,
    \wbm_dat_o[4] , \wbm_dat_o[5] , \wbm_dat_o[6] , \wbm_dat_o[7] ,
    \wbm_dat_o[8] , \wbm_dat_o[9] , \wbm_dat_o[10] , \wbm_dat_o[11] ,
    \wbm_dat_o[12] , \wbm_dat_o[13] , \wbm_dat_o[14] , \wbm_dat_o[15] ,
    \wbm_dat_o[16] , \wbm_dat_o[17] , \wbm_dat_o[18] , \wbm_dat_o[19] ,
    \wbm_dat_o[20] , \wbm_dat_o[21] , \wbm_dat_o[22] , \wbm_dat_o[23] ,
    \wbm_dat_o[24] , \wbm_dat_o[25] , \wbm_dat_o[26] , \wbm_dat_o[27] ,
    \wbm_dat_o[28] , \wbm_dat_o[29] , \wbm_dat_o[30] , \wbm_dat_o[31] ,
    \pci_ad_oe_o[0] , \pci_ad_oe_o[1] , \pci_ad_oe_o[2] , \pci_ad_oe_o[3] ,
    \pci_ad_oe_o[4] , \pci_ad_oe_o[5] , \pci_ad_oe_o[6] , \pci_ad_oe_o[7] ,
    \pci_ad_oe_o[8] , \pci_ad_oe_o[9] , \pci_ad_oe_o[10] ,
    \pci_ad_oe_o[11] , \pci_ad_oe_o[12] , \pci_ad_oe_o[13] ,
    \pci_ad_oe_o[14] , \pci_ad_oe_o[15] , \pci_ad_oe_o[16] ,
    \pci_ad_oe_o[17] , \pci_ad_oe_o[18] , \pci_ad_oe_o[19] ,
    \pci_ad_oe_o[20] , \pci_ad_oe_o[21] , \pci_ad_oe_o[22] ,
    \pci_ad_oe_o[23] , \pci_ad_oe_o[24] , \pci_ad_oe_o[25] ,
    \pci_ad_oe_o[26] , \pci_ad_oe_o[27] , \pci_ad_oe_o[28] ,
    \pci_ad_oe_o[29] , \pci_ad_oe_o[30] , \pci_ad_oe_o[31] , \pci_ad_o[0] ,
    \pci_ad_o[1] , \pci_ad_o[2] , \pci_ad_o[3] , \pci_ad_o[4] ,
    \pci_ad_o[5] , \pci_ad_o[6] , \pci_ad_o[7] , \pci_ad_o[8] ,
    \pci_ad_o[9] , \pci_ad_o[10] , \pci_ad_o[11] , \pci_ad_o[12] ,
    \pci_ad_o[13] , \pci_ad_o[14] , \pci_ad_o[15] , \pci_ad_o[16] ,
    \pci_ad_o[17] , \pci_ad_o[18] , \pci_ad_o[19] , \pci_ad_o[20] ,
    \pci_ad_o[21] , \pci_ad_o[22] , \pci_ad_o[23] , \pci_ad_o[24] ,
    \pci_ad_o[25] , \pci_ad_o[26] , \pci_ad_o[27] , \pci_ad_o[28] ,
    \pci_ad_o[29] , \pci_ad_o[30] , \pci_ad_o[31] , \wbm_sel_o[0] ,
    \wbm_sel_o[1] , \wbm_sel_o[2] , \wbm_sel_o[3] , \pci_cbe_oe_o[0] ,
    \pci_cbe_oe_o[1] , \pci_cbe_oe_o[2] , \pci_cbe_oe_o[3] ,
    \pci_cbe_o[0] , \pci_cbe_o[1] , \pci_cbe_o[2] , \pci_cbe_o[3] ,
    \wbm_cti_o[0] , \wbm_cti_o[1] , \wbm_cti_o[2] , \wbm_bte_o[0] ,
    \wbm_bte_o[1]   );
  input  clock;
  input  wb_clk_i, wb_rst_i, wb_int_i, wbs_cyc_i, wbs_stb_i, wbs_we_i,
    wbm_ack_i, wbm_rty_i, wbm_err_i, pci_clk_i, pci_rst_i, pci_inta_i,
    pci_gnt_i, pci_frame_i, pci_irdy_i, pci_idsel_i, pci_devsel_i,
    pci_trdy_i, pci_stop_i, pci_par_i, pci_perr_i, \wbs_adr_i[0] ,
    \wbs_adr_i[1] , \wbs_adr_i[2] , \wbs_adr_i[3] , \wbs_adr_i[4] ,
    \wbs_adr_i[5] , \wbs_adr_i[6] , \wbs_adr_i[7] , \wbs_adr_i[8] ,
    \wbs_adr_i[9] , \wbs_adr_i[10] , \wbs_adr_i[11] , \wbs_adr_i[12] ,
    \wbs_adr_i[13] , \wbs_adr_i[14] , \wbs_adr_i[15] , \wbs_adr_i[16] ,
    \wbs_adr_i[17] , \wbs_adr_i[18] , \wbs_adr_i[19] , \wbs_adr_i[20] ,
    \wbs_adr_i[21] , \wbs_adr_i[22] , \wbs_adr_i[23] , \wbs_adr_i[24] ,
    \wbs_adr_i[25] , \wbs_adr_i[26] , \wbs_adr_i[27] , \wbs_adr_i[28] ,
    \wbs_adr_i[29] , \wbs_adr_i[30] , \wbs_adr_i[31] , \wbs_dat_i[0] ,
    \wbs_dat_i[1] , \wbs_dat_i[2] , \wbs_dat_i[3] , \wbs_dat_i[4] ,
    \wbs_dat_i[5] , \wbs_dat_i[6] , \wbs_dat_i[7] , \wbs_dat_i[8] ,
    \wbs_dat_i[9] , \wbs_dat_i[10] , \wbs_dat_i[11] , \wbs_dat_i[12] ,
    \wbs_dat_i[13] , \wbs_dat_i[14] , \wbs_dat_i[15] , \wbs_dat_i[16] ,
    \wbs_dat_i[17] , \wbs_dat_i[18] , \wbs_dat_i[19] , \wbs_dat_i[20] ,
    \wbs_dat_i[21] , \wbs_dat_i[22] , \wbs_dat_i[23] , \wbs_dat_i[24] ,
    \wbs_dat_i[25] , \wbs_dat_i[26] , \wbs_dat_i[27] , \wbs_dat_i[28] ,
    \wbs_dat_i[29] , \wbs_dat_i[30] , \wbs_dat_i[31] , \wbm_dat_i[0] ,
    \wbm_dat_i[1] , \wbm_dat_i[2] , \wbm_dat_i[3] , \wbm_dat_i[4] ,
    \wbm_dat_i[5] , \wbm_dat_i[6] , \wbm_dat_i[7] , \wbm_dat_i[8] ,
    \wbm_dat_i[9] , \wbm_dat_i[10] , \wbm_dat_i[11] , \wbm_dat_i[12] ,
    \wbm_dat_i[13] , \wbm_dat_i[14] , \wbm_dat_i[15] , \wbm_dat_i[16] ,
    \wbm_dat_i[17] , \wbm_dat_i[18] , \wbm_dat_i[19] , \wbm_dat_i[20] ,
    \wbm_dat_i[21] , \wbm_dat_i[22] , \wbm_dat_i[23] , \wbm_dat_i[24] ,
    \wbm_dat_i[25] , \wbm_dat_i[26] , \wbm_dat_i[27] , \wbm_dat_i[28] ,
    \wbm_dat_i[29] , \wbm_dat_i[30] , \wbm_dat_i[31] , \pci_ad_i[0] ,
    \pci_ad_i[1] , \pci_ad_i[2] , \pci_ad_i[3] , \pci_ad_i[4] ,
    \pci_ad_i[5] , \pci_ad_i[6] , \pci_ad_i[7] , \pci_ad_i[8] ,
    \pci_ad_i[9] , \pci_ad_i[10] , \pci_ad_i[11] , \pci_ad_i[12] ,
    \pci_ad_i[13] , \pci_ad_i[14] , \pci_ad_i[15] , \pci_ad_i[16] ,
    \pci_ad_i[17] , \pci_ad_i[18] , \pci_ad_i[19] , \pci_ad_i[20] ,
    \pci_ad_i[21] , \pci_ad_i[22] , \pci_ad_i[23] , \pci_ad_i[24] ,
    \pci_ad_i[25] , \pci_ad_i[26] , \pci_ad_i[27] , \pci_ad_i[28] ,
    \pci_ad_i[29] , \pci_ad_i[30] , \pci_ad_i[31] , \wbs_sel_i[0] ,
    \wbs_sel_i[1] , \wbs_sel_i[2] , \wbs_sel_i[3] , \pci_cbe_i[0] ,
    \pci_cbe_i[1] , \pci_cbe_i[2] , \pci_cbe_i[3] , \wbs_cti_i[0] ,
    \wbs_cti_i[1] , \wbs_cti_i[2] , \wbs_bte_i[0] , \wbs_bte_i[1] ;
  output wb_rst_o, wb_int_o, wbs_ack_o, wbs_rty_o, wbs_err_o, wbm_cyc_o,
    wbm_stb_o, wbm_we_o, pci_rst_o, pci_inta_o, pci_rst_oe_o,
    pci_inta_oe_o, pci_req_o, pci_req_oe_o, pci_frame_o, pci_frame_oe_o,
    pci_irdy_oe_o, pci_devsel_oe_o, pci_trdy_oe_o, pci_stop_oe_o,
    pci_irdy_o, pci_devsel_o, pci_trdy_o, pci_stop_o, pci_par_o,
    pci_par_oe_o, pci_perr_o, pci_perr_oe_o, pci_serr_o, pci_serr_oe_o,
    \wbs_dat_o[0] , \wbs_dat_o[1] , \wbs_dat_o[2] , \wbs_dat_o[3] ,
    \wbs_dat_o[4] , \wbs_dat_o[5] , \wbs_dat_o[6] , \wbs_dat_o[7] ,
    \wbs_dat_o[8] , \wbs_dat_o[9] , \wbs_dat_o[10] , \wbs_dat_o[11] ,
    \wbs_dat_o[12] , \wbs_dat_o[13] , \wbs_dat_o[14] , \wbs_dat_o[15] ,
    \wbs_dat_o[16] , \wbs_dat_o[17] , \wbs_dat_o[18] , \wbs_dat_o[19] ,
    \wbs_dat_o[20] , \wbs_dat_o[21] , \wbs_dat_o[22] , \wbs_dat_o[23] ,
    \wbs_dat_o[24] , \wbs_dat_o[25] , \wbs_dat_o[26] , \wbs_dat_o[27] ,
    \wbs_dat_o[28] , \wbs_dat_o[29] , \wbs_dat_o[30] , \wbs_dat_o[31] ,
    \wbm_adr_o[0] , \wbm_adr_o[1] , \wbm_adr_o[2] , \wbm_adr_o[3] ,
    \wbm_adr_o[4] , \wbm_adr_o[5] , \wbm_adr_o[6] , \wbm_adr_o[7] ,
    \wbm_adr_o[8] , \wbm_adr_o[9] , \wbm_adr_o[10] , \wbm_adr_o[11] ,
    \wbm_adr_o[12] , \wbm_adr_o[13] , \wbm_adr_o[14] , \wbm_adr_o[15] ,
    \wbm_adr_o[16] , \wbm_adr_o[17] , \wbm_adr_o[18] , \wbm_adr_o[19] ,
    \wbm_adr_o[20] , \wbm_adr_o[21] , \wbm_adr_o[22] , \wbm_adr_o[23] ,
    \wbm_adr_o[24] , \wbm_adr_o[25] , \wbm_adr_o[26] , \wbm_adr_o[27] ,
    \wbm_adr_o[28] , \wbm_adr_o[29] , \wbm_adr_o[30] , \wbm_adr_o[31] ,
    \wbm_dat_o[0] , \wbm_dat_o[1] , \wbm_dat_o[2] , \wbm_dat_o[3] ,
    \wbm_dat_o[4] , \wbm_dat_o[5] , \wbm_dat_o[6] , \wbm_dat_o[7] ,
    \wbm_dat_o[8] , \wbm_dat_o[9] , \wbm_dat_o[10] , \wbm_dat_o[11] ,
    \wbm_dat_o[12] , \wbm_dat_o[13] , \wbm_dat_o[14] , \wbm_dat_o[15] ,
    \wbm_dat_o[16] , \wbm_dat_o[17] , \wbm_dat_o[18] , \wbm_dat_o[19] ,
    \wbm_dat_o[20] , \wbm_dat_o[21] , \wbm_dat_o[22] , \wbm_dat_o[23] ,
    \wbm_dat_o[24] , \wbm_dat_o[25] , \wbm_dat_o[26] , \wbm_dat_o[27] ,
    \wbm_dat_o[28] , \wbm_dat_o[29] , \wbm_dat_o[30] , \wbm_dat_o[31] ,
    \pci_ad_oe_o[0] , \pci_ad_oe_o[1] , \pci_ad_oe_o[2] , \pci_ad_oe_o[3] ,
    \pci_ad_oe_o[4] , \pci_ad_oe_o[5] , \pci_ad_oe_o[6] , \pci_ad_oe_o[7] ,
    \pci_ad_oe_o[8] , \pci_ad_oe_o[9] , \pci_ad_oe_o[10] ,
    \pci_ad_oe_o[11] , \pci_ad_oe_o[12] , \pci_ad_oe_o[13] ,
    \pci_ad_oe_o[14] , \pci_ad_oe_o[15] , \pci_ad_oe_o[16] ,
    \pci_ad_oe_o[17] , \pci_ad_oe_o[18] , \pci_ad_oe_o[19] ,
    \pci_ad_oe_o[20] , \pci_ad_oe_o[21] , \pci_ad_oe_o[22] ,
    \pci_ad_oe_o[23] , \pci_ad_oe_o[24] , \pci_ad_oe_o[25] ,
    \pci_ad_oe_o[26] , \pci_ad_oe_o[27] , \pci_ad_oe_o[28] ,
    \pci_ad_oe_o[29] , \pci_ad_oe_o[30] , \pci_ad_oe_o[31] , \pci_ad_o[0] ,
    \pci_ad_o[1] , \pci_ad_o[2] , \pci_ad_o[3] , \pci_ad_o[4] ,
    \pci_ad_o[5] , \pci_ad_o[6] , \pci_ad_o[7] , \pci_ad_o[8] ,
    \pci_ad_o[9] , \pci_ad_o[10] , \pci_ad_o[11] , \pci_ad_o[12] ,
    \pci_ad_o[13] , \pci_ad_o[14] , \pci_ad_o[15] , \pci_ad_o[16] ,
    \pci_ad_o[17] , \pci_ad_o[18] , \pci_ad_o[19] , \pci_ad_o[20] ,
    \pci_ad_o[21] , \pci_ad_o[22] , \pci_ad_o[23] , \pci_ad_o[24] ,
    \pci_ad_o[25] , \pci_ad_o[26] , \pci_ad_o[27] , \pci_ad_o[28] ,
    \pci_ad_o[29] , \pci_ad_o[30] , \pci_ad_o[31] , \wbm_sel_o[0] ,
    \wbm_sel_o[1] , \wbm_sel_o[2] , \wbm_sel_o[3] , \pci_cbe_oe_o[0] ,
    \pci_cbe_oe_o[1] , \pci_cbe_oe_o[2] , \pci_cbe_oe_o[3] ,
    \pci_cbe_o[0] , \pci_cbe_o[1] , \pci_cbe_o[2] , \pci_cbe_o[3] ,
    \wbm_cti_o[0] , \wbm_cti_o[1] , \wbm_cti_o[2] , \wbm_bte_o[0] ,
    \wbm_bte_o[1] ;
  reg \\pci_target_unit_wishbone_master_wb_cti_o_reg[0] ,
    \\pci_target_unit_wishbone_master_wb_cti_o_reg[2] ,
    configuration_status_bit8_reg,
    \\pci_target_unit_wishbone_master_wb_sel_o_reg[0] ,
    \\pci_target_unit_wishbone_master_wb_sel_o_reg[1] ,
    \\pci_target_unit_wishbone_master_wb_sel_o_reg[2] ,
    \\pci_target_unit_wishbone_master_wb_sel_o_reg[3] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[0] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[10] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[11] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[12] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[13] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[16] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[17] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[19] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[1] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[20] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[21] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[22] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[23] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[24] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[25] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[26] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[27] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[28] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[29] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[2] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[31] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[3] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[4] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[5] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[6] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[8] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[9] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[30] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[14] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[18] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[7] ,
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[15] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[19] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[22] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[24] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[20] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[27] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[21] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[30] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[25] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[28] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[31] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[29] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[17] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[10] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[11] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[12] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[16] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[14] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[13] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[23] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[26] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[3] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[4] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[5] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[6] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[8] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[9] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[2] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[18] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[15] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[7] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[0] ,
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[1] ,
    parity_checker_perr_sampled_reg,
    \\pci_target_unit_wishbone_master_bc_register_reg[0] ,
    \\pci_target_unit_wishbone_master_bc_register_reg[1] ,
    \\pci_target_unit_wishbone_master_bc_register_reg[2] ,
    \\pci_target_unit_wishbone_master_bc_register_reg[3] ,
    pci_target_unit_wishbone_master_burst_chopped_reg,
    pci_target_unit_pci_target_sm_backoff_reg,
    wishbone_slave_unit_del_sync_req_done_reg_reg,
    \\wishbone_slave_unit_wishbone_slave_c_state_reg[0] ,
    \\pci_target_unit_wishbone_master_wb_cti_o_reg[1] ,
    wishbone_slave_unit_del_sync_req_comp_pending_reg,
    \\wishbone_slave_unit_wishbone_slave_c_state_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[38] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[10] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[11] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[12] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[13] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[16] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[14] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[17] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[19] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[20] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[21] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[22] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[23] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[24] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[25] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[26] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[27] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[28] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[29] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[30] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[31] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[32] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[33] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[34] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[35] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[37] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[3] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[4] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[5] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[6] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[8] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[9] ,
    output_backup_trdy_out_reg, pci_io_mux_trdy_iob_dat_out_reg,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[15] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[18] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[7] ,
    pci_io_mux_stop_iob_dat_out_reg, output_backup_stop_out_reg,
    pci_io_mux_devsel_iob_dat_out_reg, output_backup_devsel_out_reg,
    output_backup_perr_en_out_reg, \\output_backup_ad_out_reg[31] ,
    pci_io_mux_ad_iob31_dat_out_reg, pci_io_mux_perr_iob_en_out_reg,
    \\configuration_status_bit15_11_reg[15] ,
    wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg,
    \\output_backup_cbe_out_reg[0] , \\output_backup_cbe_out_reg[3] ,
    pci_io_mux_cbe_iob0_dat_out_reg, pci_io_mux_cbe_iob2_dat_out_reg,
    \\output_backup_cbe_out_reg[2] , pci_io_mux_cbe_iob3_dat_out_reg,
    \\output_backup_ad_out_reg[15] , \\output_backup_ad_out_reg[23] ,
    \\output_backup_ad_out_reg[24] , \\output_backup_ad_out_reg[27] ,
    \\output_backup_ad_out_reg[28] , \\output_backup_ad_out_reg[29] ,
    \\output_backup_ad_out_reg[2] , \\output_backup_ad_out_reg[3] ,
    \\output_backup_ad_out_reg[4] , \\output_backup_ad_out_reg[5] ,
    \\output_backup_ad_out_reg[6] , \\output_backup_ad_out_reg[7] ,
    \\output_backup_ad_out_reg[8] , pci_io_mux_ad_iob11_dat_out_reg,
    pci_io_mux_ad_iob12_dat_out_reg, pci_io_mux_ad_iob13_dat_out_reg,
    pci_io_mux_ad_iob14_dat_out_reg, pci_io_mux_ad_iob15_dat_out_reg,
    pci_io_mux_ad_iob24_dat_out_reg, pci_io_mux_ad_iob27_dat_out_reg,
    pci_io_mux_ad_iob29_dat_out_reg, pci_io_mux_ad_iob28_dat_out_reg,
    pci_io_mux_ad_iob2_dat_out_reg, pci_io_mux_ad_iob4_dat_out_reg,
    pci_io_mux_ad_iob5_dat_out_reg, pci_io_mux_ad_iob6_dat_out_reg,
    pci_io_mux_ad_iob7_dat_out_reg, pci_io_mux_ad_iob23_dat_out_reg,
    pci_io_mux_ad_iob8_dat_out_reg, pci_io_mux_ad_iob3_dat_out_reg,
    \\output_backup_ad_out_reg[13] , \\output_backup_ad_out_reg[14] ,
    \\output_backup_ad_out_reg[16] , \\output_backup_ad_out_reg[17] ,
    \\output_backup_ad_out_reg[18] , \\output_backup_ad_out_reg[19] ,
    \\output_backup_ad_out_reg[20] , \\output_backup_ad_out_reg[22] ,
    \\output_backup_ad_out_reg[9] , pci_io_mux_ad_iob10_dat_out_reg,
    pci_io_mux_ad_iob16_dat_out_reg, pci_io_mux_ad_iob17_dat_out_reg,
    pci_io_mux_ad_iob18_dat_out_reg, pci_io_mux_ad_iob19_dat_out_reg,
    pci_io_mux_ad_iob22_dat_out_reg, pci_io_mux_ad_iob20_dat_out_reg,
    \\output_backup_ad_out_reg[10] , pci_io_mux_ad_iob9_dat_out_reg,
    \\output_backup_ad_out_reg[11] , \\output_backup_ad_out_reg[12] ,
    \\output_backup_ad_out_reg[1] , \\output_backup_ad_out_reg[30] ,
    pci_io_mux_ad_iob1_dat_out_reg, pci_io_mux_ad_iob30_dat_out_reg,
    \\output_backup_ad_out_reg[21] , pci_io_mux_ad_iob21_dat_out_reg,
    \\configuration_status_bit15_11_reg[14] ,
    \\output_backup_ad_out_reg[26] , pci_io_mux_ad_iob26_dat_out_reg,
    pci_io_mux_ad_iob0_dat_out_reg, \\output_backup_ad_out_reg[0] ,
    parity_checker_perr_en_crit_gen_perr_en_reg_out_reg,
    \\output_backup_ad_out_reg[25] , pci_io_mux_ad_iob25_dat_out_reg,
    \\wishbone_slave_unit_pci_initiator_if_be_out_reg[0] ,
    \\wishbone_slave_unit_pci_initiator_if_be_out_reg[2] ,
    \\wishbone_slave_unit_pci_initiator_if_be_out_reg[3] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[10] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[11] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[16] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[18] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[19] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[1] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[21] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[22] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[30] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[5] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[6] ,
    pci_io_mux_perr_iob_dat_out_reg, pci_io_mux_serr_iob_en_out_reg,
    pci_io_mux_serr_iob_dat_out_reg,
    pci_target_unit_wishbone_master_first_wb_data_access_reg,
    output_backup_perr_out_reg, output_backup_serr_out_reg,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[15] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[24] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[25] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[27] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[2] ,
    output_backup_serr_en_out_reg,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[0] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[12] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[13] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[14] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[17] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[20] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[23] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[26] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[28] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[29] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[31] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[3] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[4] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[7] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[8] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[9] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[26] ,
    \\pci_target_unit_fifos_pciw_outTransactionCount_reg[1] ,
    \\pci_target_unit_fifos_outGreyCount_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[0] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[2] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[0] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[10] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[11] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[12] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[13] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[14] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[15] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[17] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[18] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[19] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[20] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[22] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[24] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[27] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[28] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[29] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[2] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[31] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[3] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[4] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[6] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[7] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[8] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10] ,
    \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[2] ,
    \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[3] ,
    \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[0] ,
    \\wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[0] ,
    \\pci_target_unit_fifos_pciw_outTransactionCount_reg[0] ,
    \\pci_target_unit_fifos_outGreyCount_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg[1] ,
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9] ,
    \\wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[1] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[5] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[9] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[1] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[23] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[16] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[3] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[21] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[25] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0] ,
    pci_target_unit_wishbone_master_wb_we_o_reg,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2] ,
    pci_target_unit_wishbone_master_wb_cyc_o_reg,
    pci_target_unit_wishbone_master_wb_stb_o_reg,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[6] ,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_reg[1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[9] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[15] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[25] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[7] ,
    parity_checker_check_perr_reg,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[0] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[10] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[11] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[13] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[14] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[17] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[18] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[19] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[21] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[22] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[20] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[24] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[26] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[28] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[29] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[2] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[31] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[3] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[4] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[6] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[8] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[9] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[5] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[30] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[27] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[23] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[12] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[1] ,
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26] ,
    output_backup_par_en_out_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36] ,
    pci_io_mux_par_iob_en_out_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[25] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[15] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[7] ,
    \\pci_target_unit_wishbone_master_c_state_reg[0] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[17] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[18] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[16] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[19] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[1] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[20] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[21] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[23] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[24] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[22] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[26] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[27] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[28] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[29] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[2] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[30] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[31] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[3] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[4] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[5] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[6] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[8] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[9] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[37] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[0] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[10] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[11] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[12] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[13] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[14] ,
    i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg,
    pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28] ,
    i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][19] ,
    pci_io_mux_ad_iob23_en_out_reg, pci_io_mux_ad_iob22_en_out_reg,
    pci_io_mux_ad_iob21_en_out_reg, pci_io_mux_ad_iob19_en_out_reg,
    pci_io_mux_ad_iob17_en_out_reg, pci_io_mux_ad_iob18_en_out_reg,
    pci_io_mux_ad_iob15_en_out_reg, pci_io_mux_ad_iob14_en_out_reg,
    pci_io_mux_ad_iob13_en_out_reg, pci_io_mux_ad_iob11_en_out_reg,
    pci_io_mux_ad_iob25_en_out_reg, pci_io_mux_ad_iob8_en_out_reg,
    pci_io_mux_ad_iob7_en_out_reg, pci_io_mux_ad_iob9_en_out_reg,
    pci_io_mux_ad_iob5_en_out_reg, pci_io_mux_ad_iob3_en_out_reg,
    pci_io_mux_ad_iob4_en_out_reg, pci_io_mux_ad_iob1_en_out_reg,
    pci_io_mux_ad_iob2_en_out_reg, pci_io_mux_ad_iob26_en_out_reg,
    pci_io_mux_ad_iob31_en_out_reg, pci_io_mux_ad_iob29_en_out_reg,
    pci_io_mux_ad_iob28_en_out_reg, pci_io_mux_ad_iob27_en_out_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][13] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][13] ,
    output_backup_mas_ad_en_out_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][15] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][23] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][24] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][26] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][30] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][7] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][8] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][9] ,
    output_backup_tar_ad_en_out_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][11] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][17] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][28] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][27] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][35] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][19] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][3] ,
    pci_io_mux_ad_iob30_en_out_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][29] ,
    pci_io_mux_ad_iob0_en_out_reg, pci_io_mux_ad_iob6_en_out_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][18] ,
    pci_io_mux_ad_iob12_en_out_reg, pci_io_mux_ad_iob10_en_out_reg,
    pci_io_mux_ad_iob16_en_out_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][3] ,
    pci_io_mux_ad_iob20_en_out_reg, pci_io_mux_ad_iob24_en_out_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][10] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][20] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][16] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][21] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][18] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][32] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][32] ,
    pci_target_unit_wishbone_master_first_data_is_burst_reg_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][33] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][25] ,
    i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][12] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][22] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][6] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][5] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][34] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][14] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][25] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[0] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[10] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[11] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[13] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[15] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[16] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[17] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[19] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[1] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[20] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[23] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[24] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[26] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[27] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[28] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[30] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[31] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[7] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[8] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[9] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[3] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[29] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[18] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[21] ,
    \\pci_target_unit_pci_target_sm_c_state_reg[0] ,
    \\pci_target_unit_pci_target_sm_c_state_reg[1] ,
    \\pci_target_unit_pci_target_sm_c_state_reg[2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3] ,
    \\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[1] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[12] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[22] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[2] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[5] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][36] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[25] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[6] ,
    \\wishbone_slave_unit_del_sync_addr_out_reg[14] ,
    \\wishbone_slave_unit_fifos_inGreyCount_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2] ,
    \\wishbone_slave_unit_fifos_inGreyCount_reg[1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][36] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][36] ,
    \\wishbone_slave_unit_fifos_inGreyCount_reg[2] ,
    \\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0] ,
    i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[0] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[1] ,
    wishbone_slave_unit_del_sync_burst_out_reg,
    pci_target_unit_wishbone_master_addr_into_cnt_reg_reg,
    output_backup_trdy_en_out_reg,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[2] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1] ,
    pci_io_mux_trdy_iob_en_out_reg, pci_io_mux_stop_iob_en_out_reg,
    pci_io_mux_devsel_iob_en_out_reg,
    \\pci_target_unit_wishbone_master_rty_counter_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0] ,
    \\wishbone_slave_unit_del_sync_bc_out_reg[3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0] ,
    output_backup_frame_out_reg,
    \\pci_target_unit_wishbone_master_rty_counter_reg[5] ,
    \\pci_target_unit_wishbone_master_rty_counter_reg[6] ,
    \\wishbone_slave_unit_del_sync_bc_out_reg[2] ,
    \\pci_target_unit_wishbone_master_rty_counter_reg[1] ,
    \\pci_target_unit_wishbone_master_rty_counter_reg[2] ,
    \\pci_target_unit_wishbone_master_rty_counter_reg[4] ,
    \\wishbone_slave_unit_fifos_outGreyCount_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3] ,
    \\pci_target_unit_wishbone_master_rty_counter_reg[3] ,
    \\pci_target_unit_wishbone_master_rty_counter_reg[7] ,
    pci_io_mux_frame_iob_dat_out_reg,
    pci_target_unit_pci_target_sm_rd_request_reg,
    pci_target_unit_pci_target_sm_rd_progress_reg,
    \\wishbone_slave_unit_del_sync_be_out_reg[0] ,
    \\wishbone_slave_unit_del_sync_be_out_reg[1] ,
    \\wishbone_slave_unit_del_sync_be_out_reg[2] ,
    wishbone_slave_unit_del_sync_we_out_reg,
    \\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[1] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1] ,
    \\wishbone_slave_unit_del_sync_be_out_reg[3] ,
    \\wishbone_slave_unit_del_sync_bc_out_reg[1] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[12] ,
    pci_target_unit_pci_target_if_norm_prf_en_reg,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[0] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[10] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[11] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[13] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[14] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[15] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[17] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[18] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[1] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[21] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[23] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[25] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[26] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[27] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[29] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[2] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[30] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[32] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[33] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[34] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[3] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[5] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[8] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[7] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[0] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[10] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[11] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[14] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[1] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[3] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[5] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[9] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[7] ,
    \\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0] ,
    pci_target_unit_pci_target_if_pciw_fifo_wenable_out_reg,
    \\wishbone_slave_unit_fifos_outGreyCount_reg[2] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[6] ,
    \\wishbone_slave_unit_fifos_outGreyCount_reg[1] ,
    \\wishbone_slave_unit_del_sync_bc_out_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2] ,
    i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[6] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[4] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[13] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[2] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[15] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[16] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[9] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[4] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[35] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[31] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[22] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[28] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[24] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[16] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[20] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[12] ,
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[19] ,
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[8] ,
    pci_target_unit_pci_target_sm_wr_progress_reg,
    pci_target_unit_wishbone_master_w_attempt_reg,
    \\configuration_wb_am2_reg[31] , \\configuration_wb_am1_reg[31] ,
    pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg,
    \\output_backup_cbe_out_reg[1] ,
    wishbone_slave_unit_pci_initiator_if_del_read_req_reg,
    \\configuration_pci_img_ctrl1_bit2_1_reg[1] ,
    \\configuration_pci_img_ctrl1_bit2_1_reg[2] ,
    \\configuration_wb_ta1_reg[31] , configuration_wb_err_cs_bit0_reg,
    \\configuration_wb_ta2_reg[31] , pci_io_mux_cbe_iob1_dat_out_reg,
    pci_target_unit_pci_target_sm_master_will_request_read_reg,
    wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg,
    output_backup_par_out_reg, pci_io_mux_par_iob_dat_out_reg,
    configuration_pci_err_cs_bit0_reg,
    \\configuration_wb_img_ctrl1_bit2_0_reg[2] ,
    \\configuration_interrupt_line_reg[6] ,
    \\configuration_wb_img_ctrl2_bit2_0_reg[1] ,
    \\configuration_interrupt_line_reg[2] ,
    wishbone_slave_unit_del_sync_req_req_pending_reg,
    \\configuration_wb_img_ctrl1_bit2_0_reg[0] ,
    \\configuration_wb_img_ctrl1_bit2_0_reg[1] ,
    \\configuration_interrupt_line_reg[0] ,
    \\configuration_interrupt_line_reg[1] ,
    \\configuration_wb_img_ctrl2_bit2_0_reg[0] ,
    \\configuration_wb_img_ctrl2_bit2_0_reg[2] ,
    \\configuration_command_bit2_0_reg[0] ,
    \\configuration_command_bit2_0_reg[1] ,
    \\configuration_command_bit2_0_reg[2] , configuration_wb_ba1_bit0_reg,
    configuration_wb_ba2_bit0_reg, configuration_command_bit8_reg,
    configuration_wb_err_cs_bit8_reg,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1] ,
    \\configuration_status_bit15_11_reg[11] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1] ,
    \\configuration_status_bit15_11_reg[12] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0] ,
    \\configuration_status_bit15_11_reg[13] ,
    \\configuration_isr_bit2_0_reg[1] ,
    wishbone_slave_unit_del_sync_comp_comp_pending_reg,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[0] ,
    pci_target_unit_wishbone_master_reset_rty_cnt_reg,
    \\configuration_wb_ba2_bit31_12_reg[31] ,
    \\configuration_wb_ba1_bit31_12_reg[31] ,
    configuration_command_bit6_reg,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][1] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][6] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][3] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[1] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][26] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][31] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][2] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][22] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][24] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][19] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][20] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][11] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][0] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][8] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][15] ,
    \\configuration_icr_bit2_0_reg[0] , \\configuration_icr_bit2_0_reg[1] ,
    \\configuration_icr_bit2_0_reg[2] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][4] ,
    \\configuration_interrupt_line_reg[3] ,
    \\configuration_cache_line_size_reg_reg[3] ,
    \\configuration_interrupt_line_reg[5] ,
    \\configuration_interrupt_line_reg[4] ,
    \\configuration_cache_line_size_reg_reg[5] ,
    \\configuration_cache_line_size_reg_reg[4] ,
    configuration_sync_isr_2_del_bit_reg,
    configuration_sync_pci_err_cs_8_del_bit_reg,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[0] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[2] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][0] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][10] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][12] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][14] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][16] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][18] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][1] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][20] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][21] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][23] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][25] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][27] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][29] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][30] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][37] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][4] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][5] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][6] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][8] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][0] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][11] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][12] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][13] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][15] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][16] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][17] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][19] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][1] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][20] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][22] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][24] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][26] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][28] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][2] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][31] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][3] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][4] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][5] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][7] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][8] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][9] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][10] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][11] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][12] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][14] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][16] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][18] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][19] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][1] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][21] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][23] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][25] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][26] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][27] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][29] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][30] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][37] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][3] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][4] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][6] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][7] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][8] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][0] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][10] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][11] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][13] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][15] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][17] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][18] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][19] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][20] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][22] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][24] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][25] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][26] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][28] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][29] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][2] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][31] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][37] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][3] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][5] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][7] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][9] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][14] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][15] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][16] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][18] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][1] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][21] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][22] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][23] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][25] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][27] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][29] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][2] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][30] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][37] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][4] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][6] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][7] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][8] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][0] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][11] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][13] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][14] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][15] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][17] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][18] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][19] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][20] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][22] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][24] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][26] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][28] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][29] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][2] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][31] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][3] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][5] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][7] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][9] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][10] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][12] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][13] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][14] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][16] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][17] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][18] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][1] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][21] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][23] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][25] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][27] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][28] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][29] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][30] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][37] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][4] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][5] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][6] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][8] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][9] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][0] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][11] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][13] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][15] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][17] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][19] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][1] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][20] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][22] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][24] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][26] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][27] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][28] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][2] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][31] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][3] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][4] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][5] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][7] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][9] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][10] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][12] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][30] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][37] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][25] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][27] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][23] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][21] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][1] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][16] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][9] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][10] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][12] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][26] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][21] ,
    \\configuration_cache_line_size_reg_reg[7] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][3] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][5] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][31] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][28] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][24] ,
    \\configuration_interrupt_line_reg[7] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][19] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][20] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][17] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][4] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][8] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][6] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][30] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][27] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][23] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][8] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][9] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][28] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][14] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][16] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][12] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][5] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][2] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][31] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][24] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][22] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][0] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][0] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][20] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][11] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][13] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][17] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][13] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][15] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][29] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][6] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][6] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][37] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][21] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][30] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][29] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][30] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][37] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][25] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][23] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][25] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][10] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][18] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][27] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][16] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][18] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][23] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][12] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][14] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][21] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][14] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][10] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][9] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][7] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][7] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][28] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][2] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][3] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][31] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][26] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][22] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][24] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][13] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][19] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][17] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][15] ,
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][11] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[5] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[7] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[8] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[23] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[4] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[31] ,
    \\configuration_pci_ba0_bit31_8_reg[12] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[27] ,
    \\configuration_latency_timer_reg[1] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[12] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[1] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[21] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[14] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[16] ,
    \\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1] ,
    configuration_icr_bit31_reg,
    wishbone_slave_unit_wishbone_slave_img_wallow_reg,
    wishbone_slave_unit_wishbone_slave_do_del_request_reg,
    wishbone_slave_unit_wishbone_slave_mrl_en_reg,
    wishbone_slave_unit_wishbone_slave_pref_en_reg,
    wishbone_slave_unit_wishbone_slave_del_addr_hit_reg,
    \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[1] ,
    wishbone_slave_unit_wishbone_slave_del_completion_allow_reg,
    pci_target_unit_del_sync_comp_comp_pending_reg,
    pci_target_unit_del_sync_comp_req_pending_reg,
    \\pci_target_unit_wishbone_master_c_state_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][37] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][37] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][37] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][37] ,
    wishbone_slave_unit_pci_initiator_if_intermediate_last_reg,
    \\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[1] ,
    \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1] ,
    \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0] ,
    \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2] ,
    \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3] ,
    \\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0] ,
    \\configuration_latency_timer_reg[0] ,
    \\configuration_latency_timer_reg[2] ,
    \\configuration_latency_timer_reg[3] ,
    \\configuration_latency_timer_reg[4] ,
    \\configuration_latency_timer_reg[5] ,
    \\configuration_latency_timer_reg[6] ,
    \\configuration_latency_timer_reg[7] ,
    \\configuration_cache_line_size_reg_reg[0] ,
    \\configuration_pci_ba0_bit31_8_reg[14] ,
    \\configuration_cache_line_size_reg_reg[1] ,
    \\configuration_cache_line_size_reg_reg[2] ,
    \\configuration_pci_ba0_bit31_8_reg[13] ,
    \\configuration_pci_ba0_bit31_8_reg[17] ,
    \\configuration_cache_line_size_reg_reg[6] ,
    \\configuration_pci_ba0_bit31_8_reg[16] ,
    \\configuration_pci_ba0_bit31_8_reg[20] ,
    \\configuration_pci_ba0_bit31_8_reg[23] ,
    \\configuration_pci_ba0_bit31_8_reg[18] ,
    \\configuration_pci_ba0_bit31_8_reg[15] ,
    \\configuration_pci_ba0_bit31_8_reg[19] ,
    \\configuration_pci_ba0_bit31_8_reg[25] ,
    \\configuration_pci_ba0_bit31_8_reg[27] ,
    \\configuration_pci_ba0_bit31_8_reg[28] ,
    \\configuration_pci_ba0_bit31_8_reg[30] ,
    \\configuration_pci_ba0_bit31_8_reg[29] ,
    \\pci_target_unit_wishbone_master_read_count_reg[1] ,
    \\pci_target_unit_wishbone_master_read_count_reg[2] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[0] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[10] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[11] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[13] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[15] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[17] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[18] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[19] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[20] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[22] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[24] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[25] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[26] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[28] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[29] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[2] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[3] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[6] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[9] ,
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[30] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][37] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][37] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][37] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][37] ,
    wishbone_slave_unit_del_sync_comp_req_pending_reg,
    \\configuration_pci_ba0_bit31_8_reg[31] ,
    \\configuration_pci_ba0_bit31_8_reg[26] ,
    \\configuration_pci_ba0_bit31_8_reg[24] ,
    \\configuration_pci_ba0_bit31_8_reg[21] ,
    \\configuration_pci_ba0_bit31_8_reg[22] ,
    \\configuration_pci_am1_reg[16] , \\configuration_pci_am1_reg[15] ,
    \\configuration_pci_am1_reg[24] ,
    \\configuration_pci_ba1_bit31_8_reg[11] ,
    \\configuration_pci_ba1_bit31_8_reg[15] ,
    \\wishbone_slave_unit_pci_initiator_if_read_count_reg[3] ,
    wishbone_slave_unit_wishbone_slave_map_reg,
    \\configuration_pci_ba1_bit31_8_reg[18] ,
    \\configuration_pci_ba1_bit31_8_reg[19] ,
    \\configuration_pci_ba1_bit31_8_reg[20] ,
    \\configuration_pci_ba1_bit31_8_reg[21] ,
    \\configuration_pci_ba1_bit31_8_reg[23] ,
    \\configuration_pci_ba1_bit31_8_reg[25] ,
    \\configuration_pci_ba1_bit31_8_reg[26] ,
    \\configuration_pci_ba1_bit31_8_reg[27] ,
    \\configuration_pci_ba1_bit31_8_reg[29] ,
    \\configuration_pci_ba1_bit31_8_reg[30] ,
    \\configuration_pci_ba1_bit31_8_reg[10] ,
    \\configuration_pci_ba1_bit31_8_reg[12] ,
    \\configuration_pci_ba1_bit31_8_reg[13] ,
    \\configuration_pci_ba1_bit31_8_reg[14] ,
    \\configuration_pci_ba1_bit31_8_reg[16] ,
    \\pci_target_unit_wishbone_master_c_state_reg[1] ,
    \\configuration_pci_am1_reg[21] , \\configuration_pci_am1_reg[10] ,
    \\configuration_pci_am1_reg[12] , \\configuration_pci_am1_reg[11] ,
    \\configuration_pci_am1_reg[13] , \\configuration_pci_am1_reg[18] ,
    \\configuration_pci_am1_reg[17] , \\configuration_pci_am1_reg[20] ,
    \\configuration_pci_am1_reg[14] , \\configuration_pci_am1_reg[22] ,
    \\configuration_pci_am1_reg[23] , \\configuration_pci_am1_reg[25] ,
    \\configuration_pci_am1_reg[19] , \\configuration_pci_am1_reg[29] ,
    \\configuration_pci_am1_reg[31] , \\configuration_pci_am1_reg[30] ,
    \\configuration_pci_am1_reg[28] ,
    \\pci_target_unit_wishbone_master_read_count_reg[0] ,
    \\configuration_pci_ba1_bit31_8_reg[31] ,
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[1] ,
    \\configuration_pci_ba1_bit31_8_reg[8] ,
    \\configuration_pci_ba1_bit31_8_reg[9] ,
    \\configuration_pci_ba1_bit31_8_reg[22] ,
    \\configuration_pci_ba1_bit31_8_reg[28] ,
    \\configuration_pci_ba1_bit31_8_reg[24] ,
    \\configuration_pci_ba1_bit31_8_reg[17] ,
    wishbone_slave_unit_pci_initiator_if_current_last_reg,
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[0] ,
    \\configuration_pci_am1_reg[26] , \\configuration_pci_am1_reg[8] ,
    \\configuration_pci_am1_reg[9] , \\configuration_pci_am1_reg[27] ,
    \\wishbone_slave_unit_wishbone_slave_c_state_reg[1] ,
    \\configuration_pci_ta1_reg[10] ,
    pci_target_unit_wishbone_master_read_bound_reg,
    \\configuration_pci_ta1_reg[29] , \\configuration_pci_ta1_reg[16] ,
    \\wishbone_slave_unit_pci_initiator_if_read_count_reg[2] ,
    \\configuration_pci_ta1_reg[17] , \\configuration_pci_ta1_reg[18] ,
    \\configuration_pci_ta1_reg[20] , \\configuration_pci_ta1_reg[21] ,
    \\configuration_pci_ta1_reg[24] , \\configuration_pci_ta1_reg[23] ,
    \\configuration_pci_ta1_reg[30] , \\configuration_pci_ta1_reg[28] ,
    \\configuration_pci_ta1_reg[31] , \\configuration_pci_ta1_reg[14] ,
    wishbone_slave_unit_pci_initiator_if_err_recovery_reg,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][37] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][37] ,
    \\configuration_pci_ta1_reg[11] , \\configuration_pci_ta1_reg[13] ,
    \\configuration_pci_ta1_reg[15] , \\configuration_pci_ta1_reg[12] ,
    \\configuration_pci_ta1_reg[8] , \\configuration_pci_ta1_reg[9] ,
    \\configuration_pci_ta1_reg[27] , \\configuration_pci_ta1_reg[26] ,
    \\configuration_pci_ta1_reg[25] , \\configuration_pci_ta1_reg[22] ,
    \\configuration_pci_ta1_reg[19] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][32] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][32] ,
    wishbone_slave_unit_pci_initiator_if_posted_write_req_reg,
    pci_io_mux_frame_iob_en_out_reg,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[27] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[17] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[19] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[20] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[22] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[23] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[24] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[28] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[29] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[2] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[31] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[3] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[4] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[6] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[8] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[16] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[0] ,
    output_backup_cbe_en_out_reg,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][32] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][32] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][32] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][32] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][36] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][32] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[13] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[15] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[9] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[5] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[7] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][36] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[26] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[30] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[18] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[21] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[1] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[12] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[25] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[11] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[0] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[10] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][36] ,
    \\wishbone_slave_unit_pci_initiator_if_be_out_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][32] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][0] ,
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][1] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[16] ,
    configuration_set_isr_bit2_reg,
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[2] ,
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[3] ,
    wishbone_slave_unit_wishbone_slave_wb_conf_hit_reg,
    \\configuration_wb_err_addr_reg[0] ,
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6] ,
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2] ,
    output_backup_frame_en_out_reg,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][1] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][0] ,
    pci_io_mux_cbe_iob3_en_out_reg, pci_io_mux_cbe_iob2_en_out_reg,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][9] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][36] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][14] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][36] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][7] ,
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][4] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][1] ,
    configuration_wb_err_cs_bit9_reg,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][26] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][1] ,
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][18] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][27] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][12] ,
    pci_io_mux_cbe_iob1_en_out_reg, pci_io_mux_cbe_iob0_en_out_reg,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][29] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][30] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][25] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][12] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][14] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][10] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][4] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][6] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][15] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][16] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][9] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][31] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][6] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][7] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][8] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][4] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][28] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][22] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][26] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][21] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][11] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][12] ,
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][12] ,
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][22] ,
    i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][18] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][20] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][23] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][13] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][19] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][24] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][36] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][17] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][15] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][16] ,
    \\configuration_wb_err_addr_reg[11] ,
    \\configuration_wb_err_data_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][20] ,
    \\configuration_wb_err_cs_bit31_24_reg[30] ,
    \\configuration_wb_err_addr_reg[19] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][25] ,
    \\configuration_pci_err_data_reg[28] ,
    wishbone_slave_unit_pci_initiator_if_data_source_reg,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][9] ,
    \\configuration_wb_err_cs_bit31_24_reg[28] ,
    \\configuration_wb_err_addr_reg[15] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][16] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][4] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][14] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][22] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][4] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][30] ,
    \\configuration_wb_err_data_reg[6] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][21] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][24] ,
    \\configuration_wb_err_data_reg[8] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][27] ,
    \\configuration_wb_err_data_reg[30] ,
    \\configuration_wb_err_data_reg[4] ,
    \\configuration_wb_err_data_reg[31] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][15] ,
    \\configuration_wb_err_data_reg[28] ,
    \\configuration_wb_err_data_reg[27] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][29] ,
    \\configuration_wb_err_data_reg[24] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][23] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][22] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][18] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][21] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][21] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][16] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][12] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][35] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][26] ,
    \\configuration_wb_err_data_reg[20] ,
    wishbone_slave_unit_pci_initiator_if_read_bound_reg,
    configuration_pci_err_cs_bit9_reg, configuration_pci_err_cs_bit10_reg,
    \\configuration_pci_err_cs_bit31_24_reg[30] ,
    \\configuration_pci_err_cs_bit31_24_reg[28] ,
    \\configuration_pci_err_cs_bit31_24_reg[29] ,
    \\wishbone_slave_unit_pci_initiator_if_read_count_reg[1] ,
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4] ,
    \\configuration_pci_err_addr_reg[0] ,
    \\configuration_pci_err_addr_reg[11] ,
    \\configuration_pci_err_addr_reg[12] ,
    \\configuration_pci_err_addr_reg[15] ,
    \\configuration_pci_err_addr_reg[19] ,
    \\configuration_pci_err_addr_reg[20] ,
    \\configuration_pci_err_addr_reg[22] ,
    \\configuration_pci_err_addr_reg[26] ,
    \\configuration_pci_err_addr_reg[28] ,
    \\configuration_pci_err_addr_reg[2] ,
    \\configuration_pci_err_addr_reg[31] ,
    \\configuration_pci_err_addr_reg[4] ,
    \\configuration_pci_err_addr_reg[6] ,
    \\configuration_pci_err_addr_reg[8] ,
    \\configuration_pci_err_data_reg[0] ,
    \\configuration_pci_err_data_reg[11] ,
    \\configuration_pci_err_data_reg[13] ,
    \\configuration_pci_err_data_reg[15] ,
    \\configuration_pci_err_data_reg[17] ,
    \\configuration_pci_err_data_reg[19] ,
    \\configuration_pci_err_data_reg[21] ,
    \\configuration_pci_err_data_reg[25] ,
    \\configuration_pci_err_data_reg[29] ,
    \\configuration_pci_err_data_reg[31] ,
    \\configuration_pci_err_data_reg[3] ,
    \\configuration_pci_err_data_reg[7] ,
    pci_target_unit_pci_target_sm_same_read_reg_reg,
    \\configuration_wb_err_cs_bit31_24_reg[25] ,
    \\configuration_wb_err_cs_bit31_24_reg[31] ,
    \\configuration_wb_err_data_reg[10] ,
    \\configuration_wb_err_data_reg[11] ,
    \\configuration_wb_err_data_reg[12] ,
    \\configuration_wb_err_data_reg[14] ,
    \\configuration_wb_err_data_reg[15] ,
    \\configuration_wb_err_data_reg[16] ,
    \\configuration_wb_err_data_reg[18] ,
    \\configuration_wb_err_data_reg[19] ,
    \\configuration_wb_err_data_reg[1] ,
    \\configuration_wb_err_data_reg[21] ,
    \\configuration_wb_err_data_reg[22] ,
    \\configuration_wb_err_data_reg[23] ,
    \\configuration_wb_err_data_reg[25] ,
    \\configuration_wb_err_data_reg[26] ,
    \\configuration_wb_err_data_reg[29] ,
    \\configuration_wb_err_data_reg[2] ,
    \\configuration_wb_err_data_reg[3] ,
    \\configuration_wb_err_data_reg[5] ,
    \\configuration_wb_err_data_reg[9] ,
    \\configuration_wb_err_data_reg[7] ,
    \\configuration_wb_err_addr_reg[10] ,
    \\configuration_wb_err_addr_reg[12] ,
    \\configuration_wb_err_addr_reg[13] ,
    \\configuration_wb_err_addr_reg[14] ,
    \\configuration_wb_err_addr_reg[16] ,
    \\configuration_wb_err_addr_reg[18] ,
    \\configuration_wb_err_addr_reg[20] ,
    \\configuration_wb_err_addr_reg[22] ,
    \\configuration_wb_err_addr_reg[24] ,
    \\configuration_wb_err_addr_reg[26] ,
    \\configuration_wb_err_addr_reg[28] ,
    \\configuration_wb_err_addr_reg[2] ,
    \\configuration_wb_err_addr_reg[31] ,
    \\configuration_wb_err_addr_reg[4] ,
    \\configuration_wb_err_addr_reg[6] ,
    \\configuration_wb_err_addr_reg[7] ,
    \\configuration_wb_err_addr_reg[8] ,
    \\pci_target_unit_fifos_pciw_inTransactionCount_reg[1] ,
    \\pci_target_unit_fifos_inGreyCount_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][17] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][12] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][11] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][20] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][7] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][24] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][3] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][34] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][33] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][15] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][29] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][11] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][13] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][15] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][17] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][20] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][23] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][25] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][28] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][18] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][30] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][34] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][35] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][5] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][7] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][10] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][12] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][17] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][22] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][24] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][31] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][8] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][16] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][19] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][22] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][26] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][2] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][34] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][33] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][5] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][7] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][9] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][14] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][10] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][17] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][20] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][22] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][24] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][23] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][21] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][25] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][12] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][34] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][5] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][7] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][16] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][23] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][21] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][14] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][11] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][13] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][15] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][17] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][19] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][27] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][2] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][3] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][4] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][6] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][7] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][16] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][20] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][22] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][27] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][29] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][33] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][6] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][8] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][10] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][14] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][9] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][19] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][23] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][28] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][8] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][11] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][21] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][24] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][27] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][2] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][18] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][29] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][35] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][26] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][38] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][38] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][38] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][38] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][13] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][18] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][13] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][25] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][19] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][15] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][20] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][28] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][12] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][14] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][9] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][18] ,
    \\configuration_wb_err_cs_bit31_24_reg[29] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][33] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][27] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][6] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][35] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][5] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][6] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][6] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][3] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][8] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][23] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][22] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][4] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][9] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][6] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][15] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][30] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][8] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][11] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][13] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][9] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][14] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][19] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][4] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][3] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][33] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][2] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][31] ,
    \\configuration_wb_err_data_reg[13] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][27] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][29] ,
    \\configuration_wb_err_cs_bit31_24_reg[24] ,
    \\configuration_wb_err_cs_bit31_24_reg[27] ,
    \\configuration_wb_err_cs_bit31_24_reg[26] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][12] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][3] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][10] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][7] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][4] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][29] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][11] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][28] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][5] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][16] ,
    \\configuration_wb_err_data_reg[17] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][4] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][31] ,
    \\configuration_pci_err_data_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][35] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][31] ,
    \\configuration_wb_err_addr_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][22] ,
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[7] ,
    pci_target_unit_pci_target_if_same_read_reg_reg,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][34] ,
    \\configuration_pci_err_data_reg[8] ,
    \\configuration_pci_err_data_reg[30] ,
    \\configuration_pci_err_data_reg[9] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][13] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][20] ,
    \\configuration_pci_err_data_reg[5] ,
    \\configuration_pci_err_data_reg[6] ,
    \\configuration_pci_err_data_reg[4] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][6] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][2] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][30] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][23] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][4] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][26] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][7] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][24] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][26] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][31] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][29] ,
    \\configuration_pci_err_data_reg[23] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][26] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][25] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][23] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][5] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][10] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][31] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][2] ,
    \\configuration_wb_err_addr_reg[17] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][25] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][9] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][6] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][24] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][8] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][17] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][31] ,
    \\configuration_pci_err_data_reg[24] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][33] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][9] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][18] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][21] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][19] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][33] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][10] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][15] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][3] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][15] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][14] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][34] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][11] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][12] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][34] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][13] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][8] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][19] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][25] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][17] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][30] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][5] ,
    \\configuration_pci_err_data_reg[26] ,
    \\configuration_pci_err_data_reg[27] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][34] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][35] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][28] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][35] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][38] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][28] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][16] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][26] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][27] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][10] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][7] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][8] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][18] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][18] ,
    \\configuration_pci_err_addr_reg[7] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][20] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][38] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][14] ,
    \\configuration_pci_err_addr_reg[9] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][12] ,
    \\configuration_pci_err_data_reg[18] ,
    \\configuration_pci_err_data_reg[1] ,
    \\configuration_pci_err_data_reg[20] ,
    \\configuration_pci_err_data_reg[22] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][10] ,
    \\configuration_pci_err_data_reg[14] ,
    \\configuration_pci_err_cs_bit31_24_reg[24] ,
    \\configuration_pci_err_data_reg[16] ,
    \\configuration_pci_err_cs_bit31_24_reg[25] ,
    \\configuration_pci_err_data_reg[10] ,
    \\configuration_pci_err_data_reg[12] ,
    \\configuration_pci_err_cs_bit31_24_reg[26] ,
    \\configuration_pci_err_cs_bit31_24_reg[27] ,
    \\configuration_pci_err_addr_reg[3] ,
    \\configuration_pci_err_addr_reg[10] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][5] ,
    \\configuration_wb_err_addr_reg[21] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][38] ,
    \\configuration_pci_err_addr_reg[5] ,
    \\configuration_pci_err_addr_reg[30] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][11] ,
    \\configuration_pci_err_addr_reg[27] ,
    \\configuration_pci_err_addr_reg[29] ,
    \\configuration_pci_err_addr_reg[25] ,
    \\configuration_pci_err_addr_reg[1] ,
    \\configuration_pci_err_addr_reg[23] ,
    \\configuration_pci_err_addr_reg[24] ,
    \\configuration_pci_err_addr_reg[21] ,
    \\configuration_pci_err_addr_reg[13] ,
    \\configuration_pci_err_addr_reg[18] ,
    \\configuration_pci_err_addr_reg[17] ,
    \\configuration_pci_err_addr_reg[14] ,
    \\configuration_pci_err_addr_reg[16] ,
    \\configuration_pci_err_cs_bit31_24_reg[31] ,
    \\wishbone_slave_unit_pci_initiator_if_read_count_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][3] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][25] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][33] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][31] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][2] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][24] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][13] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][21] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][26] ,
    \\configuration_wb_err_addr_reg[9] ,
    \\configuration_wb_err_addr_reg[5] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][30] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][30] ,
    \\configuration_wb_err_addr_reg[3] ,
    \\configuration_wb_err_addr_reg[23] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][27] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][30] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][28] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][29] ,
    \\configuration_wb_err_addr_reg[30] ,
    \\configuration_wb_err_addr_reg[29] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][19] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][35] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][16] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][28] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][17] ,
    \\configuration_wb_err_addr_reg[25] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][2] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][3] ,
    \\configuration_wb_err_addr_reg[27] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][38] ,
    \\pci_target_unit_fifos_pciw_inTransactionCount_reg[0] ,
    \\pci_target_unit_fifos_inGreyCount_reg[1] ,
    pci_target_unit_del_sync_comp_rty_exp_reg_reg,
    \\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2] ,
    configuration_set_pci_err_cs_bit8_reg,
    wishbone_slave_unit_pci_initiator_if_del_write_req_reg,
    pci_target_unit_wishbone_master_wb_read_done_out_reg,
    pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0] ,
    pci_target_unit_del_sync_req_done_reg_reg,
    \\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1] ,
    \\pci_target_unit_pci_target_if_strd_address_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1] ,
    wishbone_slave_unit_pci_initiator_sm_timeout_reg,
    \\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][39] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][39] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][39] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][39] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][39] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][39] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][39] ,
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][39] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[2] ,
    pci_target_unit_pci_target_sm_wr_to_fifo_reg,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[15] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[2] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[2] ,
    pci_target_unit_del_sync_req_comp_pending_reg,
    wishbone_slave_unit_pci_initiator_sm_transfer_reg,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[1] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[1] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[14] ,
    wishbone_slave_unit_del_sync_comp_rty_exp_reg_reg,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2] ,
    parity_checker_check_for_serr_on_second_reg,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[1] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[1] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[0] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[12] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[1] ,
    \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[3] ,
    i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg,
    pci_target_unit_pci_target_if_target_rd_reg,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[11] ,
    pci_target_unit_pci_target_sm_rd_from_fifo_reg,
    pci_resets_and_interrupts_inta_en_out_reg,
    \\pci_target_unit_pci_target_if_norm_bc_reg[0] ,
    \\pci_target_unit_pci_target_if_strd_address_reg[3] ,
    pci_target_unit_wishbone_master_retried_reg,
    pci_target_unit_wishbone_master_pcir_fifo_wenable_out_reg,
    pci_target_unit_pci_target_sm_rw_cbe0_reg,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[10] ,
    \\pci_target_unit_del_sync_be_out_reg[0] ,
    \\input_register_pci_cbe_reg_out_reg[0] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[8] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[13] ,
    wishbone_slave_unit_pci_initiator_if_last_transfered_reg,
    \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[0] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[7] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[9] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[4] ,
    \\pci_target_unit_pci_target_if_strd_address_reg[1] ,
    \\pci_target_unit_pci_target_if_strd_address_reg[8] ,
    \\pci_target_unit_pci_target_if_strd_address_reg[6] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[6] ,
    pci_target_unit_pci_target_sm_cnf_progress_reg,
    wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[3] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[0] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[1] ,
    wishbone_slave_unit_pci_initiator_if_rdy_out_reg,
    \\pci_target_unit_pci_target_if_norm_address_reg[1] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[2] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[3] ,
    \\pci_target_unit_pci_target_if_norm_bc_reg[1] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_control_out_reg[1] ,
    \\pci_target_unit_pci_target_if_strd_address_reg[4] ,
    \\pci_target_unit_pci_target_if_strd_address_reg[7] ,
    \\pci_target_unit_pci_target_if_strd_address_reg[9] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[5] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[1] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[6] ,
    \\pci_target_unit_pci_target_if_strd_address_reg[5] ,
    \\pci_target_unit_del_sync_comp_cycle_count_reg[0] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[2] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[11] ,
    \\pci_target_unit_del_sync_addr_out_reg[22] ,
    \\pci_target_unit_del_sync_addr_out_reg[21] ,
    \\pci_target_unit_del_sync_bc_out_reg[1] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[16] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[22] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[23] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[24] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[25] ,
    \\pci_target_unit_del_sync_addr_out_reg[16] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[17] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[10] ,
    \\pci_target_unit_del_sync_be_out_reg[1] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[30] ,
    \\input_register_pci_cbe_reg_out_reg[3] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[14] ,
    \\input_register_pci_cbe_reg_out_reg[2] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[28] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[27] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[13] ,
    \\pci_target_unit_pci_target_if_norm_bc_reg[3] ,
    \\pci_target_unit_pci_target_if_norm_bc_reg[2] ,
    \\pci_target_unit_del_sync_addr_out_reg[2] ,
    wishbone_slave_unit_pci_initiator_sm_mabort1_reg,
    \\pci_target_unit_del_sync_addr_out_reg[26] ,
    \\pci_target_unit_del_sync_addr_out_reg[25] ,
    \\pci_target_unit_del_sync_addr_out_reg[24] ,
    \\pci_target_unit_del_sync_addr_out_reg[23] ,
    \\pci_target_unit_del_sync_addr_out_reg[28] ,
    \\pci_target_unit_del_sync_addr_out_reg[20] ,
    pci_target_unit_del_sync_burst_out_reg,
    \\pci_target_unit_del_sync_addr_out_reg[4] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[5] ,
    \\pci_target_unit_del_sync_addr_out_reg[7] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[21] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[12] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[31] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[26] ,
    input_register_pci_trdy_reg_out_reg,
    \\pci_target_unit_pci_target_if_norm_address_reg[15] ,
    \\pci_target_unit_del_sync_addr_out_reg[27] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[13] ,
    \\pci_target_unit_del_sync_addr_out_reg[9] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[21] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[3] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[20] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[27] ,
    \\pci_target_unit_del_sync_addr_out_reg[31] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[8] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[4] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[6] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[1] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[29] ,
    \\input_register_pci_cbe_reg_out_reg[1] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[30] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[26] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[22] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[18] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[12] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[29] ,
    \\pci_target_unit_del_sync_be_out_reg[2] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[20] ,
    \\pci_target_unit_del_sync_addr_out_reg[1] ,
    \\pci_target_unit_del_sync_addr_out_reg[14] ,
    \\pci_target_unit_del_sync_addr_out_reg[6] ,
    \\pci_target_unit_del_sync_addr_out_reg[11] ,
    \\pci_target_unit_del_sync_be_out_reg[3] ,
    wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg,
    \\pci_target_unit_del_sync_addr_out_reg[19] ,
    \\pci_target_unit_del_sync_addr_out_reg[15] ,
    \\pci_target_unit_del_sync_addr_out_reg[30] ,
    \\pci_target_unit_del_sync_addr_out_reg[8] ,
    \\pci_target_unit_del_sync_addr_out_reg[3] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[19] ,
    \\pci_target_unit_del_sync_addr_out_reg[13] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[18] ,
    \\pci_target_unit_del_sync_addr_out_reg[12] ,
    \\pci_target_unit_del_sync_addr_out_reg[10] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0] ,
    pci_target_unit_pci_target_sm_state_backoff_reg_reg,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[10] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[11] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[16] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[19] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[23] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[28] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[2] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[2] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[3] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[5] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[7] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[9] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[31] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[24] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[14] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[15] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[25] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[17] ,
    \\pci_target_unit_del_sync_bc_out_reg[3] ,
    \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[2] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[9] ,
    \\pci_target_unit_del_sync_addr_out_reg[5] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[4] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[0] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[8] ,
    \\pci_target_unit_pci_target_if_strd_address_reg[0] ,
    \\pci_target_unit_pci_target_if_norm_address_reg[7] ,
    \\pci_target_unit_del_sync_bc_out_reg[0] ,
    \\pci_target_unit_del_sync_bc_out_reg[2] ,
    \\pci_target_unit_del_sync_addr_out_reg[29] ,
    \\pci_target_unit_del_sync_addr_out_reg[18] ,
    \\pci_target_unit_del_sync_addr_out_reg[0] ,
    \\pci_target_unit_del_sync_addr_out_reg[17] ,
    input_register_pci_frame_reg_out_reg,
    input_register_pci_devsel_reg_out_reg, pci_io_mux_irdy_iob_dat_out_reg,
    input_register_pci_irdy_reg_out_reg, output_backup_irdy_out_reg,
    \\wishbone_slave_unit_del_sync_rty_exp_back_prop_sync_sync_data_out_reg[0] ,
    pci_target_unit_del_sync_req_req_pending_reg,
    input_register_pci_stop_reg_out_reg,
    \\configuration_sync_cache_lsize_to_wb_bits_reg[8] ,
    configuration_interrupt_out_reg, pci_io_mux_req_iob_dat_out_reg,
    \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[3] ,
    pci_target_unit_pci_target_sm_state_transfere_reg_reg,
    pci_target_unit_pci_target_sm_previous_frame_reg,
    \\input_register_pci_ad_reg_out_reg[7] ,
    \\input_register_pci_ad_reg_out_reg[17] ,
    \\input_register_pci_ad_reg_out_reg[30] ,
    \\input_register_pci_ad_reg_out_reg[16] ,
    \\input_register_pci_ad_reg_out_reg[28] ,
    \\input_register_pci_ad_reg_out_reg[0] ,
    \\configuration_int_pin_sync_sync_data_out_reg[0] ,
    \\input_register_pci_ad_reg_out_reg[24] ,
    \\input_register_pci_ad_reg_out_reg[10] ,
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[6] ,
    \\input_register_pci_ad_reg_out_reg[12] ,
    \\input_register_pci_ad_reg_out_reg[3] ,
    \\input_register_pci_ad_reg_out_reg[13] ,
    parity_checker_master_perr_report_reg,
    \\input_register_pci_ad_reg_out_reg[4] ,
    \\input_register_pci_ad_reg_out_reg[9] ,
    \\input_register_pci_ad_reg_out_reg[14] ,
    pci_target_unit_del_sync_comp_done_reg_clr_reg,
    configuration_wb_init_complete_out_reg,
    \\input_register_pci_ad_reg_out_reg[29] ,
    \\input_register_pci_ad_reg_out_reg[25] ,
    parity_checker_frame_dec2_reg,
    \\input_register_pci_ad_reg_out_reg[15] ,
    \\input_register_pci_ad_reg_out_reg[23] ,
    \\input_register_pci_ad_reg_out_reg[20] ,
    wishbone_slave_unit_del_sync_req_rty_exp_clr_reg,
    \\input_register_pci_ad_reg_out_reg[26] ,
    \\input_register_pci_ad_reg_out_reg[31] ,
    \\input_register_pci_ad_reg_out_reg[6] ,
    configuration_init_complete_reg, input_register_pci_idsel_reg_out_reg,
    \\input_register_pci_ad_reg_out_reg[21] ,
    \\input_register_pci_ad_reg_out_reg[1] ,
    \\input_register_pci_ad_reg_out_reg[18] ,
    \\input_register_pci_ad_reg_out_reg[22] ,
    \\input_register_pci_ad_reg_out_reg[2] ,
    pci_target_unit_pci_target_sm_read_completed_reg_reg,
    \\input_register_pci_ad_reg_out_reg[11] ,
    \\input_register_pci_ad_reg_out_reg[5] ,
    \\input_register_pci_ad_reg_out_reg[8] ,
    \\input_register_pci_ad_reg_out_reg[19] ,
    \\input_register_pci_ad_reg_out_reg[27] ,
    parity_checker_frame_and_irdy_en_prev_prev_reg,
    wishbone_slave_unit_del_sync_comp_done_reg_main_reg,
    pci_target_unit_del_sync_comp_rty_exp_clr_reg,
    configuration_pci_err_cs_bit8_reg, \\configuration_isr_bit2_0_reg[2] ,
    \\configuration_isr_bit2_0_reg[0] ,
    wishbone_slave_unit_pci_initiator_if_write_req_int_reg,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[0] ,
    \\configuration_i_wb_init_complete_sync_sync_data_out_reg[0] ,
    configuration_sync_isr_2_sync_del_bit_reg,
    pci_io_mux_req_iob_en_out_reg,
    pci_target_unit_del_sync_req_rty_exp_reg_reg,
    configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg,
    configuration_sync_isr_2_delayed_bckp_bit_reg,
    wishbone_slave_unit_del_sync_req_comp_pending_sample_reg,
    \\configuration_sync_cache_lsize_to_wb_bits_reg[3] ,
    pci_target_unit_del_sync_req_comp_pending_sample_reg,
    \\pci_target_unit_del_sync_req_sync_sync_data_out_reg[0] ,
    pci_target_unit_del_sync_comp_done_reg_main_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0] ,
    pci_io_mux_irdy_iob_en_out_reg,
    \\pci_target_unit_del_sync_rty_exp_back_prop_sync_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1] ,
    \\wishbone_slave_unit_del_sync_req_sync_sync_data_out_reg[0] ,
    wishbone_slave_unit_pci_initiator_sm_mabort2_reg,
    \\wishbone_slave_unit_del_sync_done_sync_sync_data_out_reg[0] ,
    pci_target_unit_del_sync_comp_flush_out_reg,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0] ,
    wishbone_slave_unit_del_sync_comp_flush_out_reg,
    pci_target_unit_pci_target_sm_bckp_trdy_reg_reg,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3] ,
    configuration_sync_pci_err_cs_8_sync_del_bit_reg,
    parity_checker_frame_and_irdy_en_prev_reg,
    \\configuration_isr_bit0_sync_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[2] ,
    \\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[1] ,
    \\configuration_pci_err_cs_bits_sync_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[3] ,
    \\pci_target_unit_fifos_wb_clk_inGreyCount_reg[0] ,
    \\pci_target_unit_fifos_wb_clk_inGreyCount_reg[1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[2] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[1] ,
    \\configuration_isr_bit2_sync_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[1] ,
    \\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[0] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[0] ,
    output_backup_irdy_en_out_reg,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[3] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1] ,
    \\wishbone_slave_unit_del_sync_comp_sync_sync_data_out_reg[0] ,
    \\pci_target_unit_del_sync_comp_sync_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[1] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[1] ,
    \\pci_target_unit_del_sync_rty_exp_sync_sync_data_out_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2] ,
    \\configuration_sync_isr_2_delete_sync_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[2] ,
    \\pci_target_unit_del_sync_done_sync_sync_data_out_reg[0] ,
    pci_target_unit_del_sync_req_rty_exp_clr_reg,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[2] ,
    configuration_rst_inactive_reg,
    \\configuration_sync_cache_lsize_to_wb_bits_reg[2] ,
    \\configuration_sync_cache_lsize_to_wb_bits_reg[4] ,
    \\configuration_sync_cache_lsize_to_wb_bits_reg[7] ,
    \\configuration_sync_cache_lsize_to_wb_bits_reg[5] ,
    configuration_sync_command_bit_reg,
    \\configuration_sync_cache_lsize_to_wb_bits_reg[6] ,
    configuration_sync_isr_2_sync_bckp_bit_reg,
    wishbone_slave_unit_del_sync_req_rty_exp_reg_reg,
    configuration_sync_pci_err_cs_8_sync_bckp_bit_reg,
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg[1] ,
    \\wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[2] ,
    pci_target_unit_wishbone_master_burst_chopped_delayed_reg,
    \\wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[1] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[2] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg[2] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[1] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[3] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[3] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[1] ,
    \\pci_target_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[1] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg[0] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[0] ,
    \\pci_target_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[2] ,
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[2] ,
    \\configuration_sync_pci_err_cs_8_delete_sync_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[18] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[31] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[3] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[4] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[25] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[6] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[16] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[11] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[2] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[1] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[15] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[14] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg[0] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[2] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[13] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[11] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[10] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg[2] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[15] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[8] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[0] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[6] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[21] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[25] ,
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[0] ,
    \\configuration_sync_isr_2_clear_delete_sync_sync_data_out_reg[0] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[19] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[30] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[27] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[29] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[3] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[19] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[23] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[22] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[28] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[24] ,
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[4] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[2] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[5] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[4] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[13] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[8] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[16] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[17] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[1] ,
    configuration_rst_inactive_sync_reg,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[26] ,
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[5] ,
    configuration_sync_isr_2_delayed_del_bit_reg,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[22] ,
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[2] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[1] ,
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg[1] ,
    \\wishbone_slave_unit_del_sync_rty_exp_sync_sync_data_out_reg[0] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[23] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[20] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[12] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[12] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[21] ,
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[7] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[20] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[26] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[9] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[24] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[7] ,
    \\configuration_command_bit_sync_sync_data_out_reg[0] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[0] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[14] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[31] ,
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[1] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[0] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[10] ,
    \\configuration_sync_pci_err_cs_8_clear_delete_sync_sync_data_out_reg[0] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[3] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[18] ,
    wishbone_slave_unit_del_sync_comp_done_reg_clr_reg,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[27] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[28] ,
    configuration_sync_pci_err_cs_8_delayed_del_bit_reg,
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[3] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[5] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[29] ,
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[2] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[17] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[9] ,
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[30] ;
  wire \new_[3728]_ , new_configuration_rst_inactive_sync_reg_in_,
    \new_[3738]_ , \new_[3746]_ , \new_[3747]_ , \new_[3784]_ ,
    \new_[3785]_ , \new_[3786]_ , \new_[3846]_ , \new_[3861]_ ,
    \new_[3862]_ , \new_[3863]_ , \new_[3864]_ , \new_[3865]_ ,
    \new_[3883]_ , \new_[3884]_ , \new_[3885]_ , \new_[3886]_ ,
    \new_[3889]_ , \new_[3893]_ , \new_[3894]_ , \new_[3895]_ ,
    \new_[3896]_ , \new_[3897]_ , \new_[3898]_ , \new_[3899]_ ,
    \new_[3900]_ , \new_[3901]_ , \new_[3902]_ , \new_[3903]_ ,
    \new_[3904]_ , \new_[3905]_ , \new_[3906]_ , \new_[3907]_ ,
    \new_[3908]_ , \new_[3909]_ , \new_[3910]_ , \new_[3911]_ ,
    \new_[3912]_ , \new_[3913]_ , \new_[3914]_ , \new_[3915]_ ,
    \new_[3916]_ , \new_[3917]_ , \new_[3918]_ , \new_[3919]_ ,
    \new_[3921]_ , \new_[3922]_ , \new_[3923]_ , \new_[3924]_ ,
    \new_[3925]_ , \new_[3926]_ , \new_[3927]_ , \new_[3928]_ ,
    \new_[3929]_ , \new_[3930]_ , \new_[3931]_ , \new_[3932]_ ,
    \new_[3933]_ , \new_[3934]_ , \new_[3935]_ , \new_[3936]_ ,
    \new_[3937]_ , \new_[3938]_ , \new_[3939]_ , \new_[3940]_ ,
    \new_[3941]_ , \new_[3942]_ , \new_[3943]_ , \new_[3944]_ ,
    \new_[3945]_ , \new_[3946]_ , \new_[3947]_ , \new_[3948]_ ,
    \new_[3949]_ , \new_[3950]_ , \new_[3951]_ , \new_[3952]_ ,
    \new_[3953]_ , \new_[3954]_ , \new_[3955]_ , \new_[3956]_ ,
    \new_[3957]_ , \new_[3958]_ , \new_[3959]_ , \new_[3960]_ ,
    \new_[3961]_ , \new_[3962]_ , \new_[3963]_ , \new_[3964]_ ,
    \new_[3965]_ , \new_[3966]_ , \new_[3967]_ , \new_[3968]_ ,
    \new_[3969]_ , \new_[3970]_ , \new_[3971]_ , \new_[3972]_ ,
    \new_[3973]_ , \new_[3974]_ , \new_[3976]_ , \new_[3977]_ ,
    \new_[3978]_ , \new_[3983]_ , \new_[3984]_ , \new_[3985]_ ,
    \new_[3986]_ , \new_[3987]_ , \new_[3988]_ , \new_[3989]_ ,
    \new_[3990]_ , \new_[3991]_ , \new_[3992]_ , \new_[3993]_ ,
    \new_[3994]_ , \new_[3995]_ , \new_[3997]_ , \new_[3998]_ ,
    \new_[3999]_ , \new_[4000]_ , \new_[4001]_ , \new_[4002]_ ,
    \new_[4003]_ , \new_[4004]_ , \new_[4005]_ , \new_[4006]_ ,
    \new_[4007]_ , \new_[4008]_ , \new_[4009]_ , \new_[4010]_ ,
    \new_[4011]_ , \new_[4012]_ , \new_[4013]_ , \new_[4014]_ ,
    \new_[4015]_ , \new_[4016]_ , \new_[4017]_ , \new_[4018]_ ,
    \new_[4019]_ , \new_[4020]_ , \new_[4021]_ , \new_[4022]_ ,
    \new_[4023]_ , \new_[4024]_ , \new_[4025]_ , \new_[4026]_ ,
    \new_[4027]_ , \new_[4028]_ , \new_[4029]_ , \new_[4030]_ ,
    \new_[4031]_ , \new_[4032]_ , \new_[4033]_ , \new_[4034]_ ,
    \new_[4035]_ , \new_[4036]_ , \new_[4037]_ , \new_[4038]_ ,
    \new_[4040]_ , \new_[4041]_ , \new_[4042]_ , \new_[4045]_ ,
    \new_[4046]_ , \new_[4047]_ , \new_[4048]_ , \new_[4049]_ ,
    \new_[4050]_ , \new_[4051]_ , \new_[4052]_ , \new_[4053]_ ,
    \new_[4054]_ , \new_[4055]_ , \new_[4056]_ , \new_[4057]_ ,
    \new_[4058]_ , \new_[4059]_ , \new_[4060]_ , \new_[4061]_ ,
    \new_[4062]_ , \new_[4063]_ , \new_[4064]_ , \new_[4065]_ ,
    \new_[4066]_ , \new_[4067]_ , \new_[4068]_ , \new_[4069]_ ,
    \new_[4070]_ , \new_[4071]_ , \new_[4072]_ , \new_[4073]_ ,
    \new_[4074]_ , \new_[4075]_ , \new_[4076]_ , \new_[4077]_ ,
    \new_[4078]_ , \new_[4079]_ , \new_[4080]_ , \new_[4081]_ ,
    \new_[4082]_ , \new_[4084]_ , \new_[4088]_ , \new_[4089]_ ,
    \new_[4090]_ , \new_[4092]_ , \new_[4094]_ , \new_[4095]_ ,
    \new_[4096]_ , \new_[4122]_ , \new_[4130]_ , \new_[4133]_ ,
    \new_[4134]_ , \new_[4136]_ , \new_[4137]_ , \new_[4141]_ ,
    \new_[4142]_ , \new_[4143]_ , \new_[4144]_ , \new_[4145]_ ,
    \new_[4146]_ , \new_[4147]_ , \new_[4148]_ , \new_[4149]_ ,
    \new_[4150]_ , \new_[4151]_ , \new_[4152]_ , \new_[4153]_ ,
    \new_[4154]_ , \new_[4155]_ , \new_[4156]_ , \new_[4157]_ ,
    \new_[4158]_ , \new_[4159]_ , \new_[4160]_ , \new_[4161]_ ,
    \new_[4162]_ , \new_[4163]_ , \new_[4164]_ , \new_[4165]_ ,
    \new_[4166]_ , \new_[4167]_ , \new_[4168]_ , \new_[4169]_ ,
    \new_[4170]_ , \new_[4171]_ , \new_[4172]_ , \new_[4173]_ ,
    \new_[4174]_ , \new_[4175]_ , \new_[4178]_ , \new_[4180]_ ,
    \new_[4181]_ , \new_[4182]_ , \new_[4183]_ , \new_[4184]_ ,
    \new_[4185]_ , \new_[4186]_ , \new_[4187]_ , \new_[4188]_ ,
    \new_[4189]_ , \new_[4190]_ , \new_[4191]_ , \new_[4192]_ ,
    \new_[4210]_ , \new_[4211]_ , \new_[4212]_ , \new_[4213]_ ,
    \new_[4214]_ , \new_[4215]_ , \new_[4216]_ , \new_[4217]_ ,
    \new_[4218]_ , \new_[4226]_ , \new_[4228]_ , \new_[4229]_ ,
    \new_[4230]_ , \new_[4234]_ , \new_[4235]_ , \new_[4236]_ ,
    \new_[4237]_ , \new_[4238]_ , \new_[4239]_ , \new_[4240]_ ,
    \new_[4241]_ , \new_[4242]_ , \new_[4243]_ , \new_[4244]_ ,
    \new_[4245]_ , \new_[4246]_ , \new_[4247]_ , \new_[4248]_ ,
    \new_[4249]_ , \new_[4250]_ , \new_[4251]_ , \new_[4252]_ ,
    \new_[4253]_ , \new_[4254]_ , \new_[4255]_ , \new_[4256]_ ,
    \new_[4257]_ , \new_[4258]_ , \new_[4259]_ , \new_[4260]_ ,
    \new_[4261]_ , \new_[4264]_ , \new_[4265]_ , \new_[4267]_ ,
    \new_[4268]_ , \new_[4270]_ , \new_[4272]_ , \new_[4273]_ ,
    \new_[4274]_ , \new_[4275]_ , \new_[4276]_ , \new_[4278]_ ,
    \new_[4279]_ , \new_[4280]_ , \new_[4281]_ , \new_[4282]_ ,
    \new_[4283]_ , \new_[4284]_ , \new_[4285]_ , \new_[4286]_ ,
    \new_[4287]_ , \new_[4288]_ , \new_[4289]_ , \new_[4290]_ ,
    \new_[4291]_ , \new_[4292]_ , \new_[4293]_ , \new_[4294]_ ,
    \new_[4295]_ , \new_[4296]_ , \new_[4297]_ , \new_[4298]_ ,
    \new_[4299]_ , \new_[4300]_ , \new_[4301]_ , \new_[4302]_ ,
    \new_[4303]_ , \new_[4304]_ , \new_[4305]_ , \new_[4306]_ ,
    \new_[4307]_ , \new_[4308]_ , \new_[4309]_ , \new_[4310]_ ,
    \new_[4311]_ , \new_[4312]_ , \new_[4313]_ , \new_[4314]_ ,
    \new_[4315]_ , \new_[4316]_ , \new_[4317]_ , \new_[4318]_ ,
    \new_[4319]_ , \new_[4320]_ , \new_[4321]_ , \new_[4322]_ ,
    \new_[4323]_ , \new_[4324]_ , \new_[4325]_ , \new_[4326]_ ,
    \new_[4327]_ , \new_[4328]_ , \new_[4329]_ , \new_[4330]_ ,
    \new_[4331]_ , \new_[4332]_ , \new_[4333]_ , \new_[4334]_ ,
    \new_[4335]_ , \new_[4336]_ , \new_[4337]_ , \new_[4338]_ ,
    \new_[4339]_ , \new_[4340]_ , \new_[4341]_ , \new_[4342]_ ,
    \new_[4343]_ , \new_[4345]_ , \new_[4346]_ , \new_[4347]_ ,
    \new_[4354]_ , \new_[4355]_ , \new_[4356]_ , \new_[4407]_ ,
    \new_[4408]_ , \new_[4409]_ , \new_[4410]_ , \new_[4411]_ ,
    \new_[4412]_ , \new_[4413]_ , \new_[4414]_ , \new_[4415]_ ,
    \new_[4416]_ , \new_[4417]_ , \new_[4418]_ , \new_[4419]_ ,
    \new_[4420]_ , \new_[4421]_ , \new_[4422]_ , \new_[4423]_ ,
    \new_[4424]_ , \new_[4425]_ , \new_[4426]_ , \new_[4427]_ ,
    \new_[4428]_ , \new_[4429]_ , \new_[4430]_ , \new_[4431]_ ,
    \new_[4432]_ , \new_[4433]_ , \new_[4434]_ , \new_[4435]_ ,
    \new_[4436]_ , \new_[4437]_ , \new_[4438]_ , \new_[4439]_ ,
    \new_[4440]_ , \new_[4441]_ , \new_[4442]_ , \new_[4443]_ ,
    \new_[4444]_ , \new_[4445]_ , \new_[4446]_ , \new_[4447]_ ,
    \new_[4448]_ , \new_[4449]_ , \new_[4450]_ , \new_[4451]_ ,
    \new_[4452]_ , \new_[4453]_ , \new_[4454]_ , \new_[4455]_ ,
    \new_[4456]_ , \new_[4458]_ , \new_[4459]_ , \new_[4460]_ ,
    \new_[4461]_ , \new_[4462]_ , \new_[4463]_ , \new_[4464]_ ,
    \new_[4465]_ , \new_[4466]_ , \new_[4467]_ , \new_[4468]_ ,
    \new_[4469]_ , \new_[4470]_ , \new_[4471]_ , \new_[4472]_ ,
    \new_[4473]_ , \new_[4474]_ , \new_[4475]_ , \new_[4476]_ ,
    \new_[4477]_ , \new_[4478]_ , \new_[4479]_ , \new_[4480]_ ,
    \new_[4481]_ , \new_[4482]_ , \new_[4483]_ , \new_[4484]_ ,
    \new_[4485]_ , \new_[4486]_ , \new_[4487]_ , \new_[4488]_ ,
    \new_[4489]_ , \new_[4490]_ , \new_[4491]_ , \new_[4492]_ ,
    \new_[4493]_ , \new_[4494]_ , \new_[4495]_ , \new_[4496]_ ,
    \new_[4497]_ , \new_[4498]_ , \new_[4499]_ , \new_[4500]_ ,
    \new_[4501]_ , \new_[4502]_ , \new_[4503]_ , \new_[4504]_ ,
    \new_[4505]_ , \new_[4506]_ , \new_[4507]_ , \new_[4508]_ ,
    \new_[4509]_ , \new_[4510]_ , \new_[4511]_ , \new_[4512]_ ,
    \new_[4513]_ , \new_[4514]_ , \new_[4515]_ , \new_[4516]_ ,
    \new_[4517]_ , \new_[4518]_ , \new_[4519]_ , \new_[4520]_ ,
    \new_[4521]_ , \new_[4522]_ , \new_[4523]_ , \new_[4524]_ ,
    \new_[4525]_ , \new_[4526]_ , \new_[4527]_ , \new_[4528]_ ,
    \new_[4529]_ , \new_[4530]_ , \new_[4531]_ , \new_[4532]_ ,
    \new_[4533]_ , \new_[4534]_ , \new_[4535]_ , \new_[4536]_ ,
    \new_[4537]_ , \new_[4538]_ , \new_[4539]_ , \new_[4540]_ ,
    \new_[4541]_ , \new_[4542]_ , \new_[4543]_ , \new_[4544]_ ,
    \new_[4545]_ , \new_[4546]_ , \new_[4547]_ , \new_[4548]_ ,
    \new_[4549]_ , \new_[4550]_ , \new_[4551]_ , \new_[4552]_ ,
    \new_[4553]_ , \new_[4554]_ , \new_[4555]_ , \new_[4556]_ ,
    \new_[4557]_ , \new_[4558]_ , \new_[4559]_ , \new_[4560]_ ,
    \new_[4561]_ , \new_[4562]_ , \new_[4563]_ , \new_[4564]_ ,
    \new_[4565]_ , \new_[4566]_ , \new_[4567]_ , \new_[4568]_ ,
    \new_[4569]_ , \new_[4570]_ , \new_[4571]_ , \new_[4572]_ ,
    \new_[4573]_ , \new_[4574]_ , \new_[4575]_ , \new_[4576]_ ,
    \new_[4577]_ , \new_[4578]_ , \new_[4579]_ , \new_[4580]_ ,
    \new_[4581]_ , \new_[4582]_ , \new_[4583]_ , \new_[4584]_ ,
    \new_[4585]_ , \new_[4586]_ , \new_[4587]_ , \new_[4588]_ ,
    \new_[4589]_ , \new_[4590]_ , \new_[4591]_ , \new_[4592]_ ,
    \new_[4593]_ , \new_[4596]_ , \new_[4597]_ , \new_[4598]_ ,
    \new_[4599]_ , \new_[4601]_ , \new_[4606]_ , \new_[4609]_ ,
    \new_[4610]_ , \new_[4611]_ , \new_[4612]_ , \new_[4627]_ ,
    \new_[4628]_ , \new_[4629]_ , \new_[4630]_ , \new_[4631]_ ,
    \new_[4632]_ , \new_[4633]_ , \new_[4634]_ , \new_[4635]_ ,
    \new_[4636]_ , \new_[4637]_ , \new_[4638]_ , \new_[4639]_ ,
    \new_[4640]_ , \new_[4641]_ , \new_[4642]_ , \new_[4643]_ ,
    \new_[4644]_ , \new_[4645]_ , \new_[4646]_ , \new_[4647]_ ,
    \new_[4648]_ , \new_[4649]_ , \new_[4650]_ , \new_[4651]_ ,
    \new_[4652]_ , \new_[4653]_ , \new_[4654]_ , \new_[4655]_ ,
    \new_[4656]_ , \new_[4657]_ , \new_[4658]_ , \new_[4659]_ ,
    \new_[4660]_ , \new_[4661]_ , \new_[4662]_ , \new_[4663]_ ,
    \new_[4664]_ , \new_[4665]_ , \new_[4666]_ , \new_[4667]_ ,
    \new_[4668]_ , \new_[4669]_ , \new_[4670]_ , \new_[4671]_ ,
    \new_[4672]_ , \new_[4673]_ , \new_[4674]_ , \new_[4675]_ ,
    \new_[4676]_ , \new_[4677]_ , \new_[4678]_ , \new_[4679]_ ,
    \new_[4680]_ , \new_[4681]_ , \new_[4682]_ , \new_[4683]_ ,
    \new_[4684]_ , \new_[4685]_ , \new_[4686]_ , \new_[4687]_ ,
    \new_[4688]_ , \new_[4689]_ , \new_[4690]_ , \new_[4691]_ ,
    \new_[4692]_ , \new_[4693]_ , \new_[4694]_ , \new_[4695]_ ,
    \new_[4696]_ , \new_[4697]_ , \new_[4698]_ , \new_[4699]_ ,
    \new_[4700]_ , \new_[4701]_ , \new_[4702]_ , \new_[4703]_ ,
    \new_[4704]_ , \new_[4705]_ , \new_[4706]_ , \new_[4707]_ ,
    \new_[4708]_ , \new_[4709]_ , \new_[4710]_ , \new_[4711]_ ,
    \new_[4712]_ , \new_[4713]_ , \new_[4714]_ , \new_[4715]_ ,
    \new_[4716]_ , \new_[4717]_ , \new_[4718]_ , \new_[4719]_ ,
    \new_[4720]_ , \new_[4721]_ , \new_[4722]_ , \new_[4723]_ ,
    \new_[4724]_ , \new_[4725]_ , \new_[4726]_ , \new_[4727]_ ,
    \new_[4728]_ , \new_[4729]_ , \new_[4730]_ , \new_[4731]_ ,
    \new_[4732]_ , \new_[4733]_ , \new_[4734]_ , \new_[4735]_ ,
    \new_[4736]_ , \new_[4737]_ , \new_[4738]_ , \new_[4739]_ ,
    \new_[4740]_ , \new_[4741]_ , \new_[4742]_ , \new_[4743]_ ,
    \new_[4744]_ , \new_[4745]_ , \new_[4746]_ , \new_[4747]_ ,
    \new_[4748]_ , \new_[4749]_ , \new_[4750]_ , \new_[4751]_ ,
    \new_[4752]_ , \new_[4753]_ , \new_[4754]_ , \new_[4755]_ ,
    \new_[4756]_ , \new_[4757]_ , \new_[4758]_ , \new_[4759]_ ,
    \new_[4760]_ , \new_[4761]_ , \new_[4762]_ , \new_[4763]_ ,
    \new_[4764]_ , \new_[4765]_ , \new_[4766]_ , \new_[4767]_ ,
    \new_[4768]_ , \new_[4769]_ , \new_[4770]_ , \new_[4771]_ ,
    \new_[4772]_ , \new_[4773]_ , \new_[4774]_ , \new_[4775]_ ,
    \new_[4777]_ , \new_[4778]_ , \new_[4779]_ , \new_[4780]_ ,
    \new_[4781]_ , \new_[4782]_ , \new_[4783]_ , \new_[4784]_ ,
    \new_[4785]_ , \new_[4786]_ , \new_[4787]_ , \new_[4788]_ ,
    \new_[4790]_ , \new_[4792]_ , \new_[4798]_ , \new_[4799]_ ,
    \new_[4800]_ , \new_[4801]_ , \new_[4802]_ , \new_[4803]_ ,
    \new_[4804]_ , \new_[4805]_ , \new_[4806]_ , \new_[4807]_ ,
    \new_[4808]_ , \new_[4809]_ , \new_[4810]_ , \new_[4811]_ ,
    \new_[4812]_ , \new_[4813]_ , \new_[4814]_ , \new_[4815]_ ,
    \new_[4816]_ , \new_[4817]_ , \new_[4818]_ , \new_[4819]_ ,
    \new_[4820]_ , \new_[4821]_ , \new_[4822]_ , \new_[4823]_ ,
    \new_[4824]_ , \new_[4825]_ , \new_[4826]_ , \new_[4827]_ ,
    \new_[4828]_ , \new_[4829]_ , \new_[4830]_ , \new_[4831]_ ,
    \new_[4832]_ , \new_[4833]_ , \new_[4834]_ , \new_[4835]_ ,
    \new_[4836]_ , \new_[4837]_ , \new_[4838]_ , \new_[4839]_ ,
    \new_[4840]_ , \new_[4841]_ , \new_[4842]_ , \new_[4843]_ ,
    \new_[4844]_ , \new_[4845]_ , \new_[4846]_ , \new_[4847]_ ,
    \new_[4848]_ , \new_[4849]_ , \new_[4850]_ , \new_[4851]_ ,
    \new_[4852]_ , \new_[4853]_ , \new_[4854]_ , \new_[4855]_ ,
    \new_[4856]_ , \new_[4857]_ , \new_[4858]_ , \new_[4859]_ ,
    \new_[4860]_ , \new_[4861]_ , \new_[4862]_ , \new_[4863]_ ,
    \new_[4864]_ , \new_[4865]_ , \new_[4866]_ , \new_[4867]_ ,
    \new_[4868]_ , \new_[4869]_ , \new_[4871]_ , \new_[4872]_ ,
    \new_[4873]_ , \new_[4875]_ , \new_[4876]_ , \new_[4896]_ ,
    \new_[4899]_ , \new_[4900]_ , \new_[4903]_ , \new_[4905]_ ,
    \new_[4907]_ , \new_[4908]_ , \new_[4909]_ , \new_[4911]_ ,
    \new_[4912]_ , \new_[4913]_ , \new_[4914]_ , \new_[4915]_ ,
    \new_[4916]_ , \new_[4918]_ , \new_[4919]_ , \new_[4920]_ ,
    \new_[4921]_ , \new_[4922]_ , \new_[4926]_ , \new_[4928]_ ,
    \new_[4929]_ , \new_[4930]_ , \new_[4931]_ , \new_[4932]_ ,
    \new_[4933]_ , \new_[4934]_ , \new_[4935]_ , \new_[4936]_ ,
    \new_[4937]_ , \new_[4938]_ , \new_[4939]_ , \new_[4940]_ ,
    \new_[4941]_ , \new_[4942]_ , \new_[4943]_ , \new_[4944]_ ,
    \new_[4945]_ , \new_[4946]_ , \new_[4949]_ , \new_[4950]_ ,
    \new_[4951]_ , \new_[4952]_ , \new_[4953]_ , \new_[4954]_ ,
    \new_[4956]_ , \new_[4957]_ , \new_[4958]_ , \new_[4959]_ ,
    \new_[4960]_ , \new_[4961]_ , \new_[4962]_ , \new_[4963]_ ,
    \new_[4964]_ , \new_[4965]_ , \new_[4966]_ , \new_[4967]_ ,
    \new_[4968]_ , \new_[4969]_ , \new_[4970]_ , \new_[4971]_ ,
    \new_[4972]_ , \new_[4973]_ , \new_[4974]_ , \new_[4975]_ ,
    \new_[4976]_ , \new_[4977]_ , \new_[4978]_ , \new_[4979]_ ,
    \new_[4980]_ , \new_[4981]_ , \new_[4982]_ , \new_[4983]_ ,
    \new_[4984]_ , \new_[4986]_ , \new_[4987]_ , \new_[4988]_ ,
    \new_[4989]_ , \new_[4990]_ , \new_[4991]_ , \new_[4992]_ ,
    \new_[4993]_ , \new_[4995]_ , \new_[4997]_ , \new_[4998]_ ,
    \new_[4999]_ , \new_[5002]_ , \new_[5003]_ , \new_[5004]_ ,
    \new_[5005]_ , \new_[5006]_ , \new_[5008]_ , \new_[5009]_ ,
    \new_[5010]_ , \new_[5011]_ , \new_[5012]_ , \new_[5013]_ ,
    \new_[5014]_ , \new_[5015]_ , \new_[5016]_ , \new_[5017]_ ,
    \new_[5018]_ , \new_[5019]_ , \new_[5020]_ , \new_[5021]_ ,
    \new_[5022]_ , \new_[5023]_ , \new_[5024]_ , \new_[5025]_ ,
    \new_[5026]_ , \new_[5027]_ , \new_[5028]_ , \new_[5029]_ ,
    \new_[5030]_ , \new_[5031]_ , \new_[5032]_ , \new_[5033]_ ,
    \new_[5034]_ , \new_[5035]_ , \new_[5036]_ , \new_[5037]_ ,
    \new_[5038]_ , \new_[5039]_ , \new_[5040]_ , \new_[5041]_ ,
    \new_[5042]_ , \new_[5043]_ , \new_[5044]_ , \new_[5045]_ ,
    \new_[5046]_ , \new_[5047]_ , \new_[5048]_ , \new_[5049]_ ,
    \new_[5050]_ , \new_[5051]_ , \new_[5052]_ , \new_[5053]_ ,
    \new_[5054]_ , \new_[5055]_ , \new_[5056]_ , \new_[5057]_ ,
    \new_[5058]_ , \new_[5059]_ , \new_[5060]_ , \new_[5061]_ ,
    \new_[5062]_ , \new_[5063]_ , \new_[5064]_ , \new_[5066]_ ,
    \new_[5068]_ , \new_[5069]_ , \new_[5072]_ , \new_[5074]_ ,
    \new_[5075]_ , \new_[5078]_ , \new_[5079]_ , \new_[5080]_ ,
    \new_[5081]_ , \new_[5088]_ , \new_[5089]_ , \new_[5090]_ ,
    \new_[5091]_ , \new_[5096]_ , \new_[5097]_ , \new_[5099]_ ,
    \new_[5100]_ , \new_[5101]_ , \new_[5102]_ , \new_[5103]_ ,
    \new_[5104]_ , \new_[5105]_ , \new_[5106]_ , \new_[5107]_ ,
    \new_[5109]_ , \new_[5110]_ , \new_[5112]_ , \new_[5113]_ ,
    \new_[5114]_ , \new_[5115]_ , \new_[5116]_ , \new_[5117]_ ,
    \new_[5118]_ , \new_[5119]_ , \new_[5120]_ , \new_[5121]_ ,
    \new_[5122]_ , \new_[5123]_ , \new_[5124]_ , \new_[5125]_ ,
    \new_[5126]_ , \new_[5127]_ , \new_[5128]_ , \new_[5129]_ ,
    \new_[5130]_ , \new_[5131]_ , \new_[5132]_ , \new_[5133]_ ,
    \new_[5134]_ , \new_[5135]_ , \new_[5136]_ , \new_[5137]_ ,
    \new_[5138]_ , \new_[5139]_ , \new_[5140]_ , \new_[5141]_ ,
    \new_[5142]_ , \new_[5143]_ , \new_[5161]_ , \new_[5163]_ ,
    \new_[5164]_ , \new_[5165]_ , \new_[5166]_ , \new_[5167]_ ,
    \new_[5168]_ , \new_[5169]_ , \new_[5170]_ , \new_[5171]_ ,
    \new_[5172]_ , \new_[5173]_ , \new_[5174]_ , \new_[5191]_ ,
    \new_[5192]_ , \new_[5193]_ , \new_[5194]_ , \new_[5195]_ ,
    \new_[5196]_ , \new_[5197]_ , \new_[5198]_ , \new_[5199]_ ,
    \new_[5200]_ , \new_[5201]_ , \new_[5202]_ , \new_[5203]_ ,
    \new_[5204]_ , \new_[5205]_ , \new_[5206]_ , \new_[5207]_ ,
    \new_[5208]_ , \new_[5209]_ , \new_[5210]_ , \new_[5211]_ ,
    \new_[5212]_ , \new_[5213]_ , \new_[5214]_ , \new_[5215]_ ,
    \new_[5216]_ , \new_[5217]_ , \new_[5218]_ , \new_[5219]_ ,
    \new_[5220]_ , \new_[5225]_ , \new_[5226]_ , \new_[5227]_ ,
    \new_[5273]_ , \new_[5274]_ , \new_[5275]_ , \new_[5276]_ ,
    \new_[5277]_ , \new_[5278]_ , \new_[5279]_ , \new_[5280]_ ,
    \new_[5281]_ , \new_[5282]_ , \new_[5283]_ , \new_[5284]_ ,
    \new_[5285]_ , \new_[5286]_ , \new_[5287]_ , \new_[5288]_ ,
    \new_[5289]_ , \new_[5292]_ , \new_[5295]_ , \new_[5297]_ ,
    \new_[5298]_ , \new_[5299]_ , \new_[5303]_ , \new_[5304]_ ,
    \new_[5305]_ , \new_[5306]_ , \new_[5307]_ , \new_[5308]_ ,
    \new_[5309]_ , \new_[5310]_ , \new_[5311]_ , \new_[5312]_ ,
    \new_[5313]_ , \new_[5314]_ , \new_[5315]_ , \new_[5316]_ ,
    \new_[5317]_ , \new_[5318]_ , \new_[5319]_ , \new_[5320]_ ,
    \new_[5321]_ , \new_[5322]_ , \new_[5323]_ , \new_[5324]_ ,
    \new_[5325]_ , \new_[5326]_ , \new_[5327]_ , \new_[5328]_ ,
    \new_[5329]_ , \new_[5330]_ , \new_[5331]_ , \new_[5332]_ ,
    \new_[5333]_ , \new_[5334]_ , \new_[5335]_ , \new_[5336]_ ,
    \new_[5337]_ , \new_[5338]_ , \new_[5339]_ , \new_[5340]_ ,
    \new_[5341]_ , \new_[5342]_ , \new_[5343]_ , \new_[5344]_ ,
    \new_[5345]_ , \new_[5346]_ , \new_[5347]_ , \new_[5348]_ ,
    \new_[5349]_ , \new_[5350]_ , \new_[5351]_ , \new_[5352]_ ,
    \new_[5353]_ , \new_[5354]_ , \new_[5355]_ , \new_[5356]_ ,
    \new_[5357]_ , \new_[5358]_ , \new_[5359]_ , \new_[5360]_ ,
    \new_[5361]_ , \new_[5362]_ , \new_[5363]_ , \new_[5364]_ ,
    \new_[5365]_ , \new_[5366]_ , \new_[5368]_ , \new_[5369]_ ,
    \new_[5382]_ , \new_[5383]_ , \new_[5384]_ , \new_[5385]_ ,
    \new_[5386]_ , \new_[5387]_ , \new_[5388]_ , \new_[5389]_ ,
    \new_[5390]_ , \new_[5391]_ , \new_[5392]_ , \new_[5393]_ ,
    \new_[5394]_ , \new_[5395]_ , \new_[5396]_ , \new_[5397]_ ,
    \new_[5398]_ , \new_[5399]_ , \new_[5400]_ , \new_[5401]_ ,
    \new_[5402]_ , \new_[5403]_ , \new_[5404]_ , \new_[5405]_ ,
    \new_[5406]_ , \new_[5407]_ , \new_[5408]_ , \new_[5409]_ ,
    \new_[5410]_ , \new_[5411]_ , \new_[5412]_ , \new_[5413]_ ,
    \new_[5414]_ , \new_[5415]_ , \new_[5416]_ , \new_[5417]_ ,
    \new_[5418]_ , \new_[5419]_ , \new_[5420]_ , \new_[5421]_ ,
    \new_[5422]_ , \new_[5423]_ , \new_[5424]_ , \new_[5425]_ ,
    \new_[5426]_ , \new_[5427]_ , \new_[5428]_ , \new_[5429]_ ,
    \new_[5430]_ , \new_[5431]_ , \new_[5432]_ , \new_[5433]_ ,
    \new_[5434]_ , \new_[5435]_ , \new_[5436]_ , \new_[5437]_ ,
    \new_[5438]_ , \new_[5439]_ , \new_[5440]_ , \new_[5441]_ ,
    \new_[5442]_ , \new_[5443]_ , \new_[5444]_ , \new_[5445]_ ,
    \new_[5446]_ , \new_[5447]_ , \new_[5448]_ , \new_[5449]_ ,
    \new_[5450]_ , \new_[5456]_ , \new_[5457]_ , \new_[5458]_ ,
    \new_[5459]_ , \new_[5460]_ , \new_[5461]_ , \new_[5462]_ ,
    \new_[5463]_ , \new_[5464]_ , \new_[5465]_ , \new_[5466]_ ,
    \new_[5467]_ , \new_[5468]_ , \new_[5469]_ , \new_[5470]_ ,
    \new_[5471]_ , \new_[5472]_ , \new_[5473]_ , \new_[5474]_ ,
    \new_[5475]_ , \new_[5476]_ , \new_[5477]_ , \new_[5478]_ ,
    \new_[5479]_ , \new_[5480]_ , \new_[5481]_ , \new_[5482]_ ,
    \new_[5483]_ , \new_[5484]_ , \new_[5485]_ , \new_[5486]_ ,
    \new_[5487]_ , \new_[5488]_ , \new_[5489]_ , \new_[5490]_ ,
    \new_[5491]_ , \new_[5492]_ , \new_[5493]_ , \new_[5494]_ ,
    \new_[5495]_ , \new_[5496]_ , \new_[5497]_ , \new_[5498]_ ,
    \new_[5499]_ , \new_[5500]_ , \new_[5501]_ , \new_[5502]_ ,
    \new_[5503]_ , \new_[5504]_ , \new_[5505]_ , \new_[5506]_ ,
    \new_[5507]_ , \new_[5508]_ , \new_[5509]_ , \new_[5510]_ ,
    \new_[5511]_ , \new_[5512]_ , \new_[5513]_ , \new_[5514]_ ,
    \new_[5515]_ , \new_[5516]_ , \new_[5517]_ , \new_[5518]_ ,
    \new_[5519]_ , \new_[5520]_ , \new_[5521]_ , \new_[5522]_ ,
    \new_[5523]_ , \new_[5524]_ , \new_[5525]_ , \new_[5526]_ ,
    \new_[5527]_ , \new_[5528]_ , \new_[5529]_ , \new_[5530]_ ,
    \new_[5531]_ , \new_[5532]_ , \new_[5533]_ , \new_[5534]_ ,
    \new_[5535]_ , \new_[5536]_ , \new_[5537]_ , \new_[5538]_ ,
    \new_[5539]_ , \new_[5540]_ , \new_[5541]_ , \new_[5542]_ ,
    \new_[5543]_ , \new_[5544]_ , \new_[5545]_ , \new_[5546]_ ,
    \new_[5547]_ , \new_[5548]_ , \new_[5549]_ , \new_[5550]_ ,
    \new_[5551]_ , \new_[5552]_ , \new_[5553]_ , \new_[5554]_ ,
    \new_[5555]_ , \new_[5556]_ , \new_[5557]_ , \new_[5558]_ ,
    \new_[5559]_ , \new_[5560]_ , \new_[5561]_ , \new_[5562]_ ,
    \new_[5563]_ , \new_[5564]_ , \new_[5565]_ , \new_[5566]_ ,
    \new_[5567]_ , \new_[5568]_ , \new_[5569]_ , \new_[5570]_ ,
    \new_[5571]_ , \new_[5572]_ , \new_[5573]_ , \new_[5574]_ ,
    \new_[5575]_ , \new_[5576]_ , \new_[5577]_ , \new_[5578]_ ,
    \new_[5579]_ , \new_[5580]_ , \new_[5581]_ , \new_[5582]_ ,
    \new_[5583]_ , \new_[5584]_ , \new_[5585]_ , \new_[5586]_ ,
    \new_[5587]_ , \new_[5588]_ , \new_[5589]_ , \new_[5590]_ ,
    \new_[5591]_ , \new_[5592]_ , \new_[5593]_ , \new_[5594]_ ,
    \new_[5595]_ , \new_[5596]_ , \new_[5597]_ , \new_[5598]_ ,
    \new_[5599]_ , \new_[5600]_ , \new_[5601]_ , \new_[5602]_ ,
    \new_[5603]_ , \new_[5604]_ , \new_[5605]_ , \new_[5606]_ ,
    \new_[5607]_ , \new_[5626]_ , \new_[5629]_ , \new_[5630]_ ,
    \new_[5631]_ , \new_[5632]_ , \new_[5633]_ , \new_[5634]_ ,
    \new_[5635]_ , \new_[5636]_ , \new_[5637]_ , \new_[5638]_ ,
    \new_[5639]_ , \new_[5640]_ , \new_[5641]_ , \new_[5642]_ ,
    \new_[5643]_ , \new_[5644]_ , \new_[5646]_ , \new_[5647]_ ,
    \new_[5648]_ , \new_[5671]_ , \new_[5672]_ , \new_[5673]_ ,
    \new_[5674]_ , \new_[5675]_ , \new_[5676]_ , \new_[5677]_ ,
    \new_[5678]_ , \new_[5679]_ , \new_[5680]_ , \new_[5681]_ ,
    \new_[5682]_ , \new_[5683]_ , \new_[5684]_ , \new_[5685]_ ,
    \new_[5686]_ , \new_[5687]_ , \new_[5688]_ , \new_[5689]_ ,
    \new_[5690]_ , \new_[5691]_ , \new_[5692]_ , \new_[5693]_ ,
    \new_[5694]_ , \new_[5695]_ , \new_[5696]_ , \new_[5697]_ ,
    \new_[5698]_ , \new_[5699]_ , \new_[5700]_ , \new_[5701]_ ,
    \new_[5702]_ , \new_[5703]_ , \new_[5704]_ , \new_[5705]_ ,
    \new_[5706]_ , \new_[5707]_ , \new_[5708]_ , \new_[5709]_ ,
    \new_[5710]_ , \new_[5711]_ , \new_[5712]_ , \new_[5713]_ ,
    \new_[5714]_ , \new_[5715]_ , \new_[5716]_ , \new_[5717]_ ,
    \new_[5718]_ , \new_[5719]_ , \new_[5720]_ , \new_[5721]_ ,
    \new_[5722]_ , \new_[5723]_ , \new_[5724]_ , \new_[5725]_ ,
    \new_[5726]_ , \new_[5727]_ , \new_[5728]_ , \new_[5729]_ ,
    \new_[5730]_ , \new_[5731]_ , \new_[5732]_ , \new_[5733]_ ,
    \new_[5734]_ , \new_[5735]_ , \new_[5736]_ , \new_[5737]_ ,
    \new_[5738]_ , \new_[5739]_ , \new_[5748]_ , \new_[5749]_ ,
    \new_[5750]_ , \new_[5751]_ , \new_[5752]_ , \new_[5753]_ ,
    \new_[5754]_ , \new_[5755]_ , \new_[5756]_ , \new_[5757]_ ,
    \new_[5758]_ , \new_[5759]_ , \new_[5760]_ , \new_[5761]_ ,
    \new_[5762]_ , \new_[5763]_ , \new_[5764]_ , \new_[5765]_ ,
    \new_[5766]_ , \new_[5767]_ , \new_[5768]_ , \new_[5769]_ ,
    \new_[5770]_ , \new_[5771]_ , \new_[5772]_ , \new_[5773]_ ,
    \new_[5774]_ , \new_[5775]_ , \new_[5776]_ , \new_[5777]_ ,
    \new_[5778]_ , \new_[5779]_ , \new_[5780]_ , \new_[5781]_ ,
    \new_[5782]_ , \new_[5783]_ , \new_[5784]_ , \new_[5785]_ ,
    \new_[5786]_ , \new_[5787]_ , \new_[5788]_ , \new_[5789]_ ,
    \new_[5790]_ , \new_[5792]_ , \new_[5793]_ , \new_[5794]_ ,
    \new_[5796]_ , \new_[5797]_ , \new_[5798]_ , \new_[5799]_ ,
    \new_[5801]_ , \new_[5802]_ , \new_[5803]_ , \new_[5804]_ ,
    \new_[5805]_ , \new_[5806]_ , \new_[5807]_ , \new_[5808]_ ,
    \new_[5809]_ , \new_[5810]_ , \new_[5811]_ , \new_[5812]_ ,
    \new_[5813]_ , \new_[5814]_ , \new_[5815]_ , \new_[5816]_ ,
    \new_[5817]_ , \new_[5818]_ , \new_[5819]_ , \new_[5820]_ ,
    \new_[5821]_ , \new_[5822]_ , \new_[5823]_ , \new_[5824]_ ,
    \new_[5825]_ , \new_[5826]_ , \new_[5827]_ , \new_[5828]_ ,
    \new_[5829]_ , \new_[5830]_ , \new_[5831]_ , \new_[5832]_ ,
    \new_[5833]_ , \new_[5834]_ , \new_[5835]_ , \new_[5836]_ ,
    \new_[5837]_ , \new_[5838]_ , \new_[5839]_ , \new_[5840]_ ,
    \new_[5841]_ , \new_[5842]_ , \new_[5843]_ , \new_[5844]_ ,
    \new_[5845]_ , \new_[5846]_ , \new_[5847]_ , \new_[5848]_ ,
    \new_[5849]_ , \new_[5850]_ , \new_[5851]_ , \new_[5852]_ ,
    \new_[5853]_ , \new_[5854]_ , \new_[5855]_ , \new_[5856]_ ,
    \new_[5857]_ , \new_[5858]_ , \new_[5859]_ , \new_[5860]_ ,
    \new_[5861]_ , \new_[5862]_ , \new_[5863]_ , \new_[5864]_ ,
    \new_[5865]_ , \new_[5866]_ , \new_[5867]_ , \new_[5868]_ ,
    \new_[5869]_ , \new_[5870]_ , \new_[5871]_ , \new_[5872]_ ,
    \new_[5873]_ , \new_[5874]_ , \new_[5875]_ , \new_[5876]_ ,
    \new_[5877]_ , \new_[5878]_ , \new_[5879]_ , \new_[5880]_ ,
    \new_[5881]_ , \new_[5882]_ , \new_[5883]_ , \new_[5884]_ ,
    \new_[5885]_ , \new_[5886]_ , \new_[5887]_ , \new_[5888]_ ,
    \new_[5889]_ , \new_[5890]_ , \new_[5891]_ , \new_[5892]_ ,
    \new_[5893]_ , \new_[5894]_ , \new_[5895]_ , \new_[5896]_ ,
    \new_[5897]_ , \new_[5898]_ , \new_[5899]_ , \new_[5900]_ ,
    \new_[5901]_ , \new_[5902]_ , \new_[5903]_ , \new_[5904]_ ,
    \new_[5905]_ , \new_[5906]_ , \new_[5907]_ , \new_[5908]_ ,
    \new_[5909]_ , \new_[5910]_ , \new_[5911]_ , \new_[5912]_ ,
    \new_[5913]_ , \new_[5914]_ , \new_[5915]_ , \new_[5916]_ ,
    \new_[5917]_ , \new_[5918]_ , \new_[5950]_ , \new_[5951]_ ,
    \new_[5952]_ , \new_[5953]_ , \new_[5954]_ , \new_[5955]_ ,
    \new_[5956]_ , \new_[5957]_ , \new_[5958]_ , \new_[5959]_ ,
    \new_[5960]_ , \new_[5961]_ , \new_[5962]_ , \new_[5963]_ ,
    \new_[5964]_ , \new_[5965]_ , \new_[5966]_ , \new_[5967]_ ,
    \new_[5968]_ , \new_[5969]_ , \new_[5970]_ , \new_[5971]_ ,
    \new_[5972]_ , \new_[5973]_ , \new_[5974]_ , \new_[5975]_ ,
    \new_[5976]_ , \new_[5977]_ , \new_[5978]_ , \new_[5979]_ ,
    \new_[5980]_ , \new_[5981]_ , \new_[5982]_ , \new_[5983]_ ,
    \new_[5984]_ , \new_[5985]_ , \new_[5986]_ , \new_[5988]_ ,
    \new_[5989]_ , \new_[5993]_ , \new_[5997]_ , \new_[5998]_ ,
    \new_[5999]_ , \new_[6000]_ , \new_[6001]_ , \new_[6002]_ ,
    \new_[6003]_ , \new_[6004]_ , \new_[6005]_ , \new_[6006]_ ,
    \new_[6007]_ , \new_[6008]_ , \new_[6009]_ , \new_[6010]_ ,
    \new_[6011]_ , \new_[6012]_ , \new_[6013]_ , \new_[6014]_ ,
    \new_[6015]_ , \new_[6016]_ , \new_[6017]_ , \new_[6018]_ ,
    \new_[6019]_ , \new_[6020]_ , \new_[6021]_ , \new_[6022]_ ,
    \new_[6023]_ , \new_[6024]_ , \new_[6025]_ , \new_[6026]_ ,
    \new_[6027]_ , \new_[6028]_ , \new_[6029]_ , \new_[6030]_ ,
    \new_[6031]_ , \new_[6032]_ , \new_[6033]_ , \new_[6034]_ ,
    \new_[6035]_ , \new_[6036]_ , \new_[6037]_ , \new_[6038]_ ,
    \new_[6039]_ , \new_[6040]_ , \new_[6041]_ , \new_[6042]_ ,
    \new_[6043]_ , \new_[6044]_ , \new_[6045]_ , \new_[6046]_ ,
    \new_[6047]_ , \new_[6048]_ , \new_[6049]_ , \new_[6050]_ ,
    \new_[6051]_ , \new_[6052]_ , \new_[6053]_ , \new_[6054]_ ,
    \new_[6055]_ , \new_[6056]_ , \new_[6057]_ , \new_[6058]_ ,
    \new_[6059]_ , \new_[6060]_ , \new_[6061]_ , \new_[6062]_ ,
    \new_[6063]_ , \new_[6064]_ , \new_[6065]_ , \new_[6066]_ ,
    \new_[6067]_ , \new_[6068]_ , \new_[6069]_ , \new_[6070]_ ,
    \new_[6071]_ , \new_[6072]_ , \new_[6073]_ , \new_[6074]_ ,
    \new_[6075]_ , \new_[6076]_ , \new_[6077]_ , \new_[6078]_ ,
    \new_[6079]_ , \new_[6080]_ , \new_[6081]_ , \new_[6082]_ ,
    \new_[6083]_ , \new_[6084]_ , \new_[6085]_ , \new_[6086]_ ,
    \new_[6087]_ , \new_[6088]_ , \new_[6089]_ , \new_[6090]_ ,
    \new_[6091]_ , \new_[6092]_ , \new_[6093]_ , \new_[6094]_ ,
    \new_[6095]_ , \new_[6096]_ , \new_[6097]_ , \new_[6098]_ ,
    \new_[6099]_ , \new_[6100]_ , \new_[6101]_ , \new_[6102]_ ,
    \new_[6103]_ , \new_[6104]_ , \new_[6105]_ , \new_[6106]_ ,
    \new_[6107]_ , \new_[6108]_ , \new_[6109]_ , \new_[6110]_ ,
    \new_[6111]_ , \new_[6112]_ , \new_[6113]_ , \new_[6114]_ ,
    \new_[6115]_ , \new_[6116]_ , \new_[6117]_ , \new_[6118]_ ,
    \new_[6119]_ , \new_[6120]_ , \new_[6121]_ , \new_[6122]_ ,
    \new_[6123]_ , \new_[6124]_ , \new_[6125]_ , \new_[6126]_ ,
    \new_[6127]_ , \new_[6128]_ , \new_[6129]_ , \new_[6130]_ ,
    \new_[6131]_ , \new_[6132]_ , \new_[6133]_ , \new_[6134]_ ,
    \new_[6135]_ , \new_[6136]_ , \new_[6137]_ , \new_[6138]_ ,
    \new_[6139]_ , \new_[6140]_ , \new_[6141]_ , \new_[6142]_ ,
    \new_[6143]_ , \new_[6144]_ , \new_[6145]_ , \new_[6146]_ ,
    \new_[6147]_ , \new_[6148]_ , \new_[6149]_ , \new_[6150]_ ,
    \new_[6151]_ , \new_[6152]_ , \new_[6153]_ , \new_[6154]_ ,
    \new_[6155]_ , \new_[6156]_ , \new_[6157]_ , \new_[6158]_ ,
    \new_[6159]_ , \new_[6160]_ , \new_[6161]_ , \new_[6162]_ ,
    \new_[6163]_ , \new_[6164]_ , \new_[6165]_ , \new_[6166]_ ,
    \new_[6167]_ , \new_[6168]_ , \new_[6169]_ , \new_[6170]_ ,
    \new_[6171]_ , \new_[6172]_ , \new_[6173]_ , \new_[6174]_ ,
    \new_[6175]_ , \new_[6176]_ , \new_[6177]_ , \new_[6178]_ ,
    \new_[6179]_ , \new_[6180]_ , \new_[6181]_ , \new_[6182]_ ,
    \new_[6183]_ , \new_[6184]_ , \new_[6185]_ , \new_[6186]_ ,
    \new_[6187]_ , \new_[6188]_ , \new_[6189]_ , \new_[6190]_ ,
    \new_[6191]_ , \new_[6192]_ , \new_[6193]_ , \new_[6194]_ ,
    \new_[6195]_ , \new_[6196]_ , \new_[6197]_ , \new_[6228]_ ,
    \new_[6229]_ , \new_[6230]_ , \new_[6231]_ , \new_[6232]_ ,
    \new_[6233]_ , \new_[6234]_ , \new_[6235]_ , \new_[6236]_ ,
    \new_[6237]_ , \new_[6238]_ , \new_[6239]_ , \new_[6240]_ ,
    \new_[6241]_ , \new_[6242]_ , \new_[6243]_ , \new_[6244]_ ,
    \new_[6245]_ , \new_[6246]_ , \new_[6247]_ , \new_[6248]_ ,
    \new_[6249]_ , \new_[6250]_ , \new_[6251]_ , \new_[6252]_ ,
    \new_[6253]_ , \new_[6254]_ , \new_[6255]_ , \new_[6256]_ ,
    \new_[6257]_ , \new_[6258]_ , \new_[6259]_ , \new_[6260]_ ,
    \new_[6261]_ , \new_[6262]_ , \new_[6263]_ , \new_[6264]_ ,
    \new_[6265]_ , \new_[6266]_ , \new_[6267]_ , \new_[6268]_ ,
    \new_[6269]_ , \new_[6270]_ , \new_[6271]_ , \new_[6272]_ ,
    \new_[6273]_ , \new_[6274]_ , \new_[6275]_ , \new_[6276]_ ,
    \new_[6277]_ , \new_[6278]_ , \new_[6279]_ , \new_[6280]_ ,
    \new_[6281]_ , \new_[6282]_ , \new_[6283]_ , \new_[6284]_ ,
    \new_[6285]_ , \new_[6286]_ , \new_[6287]_ , \new_[6288]_ ,
    \new_[6289]_ , \new_[6290]_ , \new_[6291]_ , \new_[6292]_ ,
    \new_[6293]_ , \new_[6294]_ , \new_[6295]_ , \new_[6296]_ ,
    \new_[6297]_ , \new_[6298]_ , \new_[6299]_ , \new_[6300]_ ,
    \new_[6301]_ , \new_[6302]_ , \new_[6303]_ , \new_[6304]_ ,
    \new_[6305]_ , \new_[6306]_ , \new_[6307]_ , \new_[6308]_ ,
    \new_[6309]_ , \new_[6310]_ , \new_[6311]_ , \new_[6312]_ ,
    \new_[6313]_ , \new_[6314]_ , \new_[6315]_ , \new_[6316]_ ,
    \new_[6317]_ , \new_[6318]_ , \new_[6319]_ , \new_[6320]_ ,
    \new_[6321]_ , \new_[6322]_ , \new_[6323]_ , \new_[6324]_ ,
    \new_[6325]_ , \new_[6326]_ , \new_[6327]_ , \new_[6328]_ ,
    \new_[6329]_ , \new_[6330]_ , \new_[6331]_ , \new_[6332]_ ,
    \new_[6333]_ , \new_[6334]_ , \new_[6335]_ , \new_[6336]_ ,
    \new_[6337]_ , \new_[6338]_ , \new_[6339]_ , \new_[6340]_ ,
    \new_[6341]_ , \new_[6342]_ , \new_[6343]_ , \new_[6344]_ ,
    \new_[6345]_ , \new_[6346]_ , \new_[6347]_ , \new_[6348]_ ,
    \new_[6349]_ , \new_[6350]_ , \new_[6351]_ , \new_[6352]_ ,
    \new_[6353]_ , \new_[6354]_ , \new_[6355]_ , \new_[6356]_ ,
    \new_[6357]_ , \new_[6358]_ , \new_[6359]_ , \new_[6360]_ ,
    \new_[6361]_ , \new_[6362]_ , \new_[6363]_ , \new_[6364]_ ,
    \new_[6365]_ , \new_[6366]_ , \new_[6367]_ , \new_[6368]_ ,
    \new_[6369]_ , \new_[6370]_ , \new_[6371]_ , \new_[6372]_ ,
    \new_[6373]_ , \new_[6374]_ , \new_[6375]_ , \new_[6376]_ ,
    \new_[6377]_ , \new_[6378]_ , \new_[6379]_ , \new_[6380]_ ,
    \new_[6381]_ , \new_[6382]_ , \new_[6383]_ , \new_[6384]_ ,
    \new_[6385]_ , \new_[6386]_ , \new_[6387]_ , \new_[6388]_ ,
    \new_[6389]_ , \new_[6390]_ , \new_[6391]_ , \new_[6392]_ ,
    \new_[6393]_ , \new_[6394]_ , \new_[6395]_ , \new_[6396]_ ,
    \new_[6397]_ , \new_[6398]_ , \new_[6399]_ , \new_[6400]_ ,
    \new_[6401]_ , \new_[6402]_ , \new_[6403]_ , \new_[6404]_ ,
    \new_[6405]_ , \new_[6406]_ , \new_[6407]_ , \new_[6408]_ ,
    \new_[6409]_ , \new_[6410]_ , \new_[6411]_ , \new_[6412]_ ,
    \new_[6413]_ , \new_[6414]_ , \new_[6415]_ , \new_[6416]_ ,
    \new_[6417]_ , \new_[6418]_ , \new_[6419]_ , \new_[6420]_ ,
    \new_[6421]_ , \new_[6422]_ , \new_[6423]_ , \new_[6424]_ ,
    \new_[6425]_ , \new_[6426]_ , \new_[6427]_ , \new_[6428]_ ,
    \new_[6429]_ , \new_[6430]_ , \new_[6431]_ , \new_[6432]_ ,
    \new_[6433]_ , \new_[6434]_ , \new_[6435]_ , \new_[6436]_ ,
    \new_[6437]_ , \new_[6438]_ , \new_[6439]_ , \new_[6440]_ ,
    \new_[6441]_ , \new_[6442]_ , \new_[6443]_ , \new_[6444]_ ,
    \new_[6445]_ , \new_[6446]_ , \new_[6447]_ , \new_[6448]_ ,
    \new_[6449]_ , \new_[6450]_ , \new_[6451]_ , \new_[6452]_ ,
    \new_[6453]_ , \new_[6454]_ , \new_[6455]_ , \new_[6456]_ ,
    \new_[6457]_ , \new_[6458]_ , \new_[6459]_ , \new_[6460]_ ,
    \new_[6461]_ , \new_[6462]_ , \new_[6463]_ , \new_[6464]_ ,
    \new_[6465]_ , \new_[6466]_ , \new_[6467]_ , \new_[6468]_ ,
    \new_[6469]_ , \new_[6470]_ , \new_[6471]_ , \new_[6472]_ ,
    \new_[6473]_ , \new_[6474]_ , \new_[6475]_ , \new_[6476]_ ,
    \new_[6477]_ , \new_[6478]_ , \new_[6479]_ , \new_[6480]_ ,
    \new_[6481]_ , \new_[6482]_ , \new_[6483]_ , \new_[6484]_ ,
    \new_[6485]_ , \new_[6486]_ , \new_[6487]_ , \new_[6488]_ ,
    \new_[6489]_ , \new_[6490]_ , \new_[6491]_ , \new_[6492]_ ,
    \new_[6493]_ , \new_[6494]_ , \new_[6495]_ , \new_[6496]_ ,
    \new_[6497]_ , \new_[6498]_ , \new_[6499]_ , \new_[6500]_ ,
    \new_[6501]_ , \new_[6502]_ , \new_[6503]_ , \new_[6504]_ ,
    \new_[6505]_ , \new_[6506]_ , \new_[6507]_ , \new_[6508]_ ,
    \new_[6509]_ , \new_[6510]_ , \new_[6511]_ , \new_[6512]_ ,
    \new_[6513]_ , \new_[6514]_ , \new_[6515]_ , \new_[6516]_ ,
    \new_[6517]_ , \new_[6518]_ , \new_[6519]_ , \new_[6520]_ ,
    \new_[6521]_ , \new_[6522]_ , \new_[6523]_ , \new_[6524]_ ,
    \new_[6525]_ , \new_[6526]_ , \new_[6527]_ , \new_[6528]_ ,
    \new_[6529]_ , \new_[6530]_ , \new_[6531]_ , \new_[6532]_ ,
    \new_[6533]_ , \new_[6534]_ , \new_[6535]_ , \new_[6536]_ ,
    \new_[6537]_ , \new_[6538]_ , \new_[6539]_ , \new_[6540]_ ,
    \new_[6541]_ , \new_[6542]_ , \new_[6543]_ , \new_[6544]_ ,
    \new_[6545]_ , \new_[6546]_ , \new_[6547]_ , \new_[6548]_ ,
    \new_[6549]_ , \new_[6550]_ , \new_[6551]_ , \new_[6552]_ ,
    \new_[6553]_ , \new_[6554]_ , \new_[6555]_ , \new_[6556]_ ,
    \new_[6557]_ , \new_[6558]_ , \new_[6583]_ , \new_[6584]_ ,
    \new_[6585]_ , \new_[6586]_ , \new_[6587]_ , \new_[6588]_ ,
    \new_[6589]_ , \new_[6590]_ , \new_[6591]_ , \new_[6592]_ ,
    \new_[6593]_ , \new_[6594]_ , \new_[6595]_ , \new_[6596]_ ,
    \new_[6597]_ , \new_[6598]_ , \new_[6599]_ , \new_[6600]_ ,
    \new_[6601]_ , \new_[6602]_ , \new_[6603]_ , \new_[6604]_ ,
    \new_[6605]_ , \new_[6606]_ , \new_[6607]_ , \new_[6608]_ ,
    \new_[6609]_ , \new_[6610]_ , \new_[6611]_ , \new_[6612]_ ,
    \new_[6613]_ , \new_[6614]_ , \new_[6615]_ , \new_[6616]_ ,
    \new_[6617]_ , \new_[6618]_ , \new_[6619]_ , \new_[6620]_ ,
    \new_[6621]_ , \new_[6622]_ , \new_[6623]_ , \new_[6624]_ ,
    \new_[6625]_ , \new_[6626]_ , \new_[6627]_ , \new_[6628]_ ,
    \new_[6629]_ , \new_[6630]_ , \new_[6631]_ , \new_[6632]_ ,
    \new_[6633]_ , \new_[6634]_ , \new_[6635]_ , \new_[6636]_ ,
    \new_[6637]_ , \new_[6638]_ , \new_[6639]_ , \new_[6640]_ ,
    \new_[6641]_ , \new_[6642]_ , \new_[6643]_ , \new_[6644]_ ,
    \new_[6645]_ , \new_[6646]_ , \new_[6647]_ , \new_[6648]_ ,
    \new_[6649]_ , \new_[6650]_ , \new_[6651]_ , \new_[6652]_ ,
    \new_[6653]_ , \new_[6654]_ , \new_[6655]_ , \new_[6656]_ ,
    \new_[6657]_ , \new_[6658]_ , \new_[6659]_ , \new_[6660]_ ,
    \new_[6661]_ , \new_[6662]_ , \new_[6663]_ , \new_[6664]_ ,
    \new_[6665]_ , \new_[6666]_ , \new_[6667]_ , \new_[6668]_ ,
    \new_[6669]_ , \new_[6670]_ , \new_[6671]_ , \new_[6672]_ ,
    \new_[6673]_ , \new_[6674]_ , \new_[6675]_ , \new_[6676]_ ,
    \new_[6677]_ , \new_[6678]_ , \new_[6679]_ , \new_[6680]_ ,
    \new_[6681]_ , \new_[6682]_ , \new_[6683]_ , \new_[6684]_ ,
    \new_[6685]_ , \new_[6686]_ , \new_[6687]_ , \new_[6688]_ ,
    \new_[6689]_ , \new_[6690]_ , \new_[6691]_ , \new_[6692]_ ,
    \new_[6693]_ , \new_[6694]_ , \new_[6695]_ , \new_[6696]_ ,
    \new_[6697]_ , \new_[6698]_ , \new_[6699]_ , \new_[6700]_ ,
    \new_[6701]_ , \new_[6702]_ , \new_[6703]_ , \new_[6704]_ ,
    \new_[6705]_ , \new_[6706]_ , \new_[6707]_ , \new_[6708]_ ,
    \new_[6709]_ , \new_[6710]_ , \new_[6711]_ , \new_[6712]_ ,
    \new_[6713]_ , \new_[6714]_ , \new_[6715]_ , \new_[6716]_ ,
    \new_[6717]_ , \new_[6718]_ , \new_[6719]_ , \new_[6720]_ ,
    \new_[6721]_ , \new_[6722]_ , \new_[6723]_ , \new_[6724]_ ,
    \new_[6725]_ , \new_[6726]_ , \new_[6727]_ , \new_[6728]_ ,
    \new_[6729]_ , \new_[6730]_ , \new_[6731]_ , \new_[6732]_ ,
    \new_[6733]_ , \new_[6734]_ , \new_[6735]_ , \new_[6736]_ ,
    \new_[6737]_ , \new_[6738]_ , \new_[6739]_ , \new_[6740]_ ,
    \new_[6741]_ , \new_[6742]_ , \new_[6743]_ , \new_[6744]_ ,
    \new_[6745]_ , \new_[6746]_ , \new_[6747]_ , \new_[6748]_ ,
    \new_[6749]_ , \new_[6750]_ , \new_[6751]_ , \new_[6752]_ ,
    \new_[6753]_ , \new_[6754]_ , \new_[6755]_ , \new_[6756]_ ,
    \new_[6757]_ , \new_[6758]_ , \new_[6759]_ , \new_[6760]_ ,
    \new_[6761]_ , \new_[6762]_ , \new_[6763]_ , \new_[6764]_ ,
    \new_[6765]_ , \new_[6766]_ , \new_[6767]_ , \new_[6768]_ ,
    \new_[6769]_ , \new_[6770]_ , \new_[6771]_ , \new_[6772]_ ,
    \new_[6773]_ , \new_[6774]_ , \new_[6775]_ , \new_[6776]_ ,
    \new_[6777]_ , \new_[6778]_ , \new_[6779]_ , \new_[6780]_ ,
    \new_[6781]_ , \new_[6782]_ , \new_[6783]_ , \new_[6784]_ ,
    \new_[6785]_ , \new_[6786]_ , \new_[6787]_ , \new_[6788]_ ,
    \new_[6789]_ , \new_[6790]_ , \new_[6791]_ , \new_[6792]_ ,
    \new_[6793]_ , \new_[6794]_ , \new_[6795]_ , \new_[6796]_ ,
    \new_[6797]_ , \new_[6798]_ , \new_[6799]_ , \new_[6800]_ ,
    \new_[6801]_ , \new_[6802]_ , \new_[6803]_ , \new_[6804]_ ,
    \new_[6805]_ , \new_[6806]_ , \new_[6807]_ , \new_[6808]_ ,
    \new_[6809]_ , \new_[6810]_ , \new_[6811]_ , \new_[6812]_ ,
    \new_[6813]_ , \new_[6814]_ , \new_[6815]_ , \new_[6816]_ ,
    \new_[6817]_ , \new_[6818]_ , \new_[6819]_ , \new_[6820]_ ,
    \new_[6821]_ , \new_[6822]_ , \new_[6823]_ , \new_[6824]_ ,
    \new_[6825]_ , \new_[6826]_ , \new_[6827]_ , \new_[6828]_ ,
    \new_[6829]_ , \new_[6830]_ , \new_[6831]_ , \new_[6832]_ ,
    \new_[6833]_ , \new_[6834]_ , \new_[6835]_ , \new_[6836]_ ,
    \new_[6837]_ , \new_[6838]_ , \new_[6839]_ , \new_[6840]_ ,
    \new_[6841]_ , \new_[6842]_ , \new_[6843]_ , \new_[6844]_ ,
    \new_[6845]_ , \new_[6846]_ , \new_[6847]_ , \new_[6848]_ ,
    \new_[6849]_ , \new_[6850]_ , \new_[6851]_ , \new_[6852]_ ,
    \new_[6853]_ , \new_[6854]_ , \new_[6855]_ , \new_[6856]_ ,
    \new_[6857]_ , \new_[6858]_ , \new_[6859]_ , \new_[6860]_ ,
    \new_[6861]_ , \new_[6862]_ , \new_[6863]_ , \new_[6864]_ ,
    \new_[6865]_ , \new_[6866]_ , \new_[6867]_ , \new_[6868]_ ,
    \new_[6869]_ , \new_[6870]_ , \new_[6871]_ , \new_[6872]_ ,
    \new_[6873]_ , \new_[6874]_ , \new_[6875]_ , \new_[6876]_ ,
    \new_[6877]_ , \new_[6878]_ , \new_[6879]_ , \new_[6880]_ ,
    \new_[6881]_ , \new_[6882]_ , \new_[6883]_ , \new_[6884]_ ,
    \new_[6885]_ , \new_[6886]_ , \new_[6887]_ , \new_[6888]_ ,
    \new_[6889]_ , \new_[6890]_ , \new_[6891]_ , \new_[6892]_ ,
    \new_[6893]_ , \new_[6894]_ , \new_[6895]_ , \new_[6896]_ ,
    \new_[6897]_ , \new_[6898]_ , \new_[6899]_ , \new_[6900]_ ,
    \new_[6901]_ , \new_[6902]_ , \new_[6903]_ , \new_[6904]_ ,
    \new_[6905]_ , \new_[6906]_ , \new_[6907]_ , \new_[6908]_ ,
    \new_[6909]_ , \new_[6910]_ , \new_[6911]_ , \new_[6912]_ ,
    \new_[6913]_ , \new_[6914]_ , \new_[6915]_ , \new_[6916]_ ,
    \new_[6917]_ , \new_[6918]_ , \new_[6919]_ , \new_[6920]_ ,
    \new_[6921]_ , \new_[6922]_ , \new_[6923]_ , \new_[6924]_ ,
    \new_[6925]_ , \new_[6926]_ , \new_[6927]_ , \new_[6928]_ ,
    \new_[6929]_ , \new_[6930]_ , \new_[6931]_ , \new_[6932]_ ,
    \new_[6933]_ , \new_[6934]_ , \new_[6935]_ , \new_[6936]_ ,
    \new_[6939]_ , \new_[6940]_ , \new_[6941]_ , \new_[6942]_ ,
    \new_[6943]_ , \new_[6944]_ , \new_[6945]_ , \new_[6946]_ ,
    \new_[6947]_ , \new_[6948]_ , \new_[6949]_ , \new_[6950]_ ,
    \new_[6951]_ , \new_[6952]_ , \new_[6953]_ , \new_[6954]_ ,
    \new_[6955]_ , \new_[6956]_ , \new_[6957]_ , \new_[6958]_ ,
    \new_[6959]_ , \new_[6960]_ , \new_[6961]_ , \new_[6962]_ ,
    \new_[6963]_ , \new_[6964]_ , \new_[6965]_ , \new_[6966]_ ,
    \new_[6967]_ , \new_[6968]_ , \new_[6969]_ , \new_[6970]_ ,
    \new_[6971]_ , \new_[6972]_ , \new_[6973]_ , \new_[6974]_ ,
    \new_[6975]_ , \new_[6976]_ , \new_[6977]_ , \new_[6978]_ ,
    \new_[6979]_ , \new_[6980]_ , \new_[6981]_ , \new_[6982]_ ,
    \new_[6983]_ , \new_[6984]_ , \new_[6985]_ , \new_[6987]_ ,
    \new_[6989]_ , \new_[6990]_ , \new_[6991]_ , \new_[6992]_ ,
    \new_[6993]_ , \new_[6994]_ , \new_[6996]_ , \new_[6997]_ ,
    \new_[6998]_ , \new_[6999]_ , \new_[7001]_ , \new_[7003]_ ,
    \new_[7004]_ , \new_[7005]_ , \new_[7006]_ , \new_[7008]_ ,
    \new_[7009]_ , \new_[7010]_ , \new_[7011]_ , \new_[7012]_ ,
    \new_[7015]_ , \new_[7016]_ , \new_[7017]_ , \new_[7018]_ ,
    \new_[7019]_ , \new_[7020]_ , \new_[7021]_ , \new_[7022]_ ,
    \new_[7023]_ , \new_[7024]_ , \new_[7025]_ , \new_[7026]_ ,
    \new_[7027]_ , \new_[7028]_ , \new_[7029]_ , \new_[7030]_ ,
    \new_[7031]_ , \new_[7032]_ , \new_[7033]_ , \new_[7034]_ ,
    \new_[7035]_ , \new_[7036]_ , \new_[7037]_ , \new_[7038]_ ,
    \new_[7039]_ , \new_[7040]_ , \new_[7041]_ , \new_[7042]_ ,
    \new_[7043]_ , \new_[7044]_ , \new_[7045]_ , \new_[7046]_ ,
    \new_[7047]_ , \new_[7048]_ , \new_[7049]_ , \new_[7050]_ ,
    \new_[7051]_ , \new_[7052]_ , \new_[7053]_ , \new_[7054]_ ,
    \new_[7055]_ , \new_[7056]_ , \new_[7057]_ , \new_[7058]_ ,
    \new_[7059]_ , \new_[7060]_ , \new_[7061]_ , \new_[7062]_ ,
    \new_[7063]_ , \new_[7064]_ , \new_[7065]_ , \new_[7066]_ ,
    \new_[7067]_ , \new_[7068]_ , \new_[7069]_ , \new_[7070]_ ,
    \new_[7071]_ , \new_[7072]_ , \new_[7073]_ , \new_[7074]_ ,
    \new_[7075]_ , \new_[7076]_ , \new_[7077]_ , \new_[7078]_ ,
    \new_[7079]_ , \new_[7080]_ , \new_[7081]_ , \new_[7082]_ ,
    \new_[7083]_ , \new_[7084]_ , \new_[7085]_ , \new_[7086]_ ,
    \new_[7087]_ , \new_[7088]_ , \new_[7089]_ , \new_[7090]_ ,
    \new_[7091]_ , \new_[7092]_ , \new_[7093]_ , \new_[7094]_ ,
    \new_[7095]_ , \new_[7096]_ , \new_[7097]_ , \new_[7098]_ ,
    \new_[7099]_ , \new_[7100]_ , \new_[7101]_ , \new_[7102]_ ,
    \new_[7103]_ , \new_[7104]_ , \new_[7105]_ , \new_[7106]_ ,
    \new_[7107]_ , \new_[7108]_ , \new_[7109]_ , \new_[7110]_ ,
    \new_[7111]_ , \new_[7112]_ , \new_[7113]_ , \new_[7114]_ ,
    \new_[7115]_ , \new_[7116]_ , \new_[7117]_ , \new_[7118]_ ,
    \new_[7119]_ , \new_[7120]_ , \new_[7121]_ , \new_[7122]_ ,
    \new_[7123]_ , \new_[7124]_ , \new_[7125]_ , \new_[7126]_ ,
    \new_[7127]_ , \new_[7128]_ , \new_[7129]_ , \new_[7130]_ ,
    \new_[7131]_ , \new_[7132]_ , \new_[7133]_ , \new_[7134]_ ,
    \new_[7135]_ , \new_[7136]_ , \new_[7137]_ , \new_[7138]_ ,
    \new_[7139]_ , \new_[7140]_ , \new_[7141]_ , \new_[7142]_ ,
    \new_[7143]_ , \new_[7144]_ , \new_[7145]_ , \new_[7146]_ ,
    \new_[7147]_ , \new_[7148]_ , \new_[7149]_ , \new_[7150]_ ,
    \new_[7151]_ , \new_[7152]_ , \new_[7153]_ , \new_[7154]_ ,
    \new_[7155]_ , \new_[7156]_ , \new_[7157]_ , \new_[7158]_ ,
    \new_[7159]_ , \new_[7160]_ , \new_[7161]_ , \new_[7162]_ ,
    \new_[7163]_ , \new_[7164]_ , \new_[7165]_ , \new_[7166]_ ,
    \new_[7167]_ , \new_[7168]_ , \new_[7169]_ , \new_[7170]_ ,
    \new_[7171]_ , \new_[7172]_ , \new_[7173]_ , \new_[7174]_ ,
    \new_[7175]_ , \new_[7176]_ , \new_[7177]_ , \new_[7178]_ ,
    \new_[7179]_ , \new_[7180]_ , \new_[7181]_ , \new_[7182]_ ,
    \new_[7183]_ , \new_[7184]_ , \new_[7185]_ , \new_[7186]_ ,
    \new_[7187]_ , \new_[7188]_ , \new_[7189]_ , \new_[7190]_ ,
    \new_[7191]_ , \new_[7192]_ , \new_[7193]_ , \new_[7194]_ ,
    \new_[7195]_ , \new_[7196]_ , \new_[7197]_ , \new_[7198]_ ,
    \new_[7199]_ , \new_[7200]_ , \new_[7201]_ , \new_[7202]_ ,
    \new_[7203]_ , \new_[7204]_ , \new_[7205]_ , \new_[7206]_ ,
    \new_[7207]_ , \new_[7208]_ , \new_[7209]_ , \new_[7210]_ ,
    \new_[7211]_ , \new_[7212]_ , \new_[7213]_ , \new_[7214]_ ,
    \new_[7215]_ , \new_[7216]_ , \new_[7217]_ , \new_[7218]_ ,
    \new_[7219]_ , \new_[7220]_ , \new_[7221]_ , \new_[7222]_ ,
    \new_[7223]_ , \new_[7224]_ , \new_[7225]_ , \new_[7226]_ ,
    \new_[7227]_ , \new_[7228]_ , \new_[7229]_ , \new_[7230]_ ,
    \new_[7231]_ , \new_[7232]_ , \new_[7233]_ , \new_[7234]_ ,
    \new_[7235]_ , \new_[7236]_ , \new_[7237]_ , \new_[7238]_ ,
    \new_[7239]_ , \new_[7240]_ , \new_[7241]_ , \new_[7242]_ ,
    \new_[7243]_ , \new_[7244]_ , \new_[7245]_ , \new_[7246]_ ,
    \new_[7247]_ , \new_[7248]_ , \new_[7249]_ , \new_[7250]_ ,
    \new_[7251]_ , \new_[7252]_ , \new_[7253]_ , \new_[7254]_ ,
    \new_[7255]_ , \new_[7256]_ , \new_[7257]_ , \new_[7258]_ ,
    \new_[7259]_ , \new_[7260]_ , \new_[7261]_ , \new_[7262]_ ,
    \new_[7263]_ , \new_[7264]_ , \new_[7265]_ , \new_[7266]_ ,
    \new_[7275]_ , \new_[7281]_ , \new_[7283]_ , \new_[7288]_ ,
    \new_[7293]_ , \new_[7302]_ , \new_[7303]_ , \new_[7304]_ ,
    \new_[7306]_ , \new_[7307]_ , \new_[7308]_ , \new_[7309]_ ,
    \new_[7310]_ , \new_[7311]_ , \new_[7312]_ , \new_[7313]_ ,
    \new_[7314]_ , \new_[7315]_ , \new_[7316]_ , \new_[7317]_ ,
    \new_[7318]_ , \new_[7319]_ , \new_[7320]_ , \new_[7321]_ ,
    \new_[7322]_ , \new_[7323]_ , \new_[7324]_ , \new_[7325]_ ,
    \new_[7326]_ , \new_[7327]_ , \new_[7328]_ , \new_[7329]_ ,
    \new_[7330]_ , \new_[7331]_ , \new_[7332]_ , \new_[7333]_ ,
    \new_[7334]_ , \new_[7335]_ , \new_[7336]_ , \new_[7337]_ ,
    \new_[7338]_ , \new_[7339]_ , \new_[7340]_ , \new_[7341]_ ,
    \new_[7342]_ , \new_[7343]_ , \new_[7344]_ , \new_[7345]_ ,
    \new_[7346]_ , \new_[7347]_ , \new_[7348]_ , \new_[7349]_ ,
    \new_[7350]_ , \new_[7351]_ , \new_[7352]_ , \new_[7353]_ ,
    \new_[7354]_ , \new_[7355]_ , \new_[7356]_ , \new_[7357]_ ,
    \new_[7358]_ , \new_[7359]_ , \new_[7360]_ , \new_[7361]_ ,
    \new_[7362]_ , \new_[7363]_ , \new_[7364]_ , \new_[7365]_ ,
    \new_[7366]_ , \new_[7367]_ , \new_[7368]_ , \new_[7369]_ ,
    \new_[7370]_ , \new_[7371]_ , \new_[7372]_ , \new_[7373]_ ,
    \new_[7374]_ , \new_[7375]_ , \new_[7376]_ , \new_[7377]_ ,
    \new_[7378]_ , \new_[7379]_ , \new_[7380]_ , \new_[7381]_ ,
    \new_[7382]_ , \new_[7383]_ , \new_[7384]_ , \new_[7385]_ ,
    \new_[7386]_ , \new_[7387]_ , \new_[7388]_ , \new_[7389]_ ,
    \new_[7390]_ , \new_[7391]_ , \new_[7392]_ , \new_[7393]_ ,
    \new_[7394]_ , \new_[7395]_ , \new_[7396]_ , \new_[7397]_ ,
    \new_[7398]_ , \new_[7399]_ , \new_[7400]_ , \new_[7401]_ ,
    \new_[7402]_ , \new_[7403]_ , \new_[7404]_ , \new_[7405]_ ,
    \new_[7406]_ , \new_[7407]_ , \new_[7408]_ , \new_[7409]_ ,
    \new_[7410]_ , \new_[7411]_ , \new_[7412]_ , \new_[7413]_ ,
    \new_[7414]_ , \new_[7415]_ , \new_[7416]_ , \new_[7417]_ ,
    \new_[7418]_ , \new_[7419]_ , \new_[7420]_ , \new_[7421]_ ,
    \new_[7422]_ , \new_[7423]_ , \new_[7424]_ , \new_[7425]_ ,
    \new_[7426]_ , \new_[7427]_ , \new_[7428]_ , \new_[7429]_ ,
    \new_[7431]_ , \new_[7432]_ , \new_[7433]_ , \new_[7434]_ ,
    \new_[7435]_ , \new_[7436]_ , \new_[7437]_ , \new_[7438]_ ,
    \new_[7439]_ , \new_[7440]_ , \new_[7441]_ , \new_[7442]_ ,
    \new_[7443]_ , \new_[7444]_ , \new_[7445]_ , \new_[7446]_ ,
    \new_[7447]_ , \new_[7448]_ , \new_[7449]_ , \new_[7450]_ ,
    \new_[7451]_ , \new_[7452]_ , \new_[7453]_ , \new_[7454]_ ,
    \new_[7455]_ , \new_[7456]_ , \new_[7457]_ , \new_[7458]_ ,
    \new_[7459]_ , \new_[7460]_ , \new_[7461]_ , \new_[7462]_ ,
    \new_[7463]_ , \new_[7464]_ , \new_[7465]_ , \new_[7466]_ ,
    \new_[7467]_ , \new_[7468]_ , \new_[7469]_ , \new_[7470]_ ,
    \new_[7471]_ , \new_[7472]_ , \new_[7473]_ , \new_[7474]_ ,
    \new_[7475]_ , \new_[7476]_ , \new_[7477]_ , \new_[7478]_ ,
    \new_[7479]_ , \new_[7480]_ , \new_[7481]_ , \new_[7482]_ ,
    \new_[7483]_ , \new_[7484]_ , \new_[7486]_ , \new_[7488]_ ,
    \new_[7489]_ , \new_[7491]_ , \new_[7492]_ , \new_[7494]_ ,
    \new_[7496]_ , \new_[7497]_ , \new_[7498]_ , \new_[7499]_ ,
    \new_[7500]_ , \new_[7501]_ , \new_[7503]_ , \new_[7504]_ ,
    \new_[7505]_ , \new_[7507]_ , \new_[7508]_ , \new_[7509]_ ,
    \new_[7510]_ , \new_[7631]_ , \new_[7641]_ , \new_[7642]_ ,
    \new_[7648]_ , \new_[7658]_ , \new_[7665]_ , \new_[7669]_ ,
    \new_[7674]_ , \new_[7679]_ , \new_[7688]_ , \new_[7704]_ ,
    \new_[7705]_ , \new_[7707]_ , \new_[7730]_ , \new_[7734]_ ,
    \new_[7738]_ , \new_[7741]_ , \new_[7746]_ , \new_[7747]_ ,
    \new_[7751]_ , \new_[7764]_ , \new_[7771]_ , \new_[7777]_ ,
    \new_[7783]_ , \new_[7788]_ , \new_[7802]_ , \new_[7803]_ ,
    \new_[7806]_ , \new_[7819]_ , \new_[7822]_ , \new_[7844]_ ,
    \new_[7861]_ , \new_[7866]_ , \new_[7869]_ , \new_[7895]_ ,
    \new_[7900]_ , \new_[7910]_ , \new_[7921]_ , \new_[7926]_ ,
    \new_[7935]_ , \new_[7944]_ , \new_[7953]_ , \new_[7954]_ ,
    \new_[7960]_ , \new_[7961]_ , \new_[7962]_ , \new_[7963]_ ,
    \new_[7964]_ , \new_[7965]_ , \new_[7966]_ , \new_[7967]_ ,
    \new_[7968]_ , \new_[7969]_ , \new_[7970]_ , \new_[7971]_ ,
    \new_[7972]_ , \new_[7973]_ , \new_[7974]_ , \new_[7975]_ ,
    \new_[7976]_ , \new_[7977]_ , \new_[7978]_ , \new_[7979]_ ,
    \new_[7980]_ , \new_[7981]_ , \new_[7982]_ , \new_[7983]_ ,
    \new_[7984]_ , \new_[7985]_ , \new_[7986]_ , \new_[7987]_ ,
    \new_[7988]_ , \new_[7989]_ , \new_[7990]_ , \new_[7991]_ ,
    \new_[7992]_ , \new_[7993]_ , \new_[7994]_ , \new_[7995]_ ,
    \new_[7996]_ , \new_[7997]_ , \new_[7998]_ , \new_[7999]_ ,
    \new_[8000]_ , \new_[8001]_ , \new_[8002]_ , \new_[8003]_ ,
    \new_[8004]_ , \new_[8005]_ , \new_[8006]_ , \new_[8007]_ ,
    \new_[8008]_ , \new_[8009]_ , \new_[8010]_ , \new_[8011]_ ,
    \new_[8012]_ , \new_[8013]_ , \new_[8014]_ , \new_[8015]_ ,
    \new_[8016]_ , \new_[8017]_ , \new_[8018]_ , \new_[8019]_ ,
    \new_[8020]_ , \new_[8021]_ , \new_[8022]_ , \new_[8023]_ ,
    \new_[8024]_ , \new_[8025]_ , \new_[8026]_ , \new_[8027]_ ,
    \new_[8028]_ , \new_[8029]_ , \new_[8030]_ , \new_[8031]_ ,
    \new_[8032]_ , \new_[8033]_ , \new_[8034]_ , \new_[8035]_ ,
    \new_[8036]_ , \new_[8037]_ , \new_[8038]_ , \new_[8039]_ ,
    \new_[8040]_ , \new_[8041]_ , \new_[8042]_ , \new_[8043]_ ,
    \new_[8044]_ , \new_[8045]_ , \new_[8046]_ , \new_[8047]_ ,
    \new_[8048]_ , \new_[8049]_ , \new_[8050]_ , \new_[8051]_ ,
    \new_[8052]_ , \new_[8053]_ , \new_[8054]_ , \new_[8055]_ ,
    \new_[8056]_ , \new_[8057]_ , \new_[8058]_ , \new_[8059]_ ,
    \new_[8060]_ , \new_[8061]_ , \new_[8062]_ , \new_[8063]_ ,
    \new_[8064]_ , \new_[8065]_ , \new_[8066]_ , \new_[8067]_ ,
    \new_[8068]_ , \new_[8069]_ , \new_[8070]_ , \new_[8071]_ ,
    \new_[8072]_ , \new_[8073]_ , \new_[8074]_ , \new_[8075]_ ,
    \new_[8076]_ , \new_[8077]_ , \new_[8078]_ , \new_[8079]_ ,
    \new_[8080]_ , \new_[8081]_ , \new_[8082]_ , \new_[8083]_ ,
    \new_[8084]_ , \new_[8085]_ , \new_[8086]_ , \new_[8087]_ ,
    \new_[8088]_ , \new_[8089]_ , \new_[8090]_ , \new_[8091]_ ,
    \new_[8092]_ , \new_[8093]_ , \new_[8094]_ , \new_[8095]_ ,
    \new_[8096]_ , \new_[8097]_ , \new_[8098]_ , \new_[8099]_ ,
    \new_[8100]_ , \new_[8101]_ , \new_[8102]_ , \new_[8103]_ ,
    \new_[8104]_ , \new_[8105]_ , \new_[8106]_ , \new_[8107]_ ,
    \new_[8108]_ , \new_[8109]_ , \new_[8110]_ , \new_[8111]_ ,
    \new_[8112]_ , \new_[8113]_ , \new_[8114]_ , \new_[8115]_ ,
    \new_[8116]_ , \new_[8117]_ , \new_[8118]_ , \new_[8119]_ ,
    \new_[8120]_ , \new_[8121]_ , \new_[8122]_ , \new_[8123]_ ,
    \new_[8124]_ , \new_[8125]_ , \new_[8126]_ , \new_[8127]_ ,
    \new_[8128]_ , \new_[8129]_ , \new_[8130]_ , \new_[8131]_ ,
    \new_[8132]_ , \new_[8133]_ , \new_[8134]_ , \new_[8135]_ ,
    \new_[8136]_ , \new_[8137]_ , \new_[8138]_ , \new_[8139]_ ,
    \new_[8140]_ , \new_[8141]_ , \new_[8142]_ , \new_[8143]_ ,
    \new_[8144]_ , \new_[8145]_ , \new_[8146]_ , \new_[8147]_ ,
    \new_[8148]_ , \new_[8149]_ , \new_[8150]_ , \new_[8151]_ ,
    \new_[8152]_ , \new_[8153]_ , \new_[8154]_ , \new_[8155]_ ,
    \new_[8156]_ , \new_[8157]_ , \new_[8158]_ , \new_[8159]_ ,
    \new_[8160]_ , \new_[8161]_ , \new_[8162]_ , \new_[8163]_ ,
    \new_[8164]_ , \new_[8165]_ , \new_[8166]_ , \new_[8167]_ ,
    \new_[8168]_ , \new_[8169]_ , \new_[8170]_ , \new_[8171]_ ,
    \new_[8172]_ , \new_[8173]_ , \new_[8174]_ , \new_[8175]_ ,
    \new_[8176]_ , \new_[8177]_ , \new_[8178]_ , \new_[8179]_ ,
    \new_[8180]_ , \new_[8181]_ , \new_[8182]_ , \new_[8183]_ ,
    \new_[8184]_ , \new_[8185]_ , \new_[8186]_ , \new_[8187]_ ,
    \new_[8188]_ , \new_[8189]_ , \new_[8190]_ , \new_[8191]_ ,
    \new_[8192]_ , \new_[8193]_ , \new_[8194]_ , \new_[8195]_ ,
    \new_[8196]_ , \new_[8197]_ , \new_[8198]_ , \new_[8199]_ ,
    \new_[8200]_ , \new_[8201]_ , \new_[8202]_ , \new_[8203]_ ,
    \new_[8204]_ , \new_[8205]_ , \new_[8206]_ , \new_[8207]_ ,
    \new_[8208]_ , \new_[8209]_ , \new_[8210]_ , \new_[8211]_ ,
    \new_[8212]_ , \new_[8213]_ , \new_[8214]_ , \new_[8215]_ ,
    \new_[8216]_ , \new_[8217]_ , \new_[8218]_ , \new_[8219]_ ,
    \new_[8220]_ , \new_[8221]_ , \new_[8222]_ , \new_[8223]_ ,
    \new_[8224]_ , \new_[8226]_ , \new_[8241]_ , \new_[8242]_ ,
    \new_[8261]_ , \new_[8262]_ , \new_[8263]_ , \new_[8264]_ ,
    \new_[8265]_ , \new_[8266]_ , \new_[8268]_ , \new_[8269]_ ,
    \new_[8270]_ , \new_[8271]_ , \new_[8272]_ , \new_[8273]_ ,
    \new_[8274]_ , \new_[8275]_ , \new_[8276]_ , \new_[8277]_ ,
    \new_[8278]_ , \new_[8279]_ , \new_[8280]_ , \new_[8281]_ ,
    \new_[8282]_ , \new_[8283]_ , \new_[8284]_ , \new_[8285]_ ,
    \new_[8286]_ , \new_[8287]_ , \new_[8288]_ , \new_[8289]_ ,
    \new_[8290]_ , \new_[8291]_ , \new_[8292]_ , \new_[8293]_ ,
    \new_[8294]_ , \new_[8295]_ , \new_[8296]_ , \new_[8297]_ ,
    \new_[8298]_ , \new_[8299]_ , \new_[8300]_ , \new_[8301]_ ,
    \new_[8302]_ , \new_[8303]_ , \new_[8304]_ , \new_[8305]_ ,
    \new_[8306]_ , \new_[8307]_ , \new_[8308]_ , \new_[8309]_ ,
    \new_[8310]_ , \new_[8311]_ , \new_[8312]_ , \new_[8313]_ ,
    \new_[8314]_ , \new_[8315]_ , \new_[8316]_ , \new_[8317]_ ,
    \new_[8318]_ , \new_[8319]_ , \new_[8320]_ , \new_[8321]_ ,
    \new_[8322]_ , \new_[8323]_ , \new_[8324]_ , \new_[8325]_ ,
    \new_[8326]_ , \new_[8327]_ , \new_[8328]_ , \new_[8329]_ ,
    \new_[8330]_ , \new_[8331]_ , \new_[8332]_ , \new_[8333]_ ,
    \new_[8334]_ , \new_[8335]_ , \new_[8336]_ , \new_[8337]_ ,
    \new_[8338]_ , \new_[8339]_ , \new_[8340]_ , \new_[8341]_ ,
    \new_[8342]_ , \new_[8343]_ , \new_[8344]_ , \new_[8345]_ ,
    \new_[8346]_ , \new_[8347]_ , \new_[8348]_ , \new_[8349]_ ,
    \new_[8350]_ , \new_[8351]_ , \new_[8352]_ , \new_[8353]_ ,
    \new_[8354]_ , \new_[8355]_ , \new_[8356]_ , \new_[8357]_ ,
    \new_[8358]_ , \new_[8359]_ , \new_[8360]_ , \new_[8361]_ ,
    \new_[8362]_ , \new_[8363]_ , \new_[8364]_ , \new_[8365]_ ,
    \new_[8366]_ , \new_[8367]_ , \new_[8368]_ , \new_[8369]_ ,
    \new_[8370]_ , \new_[8371]_ , \new_[8372]_ , \new_[8373]_ ,
    \new_[8374]_ , \new_[8375]_ , \new_[8376]_ , \new_[8377]_ ,
    \new_[8378]_ , \new_[8379]_ , \new_[8380]_ , \new_[8381]_ ,
    \new_[8382]_ , \new_[8383]_ , \new_[8384]_ , \new_[8385]_ ,
    \new_[8386]_ , \new_[8387]_ , \new_[8388]_ , \new_[8389]_ ,
    \new_[8390]_ , \new_[8391]_ , \new_[8392]_ , \new_[8394]_ ,
    \new_[8395]_ , \new_[8396]_ , \new_[8397]_ , \new_[8398]_ ,
    \new_[8400]_ , \new_[8401]_ , \new_[8548]_ , \new_[8549]_ ,
    \new_[8550]_ , \new_[8551]_ , \new_[8552]_ , \new_[8553]_ ,
    \new_[8554]_ , \new_[8555]_ , \new_[8556]_ , \new_[8557]_ ,
    \new_[8558]_ , \new_[8559]_ , \new_[8560]_ , \new_[8561]_ ,
    \new_[8562]_ , \new_[8563]_ , \new_[8564]_ , \new_[8565]_ ,
    \new_[8566]_ , \new_[8567]_ , \new_[8568]_ , \new_[8569]_ ,
    \new_[8570]_ , \new_[8571]_ , \new_[8572]_ , \new_[8573]_ ,
    \new_[8574]_ , \new_[8575]_ , \new_[8576]_ , \new_[8577]_ ,
    \new_[8578]_ , \new_[8579]_ , \new_[8580]_ , \new_[8581]_ ,
    \new_[8582]_ , \new_[8583]_ , \new_[8584]_ , \new_[8585]_ ,
    \new_[8586]_ , \new_[8587]_ , \new_[8588]_ , \new_[8589]_ ,
    \new_[8590]_ , \new_[8591]_ , \new_[8592]_ , \new_[8593]_ ,
    \new_[8594]_ , \new_[8595]_ , \new_[8596]_ , \new_[8597]_ ,
    \new_[8598]_ , \new_[8599]_ , \new_[8600]_ , \new_[8601]_ ,
    \new_[8602]_ , \new_[8603]_ , \new_[8604]_ , \new_[8605]_ ,
    \new_[8606]_ , \new_[8607]_ , \new_[8608]_ , \new_[8609]_ ,
    \new_[8610]_ , \new_[8611]_ , \new_[8612]_ , \new_[8613]_ ,
    \new_[8614]_ , \new_[8615]_ , \new_[8616]_ , \new_[8617]_ ,
    \new_[8618]_ , \new_[8619]_ , \new_[8620]_ , \new_[8621]_ ,
    \new_[8622]_ , \new_[8623]_ , \new_[8624]_ , \new_[8625]_ ,
    \new_[8626]_ , \new_[8627]_ , \new_[8628]_ , \new_[8629]_ ,
    \new_[8630]_ , \new_[8631]_ , \new_[8632]_ , \new_[8633]_ ,
    \new_[8634]_ , \new_[8635]_ , \new_[8636]_ , \new_[8637]_ ,
    \new_[8638]_ , \new_[8639]_ , \new_[8640]_ , \new_[8641]_ ,
    \new_[8642]_ , \new_[8643]_ , \new_[8644]_ , \new_[8645]_ ,
    \new_[8646]_ , \new_[8647]_ , \new_[8648]_ , \new_[8649]_ ,
    \new_[8650]_ , \new_[8651]_ , \new_[8652]_ , \new_[8653]_ ,
    \new_[8654]_ , \new_[8655]_ , \new_[8656]_ , \new_[8657]_ ,
    \new_[8658]_ , \new_[8659]_ , \new_[8660]_ , \new_[8661]_ ,
    \new_[8662]_ , \new_[8663]_ , \new_[8664]_ , \new_[8665]_ ,
    \new_[8666]_ , \new_[8667]_ , \new_[8668]_ , \new_[8669]_ ,
    \new_[8670]_ , \new_[8671]_ , \new_[8672]_ , \new_[8673]_ ,
    \new_[8674]_ , \new_[8675]_ , \new_[8676]_ , \new_[8677]_ ,
    \new_[8678]_ , \new_[8679]_ , \new_[8681]_ , \new_[8682]_ ,
    \new_[8683]_ , \new_[8684]_ , \new_[8685]_ , \new_[8686]_ ,
    \new_[8687]_ , \new_[8688]_ , \new_[8689]_ , \new_[8690]_ ,
    \new_[8691]_ , \new_[8692]_ , \new_[8693]_ , \new_[8694]_ ,
    \new_[8695]_ , \new_[8696]_ , \new_[8697]_ , \new_[8698]_ ,
    \new_[8700]_ , \new_[8703]_ , \new_[8704]_ , \new_[8705]_ ,
    \new_[8706]_ , \new_[8707]_ , \new_[8708]_ , \new_[8709]_ ,
    \new_[8710]_ , \new_[8711]_ , \new_[8712]_ , \new_[8713]_ ,
    \new_[8714]_ , \new_[8715]_ , \new_[8716]_ , \new_[8717]_ ,
    \new_[8718]_ , \new_[8719]_ , \new_[8720]_ , \new_[8721]_ ,
    \new_[8722]_ , \new_[8723]_ , \new_[8724]_ , \new_[8725]_ ,
    \new_[8726]_ , \new_[8727]_ , \new_[8728]_ , \new_[8729]_ ,
    \new_[8730]_ , \new_[8731]_ , \new_[8732]_ , \new_[8733]_ ,
    \new_[8734]_ , \new_[8735]_ , \new_[8736]_ , \new_[8737]_ ,
    \new_[8738]_ , \new_[8739]_ , \new_[8740]_ , \new_[8741]_ ,
    \new_[8742]_ , \new_[8743]_ , \new_[8744]_ , \new_[8745]_ ,
    \new_[8746]_ , \new_[8747]_ , \new_[8748]_ , \new_[8749]_ ,
    \new_[8750]_ , \new_[8751]_ , \new_[8752]_ , \new_[8753]_ ,
    \new_[8754]_ , \new_[8755]_ , \new_[8756]_ , \new_[8757]_ ,
    \new_[8758]_ , \new_[8759]_ , \new_[8760]_ , \new_[8761]_ ,
    \new_[8762]_ , \new_[8763]_ , \new_[8764]_ , \new_[8765]_ ,
    \new_[8766]_ , \new_[8767]_ , \new_[8768]_ , \new_[8769]_ ,
    \new_[8770]_ , \new_[8771]_ , \new_[8772]_ , \new_[8773]_ ,
    \new_[8774]_ , \new_[8775]_ , \new_[8776]_ , \new_[8777]_ ,
    \new_[8778]_ , \new_[8779]_ , \new_[8780]_ , \new_[8781]_ ,
    \new_[8782]_ , \new_[8783]_ , \new_[8784]_ , \new_[8785]_ ,
    \new_[8786]_ , \new_[8787]_ , \new_[8788]_ , \new_[8789]_ ,
    \new_[8790]_ , \new_[8791]_ , \new_[8792]_ , \new_[8793]_ ,
    \new_[8794]_ , \new_[8795]_ , \new_[8796]_ , \new_[8797]_ ,
    \new_[8798]_ , \new_[8799]_ , \new_[8800]_ , \new_[8801]_ ,
    \new_[8802]_ , \new_[8803]_ , \new_[8804]_ , \new_[8805]_ ,
    \new_[8806]_ , \new_[8807]_ , \new_[8808]_ , \new_[8809]_ ,
    \new_[8810]_ , \new_[8811]_ , \new_[8812]_ , \new_[8813]_ ,
    \new_[8814]_ , \new_[8815]_ , \new_[8816]_ , \new_[8817]_ ,
    \new_[8818]_ , \new_[8819]_ , \new_[8820]_ , \new_[8821]_ ,
    \new_[8822]_ , \new_[8823]_ , \new_[8824]_ , \new_[8825]_ ,
    \new_[8826]_ , \new_[8827]_ , \new_[8828]_ , \new_[8829]_ ,
    \new_[8830]_ , \new_[8831]_ , \new_[8832]_ , \new_[8833]_ ,
    \new_[8834]_ , \new_[8835]_ , \new_[8836]_ , \new_[8837]_ ,
    \new_[8838]_ , \new_[8839]_ , \new_[8840]_ , \new_[8841]_ ,
    \new_[8842]_ , \new_[8843]_ , \new_[8844]_ , \new_[8845]_ ,
    \new_[8846]_ , \new_[8847]_ , \new_[8848]_ , \new_[8849]_ ,
    \new_[8850]_ , \new_[8851]_ , \new_[8852]_ , \new_[8853]_ ,
    \new_[8854]_ , \new_[8855]_ , \new_[8856]_ , \new_[8857]_ ,
    \new_[8858]_ , \new_[8859]_ , \new_[8860]_ , \new_[8861]_ ,
    \new_[8862]_ , \new_[8863]_ , \new_[8864]_ , \new_[8865]_ ,
    \new_[8866]_ , \new_[8867]_ , \new_[8868]_ , \new_[8869]_ ,
    \new_[8870]_ , \new_[8871]_ , \new_[8872]_ , \new_[8873]_ ,
    \new_[8874]_ , \new_[8875]_ , \new_[8876]_ , \new_[8877]_ ,
    \new_[8878]_ , \new_[8879]_ , \new_[8880]_ , \new_[8881]_ ,
    \new_[8882]_ , \new_[8883]_ , \new_[8884]_ , \new_[8885]_ ,
    \new_[8886]_ , \new_[8887]_ , \new_[8888]_ , \new_[8889]_ ,
    \new_[8890]_ , \new_[8891]_ , \new_[8892]_ , \new_[8893]_ ,
    \new_[8894]_ , \new_[8895]_ , \new_[8896]_ , \new_[8897]_ ,
    \new_[8898]_ , \new_[8899]_ , \new_[8900]_ , \new_[8901]_ ,
    \new_[8902]_ , \new_[8903]_ , \new_[8904]_ , \new_[8905]_ ,
    \new_[8906]_ , \new_[8907]_ , \new_[8908]_ , \new_[8909]_ ,
    \new_[8910]_ , \new_[8911]_ , \new_[8912]_ , \new_[8913]_ ,
    \new_[8914]_ , \new_[8915]_ , \new_[8916]_ , \new_[8917]_ ,
    \new_[8918]_ , \new_[8919]_ , \new_[8920]_ , \new_[8921]_ ,
    \new_[8922]_ , \new_[8923]_ , \new_[8924]_ , \new_[8925]_ ,
    \new_[8926]_ , \new_[8927]_ , \new_[8928]_ , \new_[8929]_ ,
    \new_[8930]_ , \new_[8931]_ , \new_[8932]_ , \new_[8933]_ ,
    \new_[8934]_ , \new_[8935]_ , \new_[8936]_ , \new_[8937]_ ,
    \new_[8938]_ , \new_[8939]_ , \new_[8940]_ , \new_[8941]_ ,
    \new_[8942]_ , \new_[8943]_ , \new_[8944]_ , \new_[8945]_ ,
    \new_[8946]_ , \new_[8947]_ , \new_[8948]_ , \new_[8949]_ ,
    \new_[8950]_ , \new_[8951]_ , \new_[8952]_ , \new_[8953]_ ,
    \new_[8954]_ , \new_[8955]_ , \new_[8956]_ , \new_[8957]_ ,
    \new_[8958]_ , \new_[8959]_ , \new_[8960]_ , \new_[8961]_ ,
    \new_[8962]_ , \new_[8963]_ , \new_[8964]_ , \new_[8965]_ ,
    \new_[8966]_ , \new_[8967]_ , \new_[8968]_ , \new_[8969]_ ,
    \new_[8970]_ , \new_[8971]_ , \new_[8972]_ , \new_[8973]_ ,
    \new_[8974]_ , \new_[8975]_ , \new_[8976]_ , \new_[8977]_ ,
    \new_[8978]_ , \new_[8979]_ , \new_[8980]_ , \new_[8981]_ ,
    \new_[8982]_ , \new_[8983]_ , \new_[8984]_ , \new_[8985]_ ,
    \new_[8986]_ , \new_[8987]_ , \new_[8988]_ , \new_[8989]_ ,
    \new_[8990]_ , \new_[8991]_ , \new_[8992]_ , \new_[8993]_ ,
    \new_[8994]_ , \new_[8995]_ , \new_[8996]_ , \new_[8997]_ ,
    \new_[8998]_ , \new_[8999]_ , \new_[9000]_ , \new_[9001]_ ,
    \new_[9002]_ , \new_[9003]_ , \new_[9004]_ , \new_[9005]_ ,
    \new_[9006]_ , \new_[9007]_ , \new_[9008]_ , \new_[9009]_ ,
    \new_[9010]_ , \new_[9011]_ , \new_[9012]_ , \new_[9013]_ ,
    \new_[9014]_ , \new_[9015]_ , \new_[9016]_ , \new_[9017]_ ,
    \new_[9018]_ , \new_[9019]_ , \new_[9020]_ , \new_[9021]_ ,
    \new_[9022]_ , \new_[9023]_ , \new_[9024]_ , \new_[9025]_ ,
    \new_[9026]_ , \new_[9027]_ , \new_[9028]_ , \new_[9029]_ ,
    \new_[9030]_ , \new_[9031]_ , \new_[9032]_ , \new_[9033]_ ,
    \new_[9034]_ , \new_[9035]_ , \new_[9036]_ , \new_[9037]_ ,
    \new_[9038]_ , \new_[9039]_ , \new_[9040]_ , \new_[9041]_ ,
    \new_[9042]_ , \new_[9043]_ , \new_[9044]_ , \new_[9045]_ ,
    \new_[9046]_ , \new_[9047]_ , \new_[9048]_ , \new_[9049]_ ,
    \new_[9050]_ , \new_[9051]_ , \new_[9052]_ , \new_[9053]_ ,
    \new_[9054]_ , \new_[9055]_ , \new_[9056]_ , \new_[9057]_ ,
    \new_[9058]_ , \new_[9059]_ , \new_[9060]_ , \new_[9061]_ ,
    \new_[9062]_ , \new_[9063]_ , \new_[9064]_ , \new_[9065]_ ,
    \new_[9066]_ , \new_[9067]_ , \new_[9068]_ , \new_[9069]_ ,
    \new_[9070]_ , \new_[9071]_ , \new_[9072]_ , \new_[9073]_ ,
    \new_[9074]_ , \new_[9075]_ , \new_[9076]_ , \new_[9077]_ ,
    \new_[9078]_ , \new_[9079]_ , \new_[9080]_ , \new_[9081]_ ,
    \new_[9082]_ , \new_[9083]_ , \new_[9084]_ , \new_[9085]_ ,
    \new_[9086]_ , \new_[9087]_ , \new_[9088]_ , \new_[9089]_ ,
    \new_[9090]_ , \new_[9091]_ , \new_[9092]_ , \new_[9093]_ ,
    \new_[9094]_ , \new_[9095]_ , \new_[9096]_ , \new_[9097]_ ,
    \new_[9098]_ , \new_[9099]_ , \new_[9100]_ , \new_[9101]_ ,
    \new_[9102]_ , \new_[9127]_ , \new_[9128]_ , \new_[9132]_ ,
    \new_[9133]_ , \new_[9134]_ , \new_[9135]_ , \new_[9136]_ ,
    \new_[9137]_ , \new_[9138]_ , \new_[9139]_ , \new_[9140]_ ,
    \new_[9141]_ , \new_[9142]_ , \new_[9143]_ , \new_[9144]_ ,
    \new_[9145]_ , \new_[9146]_ , \new_[9147]_ , \new_[9148]_ ,
    \new_[9149]_ , \new_[9150]_ , \new_[9151]_ , \new_[9152]_ ,
    \new_[9153]_ , \new_[9154]_ , \new_[9155]_ , \new_[9156]_ ,
    \new_[9157]_ , \new_[9158]_ , \new_[9159]_ , \new_[9160]_ ,
    \new_[9161]_ , \new_[9162]_ , \new_[9163]_ , \new_[9164]_ ,
    \new_[9165]_ , \new_[9166]_ , \new_[9167]_ , \new_[9168]_ ,
    \new_[9169]_ , \new_[9170]_ , \new_[9171]_ , \new_[9172]_ ,
    \new_[9173]_ , \new_[9174]_ , \new_[9175]_ , \new_[9176]_ ,
    \new_[9177]_ , \new_[9178]_ , \new_[9179]_ , \new_[9180]_ ,
    \new_[9181]_ , \new_[9182]_ , \new_[9183]_ , \new_[9184]_ ,
    \new_[9185]_ , \new_[9186]_ , \new_[9187]_ , \new_[9188]_ ,
    \new_[9189]_ , \new_[9190]_ , \new_[9191]_ , \new_[9192]_ ,
    \new_[9193]_ , \new_[9194]_ , \new_[9195]_ , \new_[9196]_ ,
    \new_[9197]_ , \new_[9198]_ , \new_[9199]_ , \new_[9200]_ ,
    \new_[9201]_ , \new_[9202]_ , \new_[9203]_ , \new_[9204]_ ,
    \new_[9205]_ , \new_[9206]_ , \new_[9207]_ , \new_[9208]_ ,
    \new_[9216]_ , \new_[9217]_ , \new_[9218]_ , \new_[9219]_ ,
    \new_[9220]_ , \new_[9221]_ , \new_[9222]_ , \new_[9223]_ ,
    \new_[9224]_ , \new_[9225]_ , \new_[9226]_ , \new_[9227]_ ,
    \new_[9228]_ , \new_[9229]_ , \new_[9230]_ , \new_[9231]_ ,
    \new_[9232]_ , \new_[9233]_ , \new_[9234]_ , \new_[9235]_ ,
    \new_[9236]_ , \new_[9237]_ , \new_[9238]_ , \new_[9239]_ ,
    \new_[9240]_ , \new_[9241]_ , \new_[9242]_ , \new_[9243]_ ,
    \new_[9244]_ , \new_[9245]_ , \new_[9246]_ , \new_[9247]_ ,
    \new_[9248]_ , \new_[9249]_ , \new_[9250]_ , \new_[9251]_ ,
    \new_[9252]_ , \new_[9253]_ , \new_[9268]_ , \new_[9269]_ ,
    \new_[9270]_ , \new_[9271]_ , \new_[9272]_ , \new_[9273]_ ,
    \new_[9275]_ , \new_[9276]_ , \new_[9277]_ , \new_[9280]_ ,
    \new_[9281]_ , \new_[9282]_ , \new_[9283]_ , \new_[9284]_ ,
    \new_[9285]_ , \new_[9286]_ , \new_[9287]_ , \new_[9288]_ ,
    \new_[9289]_ , \new_[9290]_ , \new_[9291]_ , \new_[9292]_ ,
    \new_[9293]_ , \new_[9294]_ , \new_[9295]_ , \new_[9296]_ ,
    \new_[9297]_ , \new_[9298]_ , \new_[9299]_ , \new_[9300]_ ,
    \new_[9301]_ , \new_[9302]_ , \new_[9303]_ , \new_[9304]_ ,
    \new_[9305]_ , \new_[9307]_ , \new_[9310]_ , \new_[9311]_ ,
    \new_[9312]_ , \new_[9313]_ , \new_[9314]_ , \new_[9315]_ ,
    \new_[9316]_ , \new_[9317]_ , \new_[9318]_ , \new_[9319]_ ,
    \new_[9320]_ , \new_[9321]_ , \new_[9322]_ , \new_[9323]_ ,
    \new_[9324]_ , \new_[9325]_ , \new_[9326]_ , \new_[9327]_ ,
    \new_[9328]_ , \new_[9329]_ , \new_[9330]_ , \new_[9331]_ ,
    \new_[9332]_ , \new_[9333]_ , \new_[9334]_ , \new_[9335]_ ,
    \new_[9336]_ , \new_[9337]_ , \new_[9338]_ , \new_[9339]_ ,
    \new_[9340]_ , \new_[9341]_ , \new_[9342]_ , \new_[9343]_ ,
    \new_[9344]_ , \new_[9345]_ , \new_[9346]_ , \new_[9347]_ ,
    \new_[9348]_ , \new_[9349]_ , \new_[9350]_ , \new_[9351]_ ,
    \new_[9352]_ , \new_[9353]_ , \new_[9354]_ , \new_[9355]_ ,
    \new_[9356]_ , \new_[9357]_ , \new_[9358]_ , \new_[9359]_ ,
    \new_[9360]_ , \new_[9361]_ , \new_[9362]_ , \new_[9363]_ ,
    \new_[9364]_ , \new_[9365]_ , \new_[9366]_ , \new_[9367]_ ,
    \new_[9368]_ , \new_[9369]_ , \new_[9370]_ , \new_[9371]_ ,
    \new_[9372]_ , \new_[9373]_ , \new_[9374]_ , \new_[9375]_ ,
    \new_[9376]_ , \new_[9377]_ , \new_[9378]_ , \new_[9379]_ ,
    \new_[9380]_ , \new_[9381]_ , \new_[9382]_ , \new_[9383]_ ,
    \new_[9384]_ , \new_[9385]_ , \new_[9386]_ , \new_[9387]_ ,
    \new_[9388]_ , \new_[9389]_ , \new_[9390]_ , \new_[9391]_ ,
    \new_[9392]_ , \new_[9393]_ , \new_[9394]_ , \new_[9395]_ ,
    \new_[9396]_ , \new_[9397]_ , \new_[9398]_ , \new_[9399]_ ,
    \new_[9400]_ , \new_[9401]_ , \new_[9402]_ , \new_[9403]_ ,
    \new_[9404]_ , \new_[9405]_ , \new_[9406]_ , \new_[9407]_ ,
    \new_[9408]_ , \new_[9409]_ , \new_[9410]_ , \new_[9411]_ ,
    \new_[9412]_ , \new_[9413]_ , \new_[9414]_ , \new_[9415]_ ,
    \new_[9416]_ , \new_[9417]_ , \new_[9418]_ , \new_[9419]_ ,
    \new_[9420]_ , \new_[9421]_ , \new_[9422]_ , \new_[9423]_ ,
    \new_[9424]_ , \new_[9425]_ , \new_[9426]_ , \new_[9427]_ ,
    \new_[9428]_ , \new_[9429]_ , \new_[9430]_ , \new_[9431]_ ,
    \new_[9432]_ , \new_[9433]_ , \new_[9434]_ , \new_[9435]_ ,
    \new_[9436]_ , \new_[9437]_ , \new_[9438]_ , \new_[9439]_ ,
    \new_[9440]_ , \new_[9441]_ , \new_[9442]_ , \new_[9443]_ ,
    \new_[9444]_ , \new_[9445]_ , \new_[9446]_ , \new_[9447]_ ,
    \new_[9448]_ , \new_[9449]_ , \new_[9450]_ , \new_[9451]_ ,
    \new_[9452]_ , \new_[9453]_ , \new_[9462]_ , \new_[9463]_ ,
    \new_[9464]_ , \new_[9465]_ , \new_[9466]_ , \new_[9467]_ ,
    \new_[9468]_ , \new_[9469]_ , \new_[9470]_ , \new_[9471]_ ,
    \new_[9472]_ , \new_[9476]_ , \new_[9477]_ , \new_[9478]_ ,
    \new_[9479]_ , \new_[9480]_ , \new_[9481]_ , \new_[9482]_ ,
    \new_[9483]_ , \new_[9484]_ , \new_[9485]_ , \new_[9487]_ ,
    \new_[9488]_ , \new_[9490]_ , \new_[9491]_ , \new_[9492]_ ,
    \new_[9493]_ , \new_[9496]_ , \new_[9497]_ , \new_[9498]_ ,
    \new_[9499]_ , \new_[9500]_ , \new_[9501]_ , \new_[9502]_ ,
    \new_[9503]_ , \new_[9504]_ , \new_[9505]_ , \new_[9506]_ ,
    \new_[9507]_ , \new_[9508]_ , \new_[9509]_ , \new_[9510]_ ,
    \new_[9511]_ , \new_[9512]_ , \new_[9513]_ , \new_[9529]_ ,
    \new_[9530]_ , \new_[9531]_ , \new_[9532]_ , \new_[9533]_ ,
    \new_[9534]_ , \new_[9535]_ , \new_[9536]_ , \new_[9537]_ ,
    \new_[9538]_ , \new_[9539]_ , \new_[9540]_ , \new_[9541]_ ,
    \new_[9542]_ , \new_[9543]_ , \new_[9544]_ , \new_[9545]_ ,
    \new_[9546]_ , \new_[9547]_ , \new_[9548]_ , \new_[9549]_ ,
    \new_[9550]_ , \new_[9551]_ , \new_[9552]_ , \new_[9553]_ ,
    \new_[9554]_ , \new_[9555]_ , \new_[9556]_ , \new_[9557]_ ,
    \new_[9558]_ , \new_[9559]_ , \new_[9560]_ , \new_[9561]_ ,
    \new_[9562]_ , \new_[9565]_ , \new_[9567]_ , \new_[9568]_ ,
    \new_[9569]_ , \new_[9570]_ , \new_[9571]_ , \new_[9572]_ ,
    \new_[9573]_ , \new_[9574]_ , \new_[9575]_ , \new_[9576]_ ,
    \new_[9587]_ , \new_[9588]_ , \new_[9590]_ , \new_[9591]_ ,
    \new_[9592]_ , \new_[9593]_ , \new_[9594]_ , \new_[9595]_ ,
    \new_[9596]_ , \new_[9597]_ , \new_[9598]_ , \new_[9599]_ ,
    \new_[9600]_ , \new_[9601]_ , \new_[9602]_ , \new_[9603]_ ,
    \new_[9604]_ , \new_[9605]_ , \new_[9606]_ , \new_[9607]_ ,
    \new_[9608]_ , \new_[9609]_ , \new_[9610]_ , \new_[9611]_ ,
    \new_[9612]_ , \new_[9613]_ , \new_[9614]_ , \new_[9615]_ ,
    \new_[9616]_ , \new_[9617]_ , \new_[9618]_ , \new_[9619]_ ,
    \new_[9620]_ , \new_[9621]_ , \new_[9622]_ , \new_[9623]_ ,
    \new_[9624]_ , \new_[9625]_ , \new_[9626]_ , \new_[9627]_ ,
    \new_[9628]_ , \new_[9629]_ , \new_[9630]_ , \new_[9631]_ ,
    \new_[9632]_ , \new_[9633]_ , \new_[9634]_ , \new_[9635]_ ,
    \new_[9636]_ , \new_[9637]_ , \new_[9638]_ , \new_[9639]_ ,
    \new_[9640]_ , \new_[9641]_ , \new_[9642]_ , \new_[9643]_ ,
    \new_[9644]_ , \new_[9646]_ , \new_[9647]_ , \new_[9650]_ ,
    \new_[9651]_ , \new_[9652]_ , \new_[9653]_ , \new_[9654]_ ,
    \new_[9655]_ , \new_[9656]_ , \new_[9657]_ , \new_[9658]_ ,
    \new_[9659]_ , \new_[9660]_ , \new_[9661]_ , \new_[9662]_ ,
    \new_[9663]_ , \new_[9664]_ , \new_[9665]_ , \new_[9666]_ ,
    \new_[9667]_ , \new_[9668]_ , \new_[9669]_ , \new_[9670]_ ,
    \new_[9671]_ , \new_[9672]_ , \new_[9673]_ , \new_[9674]_ ,
    \new_[9675]_ , \new_[9676]_ , \new_[9677]_ , \new_[9678]_ ,
    \new_[9679]_ , \new_[9680]_ , \new_[9681]_ , \new_[9682]_ ,
    \new_[9683]_ , \new_[9685]_ , \new_[9686]_ , \new_[9687]_ ,
    \new_[9688]_ , \new_[9689]_ , \new_[9690]_ , \new_[9691]_ ,
    \new_[9692]_ , \new_[9693]_ , \new_[9694]_ , \new_[9695]_ ,
    \new_[9696]_ , \new_[9697]_ , \new_[9698]_ , \new_[9699]_ ,
    \new_[9700]_ , \new_[9701]_ , \new_[9702]_ , \new_[9703]_ ,
    \new_[9704]_ , \new_[9705]_ , \new_[9706]_ , \new_[9707]_ ,
    \new_[9708]_ , \new_[9709]_ , \new_[9710]_ , \new_[9711]_ ,
    \new_[9712]_ , \new_[9713]_ , \new_[9714]_ , \new_[9715]_ ,
    \new_[9716]_ , \new_[9717]_ , \new_[9718]_ , \new_[9719]_ ,
    \new_[9720]_ , \new_[9721]_ , \new_[9722]_ , \new_[9723]_ ,
    \new_[9724]_ , \new_[9725]_ , \new_[9726]_ , \new_[9727]_ ,
    \new_[9728]_ , \new_[9729]_ , \new_[9730]_ , \new_[9731]_ ,
    \new_[9732]_ , \new_[9733]_ , \new_[9734]_ , \new_[9735]_ ,
    \new_[9736]_ , \new_[9737]_ , \new_[9738]_ , \new_[9739]_ ,
    \new_[9740]_ , \new_[9741]_ , \new_[9742]_ , \new_[9743]_ ,
    \new_[9744]_ , \new_[9745]_ , \new_[9746]_ , \new_[9747]_ ,
    \new_[9748]_ , \new_[9749]_ , \new_[9750]_ , \new_[9751]_ ,
    \new_[9752]_ , \new_[9753]_ , \new_[9754]_ , \new_[9755]_ ,
    \new_[9756]_ , \new_[9757]_ , \new_[9758]_ , \new_[9760]_ ,
    \new_[9761]_ , \new_[9762]_ , \new_[9763]_ , \new_[9764]_ ,
    \new_[9765]_ , \new_[9766]_ , \new_[9767]_ , \new_[9768]_ ,
    \new_[9769]_ , \new_[9770]_ , \new_[9771]_ , \new_[9772]_ ,
    \new_[9773]_ , \new_[9774]_ , \new_[9775]_ , \new_[9776]_ ,
    \new_[9777]_ , \new_[9778]_ , \new_[9779]_ , \new_[9780]_ ,
    \new_[9781]_ , \new_[9782]_ , \new_[9783]_ , \new_[9784]_ ,
    \new_[9785]_ , \new_[9786]_ , \new_[9787]_ , \new_[9788]_ ,
    \new_[9789]_ , \new_[9790]_ , \new_[9791]_ , \new_[9792]_ ,
    \new_[9793]_ , \new_[9794]_ , \new_[9795]_ , \new_[9796]_ ,
    \new_[9797]_ , \new_[9798]_ , \new_[9799]_ , \new_[9800]_ ,
    \new_[9801]_ , \new_[9802]_ , \new_[9803]_ , \new_[9804]_ ,
    \new_[9805]_ , \new_[9806]_ , \new_[9807]_ , \new_[9808]_ ,
    \new_[9809]_ , \new_[9810]_ , \new_[9811]_ , \new_[9812]_ ,
    \new_[9813]_ , \new_[9814]_ , \new_[9815]_ , \new_[9816]_ ,
    \new_[9817]_ , \new_[9818]_ , \new_[9819]_ , \new_[9820]_ ,
    \new_[9821]_ , \new_[9822]_ , \new_[9823]_ , \new_[9824]_ ,
    \new_[9825]_ , \new_[9826]_ , \new_[9827]_ , \new_[9828]_ ,
    \new_[9829]_ , \new_[9830]_ , \new_[9833]_ , \new_[9834]_ ,
    \new_[9836]_ , \new_[9837]_ , \new_[9838]_ , \new_[9839]_ ,
    \new_[9840]_ , \new_[9841]_ , \new_[9842]_ , \new_[9846]_ ,
    \new_[9847]_ , \new_[9853]_ , \new_[9854]_ , \new_[9855]_ ,
    \new_[9856]_ , \new_[9857]_ , \new_[9877]_ , \new_[9878]_ ,
    \new_[9879]_ , \new_[9880]_ , \new_[9881]_ , \new_[9884]_ ,
    \new_[9885]_ , \new_[9886]_ , \new_[9887]_ , \new_[9888]_ ,
    \new_[9895]_ , \new_[9896]_ , \new_[9899]_ , \new_[9900]_ ,
    \new_[9901]_ , \new_[9902]_ , \new_[9903]_ , \new_[9904]_ ,
    \new_[9905]_ , \new_[9906]_ , \new_[9907]_ , \new_[9908]_ ,
    \new_[9910]_ , \new_[9915]_ , \new_[9918]_ , \new_[9919]_ ,
    \new_[9931]_ , \new_[9968]_ , \new_[9970]_ , \new_[9971]_ ,
    \new_[9972]_ , \new_[9979]_ , \new_[9980]_ , \new_[9982]_ ,
    \new_[9983]_ , \new_[9985]_ , \new_[9986]_ , \new_[9987]_ ,
    \new_[9988]_ , \new_[9989]_ , \new_[9991]_ , \new_[9992]_ ,
    \new_[9993]_ , \new_[9994]_ , \new_[9995]_ , \new_[9996]_ ,
    \new_[9997]_ , \new_[9998]_ , \new_[10000]_ , \new_[10001]_ ,
    \new_[10002]_ , \new_[10003]_ , \new_[10004]_ , \new_[10005]_ ,
    \new_[10006]_ , \new_[10007]_ , \new_[10008]_ , \new_[10009]_ ,
    \new_[10010]_ , \new_[10011]_ , \new_[10012]_ , \new_[10013]_ ,
    \new_[10016]_ , \new_[10017]_ , \new_[10018]_ , \new_[10019]_ ,
    \new_[10020]_ , \new_[10021]_ , \new_[10022]_ , \new_[10023]_ ,
    \new_[10025]_ , \new_[10026]_ , \new_[10027]_ , \new_[10028]_ ,
    \new_[10029]_ , \new_[10030]_ , \new_[10031]_ , \new_[10032]_ ,
    \new_[10033]_ , \new_[10034]_ , \new_[10035]_ , \new_[10036]_ ,
    \new_[10037]_ , \new_[10038]_ , \new_[10039]_ , \new_[10040]_ ,
    \new_[10041]_ , \new_[10042]_ , \new_[10043]_ , \new_[10046]_ ,
    \new_[10047]_ , \new_[10048]_ , \new_[10049]_ , \new_[10050]_ ,
    \new_[10051]_ , \new_[10052]_ , \new_[10053]_ , \new_[10054]_ ,
    \new_[10055]_ , \new_[10056]_ , \new_[10057]_ , \new_[10058]_ ,
    \new_[10059]_ , \new_[10060]_ , \new_[10061]_ , \new_[10062]_ ,
    \new_[10063]_ , \new_[10064]_ , \new_[10065]_ , \new_[10066]_ ,
    \new_[10068]_ , \new_[10069]_ , \new_[10072]_ , \new_[10073]_ ,
    \new_[10074]_ , \new_[10075]_ , \new_[10076]_ , \new_[10077]_ ,
    \new_[10078]_ , \new_[10079]_ , \new_[10080]_ , \new_[10081]_ ,
    \new_[10082]_ , \new_[10083]_ , \new_[10084]_ , \new_[10085]_ ,
    \new_[10086]_ , \new_[10087]_ , \new_[10088]_ , \new_[10089]_ ,
    \new_[10090]_ , \new_[10091]_ , \new_[10092]_ , \new_[10093]_ ,
    \new_[10094]_ , \new_[10095]_ , \new_[10096]_ , \new_[10097]_ ,
    \new_[10098]_ , \new_[10099]_ , \new_[10100]_ , \new_[10101]_ ,
    \new_[10102]_ , \new_[10103]_ , \new_[10104]_ , \new_[10105]_ ,
    \new_[10106]_ , \new_[10107]_ , \new_[10108]_ , \new_[10109]_ ,
    \new_[10110]_ , \new_[10111]_ , \new_[10112]_ , \new_[10113]_ ,
    \new_[10114]_ , \new_[10115]_ , \new_[10116]_ , \new_[10117]_ ,
    \new_[10118]_ , \new_[10119]_ , \new_[10120]_ , \new_[10121]_ ,
    \new_[10122]_ , \new_[10123]_ , \new_[10124]_ , \new_[10125]_ ,
    \new_[10126]_ , \new_[10127]_ , \new_[10128]_ , \new_[10129]_ ,
    \new_[10130]_ , \new_[10131]_ , \new_[10132]_ , \new_[10133]_ ,
    \new_[10134]_ , \new_[10135]_ , \new_[10136]_ , \new_[10137]_ ,
    \new_[10138]_ , \new_[10139]_ , \new_[10140]_ , \new_[10141]_ ,
    \new_[10142]_ , \new_[10143]_ , \new_[10144]_ , \new_[10145]_ ,
    \new_[10146]_ , \new_[10147]_ , \new_[10148]_ , \new_[10149]_ ,
    \new_[10150]_ , \new_[10151]_ , \new_[10152]_ , \new_[10153]_ ,
    \new_[10154]_ , \new_[10155]_ , \new_[10156]_ , \new_[10157]_ ,
    \new_[10158]_ , \new_[10159]_ , \new_[10160]_ , \new_[10161]_ ,
    \new_[10162]_ , \new_[10163]_ , \new_[10164]_ , \new_[10165]_ ,
    \new_[10166]_ , \new_[10167]_ , \new_[10168]_ , \new_[10169]_ ,
    \new_[10170]_ , \new_[10171]_ , \new_[10172]_ , \new_[10173]_ ,
    \new_[10174]_ , \new_[10175]_ , \new_[10176]_ , \new_[10177]_ ,
    \new_[10178]_ , \new_[10179]_ , \new_[10180]_ , \new_[10181]_ ,
    \new_[10182]_ , \new_[10183]_ , \new_[10184]_ , \new_[10185]_ ,
    \new_[10186]_ , \new_[10187]_ , \new_[10188]_ , \new_[10189]_ ,
    \new_[10190]_ , \new_[10191]_ , \new_[10192]_ , \new_[10193]_ ,
    \new_[10194]_ , \new_[10195]_ , \new_[10196]_ , \new_[10197]_ ,
    \new_[10198]_ , \new_[10199]_ , \new_[10200]_ , \new_[10201]_ ,
    \new_[10202]_ , \new_[10203]_ , \new_[10204]_ , \new_[10205]_ ,
    \new_[10206]_ , \new_[10207]_ , \new_[10208]_ , \new_[10209]_ ,
    \new_[10210]_ , \new_[10211]_ , \new_[10212]_ , \new_[10213]_ ,
    \new_[10214]_ , \new_[10215]_ , \new_[10216]_ , \new_[10217]_ ,
    \new_[10218]_ , \new_[10219]_ , \new_[10220]_ , \new_[10221]_ ,
    \new_[10222]_ , \new_[10223]_ , \new_[10224]_ , \new_[10225]_ ,
    \new_[10226]_ , \new_[10227]_ , \new_[10228]_ , \new_[10229]_ ,
    \new_[10230]_ , \new_[10231]_ , \new_[10232]_ , \new_[10233]_ ,
    \new_[10234]_ , \new_[10235]_ , \new_[10236]_ , \new_[10237]_ ,
    \new_[10238]_ , \new_[10239]_ , \new_[10240]_ , \new_[10241]_ ,
    \new_[10242]_ , \new_[10243]_ , \new_[10244]_ , \new_[10245]_ ,
    \new_[10246]_ , \new_[10247]_ , \new_[10249]_ , \new_[10250]_ ,
    \new_[10251]_ , \new_[10252]_ , \new_[10253]_ , \new_[10254]_ ,
    \new_[10255]_ , \new_[10256]_ , \new_[10258]_ , \new_[10259]_ ,
    \new_[10260]_ , \new_[10261]_ , \new_[10262]_ , \new_[10263]_ ,
    \new_[10264]_ , \new_[10265]_ , \new_[10266]_ , \new_[10267]_ ,
    \new_[10268]_ , \new_[10269]_ , \new_[10270]_ , \new_[10271]_ ,
    \new_[10272]_ , \new_[10273]_ , \new_[10274]_ , \new_[10275]_ ,
    \new_[10276]_ , \new_[10277]_ , \new_[10278]_ , \new_[10279]_ ,
    \new_[10280]_ , \new_[10281]_ , \new_[10282]_ , \new_[10283]_ ,
    \new_[10284]_ , \new_[10285]_ , \new_[10286]_ , \new_[10287]_ ,
    \new_[10288]_ , \new_[10289]_ , \new_[10290]_ , \new_[10291]_ ,
    \new_[10292]_ , \new_[10293]_ , \new_[10294]_ , \new_[10295]_ ,
    \new_[10296]_ , \new_[10297]_ , \new_[10298]_ , \new_[10299]_ ,
    \new_[10300]_ , \new_[10301]_ , \new_[10302]_ , \new_[10303]_ ,
    \new_[10304]_ , \new_[10305]_ , \new_[10306]_ , \new_[10307]_ ,
    \new_[10308]_ , \new_[10309]_ , \new_[10310]_ , \new_[10311]_ ,
    \new_[10312]_ , \new_[10313]_ , \new_[10315]_ , \new_[10316]_ ,
    \new_[10317]_ , \new_[10318]_ , \new_[10319]_ , \new_[10320]_ ,
    \new_[10321]_ , \new_[10324]_ , \new_[10325]_ , \new_[10327]_ ,
    \new_[10328]_ , \new_[10329]_ , \new_[10331]_ , \new_[10332]_ ,
    \new_[10335]_ , \new_[10336]_ , \new_[10337]_ , \new_[10338]_ ,
    \new_[10339]_ , \new_[10340]_ , \new_[10341]_ , \new_[10342]_ ,
    \new_[10343]_ , \new_[10344]_ , \new_[10349]_ , \new_[10350]_ ,
    \new_[10351]_ , \new_[10352]_ , \new_[10353]_ , \new_[10354]_ ,
    \new_[10355]_ , \new_[10356]_ , \new_[10357]_ , \new_[10358]_ ,
    \new_[10359]_ , \new_[10360]_ , \new_[10361]_ , \new_[10362]_ ,
    \new_[10363]_ , \new_[10364]_ , \new_[10365]_ , \new_[10366]_ ,
    \new_[10367]_ , \new_[10368]_ , \new_[10369]_ , \new_[10370]_ ,
    \new_[10371]_ , \new_[10372]_ , \new_[10374]_ , \new_[10375]_ ,
    \new_[10376]_ , \new_[10377]_ , \new_[10378]_ , \new_[10379]_ ,
    \new_[10380]_ , \new_[10381]_ , \new_[10382]_ , \new_[10383]_ ,
    \new_[10384]_ , \new_[10385]_ , \new_[10386]_ , \new_[10387]_ ,
    \new_[10388]_ , \new_[10389]_ , \new_[10390]_ , \new_[10391]_ ,
    \new_[10392]_ , \new_[10393]_ , \new_[10394]_ , \new_[10395]_ ,
    \new_[10396]_ , \new_[10398]_ , \new_[10399]_ , \new_[10401]_ ,
    \new_[10402]_ , \new_[10403]_ , \new_[10404]_ , \new_[10405]_ ,
    \new_[10406]_ , \new_[10407]_ , \new_[10408]_ , \new_[10409]_ ,
    \new_[10410]_ , \new_[10411]_ , \new_[10412]_ , \new_[10413]_ ,
    \new_[10414]_ , \new_[10415]_ , \new_[10416]_ , \new_[10417]_ ,
    \new_[10418]_ , \new_[10419]_ , \new_[10420]_ , \new_[10421]_ ,
    \new_[10422]_ , \new_[10423]_ , \new_[10424]_ , \new_[10425]_ ,
    \new_[10426]_ , \new_[10427]_ , \new_[10428]_ , \new_[10429]_ ,
    \new_[10430]_ , \new_[10431]_ , \new_[10432]_ , \new_[10433]_ ,
    \new_[10434]_ , \new_[10435]_ , \new_[10444]_ , \new_[10445]_ ,
    \new_[10446]_ , \new_[10447]_ , \new_[10448]_ , \new_[10449]_ ,
    \new_[10450]_ , \new_[10453]_ , \new_[10455]_ , \new_[10456]_ ,
    \new_[10457]_ , \new_[10458]_ , \new_[10459]_ , \new_[10460]_ ,
    \new_[10461]_ , \new_[10462]_ , \new_[10463]_ , \new_[10464]_ ,
    \new_[10465]_ , \new_[10481]_ , \new_[10483]_ , \new_[10484]_ ,
    \new_[10485]_ , \new_[10486]_ , \new_[10491]_ , \new_[10492]_ ,
    \new_[10493]_ , \new_[10494]_ , \new_[10495]_ , \new_[10496]_ ,
    \new_[10497]_ , \new_[10498]_ , \new_[10499]_ , \new_[10500]_ ,
    \new_[10501]_ , \new_[10502]_ , \new_[10503]_ , \new_[10504]_ ,
    \new_[10505]_ , \new_[10506]_ , \new_[10507]_ , \new_[10508]_ ,
    \new_[10509]_ , \new_[10510]_ , \new_[10511]_ , \new_[10512]_ ,
    \new_[10513]_ , \new_[10514]_ , \new_[10515]_ , \new_[10516]_ ,
    \new_[10517]_ , \new_[10518]_ , \new_[10519]_ , \new_[10520]_ ,
    \new_[10521]_ , \new_[10522]_ , \new_[10523]_ , \new_[10524]_ ,
    \new_[10525]_ , \new_[10526]_ , \new_[10527]_ , \new_[10528]_ ,
    \new_[10529]_ , \new_[10530]_ , \new_[10531]_ , \new_[10532]_ ,
    \new_[10533]_ , \new_[10534]_ , \new_[10535]_ , \new_[10744]_ ,
    \new_[10759]_ , \new_[10773]_ , \new_[10774]_ , \new_[10775]_ ,
    \new_[10794]_ , \new_[10816]_ , \new_[10822]_ , \new_[10823]_ ,
    \new_[10824]_ , \new_[10825]_ , \new_[10826]_ , \new_[10827]_ ,
    \new_[10828]_ , \new_[10829]_ , \new_[10830]_ , \new_[10831]_ ,
    \new_[10835]_ , \new_[10836]_ , \new_[10837]_ , \new_[10838]_ ,
    \new_[10839]_ , \new_[10840]_ , \new_[10841]_ , \new_[10842]_ ,
    \new_[10843]_ , \new_[10844]_ , \new_[10845]_ , \new_[10846]_ ,
    \new_[10847]_ , \new_[10848]_ , \new_[10849]_ , \new_[10850]_ ,
    \new_[10851]_ , \new_[10852]_ , \new_[10853]_ , \new_[10854]_ ,
    \new_[10855]_ , \new_[10857]_ , \new_[10858]_ , \new_[10859]_ ,
    \new_[10860]_ , \new_[10861]_ , \new_[10862]_ , \new_[10863]_ ,
    \new_[10864]_ , \new_[10865]_ , \new_[10866]_ , \new_[10867]_ ,
    \new_[10868]_ , \new_[10869]_ , \new_[10870]_ , \new_[10871]_ ,
    \new_[10872]_ , \new_[10873]_ , \new_[10874]_ , \new_[10875]_ ,
    \new_[10876]_ , \new_[10877]_ , \new_[10878]_ , \new_[10879]_ ,
    \new_[10880]_ , \new_[10881]_ , \new_[10882]_ , \new_[10883]_ ,
    \new_[10884]_ , \new_[10885]_ , \new_[10886]_ , \new_[10887]_ ,
    \new_[10888]_ , \new_[10921]_ , \new_[10922]_ , \new_[10923]_ ,
    \new_[10924]_ , \new_[10925]_ , \new_[10926]_ , \new_[10927]_ ,
    \new_[10928]_ , \new_[10929]_ , \new_[10930]_ , \new_[10931]_ ,
    \new_[10932]_ , \new_[10933]_ , \new_[10934]_ , \new_[10935]_ ,
    \new_[10936]_ , \new_[10937]_ , \new_[10938]_ , \new_[10942]_ ,
    \new_[10947]_ , \new_[10948]_ , \new_[10949]_ , \new_[10950]_ ,
    \new_[10951]_ , \new_[10952]_ , \new_[10954]_ , \new_[10955]_ ,
    \new_[10956]_ , \new_[10958]_ , \new_[10960]_ , \new_[10961]_ ,
    \new_[10962]_ , \new_[10967]_ , \new_[10972]_ , \new_[10973]_ ,
    \new_[10974]_ , \new_[10975]_ , \new_[10976]_ , \new_[10977]_ ,
    \new_[10978]_ , \new_[10979]_ , \new_[10980]_ , \new_[10981]_ ,
    \new_[10982]_ , \new_[10983]_ , \new_[10984]_ , \new_[10985]_ ,
    \new_[10986]_ , \new_[10987]_ , \new_[10988]_ , \new_[10989]_ ,
    \new_[10990]_ , \new_[10991]_ , \new_[10992]_ , \new_[10993]_ ,
    \new_[10994]_ , \new_[10995]_ , \new_[10996]_ , \new_[10997]_ ,
    \new_[10998]_ , \new_[10999]_ , \new_[11000]_ , \new_[11001]_ ,
    \new_[11002]_ , \new_[11003]_ , \new_[11004]_ , \new_[11005]_ ,
    \new_[11006]_ , \new_[11007]_ , \new_[11008]_ , \new_[11009]_ ,
    \new_[11010]_ , \new_[11011]_ , \new_[11012]_ , \new_[11013]_ ,
    \new_[11014]_ , \new_[11016]_ , \new_[11018]_ , \new_[11026]_ ,
    \new_[11027]_ , \new_[11028]_ , \new_[11029]_ , \new_[11031]_ ,
    \new_[11036]_ , \new_[11046]_ , \new_[11047]_ , \new_[11067]_ ,
    \new_[11068]_ , \new_[11069]_ , \new_[11070]_ , \new_[11071]_ ,
    \new_[11072]_ , \new_[11074]_ , \new_[11075]_ , \new_[11077]_ ,
    \new_[11078]_ , \new_[11079]_ , \new_[11080]_ , \new_[11081]_ ,
    \new_[11082]_ , \new_[11083]_ , \new_[11084]_ , \new_[11085]_ ,
    \new_[11086]_ , \new_[11087]_ , \new_[11088]_ , \new_[11089]_ ,
    \new_[11090]_ , \new_[11091]_ , \new_[11092]_ , \new_[11093]_ ,
    \new_[11094]_ , \new_[11095]_ , \new_[11096]_ , \new_[11097]_ ,
    \new_[11098]_ , \new_[11099]_ , \new_[11100]_ , \new_[11101]_ ,
    \new_[11102]_ , \new_[11103]_ , \new_[11104]_ , \new_[11105]_ ,
    \new_[11106]_ , \new_[11107]_ , \new_[11108]_ , \new_[11109]_ ,
    \new_[11110]_ , \new_[11111]_ , \new_[11112]_ , \new_[11113]_ ,
    \new_[11114]_ , \new_[11115]_ , \new_[11116]_ , \new_[11117]_ ,
    \new_[11118]_ , \new_[11119]_ , \new_[11120]_ , \new_[11121]_ ,
    \new_[11122]_ , \new_[11123]_ , \new_[11124]_ , \new_[11125]_ ,
    \new_[11126]_ , \new_[11127]_ , \new_[11128]_ , \new_[11129]_ ,
    \new_[11130]_ , \new_[11131]_ , \new_[11132]_ , \new_[11133]_ ,
    \new_[11134]_ , \new_[11135]_ , \new_[11136]_ , \new_[11137]_ ,
    \new_[11138]_ , \new_[11139]_ , \new_[11140]_ , \new_[11141]_ ,
    \new_[11142]_ , \new_[11143]_ , \new_[11145]_ , \new_[11150]_ ,
    \new_[11151]_ , \new_[11152]_ , \new_[11153]_ , \new_[11154]_ ,
    \new_[11155]_ , \new_[11156]_ , \new_[11157]_ , \new_[11158]_ ,
    \new_[11159]_ , \new_[11160]_ , \new_[11161]_ , \new_[11162]_ ,
    \new_[11163]_ , \new_[11164]_ , \new_[11165]_ , \new_[11166]_ ,
    \new_[11167]_ , \new_[11168]_ , \new_[11169]_ , \new_[11170]_ ,
    \new_[11171]_ , \new_[11172]_ , \new_[11173]_ , \new_[11175]_ ,
    \new_[11176]_ , \new_[11177]_ , \new_[11178]_ , \new_[11203]_ ,
    \new_[11204]_ , \new_[11205]_ , \new_[11206]_ , \new_[11208]_ ,
    \new_[11209]_ , \new_[11210]_ , \new_[11212]_ , \new_[11213]_ ,
    \new_[11214]_ , \new_[11216]_ , \new_[11218]_ , \new_[11220]_ ,
    \new_[11221]_ , \new_[11233]_ , \new_[11235]_ , \new_[11238]_ ,
    \new_[11244]_ , \new_[11245]_ , \new_[11246]_ , \new_[11247]_ ,
    \new_[11248]_ , \new_[11249]_ , \new_[11250]_ , \new_[11251]_ ,
    \new_[11252]_ , \new_[11253]_ , \new_[11254]_ , \new_[11255]_ ,
    \new_[11256]_ , \new_[11257]_ , \new_[11258]_ , \new_[11259]_ ,
    \new_[11260]_ , \new_[11261]_ , \new_[11262]_ , \new_[11263]_ ,
    \new_[11264]_ , \new_[11265]_ , \new_[11266]_ , \new_[11267]_ ,
    \new_[11268]_ , \new_[11269]_ , \new_[11270]_ , \new_[11271]_ ,
    \new_[11272]_ , \new_[11273]_ , \new_[11274]_ , \new_[11275]_ ,
    \new_[11276]_ , \new_[11277]_ , \new_[11278]_ , \new_[11279]_ ,
    \new_[11280]_ , \new_[11281]_ , \new_[11282]_ , \new_[11283]_ ,
    \new_[11284]_ , \new_[11285]_ , \new_[11286]_ , \new_[11287]_ ,
    \new_[11288]_ , \new_[11289]_ , \new_[11290]_ , \new_[11291]_ ,
    \new_[11292]_ , \new_[11293]_ , \new_[11294]_ , \new_[11295]_ ,
    \new_[11296]_ , \new_[11297]_ , \new_[11298]_ , \new_[11299]_ ,
    \new_[11300]_ , \new_[11301]_ , \new_[11302]_ , \new_[11303]_ ,
    \new_[11304]_ , \new_[11305]_ , \new_[11306]_ , \new_[11307]_ ,
    \new_[11308]_ , \new_[11309]_ , \new_[11310]_ , \new_[11311]_ ,
    \new_[11312]_ , \new_[11313]_ , \new_[11314]_ , \new_[11315]_ ,
    \new_[11316]_ , \new_[11317]_ , \new_[11318]_ , \new_[11319]_ ,
    \new_[11320]_ , \new_[11321]_ , \new_[11322]_ , \new_[11323]_ ,
    \new_[11324]_ , \new_[11325]_ , \new_[11326]_ , \new_[11327]_ ,
    \new_[11328]_ , \new_[11329]_ , \new_[11330]_ , \new_[11331]_ ,
    \new_[11332]_ , \new_[11333]_ , \new_[11334]_ , \new_[11336]_ ,
    \new_[11337]_ , \new_[11338]_ , \new_[11339]_ , \new_[11340]_ ,
    \new_[11343]_ , \new_[11344]_ , \new_[11345]_ , \new_[11346]_ ,
    \new_[11347]_ , \new_[11348]_ , \new_[11349]_ , \new_[11350]_ ,
    \new_[11351]_ , \new_[11352]_ , \new_[11353]_ , \new_[11354]_ ,
    \new_[11355]_ , \new_[11356]_ , \new_[11357]_ , \new_[11358]_ ,
    \new_[11359]_ , \new_[11360]_ , \new_[11361]_ , \new_[11362]_ ,
    \new_[11363]_ , \new_[11364]_ , \new_[11365]_ , \new_[11366]_ ,
    \new_[11367]_ , \new_[11368]_ , \new_[11369]_ , \new_[11370]_ ,
    \new_[11371]_ , \new_[11372]_ , \new_[11373]_ , \new_[11374]_ ,
    \new_[11375]_ , \new_[11376]_ , \new_[11377]_ , \new_[11378]_ ,
    \new_[11379]_ , \new_[11380]_ , \new_[11381]_ , \new_[11382]_ ,
    \new_[11383]_ , \new_[11384]_ , \new_[11385]_ , \new_[11386]_ ,
    \new_[11387]_ , \new_[11388]_ , \new_[11389]_ , \new_[11390]_ ,
    \new_[11391]_ , \new_[11392]_ , \new_[11393]_ , \new_[11394]_ ,
    \new_[11395]_ , \new_[11396]_ , \new_[11397]_ , \new_[11398]_ ,
    \new_[11399]_ , \new_[11400]_ , \new_[11401]_ , \new_[11402]_ ,
    \new_[11403]_ , \new_[11404]_ , \new_[11405]_ , \new_[11406]_ ,
    \new_[11407]_ , \new_[11408]_ , \new_[11409]_ , \new_[11410]_ ,
    \new_[11411]_ , \new_[11412]_ , \new_[11413]_ , \new_[11414]_ ,
    \new_[11415]_ , \new_[11416]_ , \new_[11417]_ , \new_[11418]_ ,
    \new_[11419]_ , \new_[11420]_ , \new_[11421]_ , \new_[11422]_ ,
    \new_[11423]_ , \new_[11424]_ , \new_[11425]_ , \new_[11426]_ ,
    \new_[11427]_ , \new_[11428]_ , \new_[11429]_ , \new_[11430]_ ,
    \new_[11431]_ , \new_[11432]_ , \new_[11433]_ , \new_[11434]_ ,
    \new_[11435]_ , \new_[11436]_ , \new_[11437]_ , \new_[11438]_ ,
    \new_[11439]_ , \new_[11440]_ , \new_[11441]_ , \new_[11442]_ ,
    \new_[11443]_ , \new_[11444]_ , \new_[11445]_ , \new_[11446]_ ,
    \new_[11447]_ , \new_[11448]_ , \new_[11449]_ , \new_[11450]_ ,
    \new_[11451]_ , \new_[11452]_ , \new_[11453]_ , \new_[11454]_ ,
    \new_[11455]_ , \new_[11456]_ , \new_[11457]_ , \new_[11458]_ ,
    \new_[11459]_ , \new_[11460]_ , \new_[11461]_ , \new_[11462]_ ,
    \new_[11463]_ , \new_[11464]_ , \new_[11465]_ , \new_[11466]_ ,
    \new_[11467]_ , \new_[11468]_ , \new_[11469]_ , \new_[11470]_ ,
    \new_[11471]_ , \new_[11472]_ , \new_[11473]_ , \new_[11474]_ ,
    \new_[11475]_ , \new_[11476]_ , \new_[11477]_ , \new_[11478]_ ,
    \new_[11479]_ , \new_[11480]_ , \new_[11481]_ , \new_[11482]_ ,
    \new_[11483]_ , \new_[11484]_ , \new_[11485]_ , \new_[11486]_ ,
    \new_[11487]_ , \new_[11488]_ , \new_[11489]_ , \new_[11490]_ ,
    \new_[11491]_ , \new_[11492]_ , \new_[11493]_ , \new_[11494]_ ,
    \new_[11495]_ , \new_[11496]_ , \new_[11497]_ , \new_[11498]_ ,
    \new_[11499]_ , \new_[11500]_ , \new_[11501]_ , \new_[11502]_ ,
    \new_[11503]_ , \new_[11504]_ , \new_[11505]_ , \new_[11506]_ ,
    \new_[11507]_ , \new_[11508]_ , \new_[11509]_ , \new_[11510]_ ,
    \new_[11511]_ , \new_[11512]_ , \new_[11513]_ , \new_[11514]_ ,
    \new_[11515]_ , \new_[11516]_ , \new_[11517]_ , \new_[11518]_ ,
    \new_[11519]_ , \new_[11520]_ , \new_[11521]_ , \new_[11522]_ ,
    \new_[11523]_ , \new_[11524]_ , \new_[11525]_ , \new_[11526]_ ,
    \new_[11527]_ , \new_[11528]_ , \new_[11529]_ , \new_[11530]_ ,
    \new_[11531]_ , \new_[11532]_ , \new_[11533]_ , \new_[11534]_ ,
    \new_[11535]_ , \new_[11536]_ , \new_[11537]_ , \new_[11538]_ ,
    \new_[11539]_ , \new_[11540]_ , \new_[11541]_ , \new_[11542]_ ,
    \new_[11543]_ , \new_[11544]_ , \new_[11545]_ , \new_[11546]_ ,
    \new_[11547]_ , \new_[11548]_ , \new_[11549]_ , \new_[11550]_ ,
    \new_[11551]_ , \new_[11552]_ , \new_[11553]_ , \new_[11554]_ ,
    \new_[11555]_ , \new_[11556]_ , \new_[11557]_ , \new_[11558]_ ,
    \new_[11559]_ , \new_[11560]_ , \new_[11561]_ , \new_[11562]_ ,
    \new_[11563]_ , \new_[11564]_ , \new_[11565]_ , \new_[11566]_ ,
    \new_[11567]_ , \new_[11568]_ , \new_[11569]_ , \new_[11570]_ ,
    \new_[11571]_ , \new_[11572]_ , \new_[11573]_ , \new_[11574]_ ,
    \new_[11575]_ , \new_[11576]_ , \new_[11577]_ , \new_[11578]_ ,
    \new_[11579]_ , \new_[11580]_ , \new_[11581]_ , \new_[11582]_ ,
    \new_[11583]_ , \new_[11584]_ , \new_[11585]_ , \new_[11586]_ ,
    \new_[11587]_ , \new_[11588]_ , \new_[11589]_ , \new_[11590]_ ,
    \new_[11591]_ , \new_[11592]_ , \new_[11593]_ , \new_[11594]_ ,
    \new_[11595]_ , \new_[11596]_ , \new_[11597]_ , \new_[11598]_ ,
    \new_[11599]_ , \new_[11600]_ , \new_[11601]_ , \new_[11602]_ ,
    \new_[11603]_ , \new_[11604]_ , \new_[11605]_ , \new_[11606]_ ,
    \new_[11607]_ , \new_[11608]_ , \new_[11609]_ , \new_[11610]_ ,
    \new_[11611]_ , \new_[11612]_ , \new_[11613]_ , \new_[11614]_ ,
    \new_[11616]_ , \new_[11617]_ , \new_[11622]_ , \new_[11624]_ ,
    \new_[11630]_ , \new_[11633]_ , \new_[11634]_ , \new_[11636]_ ,
    \new_[11637]_ , \new_[11638]_ , \new_[11640]_ , \new_[11641]_ ,
    \new_[11644]_ , \new_[11645]_ , \new_[11646]_ , \new_[11647]_ ,
    \new_[11648]_ , \new_[11649]_ , \new_[11650]_ , \new_[11651]_ ,
    \new_[11652]_ , \new_[11653]_ , \new_[11654]_ , \new_[11655]_ ,
    \new_[11656]_ , \new_[11657]_ , \new_[11658]_ , \new_[11659]_ ,
    \new_[11660]_ , \new_[11661]_ , \new_[11662]_ , \new_[11663]_ ,
    \new_[11664]_ , \new_[11665]_ , \new_[11666]_ , \new_[11667]_ ,
    \new_[11668]_ , \new_[11669]_ , \new_[11670]_ , \new_[11671]_ ,
    \new_[11672]_ , \new_[11673]_ , \new_[11674]_ , \new_[11675]_ ,
    \new_[11676]_ , \new_[11677]_ , \new_[11678]_ , \new_[11679]_ ,
    \new_[11680]_ , \new_[11681]_ , \new_[11682]_ , \new_[11683]_ ,
    \new_[11684]_ , \new_[11685]_ , \new_[11686]_ , \new_[11687]_ ,
    \new_[11688]_ , \new_[11689]_ , \new_[11690]_ , \new_[11691]_ ,
    \new_[11692]_ , \new_[11693]_ , \new_[11694]_ , \new_[11695]_ ,
    \new_[11696]_ , \new_[11697]_ , \new_[11698]_ , \new_[11699]_ ,
    \new_[11700]_ , \new_[11701]_ , \new_[11702]_ , \new_[11703]_ ,
    \new_[11704]_ , \new_[11705]_ , \new_[11706]_ , \new_[11707]_ ,
    \new_[11708]_ , \new_[11709]_ , \new_[11710]_ , \new_[11711]_ ,
    \new_[11712]_ , \new_[11713]_ , \new_[11714]_ , \new_[11715]_ ,
    \new_[11716]_ , \new_[11717]_ , \new_[11718]_ , \new_[11719]_ ,
    \new_[11720]_ , \new_[11721]_ , \new_[11722]_ , \new_[11723]_ ,
    \new_[11724]_ , \new_[11725]_ , \new_[11726]_ , \new_[11727]_ ,
    \new_[11728]_ , \new_[11729]_ , \new_[11730]_ , \new_[11731]_ ,
    \new_[11732]_ , \new_[11733]_ , \new_[11734]_ , \new_[11735]_ ,
    \new_[11736]_ , \new_[11737]_ , \new_[11738]_ , \new_[11739]_ ,
    \new_[11740]_ , \new_[11741]_ , \new_[11742]_ , \new_[11743]_ ,
    \new_[11744]_ , \new_[11745]_ , \new_[11746]_ , \new_[11747]_ ,
    \new_[11748]_ , \new_[11749]_ , \new_[11750]_ , \new_[11751]_ ,
    \new_[11752]_ , \new_[11753]_ , \new_[11754]_ , \new_[11755]_ ,
    \new_[11756]_ , \new_[11757]_ , \new_[11758]_ , \new_[11759]_ ,
    \new_[11760]_ , \new_[11761]_ , \new_[11762]_ , \new_[11763]_ ,
    \new_[11764]_ , \new_[11765]_ , \new_[11766]_ , \new_[11767]_ ,
    \new_[11768]_ , \new_[11769]_ , \new_[11770]_ , \new_[11771]_ ,
    \new_[11772]_ , \new_[11773]_ , \new_[11774]_ , \new_[11775]_ ,
    \new_[11776]_ , \new_[11777]_ , \new_[11778]_ , \new_[11779]_ ,
    \new_[11780]_ , \new_[11781]_ , \new_[11782]_ , \new_[11783]_ ,
    \new_[11784]_ , \new_[11785]_ , \new_[11786]_ , \new_[11787]_ ,
    \new_[11788]_ , \new_[11789]_ , \new_[11790]_ , \new_[11791]_ ,
    \new_[11792]_ , \new_[11793]_ , \new_[11794]_ , \new_[11795]_ ,
    \new_[11796]_ , \new_[11797]_ , \new_[11798]_ , \new_[11799]_ ,
    \new_[11800]_ , \new_[11801]_ , \new_[11804]_ , \new_[11805]_ ,
    \new_[11806]_ , \new_[11807]_ , \new_[11808]_ , \new_[11809]_ ,
    \new_[11810]_ , \new_[11811]_ , \new_[11812]_ , \new_[11813]_ ,
    \new_[11814]_ , \new_[11815]_ , \new_[11816]_ , \new_[11817]_ ,
    \new_[11818]_ , \new_[11819]_ , \new_[11820]_ , \new_[11821]_ ,
    \new_[11822]_ , \new_[11823]_ , \new_[11824]_ , \new_[11825]_ ,
    \new_[11826]_ , \new_[11827]_ , \new_[11828]_ , \new_[11829]_ ,
    \new_[11830]_ , \new_[11831]_ , \new_[11832]_ , \new_[11833]_ ,
    \new_[11834]_ , \new_[11835]_ , \new_[11836]_ , \new_[11837]_ ,
    \new_[11838]_ , \new_[11839]_ , \new_[11840]_ , \new_[11841]_ ,
    \new_[11842]_ , \new_[11843]_ , \new_[11844]_ , \new_[11845]_ ,
    \new_[11846]_ , \new_[11847]_ , \new_[11848]_ , \new_[11849]_ ,
    \new_[11850]_ , \new_[11851]_ , \new_[11852]_ , \new_[11853]_ ,
    \new_[11854]_ , \new_[11855]_ , \new_[11856]_ , \new_[11857]_ ,
    \new_[11858]_ , \new_[11859]_ , \new_[11860]_ , \new_[11861]_ ,
    \new_[11862]_ , \new_[11864]_ , \new_[11865]_ , \new_[11867]_ ,
    \new_[11868]_ , \new_[11869]_ , \new_[11870]_ , \new_[11871]_ ,
    \new_[11872]_ , \new_[11873]_ , \new_[11874]_ , \new_[11875]_ ,
    \new_[11876]_ , \new_[11877]_ , \new_[11878]_ , \new_[11879]_ ,
    \new_[11880]_ , \new_[11881]_ , \new_[11882]_ , \new_[11883]_ ,
    \new_[11884]_ , \new_[11885]_ , \new_[11886]_ , \new_[11887]_ ,
    \new_[11888]_ , \new_[11889]_ , \new_[11890]_ , \new_[11891]_ ,
    \new_[11892]_ , \new_[11893]_ , \new_[11894]_ , \new_[11896]_ ,
    \new_[11899]_ , \new_[11900]_ , \new_[11901]_ , \new_[11902]_ ,
    \new_[11903]_ , \new_[11904]_ , \new_[11905]_ , \new_[11906]_ ,
    \new_[11908]_ , \new_[11909]_ , \new_[11910]_ , \new_[11911]_ ,
    \new_[11912]_ , \new_[11913]_ , \new_[11914]_ , \new_[11916]_ ,
    \new_[11917]_ , \new_[11918]_ , \new_[11923]_ , \new_[11927]_ ,
    \new_[11931]_ , \new_[11934]_ , \new_[11936]_ , \new_[11938]_ ,
    \new_[11939]_ , \new_[11940]_ , \new_[11944]_ , \new_[11945]_ ,
    \new_[11946]_ , \new_[11947]_ , \new_[11948]_ , \new_[11949]_ ,
    \new_[11953]_ , \new_[11954]_ , \new_[11955]_ , \new_[11956]_ ,
    \new_[11957]_ , \new_[11958]_ , \new_[11959]_ , \new_[11960]_ ,
    \new_[11961]_ , \new_[11962]_ , \new_[11963]_ , \new_[11964]_ ,
    \new_[11965]_ , \new_[11966]_ , \new_[11967]_ , \new_[11968]_ ,
    \new_[11969]_ , \new_[11970]_ , \new_[11971]_ , \new_[11972]_ ,
    \new_[11973]_ , \new_[11974]_ , \new_[11975]_ , \new_[11976]_ ,
    \new_[11977]_ , \new_[11978]_ , \new_[11979]_ , \new_[11980]_ ,
    \new_[11981]_ , \new_[11982]_ , \new_[11983]_ , \new_[11984]_ ,
    \new_[11985]_ , \new_[11986]_ , \new_[11987]_ , \new_[11988]_ ,
    \new_[11989]_ , \new_[11990]_ , \new_[11991]_ , \new_[11992]_ ,
    \new_[11993]_ , \new_[11994]_ , \new_[11995]_ , \new_[11996]_ ,
    \new_[11997]_ , \new_[11998]_ , \new_[11999]_ , \new_[12000]_ ,
    \new_[12001]_ , \new_[12002]_ , \new_[12003]_ , \new_[12004]_ ,
    \new_[12005]_ , \new_[12006]_ , \new_[12007]_ , \new_[12008]_ ,
    \new_[12009]_ , \new_[12010]_ , \new_[12011]_ , \new_[12012]_ ,
    \new_[12013]_ , \new_[12014]_ , \new_[12015]_ , \new_[12016]_ ,
    \new_[12017]_ , \new_[12018]_ , \new_[12019]_ , \new_[12020]_ ,
    \new_[12021]_ , \new_[12022]_ , \new_[12023]_ , \new_[12024]_ ,
    \new_[12025]_ , \new_[12026]_ , \new_[12027]_ , \new_[12028]_ ,
    \new_[12029]_ , \new_[12030]_ , \new_[12031]_ , \new_[12032]_ ,
    \new_[12033]_ , \new_[12034]_ , \new_[12035]_ , \new_[12036]_ ,
    \new_[12037]_ , \new_[12038]_ , \new_[12039]_ , \new_[12040]_ ,
    \new_[12041]_ , \new_[12042]_ , \new_[12043]_ , \new_[12044]_ ,
    \new_[12045]_ , \new_[12046]_ , \new_[12047]_ , \new_[12048]_ ,
    \new_[12049]_ , \new_[12050]_ , \new_[12051]_ , \new_[12052]_ ,
    \new_[12053]_ , \new_[12054]_ , \new_[12055]_ , \new_[12056]_ ,
    \new_[12057]_ , \new_[12058]_ , \new_[12059]_ , \new_[12060]_ ,
    \new_[12061]_ , \new_[12062]_ , \new_[12063]_ , \new_[12064]_ ,
    \new_[12065]_ , \new_[12066]_ , \new_[12067]_ , \new_[12068]_ ,
    \new_[12069]_ , \new_[12070]_ , \new_[12071]_ , \new_[12072]_ ,
    \new_[12073]_ , \new_[12074]_ , \new_[12075]_ , \new_[12076]_ ,
    \new_[12077]_ , \new_[12078]_ , \new_[12079]_ , \new_[12080]_ ,
    \new_[12081]_ , \new_[12082]_ , \new_[12083]_ , \new_[12084]_ ,
    \new_[12085]_ , \new_[12086]_ , \new_[12087]_ , \new_[12088]_ ,
    \new_[12089]_ , \new_[12090]_ , \new_[12091]_ , \new_[12092]_ ,
    \new_[12093]_ , \new_[12094]_ , \new_[12095]_ , \new_[12096]_ ,
    \new_[12097]_ , \new_[12098]_ , \new_[12099]_ , \new_[12100]_ ,
    \new_[12101]_ , \new_[12102]_ , \new_[12103]_ , \new_[12104]_ ,
    \new_[12105]_ , \new_[12106]_ , \new_[12107]_ , \new_[12108]_ ,
    \new_[12109]_ , \new_[12110]_ , \new_[12111]_ , \new_[12112]_ ,
    \new_[12113]_ , \new_[12114]_ , \new_[12115]_ , \new_[12116]_ ,
    \new_[12117]_ , \new_[12118]_ , \new_[12119]_ , \new_[12120]_ ,
    \new_[12121]_ , \new_[12122]_ , \new_[12123]_ , \new_[12124]_ ,
    \new_[12125]_ , \new_[12126]_ , \new_[12127]_ , \new_[12128]_ ,
    \new_[12129]_ , \new_[12130]_ , \new_[12131]_ , \new_[12132]_ ,
    \new_[12133]_ , \new_[12134]_ , \new_[12135]_ , \new_[12136]_ ,
    \new_[12137]_ , \new_[12138]_ , \new_[12139]_ , \new_[12140]_ ,
    \new_[12141]_ , \new_[12142]_ , \new_[12143]_ , \new_[12144]_ ,
    \new_[12145]_ , \new_[12146]_ , \new_[12147]_ , \new_[12148]_ ,
    \new_[12149]_ , \new_[12150]_ , \new_[12151]_ , \new_[12152]_ ,
    \new_[12153]_ , \new_[12154]_ , \new_[12155]_ , \new_[12156]_ ,
    \new_[12157]_ , \new_[12158]_ , \new_[12159]_ , \new_[12160]_ ,
    \new_[12161]_ , \new_[12162]_ , \new_[12163]_ , \new_[12164]_ ,
    \new_[12165]_ , \new_[12166]_ , \new_[12167]_ , \new_[12168]_ ,
    \new_[12169]_ , \new_[12170]_ , \new_[12171]_ , \new_[12172]_ ,
    \new_[12173]_ , \new_[12174]_ , \new_[12175]_ , \new_[12176]_ ,
    \new_[12177]_ , \new_[12178]_ , \new_[12179]_ , \new_[12180]_ ,
    \new_[12181]_ , \new_[12182]_ , \new_[12183]_ , \new_[12184]_ ,
    \new_[12185]_ , \new_[12186]_ , \new_[12189]_ , \new_[12190]_ ,
    \new_[12192]_ , \new_[12194]_ , \new_[12195]_ , \new_[12196]_ ,
    \new_[12197]_ , \new_[12198]_ , \new_[12199]_ , \new_[12201]_ ,
    \new_[12202]_ , \new_[12205]_ , \new_[12212]_ , \new_[12223]_ ,
    \new_[12234]_ , \new_[12235]_ , \new_[12236]_ , \new_[12238]_ ,
    \new_[12241]_ , \new_[12242]_ , \new_[12243]_ , \new_[12244]_ ,
    \new_[12245]_ , \new_[12246]_ , \new_[12247]_ , \new_[12248]_ ,
    \new_[12249]_ , \new_[12250]_ , \new_[12251]_ , \new_[12252]_ ,
    \new_[12253]_ , \new_[12254]_ , \new_[12255]_ , \new_[12256]_ ,
    \new_[12257]_ , \new_[12258]_ , \new_[12259]_ , \new_[12260]_ ,
    \new_[12261]_ , \new_[12266]_ , \new_[12267]_ , \new_[12268]_ ,
    \new_[12269]_ , \new_[12270]_ , \new_[12271]_ , \new_[12272]_ ,
    \new_[12273]_ , \new_[12274]_ , \new_[12277]_ , \new_[12278]_ ,
    \new_[12281]_ , \new_[12282]_ , \new_[12286]_ , \new_[12287]_ ,
    \new_[12289]_ , \new_[12290]_ , \new_[12291]_ , \new_[12292]_ ,
    \new_[12293]_ , \new_[12294]_ , \new_[12295]_ , \new_[12296]_ ,
    \new_[12297]_ , \new_[12298]_ , \new_[12299]_ , \new_[12300]_ ,
    \new_[12301]_ , \new_[12302]_ , \new_[12303]_ , \new_[12304]_ ,
    \new_[12305]_ , \new_[12306]_ , \new_[12307]_ , \new_[12308]_ ,
    \new_[12309]_ , \new_[12310]_ , \new_[12311]_ , \new_[12312]_ ,
    \new_[12313]_ , \new_[12314]_ , \new_[12315]_ , \new_[12316]_ ,
    \new_[12317]_ , \new_[12318]_ , \new_[12319]_ , \new_[12320]_ ,
    \new_[12321]_ , \new_[12322]_ , \new_[12323]_ , \new_[12324]_ ,
    \new_[12325]_ , \new_[12326]_ , \new_[12327]_ , \new_[12328]_ ,
    \new_[12329]_ , \new_[12330]_ , \new_[12331]_ , \new_[12332]_ ,
    \new_[12333]_ , \new_[12334]_ , \new_[12335]_ , \new_[12336]_ ,
    \new_[12337]_ , \new_[12338]_ , \new_[12339]_ , \new_[12340]_ ,
    \new_[12341]_ , \new_[12342]_ , \new_[12343]_ , \new_[12344]_ ,
    \new_[12345]_ , \new_[12346]_ , \new_[12347]_ , \new_[12348]_ ,
    \new_[12349]_ , \new_[12350]_ , \new_[12351]_ , \new_[12352]_ ,
    \new_[12353]_ , \new_[12354]_ , \new_[12355]_ , \new_[12356]_ ,
    \new_[12357]_ , \new_[12358]_ , \new_[12359]_ , \new_[12360]_ ,
    \new_[12361]_ , \new_[12362]_ , \new_[12363]_ , \new_[12364]_ ,
    \new_[12365]_ , \new_[12366]_ , \new_[12367]_ , \new_[12368]_ ,
    \new_[12369]_ , \new_[12370]_ , \new_[12371]_ , \new_[12372]_ ,
    \new_[12373]_ , \new_[12374]_ , \new_[12375]_ , \new_[12376]_ ,
    \new_[12377]_ , \new_[12378]_ , \new_[12379]_ , \new_[12380]_ ,
    \new_[12381]_ , \new_[12382]_ , \new_[12383]_ , \new_[12384]_ ,
    \new_[12385]_ , \new_[12386]_ , \new_[12387]_ , \new_[12388]_ ,
    \new_[12389]_ , \new_[12390]_ , \new_[12391]_ , \new_[12392]_ ,
    \new_[12393]_ , \new_[12394]_ , \new_[12395]_ , \new_[12396]_ ,
    \new_[12397]_ , \new_[12398]_ , \new_[12399]_ , \new_[12400]_ ,
    \new_[12401]_ , \new_[12402]_ , \new_[12403]_ , \new_[12404]_ ,
    \new_[12405]_ , \new_[12406]_ , \new_[12407]_ , \new_[12408]_ ,
    \new_[12409]_ , \new_[12410]_ , \new_[12411]_ , \new_[12412]_ ,
    \new_[12413]_ , \new_[12414]_ , \new_[12415]_ , \new_[12416]_ ,
    \new_[12417]_ , \new_[12418]_ , \new_[12419]_ , \new_[12420]_ ,
    \new_[12421]_ , \new_[12422]_ , \new_[12423]_ , \new_[12424]_ ,
    \new_[12425]_ , \new_[12426]_ , \new_[12427]_ , \new_[12428]_ ,
    \new_[12429]_ , \new_[12430]_ , \new_[12431]_ , \new_[12432]_ ,
    \new_[12433]_ , \new_[12434]_ , \new_[12435]_ , \new_[12436]_ ,
    \new_[12437]_ , \new_[12438]_ , \new_[12439]_ , \new_[12440]_ ,
    \new_[12441]_ , \new_[12442]_ , \new_[12443]_ , \new_[12444]_ ,
    \new_[12445]_ , \new_[12446]_ , \new_[12447]_ , \new_[12448]_ ,
    \new_[12449]_ , \new_[12450]_ , \new_[12451]_ , \new_[12452]_ ,
    \new_[12453]_ , \new_[12454]_ , \new_[12455]_ , \new_[12456]_ ,
    \new_[12457]_ , \new_[12458]_ , \new_[12459]_ , \new_[12460]_ ,
    \new_[12461]_ , \new_[12462]_ , \new_[12463]_ , \new_[12464]_ ,
    \new_[12465]_ , \new_[12466]_ , \new_[12467]_ , \new_[12468]_ ,
    \new_[12469]_ , \new_[12470]_ , \new_[12471]_ , \new_[12472]_ ,
    \new_[12473]_ , \new_[12474]_ , \new_[12475]_ , \new_[12476]_ ,
    \new_[12477]_ , \new_[12478]_ , \new_[12479]_ , \new_[12481]_ ,
    \new_[12482]_ , \new_[12483]_ , \new_[12484]_ , \new_[12485]_ ,
    \new_[12486]_ , \new_[12487]_ , \new_[12488]_ , \new_[12489]_ ,
    \new_[12490]_ , \new_[12491]_ , \new_[12492]_ , \new_[12493]_ ,
    \new_[12494]_ , \new_[12495]_ , \new_[12496]_ , \new_[12497]_ ,
    \new_[12498]_ , \new_[12499]_ , \new_[12500]_ , \new_[12501]_ ,
    \new_[12502]_ , \new_[12503]_ , \new_[12504]_ , \new_[12505]_ ,
    \new_[12506]_ , \new_[12507]_ , \new_[12508]_ , \new_[12509]_ ,
    \new_[12510]_ , \new_[12511]_ , \new_[12512]_ , \new_[12513]_ ,
    \new_[12514]_ , \new_[12515]_ , \new_[12516]_ , \new_[12517]_ ,
    \new_[12518]_ , \new_[12519]_ , \new_[12520]_ , \new_[12521]_ ,
    \new_[12522]_ , \new_[12523]_ , \new_[12524]_ , \new_[12525]_ ,
    \new_[12526]_ , \new_[12527]_ , \new_[12528]_ , \new_[12529]_ ,
    \new_[12530]_ , \new_[12531]_ , \new_[12532]_ , \new_[12533]_ ,
    \new_[12534]_ , \new_[12535]_ , \new_[12536]_ , \new_[12537]_ ,
    \new_[12538]_ , \new_[12542]_ , \new_[12543]_ , \new_[12545]_ ,
    \new_[12547]_ , \new_[12548]_ , \new_[12549]_ , \new_[12565]_ ,
    \new_[12566]_ , \new_[12567]_ , \new_[12568]_ , \new_[12569]_ ,
    \new_[12570]_ , \new_[12571]_ , \new_[12572]_ , \new_[12573]_ ,
    \new_[12574]_ , \new_[12575]_ , \new_[12576]_ , \new_[13117]_ ,
    \new_[13118]_ , \new_[13119]_ , \new_[13120]_ , \new_[13121]_ ,
    \new_[13122]_ , \new_[13123]_ , \new_[13125]_ , \new_[13126]_ ,
    \new_[13127]_ , \new_[13128]_ , \new_[13129]_ , \new_[13130]_ ,
    \new_[13131]_ , \new_[13132]_ , \new_[13134]_ , \new_[13135]_ ,
    \new_[13136]_ , \new_[13138]_ , \new_[13141]_ , \new_[13142]_ ,
    \new_[13144]_ , \new_[13146]_ , \new_[13147]_ , \new_[13149]_ ,
    \new_[13150]_ , \new_[13151]_ , \new_[13152]_ , \new_[13153]_ ,
    \new_[13154]_ , \new_[13155]_ , \new_[13157]_ , \new_[13158]_ ,
    \new_[13160]_ , \new_[13208]_ , \new_[13210]_ , \new_[13212]_ ,
    \new_[13213]_ , \new_[13214]_ , \new_[13215]_ , \new_[13216]_ ,
    \new_[13217]_ , \new_[13218]_ , \new_[13219]_ , \new_[13221]_ ,
    \new_[13222]_ , \new_[13223]_ , \new_[13295]_ , \new_[13296]_ ,
    \new_[13297]_ , \new_[13298]_ , \new_[13299]_ , \new_[13434]_ ,
    \new_[13435]_ , \new_[13436]_ , \new_[13437]_ , \new_[13490]_ ,
    \new_[13571]_ , \new_[13572]_ , \new_[13577]_ , \new_[13582]_ ,
    \new_[13583]_ , \new_[13584]_ , \new_[13585]_ , \new_[13586]_ ,
    \new_[13587]_ , \new_[13588]_ , \new_[13589]_ , \new_[13590]_ ,
    \new_[13591]_ , \new_[13592]_ , \new_[13593]_ , \new_[13594]_ ,
    \new_[13595]_ , \new_[13596]_ , \new_[13597]_ , \new_[13598]_ ,
    \new_[13599]_ , \new_[13600]_ , \new_[13601]_ , \new_[13603]_ ,
    \new_[13606]_ , \new_[13607]_ , \new_[13608]_ , \new_[13609]_ ,
    \new_[13610]_ , \new_[13611]_ , \new_[13612]_ , \new_[13613]_ ,
    \new_[13614]_ , \new_[13615]_ , \new_[13616]_ , \new_[13617]_ ,
    \new_[13618]_ , \new_[13620]_ , \new_[13621]_ , \new_[13622]_ ,
    \new_[13623]_ , \new_[13624]_ , \new_[13625]_ , \new_[13626]_ ,
    \new_[13627]_ , \new_[13628]_ , \new_[13629]_ , \new_[13630]_ ,
    \new_[13633]_ , \new_[13635]_ , \new_[13640]_ , \new_[13643]_ ,
    \new_[13644]_ , \new_[13645]_ , \new_[13646]_ , \new_[13647]_ ,
    \new_[13648]_ , \new_[13649]_ , \new_[13672]_ , \new_[13674]_ ,
    \new_[13676]_ , \new_[13677]_ , \new_[13678]_ , \new_[13679]_ ,
    \new_[13680]_ , \new_[13681]_ , \new_[13682]_ , \new_[13683]_ ,
    \new_[13684]_ , \new_[13685]_ , \new_[13686]_ , \new_[13687]_ ,
    \new_[13688]_ , \new_[13689]_ , \new_[13690]_ , \new_[13692]_ ,
    \new_[13693]_ , \new_[13694]_ , \new_[13695]_ , \new_[13696]_ ,
    \new_[13697]_ , \new_[13698]_ , \new_[13699]_ , \new_[13700]_ ,
    \new_[13701]_ , \new_[13702]_ , \new_[13703]_ , \new_[13704]_ ,
    \new_[13705]_ , \new_[13706]_ , \new_[13707]_ , \new_[13709]_ ,
    \new_[13710]_ , \new_[13711]_ , \new_[13714]_ , \new_[13715]_ ,
    \new_[13716]_ , \new_[13717]_ , \new_[13718]_ , \new_[13719]_ ,
    \new_[13720]_ , \new_[13721]_ , \new_[13722]_ , \new_[13723]_ ,
    \new_[13724]_ , \new_[13725]_ , \new_[13726]_ , \new_[13727]_ ,
    \new_[13728]_ , \new_[13729]_ , \new_[13730]_ , \new_[13731]_ ,
    \new_[13732]_ , \new_[13733]_ , \new_[13734]_ , \new_[13735]_ ,
    \new_[13736]_ , \new_[13737]_ , \new_[13738]_ , \new_[13739]_ ,
    \new_[13740]_ , \new_[13741]_ , \new_[13742]_ , \new_[13743]_ ,
    \new_[13744]_ , \new_[13745]_ , \new_[13746]_ , \new_[13747]_ ,
    \new_[13748]_ , \new_[13749]_ , \new_[13750]_ , \new_[13751]_ ,
    \new_[13752]_ , \new_[13753]_ , \new_[13754]_ , \new_[13755]_ ,
    \new_[13756]_ , \new_[13757]_ , \new_[13758]_ , \new_[13759]_ ,
    \new_[13761]_ , \new_[13762]_ , \new_[13763]_ , \new_[13764]_ ,
    \new_[13765]_ , \new_[13766]_ , \new_[13767]_ , \new_[13768]_ ,
    \new_[13769]_ , \new_[13770]_ , \new_[13771]_ , \new_[13772]_ ,
    \new_[13773]_ , \new_[13774]_ , \new_[13775]_ , \new_[13776]_ ,
    \new_[13777]_ , \new_[13778]_ , \new_[13779]_ , \new_[13780]_ ,
    \new_[13781]_ , \new_[13782]_ , \new_[13783]_ , \new_[13784]_ ,
    \new_[13785]_ , \new_[13787]_ , \new_[13788]_ , \new_[13789]_ ,
    \new_[13790]_ , \new_[13791]_ , \new_[13792]_ , \new_[13793]_ ,
    \new_[13794]_ , \new_[13795]_ , \new_[13796]_ , \new_[13797]_ ,
    \new_[13798]_ , \new_[13799]_ , \new_[13800]_ , \new_[13801]_ ,
    \new_[13802]_ , \new_[13803]_ , \new_[13804]_ , \new_[13807]_ ,
    \new_[13808]_ , \new_[13809]_ , \new_[13810]_ , \new_[13811]_ ,
    \new_[13812]_ , \new_[13813]_ , \new_[13814]_ , \new_[13815]_ ,
    \new_[13816]_ , \new_[13817]_ , \new_[13818]_ , \new_[13819]_ ,
    \new_[13820]_ , \new_[13821]_ , \new_[13822]_ , \new_[13823]_ ,
    \new_[13826]_ , \new_[13827]_ , \new_[13828]_ , \new_[13829]_ ,
    \new_[13830]_ , \new_[13832]_ , \new_[13833]_ , \new_[13834]_ ,
    \new_[13835]_ , \new_[13836]_ , \new_[13837]_ , \new_[13838]_ ,
    \new_[13839]_ , \new_[13840]_ , \new_[13841]_ , \new_[13842]_ ,
    \new_[13843]_ , \new_[13844]_ , \new_[13845]_ , \new_[13846]_ ,
    \new_[13847]_ , \new_[13848]_ , \new_[13849]_ , \new_[13850]_ ,
    \new_[13851]_ , \new_[13852]_ , \new_[13853]_ , \new_[13854]_ ,
    \new_[13858]_ , \new_[13860]_ , \new_[13862]_ , \new_[13863]_ ,
    \new_[13864]_ , \new_[13869]_ , \new_[13870]_ , \new_[13871]_ ,
    \new_[13872]_ , \new_[13875]_ , \new_[13876]_ , \new_[13877]_ ,
    \new_[13878]_ , \new_[13879]_ , \new_[13880]_ , \new_[13885]_ ,
    \new_[13886]_ , \new_[13887]_ , \new_[13888]_ , \new_[13889]_ ,
    \new_[13890]_ , \new_[13891]_ , \new_[13892]_ , \new_[13893]_ ,
    \new_[13894]_ , \new_[13895]_ , \new_[13896]_ , \new_[13897]_ ,
    \new_[13898]_ , \new_[13899]_ , \new_[13900]_ , \new_[13901]_ ,
    \new_[13902]_ , \new_[13903]_ , \new_[13904]_ , \new_[13905]_ ,
    \new_[13906]_ , \new_[13907]_ , \new_[13908]_ , \new_[13909]_ ,
    \new_[13910]_ , \new_[13911]_ , \new_[13912]_ , \new_[13913]_ ,
    \new_[13915]_ , \new_[13918]_ , \new_[13919]_ , \new_[13920]_ ,
    \new_[13921]_ , \new_[13922]_ , \new_[13923]_ , \new_[13924]_ ,
    \new_[13925]_ , \new_[13926]_ , \new_[13927]_ , \new_[13928]_ ,
    \new_[13929]_ , \new_[13930]_ , \new_[13931]_ , \new_[13932]_ ,
    \new_[13933]_ , \new_[13934]_ , \new_[13935]_ , \new_[13936]_ ,
    \new_[13937]_ , \new_[13938]_ , \new_[13939]_ , \new_[13940]_ ,
    \new_[13941]_ , \new_[13942]_ , \new_[13943]_ , \new_[13944]_ ,
    \new_[13945]_ , \new_[13946]_ , \new_[13947]_ , \new_[13948]_ ,
    \new_[13949]_ , \new_[13950]_ , \new_[13951]_ , \new_[13952]_ ,
    \new_[13953]_ , \new_[13954]_ , \new_[13955]_ , \new_[13956]_ ,
    \new_[13957]_ , \new_[13958]_ , \new_[13959]_ , \new_[13960]_ ,
    \new_[13961]_ , \new_[13962]_ , \new_[13963]_ , \new_[13964]_ ,
    \new_[13965]_ , \new_[13966]_ , \new_[13967]_ , \new_[13968]_ ,
    \new_[13969]_ , \new_[13970]_ , \new_[13971]_ , \new_[13972]_ ,
    \new_[13973]_ , \new_[13974]_ , \new_[13975]_ , \new_[13976]_ ,
    \new_[13977]_ , \new_[13978]_ , \new_[13979]_ , \new_[13980]_ ,
    \new_[13981]_ , \new_[13982]_ , \new_[13983]_ , \new_[13984]_ ,
    \new_[13985]_ , \new_[13986]_ , \new_[13987]_ , \new_[13988]_ ,
    \new_[13989]_ , \new_[13990]_ , \new_[13991]_ , \new_[13992]_ ,
    \new_[13993]_ , \new_[13994]_ , \new_[13995]_ , \new_[13996]_ ,
    \new_[13997]_ , \new_[13998]_ , \new_[13999]_ , \new_[14000]_ ,
    \new_[14001]_ , \new_[14002]_ , \new_[14003]_ , \new_[14004]_ ,
    \new_[14005]_ , \new_[14006]_ , \new_[14007]_ , \new_[14008]_ ,
    \new_[14009]_ , \new_[14010]_ , \new_[14011]_ , \new_[14012]_ ,
    \new_[14013]_ , \new_[14014]_ , \new_[14015]_ , \new_[14016]_ ,
    \new_[14017]_ , \new_[14018]_ , \new_[14019]_ , \new_[14020]_ ,
    \new_[14021]_ , \new_[14022]_ , \new_[14023]_ , \new_[14024]_ ,
    \new_[14025]_ , \new_[14026]_ , \new_[14027]_ , \new_[14028]_ ,
    \new_[14029]_ , \new_[14030]_ , \new_[14031]_ , \new_[14032]_ ,
    \new_[14033]_ , \new_[14034]_ , \new_[14035]_ , \new_[14036]_ ,
    \new_[14037]_ , \new_[14038]_ , \new_[14039]_ , \new_[14040]_ ,
    \new_[14041]_ , \new_[14042]_ , \new_[14043]_ , \new_[14044]_ ,
    \new_[14045]_ , \new_[14046]_ , \new_[14047]_ , \new_[14048]_ ,
    \new_[14049]_ , \new_[14050]_ , \new_[14051]_ , \new_[14052]_ ,
    \new_[14053]_ , \new_[14054]_ , \new_[14055]_ , \new_[14056]_ ,
    \new_[14057]_ , \new_[14058]_ , \new_[14059]_ , \new_[14060]_ ,
    \new_[14061]_ , \new_[14062]_ , \new_[14063]_ , \new_[14064]_ ,
    \new_[14065]_ , \new_[14066]_ , \new_[14067]_ , \new_[14068]_ ,
    \new_[14069]_ , \new_[14070]_ , \new_[14071]_ , \new_[14072]_ ,
    \new_[14073]_ , \new_[14074]_ , \new_[14075]_ , \new_[14076]_ ,
    \new_[14077]_ , \new_[14078]_ , \new_[14079]_ , \new_[14080]_ ,
    \new_[14081]_ , \new_[14082]_ , \new_[14083]_ , \new_[14084]_ ,
    \new_[14085]_ , \new_[14086]_ , \new_[14087]_ , \new_[14088]_ ,
    \new_[14089]_ , \new_[14090]_ , \new_[14091]_ , \new_[14092]_ ,
    \new_[14093]_ , \new_[14094]_ , \new_[14095]_ , \new_[14096]_ ,
    \new_[14097]_ , \new_[14098]_ , \new_[14099]_ , \new_[14100]_ ,
    \new_[14101]_ , \new_[14102]_ , \new_[14103]_ , \new_[14104]_ ,
    \new_[14105]_ , \new_[14106]_ , \new_[14107]_ , \new_[14108]_ ,
    \new_[14109]_ , \new_[14110]_ , \new_[14111]_ , \new_[14112]_ ,
    \new_[14113]_ , \new_[14114]_ , \new_[14115]_ , \new_[14116]_ ,
    \new_[14117]_ , \new_[14118]_ , \new_[14119]_ , \new_[14120]_ ,
    \new_[14121]_ , \new_[14122]_ , \new_[14123]_ , \new_[14124]_ ,
    \new_[14125]_ , \new_[14126]_ , \new_[14127]_ , \new_[14128]_ ,
    \new_[14129]_ , \new_[14130]_ , \new_[14131]_ , \new_[14132]_ ,
    \new_[14133]_ , \new_[14134]_ , \new_[14135]_ , \new_[14136]_ ,
    \new_[14137]_ , \new_[14138]_ , \new_[14139]_ , \new_[14140]_ ,
    \new_[14141]_ , \new_[14142]_ , \new_[14143]_ , \new_[14144]_ ,
    \new_[14145]_ , \new_[14146]_ , \new_[14147]_ , \new_[14148]_ ,
    \new_[14149]_ , \new_[14150]_ , \new_[14151]_ , \new_[14152]_ ,
    \new_[14153]_ , \new_[14154]_ , \new_[14155]_ , \new_[14156]_ ,
    \new_[14157]_ , \new_[14158]_ , \new_[14159]_ , \new_[14160]_ ,
    \new_[14161]_ , \new_[14162]_ , \new_[14163]_ , \new_[14164]_ ,
    \new_[14165]_ , \new_[14166]_ , \new_[14167]_ , \new_[14168]_ ,
    \new_[14169]_ , \new_[14170]_ , \new_[14171]_ , \new_[14172]_ ,
    \new_[14173]_ , \new_[14174]_ , \new_[14175]_ , \new_[14176]_ ,
    \new_[14177]_ , \new_[14178]_ , \new_[14179]_ , \new_[14180]_ ,
    \new_[14181]_ , \new_[14182]_ , \new_[14183]_ , \new_[14184]_ ,
    \new_[14185]_ , \new_[14186]_ , \new_[14187]_ , \new_[14188]_ ,
    \new_[14190]_ , \new_[14191]_ , \new_[14192]_ , \new_[14193]_ ,
    \new_[14194]_ , \new_[14195]_ , \new_[14196]_ , \new_[14197]_ ,
    \new_[14198]_ , \new_[14199]_ , \new_[14200]_ , \new_[14201]_ ,
    \new_[14202]_ , \new_[14203]_ , \new_[14204]_ , \new_[14205]_ ,
    \new_[14207]_ , \new_[14208]_ , \new_[14209]_ , \new_[14210]_ ,
    \new_[14211]_ , \new_[14212]_ , \new_[14213]_ , \new_[14214]_ ,
    \new_[14215]_ , \new_[14216]_ , \new_[14217]_ , \new_[14218]_ ,
    \new_[14219]_ , \new_[14220]_ , \new_[14221]_ , \new_[14222]_ ,
    \new_[14223]_ , \new_[14224]_ , \new_[14225]_ , \new_[14226]_ ,
    \new_[14227]_ , \new_[14228]_ , \new_[14229]_ , \new_[14230]_ ,
    \new_[14231]_ , \new_[14232]_ , \new_[14233]_ , \new_[14234]_ ,
    \new_[14235]_ , \new_[14236]_ , \new_[14237]_ , \new_[14238]_ ,
    \new_[14239]_ , \new_[14241]_ , \new_[14242]_ , \new_[14243]_ ,
    \new_[14244]_ , \new_[14245]_ , \new_[14246]_ , \new_[14247]_ ,
    \new_[14250]_ , \new_[14252]_ , \new_[14253]_ , \new_[14254]_ ,
    \new_[14256]_ , \new_[14258]_ , \new_[14259]_ , \new_[14260]_ ,
    \new_[14261]_ , \new_[14262]_ , \new_[14278]_ , \new_[14279]_ ,
    \new_[14280]_ , \new_[14281]_ , \new_[14282]_ , \new_[14283]_ ,
    \new_[14284]_ , \new_[14285]_ , \new_[14286]_ , \new_[14287]_ ,
    \new_[14288]_ , \new_[14289]_ , \new_[14290]_ , \new_[14291]_ ,
    \new_[14292]_ , \new_[14293]_ , \new_[14294]_ , \new_[14295]_ ,
    \new_[14296]_ , \new_[14297]_ , \new_[14298]_ , \new_[14299]_ ,
    \new_[14300]_ , \new_[14301]_ , \new_[14302]_ , \new_[14303]_ ,
    \new_[14304]_ , \new_[14305]_ , \new_[14306]_ , \new_[14307]_ ,
    \new_[14308]_ , \new_[14309]_ , \new_[14310]_ , \new_[14311]_ ,
    \new_[14312]_ , \new_[14313]_ , \new_[14314]_ , \new_[14315]_ ,
    \new_[14316]_ , \new_[14317]_ , \new_[14318]_ , \new_[14319]_ ,
    \new_[14320]_ , \new_[14321]_ , \new_[14322]_ , \new_[14323]_ ,
    \new_[14324]_ , \new_[14325]_ , \new_[14326]_ , \new_[14327]_ ,
    \new_[14328]_ , \new_[14329]_ , \new_[14330]_ , \new_[14331]_ ,
    \new_[14332]_ , \new_[14333]_ , \new_[14334]_ , \new_[14335]_ ,
    \new_[14336]_ , \new_[14337]_ , \new_[14338]_ , \new_[14339]_ ,
    \new_[14340]_ , \new_[14341]_ , \new_[14342]_ , \new_[14343]_ ,
    \new_[14344]_ , \new_[14345]_ , \new_[14346]_ , \new_[14347]_ ,
    \new_[14348]_ , \new_[14349]_ , \new_[14350]_ , \new_[14351]_ ,
    \new_[14352]_ , \new_[14353]_ , \new_[14354]_ , \new_[14355]_ ,
    \new_[14356]_ , \new_[14357]_ , \new_[14358]_ , \new_[14359]_ ,
    \new_[14360]_ , \new_[14361]_ , \new_[14362]_ , \new_[14363]_ ,
    \new_[14364]_ , \new_[14365]_ , \new_[14366]_ , \new_[14367]_ ,
    \new_[14368]_ , \new_[14369]_ , \new_[14370]_ , \new_[14371]_ ,
    \new_[14372]_ , \new_[14373]_ , \new_[14374]_ , \new_[14375]_ ,
    \new_[14376]_ , \new_[14377]_ , \new_[14378]_ , \new_[14379]_ ,
    \new_[14380]_ , \new_[14381]_ , \new_[14382]_ , \new_[14383]_ ,
    \new_[14384]_ , \new_[14385]_ , \new_[14386]_ , \new_[14387]_ ,
    \new_[14388]_ , \new_[14389]_ , \new_[14390]_ , \new_[14391]_ ,
    \new_[14392]_ , \new_[14393]_ , \new_[14394]_ , \new_[14395]_ ,
    \new_[14396]_ , \new_[14397]_ , \new_[14398]_ , \new_[14399]_ ,
    \new_[14400]_ , \new_[14401]_ , \new_[14402]_ , \new_[14403]_ ,
    \new_[14404]_ , \new_[14405]_ , \new_[14406]_ , \new_[14407]_ ,
    \new_[14408]_ , \new_[14409]_ , \new_[14410]_ , \new_[14411]_ ,
    \new_[14412]_ , \new_[14413]_ , \new_[14414]_ , \new_[14415]_ ,
    \new_[14416]_ , \new_[14417]_ , \new_[14418]_ , \new_[14419]_ ,
    \new_[14420]_ , \new_[14421]_ , \new_[14422]_ , \new_[14423]_ ,
    \new_[14424]_ , \new_[14425]_ , \new_[14426]_ , \new_[14427]_ ,
    \new_[14428]_ , \new_[14429]_ , \new_[14430]_ , \new_[14431]_ ,
    \new_[14432]_ , \new_[14433]_ , \new_[14434]_ , \new_[14435]_ ,
    \new_[14436]_ , \new_[14437]_ , \new_[14438]_ , \new_[14439]_ ,
    \new_[14440]_ , \new_[14441]_ , \new_[14442]_ , \new_[14443]_ ,
    \new_[14444]_ , \new_[14445]_ , \new_[14446]_ , \new_[14447]_ ,
    \new_[14448]_ , \new_[14449]_ , \new_[14450]_ , \new_[14451]_ ,
    \new_[14452]_ , \new_[14453]_ , \new_[14454]_ , \new_[14455]_ ,
    \new_[14456]_ , \new_[14457]_ , \new_[14458]_ , \new_[14459]_ ,
    \new_[14460]_ , \new_[14461]_ , \new_[14462]_ , \new_[14463]_ ,
    \new_[14464]_ , \new_[14465]_ , \new_[14466]_ , \new_[14467]_ ,
    \new_[14468]_ , \new_[14469]_ , \new_[14470]_ , \new_[14471]_ ,
    \new_[14472]_ , \new_[14473]_ , \new_[14474]_ , \new_[14475]_ ,
    \new_[14476]_ , \new_[14477]_ , \new_[14478]_ , \new_[14479]_ ,
    \new_[14480]_ , \new_[14481]_ , \new_[14482]_ , \new_[14483]_ ,
    \new_[14484]_ , \new_[14485]_ , \new_[14486]_ , \new_[14487]_ ,
    \new_[14488]_ , \new_[14489]_ , \new_[14490]_ , \new_[14491]_ ,
    \new_[14492]_ , \new_[14493]_ , \new_[14494]_ , \new_[14495]_ ,
    \new_[14496]_ , \new_[14497]_ , \new_[14498]_ , \new_[14499]_ ,
    \new_[14500]_ , \new_[14501]_ , \new_[14502]_ , \new_[14503]_ ,
    \new_[14504]_ , \new_[14505]_ , \new_[14506]_ , \new_[14507]_ ,
    \new_[14508]_ , \new_[14509]_ , \new_[14510]_ , \new_[14511]_ ,
    \new_[14512]_ , \new_[14513]_ , \new_[14514]_ , \new_[14515]_ ,
    \new_[14516]_ , \new_[14517]_ , \new_[14518]_ , \new_[14519]_ ,
    \new_[14520]_ , \new_[14521]_ , \new_[14522]_ , \new_[14523]_ ,
    \new_[14524]_ , \new_[14525]_ , \new_[14526]_ , \new_[14527]_ ,
    \new_[14528]_ , \new_[14529]_ , \new_[14530]_ , \new_[14531]_ ,
    \new_[14532]_ , \new_[14533]_ , \new_[14534]_ , \new_[14535]_ ,
    \new_[14536]_ , \new_[14537]_ , \new_[14538]_ , \new_[14539]_ ,
    \new_[14540]_ , \new_[14541]_ , \new_[14542]_ , \new_[14543]_ ,
    \new_[14544]_ , \new_[14545]_ , \new_[14546]_ , \new_[14547]_ ,
    \new_[14548]_ , \new_[14549]_ , \new_[14550]_ , \new_[14551]_ ,
    \new_[14552]_ , \new_[14553]_ , \new_[14554]_ , \new_[14555]_ ,
    \new_[14556]_ , \new_[14557]_ , \new_[14558]_ , \new_[14559]_ ,
    \new_[14560]_ , \new_[14562]_ , \new_[14563]_ , \new_[14564]_ ,
    \new_[14565]_ , \new_[14566]_ , \new_[14567]_ , \new_[14568]_ ,
    \new_[14569]_ , \new_[14572]_ , \new_[14573]_ , \new_[14574]_ ,
    \new_[14575]_ , \new_[14576]_ , \new_[14577]_ , \new_[14578]_ ,
    \new_[14579]_ , \new_[14580]_ , \new_[14581]_ , \new_[14582]_ ,
    \new_[14583]_ , \new_[14584]_ , \new_[14585]_ , \new_[14586]_ ,
    \new_[14587]_ , \new_[14588]_ , \new_[14589]_ , \new_[14590]_ ,
    \new_[14591]_ , \new_[14592]_ , \new_[14593]_ , \new_[14594]_ ,
    \new_[14595]_ , \new_[14596]_ , \new_[14597]_ , \new_[14598]_ ,
    \new_[14599]_ , \new_[14600]_ , \new_[14601]_ , \new_[14602]_ ,
    \new_[14603]_ , \new_[14604]_ , \new_[14605]_ , \new_[14606]_ ,
    \new_[14607]_ , \new_[14608]_ , \new_[14609]_ , \new_[14610]_ ,
    \new_[14611]_ , \new_[14612]_ , \new_[14613]_ , \new_[14614]_ ,
    \new_[14615]_ , \new_[14616]_ , \new_[14617]_ , \new_[14618]_ ,
    \new_[14619]_ , \new_[14620]_ , \new_[14621]_ , \new_[14622]_ ,
    \new_[14623]_ , \new_[14624]_ , \new_[14625]_ , \new_[14626]_ ,
    \new_[14627]_ , \new_[14628]_ , \new_[14629]_ , \new_[14630]_ ,
    \new_[14631]_ , \new_[14632]_ , \new_[14633]_ , \new_[14634]_ ,
    \new_[14635]_ , \new_[14636]_ , \new_[14637]_ , \new_[14638]_ ,
    \new_[14639]_ , \new_[14640]_ , \new_[14641]_ , \new_[14642]_ ,
    \new_[14643]_ , \new_[14644]_ , \new_[14645]_ , \new_[14646]_ ,
    \new_[14647]_ , \new_[14648]_ , \new_[14649]_ , \new_[14650]_ ,
    \new_[14651]_ , \new_[14652]_ , \new_[14653]_ , \new_[14654]_ ,
    \new_[14655]_ , \new_[14656]_ , \new_[14657]_ , \new_[14658]_ ,
    \new_[14659]_ , \new_[14660]_ , \new_[14661]_ , \new_[14662]_ ,
    \new_[14663]_ , \new_[14664]_ , \new_[14665]_ , \new_[14666]_ ,
    \new_[14667]_ , \new_[14668]_ , \new_[14669]_ , \new_[14670]_ ,
    \new_[14671]_ , \new_[14672]_ , \new_[14673]_ , \new_[14674]_ ,
    \new_[14675]_ , \new_[14676]_ , \new_[14677]_ , \new_[14678]_ ,
    \new_[14679]_ , \new_[14680]_ , \new_[14681]_ , \new_[14682]_ ,
    \new_[14683]_ , \new_[14684]_ , \new_[14685]_ , \new_[14686]_ ,
    \new_[14687]_ , \new_[14688]_ , \new_[14689]_ , \new_[14690]_ ,
    \new_[14691]_ , \new_[14692]_ , \new_[14693]_ , \new_[14694]_ ,
    \new_[14695]_ , \new_[14696]_ , \new_[14697]_ , \new_[14698]_ ,
    \new_[14699]_ , \new_[14700]_ , \new_[14701]_ , \new_[14702]_ ,
    \new_[14703]_ , \new_[14704]_ , \new_[14705]_ , \new_[14706]_ ,
    \new_[14707]_ , \new_[14708]_ , \new_[14709]_ , \new_[14710]_ ,
    \new_[14711]_ , \new_[14712]_ , \new_[14713]_ , \new_[14714]_ ,
    \new_[14715]_ , \new_[14716]_ , \new_[14717]_ , \new_[14718]_ ,
    \new_[14719]_ , \new_[14720]_ , \new_[14721]_ , \new_[14722]_ ,
    \new_[14723]_ , \new_[14724]_ , \new_[14725]_ , \new_[14726]_ ,
    \new_[14727]_ , \new_[14728]_ , \new_[14729]_ , \new_[14730]_ ,
    \new_[14731]_ , \new_[14732]_ , \new_[14733]_ , \new_[14734]_ ,
    \new_[14735]_ , \new_[14736]_ , \new_[14737]_ , \new_[14738]_ ,
    \new_[14739]_ , \new_[14740]_ , \new_[14741]_ , \new_[14742]_ ,
    \new_[14743]_ , \new_[14744]_ , \new_[14745]_ , \new_[14746]_ ,
    \new_[14747]_ , \new_[14748]_ , \new_[14749]_ , \new_[14750]_ ,
    \new_[14751]_ , \new_[14752]_ , \new_[14753]_ , \new_[14754]_ ,
    \new_[14755]_ , \new_[14756]_ , \new_[14757]_ , \new_[14758]_ ,
    \new_[14759]_ , \new_[14760]_ , \new_[14761]_ , \new_[14762]_ ,
    \new_[14763]_ , \new_[14764]_ , \new_[14765]_ , \new_[14766]_ ,
    \new_[14767]_ , \new_[14768]_ , \new_[14769]_ , \new_[14770]_ ,
    \new_[14771]_ , \new_[14772]_ , \new_[14773]_ , \new_[14774]_ ,
    \new_[14775]_ , \new_[14776]_ , \new_[14777]_ , \new_[14778]_ ,
    \new_[14779]_ , \new_[14780]_ , \new_[14781]_ , \new_[14782]_ ,
    \new_[14783]_ , \new_[14784]_ , \new_[14785]_ , \new_[14786]_ ,
    \new_[14787]_ , \new_[14788]_ , \new_[14789]_ , \new_[14790]_ ,
    \new_[14791]_ , \new_[14792]_ , \new_[14793]_ , \new_[14794]_ ,
    \new_[14795]_ , \new_[14796]_ , \new_[14797]_ , \new_[14798]_ ,
    \new_[14799]_ , \new_[14800]_ , \new_[14801]_ , \new_[14802]_ ,
    \new_[14803]_ , \new_[14804]_ , \new_[14805]_ , \new_[14806]_ ,
    \new_[14807]_ , \new_[14808]_ , \new_[14809]_ , \new_[14810]_ ,
    \new_[14811]_ , \new_[14812]_ , \new_[14813]_ , \new_[14814]_ ,
    \new_[14815]_ , \new_[14816]_ , \new_[14817]_ , \new_[14818]_ ,
    \new_[14819]_ , \new_[14820]_ , \new_[14821]_ , \new_[14822]_ ,
    \new_[14823]_ , \new_[14824]_ , \new_[14825]_ , \new_[14826]_ ,
    \new_[14827]_ , \new_[14828]_ , \new_[14829]_ , \new_[14830]_ ,
    \new_[14831]_ , \new_[14832]_ , \new_[14833]_ , \new_[14834]_ ,
    \new_[14835]_ , \new_[14836]_ , \new_[14837]_ , \new_[14838]_ ,
    \new_[14839]_ , \new_[14840]_ , \new_[14843]_ , \new_[14844]_ ,
    \new_[14845]_ , \new_[14846]_ , \new_[14847]_ , \new_[14849]_ ,
    \new_[14850]_ , \new_[14851]_ , \new_[14852]_ , \new_[14853]_ ,
    \new_[14854]_ , \new_[14855]_ , \new_[14856]_ , \new_[14857]_ ,
    \new_[14858]_ , \new_[14859]_ , \new_[14860]_ , \new_[14861]_ ,
    \new_[14862]_ , \new_[14863]_ , \new_[14864]_ , \new_[14865]_ ,
    \new_[14866]_ , \new_[14867]_ , \new_[14868]_ , \new_[14869]_ ,
    \new_[14870]_ , \new_[14871]_ , \new_[14872]_ , \new_[14873]_ ,
    \new_[14874]_ , \new_[14875]_ , \new_[14876]_ , \new_[14877]_ ,
    \new_[14878]_ , \new_[14879]_ , \new_[14880]_ , \new_[14881]_ ,
    \new_[14882]_ , \new_[14883]_ , \new_[14884]_ , \new_[14885]_ ,
    \new_[14886]_ , \new_[14887]_ , \new_[14888]_ , \new_[14889]_ ,
    \new_[14890]_ , \new_[14891]_ , \new_[14892]_ , \new_[14893]_ ,
    \new_[14894]_ , \new_[14895]_ , \new_[14896]_ , \new_[14897]_ ,
    \new_[14898]_ , \new_[14899]_ , \new_[14900]_ , \new_[14901]_ ,
    \new_[14902]_ , \new_[14903]_ , \new_[14904]_ , \new_[14905]_ ,
    \new_[14906]_ , \new_[14907]_ , \new_[14908]_ , \new_[14909]_ ,
    \new_[14910]_ , \new_[14911]_ , \new_[14912]_ , \new_[14913]_ ,
    \new_[14914]_ , \new_[14915]_ , \new_[14916]_ , \new_[14917]_ ,
    \new_[14918]_ , \new_[14919]_ , \new_[14920]_ , \new_[14921]_ ,
    \new_[14922]_ , \new_[14923]_ , \new_[14924]_ , \new_[14925]_ ,
    \new_[14926]_ , \new_[14927]_ , \new_[14928]_ , \new_[14929]_ ,
    \new_[14930]_ , \new_[14931]_ , \new_[14932]_ , \new_[14933]_ ,
    \new_[14934]_ , \new_[14935]_ , \new_[14936]_ , \new_[14937]_ ,
    \new_[14938]_ , \new_[14939]_ , \new_[14940]_ , \new_[14941]_ ,
    \new_[14942]_ , \new_[14943]_ , \new_[14944]_ , \new_[14945]_ ,
    \new_[14946]_ , \new_[14947]_ , \new_[14948]_ , \new_[14949]_ ,
    \new_[14950]_ , \new_[14951]_ , \new_[14952]_ , \new_[14953]_ ,
    \new_[14955]_ , \new_[14956]_ , \new_[14957]_ , \new_[14958]_ ,
    \new_[14959]_ , \new_[14960]_ , \new_[14961]_ , \new_[14962]_ ,
    \new_[14963]_ , \new_[14964]_ , \new_[14965]_ , \new_[14966]_ ,
    \new_[14967]_ , \new_[14969]_ , \new_[14970]_ , \new_[14971]_ ,
    \new_[14972]_ , \new_[14973]_ , \new_[14974]_ , \new_[14975]_ ,
    \new_[14976]_ , \new_[14978]_ , \new_[14979]_ , \new_[14980]_ ,
    \new_[14981]_ , \new_[14982]_ , \new_[14983]_ , \new_[14984]_ ,
    \new_[14985]_ , \new_[14986]_ , \new_[14987]_ , \new_[14988]_ ,
    \new_[14989]_ , \new_[14990]_ , \new_[14991]_ , \new_[14992]_ ,
    \new_[14993]_ , \new_[14994]_ , \new_[14995]_ , \new_[14996]_ ,
    \new_[14997]_ , \new_[14998]_ , \new_[14999]_ , \new_[15000]_ ,
    \new_[15001]_ , \new_[15002]_ , \new_[15003]_ , \new_[15004]_ ,
    \new_[15005]_ , \new_[15006]_ , \new_[15007]_ , \new_[15008]_ ,
    \new_[15009]_ , \new_[15010]_ , \new_[15011]_ , \new_[15012]_ ,
    \new_[15013]_ , \new_[15014]_ , \new_[15015]_ , \new_[15016]_ ,
    \new_[15017]_ , \new_[15018]_ , \new_[15019]_ , \new_[15020]_ ,
    \new_[15021]_ , \new_[15022]_ , \new_[15024]_ , \new_[15025]_ ,
    \new_[15026]_ , \new_[15027]_ , \new_[15028]_ , \new_[15029]_ ,
    \new_[15030]_ , \new_[15031]_ , \new_[15032]_ , \new_[15033]_ ,
    \new_[15034]_ , \new_[15035]_ , \new_[15036]_ , \new_[15037]_ ,
    \new_[15038]_ , \new_[15039]_ , \new_[15040]_ , \new_[15041]_ ,
    \new_[15042]_ , \new_[15043]_ , \new_[15044]_ , \new_[15045]_ ,
    \new_[15046]_ , \new_[15047]_ , \new_[15048]_ , \new_[15049]_ ,
    \new_[15050]_ , \new_[15051]_ , \new_[15052]_ , \new_[15053]_ ,
    \new_[15054]_ , \new_[15055]_ , \new_[15056]_ , \new_[15057]_ ,
    \new_[15059]_ , \new_[15060]_ , \new_[15061]_ , \new_[15062]_ ,
    \new_[15063]_ , \new_[15064]_ , \new_[15065]_ , \new_[15066]_ ,
    \new_[15067]_ , \new_[15068]_ , \new_[15069]_ , \new_[15070]_ ,
    \new_[15071]_ , \new_[15072]_ , \new_[15073]_ , \new_[15074]_ ,
    \new_[15075]_ , \new_[15076]_ , \new_[15077]_ , \new_[15078]_ ,
    \new_[15079]_ , \new_[15080]_ , \new_[15081]_ , \new_[15082]_ ,
    \new_[15083]_ , \new_[15084]_ , \new_[15085]_ , \new_[15086]_ ,
    \new_[15087]_ , \new_[15088]_ , \new_[15089]_ , \new_[15090]_ ,
    \new_[15091]_ , \new_[15092]_ , \new_[15093]_ , \new_[15094]_ ,
    \new_[15095]_ , \new_[15096]_ , \new_[15097]_ , \new_[15098]_ ,
    \new_[15100]_ , \new_[15104]_ , \new_[15105]_ , \new_[15106]_ ,
    \new_[15107]_ , \new_[15108]_ , \new_[15109]_ , \new_[15110]_ ,
    \new_[15111]_ , \new_[15112]_ , \new_[15113]_ , \new_[15114]_ ,
    \new_[15115]_ , \new_[15116]_ , \new_[15117]_ , \new_[15118]_ ,
    \new_[15119]_ , \new_[15120]_ , \new_[15121]_ , \new_[15122]_ ,
    \new_[15123]_ , \new_[15124]_ , \new_[15125]_ , \new_[15126]_ ,
    \new_[15127]_ , \new_[15128]_ , \new_[15129]_ , \new_[15130]_ ,
    \new_[15131]_ , \new_[15132]_ , \new_[15133]_ , \new_[15134]_ ,
    \new_[15135]_ , \new_[15136]_ , \new_[15137]_ , \new_[15138]_ ,
    \new_[15139]_ , \new_[15140]_ , \new_[15141]_ , \new_[15142]_ ,
    \new_[15143]_ , \new_[15144]_ , \new_[15145]_ , \new_[15146]_ ,
    \new_[15147]_ , \new_[15148]_ , \new_[15149]_ , \new_[15150]_ ,
    \new_[15151]_ , \new_[15152]_ , \new_[15153]_ , \new_[15154]_ ,
    \new_[15156]_ , \new_[15157]_ , \new_[15158]_ , \new_[15159]_ ,
    \new_[15160]_ , \new_[15161]_ , \new_[15162]_ , \new_[15163]_ ,
    \new_[15164]_ , \new_[15165]_ , \new_[15166]_ , \new_[15167]_ ,
    \new_[15168]_ , \new_[15169]_ , \new_[15170]_ , \new_[15171]_ ,
    \new_[15172]_ , \new_[15173]_ , \new_[15174]_ , \new_[15175]_ ,
    \new_[15176]_ , \new_[15177]_ , \new_[15178]_ , \new_[15179]_ ,
    \new_[15180]_ , \new_[15181]_ , \new_[15182]_ , \new_[15183]_ ,
    \new_[15185]_ , \new_[15186]_ , \new_[15187]_ , \new_[15188]_ ,
    \new_[15189]_ , \new_[15190]_ , \new_[15191]_ , \new_[15192]_ ,
    \new_[15193]_ , \new_[15194]_ , \new_[15195]_ , \new_[15196]_ ,
    \new_[15197]_ , \new_[15198]_ , \new_[15199]_ , \new_[15200]_ ,
    \new_[15201]_ , \new_[15202]_ , \new_[15203]_ , \new_[15204]_ ,
    \new_[15205]_ , \new_[15206]_ , \new_[15207]_ , \new_[15208]_ ,
    \new_[15209]_ , \new_[15210]_ , \new_[15211]_ , \new_[15212]_ ,
    \new_[15213]_ , \new_[15214]_ , \new_[15215]_ , \new_[15216]_ ,
    \new_[15217]_ , \new_[15218]_ , \new_[15219]_ , \new_[15220]_ ,
    \new_[15221]_ , \new_[15222]_ , \new_[15224]_ , \new_[15225]_ ,
    \new_[15226]_ , \new_[15227]_ , \new_[15228]_ , \new_[15229]_ ,
    \new_[15230]_ , \new_[15231]_ , \new_[15232]_ , \new_[15233]_ ,
    \new_[15234]_ , \new_[15235]_ , \new_[15236]_ , \new_[15237]_ ,
    \new_[15238]_ , \new_[15239]_ , \new_[15240]_ , \new_[15241]_ ,
    \new_[15242]_ , \new_[15243]_ , \new_[15244]_ , \new_[15245]_ ,
    \new_[15246]_ , \new_[15247]_ , \new_[15248]_ , \new_[15249]_ ,
    \new_[15250]_ , \new_[15251]_ , \new_[15252]_ , \new_[15253]_ ,
    \new_[15254]_ , \new_[15255]_ , \new_[15256]_ , \new_[15257]_ ,
    \new_[15258]_ , \new_[15259]_ , \new_[15261]_ , \new_[15262]_ ,
    \new_[15263]_ , \new_[15264]_ , \new_[15265]_ , \new_[15266]_ ,
    \new_[15267]_ , \new_[15268]_ , \new_[15269]_ , \new_[15270]_ ,
    \new_[15271]_ , \new_[15272]_ , \new_[15273]_ , \new_[15274]_ ,
    \new_[15275]_ , \new_[15276]_ , \new_[15277]_ , \new_[15278]_ ,
    \new_[15279]_ , \new_[15281]_ , \new_[15282]_ , \new_[15283]_ ,
    \new_[15284]_ , \new_[15285]_ , \new_[15286]_ , \new_[15287]_ ,
    \new_[15288]_ , \new_[15289]_ , \new_[15290]_ , \new_[15291]_ ,
    \new_[15292]_ , \new_[15293]_ , \new_[15294]_ , \new_[15295]_ ,
    \new_[15296]_ , \new_[15297]_ , \new_[15298]_ , \new_[15299]_ ,
    \new_[15300]_ , \new_[15301]_ , \new_[15302]_ , \new_[15303]_ ,
    \new_[15304]_ , \new_[15305]_ , \new_[15306]_ , \new_[15307]_ ,
    \new_[15308]_ , \new_[15309]_ , \new_[15310]_ , \new_[15311]_ ,
    \new_[15312]_ , \new_[15313]_ , \new_[15314]_ , \new_[15315]_ ,
    \new_[15316]_ , \new_[15317]_ , \new_[15318]_ , \new_[15319]_ ,
    \new_[15320]_ , \new_[15321]_ , \new_[15322]_ , \new_[15323]_ ,
    \new_[15324]_ , \new_[15325]_ , \new_[15326]_ , \new_[15327]_ ,
    \new_[15329]_ , \new_[15330]_ , \new_[15331]_ , \new_[15332]_ ,
    \new_[15333]_ , \new_[15334]_ , \new_[15335]_ , \new_[15336]_ ,
    \new_[15337]_ , \new_[15338]_ , \new_[15339]_ , \new_[15340]_ ,
    \new_[15341]_ , \new_[15342]_ , \new_[15343]_ , \new_[15344]_ ,
    \new_[15345]_ , \new_[15346]_ , \new_[15347]_ , \new_[15348]_ ,
    \new_[15349]_ , \new_[15351]_ , \new_[15352]_ , \new_[15353]_ ,
    \new_[15354]_ , \new_[15355]_ , \new_[15356]_ , \new_[15357]_ ,
    \new_[15358]_ , \new_[15359]_ , \new_[15360]_ , \new_[15361]_ ,
    \new_[15362]_ , \new_[15363]_ , \new_[15364]_ , \new_[15365]_ ,
    \new_[15366]_ , \new_[15367]_ , \new_[15368]_ , \new_[15369]_ ,
    \new_[15370]_ , \new_[15371]_ , \new_[15372]_ , \new_[15373]_ ,
    \new_[15374]_ , \new_[15375]_ , \new_[15376]_ , \new_[15377]_ ,
    \new_[15378]_ , \new_[15379]_ , \new_[15380]_ , \new_[15381]_ ,
    \new_[15382]_ , \new_[15383]_ , \new_[15384]_ , \new_[15385]_ ,
    \new_[15387]_ , \new_[15388]_ , \new_[15389]_ , \new_[15390]_ ,
    \new_[15391]_ , \new_[15392]_ , \new_[15393]_ , \new_[15394]_ ,
    \new_[15395]_ , \new_[15396]_ , \new_[15397]_ , \new_[15398]_ ,
    \new_[15399]_ , \new_[15400]_ , \new_[15401]_ , \new_[15402]_ ,
    \new_[15403]_ , \new_[15404]_ , \new_[15405]_ , \new_[15406]_ ,
    \new_[15407]_ , \new_[15408]_ , \new_[15409]_ , \new_[15410]_ ,
    \new_[15411]_ , \new_[15412]_ , \new_[15413]_ , \new_[15414]_ ,
    \new_[15415]_ , \new_[15417]_ , \new_[15418]_ , \new_[15420]_ ,
    \new_[15422]_ , \new_[15423]_ , \new_[15424]_ , \new_[15425]_ ,
    \new_[15426]_ , \new_[15427]_ , \new_[15428]_ , \new_[15429]_ ,
    \new_[15430]_ , \new_[15431]_ , \new_[15432]_ , \new_[15433]_ ,
    \new_[15434]_ , \new_[15435]_ , \new_[15438]_ , \new_[15439]_ ,
    \new_[15440]_ , \new_[15442]_ , \new_[15443]_ , \new_[15444]_ ,
    \new_[15445]_ , \new_[15446]_ , \new_[15447]_ , \new_[15450]_ ,
    \new_[15451]_ , \new_[15453]_ , \new_[15454]_ , \new_[15455]_ ,
    \new_[15456]_ , \new_[15457]_ , \new_[15458]_ , \new_[15459]_ ,
    \new_[15460]_ , \new_[15461]_ , \new_[15462]_ , \new_[15463]_ ,
    \new_[15464]_ , \new_[15465]_ , \new_[15466]_ , \new_[15467]_ ,
    \new_[15468]_ , \new_[15469]_ , \new_[15470]_ , \new_[15471]_ ,
    \new_[15472]_ , \new_[15473]_ , \new_[15474]_ , \new_[15475]_ ,
    \new_[15476]_ , \new_[15477]_ , \new_[15478]_ , \new_[15479]_ ,
    \new_[15480]_ , \new_[15482]_ , \new_[15483]_ , \new_[15484]_ ,
    \new_[15485]_ , \new_[15486]_ , \new_[15487]_ , \new_[15488]_ ,
    \new_[15489]_ , \new_[15491]_ , \new_[15492]_ , \new_[15493]_ ,
    \new_[15494]_ , \new_[15495]_ , \new_[15496]_ , \new_[15497]_ ,
    \new_[15498]_ , \new_[15499]_ , \new_[15500]_ , \new_[15501]_ ,
    \new_[15502]_ , \new_[15503]_ , \new_[15504]_ , \new_[15505]_ ,
    \new_[15506]_ , \new_[15507]_ , \new_[15508]_ , \new_[15509]_ ,
    \new_[15510]_ , \new_[15511]_ , \new_[15512]_ , \new_[15513]_ ,
    \new_[15514]_ , \new_[15515]_ , \new_[15516]_ , \new_[15517]_ ,
    \new_[15518]_ , \new_[15519]_ , \new_[15520]_ , \new_[15521]_ ,
    \new_[15522]_ , \new_[15523]_ , \new_[15524]_ , \new_[15525]_ ,
    \new_[15526]_ , \new_[15527]_ , \new_[15528]_ , \new_[15529]_ ,
    \new_[15530]_ , \new_[15531]_ , \new_[15532]_ , \new_[15533]_ ,
    \new_[15534]_ , \new_[15535]_ , \new_[15536]_ , \new_[15537]_ ,
    \new_[15538]_ , \new_[15539]_ , \new_[15540]_ , \new_[15541]_ ,
    \new_[15542]_ , \new_[15543]_ , \new_[15544]_ , \new_[15545]_ ,
    \new_[15547]_ , \new_[15548]_ , \new_[15549]_ , \new_[15550]_ ,
    \new_[15561]_ , \new_[15563]_ , \new_[15564]_ , \new_[15566]_ ,
    \new_[15568]_ , \new_[15569]_ , \new_[15570]_ , \new_[15572]_ ,
    \new_[15573]_ , \new_[15574]_ , \new_[15575]_ , \new_[15576]_ ,
    \new_[15577]_ , \new_[15578]_ , \new_[15579]_ , \new_[15580]_ ,
    \new_[15582]_ , \new_[15583]_ , \new_[15584]_ , \new_[15585]_ ,
    \new_[15586]_ , \new_[15588]_ , \new_[15590]_ , \new_[15591]_ ,
    \new_[15592]_ , \new_[15593]_ , \new_[15594]_ , \new_[15595]_ ,
    \new_[15596]_ , \new_[15598]_ , \new_[15599]_ , \new_[15601]_ ,
    \new_[15602]_ , \new_[15603]_ , \new_[15604]_ , \new_[15605]_ ,
    \new_[15606]_ , \new_[15607]_ , \new_[15608]_ , \new_[15609]_ ,
    \new_[15610]_ , \new_[15612]_ , \new_[15613]_ , \new_[15614]_ ,
    \new_[15615]_ , \new_[15616]_ , \new_[15617]_ , \new_[15618]_ ,
    \new_[15619]_ , \new_[15620]_ , \new_[15621]_ , \new_[15622]_ ,
    \new_[15623]_ , \new_[15624]_ , \new_[15625]_ , \new_[15626]_ ,
    \new_[15627]_ , \new_[15628]_ , \new_[15629]_ , \new_[15630]_ ,
    \new_[15631]_ , \new_[15632]_ , \new_[15633]_ , \new_[15634]_ ,
    \new_[15637]_ , \new_[15638]_ , \new_[15679]_ , \new_[15680]_ ,
    \new_[15681]_ , \new_[15682]_ , \new_[15683]_ , \new_[15684]_ ,
    \new_[15685]_ , \new_[15686]_ , \new_[15687]_ , \new_[15688]_ ,
    \new_[15689]_ , \new_[15690]_ , \new_[15691]_ , \new_[15692]_ ,
    \new_[15693]_ , \new_[15694]_ , \new_[15695]_ , \new_[15696]_ ,
    \new_[15699]_ , \new_[15704]_ , \new_[15706]_ , \new_[15720]_ ,
    \new_[15734]_ , \new_[15735]_ , \new_[15736]_ , \new_[15737]_ ,
    \new_[15738]_ , \new_[15739]_ , \new_[15740]_ , \new_[15741]_ ,
    \new_[15742]_ , \new_[15743]_ , \new_[15744]_ , \new_[15745]_ ,
    \new_[15746]_ , \new_[15747]_ , \new_[15749]_ , \new_[15783]_ ,
    \new_[15784]_ , \new_[15785]_ , \new_[15786]_ , \new_[15787]_ ,
    \new_[15788]_ , \new_[15789]_ , \new_[15790]_ , \new_[15791]_ ,
    \new_[15792]_ , \new_[15794]_ , \new_[15795]_ , \new_[15796]_ ,
    \new_[15797]_ , \new_[15798]_ , \new_[15800]_ , \new_[15801]_ ,
    \new_[15802]_ , \new_[15803]_ , \new_[15804]_ , \new_[15805]_ ,
    \new_[15806]_ , \new_[15807]_ , \new_[15808]_ , \new_[15809]_ ,
    \new_[15810]_ , \new_[15811]_ , \new_[15812]_ , \new_[15814]_ ,
    \new_[15815]_ , \new_[15816]_ , \new_[15817]_ , \new_[15818]_ ,
    \new_[15819]_ , \new_[15820]_ , \new_[15821]_ , \new_[15822]_ ,
    \new_[15823]_ , \new_[15824]_ , \new_[15825]_ , \new_[15826]_ ,
    \new_[15827]_ , \new_[15828]_ , \new_[15829]_ , \new_[15830]_ ,
    \new_[15831]_ , \new_[15832]_ , \new_[15833]_ , \new_[15834]_ ,
    \new_[15835]_ , \new_[15836]_ , \new_[15837]_ , \new_[15838]_ ,
    \new_[15840]_ , \new_[15841]_ , \new_[15842]_ , \new_[15843]_ ,
    \new_[15844]_ , \new_[15845]_ , \new_[15846]_ , \new_[15847]_ ,
    \new_[15848]_ , \new_[15849]_ , \new_[15850]_ , \new_[15851]_ ,
    \new_[15852]_ , \new_[15853]_ , \new_[15854]_ , \new_[15855]_ ,
    \new_[15856]_ , \new_[15857]_ , \new_[15859]_ , \new_[15860]_ ,
    \new_[15861]_ , \new_[15862]_ , \new_[15863]_ , \new_[15866]_ ,
    \new_[15867]_ , \new_[15868]_ , \new_[15869]_ , \new_[15870]_ ,
    \new_[15871]_ , \new_[15872]_ , \new_[15873]_ , \new_[15874]_ ,
    \new_[15875]_ , \new_[15876]_ , \new_[15877]_ , \new_[15878]_ ,
    \new_[15879]_ , \new_[15880]_ , \new_[15881]_ , \new_[15882]_ ,
    \new_[15883]_ , \new_[15884]_ , \new_[15885]_ , \new_[15886]_ ,
    \new_[15887]_ , \new_[15888]_ , \new_[15889]_ , \new_[15890]_ ,
    \new_[15891]_ , \new_[15892]_ , \new_[15893]_ , \new_[15894]_ ,
    \new_[15895]_ , \new_[15896]_ , \new_[15897]_ , \new_[15898]_ ,
    \new_[15899]_ , \new_[15900]_ , \new_[15901]_ , \new_[15902]_ ,
    \new_[15903]_ , \new_[15904]_ , \new_[15905]_ , \new_[15906]_ ,
    \new_[15907]_ , \new_[15908]_ , \new_[15909]_ , \new_[15910]_ ,
    \new_[15911]_ , \new_[15912]_ , \new_[15913]_ , \new_[15914]_ ,
    \new_[15915]_ , \new_[15916]_ , \new_[15917]_ , \new_[15918]_ ,
    \new_[15919]_ , \new_[15920]_ , \new_[15921]_ , \new_[15922]_ ,
    \new_[15923]_ , \new_[15924]_ , \new_[15925]_ , \new_[15926]_ ,
    \new_[15927]_ , \new_[15928]_ , \new_[15929]_ , \new_[15930]_ ,
    \new_[15931]_ , \new_[15932]_ , \new_[15933]_ , \new_[15934]_ ,
    \new_[15935]_ , \new_[15937]_ , \new_[15938]_ , \new_[15939]_ ,
    \new_[15940]_ , \new_[15941]_ , \new_[15942]_ , \new_[15943]_ ,
    \new_[15944]_ , \new_[15945]_ , \new_[15946]_ , \new_[15947]_ ,
    \new_[15948]_ , \new_[15949]_ , \new_[15950]_ , \new_[15951]_ ,
    \new_[15952]_ , \new_[15953]_ , \new_[15954]_ , \new_[15955]_ ,
    \new_[15956]_ , \new_[15957]_ , \new_[15958]_ , \new_[15959]_ ,
    \new_[15960]_ , \new_[15961]_ , \new_[15962]_ , \new_[15963]_ ,
    \new_[15964]_ , \new_[15965]_ , \new_[15967]_ , \new_[15968]_ ,
    \new_[15970]_ , \new_[15971]_ , \new_[15972]_ , \new_[15973]_ ,
    \new_[15974]_ , \new_[15975]_ , \new_[15976]_ , \new_[15977]_ ,
    \new_[15978]_ , \new_[15979]_ , \new_[15980]_ , \new_[15981]_ ,
    \new_[15982]_ , \new_[15983]_ , \new_[15984]_ , \new_[15985]_ ,
    \new_[15986]_ , \new_[15987]_ , \new_[15988]_ , \new_[15989]_ ,
    \new_[15990]_ , \new_[15991]_ , \new_[15992]_ , \new_[15993]_ ,
    \new_[15994]_ , \new_[15995]_ , \new_[15996]_ , \new_[15997]_ ,
    \new_[15998]_ , \new_[15999]_ , \new_[16000]_ , \new_[16001]_ ,
    \new_[16002]_ , \new_[16003]_ , \new_[16004]_ , \new_[16005]_ ,
    \new_[16006]_ , \new_[16007]_ , \new_[16008]_ , \new_[16009]_ ,
    \new_[16010]_ , \new_[16011]_ , \new_[16012]_ , \new_[16013]_ ,
    \new_[16014]_ , \new_[16015]_ , \new_[16016]_ , \new_[16017]_ ,
    \new_[16018]_ , \new_[16019]_ , \new_[16020]_ , \new_[16021]_ ,
    \new_[16022]_ , \new_[16023]_ , \new_[16024]_ , \new_[16025]_ ,
    \new_[16026]_ , \new_[16027]_ , \new_[16028]_ , \new_[16029]_ ,
    \new_[16030]_ , \new_[16031]_ , \new_[16032]_ , \new_[16033]_ ,
    \new_[16034]_ , \new_[16035]_ , \new_[16036]_ , \new_[16037]_ ,
    \new_[16038]_ , \new_[16039]_ , \new_[16040]_ , \new_[16041]_ ,
    \new_[16042]_ , \new_[16043]_ , \new_[16044]_ , \new_[16045]_ ,
    \new_[16046]_ , \new_[16047]_ , \new_[16048]_ , \new_[16049]_ ,
    \new_[16050]_ , \new_[16051]_ , \new_[16052]_ , \new_[16053]_ ,
    \new_[16054]_ , \new_[16055]_ , \new_[16056]_ , \new_[16057]_ ,
    \new_[16058]_ , \new_[16059]_ , \new_[16061]_ , \new_[16062]_ ,
    \new_[16063]_ , \new_[16064]_ , \new_[16065]_ , \new_[16066]_ ,
    \new_[16067]_ , \new_[16068]_ , \new_[16069]_ , \new_[16070]_ ,
    \new_[16071]_ , \new_[16072]_ , \new_[16073]_ , \new_[16074]_ ,
    \new_[16075]_ , \new_[16076]_ , \new_[16077]_ , \new_[16078]_ ,
    \new_[16079]_ , \new_[16080]_ , \new_[16081]_ , \new_[16082]_ ,
    \new_[16083]_ , \new_[16084]_ , \new_[16085]_ , \new_[16086]_ ,
    \new_[16087]_ , \new_[16088]_ , \new_[16089]_ , \new_[16090]_ ,
    \new_[16091]_ , \new_[16092]_ , \new_[16093]_ , \new_[16094]_ ,
    \new_[16095]_ , \new_[16096]_ , \new_[16097]_ , \new_[16098]_ ,
    \new_[16099]_ , \new_[16100]_ , \new_[16101]_ , \new_[16102]_ ,
    \new_[16103]_ , \new_[16104]_ , \new_[16105]_ , \new_[16106]_ ,
    \new_[16107]_ , \new_[16108]_ , \new_[16109]_ , \new_[16110]_ ,
    \new_[16111]_ , \new_[16112]_ , \new_[16113]_ , \new_[16114]_ ,
    \new_[16115]_ , \new_[16116]_ , \new_[16117]_ , \new_[16118]_ ,
    \new_[16119]_ , \new_[16120]_ , \new_[16121]_ , \new_[16122]_ ,
    \new_[16123]_ , \new_[16124]_ , \new_[16125]_ , \new_[16126]_ ,
    \new_[16127]_ , \new_[16128]_ , \new_[16129]_ , \new_[16130]_ ,
    \new_[16131]_ , \new_[16132]_ , \new_[16133]_ , \new_[16134]_ ,
    \new_[16135]_ , \new_[16136]_ , \new_[16137]_ , \new_[16139]_ ,
    \new_[16140]_ , \new_[16141]_ , \new_[16142]_ , \new_[16143]_ ,
    \new_[16144]_ , \new_[16145]_ , \new_[16146]_ , \new_[16147]_ ,
    \new_[16148]_ , \new_[16149]_ , \new_[16150]_ , \new_[16151]_ ,
    \new_[16152]_ , \new_[16153]_ , \new_[16154]_ , \new_[16155]_ ,
    \new_[16156]_ , \new_[16157]_ , \new_[16158]_ , \new_[16159]_ ,
    \new_[16160]_ , \new_[16161]_ , \new_[16162]_ , \new_[16163]_ ,
    \new_[16164]_ , \new_[16165]_ , \new_[16166]_ , \new_[16167]_ ,
    \new_[16168]_ , \new_[16169]_ , \new_[16170]_ , \new_[16171]_ ,
    \new_[16172]_ , \new_[16173]_ , \new_[16174]_ , \new_[16175]_ ,
    \new_[16176]_ , \new_[16177]_ , \new_[16178]_ , \new_[16179]_ ,
    \new_[16180]_ , \new_[16181]_ , \new_[16182]_ , \new_[16183]_ ,
    \new_[16184]_ , \new_[16185]_ , \new_[16186]_ , \new_[16187]_ ,
    \new_[16188]_ , \new_[16189]_ , \new_[16190]_ , \new_[16191]_ ,
    \new_[16192]_ , \new_[16193]_ , \new_[16194]_ , \new_[16195]_ ,
    \new_[16196]_ , \new_[16197]_ , \new_[16198]_ , \new_[16199]_ ,
    \new_[16200]_ , \new_[16201]_ , \new_[16202]_ , \new_[16203]_ ,
    \new_[16204]_ , \new_[16205]_ , \new_[16206]_ , \new_[16207]_ ,
    \new_[16208]_ , \new_[16209]_ , \new_[16210]_ , \new_[16211]_ ,
    \new_[16212]_ , \new_[16213]_ , \new_[16214]_ , \new_[16215]_ ,
    \new_[16216]_ , \new_[16217]_ , \new_[16218]_ , \new_[16219]_ ,
    \new_[16220]_ , \new_[16221]_ , \new_[16222]_ , \new_[16223]_ ,
    \new_[16224]_ , \new_[16225]_ , \new_[16226]_ , \new_[16227]_ ,
    \new_[16228]_ , \new_[16229]_ , \new_[16230]_ , \new_[16231]_ ,
    \new_[16232]_ , \new_[16233]_ , \new_[16234]_ , \new_[16235]_ ,
    \new_[16236]_ , \new_[16237]_ , \new_[16238]_ , \new_[16239]_ ,
    \new_[16240]_ , \new_[16241]_ , \new_[16242]_ , \new_[16243]_ ,
    \new_[16244]_ , \new_[16245]_ , \new_[16246]_ , \new_[16247]_ ,
    \new_[16248]_ , \new_[16249]_ , \new_[16250]_ , \new_[16251]_ ,
    \new_[16252]_ , \new_[16253]_ , \new_[16254]_ , \new_[16255]_ ,
    \new_[16256]_ , \new_[16257]_ , \new_[16258]_ , \new_[16259]_ ,
    \new_[16260]_ , \new_[16261]_ , \new_[16262]_ , \new_[16263]_ ,
    \new_[16264]_ , \new_[16265]_ , \new_[16266]_ , \new_[16267]_ ,
    \new_[16268]_ , \new_[16269]_ , \new_[16270]_ , \new_[16271]_ ,
    \new_[16272]_ , \new_[16273]_ , \new_[16274]_ , \new_[16275]_ ,
    \new_[16276]_ , \new_[16277]_ , \new_[16278]_ , \new_[16279]_ ,
    \new_[16280]_ , \new_[16281]_ , \new_[16282]_ , \new_[16283]_ ,
    \new_[16284]_ , \new_[16285]_ , \new_[16286]_ , \new_[16287]_ ,
    \new_[16288]_ , \new_[16289]_ , \new_[16290]_ , \new_[16291]_ ,
    \new_[16292]_ , \new_[16293]_ , \new_[16294]_ , \new_[16295]_ ,
    \new_[16296]_ , \new_[16297]_ , \new_[16298]_ , \new_[16299]_ ,
    \new_[16300]_ , \new_[16301]_ , \new_[16302]_ , \new_[16303]_ ,
    \new_[16304]_ , \new_[16305]_ , \new_[16306]_ , \new_[16307]_ ,
    \new_[16308]_ , \new_[16309]_ , \new_[16310]_ , \new_[16311]_ ,
    \new_[16312]_ , \new_[16313]_ , \new_[16314]_ , \new_[16315]_ ,
    \new_[16316]_ , \new_[16317]_ , \new_[16318]_ , \new_[16319]_ ,
    \new_[16320]_ , \new_[16321]_ , \new_[16322]_ , \new_[16323]_ ,
    \new_[16324]_ , \new_[16325]_ , \new_[16326]_ , \new_[16327]_ ,
    \new_[16328]_ , \new_[16329]_ , \new_[16330]_ , \new_[16331]_ ,
    \new_[16332]_ , \new_[16333]_ , \new_[16334]_ , \new_[16335]_ ,
    \new_[16336]_ , \new_[16337]_ , \new_[16338]_ , \new_[16339]_ ,
    \new_[16340]_ , \new_[16341]_ , \new_[16342]_ , \new_[16343]_ ,
    \new_[16344]_ , \new_[16345]_ , \new_[16346]_ , \new_[16347]_ ,
    \new_[16348]_ , \new_[16349]_ , \new_[16350]_ , \new_[16351]_ ,
    \new_[16352]_ , \new_[16353]_ , \new_[16354]_ , \new_[16355]_ ,
    \new_[16356]_ , \new_[16357]_ , \new_[16358]_ , \new_[16359]_ ,
    \new_[16360]_ , \new_[16361]_ , \new_[16362]_ , \new_[16363]_ ,
    \new_[16364]_ , \new_[16365]_ , \new_[16366]_ , \new_[16367]_ ,
    \new_[16368]_ , \new_[16369]_ , \new_[16370]_ , \new_[16371]_ ,
    \new_[16372]_ , \new_[16373]_ , \new_[16374]_ , \new_[16375]_ ,
    \new_[16376]_ , \new_[16377]_ , \new_[16378]_ , \new_[16379]_ ,
    \new_[16380]_ , \new_[16381]_ , \new_[16382]_ , \new_[16383]_ ,
    \new_[16384]_ , \new_[16385]_ , \new_[16386]_ , \new_[16387]_ ,
    \new_[16388]_ , \new_[16389]_ , \new_[16390]_ , \new_[16391]_ ,
    \new_[16392]_ , \new_[16393]_ , \new_[16394]_ , \new_[16395]_ ,
    \new_[16396]_ , \new_[16397]_ , \new_[16398]_ , \new_[16399]_ ,
    \new_[16400]_ , \new_[16401]_ , \new_[16402]_ , \new_[16403]_ ,
    \new_[16404]_ , \new_[16405]_ , \new_[16406]_ , \new_[16407]_ ,
    \new_[16408]_ , \new_[16409]_ , \new_[16410]_ , \new_[16411]_ ,
    \new_[16412]_ , \new_[16413]_ , \new_[16414]_ , \new_[16415]_ ,
    \new_[16416]_ , \new_[16417]_ , \new_[16418]_ , \new_[16419]_ ,
    \new_[16420]_ , \new_[16421]_ , \new_[16422]_ , \new_[16423]_ ,
    \new_[16424]_ , \new_[16425]_ , \new_[16426]_ , \new_[16427]_ ,
    \new_[16428]_ , \new_[16429]_ , \new_[16430]_ , \new_[16431]_ ,
    \new_[16432]_ , \new_[16433]_ , \new_[16434]_ , \new_[16435]_ ,
    \new_[16436]_ , \new_[16437]_ , \new_[16438]_ , \new_[16440]_ ,
    \new_[16441]_ , \new_[16442]_ , \new_[16443]_ , \new_[16444]_ ,
    \new_[16445]_ , \new_[16446]_ , \new_[16447]_ , \new_[16448]_ ,
    \new_[16449]_ , \new_[16451]_ , \new_[16454]_ , \new_[16455]_ ,
    \new_[16456]_ , \new_[16457]_ , \new_[16458]_ , \new_[16459]_ ,
    \new_[16460]_ , \new_[16461]_ , \new_[16462]_ , \new_[16463]_ ,
    \new_[16464]_ , \new_[16465]_ , \new_[16469]_ , \new_[16470]_ ,
    \new_[16472]_ , \new_[16473]_ , \new_[16474]_ , \new_[16475]_ ,
    \new_[16476]_ , \new_[16477]_ , \new_[16478]_ , \new_[16479]_ ,
    \new_[16480]_ , \new_[16481]_ , \new_[16482]_ , \new_[16483]_ ,
    \new_[16484]_ , \new_[16485]_ , \new_[16486]_ , \new_[16487]_ ,
    \new_[16488]_ , \new_[16490]_ , \new_[16492]_ , \new_[16494]_ ,
    \new_[16496]_ , \new_[16497]_ , \new_[16498]_ , \new_[16499]_ ,
    \new_[16500]_ , \new_[16503]_ , \new_[16504]_ , \new_[16505]_ ,
    \new_[16506]_ , \new_[16508]_ , \new_[16509]_ , \new_[16510]_ ,
    \new_[16511]_ , \new_[16513]_ , \new_[16514]_ , \new_[16515]_ ,
    \new_[16516]_ , \new_[16517]_ , \new_[16519]_ , \new_[16520]_ ,
    \new_[16521]_ , \new_[16522]_ , \new_[16523]_ , \new_[16524]_ ,
    \new_[16525]_ , \new_[16526]_ , \new_[16527]_ , \new_[16528]_ ,
    \new_[16529]_ , \new_[16530]_ , \new_[16531]_ , \new_[16532]_ ,
    \new_[16533]_ , \new_[16534]_ , \new_[16535]_ , \new_[16536]_ ,
    \new_[16537]_ , \new_[16538]_ , \new_[16539]_ , \new_[16540]_ ,
    \new_[16541]_ , \new_[16542]_ , \new_[16543]_ , \new_[16544]_ ,
    \new_[16545]_ , \new_[16546]_ , \new_[16547]_ , \new_[16548]_ ,
    \new_[16549]_ , \new_[16550]_ , \new_[16551]_ , \new_[16552]_ ,
    \new_[16553]_ , \new_[16554]_ , \new_[16555]_ , \new_[16556]_ ,
    \new_[16557]_ , \new_[16558]_ , \new_[16559]_ , \new_[16560]_ ,
    \new_[16561]_ , \new_[16562]_ , \new_[16563]_ , \new_[16564]_ ,
    \new_[16565]_ , \new_[16566]_ , \new_[16567]_ , \new_[16568]_ ,
    \new_[16569]_ , \new_[16570]_ , \new_[16571]_ , \new_[16572]_ ,
    \new_[16573]_ , \new_[16574]_ , \new_[16575]_ , \new_[16576]_ ,
    \new_[16577]_ , \new_[16578]_ , \new_[16579]_ , \new_[16580]_ ,
    \new_[16581]_ , \new_[16582]_ , \new_[16583]_ , \new_[16584]_ ,
    \new_[16585]_ , \new_[16586]_ , \new_[16587]_ , \new_[16589]_ ,
    \new_[16590]_ , \new_[16591]_ , \new_[16592]_ , \new_[16593]_ ,
    \new_[16594]_ , \new_[16595]_ , \new_[16596]_ , \new_[16597]_ ,
    \new_[16598]_ , \new_[16599]_ , \new_[16600]_ , \new_[16602]_ ,
    \new_[16603]_ , \new_[16604]_ , \new_[16605]_ , \new_[16606]_ ,
    \new_[16607]_ , \new_[16608]_ , \new_[16609]_ , \new_[16610]_ ,
    \new_[16611]_ , \new_[16612]_ , \new_[16613]_ , \new_[16614]_ ,
    \new_[16615]_ , \new_[16616]_ , \new_[16617]_ , \new_[16618]_ ,
    \new_[16619]_ , \new_[16620]_ , \new_[16621]_ , \new_[16630]_ ,
    \new_[16631]_ , \new_[16632]_ , \new_[16633]_ , \new_[16634]_ ,
    \new_[16635]_ , \new_[16636]_ , \new_[16637]_ , \new_[16638]_ ,
    \new_[16639]_ , \new_[16640]_ , \new_[16641]_ , \new_[16642]_ ,
    \new_[16644]_ , \new_[16645]_ , \new_[16646]_ , \new_[16647]_ ,
    \new_[16648]_ , \new_[16649]_ , \new_[16650]_ , \new_[16654]_ ,
    \new_[16655]_ , \new_[16657]_ , \new_[16658]_ , \new_[16659]_ ,
    \new_[16660]_ , \new_[16661]_ , \new_[16662]_ , \new_[16663]_ ,
    \new_[16664]_ , \new_[16665]_ , \new_[16666]_ , \new_[16668]_ ,
    \new_[16669]_ , \new_[16670]_ , \new_[16671]_ , \new_[16672]_ ,
    \new_[16673]_ , \new_[16674]_ , \new_[16676]_ , \new_[16677]_ ,
    \new_[16678]_ , \new_[16679]_ , \new_[16680]_ , \new_[16681]_ ,
    \new_[16682]_ , \new_[16683]_ , \new_[16684]_ , \new_[16685]_ ,
    \new_[16686]_ , \new_[16687]_ , \new_[16691]_ , \new_[16692]_ ,
    \new_[16693]_ , \new_[16694]_ , \new_[16695]_ , \new_[16696]_ ,
    \new_[16697]_ , \new_[16699]_ , \new_[16700]_ , \new_[16701]_ ,
    \new_[16702]_ , \new_[16703]_ , \new_[16704]_ , \new_[16705]_ ,
    \new_[16706]_ , \new_[16708]_ , \new_[16709]_ , \new_[16710]_ ,
    \new_[16711]_ , \new_[16712]_ , \new_[16713]_ , \new_[16714]_ ,
    \new_[16715]_ , \new_[16716]_ , \new_[16717]_ , \new_[16718]_ ,
    \new_[16719]_ , \new_[16720]_ , \new_[16721]_ , \new_[16722]_ ,
    \new_[16723]_ , \new_[16724]_ , \new_[16725]_ , \new_[16726]_ ,
    \new_[16727]_ , \new_[16728]_ , \new_[16729]_ , \new_[16730]_ ,
    \new_[16731]_ , \new_[16732]_ , \new_[16734]_ , \new_[16735]_ ,
    \new_[16736]_ , \new_[16737]_ , \new_[16738]_ , \new_[16739]_ ,
    \new_[16740]_ , \new_[16741]_ , \new_[16742]_ , \new_[16743]_ ,
    \new_[16744]_ , \new_[16745]_ , \new_[16746]_ , \new_[16747]_ ,
    \new_[16748]_ , \new_[16749]_ , \new_[16750]_ , \new_[16751]_ ,
    \new_[16752]_ , \new_[16753]_ , \new_[16754]_ , \new_[16755]_ ,
    \new_[16756]_ , \new_[16757]_ , \new_[16758]_ , \new_[16759]_ ,
    \new_[16760]_ , \new_[16761]_ , \new_[16762]_ , \new_[16763]_ ,
    \new_[16764]_ , \new_[16765]_ , \new_[16766]_ , \new_[16767]_ ,
    \new_[16768]_ , \new_[16769]_ , \new_[16770]_ , \new_[16771]_ ,
    \new_[16772]_ , \new_[16773]_ , \new_[16774]_ , \new_[16775]_ ,
    \new_[16776]_ , \new_[16777]_ , \new_[16778]_ , \new_[16779]_ ,
    \new_[16780]_ , \new_[16781]_ , \new_[16782]_ , \new_[16783]_ ,
    \new_[16784]_ , \new_[16785]_ , \new_[16786]_ , \new_[16787]_ ,
    \new_[16788]_ , \new_[16789]_ , \new_[16790]_ , \new_[16791]_ ,
    \new_[16792]_ , \new_[16793]_ , \new_[16794]_ , \new_[16795]_ ,
    \new_[16796]_ , \new_[16797]_ , \new_[16798]_ , \new_[16799]_ ,
    \new_[16800]_ , \new_[16801]_ , \new_[16802]_ , \new_[16803]_ ,
    \new_[16804]_ , \new_[16805]_ , \new_[16806]_ , \new_[16807]_ ,
    \new_[16808]_ , \new_[16809]_ , \new_[16810]_ , \new_[16811]_ ,
    \new_[16816]_ , \new_[16818]_ , \new_[16819]_ , \new_[16820]_ ,
    \new_[16821]_ , \new_[16822]_ , \new_[16823]_ , \new_[16824]_ ,
    \new_[16825]_ , \new_[16826]_ , \new_[16827]_ , \new_[16828]_ ,
    \new_[16829]_ , \new_[16830]_ , \new_[16831]_ , \new_[16832]_ ,
    \new_[16833]_ , \new_[16834]_ , \new_[16835]_ , \new_[16836]_ ,
    \new_[16837]_ , \new_[16838]_ , \new_[16839]_ , \new_[16840]_ ,
    \new_[16841]_ , \new_[16842]_ , \new_[16843]_ , \new_[16844]_ ,
    \new_[16845]_ , \new_[16846]_ , \new_[16847]_ , \new_[16848]_ ,
    \new_[16849]_ , \new_[16850]_ , \new_[16851]_ , \new_[16852]_ ,
    \new_[16853]_ , \new_[16855]_ , \new_[16857]_ , \new_[16858]_ ,
    \new_[16859]_ , \new_[16860]_ , \new_[16861]_ , \new_[16863]_ ,
    \new_[16864]_ , \new_[16865]_ , \new_[16866]_ , \new_[16867]_ ,
    \new_[16868]_ , \new_[16869]_ , \new_[16870]_ , \new_[16871]_ ,
    \new_[16873]_ , \new_[16874]_ , \new_[16875]_ , \new_[16876]_ ,
    \new_[16877]_ , \new_[16878]_ , \new_[16879]_ , \new_[16880]_ ,
    \new_[16881]_ , \new_[16882]_ , \new_[16883]_ , \new_[16884]_ ,
    \new_[16885]_ , \new_[16886]_ , \new_[16887]_ , \new_[16888]_ ,
    \new_[16889]_ , \new_[16890]_ , \new_[16891]_ , \new_[16892]_ ,
    \new_[16893]_ , \new_[16894]_ , \new_[16895]_ , \new_[16896]_ ,
    \new_[16897]_ , \new_[16898]_ , \new_[16899]_ , \new_[16900]_ ,
    \new_[16901]_ , \new_[16903]_ , \new_[16904]_ , \new_[16905]_ ,
    \new_[16906]_ , \new_[16907]_ , \new_[16908]_ , \new_[16909]_ ,
    \new_[16910]_ , \new_[16911]_ , \new_[16912]_ , \new_[16913]_ ,
    \new_[16914]_ , \new_[16915]_ , \new_[16916]_ , \new_[16917]_ ,
    \new_[16918]_ , \new_[16919]_ , \new_[16920]_ , \new_[16921]_ ,
    \new_[16922]_ , \new_[16923]_ , \new_[16924]_ , \new_[16925]_ ,
    \new_[16926]_ , \new_[16927]_ , \new_[16928]_ , \new_[16929]_ ,
    \new_[16930]_ , \new_[16931]_ , \new_[16932]_ , \new_[16933]_ ,
    \new_[16934]_ , \new_[16935]_ , \new_[16936]_ , \new_[16937]_ ,
    \new_[16938]_ , \new_[16939]_ , \new_[16940]_ , \new_[16941]_ ,
    \new_[16942]_ , \new_[16943]_ , \new_[16944]_ , \new_[16945]_ ,
    \new_[16946]_ , \new_[16947]_ , \new_[16948]_ , \new_[16949]_ ,
    \new_[16950]_ , \new_[16951]_ , \new_[16954]_ , \new_[16955]_ ,
    \new_[16956]_ , \new_[16958]_ , \new_[16959]_ , \new_[16960]_ ,
    \new_[16961]_ , \new_[16962]_ , \new_[16963]_ , \new_[16964]_ ,
    \new_[16965]_ , \new_[16966]_ , \new_[16967]_ , \new_[16968]_ ,
    \new_[16969]_ , \new_[16970]_ , \new_[16971]_ , \new_[16972]_ ,
    \new_[16973]_ , \new_[16974]_ , \new_[16975]_ , \new_[16976]_ ,
    \new_[16977]_ , \new_[16978]_ , \new_[16979]_ , \new_[16980]_ ,
    \new_[16981]_ , \new_[16982]_ , \new_[16983]_ , \new_[16984]_ ,
    \new_[16985]_ , \new_[16986]_ , \new_[16987]_ , \new_[16988]_ ,
    \new_[16989]_ , \new_[16990]_ , \new_[16991]_ , \new_[16992]_ ,
    \new_[16993]_ , \new_[16994]_ , \new_[16995]_ , \new_[16996]_ ,
    \new_[16997]_ , \new_[16998]_ , \new_[16999]_ , \new_[17000]_ ,
    \new_[17001]_ , \new_[17002]_ , \new_[17003]_ , \new_[17004]_ ,
    \new_[17005]_ , \new_[17006]_ , \new_[17007]_ , \new_[17008]_ ,
    \new_[17009]_ , \new_[17011]_ , \new_[17012]_ , \new_[17013]_ ,
    \new_[17014]_ , \new_[17015]_ , \new_[17016]_ , \new_[17017]_ ,
    \new_[17018]_ , \new_[17019]_ , \new_[17020]_ , \new_[17021]_ ,
    \new_[17022]_ , \new_[17023]_ , \new_[17024]_ , \new_[17025]_ ,
    \new_[17026]_ , \new_[17027]_ , \new_[17028]_ , \new_[17029]_ ,
    \new_[17030]_ , \new_[17031]_ , \new_[17032]_ , \new_[17033]_ ,
    \new_[17034]_ , \new_[17035]_ , \new_[17036]_ , \new_[17037]_ ,
    \new_[17038]_ , \new_[17039]_ , \new_[17040]_ , \new_[17041]_ ,
    \new_[17042]_ , \new_[17043]_ , \new_[17044]_ , \new_[17045]_ ,
    \new_[17046]_ , \new_[17047]_ , \new_[17048]_ , \new_[17049]_ ,
    \new_[17050]_ , \new_[17051]_ , \new_[17052]_ , \new_[17053]_ ,
    \new_[17054]_ , \new_[17055]_ , \new_[17056]_ , \new_[17057]_ ,
    \new_[17058]_ , \new_[17059]_ , \new_[17060]_ , \new_[17061]_ ,
    \new_[17062]_ , \new_[17063]_ , \new_[17064]_ , \new_[17065]_ ,
    \new_[17066]_ , \new_[17067]_ , \new_[17068]_ , \new_[17070]_ ,
    \new_[17072]_ , \new_[17073]_ , \new_[17074]_ , \new_[17075]_ ,
    \new_[17076]_ , \new_[17077]_ , \new_[17078]_ , \new_[17080]_ ,
    \new_[17081]_ , \new_[17082]_ , \new_[17083]_ , \new_[17084]_ ,
    \new_[17086]_ , \new_[17087]_ , \new_[17089]_ , \new_[17090]_ ,
    \new_[17091]_ , \new_[17092]_ , \new_[17093]_ , \new_[17094]_ ,
    \new_[17095]_ , \new_[17096]_ , \new_[17097]_ , \new_[17098]_ ,
    \new_[17099]_ , \new_[17100]_ , \new_[17101]_ , \new_[17102]_ ,
    \new_[17103]_ , \new_[17104]_ , \new_[17105]_ , \new_[17106]_ ,
    \new_[17107]_ , \new_[17108]_ , \new_[17109]_ , \new_[17110]_ ,
    \new_[17111]_ , \new_[17112]_ , \new_[17113]_ , \new_[17114]_ ,
    \new_[17115]_ , \new_[17116]_ , \new_[17117]_ , \new_[17118]_ ,
    \new_[17119]_ , \new_[17120]_ , \new_[17121]_ , \new_[17122]_ ,
    \new_[17123]_ , \new_[17124]_ , \new_[17125]_ , \new_[17126]_ ,
    \new_[17127]_ , \new_[17128]_ , \new_[17129]_ , \new_[17130]_ ,
    \new_[17131]_ , \new_[17132]_ , \new_[17133]_ , \new_[17134]_ ,
    \new_[17135]_ , \new_[17136]_ , \new_[17137]_ , \new_[17138]_ ,
    \new_[17139]_ , \new_[17140]_ , \new_[17141]_ , \new_[17142]_ ,
    \new_[17143]_ , \new_[17144]_ , \new_[17145]_ , \new_[17146]_ ,
    \new_[17147]_ , \new_[17148]_ , \new_[17149]_ , \new_[17150]_ ,
    \new_[17151]_ , \new_[17152]_ , \new_[17153]_ , \new_[17154]_ ,
    \new_[17155]_ , \new_[17156]_ , \new_[17157]_ , \new_[17158]_ ,
    \new_[17159]_ , \new_[17160]_ , \new_[17161]_ , \new_[17162]_ ,
    \new_[17163]_ , \new_[17164]_ , \new_[17165]_ , \new_[17166]_ ,
    \new_[17167]_ , \new_[17168]_ , \new_[17169]_ , \new_[17170]_ ,
    \new_[17171]_ , \new_[17172]_ , \new_[17173]_ , \new_[17174]_ ,
    \new_[17175]_ , \new_[17176]_ , \new_[17177]_ , \new_[17178]_ ,
    \new_[17179]_ , \new_[17180]_ , \new_[17181]_ , \new_[17182]_ ,
    \new_[17183]_ , \new_[17184]_ , \new_[17185]_ , \new_[17186]_ ,
    \new_[17187]_ , \new_[17188]_ , \new_[17189]_ , \new_[17190]_ ,
    \new_[17191]_ , \new_[17192]_ , \new_[17193]_ , \new_[17194]_ ,
    \new_[17195]_ , \new_[17196]_ , \new_[17197]_ , \new_[17198]_ ,
    \new_[17199]_ , \new_[17200]_ , \new_[17201]_ , \new_[17202]_ ,
    \new_[17203]_ , \new_[17204]_ , \new_[17205]_ , \new_[17206]_ ,
    \new_[17207]_ , \new_[17208]_ , \new_[17209]_ , \new_[17210]_ ,
    \new_[17211]_ , \new_[17212]_ , \new_[17213]_ , \new_[17214]_ ,
    \new_[17215]_ , \new_[17216]_ , \new_[17217]_ , \new_[17218]_ ,
    \new_[17219]_ , \new_[17220]_ , \new_[17221]_ , \new_[17222]_ ,
    \new_[17223]_ , \new_[17224]_ , \new_[17225]_ , \new_[17226]_ ,
    \new_[17227]_ , \new_[17228]_ , \new_[17229]_ , \new_[17230]_ ,
    \new_[17231]_ , \new_[17232]_ , \new_[17233]_ , \new_[17234]_ ,
    \new_[17235]_ , \new_[17236]_ , \new_[17237]_ , \new_[17238]_ ,
    \new_[17239]_ , \new_[17240]_ , \new_[17241]_ , \new_[17243]_ ,
    \new_[17244]_ , \new_[17247]_ , \new_[17249]_ , \new_[17250]_ ,
    \new_[17251]_ , \new_[17252]_ , \new_[17253]_ , \new_[17254]_ ,
    \new_[17255]_ , \new_[17256]_ , \new_[17257]_ , \new_[17258]_ ,
    \new_[17259]_ , \new_[17260]_ , \new_[17261]_ , \new_[17262]_ ,
    \new_[17263]_ , \new_[17264]_ , \new_[17265]_ , \new_[17266]_ ,
    \new_[17267]_ , \new_[17268]_ , \new_[17269]_ , \new_[17270]_ ,
    \new_[17271]_ , \new_[17272]_ , \new_[17273]_ , \new_[17274]_ ,
    \new_[17275]_ , \new_[17276]_ , \new_[17277]_ , \new_[17278]_ ,
    \new_[17279]_ , \new_[17280]_ , \new_[17281]_ , \new_[17282]_ ,
    \new_[17283]_ , \new_[17284]_ , \new_[17285]_ , \new_[17286]_ ,
    \new_[17288]_ , \new_[17290]_ , \new_[17291]_ , \new_[17292]_ ,
    \new_[17293]_ , \new_[17294]_ , \new_[17296]_ , \new_[17298]_ ,
    \new_[17299]_ , \new_[17300]_ , \new_[17301]_ , \new_[17302]_ ,
    \new_[17303]_ , \new_[17304]_ , \new_[17305]_ , \new_[17306]_ ,
    \new_[17307]_ , \new_[17308]_ , \new_[17309]_ , \new_[17310]_ ,
    \new_[17311]_ , \new_[17312]_ , \new_[17313]_ , \new_[17314]_ ,
    \new_[17317]_ , \new_[17318]_ , \new_[17319]_ , \new_[17323]_ ,
    \new_[17324]_ , \new_[17334]_ , \new_[17339]_ , \new_[17340]_ ,
    \new_[17341]_ , \new_[17342]_ , \new_[17343]_ , \new_[17344]_ ,
    \new_[17345]_ , \new_[17346]_ , \new_[17347]_ , \new_[17348]_ ,
    \new_[17349]_ , \new_[17350]_ , \new_[17351]_ , \new_[17352]_ ,
    \new_[17353]_ , \new_[17354]_ , \new_[17355]_ , \new_[17356]_ ,
    \new_[17357]_ , \new_[17358]_ , \new_[17359]_ , \new_[17360]_ ,
    \new_[17361]_ , \new_[17362]_ , \new_[17363]_ , \new_[17364]_ ,
    \new_[17365]_ , \new_[17366]_ , \new_[17367]_ , \new_[17368]_ ,
    \new_[17369]_ , \new_[17370]_ , \new_[17371]_ , \new_[17372]_ ,
    \new_[17374]_ , \new_[17375]_ , \new_[17377]_ , \new_[17378]_ ,
    \new_[17379]_ , \new_[17380]_ , \new_[17381]_ , \new_[17382]_ ,
    \new_[17383]_ , \new_[17384]_ , \new_[17385]_ , \new_[17386]_ ,
    \new_[17387]_ , \new_[17388]_ , \new_[17389]_ , \new_[17390]_ ,
    \new_[17391]_ , \new_[17392]_ , \new_[17393]_ , \new_[17394]_ ,
    \new_[17395]_ , \new_[17396]_ , \new_[17397]_ , \new_[17398]_ ,
    \new_[17399]_ , \new_[17400]_ , \new_[17401]_ , \new_[17402]_ ,
    \new_[17403]_ , \new_[17404]_ , \new_[17405]_ , \new_[17406]_ ,
    \new_[17407]_ , \new_[17408]_ , \new_[17409]_ , \new_[17410]_ ,
    \new_[17411]_ , \new_[17412]_ , \new_[17413]_ , \new_[17414]_ ,
    \new_[17415]_ , \new_[17416]_ , \new_[17417]_ , \new_[17418]_ ,
    \new_[17419]_ , \new_[17420]_ , \new_[17421]_ , \new_[17422]_ ,
    \new_[17423]_ , \new_[17424]_ , \new_[17425]_ , \new_[17426]_ ,
    \new_[17427]_ , \new_[17428]_ , \new_[17429]_ , \new_[17430]_ ,
    \new_[17431]_ , \new_[17433]_ , \new_[17434]_ , \new_[17435]_ ,
    \new_[17436]_ , \new_[17437]_ , \new_[17438]_ , \new_[17439]_ ,
    \new_[17440]_ , \new_[17441]_ , \new_[17442]_ , \new_[17443]_ ,
    \new_[17444]_ , \new_[17445]_ , \new_[17446]_ , \new_[17447]_ ,
    \new_[17448]_ , \new_[17449]_ , \new_[17450]_ , \new_[17451]_ ,
    \new_[17452]_ , \new_[17453]_ , \new_[17454]_ , \new_[17455]_ ,
    \new_[17456]_ , \new_[17457]_ , \new_[17459]_ , \new_[17460]_ ,
    \new_[17461]_ , \new_[17462]_ , \new_[17463]_ , \new_[17464]_ ,
    \new_[17465]_ , \new_[17466]_ , \new_[17467]_ , \new_[17468]_ ,
    \new_[17469]_ , \new_[17470]_ , \new_[17471]_ , \new_[17472]_ ,
    \new_[17473]_ , \new_[17474]_ , \new_[17475]_ , \new_[17476]_ ,
    \new_[17478]_ , \new_[17479]_ , \new_[17480]_ , \new_[17481]_ ,
    \new_[17482]_ , \new_[17483]_ , \new_[17484]_ , \new_[17485]_ ,
    \new_[17486]_ , \new_[17487]_ , \new_[17488]_ , \new_[17489]_ ,
    \new_[17490]_ , \new_[17491]_ , \new_[17492]_ , \new_[17493]_ ,
    \new_[17494]_ , \new_[17495]_ , \new_[17504]_ , \new_[17505]_ ,
    \new_[17506]_ , \new_[17507]_ , \new_[17508]_ , \new_[17509]_ ,
    \new_[17510]_ , \new_[17512]_ , \new_[17513]_ , \new_[17514]_ ,
    \new_[17515]_ , \new_[17516]_ , \new_[17517]_ , \new_[17518]_ ,
    \new_[17519]_ , \new_[17520]_ , \new_[17521]_ , \new_[17522]_ ,
    \new_[17523]_ , \new_[17524]_ , \new_[17525]_ , \new_[17526]_ ,
    \new_[17527]_ , \new_[17528]_ , \new_[17529]_ , \new_[17530]_ ,
    \new_[17531]_ , \new_[17532]_ , \new_[17533]_ , \new_[17535]_ ,
    \new_[17536]_ , \new_[17537]_ , \new_[17539]_ , \new_[17540]_ ,
    \new_[17541]_ , \new_[17542]_ , \new_[17543]_ , \new_[17544]_ ,
    \new_[17545]_ , \new_[17546]_ , \new_[17547]_ , \new_[17548]_ ,
    \new_[17549]_ , \new_[17550]_ , \new_[17551]_ , \new_[17553]_ ,
    \new_[17554]_ , \new_[17555]_ , \new_[17556]_ , \new_[17557]_ ,
    \new_[17558]_ , \new_[17560]_ , \new_[17561]_ , \new_[17562]_ ,
    \new_[17563]_ , \new_[17564]_ , \new_[17565]_ , \new_[17566]_ ,
    \new_[17567]_ , \new_[17568]_ , \new_[17569]_ , \new_[17570]_ ,
    \new_[17571]_ , \new_[17572]_ , \new_[17573]_ , \new_[17574]_ ,
    \new_[17575]_ , \new_[17576]_ , \new_[17577]_ , \new_[17578]_ ,
    \new_[17579]_ , \new_[17580]_ , \new_[17581]_ , \new_[17582]_ ,
    \new_[17583]_ , \new_[17584]_ , \new_[17585]_ , \new_[17587]_ ,
    \new_[17588]_ , \new_[17589]_ , \new_[17590]_ , \new_[17591]_ ,
    \new_[17592]_ , \new_[17593]_ , \new_[17594]_ , \new_[17597]_ ,
    \new_[17598]_ , \new_[17599]_ , \new_[17601]_ , \new_[17602]_ ,
    \new_[17603]_ , \new_[17604]_ , \new_[17605]_ , \new_[17606]_ ,
    \new_[17607]_ , \new_[17608]_ , \new_[17611]_ , \new_[17612]_ ,
    \new_[17613]_ , \new_[17620]_ , \new_[17622]_ , \new_[17627]_ ,
    \new_[17628]_ , \new_[17630]_ , \new_[17631]_ , \new_[17632]_ ,
    \new_[17633]_ , \new_[17635]_ , \new_[17636]_ , \new_[17637]_ ,
    \new_[17638]_ , \new_[17639]_ , \new_[17640]_ , \new_[17641]_ ,
    \new_[17642]_ , \new_[17645]_ , \new_[17646]_ , \new_[17648]_ ,
    \new_[17649]_ , \new_[17650]_ , \new_[17652]_ , \new_[17653]_ ,
    \new_[17654]_ , \new_[17655]_ , \new_[17656]_ , \new_[17659]_ ,
    \new_[17661]_ , \new_[17662]_ , \new_[17663]_ , \new_[17664]_ ,
    \new_[17665]_ , \new_[17666]_ , \new_[17667]_ , \new_[17668]_ ,
    \new_[17669]_ , \new_[17670]_ , \new_[17671]_ , \new_[17672]_ ,
    \new_[17673]_ , \new_[17674]_ , \new_[17675]_ , \new_[17676]_ ,
    \new_[17677]_ , \new_[17678]_ , \new_[17679]_ , \new_[17680]_ ,
    \new_[17681]_ , \new_[17682]_ , \new_[17683]_ , \new_[17684]_ ,
    \new_[17685]_ , \new_[17686]_ , \new_[17687]_ , \new_[17688]_ ,
    \new_[17690]_ , \new_[17691]_ , \new_[17692]_ , \new_[17694]_ ,
    \new_[17697]_ , \new_[17698]_ , \new_[17699]_ , \new_[17700]_ ,
    \new_[17702]_ , \new_[17703]_ , \new_[17704]_ , \new_[17705]_ ,
    \new_[17706]_ , \new_[17707]_ , \new_[17708]_ , \new_[17709]_ ,
    \new_[17712]_ , \new_[17713]_ , \new_[17714]_ , \new_[17715]_ ,
    \new_[17716]_ , \new_[17717]_ , \new_[17718]_ , \new_[17719]_ ,
    \new_[17721]_ , \new_[17722]_ , \new_[17723]_ , \new_[17726]_ ,
    \new_[17727]_ , \new_[17728]_ , \new_[17729]_ , \new_[17730]_ ,
    \new_[17731]_ , \new_[17732]_ , \new_[17733]_ , \new_[17734]_ ,
    \new_[17735]_ , \new_[17736]_ , \new_[17737]_ , \new_[17738]_ ,
    \new_[17739]_ , \new_[17740]_ , \new_[17741]_ , \new_[17742]_ ,
    \new_[17743]_ , \new_[17744]_ , \new_[17746]_ , \new_[17747]_ ,
    \new_[17748]_ , \new_[17749]_ , \new_[17750]_ , \new_[17751]_ ,
    \new_[17752]_ , \new_[17753]_ , \new_[17755]_ , \new_[17756]_ ,
    \new_[17758]_ , \new_[17759]_ , \new_[17760]_ , \new_[17761]_ ,
    \new_[17762]_ , \new_[17763]_ , \new_[17764]_ , \new_[17765]_ ,
    \new_[17766]_ , \new_[17767]_ , \new_[17768]_ , \new_[17769]_ ,
    \new_[17770]_ , \new_[17771]_ , \new_[17772]_ , \new_[17773]_ ,
    \new_[17774]_ , \new_[17775]_ , \new_[17776]_ , \new_[17777]_ ,
    \new_[17778]_ , \new_[17779]_ , \new_[17780]_ , \new_[17781]_ ,
    \new_[17782]_ , \new_[17783]_ , \new_[17784]_ , \new_[17785]_ ,
    \new_[17786]_ , \new_[17787]_ , \new_[17788]_ , \new_[17789]_ ,
    \new_[17791]_ , \new_[17792]_ , \new_[17793]_ , \new_[17794]_ ,
    \new_[17795]_ , \new_[17797]_ , \new_[17798]_ , \new_[17799]_ ,
    \new_[17800]_ , \new_[17801]_ , \new_[17802]_ , \new_[17803]_ ,
    \new_[17805]_ , \new_[17806]_ , \new_[17807]_ , \new_[17808]_ ,
    \new_[17809]_ , \new_[17810]_ , \new_[17811]_ , \new_[17812]_ ,
    \new_[17813]_ , \new_[17814]_ , \new_[17815]_ , \new_[17816]_ ,
    \new_[17817]_ , \new_[17818]_ , \new_[17819]_ , \new_[17820]_ ,
    \new_[17821]_ , \new_[17822]_ , \new_[17823]_ , \new_[17824]_ ,
    \new_[17825]_ , \new_[17826]_ , \new_[17827]_ , \new_[17828]_ ,
    \new_[17829]_ , \new_[17831]_ , \new_[17832]_ , \new_[17833]_ ,
    \new_[17834]_ , \new_[17835]_ , \new_[17836]_ , \new_[17837]_ ,
    \new_[17838]_ , \new_[17839]_ , \new_[17840]_ , \new_[17841]_ ,
    \new_[17842]_ , \new_[17843]_ , \new_[17844]_ , \new_[17845]_ ,
    \new_[17846]_ , \new_[17847]_ , \new_[17848]_ , \new_[17849]_ ,
    \new_[17850]_ , \new_[17851]_ , \new_[17852]_ , \new_[17853]_ ,
    \new_[17854]_ , \new_[17855]_ , \new_[17856]_ , \new_[17857]_ ,
    \new_[17858]_ , \new_[17859]_ , \new_[17860]_ , \new_[17861]_ ,
    \new_[17862]_ , \new_[17863]_ , \new_[17864]_ , \new_[17865]_ ,
    \new_[17866]_ , \new_[17867]_ , \new_[17868]_ , \new_[17869]_ ,
    \new_[17870]_ , \new_[17871]_ , \new_[17872]_ , \new_[17873]_ ,
    \new_[17874]_ , \new_[17875]_ , \new_[17876]_ , \new_[17877]_ ,
    \new_[17878]_ , \new_[17879]_ , \new_[17880]_ , \new_[17881]_ ,
    \new_[17882]_ , \new_[17883]_ , \new_[17884]_ , \new_[17885]_ ,
    \new_[17886]_ , \new_[17887]_ , \new_[17888]_ , \new_[17889]_ ,
    \new_[17890]_ , \new_[17891]_ , \new_[17892]_ , \new_[17893]_ ,
    \new_[17894]_ , \new_[17895]_ , \new_[17896]_ , \new_[17897]_ ,
    \new_[17898]_ , \new_[17899]_ , \new_[17900]_ , \new_[17901]_ ,
    \new_[17902]_ , \new_[17903]_ , \new_[17904]_ , \new_[17905]_ ,
    \new_[17906]_ , \new_[17907]_ , \new_[17908]_ , \new_[17909]_ ,
    \new_[17910]_ , \new_[17911]_ , \new_[17912]_ , \new_[17913]_ ,
    \new_[17914]_ , \new_[17915]_ , \new_[17916]_ , \new_[17917]_ ,
    \new_[17918]_ , \new_[17919]_ , \new_[17920]_ , \new_[17921]_ ,
    \new_[17922]_ , \new_[17923]_ , \new_[17924]_ , \new_[17925]_ ,
    \new_[17926]_ , \new_[17927]_ , \new_[17928]_ , \new_[17929]_ ,
    \new_[17930]_ , \new_[17931]_ , \new_[17932]_ , \new_[17933]_ ,
    \new_[17934]_ , \new_[17935]_ , \new_[17936]_ , \new_[17937]_ ,
    \new_[17938]_ , \new_[17939]_ , \new_[17940]_ , \new_[17941]_ ,
    \new_[17942]_ , \new_[17943]_ , \new_[17944]_ , \new_[17945]_ ,
    \new_[17946]_ , \new_[17947]_ , \new_[17948]_ , \new_[17949]_ ,
    \new_[17950]_ , \new_[17951]_ , \new_[17952]_ , \new_[17953]_ ,
    \new_[17954]_ , \new_[17955]_ , \new_[17956]_ , \new_[17957]_ ,
    \new_[17958]_ , \new_[17959]_ , \new_[17960]_ , \new_[17961]_ ,
    \new_[17962]_ , \new_[17963]_ , \new_[17964]_ , \new_[17965]_ ,
    \new_[17966]_ , \new_[17967]_ , \new_[17968]_ , \new_[17969]_ ,
    \new_[17970]_ , \new_[17971]_ , \new_[17972]_ , \new_[17973]_ ,
    \new_[17974]_ , \new_[17975]_ , \new_[17976]_ , \new_[17977]_ ,
    \new_[17978]_ , \new_[17979]_ , \new_[17980]_ , \new_[17981]_ ,
    \new_[17982]_ , \new_[17983]_ , \new_[17984]_ , \new_[17985]_ ,
    \new_[17986]_ , \new_[17987]_ , \new_[17988]_ , \new_[17989]_ ,
    \new_[17990]_ , \new_[17991]_ , \new_[17992]_ , \new_[17993]_ ,
    \new_[17994]_ , \new_[17995]_ , \new_[17996]_ , \new_[17997]_ ,
    \new_[17998]_ , \new_[17999]_ , \new_[18000]_ , \new_[18001]_ ,
    \new_[18002]_ , \new_[18003]_ , \new_[18004]_ , \new_[18005]_ ,
    \new_[18006]_ , \new_[18007]_ , \new_[18008]_ , \new_[18009]_ ,
    \new_[18010]_ , \new_[18011]_ , \new_[18012]_ , \new_[18013]_ ,
    \new_[18014]_ , \new_[18015]_ , \new_[18016]_ , \new_[18017]_ ,
    \new_[18018]_ , \new_[18019]_ , \new_[18020]_ , \new_[18021]_ ,
    \new_[18022]_ , \new_[18023]_ , \new_[18024]_ , \new_[18025]_ ,
    \new_[18026]_ , \new_[18027]_ , \new_[18028]_ , \new_[18029]_ ,
    \new_[18030]_ , \new_[18031]_ , \new_[18032]_ , \new_[18033]_ ,
    \new_[18034]_ , \new_[18035]_ , \new_[18036]_ , \new_[18037]_ ,
    \new_[18038]_ , \new_[18039]_ , \new_[18040]_ , \new_[18041]_ ,
    \new_[18042]_ , \new_[18043]_ , \new_[18044]_ , \new_[18045]_ ,
    \new_[18046]_ , \new_[18047]_ , \new_[18048]_ , \new_[18049]_ ,
    \new_[18050]_ , \new_[18051]_ , \new_[18052]_ , \new_[18053]_ ,
    \new_[18054]_ , \new_[18055]_ , \new_[18056]_ , \new_[18057]_ ,
    \new_[18058]_ , \new_[18059]_ , \new_[18060]_ , \new_[18061]_ ,
    \new_[18062]_ , \new_[18063]_ , \new_[18064]_ , \new_[18066]_ ,
    \new_[18067]_ , \new_[18068]_ , \new_[18069]_ , \new_[18070]_ ,
    \new_[18071]_ , \new_[18072]_ , \new_[18073]_ , \new_[18074]_ ,
    \new_[18075]_ , \new_[18076]_ , \new_[18077]_ , \new_[18078]_ ,
    \new_[18079]_ , \new_[18080]_ , \new_[18081]_ , \new_[18082]_ ,
    \new_[18083]_ , \new_[18084]_ , \new_[18085]_ , \new_[18086]_ ,
    \new_[18087]_ , \new_[18088]_ , \new_[18089]_ , \new_[18090]_ ,
    \new_[18091]_ , \new_[18092]_ , \new_[18093]_ , \new_[18094]_ ,
    \new_[18095]_ , \new_[18096]_ , \new_[18097]_ , \new_[18098]_ ,
    \new_[18099]_ , \new_[18100]_ , \new_[18101]_ , \new_[18102]_ ,
    \new_[18103]_ , \new_[18104]_ , \new_[18105]_ , \new_[18106]_ ,
    \new_[18107]_ , \new_[18108]_ , \new_[18109]_ , \new_[18110]_ ,
    \new_[18111]_ , \new_[18112]_ , \new_[18113]_ , \new_[18114]_ ,
    \new_[18115]_ , \new_[18116]_ , \new_[18117]_ , \new_[18118]_ ,
    \new_[18120]_ , \new_[18121]_ , \new_[18122]_ , \new_[18123]_ ,
    \new_[18124]_ , \new_[18125]_ , \new_[18126]_ , \new_[18127]_ ,
    \new_[18128]_ , \new_[18129]_ , \new_[18130]_ , \new_[18131]_ ,
    \new_[18132]_ , \new_[18135]_ , \new_[18136]_ , \new_[18137]_ ,
    \new_[18138]_ , \new_[18139]_ , \new_[18140]_ , \new_[18141]_ ,
    \new_[18142]_ , \new_[18143]_ , \new_[18144]_ , \new_[18145]_ ,
    \new_[18146]_ , \new_[18147]_ , \new_[18148]_ , \new_[18149]_ ,
    \new_[18150]_ , \new_[18151]_ , \new_[18152]_ , \new_[18153]_ ,
    \new_[18154]_ , \new_[18155]_ , \new_[18156]_ , \new_[18157]_ ,
    \new_[18158]_ , \new_[18159]_ , \new_[18160]_ , \new_[18161]_ ,
    \new_[18162]_ , \new_[18163]_ , \new_[18164]_ , \new_[18165]_ ,
    \new_[18166]_ , \new_[18167]_ , \new_[18168]_ , \new_[18169]_ ,
    \new_[18170]_ , \new_[18171]_ , \new_[18172]_ , \new_[18173]_ ,
    \new_[18174]_ , \new_[18175]_ , \new_[18176]_ , \new_[18177]_ ,
    \new_[18178]_ , \new_[18179]_ , \new_[18180]_ , \new_[18181]_ ,
    \new_[18182]_ , \new_[18183]_ , \new_[18184]_ , \new_[18185]_ ,
    \new_[18186]_ , \new_[18187]_ , \new_[18188]_ , \new_[18189]_ ,
    \new_[18190]_ , \new_[18191]_ , \new_[18192]_ , \new_[18193]_ ,
    \new_[18194]_ , \new_[18195]_ , \new_[18196]_ , \new_[18197]_ ,
    \new_[18198]_ , \new_[18199]_ , \new_[18200]_ , \new_[18201]_ ,
    \new_[18202]_ , \new_[18203]_ , \new_[18204]_ , \new_[18205]_ ,
    \new_[18206]_ , \new_[18207]_ , \new_[18208]_ , \new_[18209]_ ,
    \new_[18210]_ , \new_[18211]_ , \new_[18212]_ , \new_[18213]_ ,
    \new_[18214]_ , \new_[18215]_ , \new_[18216]_ , \new_[18217]_ ,
    \new_[18218]_ , \new_[18219]_ , \new_[18220]_ , \new_[18221]_ ,
    \new_[18222]_ , \new_[18223]_ , \new_[18224]_ , \new_[18225]_ ,
    \new_[18226]_ , \new_[18227]_ , \new_[18228]_ , \new_[18229]_ ,
    \new_[18230]_ , \new_[18231]_ , \new_[18232]_ , \new_[18233]_ ,
    \new_[18234]_ , \new_[18235]_ , \new_[18236]_ , \new_[18237]_ ,
    \new_[18238]_ , \new_[18239]_ , \new_[18240]_ , \new_[18241]_ ,
    \new_[18242]_ , \new_[18243]_ , \new_[18244]_ , \new_[18245]_ ,
    \new_[18246]_ , \new_[18247]_ , \new_[18248]_ , \new_[18249]_ ,
    \new_[18250]_ , \new_[18251]_ , \new_[18252]_ , \new_[18253]_ ,
    \new_[18255]_ , \new_[18256]_ , \new_[18257]_ , \new_[18258]_ ,
    \new_[18259]_ , \new_[18260]_ , \new_[18261]_ , \new_[18262]_ ,
    \new_[18263]_ , \new_[18264]_ , \new_[18265]_ , \new_[18266]_ ,
    \new_[18267]_ , \new_[18268]_ , \new_[18269]_ , \new_[18270]_ ,
    \new_[18271]_ , \new_[18272]_ , \new_[18273]_ , \new_[18274]_ ,
    \new_[18275]_ , \new_[18276]_ , \new_[18277]_ , \new_[18278]_ ,
    \new_[18279]_ , \new_[18280]_ , \new_[18281]_ , \new_[18282]_ ,
    \new_[18283]_ , \new_[18284]_ , \new_[18285]_ , \new_[18286]_ ,
    \new_[18287]_ , \new_[18288]_ , \new_[18289]_ , \new_[18290]_ ,
    \new_[18291]_ , \new_[18292]_ , \new_[18293]_ , \new_[18294]_ ,
    \new_[18295]_ , \new_[18296]_ , \new_[18297]_ , \new_[18299]_ ,
    \new_[18300]_ , \new_[18301]_ , \new_[18302]_ , \new_[18303]_ ,
    \new_[18304]_ , \new_[18305]_ , \new_[18306]_ , \new_[18307]_ ,
    \new_[18308]_ , \new_[18309]_ , \new_[18310]_ , \new_[18311]_ ,
    \new_[18312]_ , \new_[18313]_ , \new_[18314]_ , \new_[18315]_ ,
    \new_[18316]_ , \new_[18317]_ , \new_[18318]_ , \new_[18319]_ ,
    \new_[18320]_ , \new_[18321]_ , \new_[18322]_ , \new_[18323]_ ,
    \new_[18324]_ , \new_[18325]_ , \new_[18326]_ , \new_[18327]_ ,
    \new_[18329]_ , \new_[18330]_ , \new_[18331]_ , \new_[18332]_ ,
    \new_[18333]_ , \new_[18334]_ , \new_[18335]_ , \new_[18336]_ ,
    \new_[18337]_ , \new_[18338]_ , \new_[18339]_ , \new_[18340]_ ,
    \new_[18341]_ , \new_[18342]_ , \new_[18343]_ , \new_[18344]_ ,
    \new_[18345]_ , \new_[18346]_ , \new_[18347]_ , \new_[18348]_ ,
    \new_[18349]_ , \new_[18350]_ , \new_[18351]_ , \new_[18352]_ ,
    \new_[18353]_ , \new_[18354]_ , \new_[18355]_ , \new_[18356]_ ,
    \new_[18357]_ , \new_[18358]_ , \new_[18359]_ , \new_[18360]_ ,
    \new_[18361]_ , \new_[18362]_ , \new_[18363]_ , \new_[18364]_ ,
    \new_[18365]_ , \new_[18366]_ , \new_[18367]_ , \new_[18368]_ ,
    \new_[18369]_ , \new_[18370]_ , \new_[18371]_ , \new_[18372]_ ,
    \new_[18373]_ , \new_[18374]_ , \new_[18375]_ , \new_[18376]_ ,
    \new_[18377]_ , \new_[18378]_ , \new_[18379]_ , \new_[18380]_ ,
    \new_[18381]_ , \new_[18382]_ , \new_[18383]_ , \new_[18384]_ ,
    \new_[18385]_ , \new_[18386]_ , \new_[18387]_ , \new_[18388]_ ,
    \new_[18389]_ , \new_[18390]_ , \new_[18391]_ , \new_[18392]_ ,
    \new_[18393]_ , \new_[18394]_ , \new_[18395]_ , \new_[18396]_ ,
    \new_[18397]_ , \new_[18398]_ , \new_[18399]_ , \new_[18400]_ ,
    \new_[18401]_ , \new_[18402]_ , \new_[18403]_ , \new_[18404]_ ,
    \new_[18405]_ , \new_[18406]_ , \new_[18407]_ , \new_[18408]_ ,
    \new_[18409]_ , \new_[18410]_ , \new_[18411]_ , \new_[18412]_ ,
    \new_[18413]_ , \new_[18414]_ , \new_[18415]_ , \new_[18416]_ ,
    \new_[18417]_ , \new_[18418]_ , \new_[18419]_ , \new_[18420]_ ,
    \new_[18421]_ , \new_[18422]_ , \new_[18423]_ , \new_[18424]_ ,
    \new_[18425]_ , \new_[18426]_ , \new_[18427]_ , \new_[18428]_ ,
    \new_[18429]_ , \new_[18430]_ , \new_[18431]_ , \new_[18432]_ ,
    \new_[18433]_ , \new_[18434]_ , \new_[18435]_ , \new_[18436]_ ,
    \new_[18437]_ , \new_[18438]_ , \new_[18439]_ , \new_[18440]_ ,
    \new_[18441]_ , \new_[18442]_ , \new_[18443]_ , \new_[18444]_ ,
    \new_[18445]_ , \new_[18446]_ , \new_[18447]_ , \new_[18448]_ ,
    \new_[18449]_ , \new_[18450]_ , \new_[18451]_ , \new_[18452]_ ,
    \new_[18453]_ , \new_[18454]_ , \new_[18455]_ , \new_[18456]_ ,
    \new_[18457]_ , \new_[18458]_ , \new_[18459]_ , \new_[18460]_ ,
    \new_[18461]_ , \new_[18462]_ , \new_[18463]_ , \new_[18464]_ ,
    \new_[18465]_ , \new_[18466]_ , \new_[18467]_ , \new_[18468]_ ,
    \new_[18469]_ , \new_[18470]_ , \new_[18472]_ , \new_[18473]_ ,
    \new_[18474]_ , \new_[18475]_ , \new_[18476]_ , \new_[18477]_ ,
    \new_[18478]_ , \new_[18479]_ , \new_[18480]_ , \new_[18481]_ ,
    \new_[18482]_ , \new_[18483]_ , \new_[18484]_ , \new_[18485]_ ,
    \new_[18486]_ , \new_[18487]_ , \new_[18488]_ , \new_[18489]_ ,
    \new_[18490]_ , \new_[18491]_ , \new_[18492]_ , \new_[18493]_ ,
    \new_[18494]_ , \new_[18495]_ , \new_[18496]_ , \new_[18497]_ ,
    \new_[18498]_ , \new_[18499]_ , \new_[18500]_ , \new_[18501]_ ,
    \new_[18502]_ , \new_[18503]_ , \new_[18504]_ , \new_[18505]_ ,
    \new_[18506]_ , \new_[18507]_ , \new_[18508]_ , \new_[18509]_ ,
    \new_[18510]_ , \new_[18511]_ , \new_[18512]_ , \new_[18513]_ ,
    \new_[18514]_ , \new_[18515]_ , \new_[18516]_ , \new_[18517]_ ,
    \new_[18518]_ , \new_[18519]_ , \new_[18520]_ , \new_[18521]_ ,
    \new_[18522]_ , \new_[18523]_ , \new_[18524]_ , \new_[18525]_ ,
    \new_[18526]_ , \new_[18527]_ , \new_[18528]_ , \new_[18529]_ ,
    \new_[18530]_ , \new_[18531]_ , \new_[18532]_ , \new_[18533]_ ,
    \new_[18534]_ , \new_[18535]_ , \new_[18536]_ , \new_[18537]_ ,
    \new_[18538]_ , \new_[18539]_ , \new_[18540]_ , \new_[18541]_ ,
    \new_[18542]_ , \new_[18543]_ , \new_[18544]_ , \new_[18545]_ ,
    \new_[18546]_ , \new_[18547]_ , \new_[18548]_ , \new_[18549]_ ,
    \new_[18550]_ , \new_[18551]_ , \new_[18552]_ , \new_[18553]_ ,
    \new_[18554]_ , \new_[18555]_ , \new_[18556]_ , \new_[18557]_ ,
    \new_[18558]_ , \new_[18559]_ , \new_[18560]_ , \new_[18561]_ ,
    \new_[18562]_ , \new_[18563]_ , \new_[18564]_ , \new_[18565]_ ,
    \new_[18566]_ , \new_[18567]_ , \new_[18568]_ , \new_[18569]_ ,
    \new_[18570]_ , \new_[18571]_ , \new_[18572]_ , \new_[18573]_ ,
    \new_[18574]_ , \new_[18575]_ , \new_[18576]_ , \new_[18577]_ ,
    \new_[18578]_ , \new_[18579]_ , \new_[18580]_ , \new_[18581]_ ,
    \new_[18582]_ , \new_[18583]_ , \new_[18584]_ , \new_[18585]_ ,
    \new_[18586]_ , \new_[18587]_ , \new_[18588]_ , \new_[18589]_ ,
    \new_[18590]_ , \new_[18591]_ , \new_[18592]_ , \new_[18593]_ ,
    \new_[18594]_ , \new_[18595]_ , \new_[18596]_ , \new_[18597]_ ,
    \new_[18598]_ , \new_[18599]_ , \new_[18600]_ , \new_[18601]_ ,
    \new_[18602]_ , \new_[18603]_ , \new_[18604]_ , \new_[18605]_ ,
    \new_[18606]_ , \new_[18607]_ , \new_[18608]_ , \new_[18609]_ ,
    \new_[18610]_ , \new_[18611]_ , \new_[18612]_ , \new_[18613]_ ,
    \new_[18614]_ , \new_[18615]_ , \new_[18616]_ , \new_[18617]_ ,
    \new_[18618]_ , \new_[18619]_ , \new_[18620]_ , \new_[18621]_ ,
    \new_[18622]_ , \new_[18623]_ , \new_[18624]_ , \new_[18625]_ ,
    \new_[18626]_ , \new_[18627]_ , \new_[18628]_ , \new_[18629]_ ,
    \new_[18630]_ , \new_[18631]_ , \new_[18632]_ , \new_[18633]_ ,
    \new_[18634]_ , \new_[18635]_ , \new_[18636]_ , \new_[18637]_ ,
    \new_[18638]_ , \new_[18639]_ , \new_[18640]_ , \new_[18641]_ ,
    \new_[18642]_ , \new_[18643]_ , \new_[18644]_ , \new_[18645]_ ,
    \new_[18646]_ , \new_[18647]_ , \new_[18648]_ , \new_[18649]_ ,
    \new_[18650]_ , \new_[18651]_ , \new_[18652]_ , \new_[18653]_ ,
    \new_[18654]_ , \new_[18655]_ , \new_[18656]_ , \new_[18657]_ ,
    \new_[18658]_ , \new_[18659]_ , \new_[18660]_ , \new_[18661]_ ,
    \new_[18662]_ , \new_[18663]_ , \new_[18664]_ , \new_[18665]_ ,
    \new_[18666]_ , \new_[18667]_ , \new_[18668]_ , \new_[18669]_ ,
    \new_[18670]_ , \new_[18672]_ , \new_[18673]_ , \new_[18674]_ ,
    \new_[18675]_ , \new_[18676]_ , \new_[18677]_ , \new_[18678]_ ,
    \new_[18679]_ , \new_[18680]_ , \new_[18681]_ , \new_[18682]_ ,
    \new_[18683]_ , \new_[18684]_ , \new_[18685]_ , \new_[18686]_ ,
    \new_[18687]_ , \new_[18688]_ , \new_[18689]_ , \new_[18690]_ ,
    \new_[18691]_ , \new_[18692]_ , \new_[18693]_ , \new_[18694]_ ,
    \new_[18695]_ , \new_[18696]_ , \new_[18697]_ , \new_[18698]_ ,
    \new_[18699]_ , \new_[18700]_ , \new_[18701]_ , \new_[18702]_ ,
    \new_[18703]_ , \new_[18704]_ , \new_[18705]_ , \new_[18706]_ ,
    \new_[18707]_ , \new_[18708]_ , \new_[18709]_ , \new_[18710]_ ,
    \new_[18711]_ , \new_[18712]_ , \new_[18713]_ , \new_[18714]_ ,
    \new_[18715]_ , \new_[18716]_ , \new_[18717]_ , \new_[18718]_ ,
    \new_[18719]_ , \new_[18720]_ , \new_[18721]_ , \new_[18722]_ ,
    \new_[18723]_ , \new_[18724]_ , \new_[18725]_ , \new_[18727]_ ,
    \new_[18728]_ , \new_[18729]_ , \new_[18730]_ , \new_[18731]_ ,
    \new_[18732]_ , \new_[18733]_ , \new_[18734]_ , \new_[18735]_ ,
    \new_[18736]_ , \new_[18737]_ , \new_[18738]_ , \new_[18739]_ ,
    \new_[18740]_ , \new_[18741]_ , \new_[18742]_ , \new_[18743]_ ,
    \new_[18744]_ , \new_[18745]_ , \new_[18746]_ , \new_[18747]_ ,
    \new_[18748]_ , \new_[18749]_ , \new_[18750]_ , \new_[18751]_ ,
    \new_[18752]_ , \new_[18753]_ , \new_[18754]_ , \new_[18755]_ ,
    \new_[18756]_ , \new_[18757]_ , \new_[18758]_ , \new_[18759]_ ,
    \new_[18760]_ , \new_[18761]_ , \new_[18762]_ , \new_[18763]_ ,
    \new_[18764]_ , \new_[18765]_ , \new_[18766]_ , \new_[18767]_ ,
    \new_[18768]_ , \new_[18769]_ , \new_[18770]_ , \new_[18771]_ ,
    \new_[18772]_ , \new_[18773]_ , \new_[18774]_ , \new_[18775]_ ,
    \new_[18776]_ , \new_[18777]_ , \new_[18778]_ , \new_[18779]_ ,
    \new_[18780]_ , \new_[18781]_ , \new_[18782]_ , \new_[18783]_ ,
    \new_[18784]_ , \new_[18785]_ , \new_[18786]_ , \new_[18787]_ ,
    \new_[18788]_ , \new_[18789]_ , \new_[18790]_ , \new_[18791]_ ,
    \new_[18792]_ , \new_[18793]_ , \new_[18794]_ , \new_[18795]_ ,
    \new_[18796]_ , \new_[18797]_ , \new_[18798]_ , \new_[18799]_ ,
    \new_[18800]_ , \new_[18801]_ , \new_[18802]_ , \new_[18803]_ ,
    \new_[18804]_ , \new_[18805]_ , \new_[18806]_ , \new_[18807]_ ,
    \new_[18809]_ , \new_[18810]_ , \new_[18811]_ , \new_[18812]_ ,
    \new_[18813]_ , \new_[18814]_ , \new_[18815]_ , \new_[18816]_ ,
    \new_[18817]_ , \new_[18818]_ , \new_[18819]_ , \new_[18820]_ ,
    \new_[18821]_ , \new_[18824]_ , \new_[18825]_ , \new_[18826]_ ,
    \new_[18827]_ , \new_[18828]_ , \new_[18829]_ , \new_[18830]_ ,
    \new_[18831]_ , \new_[18832]_ , \new_[18833]_ , \new_[18834]_ ,
    \new_[18835]_ , \new_[18836]_ , \new_[18837]_ , \new_[18838]_ ,
    \new_[18839]_ , \new_[18840]_ , \new_[18841]_ , \new_[18842]_ ,
    \new_[18843]_ , \new_[18844]_ , \new_[18845]_ , \new_[18846]_ ,
    \new_[18847]_ , \new_[18848]_ , \new_[18849]_ , \new_[18850]_ ,
    \new_[18851]_ , \new_[18852]_ , \new_[18853]_ , \new_[18854]_ ,
    \new_[18855]_ , \new_[18856]_ , \new_[18857]_ , \new_[18858]_ ,
    \new_[18859]_ , \new_[18860]_ , \new_[18862]_ , \new_[18863]_ ,
    \new_[18864]_ , \new_[18865]_ , \new_[18866]_ , \new_[18867]_ ,
    \new_[18868]_ , \new_[18869]_ , \new_[18870]_ , \new_[18871]_ ,
    \new_[18872]_ , \new_[18873]_ , \new_[18874]_ , \new_[18875]_ ,
    \new_[18876]_ , \new_[18877]_ , \new_[18878]_ , \new_[18879]_ ,
    \new_[18880]_ , \new_[18881]_ , \new_[18882]_ , \new_[18883]_ ,
    \new_[18884]_ , \new_[18885]_ , \new_[18886]_ , \new_[18887]_ ,
    \new_[18888]_ , \new_[18889]_ , \new_[18890]_ , \new_[18891]_ ,
    \new_[18892]_ , \new_[18893]_ , \new_[18894]_ , \new_[18895]_ ,
    \new_[18896]_ , \new_[18897]_ , \new_[18898]_ , \new_[18899]_ ,
    \new_[18900]_ , \new_[18901]_ , \new_[18902]_ , \new_[18903]_ ,
    \new_[18904]_ , \new_[18905]_ , \new_[18906]_ , \new_[18907]_ ,
    \new_[18908]_ , \new_[18909]_ , \new_[18910]_ , \new_[18911]_ ,
    \new_[18912]_ , \new_[18913]_ , \new_[18914]_ , \new_[18916]_ ,
    \new_[18917]_ , \new_[18918]_ , \new_[18919]_ , \new_[18920]_ ,
    \new_[18921]_ , \new_[18922]_ , \new_[18923]_ , \new_[18924]_ ,
    \new_[18925]_ , \new_[18926]_ , \new_[18927]_ , \new_[18928]_ ,
    \new_[18929]_ , \new_[18930]_ , \new_[18931]_ , \new_[18932]_ ,
    \new_[18933]_ , \new_[18934]_ , \new_[18935]_ , \new_[18936]_ ,
    \new_[18937]_ , \new_[18938]_ , \new_[18939]_ , \new_[18940]_ ,
    \new_[18941]_ , \new_[18942]_ , \new_[18943]_ , \new_[18944]_ ,
    \new_[18945]_ , \new_[18946]_ , \new_[18947]_ , \new_[18948]_ ,
    \new_[18949]_ , \new_[18950]_ , \new_[18951]_ , \new_[18952]_ ,
    \new_[18953]_ , \new_[18954]_ , \new_[18955]_ , \new_[18956]_ ,
    \new_[18957]_ , \new_[18958]_ , \new_[18959]_ , \new_[18960]_ ,
    \new_[18961]_ , \new_[18962]_ , \new_[18963]_ , \new_[18964]_ ,
    \new_[18965]_ , \new_[18966]_ , \new_[18967]_ , \new_[18968]_ ,
    \new_[18969]_ , \new_[18970]_ , \new_[18971]_ , \new_[18972]_ ,
    \new_[18973]_ , \new_[18974]_ , \new_[18975]_ , \new_[18976]_ ,
    \new_[18977]_ , \new_[18978]_ , \new_[18979]_ , \new_[18980]_ ,
    \new_[18981]_ , \new_[18982]_ , \new_[18983]_ , \new_[18984]_ ,
    \new_[18985]_ , \new_[18986]_ , \new_[18987]_ , \new_[18988]_ ,
    \new_[18989]_ , \new_[18990]_ , \new_[18991]_ , \new_[18992]_ ,
    \new_[18993]_ , \new_[18994]_ , \new_[18995]_ , \new_[18996]_ ,
    \new_[18997]_ , \new_[18998]_ , \new_[18999]_ , \new_[19000]_ ,
    \new_[19001]_ , \new_[19002]_ , \new_[19003]_ , \new_[19004]_ ,
    \new_[19005]_ , \new_[19006]_ , \new_[19007]_ , \new_[19008]_ ,
    \new_[19009]_ , \new_[19010]_ , \new_[19011]_ , \new_[19012]_ ,
    \new_[19013]_ , \new_[19014]_ , \new_[19015]_ , \new_[19016]_ ,
    \new_[19017]_ , \new_[19018]_ , \new_[19019]_ , \new_[19020]_ ,
    \new_[19021]_ , \new_[19022]_ , \new_[19023]_ , \new_[19024]_ ,
    \new_[19025]_ , \new_[19026]_ , \new_[19027]_ , \new_[19028]_ ,
    \new_[19029]_ , \new_[19030]_ , \new_[19031]_ , \new_[19032]_ ,
    \new_[19033]_ , \new_[19034]_ , \new_[19035]_ , \new_[19036]_ ,
    \new_[19037]_ , \new_[19038]_ , \new_[19039]_ , \new_[19040]_ ,
    \new_[19042]_ , \new_[19043]_ , \new_[19044]_ , \new_[19045]_ ,
    \new_[19046]_ , \new_[19047]_ , \new_[19048]_ , \new_[19049]_ ,
    \new_[19050]_ , \new_[19052]_ , \new_[19053]_ , \new_[19054]_ ,
    \new_[19055]_ , \new_[19056]_ , \new_[19057]_ , \new_[19058]_ ,
    \new_[19059]_ , \new_[19060]_ , \new_[19061]_ , \new_[19062]_ ,
    \new_[19063]_ , \new_[19064]_ , \new_[19065]_ , \new_[19066]_ ,
    \new_[19067]_ , \new_[19068]_ , \new_[19069]_ , \new_[19070]_ ,
    \new_[19071]_ , \new_[19072]_ , \new_[19073]_ , \new_[19074]_ ,
    \new_[19075]_ , \new_[19076]_ , \new_[19077]_ , \new_[19078]_ ,
    \new_[19079]_ , \new_[19080]_ , \new_[19081]_ , \new_[19082]_ ,
    \new_[19083]_ , \new_[19084]_ , \new_[19085]_ , \new_[19086]_ ,
    \new_[19087]_ , \new_[19088]_ , \new_[19089]_ , \new_[19090]_ ,
    \new_[19091]_ , \new_[19092]_ , \new_[19093]_ , \new_[19094]_ ,
    \new_[19095]_ , \new_[19096]_ , \new_[19097]_ , \new_[19098]_ ,
    \new_[19099]_ , \new_[19100]_ , \new_[19101]_ , \new_[19102]_ ,
    \new_[19103]_ , \new_[19104]_ , \new_[19105]_ , \new_[19106]_ ,
    \new_[19107]_ , \new_[19108]_ , \new_[19109]_ , \new_[19110]_ ,
    \new_[19111]_ , \new_[19112]_ , \new_[19113]_ , \new_[19114]_ ,
    \new_[19115]_ , \new_[19116]_ , \new_[19117]_ , \new_[19118]_ ,
    \new_[19119]_ , \new_[19120]_ , \new_[19121]_ , \new_[19122]_ ,
    \new_[19123]_ , \new_[19124]_ , \new_[19125]_ , \new_[19126]_ ,
    \new_[19127]_ , \new_[19128]_ , \new_[19129]_ , \new_[19130]_ ,
    \new_[19131]_ , \new_[19132]_ , \new_[19133]_ , \new_[19134]_ ,
    \new_[19135]_ , \new_[19136]_ , \new_[19137]_ , \new_[19138]_ ,
    \new_[19139]_ , \new_[19140]_ , \new_[19142]_ , \new_[19143]_ ,
    \new_[19144]_ , \new_[19145]_ , \new_[19146]_ , \new_[19147]_ ,
    \new_[19148]_ , \new_[19149]_ , \new_[19150]_ , \new_[19151]_ ,
    \new_[19152]_ , \new_[19153]_ , \new_[19154]_ , \new_[19155]_ ,
    \new_[19156]_ , \new_[19157]_ , \new_[19158]_ , \new_[19159]_ ,
    \new_[19160]_ , \new_[19161]_ , \new_[19162]_ , \new_[19163]_ ,
    \new_[19164]_ , \new_[19165]_ , \new_[19166]_ , \new_[19167]_ ,
    \new_[19168]_ , \new_[19169]_ , \new_[19170]_ , \new_[19171]_ ,
    \new_[19172]_ , \new_[19173]_ , \new_[19174]_ , \new_[19175]_ ,
    \new_[19176]_ , \new_[19177]_ , \new_[19178]_ , \new_[19179]_ ,
    \new_[19180]_ , \new_[19181]_ , \new_[19182]_ , \new_[19183]_ ,
    \new_[19184]_ , \new_[19185]_ , \new_[19186]_ , \new_[19187]_ ,
    \new_[19188]_ , \new_[19189]_ , \new_[19190]_ , \new_[19191]_ ,
    \new_[19192]_ , \new_[19193]_ , \new_[19194]_ , \new_[19195]_ ,
    \new_[19196]_ , \new_[19197]_ , \new_[19198]_ , \new_[19199]_ ,
    \new_[19200]_ , \new_[19201]_ , \new_[19202]_ , \new_[19203]_ ,
    \new_[19204]_ , \new_[19205]_ , \new_[19206]_ , \new_[19207]_ ,
    \new_[19208]_ , \new_[19209]_ , \new_[19210]_ , \new_[19211]_ ,
    \new_[19212]_ , \new_[19213]_ , \new_[19214]_ , \new_[19215]_ ,
    \new_[19217]_ , \new_[19218]_ , \new_[19219]_ , \new_[19220]_ ,
    \new_[19221]_ , \new_[19223]_ , \new_[19224]_ , \new_[19225]_ ,
    \new_[19226]_ , \new_[19227]_ , \new_[19228]_ , \new_[19229]_ ,
    \new_[19230]_ , \new_[19231]_ , \new_[19232]_ , \new_[19233]_ ,
    \new_[19234]_ , \new_[19235]_ , \new_[19236]_ , \new_[19237]_ ,
    \new_[19238]_ , \new_[19239]_ , \new_[19240]_ , \new_[19241]_ ,
    \new_[19242]_ , \new_[19243]_ , \new_[19244]_ , \new_[19245]_ ,
    \new_[19246]_ , \new_[19247]_ , \new_[19248]_ , \new_[19249]_ ,
    \new_[19250]_ , \new_[19251]_ , \new_[19252]_ , \new_[19253]_ ,
    \new_[19254]_ , \new_[19255]_ , \new_[19256]_ , \new_[19257]_ ,
    \new_[19258]_ , \new_[19259]_ , \new_[19260]_ , \new_[19261]_ ,
    \new_[19262]_ , \new_[19263]_ , \new_[19265]_ , \new_[19266]_ ,
    \new_[19267]_ , \new_[19268]_ , \new_[19269]_ , \new_[19270]_ ,
    \new_[19271]_ , \new_[19272]_ , \new_[19273]_ , \new_[19274]_ ,
    \new_[19275]_ , \new_[19276]_ , \new_[19277]_ , \new_[19278]_ ,
    \new_[19279]_ , \new_[19280]_ , \new_[19281]_ , \new_[19282]_ ,
    \new_[19283]_ , \new_[19284]_ , \new_[19285]_ , \new_[19286]_ ,
    \new_[19287]_ , \new_[19288]_ , \new_[19289]_ , \new_[19290]_ ,
    \new_[19291]_ , \new_[19292]_ , \new_[19293]_ , \new_[19294]_ ,
    \new_[19295]_ , \new_[19296]_ , \new_[19297]_ , \new_[19298]_ ,
    \new_[19299]_ , \new_[19300]_ , \new_[19301]_ , \new_[19302]_ ,
    \new_[19303]_ , \new_[19304]_ , \new_[19305]_ , \new_[19306]_ ,
    \new_[19307]_ , \new_[19308]_ , \new_[19309]_ , \new_[19310]_ ,
    \new_[19311]_ , \new_[19312]_ , \new_[19313]_ , \new_[19314]_ ,
    \new_[19315]_ , \new_[19316]_ , \new_[19317]_ , \new_[19318]_ ,
    \new_[19319]_ , \new_[19320]_ , \new_[19321]_ , \new_[19322]_ ,
    \new_[19323]_ , \new_[19324]_ , \new_[19325]_ , \new_[19326]_ ,
    \new_[19327]_ , \new_[19328]_ , \new_[19329]_ , \new_[19330]_ ,
    \new_[19331]_ , \new_[19332]_ , \new_[19333]_ , \new_[19334]_ ,
    \new_[19335]_ , \new_[19336]_ , \new_[19337]_ , \new_[19338]_ ,
    \new_[19339]_ , \new_[19340]_ , \new_[19341]_ , \new_[19342]_ ,
    \new_[19343]_ , \new_[19344]_ , \new_[19345]_ , \new_[19346]_ ,
    \new_[19347]_ , \new_[19348]_ , \new_[19349]_ , \new_[19350]_ ,
    \new_[19351]_ , \new_[19352]_ , \new_[19353]_ , \new_[19354]_ ,
    \new_[19355]_ , \new_[19356]_ , \new_[19357]_ , \new_[19358]_ ,
    \new_[19359]_ , \new_[19360]_ , \new_[19361]_ , \new_[19362]_ ,
    \new_[19363]_ , \new_[19364]_ , \new_[19365]_ , \new_[19366]_ ,
    \new_[19367]_ , \new_[19368]_ , \new_[19369]_ , \new_[19370]_ ,
    \new_[19371]_ , \new_[19372]_ , \new_[19373]_ , \new_[19374]_ ,
    \new_[19375]_ , \new_[19376]_ , \new_[19377]_ , \new_[19378]_ ,
    \new_[19379]_ , \new_[19380]_ , \new_[19381]_ , \new_[19382]_ ,
    \new_[19383]_ , \new_[19384]_ , \new_[19385]_ , \new_[19386]_ ,
    \new_[19387]_ , \new_[19388]_ , \new_[19389]_ , \new_[19390]_ ,
    \new_[19391]_ , \new_[19392]_ , \new_[19393]_ , \new_[19394]_ ,
    \new_[19395]_ , \new_[19396]_ , \new_[19397]_ , \new_[19398]_ ,
    \new_[19399]_ , \new_[19400]_ , \new_[19401]_ , \new_[19402]_ ,
    \new_[19403]_ , \new_[19404]_ , \new_[19405]_ , \new_[19406]_ ,
    \new_[19407]_ , \new_[19408]_ , \new_[19409]_ , \new_[19410]_ ,
    \new_[19411]_ , \new_[19412]_ , \new_[19413]_ , \new_[19414]_ ,
    \new_[19415]_ , \new_[19416]_ , \new_[19417]_ , \new_[19418]_ ,
    \new_[19419]_ , \new_[19420]_ , \new_[19421]_ , \new_[19422]_ ,
    \new_[19423]_ , \new_[19424]_ , \new_[19425]_ , \new_[19426]_ ,
    \new_[19427]_ , \new_[19428]_ , \new_[19429]_ , \new_[19430]_ ,
    \new_[19431]_ , \new_[19432]_ , \new_[19433]_ , \new_[19434]_ ,
    \new_[19435]_ , \new_[19436]_ , \new_[19437]_ , \new_[19438]_ ,
    \new_[19439]_ , \new_[19440]_ , \new_[19441]_ , \new_[19442]_ ,
    \new_[19443]_ , \new_[19444]_ , \new_[19445]_ , \new_[19446]_ ,
    \new_[19447]_ , \new_[19448]_ , \new_[19449]_ , \new_[19450]_ ,
    \new_[19451]_ , \new_[19452]_ , \new_[19453]_ , \new_[19454]_ ,
    \new_[19455]_ , \new_[19456]_ , \new_[19457]_ , \new_[19458]_ ,
    \new_[19459]_ , \new_[19460]_ , \new_[19461]_ , \new_[19462]_ ,
    \new_[19463]_ , \new_[19464]_ , \new_[19465]_ , \new_[19466]_ ,
    \new_[19467]_ , \new_[19468]_ , \new_[19469]_ , \new_[19470]_ ,
    \new_[19471]_ , \new_[19472]_ , \new_[19473]_ , \new_[19474]_ ,
    \new_[19475]_ , \new_[19476]_ , \new_[19477]_ , \new_[19478]_ ,
    \new_[19479]_ , \new_[19480]_ , \new_[19481]_ , \new_[19482]_ ,
    \new_[19483]_ , \new_[19484]_ , \new_[19485]_ , \new_[19486]_ ,
    \new_[19487]_ , \new_[19488]_ , \new_[19489]_ , \new_[19490]_ ,
    \new_[19491]_ , \new_[19492]_ , \new_[19493]_ , \new_[19494]_ ,
    \new_[19495]_ , \new_[19496]_ , \new_[19497]_ , \new_[19498]_ ,
    \new_[19499]_ , \new_[19500]_ , \new_[19501]_ , \new_[19502]_ ,
    \new_[19503]_ , \new_[19504]_ , \new_[19505]_ , \new_[19506]_ ,
    \new_[19507]_ , \new_[19508]_ , \new_[19509]_ , \new_[19510]_ ,
    \new_[19511]_ , \new_[19512]_ , \new_[19513]_ , \new_[19514]_ ,
    \new_[19515]_ , \new_[19516]_ , \new_[19517]_ , \new_[19518]_ ,
    \new_[19519]_ , \new_[19520]_ , \new_[19521]_ , \new_[19522]_ ,
    \new_[19523]_ , \new_[19524]_ , \new_[19525]_ , \new_[19526]_ ,
    \new_[19527]_ , \new_[19528]_ , \new_[19529]_ , \new_[19530]_ ,
    \new_[19531]_ , \new_[19532]_ , \new_[19533]_ , \new_[19534]_ ,
    \new_[19535]_ , \new_[19536]_ , \new_[19537]_ , \new_[19538]_ ,
    \new_[19539]_ , \new_[19540]_ , \new_[19541]_ , \new_[19542]_ ,
    \new_[19543]_ , \new_[19544]_ , \new_[19545]_ , \new_[19546]_ ,
    \new_[19547]_ , \new_[19548]_ , \new_[19549]_ , \new_[19550]_ ,
    \new_[19551]_ , \new_[19553]_ , \new_[19554]_ , \new_[19555]_ ,
    \new_[19556]_ , \new_[19557]_ , \new_[19558]_ , \new_[19559]_ ,
    \new_[19560]_ , \new_[19561]_ , \new_[19562]_ , \new_[19563]_ ,
    \new_[19564]_ , \new_[19565]_ , \new_[19566]_ , \new_[19567]_ ,
    \new_[19568]_ , \new_[19569]_ , \new_[19570]_ , \new_[19571]_ ,
    \new_[19572]_ , \new_[19573]_ , \new_[19574]_ , \new_[19575]_ ,
    \new_[19576]_ , \new_[19577]_ , \new_[19578]_ , \new_[19579]_ ,
    \new_[19580]_ , \new_[19581]_ , \new_[19582]_ , \new_[19583]_ ,
    \new_[19584]_ , \new_[19585]_ , \new_[19586]_ , \new_[19587]_ ,
    \new_[19588]_ , \new_[19589]_ , \new_[19590]_ , \new_[19591]_ ,
    \new_[19592]_ , \new_[19593]_ , \new_[19594]_ , \new_[19595]_ ,
    \new_[19596]_ , \new_[19597]_ , \new_[19598]_ , \new_[19599]_ ,
    \new_[19600]_ , \new_[19601]_ , \new_[19602]_ , \new_[19603]_ ,
    \new_[19604]_ , \new_[19605]_ , \new_[19606]_ , \new_[19607]_ ,
    \new_[19608]_ , \new_[19609]_ , \new_[19610]_ , \new_[19611]_ ,
    \new_[19612]_ , \new_[19613]_ , \new_[19614]_ , \new_[19615]_ ,
    \new_[19616]_ , \new_[19617]_ , \new_[19618]_ , \new_[19619]_ ,
    \new_[19620]_ , \new_[19621]_ , \new_[19622]_ , \new_[19623]_ ,
    \new_[19624]_ , \new_[19625]_ , \new_[19626]_ , \new_[19628]_ ,
    \new_[19629]_ , \new_[19630]_ , \new_[19631]_ , \new_[19632]_ ,
    \new_[19633]_ , \new_[19634]_ , \new_[19635]_ , \new_[19636]_ ,
    \new_[19637]_ , \new_[19638]_ , \new_[19639]_ , \new_[19640]_ ,
    \new_[19641]_ , \new_[19642]_ , \new_[19643]_ , \new_[19644]_ ,
    \new_[19645]_ , \new_[19646]_ , \new_[19647]_ , \new_[19648]_ ,
    \new_[19649]_ , \new_[19650]_ , \new_[19651]_ , \new_[19652]_ ,
    \new_[19653]_ , \new_[19654]_ , \new_[19655]_ , \new_[19656]_ ,
    \new_[19657]_ , \new_[19658]_ , \new_[19659]_ , \new_[19660]_ ,
    \new_[19661]_ , \new_[19662]_ , \new_[19663]_ , \new_[19664]_ ,
    \new_[19665]_ , \new_[19666]_ , \new_[19667]_ , \new_[19668]_ ,
    \new_[19669]_ , \new_[19670]_ , \new_[19671]_ , \new_[19672]_ ,
    \new_[19673]_ , \new_[19674]_ , \new_[19675]_ , \new_[19676]_ ,
    \new_[19677]_ , \new_[19678]_ , \new_[19679]_ , \new_[19680]_ ,
    \new_[19681]_ , \new_[19682]_ , \new_[19683]_ , \new_[19684]_ ,
    \new_[19685]_ , \new_[19686]_ , \new_[19687]_ , \new_[19688]_ ,
    \new_[19689]_ , \new_[19690]_ , \new_[19691]_ , \new_[19692]_ ,
    \new_[19693]_ , \new_[19694]_ , \new_[19695]_ , \new_[19696]_ ,
    \new_[19697]_ , \new_[19698]_ , \new_[19699]_ , \new_[19700]_ ,
    \new_[19701]_ , \new_[19702]_ , \new_[19703]_ , \new_[19704]_ ,
    \new_[19705]_ , \new_[19706]_ , \new_[19707]_ , \new_[19708]_ ,
    \new_[19709]_ , \new_[19710]_ , \new_[19711]_ , \new_[19712]_ ,
    \new_[19713]_ , \new_[19714]_ , \new_[19715]_ , \new_[19716]_ ,
    \new_[19717]_ , \new_[19718]_ , \new_[19719]_ , \new_[19720]_ ,
    \new_[19721]_ , \new_[19722]_ , \new_[19723]_ , \new_[19724]_ ,
    \new_[19725]_ , \new_[19726]_ , \new_[19727]_ , \new_[19729]_ ,
    \new_[19730]_ , \new_[19731]_ , \new_[19732]_ , \new_[19733]_ ,
    \new_[19734]_ , \new_[19735]_ , \new_[19736]_ , \new_[19737]_ ,
    \new_[19738]_ , \new_[19739]_ , \new_[19740]_ , \new_[19741]_ ,
    \new_[19742]_ , \new_[19743]_ , \new_[19744]_ , \new_[19745]_ ,
    \new_[19746]_ , \new_[19747]_ , \new_[19748]_ , \new_[19749]_ ,
    \new_[19750]_ , \new_[19751]_ , \new_[19752]_ , \new_[19753]_ ,
    \new_[19754]_ , \new_[19755]_ , \new_[19756]_ , \new_[19757]_ ,
    \new_[19759]_ , \new_[19760]_ , \new_[19761]_ , \new_[19762]_ ,
    \new_[19763]_ , \new_[19764]_ , \new_[19765]_ , \new_[19766]_ ,
    \new_[19767]_ , \new_[19768]_ , \new_[19769]_ , \new_[19770]_ ,
    \new_[19771]_ , \new_[19772]_ , \new_[19773]_ , \new_[19774]_ ,
    \new_[19775]_ , \new_[19776]_ , \new_[19777]_ , \new_[19778]_ ,
    \new_[19779]_ , \new_[19780]_ , \new_[19781]_ , \new_[19782]_ ,
    \new_[19783]_ , \new_[19784]_ , \new_[19785]_ , \new_[19786]_ ,
    \new_[19787]_ , \new_[19788]_ , \new_[19789]_ , \new_[19790]_ ,
    \new_[19791]_ , \new_[19792]_ , \new_[19793]_ , \new_[19794]_ ,
    \new_[19795]_ , \new_[19796]_ , \new_[19797]_ , \new_[19798]_ ,
    \new_[19799]_ , \new_[19800]_ , \new_[19801]_ , \new_[19802]_ ,
    \new_[19803]_ , \new_[19804]_ , \new_[19805]_ , \new_[19806]_ ,
    \new_[19807]_ , \new_[19808]_ , \new_[19809]_ , \new_[19810]_ ,
    \new_[19811]_ , \new_[19812]_ , \new_[19813]_ , \new_[19814]_ ,
    \new_[19815]_ , \new_[19816]_ , \new_[19817]_ , \new_[19818]_ ,
    \new_[19819]_ , \new_[19820]_ , \new_[19821]_ , \new_[19822]_ ,
    \new_[19823]_ , \new_[19824]_ , \new_[19825]_ , \new_[19826]_ ,
    \new_[19827]_ , \new_[19828]_ , \new_[19831]_ , \new_[19832]_ ,
    \new_[19833]_ , \new_[19834]_ , \new_[19835]_ , \new_[19836]_ ,
    \new_[19837]_ , \new_[19838]_ , \new_[19839]_ , \new_[19840]_ ,
    \new_[19841]_ , \new_[19842]_ , \new_[19843]_ , \new_[19844]_ ,
    \new_[19845]_ , \new_[19846]_ , \new_[19847]_ , \new_[19848]_ ,
    \new_[19849]_ , \new_[19850]_ , \new_[19851]_ , \new_[19852]_ ,
    \new_[19853]_ , \new_[19854]_ , \new_[19855]_ , \new_[19856]_ ,
    \new_[19857]_ , \new_[19858]_ , \new_[19859]_ , \new_[19860]_ ,
    \new_[19861]_ , \new_[19862]_ , \new_[19863]_ , \new_[19864]_ ,
    \new_[19865]_ , \new_[19866]_ , \new_[19867]_ , \new_[19868]_ ,
    \new_[19869]_ , \new_[19870]_ , \new_[19871]_ , \new_[19872]_ ,
    \new_[19873]_ , \new_[19874]_ , \new_[19875]_ , \new_[19876]_ ,
    \new_[19877]_ , \new_[19878]_ , \new_[19879]_ , \new_[19880]_ ,
    \new_[19881]_ , \new_[19882]_ , \new_[19883]_ , \new_[19884]_ ,
    \new_[19885]_ , \new_[19886]_ , \new_[19887]_ , \new_[19888]_ ,
    \new_[19889]_ , \new_[19890]_ , \new_[19891]_ , \new_[19892]_ ,
    \new_[19893]_ , \new_[19895]_ , \new_[19896]_ , \new_[19897]_ ,
    \new_[19899]_ , \new_[19900]_ , \new_[19901]_ , \new_[19902]_ ,
    \new_[19903]_ , \new_[19904]_ , \new_[19905]_ , \new_[19906]_ ,
    \new_[19907]_ , \new_[19908]_ , \new_[19909]_ , \new_[19910]_ ,
    \new_[19911]_ , \new_[19912]_ , \new_[19913]_ , \new_[19914]_ ,
    \new_[19916]_ , \new_[19917]_ , \new_[19918]_ , \new_[19919]_ ,
    \new_[19920]_ , \new_[19921]_ , \new_[19922]_ , \new_[19923]_ ,
    \new_[19924]_ , \new_[19925]_ , \new_[19926]_ , \new_[19927]_ ,
    \new_[19928]_ , \new_[19929]_ , \new_[19930]_ , \new_[19931]_ ,
    \new_[19932]_ , \new_[19933]_ , \new_[19934]_ , \new_[19935]_ ,
    \new_[19936]_ , \new_[19937]_ , \new_[19938]_ , \new_[19939]_ ,
    \new_[19940]_ , \new_[19941]_ , \new_[19942]_ , \new_[19943]_ ,
    \new_[19944]_ , \new_[19945]_ , \new_[19946]_ , \new_[19947]_ ,
    \new_[19948]_ , \new_[19949]_ , \new_[19950]_ , \new_[19951]_ ,
    \new_[19952]_ , \new_[19953]_ , \new_[19954]_ , \new_[19955]_ ,
    \new_[19956]_ , \new_[19957]_ , \new_[19958]_ , \new_[19959]_ ,
    \new_[19960]_ , \new_[19961]_ , \new_[19962]_ , \new_[19963]_ ,
    \new_[19964]_ , \new_[19965]_ , \new_[19966]_ , \new_[19967]_ ,
    \new_[19968]_ , \new_[19969]_ , \new_[19970]_ , \new_[19971]_ ,
    \new_[19972]_ , \new_[19973]_ , \new_[19974]_ , \new_[19975]_ ,
    \new_[19977]_ , \new_[19978]_ , \new_[19979]_ , \new_[19980]_ ,
    \new_[19981]_ , \new_[19982]_ , \new_[19983]_ , \new_[19984]_ ,
    \new_[19985]_ , \new_[19986]_ , \new_[19987]_ , \new_[19988]_ ,
    \new_[19989]_ , \new_[19990]_ , \new_[19991]_ , \new_[19992]_ ,
    \new_[19993]_ , \new_[19995]_ , \new_[19996]_ , \new_[19997]_ ,
    \new_[19998]_ , \new_[19999]_ , \new_[20000]_ , \new_[20001]_ ,
    \new_[20002]_ , \new_[20003]_ , \new_[20004]_ , \new_[20005]_ ,
    \new_[20006]_ , \new_[20007]_ , \new_[20008]_ , \new_[20009]_ ,
    \new_[20010]_ , \new_[20011]_ , \new_[20012]_ , \new_[20013]_ ,
    \new_[20014]_ , \new_[20015]_ , \new_[20016]_ , \new_[20017]_ ,
    \new_[20018]_ , \new_[20019]_ , \new_[20020]_ , \new_[20021]_ ,
    \new_[20022]_ , \new_[20023]_ , \new_[20024]_ , \new_[20025]_ ,
    \new_[20026]_ , \new_[20027]_ , \new_[20028]_ , \new_[20029]_ ,
    \new_[20030]_ , \new_[20031]_ , \new_[20032]_ , \new_[20033]_ ,
    \new_[20034]_ , \new_[20035]_ , \new_[20036]_ , \new_[20037]_ ,
    \new_[20038]_ , \new_[20039]_ , \new_[20040]_ , \new_[20041]_ ,
    \new_[20042]_ , \new_[20043]_ , \new_[20044]_ , \new_[20045]_ ,
    \new_[20046]_ , \new_[20047]_ , \new_[20048]_ , \new_[20049]_ ,
    \new_[20050]_ , \new_[20051]_ , \new_[20052]_ , \new_[20053]_ ,
    \new_[20054]_ , \new_[20055]_ , \new_[20056]_ , \new_[20057]_ ,
    \new_[20058]_ , \new_[20059]_ , \new_[20060]_ , \new_[20061]_ ,
    \new_[20062]_ , \new_[20063]_ , \new_[20064]_ , \new_[20065]_ ,
    \new_[20066]_ , \new_[20067]_ , \new_[20068]_ , \new_[20069]_ ,
    \new_[20070]_ , \new_[20071]_ , \new_[20072]_ , \new_[20073]_ ,
    \new_[20074]_ , \new_[20075]_ , \new_[20076]_ , \new_[20077]_ ,
    \new_[20078]_ , \new_[20079]_ , \new_[20080]_ , \new_[20081]_ ,
    \new_[20082]_ , \new_[20083]_ , \new_[20084]_ , \new_[20085]_ ,
    \new_[20086]_ , \new_[20087]_ , \new_[20088]_ , \new_[20089]_ ,
    \new_[20090]_ , \new_[20091]_ , \new_[20092]_ , \new_[20093]_ ,
    \new_[20094]_ , \new_[20095]_ , \new_[20096]_ , \new_[20097]_ ,
    \new_[20098]_ , \new_[20099]_ , \new_[20100]_ , \new_[20101]_ ,
    \new_[20103]_ , \new_[20104]_ , \new_[20105]_ , \new_[20106]_ ,
    \new_[20107]_ , \new_[20108]_ , \new_[20109]_ , \new_[20110]_ ,
    \new_[20111]_ , \new_[20112]_ , \new_[20113]_ , \new_[20114]_ ,
    \new_[20115]_ , \new_[20116]_ , \new_[20117]_ , \new_[20118]_ ,
    \new_[20119]_ , \new_[20120]_ , \new_[20121]_ , \new_[20122]_ ,
    \new_[20123]_ , \new_[20124]_ , \new_[20125]_ , \new_[20126]_ ,
    \new_[20127]_ , \new_[20128]_ , \new_[20129]_ , \new_[20130]_ ,
    \new_[20131]_ , \new_[20133]_ , \new_[20134]_ , \new_[20135]_ ,
    \new_[20136]_ , \new_[20137]_ , \new_[20138]_ , \new_[20139]_ ,
    \new_[20140]_ , \new_[20141]_ , \new_[20142]_ , \new_[20143]_ ,
    \new_[20144]_ , \new_[20145]_ , \new_[20146]_ , \new_[20147]_ ,
    \new_[20148]_ , \new_[20149]_ , \new_[20150]_ , \new_[20151]_ ,
    \new_[20152]_ , \new_[20153]_ , \new_[20154]_ , \new_[20155]_ ,
    \new_[20156]_ , \new_[20157]_ , \new_[20158]_ , \new_[20159]_ ,
    \new_[20160]_ , \new_[20161]_ , \new_[20162]_ , \new_[20163]_ ,
    \new_[20164]_ , \new_[20165]_ , \new_[20166]_ , \new_[20167]_ ,
    \new_[20168]_ , \new_[20169]_ , \new_[20170]_ , \new_[20171]_ ,
    \new_[20172]_ , \new_[20173]_ , \new_[20174]_ , \new_[20175]_ ,
    \new_[20176]_ , \new_[20177]_ , \new_[20178]_ , \new_[20179]_ ,
    \new_[20180]_ , \new_[20181]_ , \new_[20182]_ , \new_[20183]_ ,
    \new_[20184]_ , \new_[20185]_ , \new_[20186]_ , \new_[20187]_ ,
    \new_[20188]_ , \new_[20189]_ , \new_[20190]_ , \new_[20191]_ ,
    \new_[20192]_ , \new_[20193]_ , \new_[20194]_ , \new_[20195]_ ,
    \new_[20196]_ , \new_[20197]_ , \new_[20198]_ , \new_[20199]_ ,
    \new_[20200]_ , \new_[20201]_ , \new_[20202]_ , \new_[20203]_ ,
    \new_[20204]_ , \new_[20205]_ , \new_[20206]_ , \new_[20207]_ ,
    \new_[20209]_ , \new_[20210]_ , \new_[20211]_ , \new_[20212]_ ,
    \new_[20213]_ , \new_[20214]_ , \new_[20215]_ , \new_[20216]_ ,
    \new_[20217]_ , \new_[20218]_ , \new_[20220]_ , \new_[20221]_ ,
    \new_[20222]_ , \new_[20223]_ , \new_[20224]_ , \new_[20225]_ ,
    \new_[20226]_ , \new_[20227]_ , \new_[20228]_ , \new_[20229]_ ,
    \new_[20230]_ , \new_[20231]_ , \new_[20233]_ , \new_[20234]_ ,
    \new_[20235]_ , \new_[20236]_ , \new_[20237]_ , \new_[20238]_ ,
    \new_[20240]_ , \new_[20241]_ , \new_[20242]_ , \new_[20243]_ ,
    \new_[20245]_ , \new_[20246]_ , \new_[20247]_ , \new_[20248]_ ,
    \new_[20249]_ , \new_[20250]_ , \new_[20252]_ , \new_[20253]_ ,
    \new_[20254]_ , \new_[20255]_ , \new_[20256]_ , \new_[20257]_ ,
    \new_[20258]_ , \new_[20259]_ , \new_[20261]_ , \new_[20262]_ ,
    \new_[20263]_ , \new_[20264]_ , \new_[20265]_ , \new_[20266]_ ,
    \new_[20268]_ , \new_[20269]_ , \new_[20270]_ , \new_[20271]_ ,
    \new_[20272]_ , \new_[20273]_ , \new_[20275]_ , \new_[20276]_ ,
    \new_[20277]_ , \new_[20278]_ , \new_[20279]_ , \new_[20280]_ ,
    \new_[20281]_ , \new_[20282]_ , \new_[20283]_ , \new_[20284]_ ,
    \new_[20285]_ , \new_[20286]_ , \new_[20287]_ , \new_[20288]_ ,
    \new_[20289]_ , \new_[20290]_ , \new_[20291]_ , \new_[20292]_ ,
    \new_[20293]_ , \new_[20294]_ , \new_[20295]_ , \new_[20296]_ ,
    \new_[20297]_ , \new_[20298]_ , \new_[20299]_ , \new_[20300]_ ,
    \new_[20301]_ , \new_[20302]_ , \new_[20303]_ , \new_[20304]_ ,
    \new_[20305]_ , \new_[20307]_ , \new_[20308]_ , \new_[20309]_ ,
    \new_[20310]_ , \new_[20311]_ , \new_[20312]_ , \new_[20313]_ ,
    \new_[20314]_ , \new_[20315]_ , \new_[20316]_ , \new_[20317]_ ,
    \new_[20318]_ , \new_[20319]_ , \new_[20320]_ , \new_[20321]_ ,
    \new_[20322]_ , \new_[20323]_ , \new_[20324]_ , \new_[20325]_ ,
    \new_[20326]_ , \new_[20327]_ , \new_[20328]_ , \new_[20329]_ ,
    \new_[20330]_ , \new_[20331]_ , \new_[20332]_ , \new_[20333]_ ,
    \new_[20334]_ , \new_[20335]_ , \new_[20336]_ , \new_[20337]_ ,
    \new_[20338]_ , \new_[20339]_ , \new_[20340]_ , \new_[20341]_ ,
    \new_[20342]_ , \new_[20343]_ , \new_[20344]_ , \new_[20345]_ ,
    \new_[20346]_ , \new_[20347]_ , \new_[20348]_ , \new_[20349]_ ,
    \new_[20350]_ , \new_[20351]_ , \new_[20352]_ , \new_[20353]_ ,
    \new_[20354]_ , \new_[20355]_ , \new_[20356]_ , \new_[20357]_ ,
    \new_[20358]_ , \new_[20359]_ , \new_[20360]_ , \new_[20361]_ ,
    \new_[20362]_ , \new_[20363]_ , \new_[20364]_ , \new_[20365]_ ,
    \new_[20366]_ , \new_[20367]_ , \new_[20368]_ , \new_[20369]_ ,
    \new_[20370]_ , \new_[20371]_ , \new_[20372]_ , \new_[20373]_ ,
    \new_[20374]_ , \new_[20375]_ , \new_[20376]_ , \new_[20377]_ ,
    \new_[20378]_ , \new_[20379]_ , \new_[20380]_ , \new_[20381]_ ,
    \new_[20382]_ , \new_[20383]_ , \new_[20384]_ , \new_[20385]_ ,
    \new_[20386]_ , \new_[20387]_ , \new_[20388]_ , \new_[20389]_ ,
    \new_[20390]_ , \new_[20391]_ , \new_[20392]_ , \new_[20393]_ ,
    \new_[20394]_ , \new_[20395]_ , \new_[20396]_ , \new_[20397]_ ,
    \new_[20398]_ , \new_[20399]_ , \new_[20400]_ , \new_[20401]_ ,
    \new_[20402]_ , \new_[20403]_ , \new_[20404]_ , \new_[20405]_ ,
    \new_[20406]_ , \new_[20407]_ , \new_[20408]_ , \new_[20409]_ ,
    \new_[20410]_ , \new_[20411]_ , \new_[20412]_ , \new_[20413]_ ,
    \new_[20414]_ , \new_[20415]_ , \new_[20416]_ , \new_[20417]_ ,
    \new_[20418]_ , \new_[20419]_ , \new_[20420]_ , \new_[20421]_ ,
    \new_[20422]_ , \new_[20423]_ , \new_[20424]_ , \new_[20425]_ ,
    \new_[20426]_ , \new_[20427]_ , \new_[20428]_ , \new_[20429]_ ,
    \new_[20430]_ , \new_[20431]_ , \new_[20432]_ , \new_[20433]_ ,
    \new_[20434]_ , \new_[20435]_ , \new_[20436]_ , \new_[20437]_ ,
    \new_[20438]_ , \new_[20439]_ , \new_[20440]_ , \new_[20441]_ ,
    \new_[20442]_ , \new_[20443]_ , \new_[20444]_ , \new_[20445]_ ,
    \new_[20446]_ , \new_[20447]_ , \new_[20448]_ , \new_[20449]_ ,
    \new_[20450]_ , \new_[20451]_ , \new_[20452]_ , \new_[20453]_ ,
    \new_[20454]_ , \new_[20455]_ , \new_[20456]_ , \new_[20457]_ ,
    \new_[20458]_ , \new_[20459]_ , \new_[20460]_ , \new_[20461]_ ,
    \new_[20462]_ , \new_[20463]_ , \new_[20464]_ , \new_[20465]_ ,
    \new_[20466]_ , \new_[20467]_ , \new_[20468]_ , \new_[20469]_ ,
    \new_[20470]_ , \new_[20471]_ , \new_[20472]_ , \new_[20473]_ ,
    \new_[20474]_ , \new_[20475]_ , \new_[20476]_ , \new_[20477]_ ,
    \new_[20478]_ , \new_[20479]_ , \new_[20480]_ , \new_[20481]_ ,
    \new_[20482]_ , \new_[20483]_ , \new_[20484]_ , \new_[20485]_ ,
    \new_[20486]_ , \new_[20487]_ , \new_[20488]_ , \new_[20489]_ ,
    \new_[20490]_ , \new_[20491]_ , \new_[20492]_ , \new_[20493]_ ,
    \new_[20494]_ , \new_[20495]_ , \new_[20496]_ , \new_[20497]_ ,
    \new_[20498]_ , \new_[20499]_ , \new_[20500]_ , \new_[20501]_ ,
    \new_[20502]_ , \new_[20503]_ , \new_[20504]_ , \new_[20505]_ ,
    \new_[20506]_ , \new_[20507]_ , \new_[20508]_ , \new_[20509]_ ,
    \new_[20510]_ , \new_[20511]_ , \new_[20512]_ , \new_[20513]_ ,
    \new_[20514]_ , \new_[20515]_ , \new_[20516]_ , \new_[20517]_ ,
    \new_[20518]_ , \new_[20519]_ , \new_[20520]_ , \new_[20521]_ ,
    \new_[20523]_ , \new_[20524]_ , \new_[20525]_ , \new_[20526]_ ,
    \new_[20527]_ , \new_[20528]_ , \new_[20529]_ , \new_[20530]_ ,
    \new_[20531]_ , \new_[20532]_ , \new_[20533]_ , \new_[20534]_ ,
    \new_[20535]_ , \new_[20536]_ , \new_[20537]_ , \new_[20538]_ ,
    \new_[20539]_ , \new_[20540]_ , \new_[20541]_ , \new_[20542]_ ,
    \new_[20543]_ , \new_[20544]_ , \new_[20545]_ , \new_[20546]_ ,
    \new_[20547]_ , \new_[20548]_ , \new_[20549]_ , \new_[20550]_ ,
    \new_[20551]_ , \new_[20552]_ , \new_[20553]_ , \new_[20554]_ ,
    \new_[20555]_ , n740, n745, n750, n755, n760, n765, n770, n775, n780,
    n785, n790, n795, n800, n805, n810, n815, n820, n825, n830, n835, n840,
    n845, n850, n855, n860, n865, n870, n875, n880, n885, n890, n895, n900,
    n905, n910, n915, n920, n925, n930, n935, n940, n945, n950, n955, n960,
    n965, n970, n975, n980, n985, n990, n995, n1000, n1005, n1010, n1015,
    n1020, n1025, n1030, n1035, n1040, n1045, n1050, n1055, n1060, n1065,
    n1070, n1075, n1080, n1085, n1090, n1095, n1100, n1105, n1110, n1115,
    n1120, n1125, n1130, n1135, n1140, n1145, n1150, n1155, n1160, n1165,
    n1170, n1175, n1180, n1185, n1190, n1195, n1200, n1205, n1210, n1215,
    n1220, n1225, n1230, n1235, n1240, n1245, n1250, n1255, n1260, n1265,
    n1270, n1275, n1280, n1285, n1290, n1295, n1300, n1305, n1310, n1315,
    n1320, n1325, n1330, n1335, n1340, n1345, n1350, n1355, n1360, n1365,
    n1370, n1375, n1380, n1385, n1390, n1395, n1400, n1405, n1410, n1415,
    n1420, n1425, n1430, n1435, n1440, n1445, n1450, n1455, n1460, n1465,
    n1470, n1475, n1480, n1485, n1490, n1495, n1500, n1505, n1510, n1515,
    n1520, n1525, n1530, n1535, n1540, n1545, n1550, n1555, n1560, n1565,
    n1570, n1575, n1580, n1585, n1590, n1595, n1600, n1605, n1610, n1615,
    n1620, n1625, n1630, n1635, n1640, n1645, n1650, n1655, n1660, n1665,
    n1670, n1675, n1680, n1685, n1690, n1695, n1700, n1705, n1710, n1715,
    n1720, n1725, n1730, n1735, n1740, n1745, n1750, n1755, n1760, n1765,
    n1770, n1775, n1780, n1785, n1790, n1795, n1800, n1805, n1810, n1815,
    n1820, n1825, n1830, n1835, n1840, n1845, n1850, n1855, n1860, n1865,
    n1870, n1875, n1880, n1885, n1890, n1895, n1900, n1905, n1910, n1915,
    n1920, n1925, n1930, n1935, n1940, n1945, n1950, n1955, n1960, n1965,
    n1970, n1975, n1980, n1985, n1990, n1995, n2000, n2005, n2010, n2015,
    n2020, n2025, n2030, n2035, n2040, n2045, n2050, n2055, n2060, n2065,
    n2070, n2075, n2080, n2085, n2090, n2095, n2100, n2105, n2110, n2115,
    n2120, n2125, n2130, n2135, n2140, n2145, n2150, n2155, n2160, n2165,
    n2170, n2175, n2180, n2185, n2190, n2195, n2200, n2205, n2210, n2215,
    n2220, n2225, n2230, n2235, n2240, n2245, n2250, n2255, n2260, n2265,
    n2270, n2275, n2280, n2285, n2290, n2295, n2300, n2305, n2310, n2315,
    n2320, n2325, n2330, n2335, n2340, n2345, n2350, n2355, n2360, n2365,
    n2370, n2375, n2380, n2385, n2390, n2395, n2400, n2405, n2410, n2415,
    n2420, n2425, n2430, n2435, n2440, n2445, n2450, n2455, n2460, n2465,
    n2470, n2475, n2480, n2485, n2490, n2495, n2500, n2505, n2510, n2515,
    n2520, n2525, n2530, n2535, n2540, n2545, n2550, n2555, n2560, n2565,
    n2570, n2575, n2580, n2585, n2590, n2595, n2600, n2605, n2610, n2615,
    n2620, n2625, n2630, n2635, n2640, n2645, n2650, n2655, n2660, n2665,
    n2670, n2675, n2680, n2685, n2690, n2695, n2700, n2705, n2710, n2715,
    n2720, n2725, n2730, n2735, n2740, n2745, n2750, n2755, n2760, n2765,
    n2770, n2775, n2780, n2785, n2790, n2795, n2800, n2805, n2810, n2815,
    n2820, n2825, n2830, n2835, n2840, n2845, n2850, n2855, n2860, n2865,
    n2870, n2875, n2880, n2885, n2890, n2895, n2900, n2905, n2910, n2915,
    n2920, n2925, n2930, n2935, n2940, n2945, n2950, n2955, n2960, n2965,
    n2970, n2975, n2980, n2985, n2990, n2995, n3000, n3005, n3010, n3015,
    n3020, n3025, n3030, n3035, n3040, n3045, n3050, n3055, n3060, n3065,
    n3070, n3075, n3080, n3085, n3090, n3095, n3100, n3105, n3110, n3115,
    n3120, n3125, n3130, n3135, n3140, n3145, n3150, n3155, n3160, n3165,
    n3170, n3175, n3180, n3185, n3190, n3195, n3200, n3205, n3210, n3215,
    n3220, n3225, n3230, n3235, n3240, n3245, n3250, n3255, n3260, n3265,
    n3270, n3275, n3280, n3285, n3290, n3295, n3300, n3305, n3310, n3315,
    n3320, n3325, n3330, n3335, n3340, n3345, n3350, n3355, n3360, n3365,
    n3370, n3375, n3380, n3385, n3390, n3395, n3400, n3405, n3410, n3415,
    n3420, n3425, n3430, n3435, n3440, n3445, n3450, n3455, n3460, n3465,
    n3470, n3475, n3480, n3485, n3490, n3495, n3500, n3505, n3510, n3515,
    n3520, n3525, n3530, n3535, n3540, n3545, n3550, n3555, n3560, n3565,
    n3570, n3575, n3580, n3585, n3590, n3595, n3600, n3605, n3610, n3615,
    n3620, n3625, n3630, n3635, n3640, n3645, n3650, n3655, n3660, n3665,
    n3670, n3675, n3680, n3685, n3690, n3695, n3700, n3705, n3710, n3715,
    n3720, n3725, n3730, n3735, n3740, n3745, n3750, n3755, n3760, n3765,
    n3770, n3775, n3780, n3785, n3790, n3795, n3800, n3805, n3810, n3815,
    n3820, n3825, n3830, n3835, n3840, n3845, n3850, n3855, n3860, n3865,
    n3870, n3875, n3880, n3885, n3890, n3895, n3900, n3905, n3910, n3915,
    n3920, n3925, n3930, n3935, n3940, n3945, n3950, n3955, n3960, n3965,
    n3970, n3975, n3980, n3985, n3990, n3995, n4000, n4005, n4010, n4015,
    n4020, n4025, n4030, n4035, n4040, n4045, n4050, n4055, n4060, n4065,
    n4070, n4075, n4080, n4085, n4090, n4095, n4100, n4105, n4110, n4115,
    n4120, n4125, n4130, n4135, n4140, n4145, n4150, n4155, n4160, n4165,
    n4170, n4175, n4180, n4185, n4190, n4195, n4200, n4205, n4210, n4215,
    n4220, n4225, n4230, n4235, n4240, n4245, n4250, n4255, n4260, n4265,
    n4270, n4275, n4280, n4285, n4290, n4295, n4300, n4305, n4310, n4315,
    n4320, n4325, n4330, n4335, n4340, n4345, n4350, n4355, n4360, n4365,
    n4370, n4375, n4380, n4385, n4390, n4395, n4400, n4405, n4410, n4415,
    n4420, n4425, n4430, n4435, n4440, n4445, n4450, n4455, n4460, n4465,
    n4470, n4475, n4480, n4485, n4490, n4495, n4500, n4505, n4510, n4515,
    n4520, n4525, n4530, n4535, n4540, n4545, n4550, n4555, n4560, n4565,
    n4570, n4575, n4580, n4585, n4590, n4595, n4600, n4605, n4610, n4615,
    n4620, n4625, n4630, n4635, n4640, n4645, n4650, n4655, n4660, n4665,
    n4670, n4675, n4680, n4685, n4690, n4695, n4700, n4705, n4710, n4715,
    n4720, n4725, n4730, n4735, n4740, n4745, n4750, n4755, n4760, n4765,
    n4770, n4775, n4780, n4785, n4790, n4795, n4800, n4805, n4810, n4815,
    n4820, n4825, n4830, n4835, n4840, n4845, n4850, n4855, n4860, n4865,
    n4870, n4875, n4880, n4885, n4890, n4895, n4900, n4905, n4910, n4915,
    n4920, n4925, n4930, n4935, n4940, n4945, n4950, n4955, n4960, n4965,
    n4970, n4975, n4980, n4985, n4990, n4995, n5000, n5005, n5010, n5015,
    n5020, n5025, n5030, n5035, n5040, n5045, n5050, n5055, n5060, n5065,
    n5070, n5075, n5080, n5085, n5090, n5095, n5100, n5105, n5110, n5115,
    n5120, n5125, n5130, n5135, n5140, n5145, n5150, n5155, n5160, n5165,
    n5170, n5175, n5180, n5185, n5190, n5195, n5200, n5205, n5210, n5215,
    n5220, n5225, n5230, n5235, n5240, n5245, n5250, n5255, n5260, n5265,
    n5270, n5275, n5280, n5285, n5290, n5295, n5300, n5305, n5310, n5315,
    n5320, n5325, n5330, n5335, n5340, n5345, n5350, n5355, n5360, n5365,
    n5370, n5375, n5380, n5385, n5390, n5395, n5400, n5405, n5410, n5415,
    n5420, n5425, n5430, n5435, n5440, n5445, n5450, n5455, n5460, n5465,
    n5470, n5475, n5480, n5485, n5490, n5495, n5500, n5505, n5510, n5515,
    n5520, n5525, n5530, n5535, n5540, n5545, n5550, n5555, n5560, n5565,
    n5570, n5575, n5580, n5585, n5590, n5595, n5600, n5605, n5610, n5615,
    n5620, n5625, n5630, n5635, n5640, n5645, n5650, n5655, n5660, n5665,
    n5670, n5675, n5680, n5685, n5690, n5695, n5700, n5705, n5710, n5715,
    n5720, n5725, n5730, n5735, n5740, n5745, n5750, n5755, n5760, n5765,
    n5770, n5775, n5780, n5785, n5790, n5795, n5800, n5805, n5810, n5815,
    n5820, n5825, n5830, n5835, n5840, n5845, n5850, n5855, n5860, n5865,
    n5870, n5875, n5880, n5885, n5890, n5895, n5900, n5905, n5910, n5915,
    n5920, n5925, n5930, n5935, n5940, n5945, n5950, n5955, n5960, n5965,
    n5970, n5975, n5980, n5985, n5990, n5995, n6000, n6005, n6010, n6015,
    n6020, n6025, n6030, n6035, n6040, n6045, n6050, n6055, n6060, n6065,
    n6070, n6075, n6080, n6085, n6090, n6095, n6100, n6105, n6110, n6115,
    n6120, n6125, n6130, n6135, n6140, n6145, n6150, n6155, n6160, n6165,
    n6170, n6175, n6180, n6185, n6190, n6195, n6200, n6205, n6210, n6215,
    n6220, n6225, n6230, n6235, n6240, n6245, n6250, n6255, n6260, n6265,
    n6270, n6275, n6280, n6285, n6290, n6295, n6300, n6305, n6310, n6315,
    n6320, n6325, n6330, n6335, n6340, n6345, n6350, n6355, n6360, n6365,
    n6370, n6375, n6380, n6385, n6390, n6395, n6400, n6405, n6410, n6415,
    n6420, n6425, n6430, n6435, n6440, n6445, n6450, n6455, n6460, n6465,
    n6470, n6475, n6480, n6485, n6490, n6495, n6500, n6505, n6510, n6515,
    n6520, n6525, n6530, n6535, n6540, n6545, n6550, n6555, n6560, n6565,
    n6570, n6575, n6580, n6585, n6590, n6595, n6600, n6605, n6610, n6615,
    n6620, n6625, n6630, n6635, n6640, n6645, n6650, n6655, n6660, n6665,
    n6670, n6675, n6680, n6685, n6690, n6695, n6700, n6705, n6710, n6715,
    n6720, n6725, n6730, n6735, n6740, n6745, n6750, n6755, n6760, n6765,
    n6770, n6775, n6780, n6785, n6790, n6795, n6800, n6805, n6810, n6815,
    n6820, n6825, n6830, n6835, n6840, n6845, n6850, n6855, n6860, n6865,
    n6870, n6875, n6880, n6885, n6890, n6895, n6900, n6905, n6910, n6915,
    n6920, n6925, n6930, n6935, n6940, n6945, n6950, n6955, n6960, n6965,
    n6970, n6975, n6980, n6985, n6990, n6995, n7000, n7005, n7010, n7015,
    n7020, n7025, n7030, n7035, n7040, n7045, n7050, n7055, n7060, n7065,
    n7070, n7075, n7080, n7085, n7090, n7095, n7100, n7105, n7110, n7115,
    n7120, n7125, n7130, n7135, n7140, n7145, n7150, n7155, n7160, n7165,
    n7170, n7175, n7180, n7185, n7190, n7195, n7200, n7205, n7210, n7215,
    n7220, n7225, n7230, n7235, n7240, n7245, n7250, n7255, n7260, n7265,
    n7270, n7275, n7280, n7285, n7290, n7295, n7300, n7305, n7310, n7315,
    n7320, n7325, n7330, n7335, n7340, n7345, n7350, n7355, n7360, n7365,
    n7370, n7375, n7380, n7385, n7390, n7395, n7400, n7405, n7410, n7415,
    n7420, n7425, n7430, n7435, n7440, n7445, n7450, n7455, n7460, n7465,
    n7470, n7475, n7480, n7485, n7490, n7495, n7500, n7505, n7510, n7515,
    n7520, n7525, n7530, n7535, n7540, n7545, n7550, n7555, n7560, n7565,
    n7570, n7575, n7580, n7585, n7590, n7595, n7600, n7605, n7610, n7615,
    n7620, n7625, n7630, n7635, n7640, n7645, n7650, n7655, n7660, n7665,
    n7670, n7675, n7680, n7685, n7690, n7695, n7700, n7705, n7710, n7715,
    n7720, n7725, n7730, n7735, n7740, n7745, n7750, n7755, n7760, n7765,
    n7770, n7775, n7780, n7785, n7790, n7795, n7800, n7805, n7810, n7815,
    n7820, n7825, n7830, n7835, n7840, n7845, n7850, n7855, n7860, n7865,
    n7870, n7875, n7880, n7885, n7890, n7895, n7900, n7905, n7910, n7915,
    n7920, n7925, n7930, n7935, n7940, n7945, n7950, n7955, n7960, n7965,
    n7970, n7975, n7980, n7985, n7990, n7995, n8000, n8005, n8010, n8015,
    n8020, n8025, n8030, n8035, n8040, n8045, n8050, n8055, n8060, n8065,
    n8070, n8075, n8080, n8085, n8090, n8095, n8100, n8105, n8110, n8115,
    n8120, n8125, n8130, n8135, n8140, n8145, n8150, n8155, n8160, n8165,
    n8170, n8175, n8180, n8185, n8190, n8195, n8200, n8205, n8210, n8215,
    n8220, n8225, n8230, n8235, n8240, n8245, n8250, n8255, n8260, n8265,
    n8270, n8275, n8280, n8285, n8290, n8295, n8300, n8305, n8310, n8315,
    n8320, n8325, n8330, n8335, n8340, n8345, n8350, n8355, n8360, n8365,
    n8370, n8375, n8380, n8385, n8390, n8395, n8400, n8405, n8410, n8415,
    n8420, n8425, n8430, n8435, n8440, n8445, n8450, n8455, n8460, n8465,
    n8470, n8475, n8480, n8485, n8490, n8495, n8500, n8505, n8510, n8515,
    n8520, n8525, n8530, n8535, n8540, n8545, n8550, n8555, n8560, n8565,
    n8570, n8575, n8580, n8585, n8590, n8595, n8600, n8605, n8610, n8615,
    n8620, n8625, n8630, n8635, n8640, n8645, n8650, n8655, n8660, n8665,
    n8670, n8675, n8680, n8685, n8690, n8695, n8700, n8705, n8710, n8715,
    n8720, n8725, n8730, n8735, n8740, n8745, n8750, n8755, n8760, n8765,
    n8770, n8775, n8780, n8785, n8790, n8795, n8800, n8805, n8810, n8815,
    n8820, n8825, n8830, n8835, n8840, n8845, n8850, n8855, n8860, n8865,
    n8870, n8875, n8880, n8885, n8890, n8895, n8900, n8905, n8910, n8915,
    n8920, n8925, n8930, n8935, n8940, n8945, n8950, n8955, n8960, n8965,
    n8970, n8975, n8980, n8985, n8990, n8995, n9000, n9005, n9010, n9015,
    n9020, n9025, n9030, n9035, n9040, n9045, n9050, n9055, n9060, n9065,
    n9070, n9075, n9080, n9085, n9090, n9095, n9100, n9105, n9110, n9115,
    n9120, n9125, n9130, n9135, n9140, n9145, n9150, n9155, n9160, n9165,
    n9170, n9175, n9180, n9185, n9190, n9195, n9200, n9205, n9210, n9215,
    n9220, n9225, n9230, n9235, n9240, n9245, n9250, n9255, n9260, n9265,
    n9270, n9275, n9280, n9285, n9290, n9295, n9300, n9305, n9310, n9315,
    n9320, n9325, n9330, n9335, n9340, n9345, n9350, n9355, n9360, n9365,
    n9370, n9375, n9380, n9385, n9390, n9395, n9400, n9405, n9410, n9415,
    n9420, n9425, n9430, n9435, n9440, n9445, n9450, n9455, n9460, n9465,
    n9470, n9475, n9480, n9485, n9490, n9495, n9500, n9505, n9510, n9515,
    n9520, n9525, n9530, n9535, n9540, n9545, n9550, n9555, n9560, n9565,
    n9570, n9575, n9580, n9585, n9590, n9595, n9600, n9605, n9610, n9615,
    n9620, n9625, n9630, n9635, n9640, n9645, n9650, n9655, n9660, n9665,
    n9670, n9675, n9680, n9685, n9690, n9695, n9700, n9705, n9710, n9715,
    n9720, n9725, n9730, n9735, n9740, n9745, n9750, n9755, n9760, n9765,
    n9770, n9775, n9780, n9785, n9790, n9795, n9800, n9805, n9810, n9815,
    n9820, n9825, n9830, n9835, n9840, n9845, n9850, n9855, n9860, n9865,
    n9870, n9875, n9880, n9885, n9890, n9895, n9900, n9905, n9910, n9915,
    n9920, n9925, n9930, n9935, n9940, n9945, n9950, n9955, n9960, n9965,
    n9970, n9975, n9980, n9985, n9990, n9995, n10000, n10005, n10010,
    n10015, n10020, n10025, n10030, n10035, n10040, n10045, n10050, n10055,
    n10060, n10065, n10070, n10075, n10080, n10085, n10090, n10095, n10100,
    n10105, n10110, n10115, n10120, n10125, n10130, n10135, n10140, n10145,
    n10150, n10155, n10160, n10165, n10170, n10175, n10180, n10185, n10190,
    n10195, n10200, n10205, n10210, n10215, n10220, n10225, n10230, n10235,
    n10240, n10245, n10250, n10255, n10260, n10265, n10270, n10275, n10280,
    n10285, n10290, n10295, n10300, n10305, n10310, n10315, n10320, n10325,
    n10330, n10335, n10340, n10345, n10350, n10355, n10360, n10365, n10370,
    n10375, n10380, n10385, n10390, n10395, n10400, n10405, n10410, n10415,
    n10420, n10425, n10430, n10435, n10440, n10445, n10450, n10455, n10460,
    n10465, n10470, n10475, n10480, n10485, n10490, n10495, n10500, n10505,
    n10510, n10515, n10520, n10525, n10530, n10535, n10540, n10545, n10550,
    n10555, n10560, n10565, n10570, n10575, n10580, n10585, n10590, n10595,
    n10600, n10605, n10610, n10615, n10620, n10625, n10630, n10635, n10640,
    n10645, n10650, n10655, n10660, n10665, n10670, n10675, n10680, n10685,
    n10690, n10695, n10700, n10705, n10710, n10715, n10720, n10725, n10730,
    n10735, n10740, n10745, n10750, n10755, n10760, n10765, n10770, n10775,
    n10780, n10785, n10790, n10795, n10800, n10805, n10810, n10815, n10820,
    n10825, n10830, n10835, n10840, n10845, n10850, n10855, n10860, n10865,
    n10870, n10875, n10880, n10885, n10890, n10895, n10900, n10905, n10910,
    n10915, n10920, n10925, n10930, n10935, n10940, n10945, n10950, n10955,
    n10960, n10965, n10970, n10975, n10980, n10985, n10990, n10995, n11000,
    n11005, n11010, n11015, n11020, n11025, n11030, n11035, n11040, n11045,
    n11050, n11055, n11060, n11065, n11070, n11075, n11080, n11085, n11090,
    n11095, n11100, n11105, n11110, n11115, n11120, n11125, n11130, n11135,
    n11140, n11145, n11150, n11155, n11160, n11165, n11170, n11175, n11180,
    n11185, n11190, n11195, n11200, n11205, n11210, n11215, n11220, n11225,
    n11230, n11235, n11240, n11245, n11250, n11255, n11260, n11265, n11270,
    n11275, n11280, n11285, n11290, n11295, n11300, n11305, n11310, n11315,
    n11320, n11325, n11330, n11335, n11340, n11345, n11350, n11355, n11360,
    n11365, n11370, n11375, n11380, n11385, n11390, n11395, n11400, n11405,
    n11410, n11415, n11420, n11425, n11430, n11435, n11440, n11445, n11450,
    n11455, n11460, n11465, n11470, n11475, n11480, n11485, n11490, n11495,
    n11500, n11505, n11510, n11515, n11520, n11525, n11530, n11535, n11540,
    n11545, n11550, n11555, n11560, n11565, n11570, n11575, n11580, n11585,
    n11590, n11595, n11600, n11605, n11610, n11615, n11620, n11625, n11630,
    n11635, n11640, n11645, n11650, n11655, n11660, n11665, n11670, n11675,
    n11680, n11685, n11690, n11695, n11700, n11705, n11710, n11715, n11720,
    n11725, n11730, n11735, n11740, n11745, n11750, n11755, n11760, n11765,
    n11770, n11775, n11780, n11785, n11790, n11795, n11800, n11805, n11810,
    n11815, n11820, n11825, n11830, n11835, n11840, n11845, n11850, n11855,
    n11860, n11865, n11870, n11875, n11880, n11885, n11890, n11895, n11900,
    n11905, n11910, n11915, n11920, n11925, n11930, n11935, n11940, n11945,
    n11950, n11955, n11960, n11965, n11970, n11975, n11980, n11985, n11990,
    n11995, n12000, n12005, n12010, n12015, n12020, n12025, n12030, n12035,
    n12040, n12045, n12050, n12055, n12060, n12065, n12070, n12075, n12080,
    n12085, n12090, n12095, n12100, n12105, n12110, n12115, n12120, n12125,
    n12130, n12135, n12140, n12145, n12150, n12155, n12160, n12165, n12170,
    n12175, n12180, n12185, n12190, n12195, n12200, n12205, n12210, n12215,
    n12220, n12225, n12230, n12235, n12240, n12245, n12250, n12255, n12260,
    n12265, n12270, n12275, n12280, n12285, n12290, n12295, n12300, n12305,
    n12310, n12315, n12320, n12325, n12330, n12335, n12340, n12345, n12350,
    n12355, n12360, n12365, n12370, n12375, n12380, n12385, n12390, n12395,
    n12400, n12405, n12410, n12415, n12420, n12425, n12430, n12435, n12440,
    n12445, n12450, n12455, n12460, n12465, n12470, n12475, n12480, n12485,
    n12490, n12495, n12500, n12505, n12510, n12515, n12520, n12525, n12530,
    n12535, n12540, n12545, n12550, n12555, n12560, n12565, n12570, n12575,
    n12580, n12585, n12590, n12595, n12600, n12605, n12610, n12615, n12620,
    n12625, n12630, n12635, n12640, n12645, n12650, n12655, n12660, n12665,
    n12670, n12675, n12680, n12685, n12690, n12695, n12700, n12705, n12710,
    n12715, n12720, n12725, n12730, n12735, n12740, n12745, n12750, n12755,
    n12760, n12765, n12770, n12775, n12780, n12785, n12790, n12795, n12800,
    n12805, n12810, n12815, n12820, n12825, n12830, n12835, n12840, n12845,
    n12850, n12855, n12860, n12865, n12870, n12875, n12880, n12885, n12890,
    n12895, n12900, n12905, n12910, n12915, n12920, n12925, n12930, n12935,
    n12940, n12945, n12950, n12955, n12960, n12965, n12970, n12975, n12980,
    n12985, n12990, n12995, n13000, n13005, n13010, n13015, n13020, n13025,
    n13030, n13035, n13040, n13045, n13050, n13055, n13060, n13065, n13070,
    n13075, n13080, n13085, n13090, n13095, n13100, n13105, n13110, n13115,
    n13120, n13125, n13130, n13135, n13140, n13145, n13150, n13155, n13160,
    n13165, n13170, n13175, n13180, n13185, n13190, n13195, n13200, n13205,
    n13210, n13215, n13220, n13225, n13230, n13235, n13240, n13245, n13250,
    n13255, n13260, n13265, n13270, n13275, n13280, n13285, n13290, n13295,
    n13300, n13305, n13310, n13315, n13320, n13325, n13330, n13335, n13340,
    n13345, n13350, n13355, n13360, n13365, n13370, n13375, n13380, n13385,
    n13390, n13395, n13400, n13405, n13410, n13415, n13420, n13425, n13430,
    n13435, n13440, n13445, n13450, n13455, n13460, n13465, n13470, n13475,
    n13480, n13485, n13490, n13495, n13500, n13505, n13510, n13515, n13520,
    n13525, n13530, n13535, n13540, n13545, n13550, n13555, n13560, n13565,
    n13570, n13575, n13580, n13585, n13590, n13595, n13600, n13605, n13610,
    n13615, n13620, n13625, n13630, n13635, n13640, n13645, n13650, n13655,
    n13660, n13665, n13670, n13675, n13680, n13685, n13690, n13695, n13700,
    n13705, n13710, n13715, n13720, n13725, n13730, n13735, n13740, n13745,
    n13750, n13755, n13760, n13765, n13770, n13775, n13780, n13785, n13790,
    n13795, n13800, n13805, n13810, n13815, n13820, n13825, n13830, n13835,
    n13840, n13845, n13850, n13855, n13860, n13865, n13870, n13875, n13880,
    n13885, n13890, n13895, n13900, n13905, n13910, n13915, n13920, n13925,
    n13930, n13935, n13940, n13945, n13950, n13955, n13960, n13965, n13970,
    n13975, n13980, n13985, n13990, n13995, n14000, n14005, n14010, n14015,
    n14020, n14025, n14030, n14035, n14040, n14045, n14050, n14055, n14060,
    n14065, n14070, n14075, n14080, n14085, n14090, n14095, n14100, n14105,
    n14110, n14115, n14120, n14125, n14130, n14135, n14140, n14145, n14150,
    n14155, n14160, n14165, n14170, n14175, n14180, n14185, n14190, n14195,
    n14200, n14205, n14210, n14215, n14220, n14225, n14230, n14235, n14240,
    n14245, n14250, n14255, n14260, n14265, n14270, n14275, n14280, n14285,
    n14290, n14295, n14300, n14305, n14310, n14315, n14320, n14325, n14330,
    n14335, n14340, n14345, n14350, n14355, n14360, n14365, n14370, n14375,
    n14380, n14385, n14390, n14395, n14400, n14405, n14410, n14415, n14420,
    n14425, n14430, n14435, n14440, n14445, n14450, n14455, n14460, n14465,
    n14470, n14475, n14480, n14485, n14490, n14495, n14500, n14505, n14510,
    n14515, n14520, n14525, n14530, n14535, n14540, n14545, n14550, n14555,
    n14560, n14565, n14570, n14575, n14580, n14585, n14590, n14595, n14600,
    n14605, n14610, n14615, n14620, n14625, n14630, n14635, n14640, n14645,
    n14650, n14655, n14660, n14665, n14670, n14675, n14680, n14685, n14690,
    n14695, n14700, n14705, n14710, n14715, n14720, n14725, n14730, n14735,
    n14740, n14745, n14750, n14755, n14760, n14765, n14770, n14775, n14780,
    n14785, n14790, n14795, n14800, n14805, n14810, n14815, n14820, n14825,
    n14830, n14835, n14840, n14845, n14850, n14855, n14860, n14865, n14870,
    n14875, n14880, n14885, n14890, n14895, n14900, n14905, n14910, n14915,
    n14920, n14925, n14930, n14935, n14940, n14945, n14950, n14955, n14960,
    n14965, n14970, n14975, n14980, n14985, n14990, n14995, n15000, n15005,
    n15010, n15015, n15020, n15025, n15030, n15035, n15040, n15045, n15050,
    n15055, n15060, n15065, n15070, n15075, n15080, n15085, n15090, n15095,
    n15100, n15105, n15110, n15115, n15120, n15125, n15130, n15135, n15140,
    n15145, n15150, n15155, n15160, n15165, n15170, n15175, n15180, n15185,
    n15190, n15195, n15200, n15205, n15210, n15215, n15220, n15225, n15230,
    n15235, n15240, n15245, n15250, n15255, n15260, n15265, n15270, n15275,
    n15280, n15285, n15290, n15295, n15300, n15305, n15310, n15315, n15320,
    n15325, n15330, n15335, n15340, n15345, n15350, n15355, n15360, n15365,
    n15370, n15375, n15380, n15385, n15390, n15395, n15400, n15405, n15410,
    n15415, n15420, n15425, n15430, n15435, n15440, n15445, n15450, n15455,
    n15460, n15465, n15470, n15475, n15480, n15485, n15490, n15495, n15500,
    n15505, n15510, n15515, n15520, n15525, n15530, n15535, n15540, n15545,
    n15550, n15555, n15560, n15565, n15570, n15575, n15580, n15585, n15590,
    n15595, n15600, n15605, n15610, n15615, n15620, n15625, n15630, n15635,
    n15640, n15645, n15650, n15655, n15660, n15665, n15670, n15675, n15680,
    n15685, n15690, n15695, n15700, n15705, n15710, n15715, n15720, n15725,
    n15730, n15735, n15740, n15745, n15750, n15755, n15760, n15765, n15770,
    n15775, n15780, n15785, n15790, n15795, n15800, n15805, n15810, n15815,
    n15820, n15825, n15830, n15835, n15840, n15845, n15850, n15855, n15860,
    n15865, n15870, n15875, n15880, n15885, n15890, n15895, n15900, n15905,
    n15910, n15915, n15920, n15925, n15930, n15935, n15940, n15945, n15950,
    n15955, n15960, n15965, n15970, n15975, n15980, n15985, n15990, n15995,
    n16000, n16005, n16010, n16015, n16020, n16025, n16030, n16035, n16040,
    n16045, n16050, n16055, n16060, n16065, n16070, n16075, n16080, n16085,
    n16090, n16095, n16100, n16105, n16110, n16115, n16120, n16125, n16130,
    n16135, n16140, n16145, n16150, n16155, n16160, n16165, n16170, n16175,
    n16180, n16185, n16190, n16195, n16200, n16205, n16210, n16215, n16220,
    n16225, n16230, n16235, n16240, n16245, n16250, n16255, n16260, n16265,
    n16270, n16275, n16280, n16285, n16290, n16295, n16300, n16305, n16310,
    n16315, n16320, n16325, n16330, n16335, n16340, n16345, n16350, n16355,
    n16360, n16365, n16370, n16375, n16380, n16385, n16390, n16395, n16400,
    n16405, n16410, n16415, n16420, n16425, n16430, n16435, n16440, n16445,
    n16450, n16455, n16460, n16465, n16470, n16475, n16480, n16485, n16490,
    n16495, n16500, n16505, n16510, n16515, n16520, n16525, n16530, n16535,
    n16540, n16545, n16550, n16555, n16560, n16565, n16570, n16575, n16580,
    n16585, n16590, n16595, n16600, n16605, n16610, n16615, n16620, n16625,
    n16630, n16635, n16640, n16645, n16650, n16655, n16660, n16665, n16670,
    n16675, n16680, n16685, n16690, n16695, n16700, n16705, n16710, n16715,
    n16720, n16725, n16730, n16735, n16740, n16745, n16750, n16755, n16760,
    n16765, n16770, n16775, n16780, n16785, n16790, n16795, n16800, n16805,
    n16810, n16815, n16820, n16825, n16830, n16835, n16840, n16845, n16850,
    n16855, n16860, n16865, n16870, n16875, n16880, n16885, n16890, n16895,
    n16900, n16905, n16910, n16915, n16920, n16925, n16930, n16935, n16940,
    n16945, n16950, n16955, n16960, n16965, n16970, n16975, n16980, n16985,
    n16990, n16995, n17000, n17005, n17010, n17015, n17020, n17025, n17030,
    n17035, n17040, n17045, n17050, n17055, n17060, n17065, n17070, n17075,
    n17080, n17085, n17090, n17095, n17100, n17105, n17110, n17115, n17120,
    n17125, n17130, n17135, n17140, n17145, n17150, n17155, n17160, n17165,
    n17170, n17175, n17180, n17185, n17190, n17195, n17200, n17205, n17210,
    n17215, n17220, n17225, n17230, n17235, n17240, n17245, n17250, n17255,
    n17260, n17265, n17270, n17275, n17280, n17285, n17290, n17295, n17300,
    n17305, n17310, n17315, n17320, n17325, n17330, n17335, n17340, n17345,
    n17350, n17355, n17360, n17365, n17370, n17375, n17380, n17385, n17390,
    n17395, n17400, n17405, n17410, n17415, n17420, n17425, n17430, n17435,
    n17440, n17445, n17450, n17455, n17460, n17465, n17470, n17475, n17480,
    n17485, n17490, n17495, n17500, n17505, n17510, n17515, n17520, n17525,
    n17530;
  assign \new_[3728]_  = 1'b0;
  assign new_configuration_rst_inactive_sync_reg_in_ = 1'b1;
  assign pci_rst_oe_o = new_configuration_rst_inactive_sync_reg_in_;
  assign pci_inta_o = \new_[3728]_ ;
  assign pci_rst_o = \new_[3728]_ ;
  assign \wbm_bte_o[0]  = \new_[3728]_ ;
  assign \wbm_bte_o[1]  = \new_[3728]_ ;
  assign wb_int_o = \new_[3728]_ ;
  assign \wbm_cti_o[0]  = \\pci_target_unit_wishbone_master_wb_cti_o_reg[0] ;
  assign \wbm_cti_o[2]  = \\pci_target_unit_wishbone_master_wb_cti_o_reg[2] ;
  assign \new_[3738]_  = configuration_status_bit8_reg;
  assign n740 = ~\new_[4239]_  | ~\new_[3746]_  | ~\new_[4409]_ ;
  assign n745 = ~\new_[4239]_  | ~\new_[3747]_  | ~\new_[4410]_ ;
  assign n750 = ~\new_[10923]_  | (~\new_[3786]_  & ~\new_[15991]_ );
  assign \wbm_sel_o[0]  = \\pci_target_unit_wishbone_master_wb_sel_o_reg[0] ;
  assign \wbm_sel_o[1]  = \\pci_target_unit_wishbone_master_wb_sel_o_reg[1] ;
  assign \wbm_sel_o[2]  = \\pci_target_unit_wishbone_master_wb_sel_o_reg[2] ;
  assign \wbm_sel_o[3]  = \\pci_target_unit_wishbone_master_wb_sel_o_reg[3] ;
  assign \new_[3746]_  = \new_[3784]_  | \new_[5465]_ ;
  assign \new_[3747]_  = \new_[3785]_  | \new_[5465]_ ;
  assign \wbm_dat_o[0]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[0] ;
  assign \wbm_dat_o[10]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[10] ;
  assign \wbm_dat_o[11]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[11] ;
  assign \wbm_dat_o[12]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[12] ;
  assign \wbm_dat_o[13]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[13] ;
  assign \wbm_dat_o[16]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[16] ;
  assign \wbm_dat_o[17]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[17] ;
  assign \wbm_dat_o[19]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[19] ;
  assign \wbm_dat_o[1]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[1] ;
  assign \wbm_dat_o[20]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[20] ;
  assign \wbm_dat_o[21]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[21] ;
  assign \wbm_dat_o[22]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[22] ;
  assign \wbm_dat_o[23]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[23] ;
  assign \wbm_dat_o[24]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[24] ;
  assign \wbm_dat_o[25]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[25] ;
  assign \wbm_dat_o[26]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[26] ;
  assign \wbm_dat_o[27]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[27] ;
  assign \wbm_dat_o[28]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[28] ;
  assign \wbm_dat_o[29]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[29] ;
  assign \wbm_dat_o[2]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[2] ;
  assign \wbm_dat_o[31]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[31] ;
  assign \wbm_dat_o[3]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[3] ;
  assign \wbm_dat_o[4]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[4] ;
  assign \wbm_dat_o[5]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[5] ;
  assign \wbm_dat_o[6]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[6] ;
  assign \wbm_dat_o[8]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[8] ;
  assign \wbm_dat_o[9]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[9] ;
  assign \wbm_dat_o[30]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[30] ;
  assign \wbm_dat_o[14]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[14] ;
  assign \wbm_dat_o[18]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[18] ;
  assign \wbm_dat_o[7]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[7] ;
  assign \wbm_dat_o[15]  = \\pci_target_unit_wishbone_master_wb_dat_o_reg[15] ;
  assign n755 = ~\new_[5286]_  | ~\new_[5629]_  | ~\new_[3862]_ ;
  assign n765 = ~\new_[5288]_  | ~\new_[5629]_  | ~\new_[3864]_ ;
  assign n760 = ~\new_[5287]_  | ~\new_[5629]_  | ~\new_[3863]_ ;
  assign n770 = ~\new_[5289]_  | ~\new_[5629]_  | ~\new_[3865]_ ;
  assign \new_[3784]_  = ~\new_[3846]_  & (~\new_[4412]_  | ~\wbm_cti_o[0] );
  assign \new_[3785]_  = ~\new_[3846]_  & (~\new_[4412]_  | ~\wbm_cti_o[2] );
  assign \new_[3786]_  = ~\new_[4354]_  & (~\new_[3861]_  | ~\new_[17519]_ );
  assign \wbm_adr_o[19]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[19] ;
  assign \wbm_adr_o[22]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[22] ;
  assign \wbm_adr_o[24]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[24] ;
  assign \wbm_adr_o[20]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[20] ;
  assign \wbm_adr_o[27]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[27] ;
  assign \wbm_adr_o[21]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[21] ;
  assign \wbm_adr_o[30]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[30] ;
  assign \wbm_adr_o[25]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[25] ;
  assign \wbm_adr_o[28]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[28] ;
  assign \wbm_adr_o[31]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[31] ;
  assign \wbm_adr_o[29]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[29] ;
  assign \wbm_adr_o[17]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[17] ;
  assign \wbm_adr_o[10]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[10] ;
  assign \wbm_adr_o[11]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[11] ;
  assign \wbm_adr_o[12]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[12] ;
  assign \wbm_adr_o[16]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[16] ;
  assign \wbm_adr_o[14]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[14] ;
  assign \wbm_adr_o[13]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[13] ;
  assign \wbm_adr_o[23]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[23] ;
  assign \wbm_adr_o[26]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[26] ;
  assign \wbm_adr_o[3]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[3] ;
  assign \wbm_adr_o[4]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[4] ;
  assign \wbm_adr_o[5]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[5] ;
  assign \wbm_adr_o[6]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[6] ;
  assign \wbm_adr_o[8]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[8] ;
  assign \wbm_adr_o[9]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[9] ;
  assign \wbm_adr_o[2]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[2] ;
  assign n775 = ~\new_[5382]_  | (~\new_[3893]_  & ~\new_[20313]_ );
  assign n785 = ~\new_[5383]_  | (~\new_[3894]_  & ~\new_[5492]_ );
  assign n790 = ~\new_[5384]_  | (~\new_[3895]_  & ~\new_[20313]_ );
  assign n795 = ~\new_[5385]_  | (~\new_[3896]_  & ~\new_[20313]_ );
  assign n915 = ~\new_[5386]_  | (~\new_[3897]_  & ~\new_[5492]_ );
  assign n805 = ~\new_[5389]_  | (~\new_[3899]_  & ~\new_[20313]_ );
  assign n800 = ~\new_[5388]_  | (~\new_[3898]_  & ~\new_[20313]_ );
  assign n810 = ~\new_[5391]_  | (~\new_[3900]_  & ~\new_[20313]_ );
  assign n815 = ~\new_[5392]_  | (~\new_[3901]_  & ~\new_[5492]_ );
  assign n820 = ~\new_[5393]_  | (~\new_[3902]_  & ~\new_[5492]_ );
  assign n825 = ~\new_[5394]_  | (~\new_[3903]_  & ~\new_[5492]_ );
  assign n835 = ~\new_[5395]_  | (~\new_[3904]_  & ~\new_[20313]_ );
  assign n840 = ~\new_[5396]_  | (~\new_[3905]_  & ~\new_[20313]_ );
  assign n845 = ~\new_[5397]_  | (~\new_[3906]_  & ~\new_[20313]_ );
  assign n850 = ~\new_[5398]_  | (~\new_[3907]_  & ~\new_[20313]_ );
  assign n860 = ~\new_[5400]_  | (~\new_[3909]_  & ~\new_[20313]_ );
  assign n855 = ~\new_[5399]_  | (~\new_[3908]_  & ~\new_[20313]_ );
  assign n865 = ~\new_[5401]_  | (~\new_[3910]_  & ~\new_[5492]_ );
  assign n870 = ~\new_[5402]_  | (~\new_[3911]_  & ~\new_[5492]_ );
  assign n910 = ~\new_[5403]_  | (~\new_[3912]_  & ~\new_[20313]_ );
  assign n880 = ~\new_[5405]_  | (~\new_[3914]_  & ~\new_[5492]_ );
  assign n885 = ~\new_[5406]_  | (~\new_[3915]_  & ~\new_[20316]_ );
  assign n875 = ~\new_[5404]_  | (~\new_[3913]_  & ~\new_[20316]_ );
  assign n890 = ~\new_[5407]_  | (~\new_[3916]_  & ~\new_[20316]_ );
  assign n895 = ~\new_[5408]_  | (~\new_[3917]_  & ~\new_[20313]_ );
  assign n900 = ~\new_[5410]_  | (~\new_[3918]_  & ~\new_[20313]_ );
  assign n905 = ~\new_[5411]_  | (~\new_[3919]_  & ~\new_[20313]_ );
  assign \wbm_adr_o[18]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[18] ;
  assign \wbm_adr_o[15]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[15] ;
  assign \wbm_adr_o[7]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[7] ;
  assign \wbm_adr_o[0]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[0] ;
  assign \wbm_adr_o[1]  = \\pci_target_unit_wishbone_master_addr_cnt_out_reg[1] ;
  assign \new_[3846]_  = ~\new_[3889]_  & (~\new_[3921]_  | ~\new_[19874]_ );
  assign n930 = ~\new_[5387]_  | (~\new_[3922]_  & ~\new_[20316]_ );
  assign n920 = ~\new_[5390]_  | (~\new_[3923]_  & ~\new_[20313]_ );
  assign n925 = ~\new_[5409]_  | (~\new_[3924]_  & ~\new_[20313]_ );
  assign n1010 = \new_[14205]_  ? \new_[9763]_  : \new_[3988]_ ;
  assign n1015 = \new_[13787]_  ? \new_[9982]_  : \new_[3987]_ ;
  assign n1025 = \new_[14213]_  ? n6835 : \new_[3930]_ ;
  assign n1030 = \new_[13129]_  ? \new_[9763]_  : \new_[3933]_ ;
  assign n1065 = \new_[14915]_  ? \new_[9763]_  : \new_[3937]_ ;
  assign n1035 = \new_[14913]_  ? \new_[9763]_  : \new_[3940]_ ;
  assign n1040 = \new_[14886]_  ? \new_[9763]_  : \new_[3941]_ ;
  assign n1045 = \new_[14984]_  ? \new_[9763]_  : \new_[3942]_ ;
  assign n1050 = \new_[14976]_  ? \new_[9982]_  : \new_[3943]_ ;
  assign n1055 = \new_[14885]_  ? \new_[9763]_  : \new_[3945]_ ;
  assign n1060 = \new_[14983]_  ? n6835 : \new_[3946]_ ;
  assign \new_[3861]_  = parity_checker_perr_sampled_reg;
  assign \new_[3862]_  = \new_[3925]_  | \new_[20313]_ ;
  assign \new_[3863]_  = \new_[3926]_  | \new_[20313]_ ;
  assign \new_[3864]_  = \new_[3927]_  | \new_[20313]_ ;
  assign \new_[3865]_  = \new_[3928]_  | \new_[20313]_ ;
  assign n990 = \new_[13790]_  ? n6835 : \new_[3989]_ ;
  assign n935 = \new_[13816]_  ? \new_[9763]_  : \new_[3990]_ ;
  assign n950 = \new_[14211]_  ? n6835 : \new_[3991]_ ;
  assign n940 = \new_[13609]_  ? \new_[9763]_  : \new_[3929]_ ;
  assign n945 = \new_[13812]_  ? \new_[9763]_  : \new_[3931]_ ;
  assign n970 = \new_[13614]_  ? n6835 : \new_[3932]_ ;
  assign n955 = \new_[13210]_  ? \new_[9763]_  : \new_[3934]_ ;
  assign n960 = \new_[14855]_  ? n6835 : \new_[3992]_ ;
  assign n985 = \new_[13132]_  ? \new_[9982]_  : \new_[3936]_ ;
  assign n965 = \new_[11713]_  ? n6835 : \new_[3938]_ ;
  assign n975 = \new_[13798]_  ? \new_[9763]_  : \new_[3935]_ ;
  assign n980 = \new_[13149]_  ? \new_[9763]_  : \new_[3939]_ ;
  assign n995 = \new_[14845]_  ? \new_[9982]_  : \new_[3983]_ ;
  assign n1000 = \new_[14887]_  ? \new_[9763]_  : \new_[3984]_ ;
  assign n1005 = \new_[14871]_  ? \new_[9763]_  : \new_[3985]_ ;
  assign n1020 = \new_[14856]_  ? n6835 : \new_[3986]_ ;
  assign n1075 = \new_[14215]_  ? n6835 : \new_[4006]_ ;
  assign \new_[3883]_  = ~\\pci_target_unit_wishbone_master_bc_register_reg[0] ;
  assign \new_[3884]_  = ~\\pci_target_unit_wishbone_master_bc_register_reg[1] ;
  assign \new_[3885]_  = ~\\pci_target_unit_wishbone_master_bc_register_reg[2] ;
  assign \new_[3886]_  = ~\\pci_target_unit_wishbone_master_bc_register_reg[3] ;
  assign n17010 = pci_target_unit_wishbone_master_burst_chopped_reg;
  assign n1080 = \new_[14914]_  ? \new_[9763]_  : \new_[3993]_ ;
  assign \new_[3889]_  = ~\new_[3976]_  | ~\new_[4278]_ ;
  assign n1090 = ~\new_[9561]_  | ~\new_[3978]_ ;
  assign n1085 = ~\new_[9560]_  | ~\new_[3977]_ ;
  assign n1070 = \new_[13608]_  ? n6835 : \new_[4007]_ ;
  assign \new_[3893]_  = ~\new_[3947]_  & (~\new_[5299]_  | ~\wbm_dat_o[0] );
  assign \new_[3894]_  = ~\new_[3949]_  & (~\new_[20317]_  | ~\wbm_dat_o[11] );
  assign \new_[3895]_  = ~\new_[3950]_  & (~\new_[5299]_  | ~\wbm_dat_o[12] );
  assign \new_[3896]_  = ~\new_[3951]_  & (~\new_[20317]_  | ~\wbm_dat_o[13] );
  assign \new_[3897]_  = ~\new_[3952]_  & (~\new_[20317]_  | ~\wbm_dat_o[14] );
  assign \new_[3898]_  = ~\new_[3953]_  & (~\new_[5299]_  | ~\wbm_dat_o[16] );
  assign \new_[3899]_  = ~\new_[3954]_  & (~\new_[5299]_  | ~\wbm_dat_o[17] );
  assign \new_[3900]_  = ~\new_[3955]_  & (~\new_[20317]_  | ~\wbm_dat_o[19] );
  assign \new_[3901]_  = ~\new_[3956]_  & (~\new_[5299]_  | ~\wbm_dat_o[1] );
  assign \new_[3902]_  = ~\new_[3957]_  & (~\new_[20317]_  | ~\wbm_dat_o[20] );
  assign \new_[3903]_  = ~\new_[3958]_  & (~\new_[5299]_  | ~\wbm_dat_o[21] );
  assign \new_[3904]_  = ~\new_[3959]_  & (~\new_[5299]_  | ~\wbm_dat_o[23] );
  assign \new_[3905]_  = ~\new_[3960]_  & (~\new_[5299]_  | ~\wbm_dat_o[24] );
  assign \new_[3906]_  = ~\new_[3961]_  & (~\new_[20317]_  | ~\wbm_dat_o[25] );
  assign \new_[3907]_  = ~\new_[3962]_  & (~\new_[20317]_  | ~\wbm_dat_o[26] );
  assign \new_[3908]_  = ~\new_[3963]_  & (~\new_[20317]_  | ~\wbm_dat_o[27] );
  assign \new_[3909]_  = ~\new_[3964]_  & (~\new_[20317]_  | ~\wbm_dat_o[28] );
  assign \new_[3910]_  = ~\new_[3965]_  & (~\new_[20317]_  | ~\wbm_dat_o[29] );
  assign \new_[3911]_  = ~\new_[3966]_  & (~\new_[20317]_  | ~\wbm_dat_o[2] );
  assign \new_[3912]_  = ~\new_[3967]_  & (~\new_[20317]_  | ~\wbm_dat_o[30] );
  assign \new_[3913]_  = ~\new_[3968]_  & (~\new_[20317]_  | ~\wbm_dat_o[31] );
  assign \new_[3914]_  = ~\new_[3969]_  & (~\new_[5299]_  | ~\wbm_dat_o[3] );
  assign \new_[3915]_  = ~\new_[3970]_  & (~\new_[5299]_  | ~\wbm_dat_o[4] );
  assign \new_[3916]_  = ~\new_[3971]_  & (~\new_[5299]_  | ~\wbm_dat_o[5] );
  assign \new_[3917]_  = ~\new_[3972]_  & (~\new_[5299]_  | ~\wbm_dat_o[6] );
  assign \new_[3918]_  = ~\new_[3973]_  & (~\new_[20317]_  | ~\wbm_dat_o[8] );
  assign \new_[3919]_  = ~\new_[3974]_  & (~\new_[5299]_  | ~\wbm_dat_o[9] );
  assign n1095 = ~\new_[4005]_  & ~\new_[5443]_ ;
  assign \new_[3921]_  = ~\new_[4004]_  & ~\new_[4040]_ ;
  assign \new_[3922]_  = ~\new_[3997]_  & (~\new_[5299]_  | ~\wbm_dat_o[15] );
  assign \new_[3923]_  = ~\new_[3998]_  & (~\new_[20317]_  | ~\wbm_dat_o[18] );
  assign \new_[3924]_  = ~\new_[3999]_  & (~\new_[20317]_  | ~\wbm_dat_o[7] );
  assign \new_[3925]_  = ~\new_[4000]_  & (~\new_[20317]_  | ~\wbm_sel_o[0] );
  assign \new_[3926]_  = ~\new_[4001]_  & (~\new_[20317]_  | ~\wbm_sel_o[1] );
  assign \new_[3927]_  = ~\new_[4002]_  & (~\new_[20317]_  | ~\wbm_sel_o[2] );
  assign \new_[3928]_  = ~\new_[4003]_  & (~\new_[20317]_  | ~\wbm_sel_o[3] );
  assign \new_[3929]_  = \new_[15161]_  ? \new_[20499]_  : \new_[4059]_ ;
  assign \new_[3930]_  = \new_[15188]_  ? \new_[20499]_  : \new_[4060]_ ;
  assign \new_[3931]_  = \new_[15187]_  ? \new_[20499]_  : \new_[4061]_ ;
  assign \new_[3932]_  = \new_[15186]_  ? \new_[20499]_  : \new_[4062]_ ;
  assign \new_[3933]_  = \new_[15185]_  ? \new_[20499]_  : \new_[4063]_ ;
  assign \new_[3934]_  = \new_[15201]_  ? \new_[20499]_  : \new_[4064]_ ;
  assign \new_[3935]_  = \new_[15189]_  ? \new_[20498]_  : \new_[4065]_ ;
  assign \new_[3936]_  = \new_[15400]_  ? \new_[20498]_  : \new_[4066]_ ;
  assign \new_[3937]_  = \new_[15183]_  ? \new_[20498]_  : \new_[4067]_ ;
  assign \new_[3938]_  = \new_[15272]_  ? \new_[20498]_  : \new_[4068]_ ;
  assign \new_[3939]_  = \new_[15210]_  ? \new_[20498]_  : \new_[4069]_ ;
  assign \new_[3940]_  = \new_[15285]_  ? \new_[20499]_  : \new_[4075]_ ;
  assign \new_[3941]_  = \new_[15192]_  ? \new_[20498]_  : \new_[4076]_ ;
  assign \new_[3942]_  = \new_[15387]_  ? \new_[20499]_  : \new_[4077]_ ;
  assign \new_[3943]_  = \new_[15233]_  ? \new_[20498]_  : \new_[4079]_ ;
  assign \new_[3944]_  = pci_target_unit_pci_target_sm_backoff_reg;
  assign \new_[3945]_  = \new_[15284]_  ? \new_[20499]_  : \new_[4080]_ ;
  assign \new_[3946]_  = \new_[15204]_  ? \new_[20498]_  : \new_[4081]_ ;
  assign \new_[3947]_  = ~\new_[5416]_  & ~\new_[4010]_ ;
  assign \new_[3948]_  = ~\new_[5416]_  & ~\new_[4011]_ ;
  assign \new_[3949]_  = ~\new_[5416]_  & ~\new_[4012]_ ;
  assign \new_[3950]_  = ~\new_[5416]_  & ~\new_[4013]_ ;
  assign \new_[3951]_  = ~\new_[5416]_  & ~\new_[4014]_ ;
  assign \new_[3952]_  = ~\new_[5416]_  & ~\new_[4015]_ ;
  assign \new_[3953]_  = ~\new_[5416]_  & ~\new_[4016]_ ;
  assign \new_[3954]_  = ~\new_[5416]_  & ~\new_[4017]_ ;
  assign \new_[3955]_  = ~\new_[5416]_  & ~\new_[4018]_ ;
  assign \new_[3956]_  = ~\new_[5416]_  & ~\new_[4019]_ ;
  assign \new_[3957]_  = ~\new_[5416]_  & ~\new_[4020]_ ;
  assign \new_[3958]_  = ~\new_[5416]_  & ~\new_[4021]_ ;
  assign \new_[3959]_  = ~\new_[5416]_  & ~\new_[4023]_ ;
  assign \new_[3960]_  = ~\new_[5416]_  & ~\new_[4024]_ ;
  assign \new_[3961]_  = ~\new_[5416]_  & ~\new_[4025]_ ;
  assign \new_[3962]_  = ~\new_[5416]_  & ~\new_[4026]_ ;
  assign \new_[3963]_  = ~\new_[5416]_  & ~\new_[4027]_ ;
  assign \new_[3964]_  = ~\new_[5416]_  & ~\new_[4028]_ ;
  assign \new_[3965]_  = ~\new_[5416]_  & ~\new_[4029]_ ;
  assign \new_[3966]_  = ~\new_[5416]_  & ~\new_[4030]_ ;
  assign \new_[3967]_  = ~\new_[5416]_  & ~\new_[4031]_ ;
  assign \new_[3968]_  = ~\new_[5416]_  & ~\new_[4032]_ ;
  assign \new_[3969]_  = ~\new_[5416]_  & ~\new_[4033]_ ;
  assign \new_[3970]_  = ~\new_[5416]_  & ~\new_[4034]_ ;
  assign \new_[3971]_  = ~\new_[5416]_  & ~\new_[4035]_ ;
  assign \new_[3972]_  = ~\new_[5416]_  & ~\new_[4036]_ ;
  assign \new_[3973]_  = ~\new_[5416]_  & ~\new_[4037]_ ;
  assign \new_[3974]_  = ~\new_[5416]_  & ~\new_[4038]_ ;
  assign n1120 = ~\new_[15841]_  & (~\new_[16899]_  | ~\new_[4074]_ );
  assign \new_[3976]_  = ~\new_[4074]_  | ~\new_[5886]_  | ~\new_[19874]_ ;
  assign \new_[3977]_  = (~\new_[17348]_  | ~\new_[9614]_ ) & (~\new_[9762]_  | ~\new_[4048]_ );
  assign \new_[3978]_  = (~\new_[17358]_  | ~\new_[9614]_ ) & (~\new_[9762]_  | ~\new_[4056]_ );
  assign n1100 = \new_[18909]_  ? n6835 : \new_[4070]_ ;
  assign n1105 = \new_[19219]_  ? n6835 : \new_[4071]_ ;
  assign n1110 = \new_[19116]_  ? n6835 : \new_[4072]_ ;
  assign n1115 = \new_[19573]_  ? n6835 : \new_[4073]_ ;
  assign \new_[3983]_  = \new_[15329]_  ? \new_[20498]_  : \new_[4045]_ ;
  assign \new_[3984]_  = \new_[15236]_  ? \new_[20499]_  : \new_[4046]_ ;
  assign \new_[3985]_  = \new_[15309]_  ? \new_[20499]_  : \new_[4047]_ ;
  assign \new_[3986]_  = \new_[15300]_  ? \new_[20499]_  : \new_[4049]_ ;
  assign \new_[3987]_  = \new_[15232]_  ? \new_[20499]_  : \new_[4052]_ ;
  assign \new_[3988]_  = \new_[15170]_  ? \new_[20499]_  : \new_[4051]_ ;
  assign \new_[3989]_  = \new_[15406]_  ? \new_[20499]_  : \new_[4053]_ ;
  assign \new_[3990]_  = \new_[15268]_  ? \new_[20498]_  : \new_[4055]_ ;
  assign \new_[3991]_  = \new_[15190]_  ? \new_[20499]_  : \new_[4057]_ ;
  assign \new_[3992]_  = \new_[15163]_  ? \new_[20499]_  : \new_[4058]_ ;
  assign \new_[3993]_  = \new_[15194]_  ? \new_[20498]_  : \new_[4090]_ ;
  assign \new_[3994]_  = ~wishbone_slave_unit_del_sync_req_done_reg_reg;
  assign \new_[3995]_  = \\wishbone_slave_unit_wishbone_slave_c_state_reg[0] ;
  assign \wbm_cti_o[1]  = \\pci_target_unit_wishbone_master_wb_cti_o_reg[1] ;
  assign \new_[3997]_  = ~\new_[5416]_  & ~\new_[4050]_ ;
  assign \new_[3998]_  = ~\new_[5416]_  & ~\new_[4054]_ ;
  assign \new_[3999]_  = ~\new_[5416]_  & ~\new_[4078]_ ;
  assign \new_[4000]_  = ~\new_[20317]_  & ~\new_[4070]_ ;
  assign \new_[4001]_  = ~\new_[20317]_  & ~\new_[4071]_ ;
  assign \new_[4002]_  = ~\new_[20317]_  & ~\new_[4072]_ ;
  assign \new_[4003]_  = ~\new_[20317]_  & ~\new_[4073]_ ;
  assign \new_[4004]_  = ~\new_[4074]_  | (~\new_[16591]_  & ~\new_[17008]_ );
  assign \new_[4005]_  = ~\new_[4082]_  & (~\new_[4762]_  | ~\new_[4095]_ );
  assign \new_[4006]_  = \new_[15270]_  ? \new_[20498]_  : \new_[4088]_ ;
  assign \new_[4007]_  = \new_[15401]_  ? \new_[20499]_  : \new_[4089]_ ;
  assign \new_[4008]_  = wishbone_slave_unit_del_sync_req_comp_pending_reg;
  assign \new_[4009]_  = \\wishbone_slave_unit_wishbone_slave_c_state_reg[2] ;
  assign \new_[4010]_  = ~\new_[4048]_ ;
  assign \new_[4011]_  = ~\new_[4045]_ ;
  assign \new_[4012]_  = ~\new_[4046]_ ;
  assign \new_[4013]_  = ~\new_[4047]_ ;
  assign \new_[4014]_  = ~\new_[4049]_ ;
  assign \new_[4015]_  = ~\new_[4052]_ ;
  assign \new_[4016]_  = ~\new_[4051]_ ;
  assign \new_[4017]_  = ~\new_[4053]_ ;
  assign \new_[4018]_  = ~\new_[4055]_ ;
  assign \new_[4019]_  = ~\new_[4056]_ ;
  assign \new_[4020]_  = ~\new_[4057]_ ;
  assign \new_[4021]_  = ~\new_[4058]_ ;
  assign \new_[4022]_  = ~\new_[4059]_ ;
  assign \new_[4023]_  = ~\new_[4060]_ ;
  assign \new_[4024]_  = ~\new_[4061]_ ;
  assign \new_[4025]_  = ~\new_[4062]_ ;
  assign \new_[4026]_  = ~\new_[4063]_ ;
  assign \new_[4027]_  = ~\new_[4064]_ ;
  assign \new_[4028]_  = ~\new_[4065]_ ;
  assign \new_[4029]_  = ~\new_[4066]_ ;
  assign \new_[4030]_  = ~\new_[4067]_ ;
  assign \new_[4031]_  = ~\new_[4068]_ ;
  assign \new_[4032]_  = ~\new_[4069]_ ;
  assign \new_[4033]_  = ~\new_[4075]_ ;
  assign \new_[4034]_  = ~\new_[4076]_ ;
  assign \new_[4035]_  = ~\new_[4077]_ ;
  assign \new_[4036]_  = ~\new_[4079]_ ;
  assign \new_[4037]_  = ~\new_[4080]_ ;
  assign \new_[4038]_  = ~\new_[4081]_ ;
  assign n1125 = ~\new_[4407]_  | (~\new_[4122]_  & ~\new_[16800]_ );
  assign \new_[4040]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36] ;
  assign \new_[4041]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[38] ;
  assign \new_[4042]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39] ;
  assign n1140 = ~\new_[4240]_  | ~\new_[4096]_ ;
  assign n1135 = ~\new_[13804]_  | ~\new_[4276]_  | ~\new_[4134]_ ;
  assign \new_[4045]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[10] ;
  assign \new_[4046]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[11] ;
  assign \new_[4047]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[12] ;
  assign \new_[4048]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[0] ;
  assign \new_[4049]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[13] ;
  assign \new_[4050]_  = ~\new_[4088]_ ;
  assign \new_[4051]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[16] ;
  assign \new_[4052]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[14] ;
  assign \new_[4053]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[17] ;
  assign \new_[4054]_  = ~\new_[4089]_ ;
  assign \new_[4055]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[19] ;
  assign \new_[4056]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[1] ;
  assign \new_[4057]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[20] ;
  assign \new_[4058]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[21] ;
  assign \new_[4059]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[22] ;
  assign \new_[4060]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[23] ;
  assign \new_[4061]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[24] ;
  assign \new_[4062]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[25] ;
  assign \new_[4063]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[26] ;
  assign \new_[4064]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[27] ;
  assign \new_[4065]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[28] ;
  assign \new_[4066]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[29] ;
  assign \new_[4067]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[2] ;
  assign \new_[4068]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[30] ;
  assign \new_[4069]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[31] ;
  assign \new_[4070]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[32] ;
  assign \new_[4071]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[33] ;
  assign \new_[4072]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[34] ;
  assign \new_[4073]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[35] ;
  assign \new_[4074]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[37] ;
  assign \new_[4075]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[3] ;
  assign \new_[4076]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[4] ;
  assign \new_[4077]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[5] ;
  assign \new_[4078]_  = ~\new_[4090]_ ;
  assign \new_[4079]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[6] ;
  assign \new_[4080]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[8] ;
  assign \new_[4081]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[9] ;
  assign \new_[4082]_  = ~pci_perr_i & ~\new_[4095]_ ;
  assign n1130 = ~\new_[16778]_  & (~\new_[4133]_  | ~\new_[3994]_ );
  assign \new_[4084]_  = ~output_backup_trdy_out_reg;
  assign pci_trdy_o = pci_io_mux_trdy_iob_dat_out_reg;
  assign n1145 = \new_[16598]_  & \new_[4133]_ ;
  assign n1150 = ~\new_[11173]_  | ~\new_[4236]_  | ~\new_[13814]_  | ~\new_[4276]_ ;
  assign \new_[4088]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[15] ;
  assign \new_[4089]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[18] ;
  assign \new_[4090]_  = \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[7] ;
  assign pci_stop_o = pci_io_mux_stop_iob_dat_out_reg;
  assign \new_[4092]_  = ~output_backup_stop_out_reg;
  assign pci_devsel_o = pci_io_mux_devsel_iob_dat_out_reg;
  assign \new_[4094]_  = ~output_backup_devsel_out_reg;
  assign \new_[4095]_  = output_backup_perr_en_out_reg;
  assign \new_[4096]_  = ~\new_[4141]_  & (~\new_[5412]_  | ~\new_[5465]_ );
  assign n1170 = ~\new_[4282]_  | ~\new_[4143]_  | ~\new_[4416]_ ;
  assign n1185 = ~\new_[4280]_  | ~\new_[4142]_  | ~\new_[4414]_ ;
  assign n1175 = ~\new_[4419]_  | ~\new_[4144]_  | ~\new_[4418]_ ;
  assign n1180 = ~\new_[4285]_  | ~\new_[4145]_  | ~\new_[4421]_ ;
  assign n1190 = ~\new_[4287]_  | ~\new_[4146]_  | ~\new_[4423]_ ;
  assign n1200 = ~\new_[4289]_  | ~\new_[4147]_  | ~\new_[4425]_ ;
  assign n1195 = ~\new_[4291]_  | ~\new_[4148]_  | ~\new_[4426]_ ;
  assign n1205 = ~\new_[4149]_  | ~\new_[4293]_  | ~\new_[4429]_ ;
  assign n1215 = ~\new_[4432]_  | ~\new_[4150]_  | ~\new_[4431]_ ;
  assign n1220 = ~\new_[4296]_  | ~\new_[4151]_  | ~\new_[4434]_ ;
  assign n1225 = ~\new_[4436]_  | ~\new_[4152]_  | ~\new_[4435]_ ;
  assign n1230 = ~\new_[4438]_  | ~\new_[4153]_  | ~\new_[4300]_ ;
  assign n1235 = ~\new_[4440]_  | ~\new_[4154]_  | ~\new_[4302]_ ;
  assign n1245 = ~\new_[4304]_  | ~\new_[4155]_  | ~\new_[4442]_ ;
  assign n1250 = ~\new_[4444]_  | ~\new_[4443]_  | ~\new_[4156]_ ;
  assign n1255 = ~\new_[4308]_  | ~\new_[4446]_  | ~\new_[4157]_ ;
  assign n1260 = ~\new_[4448]_  | ~\new_[4158]_  | ~\new_[4447]_ ;
  assign n1265 = ~\new_[4312]_  | ~\new_[4159]_  | ~\new_[4450]_ ;
  assign n1270 = ~\new_[4452]_  | ~\new_[4160]_  | ~\new_[4314]_ ;
  assign n1275 = ~\new_[4454]_  | ~\new_[4161]_  | ~\new_[4316]_ ;
  assign n1280 = ~\new_[4319]_  | ~\new_[4162]_  | ~\new_[4455]_ ;
  assign n1285 = ~\new_[4321]_  | ~\new_[4163]_  | ~\new_[4242]_ ;
  assign n1290 = ~\new_[4244]_  | ~\new_[4164]_  | ~\new_[4323]_ ;
  assign n1295 = ~\new_[4325]_  | ~\new_[4165]_  | ~\new_[4246]_ ;
  assign n1300 = ~\new_[4328]_  | ~\new_[4166]_  | ~\new_[4327]_ ;
  assign \new_[4122]_  = ~\new_[3944]_  & (~\new_[4234]_  | ~\new_[17113]_ );
  assign n1305 = ~\new_[4331]_  | ~\new_[4167]_  | ~\new_[4330]_ ;
  assign n1165 = ~\new_[4168]_  | ~\new_[4237]_ ;
  assign n1310 = ~\new_[4169]_  | ~\new_[4253]_  | ~\new_[4336]_ ;
  assign n1320 = ~\new_[4255]_  | ~\new_[4170]_  | ~\new_[4338]_ ;
  assign n1325 = ~\new_[4257]_  | ~\new_[4171]_  | ~\new_[4340]_ ;
  assign n1330 = ~\new_[4259]_  | ~\new_[4172]_  | ~\new_[4342]_ ;
  assign n1335 = ~\new_[4173]_  | ~\new_[4270]_  | ~\new_[4346]_ ;
  assign \new_[4130]_  = \\output_backup_ad_out_reg[31] ;
  assign \pci_ad_o[31]  = pci_io_mux_ad_iob31_dat_out_reg;
  assign pci_perr_oe_o = pci_io_mux_perr_iob_en_out_reg;
  assign \new_[4133]_  = ~\new_[4235]_  & ~n16770;
  assign \new_[4134]_  = ~\new_[4238]_  | ~\new_[20398]_ ;
  assign n1345 = ~\new_[4230]_  & (~\new_[16071]_  | ~\new_[16889]_ );
  assign \new_[4136]_  = \\configuration_status_bit15_11_reg[15] ;
  assign \new_[4137]_  = ~wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg;
  assign n1370 = ~\new_[4275]_  & (~\new_[4760]_  | ~\new_[15935]_ );
  assign n1380 = \new_[4610]_  & \new_[4274]_ ;
  assign n1385 = ~n1400;
  assign \new_[4141]_  = ~\new_[5465]_  & (~\new_[4412]_  | ~\new_[18488]_ );
  assign \new_[4142]_  = ~\new_[4413]_  & ~\new_[4279]_ ;
  assign \new_[4143]_  = ~\new_[4281]_  & ~\new_[4415]_ ;
  assign \new_[4144]_  = ~\new_[4417]_  & ~\new_[4283]_ ;
  assign \new_[4145]_  = ~\new_[4284]_  & ~\new_[4420]_ ;
  assign \new_[4146]_  = ~\new_[4286]_  & ~\new_[4422]_ ;
  assign \new_[4147]_  = ~\new_[4288]_  & ~\new_[4424]_ ;
  assign \new_[4148]_  = ~\new_[4290]_  & ~\new_[4427]_ ;
  assign \new_[4149]_  = ~\new_[4428]_  & ~\new_[4292]_ ;
  assign \new_[4150]_  = ~\new_[4430]_  & ~\new_[4294]_ ;
  assign \new_[4151]_  = ~\new_[4295]_  & ~\new_[4433]_ ;
  assign \new_[4152]_  = ~\new_[4297]_  & ~\new_[4298]_ ;
  assign \new_[4153]_  = ~\new_[4299]_  & ~\new_[4437]_ ;
  assign \new_[4154]_  = ~\new_[4301]_  & ~\new_[4439]_ ;
  assign \new_[4155]_  = ~\new_[4303]_  & ~\new_[4441]_ ;
  assign \new_[4156]_  = ~\new_[4305]_  & ~\new_[4306]_ ;
  assign \new_[4157]_  = ~\new_[4307]_  & ~\new_[4445]_ ;
  assign \new_[4158]_  = ~\new_[4309]_  & ~\new_[4310]_ ;
  assign \new_[4159]_  = ~\new_[4311]_  & ~\new_[4449]_ ;
  assign \new_[4160]_  = ~\new_[4313]_  & ~\new_[4451]_ ;
  assign \new_[4161]_  = ~\new_[4453]_  & ~\new_[4315]_ ;
  assign \new_[4162]_  = ~\new_[4317]_  & ~\new_[4318]_ ;
  assign \new_[4163]_  = ~\new_[4241]_  & ~\new_[4320]_ ;
  assign \new_[4164]_  = ~\new_[4243]_  & ~\new_[4322]_ ;
  assign \new_[4165]_  = ~\new_[4245]_  & ~\new_[4324]_ ;
  assign \new_[4166]_  = ~\new_[4247]_  & ~\new_[4326]_ ;
  assign \new_[4167]_  = ~\new_[4248]_  & ~\new_[4329]_ ;
  assign \new_[4168]_  = ~\new_[4250]_  & ~\new_[4251]_ ;
  assign \new_[4169]_  = ~\new_[4335]_  & ~\new_[4252]_ ;
  assign \new_[4170]_  = ~\new_[4337]_  & ~\new_[4254]_ ;
  assign \new_[4171]_  = ~\new_[4256]_  & ~\new_[4339]_ ;
  assign \new_[4172]_  = ~\new_[4341]_  & ~\new_[4258]_ ;
  assign \new_[4173]_  = ~\new_[4343]_  & ~\new_[4264]_ ;
  assign \new_[4174]_  = \\output_backup_cbe_out_reg[0] ;
  assign \new_[4175]_  = \\output_backup_cbe_out_reg[3] ;
  assign \pci_cbe_o[0]  = pci_io_mux_cbe_iob0_dat_out_reg;
  assign \pci_cbe_o[2]  = pci_io_mux_cbe_iob2_dat_out_reg;
  assign \new_[4178]_  = \\output_backup_cbe_out_reg[2] ;
  assign \pci_cbe_o[3]  = pci_io_mux_cbe_iob3_dat_out_reg;
  assign \new_[4180]_  = \\output_backup_ad_out_reg[15] ;
  assign \new_[4181]_  = \\output_backup_ad_out_reg[23] ;
  assign \new_[4182]_  = \\output_backup_ad_out_reg[24] ;
  assign \new_[4183]_  = \\output_backup_ad_out_reg[27] ;
  assign \new_[4184]_  = \\output_backup_ad_out_reg[28] ;
  assign \new_[4185]_  = \\output_backup_ad_out_reg[29] ;
  assign \new_[4186]_  = \\output_backup_ad_out_reg[2] ;
  assign \new_[4187]_  = \\output_backup_ad_out_reg[3] ;
  assign \new_[4188]_  = \\output_backup_ad_out_reg[4] ;
  assign \new_[4189]_  = \\output_backup_ad_out_reg[5] ;
  assign \new_[4190]_  = \\output_backup_ad_out_reg[6] ;
  assign \new_[4191]_  = \\output_backup_ad_out_reg[7] ;
  assign \new_[4192]_  = \\output_backup_ad_out_reg[8] ;
  assign \pci_ad_o[11]  = pci_io_mux_ad_iob11_dat_out_reg;
  assign \pci_ad_o[12]  = pci_io_mux_ad_iob12_dat_out_reg;
  assign \pci_ad_o[13]  = pci_io_mux_ad_iob13_dat_out_reg;
  assign \pci_ad_o[14]  = pci_io_mux_ad_iob14_dat_out_reg;
  assign \pci_ad_o[15]  = pci_io_mux_ad_iob15_dat_out_reg;
  assign \pci_ad_o[24]  = pci_io_mux_ad_iob24_dat_out_reg;
  assign \pci_ad_o[27]  = pci_io_mux_ad_iob27_dat_out_reg;
  assign \pci_ad_o[29]  = pci_io_mux_ad_iob29_dat_out_reg;
  assign \pci_ad_o[28]  = pci_io_mux_ad_iob28_dat_out_reg;
  assign \pci_ad_o[2]  = pci_io_mux_ad_iob2_dat_out_reg;
  assign \pci_ad_o[4]  = pci_io_mux_ad_iob4_dat_out_reg;
  assign \pci_ad_o[5]  = pci_io_mux_ad_iob5_dat_out_reg;
  assign \pci_ad_o[6]  = pci_io_mux_ad_iob6_dat_out_reg;
  assign \pci_ad_o[7]  = pci_io_mux_ad_iob7_dat_out_reg;
  assign \pci_ad_o[23]  = pci_io_mux_ad_iob23_dat_out_reg;
  assign \pci_ad_o[8]  = pci_io_mux_ad_iob8_dat_out_reg;
  assign \pci_ad_o[3]  = pci_io_mux_ad_iob3_dat_out_reg;
  assign \new_[4210]_  = \\output_backup_ad_out_reg[13] ;
  assign \new_[4211]_  = \\output_backup_ad_out_reg[14] ;
  assign \new_[4212]_  = \\output_backup_ad_out_reg[16] ;
  assign \new_[4213]_  = \\output_backup_ad_out_reg[17] ;
  assign \new_[4214]_  = \\output_backup_ad_out_reg[18] ;
  assign \new_[4215]_  = \\output_backup_ad_out_reg[19] ;
  assign \new_[4216]_  = \\output_backup_ad_out_reg[20] ;
  assign \new_[4217]_  = \\output_backup_ad_out_reg[22] ;
  assign \new_[4218]_  = \\output_backup_ad_out_reg[9] ;
  assign \pci_ad_o[10]  = pci_io_mux_ad_iob10_dat_out_reg;
  assign \pci_ad_o[16]  = pci_io_mux_ad_iob16_dat_out_reg;
  assign \pci_ad_o[17]  = pci_io_mux_ad_iob17_dat_out_reg;
  assign \pci_ad_o[18]  = pci_io_mux_ad_iob18_dat_out_reg;
  assign \pci_ad_o[19]  = pci_io_mux_ad_iob19_dat_out_reg;
  assign \pci_ad_o[22]  = pci_io_mux_ad_iob22_dat_out_reg;
  assign \pci_ad_o[20]  = pci_io_mux_ad_iob20_dat_out_reg;
  assign \new_[4226]_  = \\output_backup_ad_out_reg[10] ;
  assign \pci_ad_o[9]  = pci_io_mux_ad_iob9_dat_out_reg;
  assign \new_[4228]_  = \\output_backup_ad_out_reg[11] ;
  assign \new_[4229]_  = \\output_backup_ad_out_reg[12] ;
  assign \new_[4230]_  = ~\new_[4628]_  | ~\new_[4356]_  | ~\new_[4601]_ ;
  assign n1400 = ~n1750 & ~\new_[4354]_ ;
  assign n1390 = ~\new_[4272]_ ;
  assign n1395 = ~\new_[4273]_ ;
  assign \new_[4234]_  = ~\new_[4355]_  & (~\new_[6944]_  | ~\new_[16436]_ );
  assign \new_[4235]_  = ~\new_[4612]_  | (~\new_[4611]_  & ~\new_[19933]_ );
  assign \new_[4236]_  = ~\new_[4759]_  | ~\new_[20397]_  | ~\new_[20398]_  | ~\new_[20396]_ ;
  assign \new_[4237]_  = ~\new_[4333]_  & ~\new_[4334]_ ;
  assign \new_[4238]_  = ~\new_[11382]_  | ~\new_[4347]_ ;
  assign \new_[4239]_  = \new_[4411]_  | \new_[5412]_ ;
  assign \new_[4240]_  = \new_[4408]_  | \new_[5412]_ ;
  assign \new_[4241]_  = ~\new_[4576]_  | ~\new_[4577]_ ;
  assign \new_[4242]_  = \new_[4506]_  & \new_[4507]_ ;
  assign \new_[4243]_  = ~\new_[4578]_  | ~\new_[4579]_ ;
  assign \new_[4244]_  = \new_[4508]_  & \new_[4661]_ ;
  assign \new_[4245]_  = ~\new_[4580]_  | ~\new_[4581]_ ;
  assign \new_[4246]_  = \new_[4509]_  & \new_[4510]_ ;
  assign \new_[4247]_  = ~\new_[4511]_  | ~\new_[4512]_ ;
  assign \new_[4248]_  = ~\new_[4515]_  | ~\new_[4516]_ ;
  assign \new_[4249]_  = ~\new_[4517]_  | ~\new_[4518]_ ;
  assign \new_[4250]_  = ~\new_[4583]_  | ~\new_[4585]_ ;
  assign \new_[4251]_  = ~\new_[4520]_  | ~\new_[4519]_ ;
  assign \new_[4252]_  = ~\new_[4587]_  | ~\new_[4586]_ ;
  assign \new_[4253]_  = \new_[4521]_  & \new_[4522]_ ;
  assign \new_[4254]_  = ~\new_[4525]_  | ~\new_[4671]_ ;
  assign \new_[4255]_  = \new_[4590]_  & \new_[4591]_ ;
  assign \new_[4256]_  = ~\new_[4526]_  | ~\new_[4527]_ ;
  assign \new_[4257]_  = \new_[4592]_  & \new_[4593]_ ;
  assign \new_[4258]_  = ~\new_[4531]_  | ~\new_[4530]_ ;
  assign \new_[4259]_  = \new_[4596]_  & \new_[4597]_ ;
  assign \new_[4260]_  = \\output_backup_ad_out_reg[1] ;
  assign \new_[4261]_  = \\output_backup_ad_out_reg[30] ;
  assign \pci_ad_o[1]  = pci_io_mux_ad_iob1_dat_out_reg;
  assign \pci_ad_o[30]  = pci_io_mux_ad_iob30_dat_out_reg;
  assign \new_[4264]_  = ~\new_[4599]_  | ~\new_[4598]_ ;
  assign \new_[4265]_  = \\output_backup_ad_out_reg[21] ;
  assign \pci_ad_o[21]  = pci_io_mux_ad_iob21_dat_out_reg;
  assign \new_[4267]_  = \\configuration_status_bit15_11_reg[14] ;
  assign \new_[4268]_  = \\output_backup_ad_out_reg[26] ;
  assign \pci_ad_o[26]  = pci_io_mux_ad_iob26_dat_out_reg;
  assign \new_[4270]_  = \new_[4532]_  & \new_[4533]_ ;
  assign n1405 = ~\new_[4763]_  | ~\new_[4606]_  | ~\new_[10924]_ ;
  assign \new_[4272]_  = ~\new_[4582]_  & (~\new_[12487]_  | ~\new_[4130]_ );
  assign \new_[4273]_  = ~\new_[4582]_  & (~\new_[12487]_  | ~\pci_ad_o[31] );
  assign \new_[4274]_  = ~\new_[4856]_  & ~\new_[4609]_ ;
  assign \new_[4275]_  = ~\new_[15940]_  | ~\new_[4854]_  | ~\new_[15057]_  | ~\new_[10962]_ ;
  assign \new_[4276]_  = ~\new_[4611]_  | ~\new_[16672]_ ;
  assign n1410 = ~\new_[13714]_  & ~\new_[4611]_ ;
  assign \new_[4278]_  = ~\new_[4412]_ ;
  assign \new_[4279]_  = ~\new_[4534]_  | ~\new_[4535]_ ;
  assign \new_[4280]_  = \new_[4461]_  & \new_[4462]_ ;
  assign \new_[4281]_  = ~\new_[4463]_  | ~\new_[4464]_ ;
  assign \new_[4282]_  = \new_[4536]_  & \new_[4537]_ ;
  assign \new_[4283]_  = ~\new_[4466]_  | ~\new_[4465]_ ;
  assign \new_[4284]_  = ~\new_[4538]_  | ~\new_[4539]_ ;
  assign \new_[4285]_  = \new_[4468]_  & \new_[4467]_ ;
  assign \new_[4286]_  = ~\new_[4540]_  | ~\new_[4541]_ ;
  assign \new_[4287]_  = \new_[4469]_  & \new_[4634]_ ;
  assign \new_[4288]_  = ~\new_[4542]_  | ~\new_[4543]_ ;
  assign \new_[4289]_  = \new_[4470]_  & \new_[4471]_ ;
  assign \new_[4290]_  = ~\new_[4544]_  | ~\new_[4545]_ ;
  assign \new_[4291]_  = \new_[4475]_  & \new_[4474]_ ;
  assign \new_[4292]_  = ~\new_[4546]_  | ~\new_[4547]_ ;
  assign \new_[4293]_  = \new_[4476]_  & \new_[4477]_ ;
  assign \new_[4294]_  = ~\new_[4481]_  | ~\new_[4482]_ ;
  assign \new_[4295]_  = ~\new_[4550]_  | ~\new_[4551]_ ;
  assign \new_[4296]_  = \new_[4483]_  & \new_[4644]_ ;
  assign \new_[4297]_  = ~\new_[4552]_  | ~\new_[4553]_ ;
  assign \new_[4298]_  = ~\new_[4484]_  | ~\new_[4645]_ ;
  assign \new_[4299]_  = ~\new_[4554]_  | ~\new_[4555]_ ;
  assign \new_[4300]_  = \new_[4485]_  & \new_[4486]_ ;
  assign \new_[4301]_  = ~\new_[4556]_  | ~\new_[4557]_ ;
  assign \new_[4302]_  = \new_[4487]_  & \new_[4488]_ ;
  assign \new_[4303]_  = ~\new_[4560]_  | ~\new_[4561]_ ;
  assign \new_[4304]_  = \new_[4492]_  & \new_[4491]_ ;
  assign \new_[4305]_  = ~\new_[4493]_  | ~\new_[4494]_ ;
  assign \new_[4306]_  = ~\new_[4562]_  | ~\new_[4563]_ ;
  assign \new_[4307]_  = ~\new_[4495]_  | ~\new_[4496]_ ;
  assign \new_[4308]_  = \new_[4564]_  & \new_[4565]_ ;
  assign \new_[4309]_  = ~\new_[4497]_  | ~\new_[4498]_ ;
  assign \new_[4310]_  = ~\new_[4567]_  | ~\new_[4566]_ ;
  assign \new_[4311]_  = ~\new_[4568]_  | ~\new_[4569]_ ;
  assign \new_[4312]_  = \new_[4499]_  & \new_[4655]_ ;
  assign \new_[4313]_  = ~\new_[4570]_  | ~\new_[4571]_ ;
  assign \new_[4314]_  = \new_[4500]_  & \new_[4501]_ ;
  assign \new_[4315]_  = ~\new_[4573]_  | ~\new_[4572]_ ;
  assign \new_[4316]_  = \new_[4502]_  & \new_[4503]_ ;
  assign \new_[4317]_  = ~\new_[4574]_  | ~\new_[4575]_ ;
  assign \new_[4318]_  = ~\new_[4504]_  | ~\new_[4505]_ ;
  assign \new_[4319]_  = \new_[4822]_  & \new_[4658]_ ;
  assign \new_[4320]_  = ~\new_[4823]_  | ~\new_[4659]_ ;
  assign \new_[4321]_  = \new_[4726]_  & \new_[4847]_ ;
  assign \new_[4322]_  = ~\new_[4728]_  | ~\new_[4727]_ ;
  assign \new_[4323]_  = \new_[4660]_  & \new_[4824]_ ;
  assign \new_[4324]_  = ~\new_[4730]_  | ~\new_[4729]_ ;
  assign \new_[4325]_  = \new_[4825]_  & \new_[4662]_ ;
  assign \new_[4326]_  = ~\new_[4826]_  | ~\new_[4663]_ ;
  assign \new_[4327]_  = \new_[4731]_  & \new_[4733]_ ;
  assign \new_[4328]_  = \new_[4732]_  & \new_[4734]_ ;
  assign \new_[4329]_  = ~\new_[4738]_  | ~\new_[4739]_ ;
  assign \new_[4330]_  = \new_[4740]_  & \new_[4741]_ ;
  assign \new_[4331]_  = \new_[4828]_  & \new_[4665]_ ;
  assign \new_[4332]_  = ~\new_[4742]_  | ~\new_[4849]_ ;
  assign \new_[4333]_  = ~\new_[4830]_  | ~\new_[4667]_ ;
  assign \new_[4334]_  = ~\new_[4745]_  | ~\new_[4746]_ ;
  assign \new_[4335]_  = ~\new_[4831]_  | ~\new_[4668]_ ;
  assign \new_[4336]_  = \new_[4747]_  & \new_[4748]_ ;
  assign \new_[4337]_  = ~\new_[4833]_  | ~\new_[4670]_ ;
  assign \new_[4338]_  = \new_[4751]_  & \new_[4850]_ ;
  assign \new_[4339]_  = ~\new_[4834]_  | ~\new_[4672]_ ;
  assign \new_[4340]_  = \new_[4752]_  & \new_[4851]_ ;
  assign \new_[4341]_  = ~\new_[4836]_  | ~\new_[4674]_ ;
  assign \new_[4342]_  = \new_[4757]_  & \new_[4852]_ ;
  assign \new_[4343]_  = ~\new_[4837]_  | ~\new_[4675]_ ;
  assign \pci_ad_o[0]  = pci_io_mux_ad_iob0_dat_out_reg;
  assign \new_[4345]_  = \\output_backup_ad_out_reg[0] ;
  assign \new_[4346]_  = \new_[4758]_  & \new_[4853]_ ;
  assign \new_[4347]_  = ~\new_[4903]_  | ~\new_[16400]_  | ~\new_[20397]_  | ~\new_[12571]_ ;
  assign n1415 = \new_[4871]_  ? \new_[12484]_  : \new_[4174]_ ;
  assign n1435 = \new_[4872]_  ? \new_[12484]_  : \new_[4178]_ ;
  assign n1420 = \new_[4873]_  ? \new_[12484]_  : \new_[4175]_ ;
  assign n1425 = \pci_cbe_o[0]  ? \new_[15613]_  : \new_[4871]_ ;
  assign n1430 = \pci_cbe_o[2]  ? \new_[15613]_  : \new_[4872]_ ;
  assign n1440 = \pci_cbe_o[3]  ? \new_[15613]_  : \new_[4873]_ ;
  assign \new_[4354]_  = parity_checker_perr_en_crit_gen_perr_en_reg_out_reg;
  assign \new_[4355]_  = ~\new_[4790]_  | ~\new_[16886]_ ;
  assign \new_[4356]_  = ~\new_[4584]_ ;
  assign n1605 = ~\new_[10975]_  | ~\new_[4782]_ ;
  assign n1610 = ~\new_[10976]_  | ~\new_[4783]_ ;
  assign n1615 = ~\new_[10977]_  | ~\new_[4784]_ ;
  assign n1620 = ~\new_[10978]_  | ~\new_[4785]_ ;
  assign n1625 = ~\new_[10980]_  | ~\new_[4786]_ ;
  assign n1630 = ~\new_[10983]_  | ~\new_[4787]_ ;
  assign n1450 = ~\new_[10984]_  | ~\new_[4764]_ ;
  assign n1455 = ~\new_[10985]_  | ~\new_[4765]_ ;
  assign n1460 = ~\new_[10988]_  | ~\new_[4766]_ ;
  assign n1465 = ~\new_[10989]_  | ~\new_[4767]_ ;
  assign n1470 = ~\new_[10990]_  | ~\new_[4768]_ ;
  assign n1475 = ~\new_[10991]_  | ~\new_[4769]_ ;
  assign n1480 = ~\new_[10993]_  | ~\new_[4770]_ ;
  assign n1485 = ~\new_[10994]_  | ~\new_[4771]_ ;
  assign n1490 = ~\new_[10995]_  | ~\new_[4772]_ ;
  assign n1495 = ~\new_[10996]_  | ~\new_[4773]_ ;
  assign n1500 = ~\new_[10997]_  | ~\new_[4774]_ ;
  assign n1505 = ~\new_[11155]_  | ~\new_[4775]_ ;
  assign n1635 = ~\new_[10998]_  | ~\new_[4788]_ ;
  assign n1640 = ~\new_[11006]_  | ~\new_[4792]_ ;
  assign n1510 = ~\new_[11172]_  | ~\new_[4777]_ ;
  assign n1515 = ~\new_[11176]_  | ~\new_[4781]_ ;
  assign n1520 = ~\new_[11160]_  | ~\new_[4778]_ ;
  assign n1525 = ~\new_[11161]_  | ~\new_[4779]_ ;
  assign n1530 = ~\new_[11162]_  | ~\new_[4780]_ ;
  assign n1645 = ~\new_[11013]_  | ~\new_[4782]_ ;
  assign n1650 = ~\new_[11163]_  | ~\new_[4783]_ ;
  assign n1655 = ~\new_[10999]_  | ~\new_[4784]_ ;
  assign n1660 = ~\new_[11000]_  | ~\new_[4785]_ ;
  assign n1670 = ~\new_[11158]_  | ~\new_[4786]_ ;
  assign n1665 = ~\new_[11166]_  | ~\new_[4787]_ ;
  assign n1535 = ~\new_[11167]_  | ~\new_[4765]_ ;
  assign n1540 = ~\new_[11002]_  | ~\new_[4766]_ ;
  assign n1580 = ~\new_[11157]_  | ~\new_[4764]_ ;
  assign n1545 = ~\new_[10981]_  | ~\new_[4768]_ ;
  assign n1550 = ~\new_[11003]_  | ~\new_[4767]_ ;
  assign n1555 = ~\new_[11153]_  | ~\new_[4769]_ ;
  assign n1590 = ~\new_[11169]_  | ~\new_[4770]_ ;
  assign n1560 = ~\new_[11152]_  | ~\new_[4771]_ ;
  assign n1565 = ~\new_[11151]_  | ~\new_[4772]_ ;
  assign n1570 = ~\new_[11170]_  | ~\new_[4773]_ ;
  assign n1575 = ~\new_[11004]_  | ~\new_[4774]_ ;
  assign n1585 = ~\new_[11171]_  | ~\new_[4775]_ ;
  assign n1680 = ~\new_[11005]_  | ~\new_[4788]_ ;
  assign n1675 = ~\new_[11008]_  | ~\new_[4792]_ ;
  assign n1690 = ~\new_[11010]_  | ~\new_[4781]_ ;
  assign n1685 = ~\new_[11009]_  | ~\new_[4777]_ ;
  assign n1595 = ~\new_[11011]_  | ~\new_[4778]_ ;
  assign n1600 = ~\new_[11012]_  | ~\new_[4779]_ ;
  assign n1445 = ~\new_[11014]_  | ~\new_[4780]_ ;
  assign \new_[4407]_  = ~\new_[10960]_  | ~\new_[16978]_  | ~\new_[4761]_  | ~\new_[16904]_ ;
  assign \new_[4408]_  = ~\new_[4676]_  & ~\wbm_cti_o[1] ;
  assign \new_[4409]_  = \new_[5368]_  | \new_[4676]_ ;
  assign \new_[4410]_  = \new_[5369]_  | \new_[4676]_ ;
  assign \new_[4411]_  = ~\new_[4676]_  | (~\new_[19873]_  & ~\new_[17455]_ );
  assign \new_[4412]_  = ~\new_[4676]_  & (~\new_[17247]_  | ~\new_[5161]_ );
  assign \new_[4413]_  = ~\new_[4798]_  | ~\new_[4629]_ ;
  assign \new_[4414]_  = \new_[4677]_  & \new_[4678]_ ;
  assign \new_[4415]_  = ~\new_[4680]_  | ~\new_[4679]_ ;
  assign \new_[4416]_  = \new_[4799]_  & \new_[4630]_ ;
  assign \new_[4417]_  = ~\new_[4800]_  | ~\new_[4631]_ ;
  assign \new_[4418]_  = \new_[4681]_  & \new_[4838]_ ;
  assign \new_[4419]_  = \new_[4682]_  & \new_[4683]_ ;
  assign \new_[4420]_  = ~\new_[4684]_  | ~\new_[4685]_ ;
  assign \new_[4421]_  = \new_[4632]_  & \new_[4801]_ ;
  assign \new_[4422]_  = ~\new_[4687]_  | ~\new_[4686]_ ;
  assign \new_[4423]_  = \new_[4633]_  & \new_[4802]_ ;
  assign \new_[4424]_  = ~\new_[4803]_  | ~\new_[4635]_ ;
  assign \new_[4425]_  = \new_[4688]_  & \new_[4839]_ ;
  assign \new_[4426]_  = \new_[4637]_  & \new_[4805]_ ;
  assign \new_[4427]_  = ~\new_[4693]_  | ~\new_[4694]_ ;
  assign \new_[4428]_  = ~\new_[4806]_  | ~\new_[4638]_ ;
  assign \new_[4429]_  = \new_[4695]_  & \new_[4696]_ ;
  assign \new_[4430]_  = ~\new_[4809]_  | ~\new_[4642]_ ;
  assign \new_[4431]_  = \new_[4703]_  & \new_[4840]_ ;
  assign \new_[4432]_  = \new_[4704]_  & \new_[4705]_ ;
  assign \new_[4433]_  = ~\new_[4706]_  | ~\new_[4707]_ ;
  assign \new_[4434]_  = \new_[4643]_  & \new_[4810]_ ;
  assign \new_[4435]_  = \new_[4646]_  & \new_[4811]_ ;
  assign \new_[4436]_  = \new_[4708]_  & \new_[4841]_ ;
  assign \new_[4437]_  = ~\new_[4710]_  | ~\new_[4709]_ ;
  assign \new_[4438]_  = \new_[4812]_  & \new_[4647]_ ;
  assign \new_[4439]_  = ~\new_[4813]_  | ~\new_[4648]_ ;
  assign \new_[4440]_  = \new_[4711]_  & \new_[4842]_ ;
  assign \new_[4441]_  = ~\new_[4815]_  | ~\new_[4650]_ ;
  assign \new_[4442]_  = \new_[4714]_  & \new_[4715]_ ;
  assign \new_[4443]_  = \new_[4816]_  & \new_[4651]_ ;
  assign \new_[4444]_  = \new_[4716]_  & \new_[4843]_ ;
  assign \new_[4445]_  = ~\new_[4718]_  | ~\new_[4717]_ ;
  assign \new_[4446]_  = \new_[4817]_  & \new_[4652]_ ;
  assign \new_[4447]_  = \new_[4818]_  & \new_[4653]_ ;
  assign \new_[4448]_  = \new_[4719]_  & \new_[4844]_ ;
  assign \new_[4449]_  = ~\new_[4721]_  | ~\new_[4720]_ ;
  assign \new_[4450]_  = \new_[4819]_  & \new_[4654]_ ;
  assign \new_[4451]_  = ~\new_[4723]_  | ~\new_[4722]_ ;
  assign \new_[4452]_  = \new_[4820]_  & \new_[4656]_ ;
  assign \new_[4453]_  = ~\new_[4821]_  | ~\new_[4657]_ ;
  assign \new_[4454]_  = \new_[4724]_  & \new_[4845]_ ;
  assign \new_[4455]_  = \new_[4725]_  & \new_[4846]_ ;
  assign \new_[4456]_  = \\output_backup_ad_out_reg[25] ;
  assign \pci_ad_o[25]  = pci_io_mux_ad_iob25_dat_out_reg;
  assign \new_[4458]_  = \\wishbone_slave_unit_pci_initiator_if_be_out_reg[0] ;
  assign \new_[4459]_  = \\wishbone_slave_unit_pci_initiator_if_be_out_reg[2] ;
  assign \new_[4460]_  = \\wishbone_slave_unit_pci_initiator_if_be_out_reg[3] ;
  assign \new_[4461]_  = ~\new_[4858]_  | ~\new_[18010]_ ;
  assign \new_[4462]_  = ~\new_[4860]_  | ~\new_[19153]_ ;
  assign \new_[4463]_  = ~\new_[4858]_  | ~\new_[18400]_ ;
  assign \new_[4464]_  = ~\new_[4861]_  | ~\new_[19384]_ ;
  assign \new_[4465]_  = ~\new_[4861]_  | ~\new_[18485]_ ;
  assign \new_[4466]_  = ~\new_[4858]_  | ~\new_[19550]_ ;
  assign \new_[4467]_  = ~\new_[4859]_  | ~\new_[18163]_ ;
  assign \new_[4468]_  = ~\new_[4862]_  | ~\new_[18764]_ ;
  assign \new_[4469]_  = ~\new_[4859]_  | ~\new_[19730]_ ;
  assign \new_[4470]_  = ~\new_[4858]_  | ~\new_[18712]_ ;
  assign \new_[4471]_  = ~\new_[4860]_  | ~\new_[19387]_ ;
  assign \new_[4472]_  = ~\new_[4859]_  | ~\new_[18418]_ ;
  assign \new_[4473]_  = ~\new_[4862]_  | ~\new_[18710]_ ;
  assign \new_[4474]_  = ~\new_[4859]_  | ~\new_[19397]_ ;
  assign \new_[4475]_  = ~\new_[4862]_  | ~\new_[18482]_ ;
  assign \new_[4476]_  = ~\new_[4859]_  | ~\new_[19356]_ ;
  assign \new_[4477]_  = ~\new_[4862]_  | ~\new_[19020]_ ;
  assign \new_[4478]_  = ~\new_[4859]_  | ~\new_[19706]_ ;
  assign \new_[4479]_  = ~\new_[4862]_  | ~\new_[18155]_ ;
  assign \new_[4480]_  = ~\new_[4858]_  | ~\new_[18432]_ ;
  assign \new_[4481]_  = ~\new_[4858]_  | ~\new_[18279]_ ;
  assign \new_[4482]_  = ~\new_[4861]_  | ~\new_[17996]_ ;
  assign \new_[4483]_  = ~\new_[4858]_  | ~\new_[19448]_ ;
  assign \new_[4484]_  = ~\new_[4858]_  | ~\new_[18433]_ ;
  assign \new_[4485]_  = ~\new_[4859]_  | ~\new_[18431]_ ;
  assign \new_[4486]_  = ~\new_[4862]_  | ~\new_[18493]_ ;
  assign \new_[4487]_  = ~\new_[4859]_  | ~\new_[18461]_ ;
  assign \new_[4488]_  = ~\new_[4862]_  | ~\new_[18494]_ ;
  assign \new_[4489]_  = ~\new_[4860]_  | ~\new_[18497]_ ;
  assign \new_[4490]_  = ~\new_[4858]_  | ~\new_[18235]_ ;
  assign \new_[4491]_  = ~\new_[4859]_  | ~\new_[18816]_ ;
  assign \new_[4492]_  = ~\new_[4862]_  | ~\new_[19496]_ ;
  assign \new_[4493]_  = ~\new_[4858]_  | ~\new_[18452]_ ;
  assign \new_[4494]_  = ~\new_[4861]_  | ~\new_[19734]_ ;
  assign \new_[4495]_  = ~\new_[4858]_  | ~\new_[19377]_ ;
  assign \new_[4496]_  = ~\new_[4860]_  | ~\new_[19076]_ ;
  assign \new_[4497]_  = ~\new_[4858]_  | ~\new_[19605]_ ;
  assign \new_[4498]_  = ~\new_[4861]_  | ~\new_[18785]_ ;
  assign \new_[4499]_  = ~\new_[4858]_  | ~\new_[18464]_ ;
  assign \new_[4500]_  = ~\new_[4859]_  | ~\new_[18477]_ ;
  assign \new_[4501]_  = ~\new_[4862]_  | ~\new_[18549]_ ;
  assign \new_[4502]_  = ~\new_[4859]_  | ~\new_[18466]_ ;
  assign \new_[4503]_  = ~\new_[4862]_  | ~\new_[19278]_ ;
  assign \new_[4504]_  = ~\new_[4858]_  | ~\new_[18255]_ ;
  assign \new_[4505]_  = ~\new_[4861]_  | ~\new_[18922]_ ;
  assign \new_[4506]_  = ~\new_[4859]_  | ~\new_[18703]_ ;
  assign \new_[4507]_  = ~\new_[4862]_  | ~\new_[17856]_ ;
  assign \new_[4508]_  = ~\new_[4858]_  | ~\new_[18465]_ ;
  assign \new_[4509]_  = ~\new_[4859]_  | ~\new_[18543]_ ;
  assign \new_[4510]_  = ~\new_[4862]_  | ~\new_[18527]_ ;
  assign \new_[4511]_  = ~\new_[4858]_  | ~\new_[18252]_ ;
  assign \new_[4512]_  = ~\new_[4861]_  | ~\new_[18706]_ ;
  assign \new_[4513]_  = ~\new_[4858]_  | ~\new_[18561]_ ;
  assign \new_[4514]_  = ~\new_[4860]_  | ~\new_[19284]_ ;
  assign \new_[4515]_  = ~\new_[4858]_  | ~\new_[19062]_ ;
  assign \new_[4516]_  = ~\new_[4860]_  | ~\new_[19071]_ ;
  assign \new_[4517]_  = ~\new_[4858]_  | ~\new_[18167]_ ;
  assign \new_[4518]_  = ~\new_[4860]_  | ~\new_[18709]_ ;
  assign \new_[4519]_  = ~\new_[4862]_  | ~\new_[18807]_ ;
  assign \new_[4520]_  = ~\new_[4859]_  | ~\new_[19274]_ ;
  assign \new_[4521]_  = ~\new_[4859]_  | ~\new_[19861]_ ;
  assign \new_[4522]_  = ~\new_[4862]_  | ~\new_[18800]_ ;
  assign \new_[4523]_  = ~\new_[4861]_  | ~\new_[18912]_ ;
  assign \new_[4524]_  = ~\new_[4858]_  | ~\new_[19385]_ ;
  assign \new_[4525]_  = ~\new_[4858]_  | ~\new_[19402]_ ;
  assign \new_[4526]_  = ~\new_[4858]_  | ~\new_[17953]_ ;
  assign \new_[4527]_  = ~\new_[4860]_  | ~\new_[18577]_ ;
  assign \new_[4528]_  = ~\new_[4859]_  | ~\new_[18626]_ ;
  assign \new_[4529]_  = ~\new_[4862]_  | ~\new_[18974]_ ;
  assign \new_[4530]_  = ~\new_[4860]_  | ~\new_[17861]_ ;
  assign \new_[4531]_  = ~\new_[4858]_  | ~\new_[18283]_ ;
  assign \new_[4532]_  = ~\new_[4858]_  | ~\new_[18708]_ ;
  assign \new_[4533]_  = ~\new_[4862]_  | ~\new_[19556]_ ;
  assign \new_[4534]_  = ~\new_[4864]_  | ~\new_[19096]_ ;
  assign \new_[4535]_  = ~\new_[4865]_  | ~\new_[18016]_ ;
  assign \new_[4536]_  = ~\new_[4864]_  | ~\new_[18913]_ ;
  assign \new_[4537]_  = ~\new_[4865]_  | ~\new_[18996]_ ;
  assign \new_[4538]_  = ~\new_[4863]_  | ~\new_[18778]_ ;
  assign \new_[4539]_  = ~\new_[4865]_  | ~\new_[17829]_ ;
  assign \new_[4540]_  = ~\new_[4863]_  | ~\new_[18651]_ ;
  assign \new_[4541]_  = ~\new_[4865]_  | ~\new_[19691]_ ;
  assign \new_[4542]_  = ~\new_[4863]_  | ~\new_[18498]_ ;
  assign \new_[4543]_  = ~\new_[4865]_  | ~\new_[19551]_ ;
  assign \new_[4544]_  = ~\new_[4863]_  | ~\new_[19744]_ ;
  assign \new_[4545]_  = ~\new_[4865]_  | ~\new_[18575]_ ;
  assign \new_[4546]_  = ~\new_[4865]_  | ~\new_[17871]_ ;
  assign \new_[4547]_  = ~\new_[4864]_  | ~\new_[19841]_ ;
  assign \new_[4548]_  = ~\new_[4864]_  | ~\new_[19769]_ ;
  assign \new_[4549]_  = ~\new_[4865]_  | ~\new_[19240]_ ;
  assign \new_[4550]_  = ~\new_[4863]_  | ~\new_[19039]_ ;
  assign \new_[4551]_  = ~\new_[4865]_  | ~\new_[19293]_ ;
  assign \new_[4552]_  = ~\new_[4863]_  | ~\new_[19102]_ ;
  assign \new_[4553]_  = ~\new_[4865]_  | ~\new_[18735]_ ;
  assign \new_[4554]_  = ~\new_[4863]_  | ~\new_[18172]_ ;
  assign \new_[4555]_  = ~\new_[4865]_  | ~\new_[19049]_ ;
  assign \new_[4556]_  = ~\new_[4863]_  | ~\new_[18210]_ ;
  assign \new_[4557]_  = ~\new_[4865]_  | ~\new_[19090]_ ;
  assign \new_[4558]_  = ~\new_[4864]_  | ~\new_[18430]_ ;
  assign \new_[4559]_  = ~\new_[4865]_  | ~\new_[17972]_ ;
  assign \new_[4560]_  = ~\new_[4863]_  | ~\new_[18760]_ ;
  assign \new_[4561]_  = ~\new_[4865]_  | ~\new_[19003]_ ;
  assign \new_[4562]_  = ~\new_[4864]_  | ~\new_[18316]_ ;
  assign \new_[4563]_  = ~\new_[4865]_  | ~\new_[19559]_ ;
  assign \new_[4564]_  = ~\new_[4864]_  | ~\new_[19100]_ ;
  assign \new_[4565]_  = ~\new_[4865]_  | ~\new_[19452]_ ;
  assign \new_[4566]_  = ~\new_[4865]_  | ~\new_[18894]_ ;
  assign \new_[4567]_  = ~\new_[4864]_  | ~\new_[19294]_ ;
  assign \new_[4568]_  = ~\new_[4863]_  | ~\new_[17979]_ ;
  assign \new_[4569]_  = ~\new_[4865]_  | ~\new_[18552]_ ;
  assign \new_[4570]_  = ~\new_[4863]_  | ~\new_[18193]_ ;
  assign \new_[4571]_  = ~\new_[4865]_  | ~\new_[19115]_ ;
  assign \new_[4572]_  = ~\new_[4865]_  | ~\new_[19528]_ ;
  assign \new_[4573]_  = ~\new_[4864]_  | ~\new_[18731]_ ;
  assign \new_[4574]_  = ~\new_[4863]_  | ~\new_[19715]_ ;
  assign \new_[4575]_  = ~\new_[4865]_  | ~\new_[18827]_ ;
  assign \new_[4576]_  = ~\new_[4863]_  | ~\new_[19470]_ ;
  assign \new_[4577]_  = ~\new_[4865]_  | ~\new_[17991]_ ;
  assign \new_[4578]_  = ~\new_[4863]_  | ~\new_[18393]_ ;
  assign \new_[4579]_  = ~\new_[4865]_  | ~\new_[17875]_ ;
  assign \new_[4580]_  = ~\new_[4863]_  | ~\new_[18833]_ ;
  assign \new_[4581]_  = ~\new_[4865]_  | ~\new_[19237]_ ;
  assign \new_[4582]_  = ~\new_[12488]_  & (~\new_[4928]_  | ~\new_[5511]_ );
  assign \new_[4583]_  = ~\new_[4863]_  | ~\new_[19261]_ ;
  assign \new_[4584]_  = ~\new_[4984]_  | ~\new_[10947]_  | ~\new_[6555]_  | ~\new_[10967]_ ;
  assign \new_[4585]_  = ~\new_[18711]_  | ~\new_[4865]_ ;
  assign \new_[4586]_  = ~\new_[4864]_  | ~\new_[19740]_ ;
  assign \new_[4587]_  = ~\new_[4865]_  | ~\new_[19723]_ ;
  assign \new_[4588]_  = ~\new_[4864]_  | ~\new_[19078]_ ;
  assign \new_[4589]_  = ~\new_[4865]_  | ~\new_[19736]_ ;
  assign \new_[4590]_  = ~\new_[4864]_  | ~\new_[19411]_ ;
  assign \new_[4591]_  = ~\new_[4865]_  | ~\new_[18854]_ ;
  assign \new_[4592]_  = ~\new_[4864]_  | ~\new_[19185]_ ;
  assign \new_[4593]_  = ~\new_[4865]_  | ~\new_[19531]_ ;
  assign n1695 = ~\new_[10979]_  | ~\new_[4867]_ ;
  assign n1715 = ~\new_[10982]_  | ~\new_[4869]_ ;
  assign \new_[4596]_  = ~\new_[4864]_  | ~\new_[18074]_ ;
  assign \new_[4597]_  = ~\new_[4865]_  | ~\new_[18980]_ ;
  assign \new_[4598]_  = ~\new_[4864]_  | ~\new_[18490]_ ;
  assign \new_[4599]_  = ~\new_[4865]_  | ~\new_[18309]_ ;
  assign n1700 = ~\new_[10992]_  | ~\new_[4868]_ ;
  assign \new_[4601]_  = ~\new_[15992]_  | ~\new_[15424]_  | ~\new_[4875]_  | ~\new_[17123]_ ;
  assign n1705 = ~\new_[11164]_  | ~\new_[4867]_ ;
  assign n1720 = ~\new_[11165]_  | ~\new_[4869]_ ;
  assign n1710 = ~\new_[11168]_  | ~\new_[4868]_ ;
  assign n1725 = ~\new_[10927]_  | ~\new_[4866]_ ;
  assign \new_[4606]_  = ~\new_[4762]_ ;
  assign n1730 = ~\new_[10987]_  | ~\new_[4876]_ ;
  assign n1735 = ~\new_[11156]_  | ~\new_[4876]_ ;
  assign \new_[4609]_  = ~\new_[20082]_  & (~\new_[15692]_  | ~\new_[4900]_ );
  assign \new_[4610]_  = ~\new_[20325]_  & (~\new_[4905]_  | ~\new_[12468]_ );
  assign \new_[4611]_  = ~\new_[4855]_  & ~\new_[19909]_ ;
  assign \new_[4612]_  = ~\new_[20397]_  | ~\new_[5002]_  | ~\new_[13681]_  | ~\new_[11974]_ ;
  assign \wbs_dat_o[10]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[10] ;
  assign \wbs_dat_o[11]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[11] ;
  assign \wbs_dat_o[16]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[16] ;
  assign \wbs_dat_o[18]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[18] ;
  assign \wbs_dat_o[19]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[19] ;
  assign \wbs_dat_o[1]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[1] ;
  assign \wbs_dat_o[21]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[21] ;
  assign \wbs_dat_o[22]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[22] ;
  assign \wbs_dat_o[30]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[30] ;
  assign \wbs_dat_o[5]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[5] ;
  assign \wbs_dat_o[6]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[6] ;
  assign pci_perr_o = pci_io_mux_perr_iob_dat_out_reg;
  assign pci_serr_oe_o = pci_io_mux_serr_iob_en_out_reg;
  assign pci_serr_o = pci_io_mux_serr_iob_dat_out_reg;
  assign \new_[4627]_  = pci_target_unit_wishbone_master_first_wb_data_access_reg;
  assign \new_[4628]_  = ~\new_[5074]_  | ~\new_[15908]_  | ~\new_[17123]_  | ~\new_[15992]_ ;
  assign \new_[4629]_  = ~\new_[4912]_  | ~\new_[19064]_ ;
  assign \new_[4630]_  = ~\new_[4912]_  | ~\new_[18377]_ ;
  assign \new_[4631]_  = ~\new_[4912]_  | ~\new_[18660]_ ;
  assign \new_[4632]_  = ~\new_[4912]_  | ~\new_[18051]_ ;
  assign \new_[4633]_  = ~\new_[4911]_  | ~\new_[18375]_ ;
  assign \new_[4634]_  = ~\new_[4914]_  | ~\new_[19401]_ ;
  assign \new_[4635]_  = ~\new_[4912]_  | ~\new_[19005]_ ;
  assign \new_[4636]_  = ~\new_[4912]_  | ~\new_[18376]_ ;
  assign \new_[4637]_  = ~\new_[4912]_  | ~\new_[19031]_ ;
  assign \new_[4638]_  = ~\new_[4912]_  | ~\new_[18053]_ ;
  assign \new_[4639]_  = ~\new_[4912]_  | ~\new_[19660]_ ;
  assign \new_[4640]_  = ~\new_[4914]_  | ~\new_[18866]_ ;
  assign \new_[4641]_  = ~\new_[4912]_  | ~\new_[18500]_ ;
  assign \new_[4642]_  = ~\new_[4912]_  | ~\new_[19805]_ ;
  assign \new_[4643]_  = ~\new_[4912]_  | ~\new_[19081]_ ;
  assign \new_[4644]_  = ~\new_[4914]_  | ~\new_[18870]_ ;
  assign \new_[4645]_  = ~\new_[4914]_  | ~\new_[18849]_ ;
  assign \new_[4646]_  = ~\new_[4911]_  | ~\new_[17811]_ ;
  assign \new_[4647]_  = ~\new_[4912]_  | ~\new_[19603]_ ;
  assign \new_[4648]_  = ~\new_[4912]_  | ~\new_[19554]_ ;
  assign \new_[4649]_  = ~\new_[4912]_  | ~\new_[19357]_ ;
  assign \new_[4650]_  = ~\new_[4912]_  | ~\new_[18761]_ ;
  assign \new_[4651]_  = ~\new_[4911]_  | ~\new_[18821]_ ;
  assign \new_[4652]_  = ~\new_[4911]_  | ~\new_[19355]_ ;
  assign \new_[4653]_  = ~\new_[4912]_  | ~\new_[18757]_ ;
  assign \new_[4654]_  = ~\new_[4912]_  | ~\new_[19299]_ ;
  assign \new_[4655]_  = ~\new_[4914]_  | ~\new_[18984]_ ;
  assign \new_[4656]_  = ~\new_[4912]_  | ~\new_[19508]_ ;
  assign \new_[4657]_  = ~\new_[4912]_  | ~\new_[19298]_ ;
  assign \new_[4658]_  = ~\new_[4912]_  | ~\new_[19618]_ ;
  assign \new_[4659]_  = ~\new_[4912]_  | ~\new_[18429]_ ;
  assign \new_[4660]_  = ~\new_[4911]_  | ~\new_[19290]_ ;
  assign \new_[4661]_  = ~\new_[4914]_  | ~\new_[18572]_ ;
  assign \new_[4662]_  = ~\new_[4911]_  | ~\new_[19286]_ ;
  assign \new_[4663]_  = ~\new_[4911]_  | ~\new_[18307]_ ;
  assign \new_[4664]_  = ~\new_[4912]_  | ~\new_[18249]_ ;
  assign \new_[4665]_  = ~\new_[4912]_  | ~\new_[19028]_ ;
  assign \new_[4666]_  = ~\new_[4911]_  | ~\new_[19209]_ ;
  assign \new_[4667]_  = ~\new_[4911]_  | ~\new_[18228]_ ;
  assign \new_[4668]_  = ~\new_[4912]_  | ~\new_[19359]_ ;
  assign \new_[4669]_  = ~\new_[4911]_  | ~\new_[19281]_ ;
  assign \new_[4670]_  = ~\new_[4912]_  | ~\new_[18398]_ ;
  assign \new_[4671]_  = ~\new_[4914]_  | ~\new_[18344]_ ;
  assign \new_[4672]_  = ~\new_[4912]_  | ~\new_[19717]_ ;
  assign \new_[4673]_  = ~\new_[4912]_  | ~\new_[18237]_ ;
  assign \new_[4674]_  = ~\new_[4912]_  | ~\new_[19134]_ ;
  assign \new_[4675]_  = ~\new_[4912]_  | ~\new_[19280]_ ;
  assign \new_[4676]_  = ~\new_[4926]_  | ~\new_[17947]_ ;
  assign \new_[4677]_  = ~\new_[4908]_  | ~\new_[17818]_ ;
  assign \new_[4678]_  = ~\new_[4922]_  | ~\new_[18017]_ ;
  assign \new_[4679]_  = ~\new_[4922]_  | ~\new_[19761]_ ;
  assign \new_[4680]_  = ~\new_[4908]_  | ~\new_[17993]_ ;
  assign \new_[4681]_  = ~\new_[4908]_  | ~\new_[17954]_ ;
  assign \new_[4682]_  = ~\new_[4919]_  | ~\new_[18408]_ ;
  assign \new_[4683]_  = ~\new_[4920]_  | ~\new_[17872]_ ;
  assign \new_[4684]_  = ~\new_[4908]_  | ~\new_[19661]_ ;
  assign \new_[4685]_  = ~\new_[4922]_  | ~\new_[19667]_ ;
  assign \new_[4686]_  = ~\new_[4922]_  | ~\new_[18094]_ ;
  assign \new_[4687]_  = ~\new_[4909]_  | ~\new_[19622]_ ;
  assign \new_[4688]_  = ~\new_[4908]_  | ~\new_[19804]_ ;
  assign \new_[4689]_  = ~\new_[4907]_  | ~\new_[19244]_ ;
  assign \new_[4690]_  = ~\new_[4922]_  | ~\new_[19426]_ ;
  assign \new_[4691]_  = ~\new_[4919]_  | ~\new_[18669]_ ;
  assign \new_[4692]_  = ~\new_[4920]_  | ~\new_[19568]_ ;
  assign \new_[4693]_  = ~\new_[4909]_  | ~\new_[18006]_ ;
  assign \new_[4694]_  = ~\new_[4922]_  | ~\new_[19570]_ ;
  assign \new_[4695]_  = ~\new_[4908]_  | ~\new_[19642]_ ;
  assign \new_[4696]_  = ~\new_[4922]_  | ~\new_[18592]_ ;
  assign \new_[4697]_  = ~\new_[4907]_  | ~\new_[18570]_ ;
  assign \new_[4698]_  = ~\new_[4922]_  | ~\new_[19465]_ ;
  assign \new_[4699]_  = ~\new_[4919]_  | ~\new_[18413]_ ;
  assign \new_[4700]_  = ~\new_[4920]_  | ~\new_[19046]_ ;
  assign \new_[4701]_  = ~\new_[4907]_  | ~\new_[18662]_ ;
  assign \new_[4702]_  = ~\new_[4922]_  | ~\new_[19492]_ ;
  assign \new_[4703]_  = ~\new_[4908]_  | ~\new_[19766]_ ;
  assign \new_[4704]_  = ~\new_[4919]_  | ~\new_[18182]_ ;
  assign \new_[4705]_  = ~\new_[4920]_  | ~\new_[18243]_ ;
  assign \new_[4706]_  = ~\new_[4908]_  | ~\new_[19442]_ ;
  assign \new_[4707]_  = ~\new_[4922]_  | ~\new_[17935]_ ;
  assign \new_[4708]_  = ~\new_[4908]_  | ~\new_[18819]_ ;
  assign \new_[4709]_  = ~\new_[4922]_  | ~\new_[19688]_ ;
  assign \new_[4710]_  = ~\new_[4909]_  | ~\new_[18005]_ ;
  assign \new_[4711]_  = ~\new_[4908]_  | ~\new_[18508]_ ;
  assign \new_[4712]_  = ~\new_[4907]_  | ~\new_[18647]_ ;
  assign \new_[4713]_  = ~\new_[4922]_  | ~\new_[18348]_ ;
  assign \new_[4714]_  = ~\new_[4908]_  | ~\new_[18524]_ ;
  assign \new_[4715]_  = ~\new_[4922]_  | ~\new_[19606]_ ;
  assign \new_[4716]_  = ~\new_[4908]_  | ~\new_[18410]_ ;
  assign \new_[4717]_  = ~\new_[4922]_  | ~\new_[19641]_ ;
  assign \new_[4718]_  = ~\new_[4908]_  | ~\new_[18233]_ ;
  assign \new_[4719]_  = ~\new_[4908]_  | ~\new_[17862]_ ;
  assign \new_[4720]_  = ~\new_[4922]_  | ~\new_[18415]_ ;
  assign \new_[4721]_  = ~\new_[4908]_  | ~\new_[19447]_ ;
  assign \new_[4722]_  = ~\new_[4922]_  | ~\new_[19843]_ ;
  assign \new_[4723]_  = ~\new_[4908]_  | ~\new_[19557]_ ;
  assign \new_[4724]_  = ~\new_[4908]_  | ~\new_[19839]_ ;
  assign \new_[4725]_  = ~\new_[4908]_  | ~\new_[19060]_ ;
  assign \new_[4726]_  = ~\new_[4908]_  | ~\new_[19731]_ ;
  assign \new_[4727]_  = ~\new_[4922]_  | ~\new_[19814]_ ;
  assign \new_[4728]_  = ~\new_[4908]_  | ~\new_[18387]_ ;
  assign \new_[4729]_  = ~\new_[4922]_  | ~\new_[19105]_ ;
  assign \new_[4730]_  = ~\new_[4909]_  | ~\new_[18841]_ ;
  assign \new_[4731]_  = ~\new_[4908]_  | ~\new_[19034]_ ;
  assign \new_[4732]_  = ~\new_[4919]_  | ~\new_[18313]_ ;
  assign \new_[4733]_  = ~\new_[4922]_  | ~\new_[18411]_ ;
  assign \new_[4734]_  = ~\new_[4920]_  | ~\new_[18809]_ ;
  assign \new_[4735]_  = ~\new_[4908]_  | ~\new_[19193]_ ;
  assign \new_[4736]_  = ~\new_[4919]_  | ~\new_[19306]_ ;
  assign \new_[4737]_  = ~\new_[4920]_  | ~\new_[18661]_ ;
  assign \new_[4738]_  = ~\new_[4909]_  | ~\new_[18732]_ ;
  assign \new_[4739]_  = ~\new_[4922]_  | ~\new_[19187]_ ;
  assign \new_[4740]_  = ~\new_[4919]_  | ~\new_[18838]_ ;
  assign \new_[4741]_  = ~\new_[4920]_  | ~\new_[18904]_ ;
  assign \new_[4742]_  = ~\new_[4908]_  | ~\new_[18806]_ ;
  assign \new_[4743]_  = ~\new_[4919]_  | ~\new_[18802]_ ;
  assign \new_[4744]_  = ~\new_[4920]_  | ~\new_[18799]_ ;
  assign \new_[4745]_  = ~\new_[4909]_  | ~\new_[18215]_ ;
  assign \new_[4746]_  = ~\new_[4922]_  | ~\new_[18188]_ ;
  assign \new_[4747]_  = ~\new_[4908]_  | ~\new_[19112]_ ;
  assign \new_[4748]_  = ~\new_[4922]_  | ~\new_[18634]_ ;
  assign \new_[4749]_  = ~\new_[4907]_  | ~\new_[18957]_ ;
  assign \new_[4750]_  = ~\new_[4922]_  | ~\new_[19597]_ ;
  assign \new_[4751]_  = ~\new_[4908]_  | ~\new_[18278]_ ;
  assign \new_[4752]_  = ~\new_[4908]_  | ~\new_[18717]_ ;
  assign \new_[4753]_  = ~\new_[4907]_  | ~\new_[18442]_ ;
  assign \new_[4754]_  = ~\new_[4922]_  | ~\new_[17820]_ ;
  assign \new_[4755]_  = ~\new_[4919]_  | ~\new_[19445]_ ;
  assign \new_[4756]_  = ~\new_[4920]_  | ~\new_[17865]_ ;
  assign \new_[4757]_  = ~\new_[4908]_  | ~\new_[18610]_ ;
  assign \new_[4758]_  = ~\new_[4908]_  | ~\new_[18858]_ ;
  assign \new_[4759]_  = \new_[20401]_  | \new_[4903]_ ;
  assign \new_[4760]_  = ~\new_[4857]_ ;
  assign \new_[4761]_  = (~\new_[11154]_  | ~\new_[5325]_ ) & (~\new_[15577]_  | ~\new_[20505]_ );
  assign \new_[4762]_  = ~output_backup_perr_out_reg;
  assign \new_[4763]_  = output_backup_serr_out_reg;
  assign \new_[4764]_  = \new_[4935]_  | \new_[11893]_ ;
  assign \new_[4765]_  = \new_[4936]_  | \new_[12487]_ ;
  assign \new_[4766]_  = \new_[4937]_  | \new_[12488]_ ;
  assign \new_[4767]_  = \new_[4938]_  | \new_[12488]_ ;
  assign \new_[4768]_  = \new_[4939]_  | \new_[12487]_ ;
  assign \new_[4769]_  = \new_[4940]_  | \new_[11893]_ ;
  assign \new_[4770]_  = \new_[4941]_  | \new_[12487]_ ;
  assign \new_[4771]_  = \new_[4956]_  | \new_[11893]_ ;
  assign \new_[4772]_  = \new_[4942]_  | \new_[12487]_ ;
  assign \new_[4773]_  = \new_[4943]_  | \new_[12487]_ ;
  assign \new_[4774]_  = \new_[4957]_  | \new_[12487]_ ;
  assign \new_[4775]_  = \new_[4944]_  | \new_[12488]_ ;
  assign n1750 = ~\new_[4946]_  & ~\new_[5513]_ ;
  assign \new_[4777]_  = \new_[4950]_  | \new_[13807]_ ;
  assign \new_[4778]_  = \new_[4952]_  | \new_[12487]_ ;
  assign \new_[4779]_  = \new_[4953]_  | \new_[13807]_ ;
  assign \new_[4780]_  = \new_[4954]_  | \new_[12487]_ ;
  assign \new_[4781]_  = \new_[4951]_  | \new_[12487]_ ;
  assign \new_[4782]_  = \new_[4929]_  | \new_[13807]_ ;
  assign \new_[4783]_  = \new_[4930]_  | \new_[13807]_ ;
  assign \new_[4784]_  = \new_[4931]_  | \new_[12488]_ ;
  assign \new_[4785]_  = \new_[13807]_  | \new_[4932]_ ;
  assign \new_[4786]_  = \new_[4933]_  | \new_[11893]_ ;
  assign \new_[4787]_  = \new_[4934]_  | \new_[12488]_ ;
  assign \new_[4788]_  = \new_[4945]_  | \new_[12488]_ ;
  assign n1740 = ~\new_[11159]_  | ~\new_[4958]_ ;
  assign \new_[4790]_  = ~\new_[20082]_  & (~\new_[4982]_  | ~\new_[20505]_ );
  assign n1745 = ~\new_[11007]_  | ~\new_[4958]_ ;
  assign \new_[4792]_  = \new_[4949]_  | \new_[12487]_ ;
  assign \wbs_dat_o[15]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[15] ;
  assign \wbs_dat_o[24]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[24] ;
  assign \wbs_dat_o[25]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[25] ;
  assign \wbs_dat_o[27]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[27] ;
  assign \wbs_dat_o[2]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[2] ;
  assign \new_[4798]_  = ~\new_[4986]_  | ~\new_[18028]_ ;
  assign \new_[4799]_  = ~\new_[4987]_  | ~\new_[18270]_ ;
  assign \new_[4800]_  = ~\new_[4986]_  | ~\new_[18032]_ ;
  assign \new_[4801]_  = ~\new_[4987]_  | ~\new_[18271]_ ;
  assign \new_[4802]_  = ~\new_[4987]_  | ~\new_[18702]_ ;
  assign \new_[4803]_  = ~\new_[4986]_  | ~\new_[18623]_ ;
  assign \new_[4804]_  = ~\new_[4986]_  | ~\new_[18273]_ ;
  assign \new_[4805]_  = ~\new_[4987]_  | ~\new_[18638]_ ;
  assign \new_[4806]_  = ~\new_[4986]_  | ~\new_[18625]_ ;
  assign \new_[4807]_  = ~\new_[4986]_  | ~\new_[18378]_ ;
  assign \new_[4808]_  = ~\new_[4988]_  | ~\new_[18853]_ ;
  assign \new_[4809]_  = ~\new_[4986]_  | ~\new_[18025]_ ;
  assign \new_[4810]_  = ~\new_[4988]_  | ~\new_[18274]_ ;
  assign \new_[4811]_  = ~\new_[4988]_  | ~\new_[19433]_ ;
  assign \new_[4812]_  = ~\new_[4987]_  | ~\new_[18612]_ ;
  assign \new_[4813]_  = ~\new_[4986]_  | ~\new_[18275]_ ;
  assign \new_[4814]_  = ~\new_[4987]_  | ~\new_[18496]_ ;
  assign \new_[4815]_  = ~\new_[4989]_  | ~\new_[18622]_ ;
  assign \new_[4816]_  = ~\new_[4988]_  | ~\new_[19379]_ ;
  assign \new_[4817]_  = ~\new_[4987]_  | ~\new_[18423]_ ;
  assign \new_[4818]_  = ~\new_[4988]_  | ~\new_[18896]_ ;
  assign \new_[4819]_  = ~\new_[4988]_  | ~\new_[18949]_ ;
  assign \new_[4820]_  = ~\new_[4987]_  | ~\new_[18713]_ ;
  assign \new_[4821]_  = ~\new_[4986]_  | ~\new_[18784]_ ;
  assign \new_[4822]_  = ~\new_[4987]_  | ~\new_[18360]_ ;
  assign \new_[4823]_  = ~\new_[4986]_  | ~\new_[18606]_ ;
  assign \new_[4824]_  = ~\new_[4988]_  | ~\new_[18652]_ ;
  assign \new_[4825]_  = ~\new_[4987]_  | ~\new_[18699]_ ;
  assign \new_[4826]_  = ~\new_[4986]_  | ~\new_[18364]_ ;
  assign \new_[4827]_  = ~\new_[4989]_  | ~\new_[19436]_ ;
  assign \new_[4828]_  = ~\new_[4987]_  | ~\new_[18715]_ ;
  assign \new_[4829]_  = ~\new_[4987]_  | ~\new_[18803]_ ;
  assign \new_[4830]_  = ~\new_[4989]_  | ~\new_[18725]_ ;
  assign \new_[4831]_  = ~\new_[4986]_  | ~\new_[18745]_ ;
  assign \new_[4832]_  = ~\new_[4988]_  | ~\new_[19301]_ ;
  assign \new_[4833]_  = ~\new_[4986]_  | ~\new_[18773]_ ;
  assign \new_[4834]_  = ~\new_[4989]_  | ~\new_[18635]_ ;
  assign \new_[4835]_  = ~\new_[4986]_  | ~\new_[18837]_ ;
  assign \new_[4836]_  = ~\new_[4989]_  | ~\new_[18269]_ ;
  assign \new_[4837]_  = ~\new_[4986]_  | ~\new_[18372]_ ;
  assign \new_[4838]_  = ~\new_[4998]_  | ~\new_[19646]_ ;
  assign \new_[4839]_  = ~\new_[4998]_  | ~\new_[18104]_ ;
  assign \new_[4840]_  = ~\new_[4998]_  | ~\new_[19095]_ ;
  assign \new_[4841]_  = ~\new_[4998]_  | ~\new_[17950]_ ;
  assign \new_[4842]_  = ~\new_[4998]_  | ~\new_[18505]_ ;
  assign \new_[4843]_  = ~\new_[4998]_  | ~\new_[19601]_ ;
  assign \new_[4844]_  = ~\new_[4998]_  | ~\new_[18599]_ ;
  assign \new_[4845]_  = ~\new_[4998]_  | ~\new_[19098]_ ;
  assign \new_[4846]_  = ~\new_[4998]_  | ~\new_[18177]_ ;
  assign \new_[4847]_  = ~\new_[4998]_  | ~\new_[19751]_ ;
  assign \new_[4848]_  = ~\new_[4998]_  | ~\new_[18346]_ ;
  assign \new_[4849]_  = ~\new_[4998]_  | ~\new_[18804]_ ;
  assign \new_[4850]_  = ~\new_[4998]_  | ~\new_[17936]_ ;
  assign \new_[4851]_  = ~\new_[4998]_  | ~\new_[18334]_ ;
  assign \new_[4852]_  = ~\new_[4998]_  | ~\new_[19195]_ ;
  assign \new_[4853]_  = ~\new_[4998]_  | ~\new_[18232]_ ;
  assign \new_[4854]_  = ~\new_[19946]_  | ~\new_[16228]_  | ~\new_[5274]_ ;
  assign \new_[4855]_  = ~\new_[13854]_  & (~\new_[14293]_  | ~\new_[5097]_ );
  assign \new_[4856]_  = ~\new_[4899]_ ;
  assign \new_[4857]_  = (~\new_[5274]_  | ~\new_[16211]_ ) & (~\new_[7283]_  | ~n16385);
  assign \new_[4858]_  = ~\new_[4913]_ ;
  assign \new_[4859]_  = ~\new_[4913]_ ;
  assign \new_[4860]_  = ~\new_[4915]_ ;
  assign \new_[4861]_  = ~\new_[4916]_ ;
  assign \new_[4862]_  = ~\new_[4916]_ ;
  assign \new_[4863]_  = ~\new_[4918]_ ;
  assign \new_[4864]_  = ~\new_[4918]_ ;
  assign \new_[4865]_  = ~\new_[4921]_ ;
  assign \new_[4866]_  = ~output_backup_serr_en_out_reg;
  assign \new_[4867]_  = \new_[5003]_  | \new_[12488]_ ;
  assign \new_[4868]_  = \new_[5005]_  | \new_[12488]_ ;
  assign \new_[4869]_  = \new_[5004]_  | \new_[12487]_ ;
  assign n1755 = ~\new_[10986]_  | ~\new_[5006]_ ;
  assign \new_[4871]_  = ~\new_[4959]_  | ~\new_[16980]_ ;
  assign \new_[4872]_  = ~\new_[4960]_  | ~\new_[16982]_ ;
  assign \new_[4873]_  = ~\new_[4961]_  | ~\new_[16880]_ ;
  assign n1760 = ~\new_[11001]_  | ~\new_[5006]_ ;
  assign \new_[4875]_  = ~\new_[16994]_  & ~\new_[4983]_ ;
  assign \new_[4876]_  = ~\new_[5199]_  & (~\new_[5887]_  | ~\new_[5078]_ );
  assign n1770 = ~\new_[12573]_  | (~\new_[5089]_  & ~\new_[13718]_ );
  assign n1775 = ~\new_[12574]_  | (~\new_[5091]_  & ~\new_[13718]_ );
  assign n1765 = ~\new_[12572]_  | (~\new_[5088]_  & ~\new_[13718]_ );
  assign \wbs_dat_o[0]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[0] ;
  assign \wbs_dat_o[12]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[12] ;
  assign \wbs_dat_o[13]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[13] ;
  assign \wbs_dat_o[14]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[14] ;
  assign \wbs_dat_o[17]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[17] ;
  assign \wbs_dat_o[20]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[20] ;
  assign \wbs_dat_o[23]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[23] ;
  assign \wbs_dat_o[26]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[26] ;
  assign \wbs_dat_o[28]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[28] ;
  assign \wbs_dat_o[29]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[29] ;
  assign \wbs_dat_o[31]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[31] ;
  assign \wbs_dat_o[3]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[3] ;
  assign \wbs_dat_o[4]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[4] ;
  assign \wbs_dat_o[7]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[7] ;
  assign \wbs_dat_o[8]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[8] ;
  assign \wbs_dat_o[9]  = \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[9] ;
  assign \new_[4896]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24] ;
  assign n1780 = \wbs_dat_o[10]  ? \new_[9284]_  : \new_[5163]_ ;
  assign n1785 = \wbs_dat_o[11]  ? \new_[9284]_  : \new_[5164]_ ;
  assign \new_[4899]_  = ~\new_[17123]_  | ~\new_[16211]_  | ~\new_[5274]_  | ~\new_[16889]_ ;
  assign \new_[4900]_  = (~\new_[16436]_  | ~n16385) & (~\new_[5325]_  | ~\new_[16211]_ );
  assign n1790 = \wbs_dat_o[16]  ? \new_[9284]_  : \new_[5165]_ ;
  assign n1795 = \wbs_dat_o[18]  ? \new_[9284]_  : \new_[5166]_ ;
  assign \new_[4903]_  = \new_[11974]_  & \new_[5097]_ ;
  assign n1800 = \wbs_dat_o[19]  ? \new_[9284]_  : \new_[5167]_ ;
  assign \new_[4905]_  = ~\new_[17467]_  | ~\new_[5274]_  | ~\new_[17797]_ ;
  assign n1805 = \wbs_dat_o[1]  ? \new_[9284]_  : \new_[5168]_ ;
  assign \new_[4907]_  = ~\new_[5118]_ ;
  assign \new_[4908]_  = ~\new_[5118]_ ;
  assign \new_[4909]_  = ~\new_[5118]_ ;
  assign n1810 = \wbs_dat_o[21]  ? \new_[9284]_  : \new_[5169]_ ;
  assign \new_[4911]_  = ~\new_[4990]_ ;
  assign \new_[4912]_  = ~\new_[4991]_ ;
  assign \new_[4913]_  = ~\new_[4992]_ ;
  assign \new_[4914]_  = \new_[4993]_ ;
  assign \new_[4915]_  = ~\new_[4993]_ ;
  assign \new_[4916]_  = ~\new_[4993]_ ;
  assign n1815 = \wbs_dat_o[22]  ? \new_[9284]_  : \new_[5170]_ ;
  assign \new_[4918]_  = ~\new_[4995]_ ;
  assign \new_[4919]_  = \new_[4995]_ ;
  assign \new_[4920]_  = \new_[4997]_ ;
  assign \new_[4921]_  = ~\new_[4997]_ ;
  assign \new_[4922]_  = ~\new_[4999]_ ;
  assign n1820 = \wbs_dat_o[30]  ? \new_[9284]_  : \new_[5171]_ ;
  assign n1825 = \wbs_dat_o[5]  ? \new_[9284]_  : \new_[5172]_ ;
  assign n1830 = \wbs_dat_o[6]  ? \new_[9284]_  : \new_[5173]_ ;
  assign \new_[4926]_  = (~\new_[14278]_  | ~\new_[5161]_ ) & (~wbm_ack_i | ~wbm_stb_o);
  assign n1850 = ~\new_[16172]_  | ~wbm_cyc_o;
  assign \new_[4928]_  = ~\new_[5066]_  & (~\new_[11884]_  | ~\new_[6162]_ );
  assign \new_[4929]_  = ~\new_[5191]_  & (~\new_[5121]_  | ~\new_[6330]_ );
  assign \new_[4930]_  = ~\new_[5192]_  & (~\new_[5122]_  | ~\new_[6330]_ );
  assign \new_[4931]_  = ~\new_[5193]_  & (~\new_[5123]_  | ~\new_[5989]_ );
  assign \new_[4932]_  = ~\new_[5194]_  & (~\new_[5124]_  | ~\new_[5989]_ );
  assign \new_[4933]_  = ~\new_[5195]_  & (~\new_[5125]_  | ~\new_[6330]_ );
  assign \new_[4934]_  = ~\new_[5197]_  & (~\new_[5126]_  | ~\new_[6330]_ );
  assign \new_[4935]_  = ~\new_[5216]_  & (~\new_[5127]_  | ~\new_[5988]_ );
  assign \new_[4936]_  = ~\new_[5198]_  & (~\new_[5128]_  | ~\new_[6330]_ );
  assign \new_[4937]_  = ~\new_[5200]_  & (~\new_[5129]_  | ~\new_[6330]_ );
  assign \new_[4938]_  = ~\new_[5201]_  & (~\new_[5130]_  | ~\new_[5989]_ );
  assign \new_[4939]_  = ~\new_[5202]_  & (~\new_[5131]_  | ~\new_[6330]_ );
  assign \new_[4940]_  = ~\new_[5203]_  & (~\new_[5132]_  | ~\new_[6330]_ );
  assign \new_[4941]_  = ~\new_[5205]_  & (~\new_[5133]_  | ~\new_[6330]_ );
  assign \new_[4942]_  = ~\new_[5206]_  & (~\new_[5134]_  | ~\new_[6330]_ );
  assign \new_[4943]_  = ~\new_[5207]_  & (~\new_[5135]_  | ~\new_[6330]_ );
  assign \new_[4944]_  = ~\new_[5208]_  & (~\new_[5136]_  | ~\new_[6330]_ );
  assign \new_[4945]_  = ~\new_[5209]_  & (~\new_[5137]_  | ~\new_[6936]_ );
  assign \new_[4946]_  = ~\new_[5072]_  | ~\new_[17519]_ ;
  assign n1855 = ~\new_[5444]_  | ~\new_[5072]_ ;
  assign n1860 = ~\new_[5072]_  | ~\new_[13120]_ ;
  assign \new_[4949]_  = ~\new_[5211]_  & (~\new_[5139]_  | ~\new_[6330]_ );
  assign \new_[4950]_  = ~\new_[5212]_  & (~\new_[5140]_  | ~\new_[5988]_ );
  assign \new_[4951]_  = ~\new_[5213]_  & (~\new_[5141]_  | ~\new_[5988]_ );
  assign \new_[4952]_  = ~\new_[5214]_  & (~\new_[5142]_  | ~\new_[6330]_ );
  assign \new_[4953]_  = ~\new_[5215]_  & (~\new_[5143]_  | ~\new_[5989]_ );
  assign \new_[4954]_  = ~\new_[5116]_  & (~\new_[5120]_  | ~\new_[6330]_ );
  assign n1840 = ~n1890;
  assign \new_[4956]_  = ~\new_[5068]_  & (~\new_[5442]_  | ~\new_[6165]_ );
  assign \new_[4957]_  = ~\new_[5069]_  & (~\new_[5350]_  | ~\new_[6165]_ );
  assign \new_[4958]_  = ~\new_[5210]_  & (~\new_[5887]_  | ~\new_[5138]_ );
  assign \new_[4959]_  = (~\new_[5225]_  | ~\new_[17279]_ ) & (~\new_[17038]_  | ~\new_[5047]_ );
  assign \new_[4960]_  = (~\new_[5226]_  | ~\new_[17279]_ ) & (~\new_[17038]_  | ~\new_[5045]_ );
  assign \new_[4961]_  = (~\new_[5227]_  | ~\new_[17279]_ ) & (~\new_[17038]_  | ~\new_[5046]_ );
  assign \new_[4962]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3] ;
  assign \new_[4963]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12] ;
  assign \new_[4964]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14] ;
  assign \new_[4965]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17] ;
  assign \new_[4966]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18] ;
  assign \new_[4967]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20] ;
  assign \new_[4968]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21] ;
  assign \new_[4969]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22] ;
  assign \new_[4970]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25] ;
  assign \new_[4971]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26] ;
  assign \new_[4972]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27] ;
  assign \new_[4973]_  = ~\\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29] ;
  assign \new_[4974]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2] ;
  assign \new_[4975]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4] ;
  assign \new_[4976]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5] ;
  assign \new_[4977]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7] ;
  assign \new_[4978]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[26] ;
  assign \new_[4979]_  = ~\\pci_target_unit_fifos_pciw_outTransactionCount_reg[1] ;
  assign \new_[4980]_  = ~\\pci_target_unit_fifos_outGreyCount_reg[0] ;
  assign \new_[4981]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0] ;
  assign \new_[4982]_  = ~\new_[5115]_  & ~\new_[16436]_ ;
  assign \new_[4983]_  = ~\new_[5113]_  | ~\new_[15682]_ ;
  assign \new_[4984]_  = ~\new_[16228]_  | ~\new_[19946]_  | ~\new_[5325]_  | ~\new_[20505]_ ;
  assign n1865 = \wbs_dat_o[15]  ? \new_[9284]_  : \new_[5280]_ ;
  assign \new_[4986]_  = ~\new_[5117]_ ;
  assign \new_[4987]_  = ~\new_[5117]_ ;
  assign \new_[4988]_  = ~\new_[5117]_ ;
  assign \new_[4989]_  = ~\new_[5117]_ ;
  assign \new_[4990]_  = ~\new_[5075]_ ;
  assign \new_[4991]_  = ~\new_[5075]_ ;
  assign \new_[4992]_  = ~\new_[19888]_ ;
  assign \new_[4993]_  = ~\new_[20538]_ ;
  assign n1870 = \wbs_dat_o[24]  ? \new_[9284]_  : \new_[5281]_ ;
  assign \new_[4995]_  = ~\new_[5079]_ ;
  assign n1875 = \wbs_dat_o[25]  ? \new_[9284]_  : \new_[5282]_ ;
  assign \new_[4997]_  = ~\new_[5080]_ ;
  assign \new_[4998]_  = \new_[5081]_ ;
  assign \new_[4999]_  = ~\new_[5081]_ ;
  assign n1880 = \wbs_dat_o[27]  ? \new_[9284]_  : \new_[5283]_ ;
  assign n1885 = \wbs_dat_o[2]  ? \new_[9284]_  : \new_[5284]_ ;
  assign \new_[5002]_  = ~\new_[5097]_ ;
  assign \new_[5003]_  = \new_[5279]_  ? \new_[6936]_  : \new_[5217]_ ;
  assign \new_[5004]_  = ~\new_[5196]_  & (~\new_[5218]_  | ~\new_[6330]_ );
  assign \new_[5005]_  = ~\new_[5204]_  & (~\new_[5220]_  | ~\new_[5988]_ );
  assign \new_[5006]_  = ~\new_[5114]_  & (~\new_[5887]_  | ~\new_[5219]_ );
  assign n1890 = ~\new_[5112]_  & ~\new_[11596]_ ;
  assign \new_[5008]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0] ;
  assign \new_[5009]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19] ;
  assign \new_[5010]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23] ;
  assign \new_[5011]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28] ;
  assign \new_[5012]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16] ;
  assign \new_[5013]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[0] ;
  assign \new_[5014]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[2] ;
  assign \new_[5015]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[0] ;
  assign \new_[5016]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[10] ;
  assign \new_[5017]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[11] ;
  assign \new_[5018]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[12] ;
  assign \new_[5019]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[13] ;
  assign \new_[5020]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[14] ;
  assign \new_[5021]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[15] ;
  assign \new_[5022]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[17] ;
  assign \new_[5023]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[18] ;
  assign \new_[5024]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[19] ;
  assign \new_[5025]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[20] ;
  assign \new_[5026]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[22] ;
  assign \new_[5027]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[24] ;
  assign \new_[5028]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[27] ;
  assign \new_[5029]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[28] ;
  assign \new_[5030]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[29] ;
  assign \new_[5031]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[2] ;
  assign \new_[5032]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[31] ;
  assign \new_[5033]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[3] ;
  assign \new_[5034]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[4] ;
  assign \new_[5035]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[6] ;
  assign \new_[5036]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[7] ;
  assign \new_[5037]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[8] ;
  assign \new_[5038]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11] ;
  assign \new_[5039]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13] ;
  assign \new_[5040]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15] ;
  assign \new_[5041]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1] ;
  assign \new_[5042]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6] ;
  assign \new_[5043]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8] ;
  assign \new_[5044]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10] ;
  assign \new_[5045]_  = \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[2] ;
  assign \new_[5046]_  = \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[3] ;
  assign \new_[5047]_  = \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[0] ;
  assign \new_[5048]_  = \\wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[0] ;
  assign \new_[5049]_  = ~\\pci_target_unit_fifos_pciw_outTransactionCount_reg[0] ;
  assign \new_[5050]_  = ~\\pci_target_unit_fifos_outGreyCount_reg[1] ;
  assign \new_[5051]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1] ;
  assign \new_[5052]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2] ;
  assign \new_[5053]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[0] ;
  assign \new_[5054]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[1] ;
  assign \new_[5055]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[2] ;
  assign \new_[5056]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg[0] ;
  assign \new_[5057]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg[2] ;
  assign \new_[5058]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg[0] ;
  assign \new_[5059]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg[1] ;
  assign \new_[5060]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg[2] ;
  assign \new_[5061]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[0] ;
  assign \new_[5062]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[1] ;
  assign \new_[5063]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[2] ;
  assign \new_[5064]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg[1] ;
  assign n1895 = \wbs_dat_o[0]  ? \new_[9284]_  : \new_[5351]_ ;
  assign \new_[5066]_  = ~\new_[6165]_  & (~\new_[5316]_  | ~\new_[16390]_ );
  assign n1900 = \wbs_dat_o[12]  ? \new_[9284]_  : \new_[5352]_ ;
  assign \new_[5068]_  = ~\new_[6165]_  & (~\new_[5318]_  | ~\new_[16393]_ );
  assign \new_[5069]_  = ~\new_[6165]_  & (~\new_[5321]_  | ~\new_[16391]_ );
  assign n1905 = \wbs_dat_o[13]  ? \new_[9284]_  : \new_[5353]_ ;
  assign n1910 = \wbs_dat_o[14]  ? \new_[9284]_  : \new_[5354]_ ;
  assign \new_[5072]_  = ~\new_[5112]_ ;
  assign n1915 = \wbs_dat_o[17]  ? \new_[9284]_  : \new_[5355]_ ;
  assign \new_[5074]_  = ~\new_[5115]_ ;
  assign \new_[5075]_  = ~\new_[5119]_ ;
  assign n1920 = \wbs_dat_o[20]  ? \new_[9284]_  : \new_[5356]_ ;
  assign n1925 = \wbs_dat_o[23]  ? \new_[9284]_  : \new_[5357]_ ;
  assign \new_[5078]_  = ~\new_[5273]_  | ~\new_[16091]_ ;
  assign \new_[5079]_  = ~\new_[20231]_  | ~\new_[5295]_  | ~\new_[20541]_ ;
  assign \new_[5080]_  = ~\new_[20231]_  | ~\new_[5295]_  | ~\new_[19889]_ ;
  assign \new_[5081]_  = ~\new_[20228]_ ;
  assign n1930 = \wbs_dat_o[26]  ? \new_[9284]_  : \new_[5358]_ ;
  assign n1935 = \wbs_dat_o[28]  ? \new_[9284]_  : \new_[5359]_ ;
  assign n1940 = \wbs_dat_o[29]  ? \new_[9284]_  : \new_[5360]_ ;
  assign n1975 = ~\new_[5278]_  | (~\new_[13128]_  & ~\new_[16782]_ );
  assign n1945 = \wbs_dat_o[31]  ? \new_[9284]_  : \new_[5361]_ ;
  assign n1950 = \wbs_dat_o[3]  ? \new_[9284]_  : \new_[5362]_ ;
  assign \new_[5088]_  = ~\new_[5275]_  & (~\new_[18491]_  | ~\new_[20153]_ );
  assign \new_[5089]_  = ~\new_[5276]_  & (~\new_[18224]_  | ~\new_[20153]_ );
  assign \new_[5090]_  = \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9] ;
  assign \new_[5091]_  = ~\new_[5277]_  & (~\new_[19636]_  | ~\new_[20153]_ );
  assign n1955 = \wbs_dat_o[4]  ? \new_[9284]_  : \new_[5363]_ ;
  assign n1960 = \wbs_dat_o[7]  ? \new_[9284]_  : \new_[5364]_ ;
  assign n1965 = \wbs_dat_o[8]  ? \new_[9284]_  : \new_[5365]_ ;
  assign n1970 = \wbs_dat_o[9]  ? \new_[9284]_  : \new_[5366]_ ;
  assign \new_[5096]_  = \\wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[1] ;
  assign \new_[5097]_  = ~\new_[5297]_  & ~\new_[5285]_ ;
  assign wbm_cyc_o = ~\new_[5161]_ ;
  assign \new_[5099]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[5] ;
  assign \new_[5100]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[9] ;
  assign \new_[5101]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[1] ;
  assign \new_[5102]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[23] ;
  assign \new_[5103]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[16] ;
  assign \new_[5104]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[3] ;
  assign \new_[5105]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[21] ;
  assign \new_[5106]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[25] ;
  assign \new_[5107]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0] ;
  assign wbm_we_o = pci_target_unit_wishbone_master_wb_we_o_reg;
  assign \new_[5109]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1] ;
  assign \new_[5110]_  = ~\\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2] ;
  assign n2075 = ~\new_[5298]_  | (~\new_[20229]_  & ~\new_[5495]_ );
  assign \new_[5112]_  = \new_[5441]_  ^ \new_[12364]_ ;
  assign \new_[5113]_  = \new_[5325]_  | \new_[16436]_ ;
  assign \new_[5114]_  = ~\new_[5349]_  & ~\new_[13807]_ ;
  assign \new_[5115]_  = ~\new_[5325]_  | ~\new_[20026]_ ;
  assign \new_[5116]_  = ~\new_[5348]_  & ~\new_[6936]_ ;
  assign \new_[5117]_  = ~\new_[20539]_  | ~\new_[20543]_  | ~\new_[19889]_ ;
  assign \new_[5118]_  = ~\new_[20539]_  | ~\new_[20231]_  | ~\new_[19889]_ ;
  assign \new_[5119]_  = ~\new_[20539]_  | ~\new_[20543]_  | ~\new_[20541]_ ;
  assign \new_[5120]_  = ~\new_[5303]_  | ~\new_[16386]_ ;
  assign \new_[5121]_  = ~\new_[5304]_  | ~\new_[16086]_ ;
  assign \new_[5122]_  = ~\new_[5305]_  | ~\new_[16392]_ ;
  assign \new_[5123]_  = ~\new_[5306]_  | ~\new_[16084]_ ;
  assign \new_[5124]_  = ~\new_[5307]_  | ~\new_[16388]_ ;
  assign \new_[5125]_  = ~\new_[5308]_  | ~\new_[16087]_ ;
  assign \new_[5126]_  = ~\new_[5309]_  | ~\new_[16085]_ ;
  assign \new_[5127]_  = ~\new_[5310]_  | ~\new_[16396]_ ;
  assign \new_[5128]_  = ~\new_[5311]_  | ~\new_[16395]_ ;
  assign \new_[5129]_  = ~\new_[5312]_  | ~\new_[16092]_ ;
  assign \new_[5130]_  = ~\new_[5313]_  | ~\new_[16387]_ ;
  assign \new_[5131]_  = ~\new_[5314]_  | ~\new_[16095]_ ;
  assign \new_[5132]_  = ~\new_[5315]_  | ~\new_[16082]_ ;
  assign \new_[5133]_  = ~\new_[5317]_  | ~\new_[16089]_ ;
  assign \new_[5134]_  = ~\new_[5319]_  | ~\new_[16081]_ ;
  assign \new_[5135]_  = ~\new_[5320]_  | ~\new_[16094]_ ;
  assign \new_[5136]_  = ~\new_[5322]_  | ~\new_[16080]_ ;
  assign \new_[5137]_  = ~\new_[5323]_  | ~\new_[16394]_ ;
  assign \new_[5138]_  = ~\new_[5326]_  | ~\new_[13808]_ ;
  assign \new_[5139]_  = ~\new_[5327]_  | ~\new_[16083]_ ;
  assign \new_[5140]_  = ~\new_[5328]_  | ~\new_[16096]_ ;
  assign \new_[5141]_  = ~\new_[5329]_  | ~\new_[16088]_ ;
  assign \new_[5142]_  = ~\new_[5330]_  | ~\new_[16097]_ ;
  assign \new_[5143]_  = ~\new_[5331]_  | ~\new_[16397]_ ;
  assign n1985 = ~\new_[5332]_  | (~\new_[13785]_  & ~\new_[16782]_ );
  assign n1990 = ~\new_[5333]_  | (~\new_[14203]_  & ~\new_[16782]_ );
  assign n1995 = ~\new_[5334]_  | (~\new_[14232]_  & ~\new_[16782]_ );
  assign n2000 = ~\new_[5335]_  | (~\new_[14864]_  & ~\new_[16782]_ );
  assign n2005 = ~\new_[5336]_  | (~\new_[13783]_  & ~\new_[16782]_ );
  assign n2010 = ~\new_[5337]_  | (~\new_[13830]_  & ~\new_[16782]_ );
  assign n2015 = ~\new_[5338]_  | (~\new_[14202]_  & ~\new_[16782]_ );
  assign n2020 = ~\new_[5339]_  | (~\new_[13640]_  & ~\new_[16782]_ );
  assign n2025 = ~\new_[5340]_  | (~\new_[13796]_  & ~\new_[16782]_ );
  assign n2030 = ~\new_[5341]_  | (~\new_[11813]_  & ~\new_[16782]_ );
  assign n2035 = ~\new_[5342]_  | (~\new_[13147]_  & ~\new_[16782]_ );
  assign n2040 = ~\new_[5343]_  | (~\new_[14235]_  & ~\new_[16782]_ );
  assign n1980 = ~\new_[5344]_  | (~\new_[14860]_  & ~\new_[16782]_ );
  assign n2045 = ~\new_[5345]_  | (~\new_[14854]_  & ~\new_[16782]_ );
  assign n2050 = ~\new_[5346]_  | (~\new_[14236]_  & ~\new_[16782]_ );
  assign n2055 = ~\new_[5347]_  | (~\new_[14858]_  & ~\new_[16782]_ );
  assign n2060 = \new_[18362]_  ? \new_[12189]_  : \new_[5450]_ ;
  assign \new_[5161]_  = ~pci_target_unit_wishbone_master_wb_cyc_o_reg;
  assign wbm_stb_o = pci_target_unit_wishbone_master_wb_stb_o_reg;
  assign \new_[5163]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[10] ;
  assign \new_[5164]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[11] ;
  assign \new_[5165]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[16] ;
  assign \new_[5166]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[18] ;
  assign \new_[5167]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[19] ;
  assign \new_[5168]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[1] ;
  assign \new_[5169]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[21] ;
  assign \new_[5170]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[22] ;
  assign \new_[5171]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[30] ;
  assign \new_[5172]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[5] ;
  assign \new_[5173]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[6] ;
  assign \new_[5174]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[30] ;
  assign n2065 = ~\new_[5292]_  | (~\new_[5493]_  & ~\new_[4979]_ );
  assign n2070 = ~\new_[5292]_  | (~\new_[5493]_  & ~\new_[4980]_ );
  assign n2295 = \new_[16847]_  ? \new_[5495]_  : \new_[17880]_ ;
  assign n2300 = \new_[15949]_  ? \new_[5495]_  : \new_[19023]_ ;
  assign n2305 = \new_[19070]_  ? \new_[5495]_  : \new_[17749]_ ;
  assign n2310 = \new_[18789]_  ? \new_[5495]_  : \new_[17529]_ ;
  assign n2315 = \new_[17866]_  ? \new_[5495]_  : \new_[5055]_ ;
  assign n2320 = \new_[17749]_  ? \new_[5495]_  : \new_[18002]_ ;
  assign n2360 = \new_[17529]_  ? \new_[5495]_  : \new_[18677]_ ;
  assign n2325 = \new_[5055]_  ? \new_[5495]_  : \new_[18512]_ ;
  assign n2330 = \new_[18002]_  ? \new_[5495]_  : n17060;
  assign n2335 = \new_[18677]_  ? \new_[5495]_  : n17000;
  assign n2340 = \new_[18512]_  ? \new_[5495]_  : n17030;
  assign n2345 = \new_[17106]_  ? \new_[5495]_  : \new_[19070]_ ;
  assign n2350 = \new_[17243]_  ? \new_[5495]_  : \new_[18789]_ ;
  assign n2355 = \new_[17826]_  ? \new_[5495]_  : \new_[17866]_ ;
  assign \new_[5191]_  = ~\new_[5423]_  & ~\new_[6936]_ ;
  assign \new_[5192]_  = ~\new_[5424]_  & ~\new_[6936]_ ;
  assign \new_[5193]_  = ~\new_[5425]_  & ~\new_[6936]_ ;
  assign \new_[5194]_  = ~\new_[5426]_  & ~\new_[6936]_ ;
  assign \new_[5195]_  = ~\new_[5427]_  & ~\new_[6936]_ ;
  assign \new_[5196]_  = ~\new_[5428]_  & ~\new_[6936]_ ;
  assign \new_[5197]_  = ~\new_[5429]_  & ~\new_[6936]_ ;
  assign \new_[5198]_  = ~\new_[6936]_  & (~\new_[5505]_  | ~\new_[11139]_ );
  assign \new_[5199]_  = ~\new_[5435]_  & ~\new_[13807]_ ;
  assign \new_[5200]_  = ~\new_[6936]_  & (~\new_[5506]_  | ~\new_[11140]_ );
  assign \new_[5201]_  = ~\new_[6936]_  & (~\new_[5507]_  | ~\new_[11141]_ );
  assign \new_[5202]_  = ~\new_[6936]_  & (~\new_[5508]_  | ~\new_[11142]_ );
  assign \new_[5203]_  = ~\new_[6936]_  & (~\new_[5509]_  | ~\new_[10831]_ );
  assign \new_[5204]_  = ~\new_[6936]_  & (~\new_[5510]_  | ~\new_[11143]_ );
  assign \new_[5205]_  = ~\new_[5437]_  & ~\new_[6936]_ ;
  assign \new_[5206]_  = ~\new_[5438]_  & ~\new_[6936]_ ;
  assign \new_[5207]_  = ~\new_[5439]_  & ~\new_[6936]_ ;
  assign \new_[5208]_  = ~\new_[6936]_  & (~\new_[5512]_  | ~\new_[11178]_ );
  assign \new_[5209]_  = ~\new_[5430]_  & ~\new_[6936]_ ;
  assign \new_[5210]_  = ~\new_[5436]_  & ~\new_[13807]_ ;
  assign \new_[5211]_  = ~\new_[5431]_  & ~\new_[6936]_ ;
  assign \new_[5212]_  = ~\new_[5440]_  & ~\new_[6936]_ ;
  assign \new_[5213]_  = ~\new_[5432]_  & ~\new_[6936]_ ;
  assign \new_[5214]_  = ~\new_[5433]_  & ~\new_[6936]_ ;
  assign \new_[5215]_  = ~\new_[5434]_  & ~\new_[6936]_ ;
  assign \new_[5216]_  = ~\new_[6936]_  & (~\new_[5504]_  | ~\new_[11889]_ );
  assign \new_[5217]_  = ~\new_[15004]_  & (~\new_[5520]_  | ~\new_[17279]_ );
  assign \new_[5218]_  = ~\new_[5417]_  | ~\new_[16093]_ ;
  assign \new_[5219]_  = ~\new_[5418]_  | ~\new_[16090]_ ;
  assign \new_[5220]_  = ~\new_[5419]_  | ~\new_[16389]_ ;
  assign n2085 = ~\new_[5420]_  | (~\new_[14197]_  & ~\new_[16782]_ );
  assign n2090 = ~\new_[5421]_  | (~\new_[13613]_  & ~\new_[16782]_ );
  assign n2095 = ~\new_[5422]_  | (~\new_[11662]_  & ~\new_[16782]_ );
  assign n2080 = \new_[14239]_  ? \new_[16782]_  : \new_[5550]_ ;
  assign \new_[5225]_  = \new_[5537]_  ? \new_[9903]_  : \new_[5538]_ ;
  assign \new_[5226]_  = \new_[5539]_  ? \new_[17323]_  : \new_[5540]_ ;
  assign \new_[5227]_  = \new_[5541]_  ? \new_[17323]_  : \new_[5542]_ ;
  assign n2100 = \new_[13603]_  ? \new_[16782]_  : \new_[5557]_ ;
  assign n2105 = \new_[18491]_  ? \new_[12189]_  : \new_[5538]_ ;
  assign n2110 = \new_[18224]_  ? \new_[12189]_  : \new_[5540]_ ;
  assign n2400 = \new_[19636]_  ? \new_[12189]_  : \new_[5542]_ ;
  assign n2115 = \new_[19517]_  ? \new_[12189]_  : \new_[5576]_ ;
  assign n2120 = \new_[18261]_  ? \new_[12189]_  : \new_[5577]_ ;
  assign n2125 = \new_[18321]_  ? \new_[12189]_  : \new_[5578]_ ;
  assign n2130 = \new_[19530]_  ? \new_[12189]_  : \new_[5579]_ ;
  assign n2135 = \new_[18951]_  ? \new_[12189]_  : \new_[5580]_ ;
  assign n2140 = \new_[19318]_  ? \new_[12189]_  : \new_[5581]_ ;
  assign n2145 = \new_[19178]_  ? \new_[12189]_  : \new_[5582]_ ;
  assign n2395 = \new_[18308]_  ? \new_[12189]_  : \new_[5583]_ ;
  assign n2150 = \new_[19111]_  ? \new_[12189]_  : \new_[5584]_ ;
  assign n2155 = \new_[17867]_  ? \new_[12189]_  : \new_[5543]_ ;
  assign n2160 = \new_[17840]_  ? \new_[12189]_  : \new_[5585]_ ;
  assign n2385 = \new_[19083]_  ? \new_[12189]_  : \new_[5586]_ ;
  assign n2165 = \new_[18946]_  ? \new_[12189]_  : \new_[5587]_ ;
  assign n2170 = \new_[18337]_  ? \new_[12189]_  : \new_[5588]_ ;
  assign n2390 = \new_[19845]_  ? \new_[12189]_  : \new_[5589]_ ;
  assign n2175 = \new_[19341]_  ? \new_[12189]_  : \new_[5590]_ ;
  assign n2180 = \new_[19381]_  ? \new_[12189]_  : \new_[5591]_ ;
  assign n2185 = \new_[19362]_  ? \new_[12189]_  : \new_[5592]_ ;
  assign n2190 = \new_[18425]_  ? \new_[12189]_  : \new_[5593]_ ;
  assign n2195 = \new_[18435]_  ? \new_[12189]_  : \new_[5594]_ ;
  assign n2200 = \new_[18565]_  ? \new_[12189]_  : \new_[5595]_ ;
  assign n2205 = \new_[18664]_  ? \new_[12189]_  : \new_[5547]_ ;
  assign n2210 = \new_[18481]_  ? \new_[12189]_  : \new_[5596]_ ;
  assign n2375 = \new_[18926]_  ? \new_[12189]_  : \new_[5597]_ ;
  assign n2215 = \new_[19226]_  ? \new_[12189]_  : \new_[5598]_ ;
  assign n2220 = \new_[18517]_  ? \new_[12189]_  : \new_[5599]_ ;
  assign n2225 = \new_[19497]_  ? \new_[12189]_  : \new_[5600]_ ;
  assign n2380 = \new_[19608]_  ? \new_[12189]_  : \new_[5601]_ ;
  assign n2260 = \new_[14870]_  ? \new_[16782]_  : \new_[5551]_ ;
  assign n2230 = \new_[14199]_  ? \new_[16782]_  : \new_[5552]_ ;
  assign n2235 = \new_[14214]_  ? \new_[16782]_  : \new_[5554]_ ;
  assign n2240 = \new_[13791]_  ? \new_[16782]_  : \new_[5556]_ ;
  assign n2245 = \new_[14883]_  ? \new_[16782]_  : \new_[5560]_ ;
  assign n2250 = \new_[14884]_  ? \new_[16782]_  : \new_[5572]_ ;
  assign n2255 = \new_[14972]_  ? \new_[16782]_  : \new_[5574]_ ;
  assign n2365 = \new_[14882]_  ? \new_[16782]_  : \new_[5575]_ ;
  assign n2265 = \new_[5045]_  ? \new_[16782]_  : \new_[5545]_ ;
  assign n2270 = \new_[5046]_  ? \new_[16782]_  : \new_[5546]_ ;
  assign n2275 = \new_[5047]_  ? \new_[16782]_  : \new_[5544]_ ;
  assign n2280 = \new_[5048]_  ? \new_[16782]_  : \new_[5548]_ ;
  assign n2370 = \new_[5096]_  ? \new_[16782]_  : \new_[5549]_ ;
  assign \new_[5273]_  = ~\new_[5445]_  | ~\new_[17646]_ ;
  assign \new_[5274]_  = ~\new_[5325]_ ;
  assign \new_[5275]_  = ~\new_[5446]_  & ~\new_[20153]_ ;
  assign \new_[5276]_  = ~\new_[5447]_  & ~\new_[20153]_ ;
  assign \new_[5277]_  = ~\new_[5448]_  & ~\new_[20153]_ ;
  assign \new_[5278]_  = ~\new_[5449]_  | ~\new_[16782]_ ;
  assign \new_[5279]_  = \new_[12057]_  ? \new_[16658]_  : \new_[5626]_ ;
  assign \new_[5280]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[15] ;
  assign \new_[5281]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[24] ;
  assign \new_[5282]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[25] ;
  assign \new_[5283]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[27] ;
  assign \new_[5284]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[2] ;
  assign \new_[5285]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[36] ;
  assign \new_[5286]_  = ~\new_[5467]_  & (~\new_[5466]_  | ~\wbm_sel_o[0] );
  assign \new_[5287]_  = ~\new_[5468]_  & (~\new_[5466]_  | ~\wbm_sel_o[1] );
  assign \new_[5288]_  = ~\new_[5469]_  & (~\new_[5466]_  | ~\wbm_sel_o[2] );
  assign \new_[5289]_  = ~\new_[5470]_  & (~\new_[5466]_  | ~\wbm_sel_o[3] );
  assign n2285 = \new_[19869]_  ^ \new_[5493]_ ;
  assign n2290 = \new_[18681]_  ? \new_[5493]_  : \new_[18046]_ ;
  assign \new_[5292]_  = ~\new_[17075]_  | ~\new_[5493]_ ;
  assign n2420 = ~\new_[20313]_  & ~n6835;
  assign n2425 = ~\new_[20539]_ ;
  assign \new_[5295]_  = ~\new_[20539]_ ;
  assign n2430 = ~\new_[20231]_ ;
  assign \new_[5297]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37] ;
  assign \new_[5298]_  = ~\new_[20229]_  | ~\new_[5495]_ ;
  assign \new_[5299]_  = ~\new_[20311]_ ;
  assign n2405 = \new_[18534]_  ? \new_[12189]_  : \new_[5642]_ ;
  assign n2410 = \new_[18934]_  ? \new_[12189]_  : \new_[5644]_ ;
  assign n2500 = \new_[18462]_  ? \new_[12189]_  : \new_[5643]_ ;
  assign \new_[5303]_  = ~\new_[5515]_  | ~\new_[17279]_ ;
  assign \new_[5304]_  = ~\new_[5516]_  | ~\new_[17279]_ ;
  assign \new_[5305]_  = ~\new_[5517]_  | ~\new_[17279]_ ;
  assign \new_[5306]_  = ~\new_[5518]_  | ~\new_[17279]_ ;
  assign \new_[5307]_  = ~\new_[5519]_  | ~\new_[17646]_ ;
  assign \new_[5308]_  = ~\new_[5521]_  | ~\new_[17279]_ ;
  assign \new_[5309]_  = ~\new_[5522]_  | ~\new_[17279]_ ;
  assign \new_[5310]_  = ~\new_[5523]_  | ~\new_[17279]_ ;
  assign \new_[5311]_  = ~\new_[5524]_  | ~\new_[17646]_ ;
  assign \new_[5312]_  = ~\new_[5525]_  | ~\new_[17279]_ ;
  assign \new_[5313]_  = ~\new_[5526]_  | ~\new_[17279]_ ;
  assign \new_[5314]_  = ~\new_[5527]_  | ~\new_[17279]_ ;
  assign \new_[5315]_  = ~\new_[5528]_  | ~\new_[17279]_ ;
  assign \new_[5316]_  = ~\new_[5529]_  | ~\new_[17279]_ ;
  assign \new_[5317]_  = ~\new_[5530]_  | ~\new_[17279]_ ;
  assign \new_[5318]_  = ~\new_[5531]_  | ~\new_[17279]_ ;
  assign \new_[5319]_  = ~\new_[5532]_  | ~\new_[17279]_ ;
  assign \new_[5320]_  = ~\new_[5533]_  | ~\new_[17279]_ ;
  assign \new_[5321]_  = ~\new_[5534]_  | ~\new_[17279]_ ;
  assign \new_[5322]_  = ~\new_[5535]_  | ~\new_[17279]_ ;
  assign \new_[5323]_  = ~\new_[5536]_  | ~\new_[17646]_ ;
  assign \new_[5324]_  = \\pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_reg[1] ;
  assign \new_[5325]_  = ~\new_[5514]_  | ~\new_[17549]_ ;
  assign \new_[5326]_  = ~\new_[5602]_  | ~\new_[17646]_ ;
  assign \new_[5327]_  = ~\new_[5603]_  | ~\new_[17279]_ ;
  assign \new_[5328]_  = ~\new_[5604]_  | ~\new_[17279]_ ;
  assign \new_[5329]_  = ~\new_[5605]_  | ~\new_[17279]_ ;
  assign \new_[5330]_  = ~\new_[5606]_  | ~\new_[17279]_ ;
  assign \new_[5331]_  = ~\new_[5607]_  | ~\new_[17279]_ ;
  assign \new_[5332]_  = ~\new_[5553]_  | ~\new_[16782]_ ;
  assign \new_[5333]_  = ~\new_[5555]_  | ~\new_[16782]_ ;
  assign \new_[5334]_  = ~\new_[5558]_  | ~\new_[16782]_ ;
  assign \new_[5335]_  = ~\new_[5559]_  | ~\new_[16782]_ ;
  assign \new_[5336]_  = ~\new_[5561]_  | ~\new_[16782]_ ;
  assign \new_[5337]_  = ~\new_[5562]_  | ~\new_[16782]_ ;
  assign \new_[5338]_  = ~\new_[5563]_  | ~\new_[16782]_ ;
  assign \new_[5339]_  = ~\new_[5564]_  | ~\new_[16782]_ ;
  assign \new_[5340]_  = ~\new_[5565]_  | ~\new_[16782]_ ;
  assign \new_[5341]_  = ~\new_[5566]_  | ~\new_[16782]_ ;
  assign \new_[5342]_  = ~\new_[5567]_  | ~\new_[16782]_ ;
  assign \new_[5343]_  = ~\new_[5568]_  | ~\new_[16782]_ ;
  assign \new_[5344]_  = ~\new_[5569]_  | ~\new_[16782]_ ;
  assign \new_[5345]_  = ~\new_[5570]_  | ~\new_[16782]_ ;
  assign \new_[5346]_  = ~\new_[5571]_  | ~\new_[16782]_ ;
  assign \new_[5347]_  = ~\new_[5573]_  | ~\new_[16782]_ ;
  assign \new_[5348]_  = ~\new_[10952]_  & (~\new_[5648]_  | ~\new_[16433]_ );
  assign \new_[5349]_  = (~\new_[11848]_  | ~\new_[6162]_ ) & (~\new_[5646]_  | ~\new_[5986]_ );
  assign \new_[5350]_  = \new_[13434]_  ? \new_[16434]_  : \new_[5647]_ ;
  assign \new_[5351]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[0] ;
  assign \new_[5352]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[12] ;
  assign \new_[5353]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[13] ;
  assign \new_[5354]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[14] ;
  assign \new_[5355]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[17] ;
  assign \new_[5356]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[20] ;
  assign \new_[5357]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[23] ;
  assign \new_[5358]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[26] ;
  assign \new_[5359]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[28] ;
  assign \new_[5360]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[29] ;
  assign \new_[5361]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[31] ;
  assign \new_[5362]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[3] ;
  assign \new_[5363]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[4] ;
  assign \new_[5364]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[7] ;
  assign \new_[5365]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[8] ;
  assign \new_[5366]_  = \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[9] ;
  assign n2415 = ~\new_[19889]_ ;
  assign \new_[5368]_  = ~\new_[5464]_  | ~\wbm_cti_o[0] ;
  assign \new_[5369]_  = ~\new_[5464]_  | ~\wbm_cti_o[2] ;
  assign n2440 = ~\new_[5466]_  & ~n6835;
  assign n2460 = ~\new_[5456]_  | ~\new_[5673]_ ;
  assign n2465 = ~\new_[20362]_  | ~\new_[5674]_ ;
  assign n2470 = ~\new_[5457]_  | ~\new_[5783]_ ;
  assign n2475 = ~\new_[5458]_  | ~\new_[5678]_ ;
  assign n2480 = ~\new_[5459]_  | ~\new_[5675]_ ;
  assign n2485 = ~\new_[20368]_  | ~\new_[5684]_ ;
  assign n2490 = ~\new_[5460]_  | ~\new_[5788]_ ;
  assign n2495 = ~\new_[5461]_  | ~\new_[5688]_ ;
  assign n2445 = ~\new_[5462]_  | ~\new_[5692]_ ;
  assign n2450 = ~\new_[5463]_  | ~\new_[5693]_ ;
  assign n2455 = ~\new_[20355]_  | ~\new_[5698]_ ;
  assign \new_[5382]_  = ~\new_[5631]_  | ~\wbm_dat_o[0] ;
  assign \new_[5383]_  = ~\new_[5631]_  | ~\wbm_dat_o[11] ;
  assign \new_[5384]_  = ~\new_[5631]_  | ~\wbm_dat_o[12] ;
  assign \new_[5385]_  = ~\new_[5631]_  | ~\wbm_dat_o[13] ;
  assign \new_[5386]_  = ~\new_[5631]_  | ~\wbm_dat_o[14] ;
  assign \new_[5387]_  = ~\new_[5631]_  | ~\wbm_dat_o[15] ;
  assign \new_[5388]_  = ~\new_[5631]_  | ~\wbm_dat_o[16] ;
  assign \new_[5389]_  = ~\new_[5631]_  | ~\wbm_dat_o[17] ;
  assign \new_[5390]_  = ~\new_[5631]_  | ~\wbm_dat_o[18] ;
  assign \new_[5391]_  = ~\new_[5632]_  | ~\wbm_dat_o[19] ;
  assign \new_[5392]_  = ~\new_[5632]_  | ~\wbm_dat_o[1] ;
  assign \new_[5393]_  = ~\new_[5632]_  | ~\wbm_dat_o[20] ;
  assign \new_[5394]_  = ~\new_[5632]_  | ~\wbm_dat_o[21] ;
  assign \new_[5395]_  = ~\new_[5632]_  | ~\wbm_dat_o[23] ;
  assign \new_[5396]_  = ~\new_[5632]_  | ~\wbm_dat_o[24] ;
  assign \new_[5397]_  = ~\new_[5632]_  | ~\wbm_dat_o[25] ;
  assign \new_[5398]_  = ~\new_[5632]_  | ~\wbm_dat_o[26] ;
  assign \new_[5399]_  = ~\new_[5632]_  | ~\wbm_dat_o[27] ;
  assign \new_[5400]_  = ~\new_[5632]_  | ~\wbm_dat_o[28] ;
  assign \new_[5401]_  = ~\new_[5632]_  | ~\wbm_dat_o[29] ;
  assign \new_[5402]_  = ~\new_[5632]_  | ~\wbm_dat_o[2] ;
  assign \new_[5403]_  = ~\new_[5632]_  | ~\wbm_dat_o[30] ;
  assign \new_[5404]_  = ~\new_[5632]_  | ~\wbm_dat_o[31] ;
  assign \new_[5405]_  = ~\new_[5632]_  | ~\wbm_dat_o[3] ;
  assign \new_[5406]_  = ~\new_[5631]_  | ~\wbm_dat_o[4] ;
  assign \new_[5407]_  = ~\new_[5631]_  | ~\wbm_dat_o[5] ;
  assign \new_[5408]_  = ~\new_[5631]_  | ~\wbm_dat_o[6] ;
  assign \new_[5409]_  = ~\new_[5631]_  | ~\wbm_dat_o[7] ;
  assign \new_[5410]_  = ~\new_[5631]_  | ~\wbm_dat_o[8] ;
  assign \new_[5411]_  = ~\new_[5631]_  | ~\wbm_dat_o[9] ;
  assign \new_[5412]_  = ~\new_[5464]_ ;
  assign \new_[5413]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[15] ;
  assign \new_[5414]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[25] ;
  assign \new_[5415]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[7] ;
  assign \new_[5416]_  = ~\new_[5494]_ ;
  assign \new_[5417]_  = ~\new_[5636]_  | ~\new_[17646]_ ;
  assign \new_[5418]_  = ~\new_[5637]_  | ~\new_[17646]_ ;
  assign \new_[5419]_  = ~\new_[5638]_  | ~\new_[17279]_ ;
  assign \new_[5420]_  = ~\new_[5639]_  | ~\new_[16782]_ ;
  assign \new_[5421]_  = ~\new_[5640]_  | ~\new_[16782]_ ;
  assign \new_[5422]_  = ~\new_[5641]_  | ~\new_[16782]_ ;
  assign \new_[5423]_  = ~\new_[10829]_  & (~\new_[5712]_  | ~\new_[16434]_ );
  assign \new_[5424]_  = ~\new_[12394]_  & (~\new_[5713]_  | ~\new_[16433]_ );
  assign \new_[5425]_  = ~\new_[12395]_  & (~\new_[5714]_  | ~\new_[16434]_ );
  assign \new_[5426]_  = ~\new_[10955]_  & (~\new_[5715]_  | ~\new_[16434]_ );
  assign \new_[5427]_  = ~\new_[12396]_  & (~\new_[5716]_  | ~\new_[16433]_ );
  assign \new_[5428]_  = ~\new_[12397]_  & (~\new_[5717]_  | ~\new_[16433]_ );
  assign \new_[5429]_  = ~\new_[12398]_  & (~\new_[5718]_  | ~\new_[16433]_ );
  assign \new_[5430]_  = ~\new_[10956]_  & (~\new_[5733]_  | ~\new_[16433]_ );
  assign \new_[5431]_  = ~\new_[11873]_  & (~\new_[5735]_  | ~\new_[16434]_ );
  assign \new_[5432]_  = ~\new_[10828]_  & (~\new_[5737]_  | ~\new_[16434]_ );
  assign \new_[5433]_  = ~\new_[10950]_  & (~\new_[5738]_  | ~\new_[16433]_ );
  assign \new_[5434]_  = ~\new_[10951]_  & (~\new_[5739]_  | ~\new_[16434]_ );
  assign \new_[5435]_  = (~\new_[11177]_  | ~\new_[6162]_ ) & (~\new_[5721]_  | ~\new_[5986]_ );
  assign \new_[5436]_  = (~\new_[5734]_  | ~\new_[5986]_ ) & (~\new_[10457]_  | ~\new_[6162]_ );
  assign \new_[5437]_  = ~\new_[12465]_  & (~\new_[5728]_  | ~\new_[16433]_ );
  assign \new_[5438]_  = ~\new_[12466]_  & (~\new_[5730]_  | ~\new_[16433]_ );
  assign \new_[5439]_  = ~\new_[12438]_  & (~\new_[5731]_  | ~\new_[16433]_ );
  assign \new_[5440]_  = ~\new_[12387]_  & (~\new_[5736]_  | ~\new_[16433]_ );
  assign \new_[5441]_  = \new_[17958]_  ? \new_[5711]_  : pci_par_i;
  assign \new_[5442]_  = \new_[13435]_  ? \new_[16658]_  : \new_[5729]_ ;
  assign \new_[5443]_  = ~parity_checker_check_perr_reg;
  assign \new_[5444]_  = ~\new_[5513]_ ;
  assign \new_[5445]_  = \new_[5671]_  ? \new_[15498]_  : \new_[18362]_ ;
  assign \new_[5446]_  = ~\new_[5538]_ ;
  assign \new_[5447]_  = ~\new_[5540]_ ;
  assign \new_[5448]_  = ~\new_[5542]_ ;
  assign \new_[5449]_  = \new_[5671]_  ? \new_[20186]_  : \new_[19366]_ ;
  assign \new_[5450]_  = \new_[5671]_  ? \new_[11961]_  : n17410;
  assign n2510 = ~\new_[5821]_  | ~\new_[5822]_  | ~\new_[5633]_  | ~\new_[6043]_ ;
  assign n2520 = ~\new_[5968]_  | ~\new_[5679]_  | ~\new_[5704]_ ;
  assign n2525 = ~\new_[5835]_  | ~\new_[5836]_  | ~\new_[5634]_  | ~\new_[5970]_ ;
  assign n2530 = ~\new_[6081]_  | ~\new_[5786]_  | ~\new_[5705]_ ;
  assign n2505 = ~\new_[5882]_  | ~\new_[5883]_  | ~\new_[5635]_  | ~\new_[5985]_ ;
  assign \new_[5456]_  = ~\new_[5700]_  & ~\new_[6006]_ ;
  assign \new_[5457]_  = ~\new_[5961]_  & ~\new_[5701]_ ;
  assign \new_[5458]_  = ~\new_[5964]_  & ~\new_[5702]_ ;
  assign \new_[5459]_  = ~\new_[5965]_  & ~\new_[5703]_ ;
  assign \new_[5460]_  = ~\new_[6101]_  & ~\new_[5706]_ ;
  assign \new_[5461]_  = ~\new_[6258]_  & ~\new_[5707]_ ;
  assign \new_[5462]_  = ~\new_[6131]_  & ~\new_[5708]_ ;
  assign \new_[5463]_  = ~\new_[5981]_  & ~\new_[5709]_ ;
  assign \new_[5464]_  = \new_[20315]_  & \new_[5790]_ ;
  assign \new_[5465]_  = \new_[20315]_  | \new_[5790]_ ;
  assign \new_[5466]_  = \new_[20315]_  & \new_[5801]_ ;
  assign \new_[5467]_  = ~\new_[5699]_  & ~\new_[18583]_ ;
  assign \new_[5468]_  = ~\new_[5699]_  & ~\new_[18300]_ ;
  assign \new_[5469]_  = ~\new_[5699]_  & ~\new_[19074]_ ;
  assign \new_[5470]_  = ~\new_[5699]_  & ~\new_[19634]_ ;
  assign \new_[5471]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[0] ;
  assign \new_[5472]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[10] ;
  assign \new_[5473]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[11] ;
  assign \new_[5474]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[13] ;
  assign \new_[5475]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[14] ;
  assign \new_[5476]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[17] ;
  assign \new_[5477]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[18] ;
  assign \new_[5478]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[19] ;
  assign \new_[5479]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[21] ;
  assign \new_[5480]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[22] ;
  assign \new_[5481]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[20] ;
  assign \new_[5482]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[24] ;
  assign \new_[5483]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[26] ;
  assign \new_[5484]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[28] ;
  assign \new_[5485]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[29] ;
  assign \new_[5486]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[2] ;
  assign \new_[5487]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[31] ;
  assign \new_[5488]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[3] ;
  assign \new_[5489]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[4] ;
  assign \new_[5490]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[6] ;
  assign \new_[5491]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[8] ;
  assign \new_[5492]_  = ~\new_[5630]_ ;
  assign \new_[5493]_  = \new_[5710]_  & \new_[4040]_ ;
  assign \new_[5494]_  = \new_[20311]_ ;
  assign \new_[5495]_  = ~\new_[5710]_ ;
  assign \new_[5496]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[9] ;
  assign \new_[5497]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[5] ;
  assign \new_[5498]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[30] ;
  assign \new_[5499]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[27] ;
  assign \new_[5500]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[23] ;
  assign \new_[5501]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[12] ;
  assign \new_[5502]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[1] ;
  assign \new_[5503]_  = ~\\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[16] ;
  assign \new_[5504]_  = ~\new_[5719]_  | ~\new_[16658]_ ;
  assign \new_[5505]_  = ~\new_[5720]_  | ~\new_[16658]_ ;
  assign \new_[5506]_  = ~\new_[5722]_  | ~\new_[16658]_ ;
  assign \new_[5507]_  = ~\new_[5723]_  | ~\new_[16658]_ ;
  assign \new_[5508]_  = ~\new_[5724]_  | ~\new_[16658]_ ;
  assign \new_[5509]_  = ~\new_[5725]_  | ~\new_[16658]_ ;
  assign \new_[5510]_  = ~\new_[5726]_  | ~\new_[16658]_ ;
  assign \new_[5511]_  = ~\new_[5727]_  | ~\new_[5986]_ ;
  assign \new_[5512]_  = ~\new_[5732]_  | ~\new_[16658]_ ;
  assign \new_[5513]_  = ~n2965 | ~\new_[5711]_  | ~\new_[17007]_ ;
  assign \new_[5514]_  = \new_[5779]_  ? \new_[20413]_  : \new_[5324]_ ;
  assign \new_[5515]_  = \new_[5748]_  ? \new_[15498]_  : \new_[19178]_ ;
  assign \new_[5516]_  = \new_[5749]_  ? \new_[15498]_  : \new_[18308]_ ;
  assign \new_[5517]_  = \new_[5750]_  ? \new_[15498]_  : \new_[19111]_ ;
  assign \new_[5518]_  = \new_[5751]_  ? \new_[15498]_  : \new_[17867]_ ;
  assign \new_[5519]_  = \new_[5752]_  ? \new_[15498]_  : \new_[17840]_ ;
  assign \new_[5520]_  = \new_[5753]_  ? \new_[15498]_  : \new_[19083]_ ;
  assign \new_[5521]_  = \new_[5754]_  ? \new_[15498]_  : \new_[18946]_ ;
  assign \new_[5522]_  = \new_[5755]_  ? \new_[15498]_  : \new_[18337]_ ;
  assign \new_[5523]_  = \new_[5756]_  ? \new_[15498]_  : \new_[19845]_ ;
  assign \new_[5524]_  = \new_[5757]_  ? \new_[15498]_  : \new_[19341]_ ;
  assign \new_[5525]_  = \new_[5758]_  ? \new_[15498]_  : \new_[19381]_ ;
  assign \new_[5526]_  = \new_[5759]_  ? \new_[15498]_  : \new_[19362]_ ;
  assign \new_[5527]_  = \new_[5760]_  ? \new_[15498]_  : \new_[18425]_ ;
  assign \new_[5528]_  = \new_[5761]_  ? \new_[15498]_  : \new_[18435]_ ;
  assign \new_[5529]_  = \new_[5762]_  ? \new_[15498]_  : \new_[18565]_ ;
  assign \new_[5530]_  = \new_[5763]_  ? \new_[15498]_  : \new_[18664]_ ;
  assign \new_[5531]_  = \new_[5764]_  ? \new_[15498]_  : \new_[18481]_ ;
  assign \new_[5532]_  = \new_[5765]_  ? \new_[15498]_  : \new_[18926]_ ;
  assign \new_[5533]_  = \new_[5766]_  ? \new_[15498]_  : \new_[19226]_ ;
  assign \new_[5534]_  = \new_[5767]_  ? \new_[15498]_  : \new_[18517]_ ;
  assign \new_[5535]_  = \new_[5768]_  ? \new_[15498]_  : \new_[19497]_ ;
  assign \new_[5536]_  = \new_[5769]_  ? \new_[15498]_  : \new_[19608]_ ;
  assign \new_[5537]_  = \new_[5770]_  ? \new_[15498]_  : \new_[18491]_ ;
  assign \new_[5538]_  = \new_[5770]_  ? \new_[11961]_  : \new_[17687]_ ;
  assign \new_[5539]_  = \new_[5771]_  ? \new_[15498]_  : \new_[18224]_ ;
  assign \new_[5540]_  = \new_[5771]_  ? \new_[11961]_  : \new_[17761]_ ;
  assign \new_[5541]_  = \new_[5772]_  ? \new_[15498]_  : \new_[19636]_ ;
  assign \new_[5542]_  = \new_[5772]_  ? \new_[11961]_  : \new_[17536]_ ;
  assign \new_[5543]_  = \new_[5751]_  ? \new_[11961]_  : n17100;
  assign \new_[5544]_  = \new_[5770]_  ? \new_[20186]_  : \new_[18190]_ ;
  assign \new_[5545]_  = \new_[5771]_  ? \new_[20186]_  : \new_[17984]_ ;
  assign \new_[5546]_  = \new_[5772]_  ? \new_[20186]_  : \new_[19048]_ ;
  assign \new_[5547]_  = \new_[5763]_  ? \new_[11961]_  : n17110;
  assign \new_[5548]_  = \new_[5773]_  ? \new_[20186]_  : \new_[18020]_ ;
  assign \new_[5549]_  = \new_[5753]_  ? \new_[20186]_  : \new_[18917]_ ;
  assign \new_[5550]_  = \new_[5761]_  ? \new_[20186]_  : \new_[19296]_ ;
  assign \new_[5551]_  = \new_[5776]_  ? \new_[20186]_  : \new_[17810]_ ;
  assign \new_[5552]_  = \new_[5777]_  ? \new_[20186]_  : \new_[19563]_ ;
  assign \new_[5553]_  = \new_[5778]_  ? \new_[20186]_  : \new_[19564]_ ;
  assign \new_[5554]_  = \new_[5748]_  ? \new_[20186]_  : \new_[17816]_ ;
  assign \new_[5555]_  = \new_[5749]_  ? \new_[20186]_  : \new_[17891]_ ;
  assign \new_[5556]_  = \new_[5750]_  ? \new_[20186]_  : \new_[18779]_ ;
  assign \new_[5557]_  = \new_[5751]_  ? \new_[20186]_  : \new_[19578]_ ;
  assign \new_[5558]_  = \new_[5752]_  ? \new_[20186]_  : \new_[18987]_ ;
  assign \new_[5559]_  = \new_[5754]_  ? \new_[20186]_  : \new_[18568]_ ;
  assign \new_[5560]_  = \new_[5763]_  ? \new_[20186]_  : \new_[18116]_ ;
  assign \new_[5561]_  = \new_[5755]_  ? \new_[20186]_  : \new_[19572]_ ;
  assign \new_[5562]_  = \new_[5756]_  ? \new_[20186]_  : \new_[19576]_ ;
  assign \new_[5563]_  = \new_[5757]_  ? \new_[20186]_  : \new_[18150]_ ;
  assign \new_[5564]_  = \new_[5758]_  ? \new_[20186]_  : \new_[19349]_ ;
  assign \new_[5565]_  = \new_[5759]_  ? \new_[20186]_  : \new_[18357]_ ;
  assign \new_[5566]_  = \new_[5760]_  ? \new_[20186]_  : \new_[19282]_ ;
  assign \new_[5567]_  = \new_[5762]_  ? \new_[20186]_  : \new_[17854]_ ;
  assign \new_[5568]_  = \new_[5764]_  ? \new_[20186]_  : \new_[19614]_ ;
  assign \new_[5569]_  = \new_[5765]_  ? \new_[20186]_  : \new_[17844]_ ;
  assign \new_[5570]_  = \new_[5766]_  ? \new_[20186]_  : \new_[18748]_ ;
  assign \new_[5571]_  = \new_[5767]_  ? \new_[20186]_  : \new_[19604]_ ;
  assign \new_[5572]_  = \new_[5768]_  ? \new_[20186]_  : \new_[17841]_ ;
  assign \new_[5573]_  = \new_[5769]_  ? \new_[20186]_  : \new_[18047]_ ;
  assign \new_[5574]_  = \new_[5774]_  ? \new_[20186]_  : \new_[17876]_ ;
  assign \new_[5575]_  = \new_[5775]_  ? \new_[20186]_  : \new_[17821]_ ;
  assign \new_[5576]_  = \new_[5773]_  ? \new_[11961]_  : n17200;
  assign \new_[5577]_  = \new_[5774]_  ? \new_[11961]_  : n17460;
  assign \new_[5578]_  = \new_[5775]_  ? \new_[11961]_  : n17135;
  assign \new_[5579]_  = \new_[5776]_  ? \new_[11961]_  : n17385;
  assign \new_[5580]_  = \new_[5777]_  ? \new_[11961]_  : n17300;
  assign \new_[5581]_  = \new_[5778]_  ? \new_[11961]_  : n17155;
  assign \new_[5582]_  = \new_[5748]_  ? \new_[11961]_  : n17150;
  assign \new_[5583]_  = \new_[5749]_  ? \new_[11961]_  : n17130;
  assign \new_[5584]_  = \new_[5750]_  ? \new_[11961]_  : n17520;
  assign \new_[5585]_  = \new_[5752]_  ? \new_[11961]_  : n17255;
  assign \new_[5586]_  = \new_[5753]_  ? \new_[11961]_  : n17145;
  assign \new_[5587]_  = \new_[5754]_  ? \new_[11961]_  : n17375;
  assign \new_[5588]_  = \new_[5755]_  ? \new_[11961]_  : n17265;
  assign \new_[5589]_  = \new_[5756]_  ? \new_[11961]_  : n17260;
  assign \new_[5590]_  = \new_[5757]_  ? \new_[11961]_  : n17275;
  assign \new_[5591]_  = \new_[5758]_  ? \new_[11961]_  : n17240;
  assign \new_[5592]_  = \new_[5759]_  ? \new_[11961]_  : n17270;
  assign \new_[5593]_  = \new_[5760]_  ? \new_[11961]_  : n17245;
  assign \new_[5594]_  = \new_[5761]_  ? \new_[11961]_  : n17140;
  assign \new_[5595]_  = \new_[5762]_  ? \new_[11961]_  : n17105;
  assign \new_[5596]_  = \new_[5764]_  ? \new_[11961]_  : n17115;
  assign \new_[5597]_  = \new_[5765]_  ? \new_[11961]_  : n17290;
  assign \new_[5598]_  = \new_[5766]_  ? \new_[11961]_  : n17125;
  assign \new_[5599]_  = \new_[5767]_  ? \new_[11961]_  : n17400;
  assign \new_[5600]_  = \new_[5768]_  ? \new_[11961]_  : n17195;
  assign \new_[5601]_  = \new_[5769]_  ? \new_[11961]_  : n17525;
  assign \new_[5602]_  = \new_[5773]_  ? \new_[15498]_  : \new_[19517]_ ;
  assign \new_[5603]_  = \new_[5774]_  ? \new_[15498]_  : \new_[18261]_ ;
  assign \new_[5604]_  = \new_[5775]_  ? \new_[15498]_  : \new_[18321]_ ;
  assign \new_[5605]_  = \new_[5776]_  ? \new_[15498]_  : \new_[19530]_ ;
  assign \new_[5606]_  = \new_[5777]_  ? \new_[15498]_  : \new_[18951]_ ;
  assign \new_[5607]_  = \new_[5778]_  ? \new_[15498]_  : \new_[19318]_ ;
  assign n2540 = \new_[5324]_  ? \new_[10827]_  : \new_[5779]_ ;
  assign n2565 = ~\new_[5802]_  | ~\new_[5803]_  | ~\new_[5782]_  | ~\new_[5960]_ ;
  assign n2570 = ~\new_[5810]_  | ~\new_[5811]_  | ~\new_[5784]_  | ~\new_[5963]_ ;
  assign n2575 = ~\new_[5818]_  | ~\new_[5819]_  | ~\new_[5676]_  | ~\new_[5966]_ ;
  assign n2580 = ~\new_[5825]_  | ~\new_[5826]_  | ~\new_[5681]_  | ~\new_[5967]_ ;
  assign n2585 = ~\new_[5830]_  | ~\new_[5831]_  | ~\new_[5680]_  | ~\new_[5969]_ ;
  assign n2590 = ~\new_[5833]_  | ~\new_[5834]_  | ~\new_[5682]_  | ~\new_[6065]_ ;
  assign n2595 = ~\new_[5839]_  | ~\new_[5840]_  | ~\new_[5685]_  | ~\new_[5971]_ ;
  assign n2535 = ~\new_[5843]_  | ~\new_[5844]_  | ~\new_[5686]_  | ~\new_[5972]_ ;
  assign n2600 = ~\new_[5846]_  | ~\new_[5847]_  | ~\new_[5687]_  | ~\new_[5973]_ ;
  assign n2605 = ~\new_[5849]_  | ~\new_[5850]_  | ~\new_[5787]_  | ~\new_[5974]_ ;
  assign n2610 = ~\new_[5856]_  | ~\new_[5857]_  | ~\new_[5689]_  | ~\new_[5976]_ ;
  assign n2615 = ~\new_[5859]_  | ~\new_[5860]_  | ~\new_[5690]_  | ~\new_[5977]_ ;
  assign n2620 = ~\new_[5862]_  | ~\new_[5863]_  | ~\new_[5691]_  | ~\new_[5978]_ ;
  assign n2545 = ~\new_[5865]_  | ~\new_[5866]_  | ~\new_[5789]_  | ~\new_[6126]_ ;
  assign n2550 = ~\new_[5873]_  | ~\new_[5874]_  | ~\new_[5694]_  | ~\new_[5982]_ ;
  assign n2555 = ~\new_[5876]_  | ~\new_[5877]_  | ~\new_[5695]_  | ~\new_[5983]_ ;
  assign n2560 = ~\new_[5879]_  | ~\new_[5880]_  | ~\new_[5696]_  | ~\new_[5984]_ ;
  assign \new_[5626]_  = ~\new_[5672]_  & (~\new_[19075]_  | ~\new_[20413]_ );
  assign n2630 = \new_[18673]_  ? \new_[10827]_  : \new_[5797]_ ;
  assign n2635 = \new_[18598]_  ? \new_[10827]_  : \new_[5799]_ ;
  assign \new_[5629]_  = ~\new_[19874]_  | ~\new_[5790]_ ;
  assign \new_[5630]_  = ~\new_[20313]_ ;
  assign \new_[5631]_  = \new_[20313]_ ;
  assign \new_[5632]_  = \new_[20313]_ ;
  assign \new_[5633]_  = ~\new_[5677]_ ;
  assign \new_[5634]_  = ~\new_[5683]_ ;
  assign \new_[5635]_  = ~\new_[5697]_ ;
  assign \new_[5636]_  = \new_[5792]_  ? \new_[15498]_  : \new_[18534]_ ;
  assign \new_[5637]_  = \new_[5793]_  ? \new_[15498]_  : \new_[18934]_ ;
  assign \new_[5638]_  = \new_[5794]_  ? \new_[15498]_  : \new_[18462]_ ;
  assign \new_[5639]_  = \new_[5792]_  ? \new_[20186]_  : \new_[17863]_ ;
  assign \new_[5640]_  = \new_[5793]_  ? \new_[20186]_  : \new_[19409]_ ;
  assign \new_[5641]_  = \new_[5794]_  ? \new_[20186]_  : \new_[19610]_ ;
  assign \new_[5642]_  = \new_[5792]_  ? \new_[11961]_  : n17210;
  assign \new_[5643]_  = \new_[5794]_  ? \new_[11961]_  : n17530;
  assign \new_[5644]_  = \new_[5793]_  ? \new_[11961]_  : n17120;
  assign n2640 = ~\new_[5711]_ ;
  assign \new_[5646]_  = \new_[5797]_  ? \new_[20413]_  : \new_[18673]_ ;
  assign \new_[5647]_  = \new_[5799]_  ? \new_[20413]_  : \new_[18598]_ ;
  assign \new_[5648]_  = \new_[5798]_  ? \new_[20413]_  : \new_[17831]_ ;
  assign n2625 = \new_[17831]_  ? \new_[10827]_  : \new_[5798]_ ;
  assign n2675 = \new_[18884]_  ? \new_[10827]_  : \new_[5890]_ ;
  assign n2680 = \new_[17882]_  ? \new_[10827]_  : \new_[5892]_ ;
  assign n2780 = \new_[19075]_  ? \new_[10827]_  : \new_[5893]_ ;
  assign n2695 = \new_[18848]_  ? \new_[10827]_  : \new_[5894]_ ;
  assign n2685 = \new_[19639]_  ? \new_[10827]_  : \new_[5895]_ ;
  assign n2690 = \new_[19844]_  ? \new_[10827]_  : \new_[5898]_ ;
  assign n2770 = \new_[18080]_  ? \new_[10827]_  : \new_[5896]_ ;
  assign n2700 = \new_[18521]_  ? \new_[10827]_  : \new_[5897]_ ;
  assign n2705 = \new_[18386]_  ? \new_[10827]_  : \new_[5899]_ ;
  assign n2765 = \new_[18105]_  ? \new_[10827]_  : \new_[5900]_ ;
  assign n2710 = \new_[18480]_  ? \new_[10827]_  : \new_[5901]_ ;
  assign n2715 = \new_[18239]_  ? \new_[10827]_  : \new_[5902]_ ;
  assign n2720 = \new_[18037]_  ? \new_[10827]_  : \new_[5903]_ ;
  assign n2760 = \new_[19849]_  ? \new_[10827]_  : \new_[5904]_ ;
  assign n2725 = \new_[18992]_  ? \new_[10827]_  : \new_[5905]_ ;
  assign n2730 = \new_[19721]_  ? \new_[10827]_  : \new_[5906]_ ;
  assign n2735 = \new_[19042]_  ? \new_[10827]_  : \new_[5907]_ ;
  assign n2755 = \new_[19009]_  ? \new_[10827]_  : \new_[5908]_ ;
  assign n2740 = \new_[18948]_  ? \new_[10827]_  : \new_[5909]_ ;
  assign n2745 = \new_[18936]_  ? \new_[10827]_  : \new_[5910]_ ;
  assign n2750 = \new_[19593]_  ? \new_[10827]_  : \new_[5911]_ ;
  assign \new_[5671]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26] ;
  assign \new_[5672]_  = ~\new_[5796]_  & ~\new_[20413]_ ;
  assign \new_[5673]_  = \new_[5806]_  & \new_[6009]_ ;
  assign \new_[5674]_  = \new_[5807]_  & \new_[6228]_ ;
  assign \new_[5675]_  = \new_[5817]_  & \new_[6034]_ ;
  assign \new_[5676]_  = \new_[5820]_  & \new_[6039]_ ;
  assign \new_[5677]_  = ~\new_[5823]_  | ~\new_[6237]_ ;
  assign \new_[5678]_  = \new_[5814]_  & \new_[6029]_ ;
  assign \new_[5679]_  = \new_[5829]_  & \new_[6056]_ ;
  assign \new_[5680]_  = \new_[5832]_  & \new_[6062]_ ;
  assign \new_[5681]_  = \new_[5827]_  & \new_[6053]_ ;
  assign \new_[5682]_  = ~\new_[5785]_ ;
  assign \new_[5683]_  = ~\new_[5837]_  | ~\new_[6071]_ ;
  assign \new_[5684]_  = \new_[5838]_  & \new_[6077]_ ;
  assign \new_[5685]_  = \new_[5841]_  & \new_[6253]_ ;
  assign \new_[5686]_  = ~\new_[5845]_  & ~\new_[6086]_ ;
  assign \new_[5687]_  = ~\new_[5848]_  & ~\new_[6091]_ ;
  assign \new_[5688]_  = \new_[5855]_  & \new_[6260]_ ;
  assign \new_[5689]_  = \new_[5858]_  & \new_[6111]_ ;
  assign \new_[5690]_  = \new_[5861]_  & \new_[6116]_ ;
  assign \new_[5691]_  = \new_[5864]_  & \new_[6122]_ ;
  assign \new_[5692]_  = ~\new_[5869]_  & ~\new_[5980]_ ;
  assign \new_[5693]_  = ~\new_[5872]_  & ~\new_[6135]_ ;
  assign \new_[5694]_  = \new_[5875]_  & \new_[6139]_ ;
  assign \new_[5695]_  = ~\new_[5878]_  & ~\new_[6144]_ ;
  assign \new_[5696]_  = \new_[5881]_  & \new_[6271]_ ;
  assign \new_[5697]_  = ~\new_[5884]_  | ~\new_[6156]_ ;
  assign \new_[5698]_  = \new_[5885]_  & \new_[6274]_ ;
  assign \new_[5699]_  = ~\new_[5790]_ ;
  assign \new_[5700]_  = ~\new_[5804]_  | ~\new_[5805]_ ;
  assign \new_[5701]_  = ~\new_[5808]_  | ~\new_[5809]_ ;
  assign \new_[5702]_  = ~\new_[5812]_  | ~\new_[5813]_ ;
  assign \new_[5703]_  = ~\new_[5815]_  | ~\new_[5816]_ ;
  assign \new_[5704]_  = ~\new_[5828]_  & ~\new_[5953]_ ;
  assign \new_[5705]_  = ~\new_[5842]_  & ~\new_[5955]_ ;
  assign \new_[5706]_  = ~\new_[5851]_  | ~\new_[5852]_ ;
  assign \new_[5707]_  = ~\new_[5853]_  | ~\new_[5854]_ ;
  assign \new_[5708]_  = ~\new_[5867]_  | ~\new_[5868]_ ;
  assign \new_[5709]_  = ~\new_[5870]_  | ~\new_[5871]_ ;
  assign \new_[5710]_  = ~\new_[20545]_ ;
  assign \new_[5711]_  = ~output_backup_par_en_out_reg;
  assign \new_[5712]_  = \new_[5891]_  ? \new_[20413]_  : \new_[18600]_ ;
  assign \new_[5713]_  = \new_[5889]_  ? \new_[20413]_  : \new_[17855]_ ;
  assign \new_[5714]_  = \new_[5890]_  ? \new_[20413]_  : \new_[18884]_ ;
  assign \new_[5715]_  = \new_[5892]_  ? \new_[20413]_  : \new_[17882]_ ;
  assign \new_[5716]_  = \new_[5894]_  ? \new_[20413]_  : \new_[18848]_ ;
  assign \new_[5717]_  = \new_[5895]_  ? \new_[20413]_  : \new_[19639]_ ;
  assign \new_[5718]_  = \new_[5898]_  ? \new_[20413]_  : \new_[19844]_ ;
  assign \new_[5719]_  = \new_[5896]_  ? \new_[20413]_  : \new_[18080]_ ;
  assign \new_[5720]_  = \new_[5897]_  ? \new_[20413]_  : \new_[18521]_ ;
  assign \new_[5721]_  = \new_[5899]_  ? \new_[20413]_  : \new_[18386]_ ;
  assign \new_[5722]_  = \new_[5900]_  ? \new_[20413]_  : \new_[18105]_ ;
  assign \new_[5723]_  = \new_[5901]_  ? \new_[20413]_  : \new_[18480]_ ;
  assign \new_[5724]_  = \new_[5902]_  ? \new_[20413]_  : \new_[18239]_ ;
  assign \new_[5725]_  = \new_[5903]_  ? \new_[20413]_  : \new_[18037]_ ;
  assign \new_[5726]_  = \new_[5904]_  ? \new_[20413]_  : \new_[19849]_ ;
  assign \new_[5727]_  = \new_[5905]_  ? \new_[20413]_  : \new_[18992]_ ;
  assign \new_[5728]_  = \new_[5906]_  ? \new_[20413]_  : \new_[19721]_ ;
  assign \new_[5729]_  = \new_[5907]_  ? \new_[20413]_  : \new_[19042]_ ;
  assign \new_[5730]_  = \new_[5908]_  ? \new_[20413]_  : \new_[19009]_ ;
  assign \new_[5731]_  = \new_[5909]_  ? \new_[20413]_  : \new_[18948]_ ;
  assign \new_[5732]_  = \new_[5910]_  ? \new_[20413]_  : \new_[18936]_ ;
  assign \new_[5733]_  = \new_[5911]_  ? \new_[20413]_  : \new_[19593]_ ;
  assign \new_[5734]_  = \new_[5913]_  ? \new_[20413]_  : \new_[18607]_ ;
  assign \new_[5735]_  = \new_[5914]_  ? \new_[20413]_  : \new_[17825]_ ;
  assign \new_[5736]_  = \new_[5915]_  ? \new_[20413]_  : \new_[19321]_ ;
  assign \new_[5737]_  = \new_[5916]_  ? \new_[20413]_  : \new_[18603]_ ;
  assign \new_[5738]_  = \new_[5917]_  ? \new_[20413]_  : \new_[19044]_ ;
  assign \new_[5739]_  = \new_[5918]_  ? \new_[20413]_  : \new_[19735]_ ;
  assign n2645 = \new_[18607]_  ? \new_[10827]_  : \new_[5913]_ ;
  assign n2650 = \new_[17825]_  ? \new_[10827]_  : \new_[5914]_ ;
  assign n2655 = \new_[19321]_  ? \new_[10827]_  : \new_[5915]_ ;
  assign n2775 = \new_[18603]_  ? \new_[10827]_  : \new_[5916]_ ;
  assign n2660 = \new_[19044]_  ? \new_[10827]_  : \new_[5917]_ ;
  assign n2665 = \new_[19735]_  ? \new_[10827]_  : \new_[5918]_ ;
  assign n2785 = \new_[18600]_  ? \new_[10827]_  : \new_[5891]_ ;
  assign n2670 = \new_[17855]_  ? \new_[10827]_  : \new_[5889]_ ;
  assign \new_[5748]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15] ;
  assign \new_[5749]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16] ;
  assign \new_[5750]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17] ;
  assign \new_[5751]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18] ;
  assign \new_[5752]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19] ;
  assign \new_[5753]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1] ;
  assign \new_[5754]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20] ;
  assign \new_[5755]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22] ;
  assign \new_[5756]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23] ;
  assign \new_[5757]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24] ;
  assign \new_[5758]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27] ;
  assign \new_[5759]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28] ;
  assign \new_[5760]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29] ;
  assign \new_[5761]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2] ;
  assign \new_[5762]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31] ;
  assign \new_[5763]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3] ;
  assign \new_[5764]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4] ;
  assign \new_[5765]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5] ;
  assign \new_[5766]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6] ;
  assign \new_[5767]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7] ;
  assign \new_[5768]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8] ;
  assign \new_[5769]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9] ;
  assign \new_[5770]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32] ;
  assign \new_[5771]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34] ;
  assign \new_[5772]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35] ;
  assign \new_[5773]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0] ;
  assign \new_[5774]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10] ;
  assign \new_[5775]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11] ;
  assign \new_[5776]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12] ;
  assign \new_[5777]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13] ;
  assign \new_[5778]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14] ;
  assign \new_[5779]_  = \new_[20415]_  & \new_[5912]_ ;
  assign \new_[5780]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33] ;
  assign \new_[5781]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36] ;
  assign \new_[5782]_  = ~\new_[5950]_  & ~\new_[6001]_ ;
  assign \new_[5783]_  = ~\new_[5951]_  & ~\new_[5962]_ ;
  assign \new_[5784]_  = ~\new_[5952]_  & ~\new_[6024]_ ;
  assign \new_[5785]_  = ~\new_[5954]_  | ~\new_[6066]_ ;
  assign \new_[5786]_  = ~\new_[5956]_  & ~\new_[6082]_ ;
  assign \new_[5787]_  = \new_[5957]_  & \new_[6096]_ ;
  assign \new_[5788]_  = ~\new_[5958]_  & ~\new_[5975]_ ;
  assign \new_[5789]_  = ~\new_[5959]_  & ~\new_[5979]_ ;
  assign \new_[5790]_  = ~\new_[5801]_ ;
  assign pci_par_oe_o = pci_io_mux_par_iob_en_out_reg;
  assign \new_[5792]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21] ;
  assign \new_[5793]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25] ;
  assign \new_[5794]_  = \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30] ;
  assign n2795 = ~n2965;
  assign \new_[5796]_  = ~\new_[5893]_ ;
  assign \new_[5797]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[25] ;
  assign \new_[5798]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[15] ;
  assign \new_[5799]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[7] ;
  assign n2790 = ~\new_[8638]_  | ~\new_[8331]_  | ~\new_[5993]_  | ~\new_[8332]_ ;
  assign \new_[5801]_  = ~n3000 | ~\new_[11137]_  | ~n9630;
  assign \new_[5802]_  = ~\new_[5997]_  & ~\new_[5998]_ ;
  assign \new_[5803]_  = ~\new_[5999]_  & ~\new_[6000]_ ;
  assign \new_[5804]_  = ~\new_[6002]_  & ~\new_[6003]_ ;
  assign \new_[5805]_  = ~\new_[6004]_  & ~\new_[6005]_ ;
  assign \new_[5806]_  = ~\new_[6007]_  & ~\new_[6008]_ ;
  assign \new_[5807]_  = ~\new_[6014]_  & ~\new_[6015]_ ;
  assign \new_[5808]_  = ~\new_[6016]_  & ~\new_[6017]_ ;
  assign \new_[5809]_  = ~\new_[6018]_  & ~\new_[6019]_ ;
  assign \new_[5810]_  = ~\new_[6020]_  & ~\new_[6021]_ ;
  assign \new_[5811]_  = ~\new_[6022]_  & ~\new_[6023]_ ;
  assign \new_[5812]_  = ~\new_[6026]_  & ~\new_[6025]_ ;
  assign \new_[5813]_  = ~\new_[6229]_  & ~\new_[6027]_ ;
  assign \new_[5814]_  = ~\new_[6028]_  & ~\new_[6230]_ ;
  assign \new_[5815]_  = ~\new_[6030]_  & ~\new_[6031]_ ;
  assign \new_[5816]_  = ~\new_[6032]_  & ~\new_[6231]_ ;
  assign \new_[5817]_  = ~\new_[6033]_  & ~\new_[6232]_ ;
  assign \new_[5818]_  = ~\new_[6233]_  & ~\new_[6035]_ ;
  assign \new_[5819]_  = ~\new_[6036]_  & ~\new_[6037]_ ;
  assign \new_[5820]_  = ~\new_[6038]_  & ~\new_[6234]_ ;
  assign \new_[5821]_  = ~\new_[6040]_  & ~\new_[6041]_ ;
  assign \new_[5822]_  = ~\new_[6042]_  & ~\new_[6235]_ ;
  assign \new_[5823]_  = ~\new_[6236]_  & ~\new_[6044]_ ;
  assign \new_[5824]_  = ~\new_[6047]_  & ~\new_[6238]_ ;
  assign \new_[5825]_  = ~\new_[6239]_  & ~\new_[6049]_ ;
  assign \new_[5826]_  = ~\new_[6050]_  & ~\new_[6051]_ ;
  assign \new_[5827]_  = ~\new_[6240]_  & ~\new_[6052]_ ;
  assign \new_[5828]_  = ~\new_[7019]_  | ~\new_[6372]_  | ~\new_[6463]_  | ~\new_[7127]_ ;
  assign \new_[5829]_  = ~\new_[6055]_  & ~\new_[6241]_ ;
  assign \new_[5830]_  = ~\new_[6057]_  & ~\new_[6058]_ ;
  assign \new_[5831]_  = ~\new_[6059]_  & ~\new_[6060]_ ;
  assign \new_[5832]_  = ~\new_[6242]_  & ~\new_[6061]_ ;
  assign \new_[5833]_  = ~\new_[6243]_  & ~\new_[6063]_ ;
  assign \new_[5834]_  = ~\new_[6064]_  & ~\new_[6244]_ ;
  assign \new_[5835]_  = ~\new_[6247]_  & ~\new_[6067]_ ;
  assign \new_[5836]_  = ~\new_[6068]_  & ~\new_[6069]_ ;
  assign \new_[5837]_  = ~\new_[6248]_  & ~\new_[6070]_ ;
  assign \new_[5838]_  = ~\new_[6075]_  & ~\new_[6076]_ ;
  assign \new_[5839]_  = ~\new_[6250]_  & ~\new_[6078]_ ;
  assign \new_[5840]_  = ~\new_[6079]_  & ~\new_[6251]_ ;
  assign \new_[5841]_  = ~\new_[6252]_  & ~\new_[6080]_ ;
  assign \new_[5842]_  = ~\new_[7023]_  | ~\new_[6382]_  | ~\new_[7152]_  | ~\new_[7153]_ ;
  assign \new_[5843]_  = ~\new_[6255]_  & ~\new_[6083]_ ;
  assign \new_[5844]_  = ~\new_[6084]_  & ~\new_[6085]_ ;
  assign \new_[5845]_  = ~\new_[7024]_  | ~\new_[6388]_  | ~\new_[6490]_  | ~\new_[6491]_ ;
  assign \new_[5846]_  = ~\new_[6087]_  & ~\new_[6088]_ ;
  assign \new_[5847]_  = ~\new_[6089]_  & ~\new_[6090]_ ;
  assign \new_[5848]_  = ~\new_[7025]_  | ~\new_[6391]_  | ~\new_[6495]_  | ~\new_[6496]_ ;
  assign \new_[5849]_  = ~\new_[6092]_  & ~\new_[6093]_ ;
  assign \new_[5850]_  = ~\new_[6094]_  & ~\new_[6095]_ ;
  assign \new_[5851]_  = ~\new_[6097]_  & ~\new_[6098]_ ;
  assign \new_[5852]_  = ~\new_[6099]_  & ~\new_[6100]_ ;
  assign \new_[5853]_  = ~\new_[6102]_  & ~\new_[6103]_ ;
  assign \new_[5854]_  = ~\new_[6104]_  & ~\new_[6105]_ ;
  assign \new_[5855]_  = ~\new_[6106]_  & ~\new_[6259]_ ;
  assign \new_[5856]_  = ~\new_[6261]_  & ~\new_[6107]_ ;
  assign \new_[5857]_  = ~\new_[6108]_  & ~\new_[6109]_ ;
  assign \new_[5858]_  = ~\new_[6110]_  & ~\new_[6262]_ ;
  assign \new_[5859]_  = ~\new_[6263]_  & ~\new_[6112]_ ;
  assign \new_[5860]_  = ~\new_[6113]_  & ~\new_[6114]_ ;
  assign \new_[5861]_  = ~\new_[6115]_  & ~\new_[6264]_ ;
  assign \new_[5862]_  = ~\new_[6117]_  & ~\new_[6118]_ ;
  assign \new_[5863]_  = ~\new_[6119]_  & ~\new_[6120]_ ;
  assign \new_[5864]_  = ~\new_[6121]_  & ~\new_[6265]_ ;
  assign \new_[5865]_  = ~\new_[6266]_  & ~\new_[6123]_ ;
  assign \new_[5866]_  = ~\new_[6124]_  & ~\new_[6125]_ ;
  assign \new_[5867]_  = ~\new_[6127]_  & ~\new_[6128]_ ;
  assign \new_[5868]_  = ~\new_[6129]_  & ~\new_[6130]_ ;
  assign \new_[5869]_  = ~\new_[6406]_  | ~\new_[7340]_  | ~\new_[6526]_  | ~\new_[7205]_ ;
  assign \new_[5870]_  = ~\new_[6132]_  & ~\new_[6133]_ ;
  assign \new_[5871]_  = ~\new_[6134]_  & ~\new_[6267]_ ;
  assign \new_[5872]_  = ~\new_[6410]_  | ~\new_[7341]_  | ~\new_[6529]_  | ~\new_[7210]_ ;
  assign \new_[5873]_  = ~\new_[6268]_  & ~\new_[6136]_ ;
  assign \new_[5874]_  = ~\new_[6269]_  & ~\new_[6137]_ ;
  assign \new_[5875]_  = ~\new_[6270]_  & ~\new_[6138]_ ;
  assign \new_[5876]_  = ~\new_[6140]_  & ~\new_[6141]_ ;
  assign \new_[5877]_  = ~\new_[6142]_  & ~\new_[6143]_ ;
  assign \new_[5878]_  = ~\new_[7028]_  | ~\new_[6414]_  | ~\new_[6537]_  | ~\new_[6536]_ ;
  assign \new_[5879]_  = ~\new_[6145]_  & ~\new_[6146]_ ;
  assign \new_[5880]_  = ~\new_[6147]_  & ~\new_[6148]_ ;
  assign \new_[5881]_  = ~\new_[6150]_  & ~\new_[6149]_ ;
  assign \new_[5882]_  = ~\new_[6151]_  & ~\new_[6152]_ ;
  assign \new_[5883]_  = ~\new_[6153]_  & ~\new_[6154]_ ;
  assign \new_[5884]_  = ~\new_[6272]_  & ~\new_[6155]_ ;
  assign \new_[5885]_  = ~\new_[6161]_  & ~\new_[6273]_ ;
  assign \new_[5886]_  = ~\new_[20199]_ ;
  assign \new_[5887]_  = ~\new_[13807]_  & ~\new_[6165]_ ;
  assign \new_[5888]_  = \\pci_target_unit_wishbone_master_c_state_reg[0] ;
  assign \new_[5889]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[17] ;
  assign \new_[5890]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[18] ;
  assign \new_[5891]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[16] ;
  assign \new_[5892]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[19] ;
  assign \new_[5893]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[1] ;
  assign \new_[5894]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[20] ;
  assign \new_[5895]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[21] ;
  assign \new_[5896]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[23] ;
  assign \new_[5897]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[24] ;
  assign \new_[5898]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[22] ;
  assign \new_[5899]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[26] ;
  assign \new_[5900]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[27] ;
  assign \new_[5901]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[28] ;
  assign \new_[5902]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[29] ;
  assign \new_[5903]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[2] ;
  assign \new_[5904]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[30] ;
  assign \new_[5905]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[31] ;
  assign \new_[5906]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[3] ;
  assign \new_[5907]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[4] ;
  assign \new_[5908]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[5] ;
  assign \new_[5909]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[6] ;
  assign \new_[5910]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[8] ;
  assign \new_[5911]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[9] ;
  assign \new_[5912]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[37] ;
  assign \new_[5913]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[0] ;
  assign \new_[5914]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[10] ;
  assign \new_[5915]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[11] ;
  assign \new_[5916]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[12] ;
  assign \new_[5917]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[13] ;
  assign \new_[5918]_  = \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[14] ;
  assign n2925 = ~\new_[8293]_  | ~\new_[8294]_  | ~\new_[6167]_  | ~\new_[8116]_ ;
  assign n2930 = ~\new_[8295]_  | ~\new_[8577]_  | ~\new_[6168]_  | ~\new_[8119]_ ;
  assign n2935 = ~\new_[8580]_  | ~\new_[8581]_  | ~\new_[6169]_  | ~\new_[8123]_ ;
  assign n2940 = ~\new_[8586]_  | ~\new_[8587]_  | ~\new_[6170]_  | ~\new_[8125]_ ;
  assign n2945 = ~\new_[8298]_  | ~\new_[8299]_  | ~\new_[6171]_  | ~\new_[8127]_ ;
  assign n2950 = ~\new_[8595]_  | ~\new_[8301]_  | ~\new_[6172]_  | ~\new_[8129]_ ;
  assign n2800 = ~\new_[8303]_  | ~\new_[8304]_  | ~\new_[6173]_  | ~\new_[8305]_ ;
  assign n2805 = ~\new_[8307]_  | ~\new_[8604]_  | ~\new_[6174]_  | ~\new_[8132]_ ;
  assign n2810 = ~\new_[8134]_  | ~\new_[8609]_  | ~\new_[6175]_  | ~\new_[8309]_ ;
  assign n2820 = ~\new_[8615]_  | ~\new_[8312]_  | ~\new_[6176]_  | ~\new_[8313]_ ;
  assign n2825 = ~\new_[8315]_  | ~\new_[8316]_  | ~\new_[6177]_  | ~\new_[8138]_ ;
  assign n2830 = ~\new_[8141]_  | ~\new_[8318]_  | ~\new_[6178]_  | ~\new_[8319]_ ;
  assign n2835 = ~\new_[8322]_  | ~\new_[8323]_  | ~\new_[6179]_  | ~\new_[8324]_ ;
  assign n2840 = ~\new_[8631]_  | ~\new_[8325]_  | ~\new_[6180]_  | ~\new_[8326]_ ;
  assign n2850 = ~\new_[8335]_  | ~\new_[8334]_  | ~\new_[6181]_  | ~\new_[8336]_ ;
  assign n2855 = ~\new_[8339]_  | ~\new_[8643]_  | ~\new_[6182]_  | ~\new_[8340]_ ;
  assign n2860 = ~\new_[8161]_  | ~\new_[8342]_  | ~\new_[6183]_  | ~\new_[8343]_ ;
  assign n2865 = ~\new_[8649]_  | ~\new_[8650]_  | ~\new_[6184]_  | ~\new_[8163]_ ;
  assign n2870 = ~\new_[7410]_  | ~\new_[8349]_  | ~\new_[6185]_  | ~\new_[8167]_ ;
  assign n2910 = ~\new_[8169]_  | ~\new_[7412]_  | ~\new_[6186]_  | ~\new_[8170]_ ;
  assign n2955 = ~\new_[7413]_  | ~\new_[8172]_  | ~\new_[6187]_  | ~\new_[8173]_ ;
  assign n2915 = ~\new_[8175]_  | ~\new_[8176]_  | ~\new_[6188]_  | ~\new_[7416]_ ;
  assign n2920 = ~\new_[8359]_  | ~\new_[7418]_  | ~\new_[6189]_  | ~\new_[8178]_ ;
  assign n2960 = ~\new_[8179]_  | ~\new_[8362]_  | ~\new_[6190]_  | ~\new_[8180]_ ;
  assign n2875 = ~\new_[7422]_  | ~\new_[8365]_  | ~\new_[6191]_  | ~\new_[8182]_ ;
  assign n2880 = ~\new_[7423]_  | ~\new_[8184]_  | ~\new_[6192]_  | ~\new_[8185]_ ;
  assign n2885 = ~\new_[8188]_  | ~\new_[8189]_  | ~\new_[6193]_  | ~\new_[8190]_ ;
  assign n2890 = ~\new_[8192]_  | ~\new_[7425]_  | ~\new_[6194]_  | ~\new_[8193]_ ;
  assign n2895 = ~\new_[8376]_  | ~\new_[8377]_  | ~\new_[6195]_  | ~\new_[7427]_ ;
  assign n2900 = ~\new_[8381]_  | ~\new_[8196]_  | ~\new_[6196]_  | ~\new_[7428]_ ;
  assign n2905 = ~\new_[7429]_  | ~\new_[8198]_  | ~\new_[6197]_  | ~\new_[8199]_ ;
  assign \new_[5950]_  = ~\new_[7079]_  | ~\new_[7080]_  | ~\new_[7077]_  | ~\new_[7078]_ ;
  assign \new_[5951]_  = ~\new_[7092]_  | ~\new_[7093]_  | ~\new_[6439]_  | ~\new_[7091]_ ;
  assign \new_[5952]_  = ~\new_[7098]_  | ~\new_[7099]_  | ~\new_[7097]_  | ~\new_[7096]_ ;
  assign \new_[5953]_  = ~\new_[7128]_  | ~\new_[7129]_  | ~\new_[6465]_  | ~\new_[6464]_ ;
  assign \new_[5954]_  = ~\new_[6245]_  & ~\new_[6246]_ ;
  assign \new_[5955]_  = ~\new_[7154]_  | ~\new_[7327]_  | ~\new_[6487]_  | ~\new_[6488]_ ;
  assign \new_[5956]_  = ~\new_[7158]_  | ~\new_[7157]_  | ~\new_[6383]_  | ~\new_[7328]_ ;
  assign \new_[5957]_  = ~\new_[6256]_  & ~\new_[6257]_ ;
  assign \new_[5958]_  = ~\new_[7057]_  | ~\new_[7332]_  | ~\new_[7175]_  | ~\new_[7176]_ ;
  assign \new_[5959]_  = ~\new_[7200]_  | ~\new_[7201]_  | ~\new_[7198]_  | ~\new_[7199]_ ;
  assign \new_[5960]_  = ~\new_[6275]_  & (~\new_[8103]_  | ~\new_[18294]_ );
  assign \new_[5961]_  = ~\new_[6282]_  | ~\new_[7309]_ ;
  assign \new_[5962]_  = ~\new_[6283]_  | ~\new_[6356]_ ;
  assign \new_[5963]_  = ~\new_[6276]_  & (~\new_[8103]_  | ~\new_[19314]_ );
  assign \new_[5964]_  = ~\new_[6284]_  | ~\new_[6359]_ ;
  assign \new_[5965]_  = ~\new_[6285]_  | ~\new_[6361]_ ;
  assign \new_[5966]_  = ~\new_[6277]_  & (~\new_[8103]_  | ~\new_[19481]_ );
  assign \new_[5967]_  = ~\new_[6291]_  & (~\new_[8284]_  | ~\new_[18211]_ );
  assign \new_[5968]_  = ~\new_[6054]_ ;
  assign \new_[5969]_  = ~\new_[6292]_  & (~\new_[7386]_  | ~\new_[19703]_ );
  assign \new_[5970]_  = ~\new_[6293]_  & (~\new_[8284]_  | ~\new_[19050]_ );
  assign \new_[5971]_  = ~\new_[6278]_  & (~\new_[8103]_  | ~\new_[19196]_ );
  assign \new_[5972]_  = ~\new_[6294]_  & (~\new_[8284]_  | ~\new_[19462]_ );
  assign \new_[5973]_  = ~\new_[6295]_  & (~\new_[8284]_  | ~\new_[19856]_ );
  assign \new_[5974]_  = ~\new_[6296]_  & (~\new_[8284]_  | ~\new_[19620]_ );
  assign \new_[5975]_  = ~\new_[6287]_  | ~\new_[6395]_ ;
  assign \new_[5976]_  = ~\new_[6279]_  & (~\new_[7387]_  | ~\new_[19483]_ );
  assign \new_[5977]_  = ~\new_[6297]_  & (~\new_[7386]_  | ~\new_[17898]_ );
  assign \new_[5978]_  = ~\new_[6298]_  & (~\new_[8284]_  | ~\new_[18352]_ );
  assign \new_[5979]_  = ~\new_[6280]_  | ~\new_[6404]_ ;
  assign \new_[5980]_  = ~\new_[6288]_  | ~\new_[6407]_ ;
  assign \new_[5981]_  = ~\new_[6289]_  | ~\new_[6409]_ ;
  assign \new_[5982]_  = ~\new_[6299]_  & (~\new_[7386]_  | ~\new_[18267]_ );
  assign \new_[5983]_  = ~\new_[6300]_  & (~\new_[8284]_  | ~\new_[18095]_ );
  assign \new_[5984]_  = ~\new_[6301]_  & (~\new_[7386]_  | ~\new_[18266]_ );
  assign \new_[5985]_  = ~\new_[6302]_  & (~\new_[8284]_  | ~\new_[19827]_ );
  assign \new_[5986]_  = \new_[6166]_  & \new_[16658]_ ;
  assign n2965 = ~\new_[6165]_  & ~\new_[6917]_ ;
  assign \new_[5988]_  = ~\new_[6166]_ ;
  assign \new_[5989]_  = ~\new_[6166]_ ;
  assign n2970 = ~\new_[8626]_  | ~\new_[8320]_  | ~\new_[6331]_  | ~\new_[8628]_ ;
  assign n2975 = ~\new_[8329]_  | ~\new_[8153]_  | ~\new_[6332]_  | ~\new_[8330]_ ;
  assign n2980 = ~\new_[8346]_  | ~\new_[8653]_  | ~\new_[6333]_  | ~\new_[8165]_ ;
  assign \new_[5993]_  = ~\new_[6334]_  & ~\new_[7408]_ ;
  assign n2990 = ~\new_[7991]_  | ~\new_[7353]_  | ~\new_[8264]_  | ~\new_[7352]_ ;
  assign n2985 = ~\new_[7356]_  | ~\new_[8029]_  | ~\new_[8269]_  | ~\new_[8028]_ ;
  assign n2995 = ~\new_[8070]_  | ~\new_[7366]_  | ~\new_[8273]_  | ~\new_[8069]_ ;
  assign \new_[5997]_  = ~\new_[6421]_  | ~\new_[7075]_ ;
  assign \new_[5998]_  = ~\new_[6350]_  | ~\new_[7306]_ ;
  assign \new_[5999]_  = ~\new_[6351]_  | ~\new_[7030]_ ;
  assign \new_[6000]_  = ~\new_[7076]_  | ~\new_[6422]_ ;
  assign \new_[6001]_  = ~\new_[7081]_  | ~\new_[6423]_ ;
  assign \new_[6002]_  = ~\new_[7082]_  | ~\new_[6424]_ ;
  assign \new_[6003]_  = ~\new_[6425]_  | ~\new_[7083]_ ;
  assign \new_[6004]_  = ~\new_[6426]_  | ~\new_[6427]_ ;
  assign \new_[6005]_  = ~\new_[6335]_  | ~\new_[7031]_ ;
  assign \new_[6006]_  = ~\new_[6428]_  | ~\new_[6429]_ ;
  assign \new_[6007]_  = ~\new_[6352]_  | ~\new_[7032]_ ;
  assign \new_[6008]_  = ~\new_[6430]_  | ~\new_[7084]_ ;
  assign \new_[6009]_  = ~\new_[6353]_  & (~\new_[8279]_  | ~\new_[18688]_ );
  assign \new_[6010]_  = ~\new_[6336]_  | ~\new_[6354]_ ;
  assign \new_[6011]_  = ~\new_[7085]_  | ~\new_[6431]_ ;
  assign \new_[6012]_  = ~\new_[6432]_  | ~\new_[7307]_ ;
  assign \new_[6013]_  = ~\new_[6433]_  | ~\new_[6434]_ ;
  assign \new_[6014]_  = ~\new_[6355]_  | ~\new_[7033]_ ;
  assign \new_[6015]_  = ~\new_[6435]_  | ~\new_[7086]_ ;
  assign \new_[6016]_  = ~\new_[6436]_  | ~\new_[7088]_ ;
  assign \new_[6017]_  = ~\new_[6437]_  | ~\new_[7089]_ ;
  assign \new_[6018]_  = ~\new_[7090]_  | ~\new_[6438]_ ;
  assign \new_[6019]_  = ~\new_[6337]_  | ~\new_[7034]_ ;
  assign \new_[6020]_  = ~\new_[6357]_  | ~\new_[7035]_ ;
  assign \new_[6021]_  = ~\new_[7094]_  | ~\new_[6440]_ ;
  assign \new_[6022]_  = ~\new_[6441]_  | ~\new_[7095]_ ;
  assign \new_[6023]_  = ~\new_[6358]_  | ~\new_[7310]_ ;
  assign \new_[6024]_  = ~\new_[7100]_  | ~\new_[6442]_ ;
  assign \new_[6025]_  = ~\new_[6443]_  | ~\new_[7311]_ ;
  assign \new_[6026]_  = ~\new_[7101]_  | ~\new_[6444]_ ;
  assign \new_[6027]_  = ~\new_[6338]_  | ~\new_[7036]_ ;
  assign \new_[6028]_  = ~\new_[7104]_  | ~\new_[6445]_ ;
  assign \new_[6029]_  = ~\new_[6446]_  & (~\new_[8094]_  | ~\new_[17902]_ );
  assign \new_[6030]_  = ~\new_[6447]_  | ~\new_[7105]_ ;
  assign \new_[6031]_  = ~\new_[7106]_  | ~\new_[6448]_ ;
  assign \new_[6032]_  = ~\new_[6339]_  | ~\new_[6360]_ ;
  assign \new_[6033]_  = ~\new_[7109]_  | ~\new_[6449]_ ;
  assign \new_[6034]_  = ~\new_[6450]_  & (~\new_[8094]_  | ~\new_[17899]_ );
  assign \new_[6035]_  = ~\new_[6362]_  | ~\new_[7039]_ ;
  assign \new_[6036]_  = ~\new_[6363]_  | ~\new_[7314]_ ;
  assign \new_[6037]_  = ~\new_[7112]_  | ~\new_[6451]_ ;
  assign \new_[6038]_  = ~\new_[6452]_  | ~\new_[7315]_ ;
  assign \new_[6039]_  = ~\new_[6453]_  & (~\new_[7386]_  | ~\new_[19275]_ );
  assign \new_[6040]_  = ~\new_[6365]_  | ~\new_[7040]_ ;
  assign \new_[6041]_  = ~\new_[6364]_  | ~\new_[7316]_ ;
  assign \new_[6042]_  = ~\new_[6454]_  | ~\new_[7115]_ ;
  assign \new_[6043]_  = ~\new_[6455]_  & (~\new_[8084]_  | ~\new_[19104]_ );
  assign \new_[6044]_  = ~\new_[6457]_  | ~\new_[6456]_ ;
  assign \new_[6045]_  = ~\new_[6367]_  | ~\new_[7042]_ ;
  assign \new_[6046]_  = ~\new_[6459]_  | ~\new_[7120]_ ;
  assign \new_[6047]_  = ~\new_[7018]_  | ~\new_[6368]_ ;
  assign \new_[6048]_  = ~\new_[6460]_  & (~\new_[8556]_  | ~\new_[18486]_ );
  assign \new_[6049]_  = ~\new_[6369]_  | ~\new_[7319]_ ;
  assign \new_[6050]_  = ~\new_[7124]_  | ~\new_[6461]_ ;
  assign \new_[6051]_  = ~\new_[6370]_  | ~\new_[7043]_ ;
  assign \new_[6052]_  = ~\new_[6340]_  | ~\new_[6371]_ ;
  assign \new_[6053]_  = ~\new_[6462]_  & (~\new_[7386]_  | ~\new_[19535]_ );
  assign \new_[6054]_  = ~\new_[6466]_  | ~\new_[6467]_ ;
  assign \new_[6055]_  = ~\new_[6373]_  | ~\new_[7044]_ ;
  assign \new_[6056]_  = ~\new_[6468]_  & (~\new_[8094]_  | ~\new_[19323]_ );
  assign \new_[6057]_  = ~\new_[7130]_  | ~\new_[6469]_ ;
  assign \new_[6058]_  = ~\new_[6374]_  | ~\new_[7321]_ ;
  assign \new_[6059]_  = ~\new_[6375]_  | ~\new_[7046]_ ;
  assign \new_[6060]_  = ~\new_[6470]_  | ~\new_[7131]_ ;
  assign \new_[6061]_  = ~\new_[6471]_  | ~\new_[7322]_ ;
  assign \new_[6062]_  = ~\new_[6341]_  & (~\new_[7387]_  | ~\new_[17846]_ );
  assign \new_[6063]_  = ~\new_[6376]_  | ~\new_[7048]_ ;
  assign \new_[6064]_  = ~\new_[6472]_  | ~\new_[7134]_ ;
  assign \new_[6065]_  = ~\new_[6473]_  & (~\new_[8084]_  | ~\new_[18127]_ );
  assign \new_[6066]_  = ~\new_[6474]_  & (~\new_[7386]_  | ~\new_[18942]_ );
  assign \new_[6067]_  = ~\new_[7138]_  | ~\new_[6475]_ ;
  assign \new_[6068]_  = ~\new_[6476]_  | ~\new_[7139]_ ;
  assign \new_[6069]_  = ~\new_[6377]_  | ~\new_[7051]_ ;
  assign \new_[6070]_  = ~\new_[6477]_  | ~\new_[6478]_ ;
  assign \new_[6071]_  = ~\new_[6479]_  & (~\new_[8082]_  | ~\new_[18318]_ );
  assign \new_[6072]_  = ~\new_[7140]_  | ~\new_[6480]_ ;
  assign \new_[6073]_  = ~\new_[6481]_  | ~\new_[6482]_ ;
  assign \new_[6074]_  = ~\new_[7022]_  | ~\new_[6378]_ ;
  assign \new_[6075]_  = ~\new_[7143]_  | ~\new_[6483]_ ;
  assign \new_[6076]_  = ~\new_[6484]_  | ~\new_[7144]_ ;
  assign \new_[6077]_  = ~\new_[6380]_  & (~\new_[8279]_  | ~\new_[18582]_ );
  assign \new_[6078]_  = ~\new_[6485]_  | ~\new_[7145]_ ;
  assign \new_[6079]_  = ~\new_[6381]_  | ~\new_[7054]_ ;
  assign \new_[6080]_  = ~\new_[6486]_  | ~\new_[7150]_ ;
  assign \new_[6081]_  = ~\new_[6254]_ ;
  assign \new_[6082]_  = ~\new_[6384]_  | ~\new_[6385]_ ;
  assign \new_[6083]_  = ~\new_[7161]_  | ~\new_[6489]_ ;
  assign \new_[6084]_  = ~\new_[6386]_  | ~\new_[20333]_ ;
  assign \new_[6085]_  = ~\new_[6387]_  | ~\new_[7329]_ ;
  assign \new_[6086]_  = ~\new_[7162]_  | ~\new_[6492]_ ;
  assign \new_[6087]_  = ~\new_[6493]_  | ~\new_[7163]_ ;
  assign \new_[6088]_  = ~\new_[6389]_  | ~\new_[7055]_ ;
  assign \new_[6089]_  = ~\new_[7164]_  | ~\new_[6494]_ ;
  assign \new_[6090]_  = ~\new_[6390]_  | ~\new_[7330]_ ;
  assign \new_[6091]_  = ~\new_[7165]_  | ~\new_[6497]_ ;
  assign \new_[6092]_  = ~\new_[7166]_  | ~\new_[6498]_ ;
  assign \new_[6093]_  = ~\new_[6392]_  | ~\new_[7331]_ ;
  assign \new_[6094]_  = ~\new_[6393]_  | ~\new_[7056]_ ;
  assign \new_[6095]_  = ~\new_[6499]_  | ~\new_[7167]_ ;
  assign \new_[6096]_  = ~\new_[6342]_  & (~\new_[7387]_  | ~\new_[17837]_ );
  assign \new_[6097]_  = ~\new_[6343]_  | ~\new_[6394]_ ;
  assign \new_[6098]_  = ~\new_[6500]_  | ~\new_[7172]_ ;
  assign \new_[6099]_  = ~\new_[7173]_  | ~\new_[6501]_ ;
  assign \new_[6100]_  = ~\new_[6502]_  | ~\new_[7174]_ ;
  assign \new_[6101]_  = ~\new_[6504]_  | ~\new_[6503]_ ;
  assign \new_[6102]_  = ~\new_[6505]_  | ~\new_[7177]_ ;
  assign \new_[6103]_  = ~\new_[6506]_  | ~\new_[7178]_ ;
  assign \new_[6104]_  = ~\new_[6344]_  | ~\new_[6396]_ ;
  assign \new_[6105]_  = ~\new_[7179]_  | ~\new_[6507]_ ;
  assign \new_[6106]_  = ~\new_[7182]_  | ~\new_[6508]_ ;
  assign \new_[6107]_  = ~\new_[6509]_  | ~\new_[7183]_ ;
  assign \new_[6108]_  = ~\new_[6397]_  | ~\new_[7061]_ ;
  assign \new_[6109]_  = ~\new_[7184]_  | ~\new_[6510]_ ;
  assign \new_[6110]_  = ~\new_[6511]_  | ~\new_[7335]_ ;
  assign \new_[6111]_  = ~\new_[6512]_  & (~\new_[7386]_  | ~\new_[18716]_ );
  assign \new_[6112]_  = ~\new_[7189]_  | ~\new_[6513]_ ;
  assign \new_[6113]_  = ~\new_[6398]_  | ~\new_[7336]_ ;
  assign \new_[6114]_  = ~\new_[6399]_  | ~\new_[7062]_ ;
  assign \new_[6115]_  = ~\new_[6514]_  | ~\new_[7337]_ ;
  assign \new_[6116]_  = ~\new_[6345]_  & (~\new_[7387]_  | ~\new_[18039]_ );
  assign \new_[6117]_  = ~\new_[6400]_  | ~\new_[7063]_ ;
  assign \new_[6118]_  = ~\new_[7192]_  | ~\new_[6515]_ ;
  assign \new_[6119]_  = ~\new_[6516]_  | ~\new_[7193]_ ;
  assign \new_[6120]_  = ~\new_[6401]_  | ~\new_[7338]_ ;
  assign \new_[6121]_  = ~\new_[7026]_  | ~\new_[6402]_ ;
  assign \new_[6122]_  = ~\new_[6517]_  & (~\new_[7386]_  | ~\new_[18368]_ );
  assign \new_[6123]_  = ~\new_[6403]_  | ~\new_[7065]_ ;
  assign \new_[6124]_  = ~\new_[6518]_  | ~\new_[7196]_ ;
  assign \new_[6125]_  = ~\new_[7197]_  | ~\new_[6519]_ ;
  assign \new_[6126]_  = ~\new_[6520]_  & (~\new_[8084]_  | ~\new_[18767]_ );
  assign \new_[6127]_  = ~\new_[6521]_  | ~\new_[7202]_ ;
  assign \new_[6128]_  = ~\new_[6522]_  | ~\new_[7203]_ ;
  assign \new_[6129]_  = ~\new_[6346]_  | ~\new_[6405]_ ;
  assign \new_[6130]_  = ~\new_[6523]_  | ~\new_[7204]_ ;
  assign \new_[6131]_  = ~\new_[6524]_  | ~\new_[6525]_ ;
  assign \new_[6132]_  = ~\new_[6527]_  | ~\new_[7206]_ ;
  assign \new_[6133]_  = ~\new_[7207]_  | ~\new_[6528]_ ;
  assign \new_[6134]_  = ~\new_[7027]_  | ~\new_[6408]_ ;
  assign \new_[6135]_  = ~\new_[6530]_  | ~\new_[6531]_ ;
  assign \new_[6136]_  = ~\new_[7213]_  | ~\new_[6532]_ ;
  assign \new_[6137]_  = ~\new_[6411]_  | ~\new_[7067]_ ;
  assign \new_[6138]_  = ~\new_[6533]_  | ~\new_[7343]_ ;
  assign \new_[6139]_  = ~\new_[6347]_  & (~\new_[7387]_  | ~\new_[18349]_ );
  assign \new_[6140]_  = ~\new_[6412]_  | ~\new_[7068]_ ;
  assign \new_[6141]_  = ~\new_[6534]_  | ~\new_[7216]_ ;
  assign \new_[6142]_  = ~\new_[6413]_  | ~\new_[7344]_ ;
  assign \new_[6143]_  = ~\new_[7217]_  | ~\new_[6535]_ ;
  assign \new_[6144]_  = ~\new_[7218]_  | ~\new_[6538]_ ;
  assign \new_[6145]_  = ~\new_[6539]_  | ~\new_[7219]_ ;
  assign \new_[6146]_  = ~\new_[7220]_  | ~\new_[6540]_ ;
  assign \new_[6147]_  = ~\new_[6415]_  | ~\new_[7069]_ ;
  assign \new_[6148]_  = ~\new_[6416]_  | ~\new_[7345]_ ;
  assign \new_[6149]_  = ~\new_[7221]_  | ~\new_[6541]_ ;
  assign \new_[6150]_  = ~\new_[6348]_  | ~\new_[6417]_ ;
  assign \new_[6151]_  = ~\new_[6542]_  | ~\new_[7223]_ ;
  assign \new_[6152]_  = ~\new_[6418]_  | ~\new_[7070]_ ;
  assign \new_[6153]_  = ~\new_[7224]_  | ~\new_[6543]_ ;
  assign \new_[6154]_  = ~\new_[6419]_  | ~\new_[7346]_ ;
  assign \new_[6155]_  = ~\new_[6544]_  | ~\new_[6545]_ ;
  assign \new_[6156]_  = ~\new_[6546]_  & (~\new_[8082]_  | ~\new_[18950]_ );
  assign \new_[6157]_  = ~\new_[6547]_  | ~\new_[7347]_ ;
  assign \new_[6158]_  = ~\new_[6548]_  | ~\new_[6549]_ ;
  assign \new_[6159]_  = ~\new_[7225]_  | ~\new_[6550]_ ;
  assign \new_[6160]_  = ~\new_[6349]_  | ~\new_[7072]_ ;
  assign \new_[6161]_  = ~\new_[6420]_  | ~\new_[7073]_ ;
  assign \new_[6162]_  = ~\new_[6936]_  & ~\new_[16658]_ ;
  assign \new_[6163]_  = i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg;
  assign \new_[6164]_  = pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg;
  assign \new_[6165]_  = ~\new_[6936]_ ;
  assign \new_[6166]_  = ~\new_[6936]_ ;
  assign \new_[6167]_  = ~\new_[6969]_  & ~\new_[8115]_ ;
  assign \new_[6168]_  = ~\new_[6970]_  & ~\new_[7401]_ ;
  assign \new_[6169]_  = ~\new_[6971]_  & ~\new_[7402]_ ;
  assign \new_[6170]_  = ~\new_[6972]_  & ~\new_[8124]_ ;
  assign \new_[6171]_  = ~\new_[6973]_  & ~\new_[8297]_ ;
  assign \new_[6172]_  = ~\new_[6974]_  & ~\new_[8128]_ ;
  assign \new_[6173]_  = ~\new_[6976]_  & ~\new_[8130]_ ;
  assign \new_[6174]_  = ~\new_[6977]_  & ~\new_[8131]_ ;
  assign \new_[6175]_  = ~\new_[6978]_  & ~\new_[8133]_ ;
  assign \new_[6176]_  = ~\new_[6979]_  & ~\new_[8136]_ ;
  assign \new_[6177]_  = ~\new_[6981]_  & ~\new_[8137]_ ;
  assign \new_[6178]_  = ~\new_[6982]_  & ~\new_[8140]_ ;
  assign \new_[6179]_  = ~\new_[6983]_  & ~\new_[8146]_ ;
  assign \new_[6180]_  = ~\new_[7407]_  & ~\new_[6984]_ ;
  assign \new_[6181]_  = ~\new_[6989]_  & ~\new_[8157]_ ;
  assign \new_[6182]_  = ~\new_[6990]_  & ~\new_[8338]_ ;
  assign \new_[6183]_  = ~\new_[6991]_  & ~\new_[8341]_ ;
  assign \new_[6184]_  = ~\new_[6992]_  & ~\new_[8162]_ ;
  assign \new_[6185]_  = ~\new_[6993]_  & ~\new_[8166]_ ;
  assign \new_[6186]_  = ~\new_[6994]_  & ~\new_[7411]_ ;
  assign \new_[6187]_  = ~\new_[6996]_  & ~\new_[8171]_ ;
  assign \new_[6188]_  = ~\new_[6997]_  & ~\new_[7414]_ ;
  assign \new_[6189]_  = ~\new_[6998]_  & ~\new_[7417]_ ;
  assign \new_[6190]_  = ~\new_[7001]_  & ~\new_[7240]_ ;
  assign \new_[6191]_  = ~\new_[7003]_  & ~\new_[7421]_ ;
  assign \new_[6192]_  = ~\new_[7004]_  & ~\new_[8183]_ ;
  assign \new_[6193]_  = ~\new_[7005]_  & ~\new_[8187]_ ;
  assign \new_[6194]_  = ~\new_[7006]_  & ~\new_[8191]_ ;
  assign \new_[6195]_  = ~\new_[7008]_  & ~\new_[7426]_ ;
  assign \new_[6196]_  = ~\new_[7010]_  & ~\new_[8195]_ ;
  assign \new_[6197]_  = ~\new_[7011]_  & ~\new_[8197]_ ;
  assign n3125 = ~\new_[7349]_  | ~\new_[7980]_  | ~\new_[7971]_  | ~\new_[7970]_ ;
  assign n3130 = ~\new_[7973]_  | ~\new_[7977]_  | ~\new_[7350]_  | ~\new_[7972]_ ;
  assign n3135 = ~\new_[7976]_  | ~\new_[7975]_  | ~\new_[7351]_  | ~\new_[7974]_ ;
  assign n3140 = ~\new_[7981]_  | ~\new_[7982]_  | ~\new_[7978]_  | ~\new_[7979]_ ;
  assign n3145 = ~\new_[7985]_  | ~\new_[7986]_  | ~\new_[7983]_  | ~\new_[7984]_ ;
  assign n3150 = ~\new_[7989]_  | ~\new_[7990]_  | ~\new_[7987]_  | ~\new_[7988]_ ;
  assign n3015 = ~\new_[8265]_  | ~\new_[7994]_  | ~\new_[7993]_  | ~\new_[7992]_ ;
  assign n3005 = ~\new_[7996]_  | ~\new_[7997]_  | ~\new_[8266]_  | ~\new_[7995]_ ;
  assign n3010 = ~\new_[8000]_  | ~\new_[8001]_  | ~\new_[7998]_  | ~\new_[7999]_ ;
  assign n3020 = ~\new_[8002]_  | ~\new_[8005]_  | ~\new_[8004]_  | ~\new_[8003]_ ;
  assign n3025 = ~\new_[8008]_  | ~\new_[8009]_  | ~\new_[8006]_  | ~\new_[8007]_ ;
  assign n3030 = ~\new_[8011]_  | ~\new_[8012]_  | ~\new_[7354]_  | ~\new_[8010]_ ;
  assign n3035 = ~\new_[8015]_  | ~\new_[8016]_  | ~\new_[8013]_  | ~\new_[8014]_ ;
  assign n3050 = ~\new_[8019]_  | ~\new_[8020]_  | ~\new_[7355]_  | ~\new_[8018]_ ;
  assign n3040 = ~\new_[8023]_  | ~\new_[8024]_  | ~\new_[8021]_  | ~\new_[8022]_ ;
  assign n3045 = ~\new_[8026]_  | ~\new_[8027]_  | ~\new_[8268]_  | ~\new_[8025]_ ;
  assign n3055 = ~\new_[8032]_  | ~\new_[8031]_  | ~\new_[7357]_  | ~\new_[8030]_ ;
  assign n3060 = ~\new_[8270]_  | ~\new_[8035]_  | ~\new_[8034]_  | ~\new_[8033]_ ;
  assign n3065 = ~\new_[8038]_  | ~\new_[8039]_  | ~\new_[8036]_  | ~\new_[8037]_ ;
  assign n3070 = ~\new_[8040]_  | ~\new_[8041]_  | ~\new_[7358]_  | ~\new_[7359]_ ;
  assign n3075 = ~\new_[8043]_  | ~\new_[8044]_  | ~\new_[7360]_  | ~\new_[8042]_ ;
  assign n3080 = ~\new_[8047]_  | ~\new_[8048]_  | ~\new_[8272]_  | ~\new_[8045]_ ;
  assign n3085 = ~\new_[8049]_  | ~\new_[8050]_  | ~\new_[7362]_  | ~\new_[7361]_ ;
  assign n3120 = ~\new_[8052]_  | ~\new_[8053]_  | ~\new_[7363]_  | ~\new_[8051]_ ;
  assign n3090 = ~\new_[8056]_  | ~\new_[8057]_  | ~\new_[7364]_  | ~\new_[8054]_ ;
  assign n3095 = ~\new_[8060]_  | ~\new_[8061]_  | ~\new_[8058]_  | ~\new_[8059]_ ;
  assign n3100 = ~\new_[8064]_  | ~\new_[8065]_  | ~\new_[8062]_  | ~\new_[8063]_ ;
  assign n3105 = ~\new_[8067]_  | ~\new_[8068]_  | ~\new_[7365]_  | ~\new_[8066]_ ;
  assign n3110 = ~\new_[8072]_  | ~\new_[8073]_  | ~\new_[7367]_  | ~\new_[8071]_ ;
  assign n3115 = ~\new_[8076]_  | ~\new_[8077]_  | ~\new_[8074]_  | ~\new_[8075]_ ;
  assign \new_[6228]_  = ~\new_[7087]_  & (~\new_[8096]_  | ~\new_[19651]_ );
  assign \new_[6229]_  = ~\new_[7102]_  | ~\new_[7103]_ ;
  assign \new_[6230]_  = ~\new_[7037]_  | ~\new_[7312]_ ;
  assign \new_[6231]_  = ~\new_[7107]_  | ~\new_[7108]_ ;
  assign \new_[6232]_  = ~\new_[7038]_  | ~\new_[7313]_ ;
  assign \new_[6233]_  = ~\new_[7111]_  | ~\new_[7110]_ ;
  assign \new_[6234]_  = ~\new_[7113]_  | ~\new_[7114]_ ;
  assign \new_[6235]_  = ~\new_[7116]_  | ~\new_[7117]_ ;
  assign \new_[6236]_  = ~\new_[7017]_  | ~\new_[7041]_ ;
  assign \new_[6237]_  = ~\new_[7118]_  & (~\new_[8285]_  | ~\new_[18576]_ );
  assign \new_[6238]_  = ~\new_[7121]_  | ~\new_[7318]_ ;
  assign \new_[6239]_  = ~\new_[7122]_  | ~\new_[7123]_ ;
  assign \new_[6240]_  = ~\new_[7125]_  | ~\new_[7126]_ ;
  assign \new_[6241]_  = ~\new_[7045]_  | ~\new_[7320]_ ;
  assign \new_[6242]_  = ~\new_[7133]_  | ~\new_[7132]_ ;
  assign \new_[6243]_  = ~\new_[7047]_  | ~\new_[7323]_ ;
  assign \new_[6244]_  = ~\new_[7135]_  | ~\new_[7136]_ ;
  assign \new_[6245]_  = ~\new_[7020]_  | ~\new_[7049]_ ;
  assign \new_[6246]_  = ~\new_[7137]_  | ~\new_[7324]_ ;
  assign \new_[6247]_  = ~\new_[7050]_  | ~\new_[7325]_ ;
  assign \new_[6248]_  = ~\new_[7021]_  | ~\new_[7052]_ ;
  assign \new_[6249]_  = ~\new_[7141]_  | ~\new_[7142]_ ;
  assign \new_[6250]_  = ~\new_[7053]_  | ~\new_[7326]_ ;
  assign \new_[6251]_  = ~\new_[7147]_  | ~\new_[7146]_ ;
  assign \new_[6252]_  = ~\new_[7148]_  | ~\new_[7149]_ ;
  assign \new_[6253]_  = ~\new_[7151]_  & (~\new_[8285]_  | ~\new_[18206]_ );
  assign \new_[6254]_  = ~\new_[7155]_  | ~\new_[7156]_ ;
  assign \new_[6255]_  = ~\new_[7159]_  | ~\new_[7160]_ ;
  assign \new_[6256]_  = ~\new_[7168]_  | ~\new_[7169]_ ;
  assign \new_[6257]_  = ~\new_[7170]_  | ~\new_[7171]_ ;
  assign \new_[6258]_  = ~\new_[7180]_  | ~\new_[7181]_ ;
  assign \new_[6259]_  = ~\new_[7058]_  | ~\new_[7333]_ ;
  assign \new_[6260]_  = ~\new_[7059]_  & (~\new_[7375]_  | ~\new_[19503]_ );
  assign \new_[6261]_  = ~\new_[7060]_  | ~\new_[7334]_ ;
  assign \new_[6262]_  = ~\new_[7185]_  | ~\new_[7186]_ ;
  assign \new_[6263]_  = ~\new_[7187]_  | ~\new_[7188]_ ;
  assign \new_[6264]_  = ~\new_[7191]_  | ~\new_[7190]_ ;
  assign \new_[6265]_  = ~\new_[7195]_  | ~\new_[7194]_ ;
  assign \new_[6266]_  = ~\new_[7064]_  | ~\new_[7339]_ ;
  assign \new_[6267]_  = ~\new_[7208]_  | ~\new_[7209]_ ;
  assign \new_[6268]_  = ~\new_[7211]_  | ~\new_[7212]_ ;
  assign \new_[6269]_  = ~\new_[7066]_  | ~\new_[7342]_ ;
  assign \new_[6270]_  = ~\new_[7214]_  | ~\new_[7215]_ ;
  assign \new_[6271]_  = ~\new_[7222]_  & (~\new_[8285]_  | ~\new_[18015]_ );
  assign \new_[6272]_  = ~\new_[7029]_  | ~\new_[7071]_ ;
  assign \new_[6273]_  = ~\new_[7074]_  | ~\new_[7348]_ ;
  assign \new_[6274]_  = ~\new_[7228]_  & (~\new_[7380]_  | ~\new_[19040]_ );
  assign \new_[6275]_  = ~\new_[19879]_  & ~\new_[11687]_ ;
  assign \new_[6276]_  = ~\new_[19879]_  & ~\new_[11727]_ ;
  assign \new_[6277]_  = ~\new_[19880]_  & ~\new_[11356]_ ;
  assign \new_[6278]_  = ~\new_[19879]_  & ~\new_[11650]_ ;
  assign \new_[6279]_  = ~\new_[19880]_  & ~\new_[11617]_ ;
  assign \new_[6280]_  = ~\new_[19877]_  | ~\new_[19030]_ ;
  assign \new_[6281]_  = ~\new_[7231]_  | ~\new_[18765]_ ;
  assign \new_[6282]_  = ~\new_[7231]_  | ~\new_[18842]_ ;
  assign \new_[6283]_  = ~\new_[7372]_  | ~\new_[19513]_ ;
  assign \new_[6284]_  = ~\new_[7372]_  | ~\new_[18470]_ ;
  assign \new_[6285]_  = ~\new_[7372]_  | ~\new_[19295]_ ;
  assign \new_[6286]_  = ~\new_[7372]_  | ~\new_[18985]_ ;
  assign \new_[6287]_  = ~\new_[7372]_  | ~\new_[19340]_ ;
  assign \new_[6288]_  = ~\new_[7372]_  | ~\new_[19374]_ ;
  assign \new_[6289]_  = ~\new_[7372]_  | ~\new_[19521]_ ;
  assign \new_[6290]_  = ~\new_[7233]_  & ~\new_[11647]_ ;
  assign \new_[6291]_  = ~\new_[7232]_  & ~\new_[11739]_ ;
  assign \new_[6292]_  = ~\new_[7233]_  & ~\new_[11510]_ ;
  assign \new_[6293]_  = ~\new_[7232]_  & ~\new_[11780]_ ;
  assign \new_[6294]_  = ~\new_[7232]_  & ~\new_[10936]_ ;
  assign \new_[6295]_  = ~\new_[7232]_  & ~\new_[11784]_ ;
  assign \new_[6296]_  = ~\new_[7232]_  & ~\new_[11493]_ ;
  assign \new_[6297]_  = ~\new_[7233]_  & ~\new_[11637]_ ;
  assign \new_[6298]_  = ~\new_[7232]_  & ~\new_[11774]_ ;
  assign \new_[6299]_  = ~\new_[7233]_  & ~\new_[11879]_ ;
  assign \new_[6300]_  = ~\new_[7232]_  & ~\new_[11723]_ ;
  assign \new_[6301]_  = ~\new_[7233]_  & ~\new_[11523]_ ;
  assign \new_[6302]_  = ~\new_[7232]_  & ~\new_[11711]_ ;
  assign \new_[6303]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11] ;
  assign \new_[6304]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10] ;
  assign \new_[6305]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13] ;
  assign \new_[6306]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14] ;
  assign \new_[6307]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15] ;
  assign \new_[6308]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16] ;
  assign \new_[6309]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17] ;
  assign \new_[6310]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19] ;
  assign \new_[6311]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20] ;
  assign \new_[6312]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21] ;
  assign \new_[6313]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23] ;
  assign \new_[6314]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24] ;
  assign \new_[6315]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25] ;
  assign \new_[6316]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27] ;
  assign \new_[6317]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12] ;
  assign \new_[6318]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29] ;
  assign \new_[6319]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30] ;
  assign \new_[6320]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31] ;
  assign \new_[6321]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3] ;
  assign \new_[6322]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5] ;
  assign \new_[6323]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6] ;
  assign \new_[6324]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7] ;
  assign \new_[6325]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9] ;
  assign \new_[6326]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28] ;
  assign \new_[6327]_  = i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg;
  assign \new_[6328]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22] ;
  assign \new_[6329]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18] ;
  assign \new_[6330]_  = \new_[6936]_ ;
  assign \new_[6331]_  = ~\new_[7302]_  & ~\new_[7405]_ ;
  assign \new_[6332]_  = ~\new_[7303]_  & ~\new_[8152]_ ;
  assign \new_[6333]_  = ~\new_[7304]_  & ~\new_[8164]_ ;
  assign \new_[6334]_  = ~\new_[9175]_  | ~\new_[8637]_  | ~\new_[9174]_  | ~\new_[8154]_ ;
  assign \new_[6335]_  = ~\new_[19877]_  | ~\new_[18141]_ ;
  assign \new_[6336]_  = ~\new_[19876]_  | ~\new_[18391]_ ;
  assign \new_[6337]_  = ~\new_[19877]_  | ~\new_[18143]_ ;
  assign \new_[6338]_  = ~\new_[19876]_  | ~\new_[18221]_ ;
  assign \new_[6339]_  = ~\new_[19876]_  | ~\new_[19231]_ ;
  assign \new_[6340]_  = ~\new_[19877]_  | ~\new_[19248]_ ;
  assign \new_[6341]_  = ~\new_[19878]_  & ~\new_[11360]_ ;
  assign \new_[6342]_  = ~\new_[19878]_  & ~\new_[11363]_ ;
  assign \new_[6343]_  = ~\new_[19876]_  | ~\new_[18250]_ ;
  assign \new_[6344]_  = ~\new_[19877]_  | ~\new_[18248]_ ;
  assign \new_[6345]_  = ~\new_[19878]_  & ~\new_[11365]_ ;
  assign \new_[6346]_  = ~\new_[19876]_  | ~\new_[18136]_ ;
  assign \new_[6347]_  = ~\new_[19878]_  & ~\new_[11349]_ ;
  assign \new_[6348]_  = ~\new_[19877]_  | ~\new_[19412]_ ;
  assign \new_[6349]_  = ~\new_[19877]_  | ~\new_[19415]_ ;
  assign \new_[6350]_  = ~\new_[7369]_  | ~\new_[19213]_ ;
  assign \new_[6351]_  = ~\new_[7372]_  | ~\new_[19382]_ ;
  assign \new_[6352]_  = ~\new_[7373]_  | ~\new_[18467]_ ;
  assign \new_[6353]_  = ~\new_[7368]_  & ~\new_[11498]_ ;
  assign \new_[6354]_  = ~\new_[7387]_  | ~\new_[19084]_ ;
  assign \new_[6355]_  = ~\new_[7373]_  | ~\new_[18479]_ ;
  assign \new_[6356]_  = ~\new_[7376]_  | ~\new_[18880]_ ;
  assign \new_[6357]_  = ~\new_[7373]_  | ~\new_[18546]_ ;
  assign \new_[6358]_  = ~\new_[7371]_  | ~\new_[19215]_ ;
  assign \new_[6359]_  = ~\new_[7376]_  | ~\new_[18643]_ ;
  assign \new_[6360]_  = ~\new_[7387]_  | ~\new_[17968]_ ;
  assign \new_[6361]_  = ~\new_[7376]_  | ~\new_[18602]_ ;
  assign \new_[6362]_  = ~\new_[7374]_  | ~\new_[18883]_ ;
  assign \new_[6363]_  = ~\new_[7370]_  | ~\new_[19220]_ ;
  assign \new_[6364]_  = ~\new_[7369]_  | ~\new_[19599]_ ;
  assign \new_[6365]_  = ~\new_[7373]_  | ~\new_[18473]_ ;
  assign \new_[6366]_  = ~\new_[7369]_  | ~\new_[18721]_ ;
  assign \new_[6367]_  = ~\new_[7372]_  | ~\new_[17932]_ ;
  assign \new_[6368]_  = ~\new_[7387]_  | ~\new_[19099]_ ;
  assign \new_[6369]_  = ~\new_[7369]_  | ~\new_[18743]_ ;
  assign \new_[6370]_  = ~\new_[7375]_  | ~\new_[18478]_ ;
  assign \new_[6371]_  = ~\new_[7387]_  | ~\new_[19093]_ ;
  assign \new_[6372]_  = ~\new_[7387]_  | ~\new_[19631]_ ;
  assign \new_[6373]_  = ~\new_[7372]_  | ~\new_[19510]_ ;
  assign \new_[6374]_  = ~\new_[7369]_  | ~\new_[18817]_ ;
  assign \new_[6375]_  = ~\new_[7372]_  | ~\new_[19511]_ ;
  assign \new_[6376]_  = ~\new_[7374]_  | ~\new_[18734]_ ;
  assign \new_[6377]_  = ~\new_[7375]_  | ~\new_[19507]_ ;
  assign \new_[6378]_  = ~\new_[7387]_  | ~\new_[17870]_ ;
  assign \new_[6379]_  = ~\new_[7376]_  | ~\new_[18793]_ ;
  assign \new_[6380]_  = ~\new_[7368]_  & ~\new_[11699]_ ;
  assign \new_[6381]_  = ~\new_[7372]_  | ~\new_[19155]_ ;
  assign \new_[6382]_  = ~\new_[7387]_  | ~\new_[18970]_ ;
  assign \new_[6383]_  = ~\new_[7371]_  | ~\new_[18414]_ ;
  assign \new_[6384]_  = ~\new_[7375]_  | ~\new_[19553]_ ;
  assign \new_[6385]_  = ~\new_[7376]_  | ~\new_[18918]_ ;
  assign \new_[6386]_  = ~\new_[7372]_  | ~\new_[17934]_ ;
  assign \new_[6387]_  = ~\new_[7371]_  | ~\new_[18144]_ ;
  assign \new_[6388]_  = ~\new_[7387]_  | ~\new_[19484]_ ;
  assign \new_[6389]_  = ~\new_[7374]_  | ~\new_[18646]_ ;
  assign \new_[6390]_  = ~\new_[7371]_  | ~\new_[19328]_ ;
  assign \new_[6391]_  = ~\new_[7387]_  | ~\new_[17974]_ ;
  assign \new_[6392]_  = ~\new_[7369]_  | ~\new_[19221]_ ;
  assign \new_[6393]_  = ~\new_[7372]_  | ~\new_[19339]_ ;
  assign \new_[6394]_  = ~\new_[7387]_  | ~\new_[17975]_ ;
  assign \new_[6395]_  = ~\new_[7376]_  | ~\new_[18593]_ ;
  assign \new_[6396]_  = ~\new_[7387]_  | ~\new_[18078]_ ;
  assign \new_[6397]_  = ~\new_[7372]_  | ~\new_[18495]_ ;
  assign \new_[6398]_  = ~\new_[7370]_  | ~\new_[18319]_ ;
  assign \new_[6399]_  = ~\new_[7375]_  | ~\new_[19024]_ ;
  assign \new_[6400]_  = ~\new_[7373]_  | ~\new_[18550]_ ;
  assign \new_[6401]_  = ~\new_[7371]_  | ~\new_[18620]_ ;
  assign \new_[6402]_  = ~\new_[7387]_  | ~\new_[19482]_ ;
  assign \new_[6403]_  = ~\new_[7374]_  | ~\new_[18449]_ ;
  assign \new_[6404]_  = ~\new_[7387]_  | ~\new_[19695]_ ;
  assign \new_[6405]_  = ~\new_[7387]_  | ~\new_[19430]_ ;
  assign \new_[6406]_  = ~\new_[7370]_  | ~\new_[18867]_ ;
  assign \new_[6407]_  = ~\new_[7376]_  | ~\new_[19505]_ ;
  assign \new_[6408]_  = ~\new_[7387]_  | ~\new_[19045]_ ;
  assign \new_[6409]_  = ~\new_[7376]_  | ~\new_[17842]_ ;
  assign \new_[6410]_  = ~\new_[7370]_  | ~\new_[18859]_ ;
  assign \new_[6411]_  = ~\new_[7375]_  | ~\new_[19376]_ ;
  assign \new_[6412]_  = ~\new_[7373]_  | ~\new_[18244]_ ;
  assign \new_[6413]_  = ~\new_[7370]_  | ~\new_[18750]_ ;
  assign \new_[6414]_  = ~\new_[7387]_  | ~\new_[17965]_ ;
  assign \new_[6415]_  = ~\new_[7372]_  | ~\new_[19516]_ ;
  assign \new_[6416]_  = ~\new_[7371]_  | ~\new_[18855]_ ;
  assign \new_[6417]_  = ~\new_[7387]_  | ~\new_[19489]_ ;
  assign \new_[6418]_  = ~\new_[7374]_  | ~\new_[18995]_ ;
  assign \new_[6419]_  = ~\new_[7371]_  | ~\new_[19464]_ ;
  assign \new_[6420]_  = ~\new_[7373]_  | ~\new_[18463]_ ;
  assign \new_[6421]_  = ~\new_[7390]_  | ~\new_[18862]_ ;
  assign \new_[6422]_  = ~\new_[7380]_  | ~\new_[18829]_ ;
  assign \new_[6423]_  = ~\new_[7385]_  | ~\new_[18850]_ ;
  assign \new_[6424]_  = ~\new_[7381]_  | ~\new_[19468]_ ;
  assign \new_[6425]_  = ~\new_[7394]_  | ~\new_[18026]_ ;
  assign \new_[6426]_  = ~\new_[7400]_  | ~\new_[18128]_ ;
  assign \new_[6427]_  = ~\new_[7386]_  | ~\new_[19327]_ ;
  assign \new_[6428]_  = ~\new_[7393]_  | ~\new_[19348]_ ;
  assign \new_[6429]_  = ~\new_[8096]_  | ~\new_[19676]_ ;
  assign \new_[6430]_  = ~\new_[7392]_  | ~\new_[19375]_ ;
  assign \new_[6431]_  = ~\new_[7381]_  | ~\new_[18447]_ ;
  assign \new_[6432]_  = ~\new_[7394]_  | ~\new_[19177]_ ;
  assign \new_[6433]_  = ~\new_[7399]_  | ~\new_[18011]_ ;
  assign \new_[6434]_  = ~\new_[7386]_  | ~\new_[19539]_ ;
  assign \new_[6435]_  = ~\new_[7392]_  | ~\new_[18336]_ ;
  assign \new_[6436]_  = ~\new_[7400]_  | ~\new_[19456]_ ;
  assign \new_[6437]_  = ~\new_[7394]_  | ~\new_[19170]_ ;
  assign \new_[6438]_  = ~\new_[18644]_  | ~\new_[7381]_ ;
  assign \new_[6439]_  = ~\new_[7389]_  | ~\new_[19871]_ ;
  assign \new_[6440]_  = ~\new_[7378]_  | ~\new_[17828]_ ;
  assign \new_[6441]_  = ~\new_[7391]_  | ~\new_[18474]_ ;
  assign \new_[6442]_  = ~\new_[7385]_  | ~\new_[18454]_ ;
  assign \new_[6443]_  = ~\new_[7394]_  | ~\new_[19644]_ ;
  assign \new_[6444]_  = ~\new_[7381]_  | ~\new_[19429]_ ;
  assign \new_[6445]_  = ~\new_[7379]_  | ~\new_[19836]_ ;
  assign \new_[6446]_  = ~\new_[7388]_  & ~\new_[11798]_ ;
  assign \new_[6447]_  = ~\new_[7399]_  | ~\new_[18013]_ ;
  assign \new_[6448]_  = ~\new_[7381]_  | ~\new_[19847]_ ;
  assign \new_[6449]_  = ~\new_[7379]_  | ~\new_[17923]_ ;
  assign \new_[6450]_  = ~\new_[7388]_  & ~\new_[11437]_ ;
  assign \new_[6451]_  = ~\new_[7380]_  | ~\new_[18728]_ ;
  assign \new_[6452]_  = ~\new_[7394]_  | ~\new_[18043]_ ;
  assign \new_[6453]_  = ~\new_[7396]_  & ~\new_[11646]_ ;
  assign \new_[6454]_  = ~\new_[7391]_  | ~\new_[19629]_ ;
  assign \new_[6455]_  = ~\new_[7382]_  & ~\new_[11860]_ ;
  assign \new_[6456]_  = ~\new_[7386]_  | ~\new_[19536]_ ;
  assign \new_[6457]_  = ~\new_[7399]_  | ~\new_[18130]_ ;
  assign \new_[6458]_  = ~\new_[7377]_  | ~\new_[19128]_ ;
  assign \new_[6459]_  = ~\new_[7389]_  | ~\new_[19654]_ ;
  assign \new_[6460]_  = ~\new_[11797]_  & ~\new_[7383]_ ;
  assign \new_[6461]_  = ~\new_[7377]_  | ~\new_[18003]_ ;
  assign \new_[6462]_  = ~\new_[7396]_  & ~\new_[11509]_ ;
  assign \new_[6463]_  = ~\new_[7395]_  | ~\new_[18048]_ ;
  assign \new_[6464]_  = ~\new_[7386]_  | ~\new_[18320]_ ;
  assign \new_[6465]_  = ~\new_[7397]_  | ~\new_[19588]_ ;
  assign \new_[6466]_  = ~\new_[7393]_  | ~\new_[18397]_ ;
  assign \new_[6467]_  = ~\new_[7380]_  | ~\new_[18824]_ ;
  assign \new_[6468]_  = ~\new_[7388]_  & ~\new_[11737]_ ;
  assign \new_[6469]_  = ~\new_[7377]_  | ~\new_[19619]_ ;
  assign \new_[6470]_  = ~\new_[7389]_  | ~\new_[17960]_ ;
  assign \new_[6471]_  = ~\new_[7394]_  | ~\new_[19135]_ ;
  assign \new_[6472]_  = ~\new_[7391]_  | ~\new_[17961]_ ;
  assign \new_[6473]_  = ~\new_[7382]_  & ~\new_[11542]_ ;
  assign \new_[6474]_  = ~\new_[7396]_  & ~\new_[11511]_ ;
  assign \new_[6475]_  = ~\new_[7378]_  | ~\new_[18658]_ ;
  assign \new_[6476]_  = ~\new_[7391]_  | ~\new_[19666]_ ;
  assign \new_[6477]_  = ~\new_[7399]_  | ~\new_[19587]_ ;
  assign \new_[6478]_  = ~\new_[7386]_  | ~\new_[19533]_ ;
  assign \new_[6479]_  = ~\new_[7384]_  & ~\new_[11854]_ ;
  assign \new_[6480]_  = ~\new_[7381]_  | ~\new_[18417]_ ;
  assign \new_[6481]_  = ~\new_[7398]_  | ~\new_[18965]_ ;
  assign \new_[6482]_  = ~\new_[7386]_  | ~\new_[18330]_ ;
  assign \new_[6483]_  = ~\new_[7379]_  | ~\new_[18690]_ ;
  assign \new_[6484]_  = ~\new_[7392]_  | ~\new_[18998]_ ;
  assign \new_[6485]_  = ~\new_[7392]_  | ~\new_[18911]_ ;
  assign \new_[6486]_  = ~\new_[7398]_  | ~\new_[18137]_ ;
  assign \new_[6487]_  = ~\new_[7397]_  | ~\new_[18739]_ ;
  assign \new_[6488]_  = ~\new_[8287]_  | ~\new_[18689]_ ;
  assign \new_[6489]_  = ~\new_[7378]_  | ~\new_[18448]_ ;
  assign \new_[6490]_  = ~\new_[7397]_  | ~\new_[19403]_ ;
  assign \new_[6491]_  = ~\new_[7386]_  | ~\new_[19277]_ ;
  assign \new_[6492]_  = ~\new_[7385]_  | ~\new_[18815]_ ;
  assign \new_[6493]_  = ~\new_[7390]_  | ~\new_[19311]_ ;
  assign \new_[6494]_  = ~\new_[7377]_  | ~\new_[17970]_ ;
  assign \new_[6495]_  = ~\new_[7397]_  | ~\new_[19831]_ ;
  assign \new_[6496]_  = ~\new_[7386]_  | ~\new_[18358]_ ;
  assign \new_[6497]_  = ~\new_[7385]_  | ~\new_[18648]_ ;
  assign \new_[6498]_  = ~\new_[7377]_  | ~\new_[19851]_ ;
  assign \new_[6499]_  = ~\new_[7389]_  | ~\new_[18872]_ ;
  assign \new_[6500]_  = ~\new_[7394]_  | ~\new_[18280]_ ;
  assign \new_[6501]_  = ~\new_[7386]_  | ~\new_[18792]_ ;
  assign \new_[6502]_  = ~\new_[7381]_  | ~\new_[19609]_ ;
  assign \new_[6503]_  = ~\new_[8096]_  | ~\new_[19351]_ ;
  assign \new_[6504]_  = ~\new_[7393]_  | ~\new_[19422]_ ;
  assign \new_[6505]_  = ~\new_[7400]_  | ~\new_[18138]_ ;
  assign \new_[6506]_  = ~\new_[7394]_  | ~\new_[18145]_ ;
  assign \new_[6507]_  = ~\new_[7381]_  | ~\new_[19628]_ ;
  assign \new_[6508]_  = ~\new_[7379]_  | ~\new_[19486]_ ;
  assign \new_[6509]_  = ~\new_[7392]_  | ~\new_[19850]_ ;
  assign \new_[6510]_  = ~\new_[7380]_  | ~\new_[19239]_ ;
  assign \new_[6511]_  = ~\new_[7394]_  | ~\new_[18109]_ ;
  assign \new_[6512]_  = ~\new_[7396]_  & ~\new_[11516]_ ;
  assign \new_[6513]_  = ~\new_[7378]_  | ~\new_[18426]_ ;
  assign \new_[6514]_  = ~\new_[7394]_  | ~\new_[18672]_ ;
  assign \new_[6515]_  = ~\new_[7378]_  | ~\new_[18087]_ ;
  assign \new_[6516]_  = ~\new_[7391]_  | ~\new_[19848]_ ;
  assign \new_[6517]_  = ~\new_[7396]_  & ~\new_[11517]_ ;
  assign \new_[6518]_  = ~\new_[7391]_  | ~\new_[19453]_ ;
  assign \new_[6519]_  = ~\new_[7380]_  | ~\new_[18813]_ ;
  assign \new_[6520]_  = ~\new_[7382]_  & ~\new_[11269]_ ;
  assign \new_[6521]_  = ~\new_[7400]_  | ~\new_[18916]_ ;
  assign \new_[6522]_  = ~\new_[7394]_  | ~\new_[18405]_ ;
  assign \new_[6523]_  = ~\new_[7381]_  | ~\new_[19130]_ ;
  assign \new_[6524]_  = ~\new_[7393]_  | ~\new_[18365]_ ;
  assign \new_[6525]_  = ~\new_[8096]_  | ~\new_[19866]_ ;
  assign \new_[6526]_  = ~\new_[7389]_  | ~\new_[18183]_ ;
  assign \new_[6527]_  = ~\new_[7400]_  | ~\new_[19458]_ ;
  assign \new_[6528]_  = ~\new_[7381]_  | ~\new_[19001]_ ;
  assign \new_[6529]_  = ~\new_[7389]_  | ~\new_[19398]_ ;
  assign \new_[6530]_  = ~\new_[7393]_  | ~\new_[18369]_ ;
  assign \new_[6531]_  = ~\new_[8096]_  | ~\new_[18875]_ ;
  assign \new_[6532]_  = ~\new_[7378]_  | ~\new_[19701]_ ;
  assign \new_[6533]_  = ~\new_[7394]_  | ~\new_[18209]_ ;
  assign \new_[6534]_  = ~\new_[7392]_  | ~\new_[17890]_ ;
  assign \new_[6535]_  = ~\new_[7380]_  | ~\new_[18154]_ ;
  assign \new_[6536]_  = ~\new_[7386]_  | ~\new_[19540]_ ;
  assign \new_[6537]_  = ~\new_[7397]_  | ~\new_[18587]_ ;
  assign \new_[6538]_  = ~\new_[7385]_  | ~\new_[19705]_ ;
  assign \new_[6539]_  = ~\new_[7390]_  | ~\new_[17827]_ ;
  assign \new_[6540]_  = ~\new_[7378]_  | ~\new_[19633]_ ;
  assign \new_[6541]_  = ~\new_[7381]_  | ~\new_[18892]_ ;
  assign \new_[6542]_  = ~\new_[7390]_  | ~\new_[17869]_ ;
  assign \new_[6543]_  = ~\new_[7379]_  | ~\new_[18451]_ ;
  assign \new_[6544]_  = ~\new_[7399]_  | ~\new_[18009]_ ;
  assign \new_[6545]_  = ~\new_[7386]_  | ~\new_[19509]_ ;
  assign \new_[6546]_  = ~\new_[7384]_  & ~\new_[11949]_ ;
  assign \new_[6547]_  = ~\new_[7394]_  | ~\new_[19586]_ ;
  assign \new_[6548]_  = ~\new_[7398]_  | ~\new_[19457]_ ;
  assign \new_[6549]_  = ~\new_[7386]_  | ~\new_[19596]_ ;
  assign \new_[6550]_  = ~\new_[7381]_  | ~\new_[19770]_ ;
  assign \new_[6551]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8] ;
  assign \new_[6552]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26] ;
  assign \new_[6553]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4] ;
  assign \new_[6554]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2] ;
  assign \new_[6555]_  = ~\new_[15904]_  | ~\new_[15992]_  | ~\new_[20026]_  | ~\new_[17123]_ ;
  assign \new_[6556]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][11] ;
  assign \new_[6557]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][19] ;
  assign \new_[6558]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][19] ;
  assign \pci_ad_oe_o[23]  = pci_io_mux_ad_iob23_en_out_reg;
  assign \pci_ad_oe_o[22]  = pci_io_mux_ad_iob22_en_out_reg;
  assign \pci_ad_oe_o[21]  = pci_io_mux_ad_iob21_en_out_reg;
  assign \pci_ad_oe_o[19]  = pci_io_mux_ad_iob19_en_out_reg;
  assign \pci_ad_oe_o[17]  = pci_io_mux_ad_iob17_en_out_reg;
  assign \pci_ad_oe_o[18]  = pci_io_mux_ad_iob18_en_out_reg;
  assign \pci_ad_oe_o[15]  = pci_io_mux_ad_iob15_en_out_reg;
  assign \pci_ad_oe_o[14]  = pci_io_mux_ad_iob14_en_out_reg;
  assign \pci_ad_oe_o[13]  = pci_io_mux_ad_iob13_en_out_reg;
  assign \pci_ad_oe_o[11]  = pci_io_mux_ad_iob11_en_out_reg;
  assign \pci_ad_oe_o[25]  = pci_io_mux_ad_iob25_en_out_reg;
  assign \pci_ad_oe_o[8]  = pci_io_mux_ad_iob8_en_out_reg;
  assign \pci_ad_oe_o[7]  = pci_io_mux_ad_iob7_en_out_reg;
  assign \pci_ad_oe_o[9]  = pci_io_mux_ad_iob9_en_out_reg;
  assign \pci_ad_oe_o[5]  = pci_io_mux_ad_iob5_en_out_reg;
  assign \pci_ad_oe_o[3]  = pci_io_mux_ad_iob3_en_out_reg;
  assign \pci_ad_oe_o[4]  = pci_io_mux_ad_iob4_en_out_reg;
  assign \pci_ad_oe_o[1]  = pci_io_mux_ad_iob1_en_out_reg;
  assign \pci_ad_oe_o[2]  = pci_io_mux_ad_iob2_en_out_reg;
  assign \pci_ad_oe_o[26]  = pci_io_mux_ad_iob26_en_out_reg;
  assign \pci_ad_oe_o[31]  = pci_io_mux_ad_iob31_en_out_reg;
  assign \pci_ad_oe_o[29]  = pci_io_mux_ad_iob29_en_out_reg;
  assign \pci_ad_oe_o[28]  = pci_io_mux_ad_iob28_en_out_reg;
  assign \pci_ad_oe_o[27]  = pci_io_mux_ad_iob27_en_out_reg;
  assign \new_[6583]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][35] ;
  assign \new_[6584]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][35] ;
  assign \new_[6585]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][35] ;
  assign \new_[6586]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][35] ;
  assign \new_[6587]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][35] ;
  assign \new_[6588]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][35] ;
  assign \new_[6589]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][35] ;
  assign \new_[6590]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][35] ;
  assign \new_[6591]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][35] ;
  assign \new_[6592]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][0] ;
  assign \new_[6593]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][10] ;
  assign \new_[6594]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][11] ;
  assign \new_[6595]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][13] ;
  assign \new_[6596]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][15] ;
  assign \new_[6597]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][16] ;
  assign \new_[6598]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][17] ;
  assign \new_[6599]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][18] ;
  assign \new_[6600]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][19] ;
  assign \new_[6601]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][20] ;
  assign \new_[6602]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][21] ;
  assign \new_[6603]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][23] ;
  assign \new_[6604]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][24] ;
  assign \new_[6605]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][26] ;
  assign \new_[6606]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][28] ;
  assign \new_[6607]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][29] ;
  assign \new_[6608]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][30] ;
  assign \new_[6609]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][31] ;
  assign \new_[6610]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][3] ;
  assign \new_[6611]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][7] ;
  assign \new_[6612]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][8] ;
  assign \new_[6613]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][9] ;
  assign \new_[6614]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][10] ;
  assign \new_[6615]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][11] ;
  assign \new_[6616]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][13] ;
  assign \new_[6617]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][15] ;
  assign \new_[6618]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][16] ;
  assign \new_[6619]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][18] ;
  assign \new_[6620]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][19] ;
  assign \new_[6621]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][20] ;
  assign \new_[6622]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][23] ;
  assign \new_[6623]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][24] ;
  assign \new_[6624]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][26] ;
  assign \new_[6625]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][27] ;
  assign \new_[6626]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][1] ;
  assign \new_[6627]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][30] ;
  assign \new_[6628]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][31] ;
  assign \new_[6629]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][3] ;
  assign \new_[6630]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][7] ;
  assign \new_[6631]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][8] ;
  assign \new_[6632]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][9] ;
  assign \new_[6633]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][0] ;
  assign \new_[6634]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][11] ;
  assign \new_[6635]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][13] ;
  assign \new_[6636]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][15] ;
  assign \new_[6637]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][16] ;
  assign \new_[6638]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][17] ;
  assign \new_[6639]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][18] ;
  assign \new_[6640]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][19] ;
  assign \new_[6641]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][1] ;
  assign \new_[6642]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][20] ;
  assign \new_[6643]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][23] ;
  assign \new_[6644]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][24] ;
  assign \new_[6645]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][26] ;
  assign \new_[6646]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][27] ;
  assign \new_[6647]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][28] ;
  assign \new_[6648]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][30] ;
  assign \new_[6649]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][31] ;
  assign \new_[6650]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][3] ;
  assign \new_[6651]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][7] ;
  assign \new_[6652]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][8] ;
  assign \new_[6653]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][9] ;
  assign \new_[6654]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][0] ;
  assign \new_[6655]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][10] ;
  assign \new_[6656]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][13] ;
  assign \new_[6657]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][15] ;
  assign \new_[6658]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][16] ;
  assign \new_[6659]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][17] ;
  assign \new_[6660]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][18] ;
  assign \new_[6661]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][1] ;
  assign \new_[6662]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][20] ;
  assign \new_[6663]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][21] ;
  assign \new_[6664]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][23] ;
  assign \new_[6665]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][24] ;
  assign \new_[6666]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][26] ;
  assign \new_[6667]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][27] ;
  assign \new_[6668]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][28] ;
  assign \new_[6669]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][29] ;
  assign \new_[6670]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][30] ;
  assign \new_[6671]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][31] ;
  assign \new_[6672]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][3] ;
  assign \new_[6673]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][7] ;
  assign \new_[6674]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][8] ;
  assign \new_[6675]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][0] ;
  assign \new_[6676]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][10] ;
  assign \new_[6677]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][11] ;
  assign \new_[6678]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][13] ;
  assign \new_[6679]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][15] ;
  assign \new_[6680]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][17] ;
  assign \new_[6681]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][18] ;
  assign \new_[6682]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][19] ;
  assign \new_[6683]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][20] ;
  assign \new_[6684]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][21] ;
  assign \new_[6685]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][23] ;
  assign \new_[6686]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][24] ;
  assign \new_[6687]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][26] ;
  assign \new_[6688]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][27] ;
  assign \new_[6689]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][28] ;
  assign \new_[6690]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][29] ;
  assign \new_[6691]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][30] ;
  assign \new_[6692]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][31] ;
  assign \new_[6693]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][3] ;
  assign \new_[6694]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][7] ;
  assign \new_[6695]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][8] ;
  assign \new_[6696]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][9] ;
  assign \new_[6697]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][10] ;
  assign \new_[6698]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][11] ;
  assign \new_[6699]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][13] ;
  assign \new_[6700]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][15] ;
  assign \new_[6701]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][16] ;
  assign \new_[6702]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][17] ;
  assign \new_[6703]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][18] ;
  assign \new_[6704]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][19] ;
  assign \new_[6705]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][1] ;
  assign \new_[6706]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][21] ;
  assign \new_[6707]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][23] ;
  assign \new_[6708]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][24] ;
  assign \new_[6709]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][26] ;
  assign \new_[6710]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][27] ;
  assign \new_[6711]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][29] ;
  assign \new_[6712]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][30] ;
  assign \new_[6713]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][31] ;
  assign \new_[6714]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][3] ;
  assign \new_[6715]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][7] ;
  assign \new_[6716]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][8] ;
  assign \new_[6717]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][9] ;
  assign \new_[6718]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][0] ;
  assign \new_[6719]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][11] ;
  assign \new_[6720]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][13] ;
  assign \new_[6721]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][15] ;
  assign \new_[6722]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][16] ;
  assign \new_[6723]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][17] ;
  assign \new_[6724]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][19] ;
  assign \new_[6725]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][1] ;
  assign \new_[6726]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][20] ;
  assign \new_[6727]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][21] ;
  assign \new_[6728]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][23] ;
  assign \new_[6729]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][24] ;
  assign \new_[6730]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][26] ;
  assign \new_[6731]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][27] ;
  assign \new_[6732]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][28] ;
  assign \new_[6733]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][30] ;
  assign \new_[6734]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][31] ;
  assign \new_[6735]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][7] ;
  assign \new_[6736]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][8] ;
  assign \new_[6737]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][9] ;
  assign \new_[6738]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][0] ;
  assign \new_[6739]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][11] ;
  assign \new_[6740]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][13] ;
  assign \new_[6741]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][15] ;
  assign \new_[6742]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][16] ;
  assign \new_[6743]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][17] ;
  assign \new_[6744]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][19] ;
  assign \new_[6745]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][1] ;
  assign \new_[6746]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][20] ;
  assign \new_[6747]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][21] ;
  assign \new_[6748]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][23] ;
  assign \new_[6749]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][24] ;
  assign \new_[6750]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][26] ;
  assign \new_[6751]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][27] ;
  assign \new_[6752]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][28] ;
  assign \new_[6753]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][30] ;
  assign \new_[6754]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][31] ;
  assign \new_[6755]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][7] ;
  assign \new_[6756]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][8] ;
  assign \new_[6757]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][9] ;
  assign \new_[6758]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][0] ;
  assign \new_[6759]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][11] ;
  assign \new_[6760]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][13] ;
  assign \new_[6761]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][15] ;
  assign \new_[6762]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][16] ;
  assign \new_[6763]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][18] ;
  assign \new_[6764]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][1] ;
  assign \new_[6765]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][20] ;
  assign \new_[6766]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][21] ;
  assign \new_[6767]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][23] ;
  assign \new_[6768]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][24] ;
  assign \new_[6769]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][26] ;
  assign \new_[6770]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][27] ;
  assign \new_[6771]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][28] ;
  assign \new_[6772]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][29] ;
  assign \new_[6773]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][30] ;
  assign \new_[6774]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][31] ;
  assign \new_[6775]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][3] ;
  assign \new_[6776]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][7] ;
  assign \new_[6777]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][8] ;
  assign \new_[6778]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][17] ;
  assign \new_[6779]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][9] ;
  assign \new_[6780]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][0] ;
  assign \new_[6781]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][11] ;
  assign \new_[6782]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][13] ;
  assign \new_[6783]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][15] ;
  assign \new_[6784]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][16] ;
  assign \new_[6785]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][17] ;
  assign \new_[6786]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][19] ;
  assign \new_[6787]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][1] ;
  assign \new_[6788]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][20] ;
  assign \new_[6789]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][23] ;
  assign \new_[6790]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][24] ;
  assign \new_[6791]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][26] ;
  assign \new_[6792]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][27] ;
  assign \new_[6793]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][28] ;
  assign \new_[6794]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][30] ;
  assign \new_[6795]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][31] ;
  assign \new_[6796]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][7] ;
  assign \new_[6797]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][8] ;
  assign \new_[6798]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][9] ;
  assign \new_[6799]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][0] ;
  assign \new_[6800]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][11] ;
  assign \new_[6801]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][13] ;
  assign \new_[6802]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][15] ;
  assign \new_[6803]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][16] ;
  assign \new_[6804]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][17] ;
  assign \new_[6805]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][19] ;
  assign \new_[6806]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][1] ;
  assign \new_[6807]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][20] ;
  assign \new_[6808]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][21] ;
  assign \new_[6809]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][23] ;
  assign \new_[6810]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][24] ;
  assign \new_[6811]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][26] ;
  assign \new_[6812]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][27] ;
  assign \new_[6813]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][28] ;
  assign \new_[6814]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][30] ;
  assign \new_[6815]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][31] ;
  assign \new_[6816]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][7] ;
  assign \new_[6817]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][8] ;
  assign \new_[6818]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][9] ;
  assign \new_[6819]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][0] ;
  assign \new_[6820]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][10] ;
  assign \new_[6821]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][11] ;
  assign \new_[6822]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][13] ;
  assign \new_[6823]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][15] ;
  assign \new_[6824]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][16] ;
  assign \new_[6825]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][17] ;
  assign \new_[6826]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][18] ;
  assign \new_[6827]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][1] ;
  assign \new_[6828]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][20] ;
  assign \new_[6829]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][21] ;
  assign \new_[6830]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][23] ;
  assign \new_[6831]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][24] ;
  assign \new_[6832]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][26] ;
  assign \new_[6833]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][27] ;
  assign \new_[6834]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][28] ;
  assign \new_[6835]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][29] ;
  assign \new_[6836]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][30] ;
  assign \new_[6837]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][31] ;
  assign \new_[6838]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][35] ;
  assign \new_[6839]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][3] ;
  assign \new_[6840]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][7] ;
  assign \new_[6841]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][9] ;
  assign \new_[6842]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][8] ;
  assign \new_[6843]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][0] ;
  assign \new_[6844]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][10] ;
  assign \new_[6845]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][13] ;
  assign \new_[6846]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][15] ;
  assign \new_[6847]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][16] ;
  assign \new_[6848]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][17] ;
  assign \new_[6849]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][18] ;
  assign \new_[6850]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][1] ;
  assign \new_[6851]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][20] ;
  assign \new_[6852]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][21] ;
  assign \new_[6853]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][23] ;
  assign \new_[6854]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][24] ;
  assign \new_[6855]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][26] ;
  assign \new_[6856]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][27] ;
  assign \new_[6857]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][28] ;
  assign \new_[6858]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][29] ;
  assign \new_[6859]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][30] ;
  assign \new_[6860]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][31] ;
  assign \new_[6861]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][35] ;
  assign \new_[6862]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][3] ;
  assign \new_[6863]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][7] ;
  assign \new_[6864]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][8] ;
  assign \new_[6865]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][9] ;
  assign \new_[6866]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][0] ;
  assign \new_[6867]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][10] ;
  assign \new_[6868]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][11] ;
  assign \new_[6869]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][13] ;
  assign \new_[6870]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][15] ;
  assign \new_[6871]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][16] ;
  assign \new_[6872]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][17] ;
  assign \new_[6873]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][18] ;
  assign \new_[6874]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][1] ;
  assign \new_[6875]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][20] ;
  assign \new_[6876]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][21] ;
  assign \new_[6877]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][23] ;
  assign \new_[6878]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][24] ;
  assign \new_[6879]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][26] ;
  assign \new_[6880]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][27] ;
  assign \new_[6881]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][28] ;
  assign \new_[6882]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][29] ;
  assign \new_[6883]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][30] ;
  assign \new_[6884]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][31] ;
  assign \new_[6885]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][35] ;
  assign \new_[6886]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][3] ;
  assign \new_[6887]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][7] ;
  assign \new_[6888]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][8] ;
  assign \new_[6889]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][9] ;
  assign \new_[6890]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][0] ;
  assign \new_[6891]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][10] ;
  assign \new_[6892]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][13] ;
  assign \new_[6893]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][15] ;
  assign \new_[6894]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][16] ;
  assign \new_[6895]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][17] ;
  assign \new_[6896]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][18] ;
  assign \new_[6897]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][1] ;
  assign \new_[6898]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][20] ;
  assign \new_[6899]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][21] ;
  assign \new_[6900]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][23] ;
  assign \new_[6901]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][24] ;
  assign \new_[6902]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][26] ;
  assign \new_[6903]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][27] ;
  assign \new_[6904]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][28] ;
  assign \new_[6905]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][29] ;
  assign \new_[6906]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][30] ;
  assign \new_[6907]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][31] ;
  assign \new_[6908]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][35] ;
  assign \new_[6909]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][3] ;
  assign \new_[6910]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][7] ;
  assign \new_[6911]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][8] ;
  assign \new_[6912]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][9] ;
  assign \new_[6913]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][0] ;
  assign \new_[6914]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][10] ;
  assign \new_[6915]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][11] ;
  assign \new_[6916]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][13] ;
  assign \new_[6917]_  = output_backup_mas_ad_en_out_reg;
  assign \new_[6918]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][15] ;
  assign \new_[6919]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][16] ;
  assign \new_[6920]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][17] ;
  assign \new_[6921]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][19] ;
  assign \new_[6922]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][1] ;
  assign \new_[6923]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][20] ;
  assign \new_[6924]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][23] ;
  assign \new_[6925]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][24] ;
  assign \new_[6926]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][26] ;
  assign \new_[6927]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][27] ;
  assign \new_[6928]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][28] ;
  assign \new_[6929]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][30] ;
  assign \new_[6930]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][31] ;
  assign \new_[6931]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][35] ;
  assign \new_[6932]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][3] ;
  assign \new_[6933]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][7] ;
  assign \new_[6934]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][8] ;
  assign \new_[6935]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][9] ;
  assign \new_[6936]_  = ~output_backup_tar_ad_en_out_reg;
  assign n3160 = ~\new_[9847]_  | (~\new_[9846]_  & ~\new_[8241]_ );
  assign n3155 = ~\new_[8150]_  | ~\new_[15279]_ ;
  assign \new_[6939]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][10] ;
  assign \new_[6940]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][19] ;
  assign \new_[6941]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][11] ;
  assign \new_[6942]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][29] ;
  assign \new_[6943]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][21] ;
  assign \new_[6944]_  = ~\new_[7283]_ ;
  assign \new_[6945]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][19] ;
  assign \new_[6946]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][11] ;
  assign \new_[6947]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][28] ;
  assign \new_[6948]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][29] ;
  assign \new_[6949]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][21] ;
  assign \new_[6950]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][17] ;
  assign \new_[6951]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][19] ;
  assign \new_[6952]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][0] ;
  assign \new_[6953]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][29] ;
  assign \new_[6954]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][3] ;
  assign \new_[6955]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][28] ;
  assign \new_[6956]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][27] ;
  assign \new_[6957]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][10] ;
  assign \new_[6958]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][18] ;
  assign \new_[6959]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][1] ;
  assign \new_[6960]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][3] ;
  assign \new_[6961]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][21] ;
  assign \new_[6962]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][29] ;
  assign \new_[6963]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][35] ;
  assign \new_[6964]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][18] ;
  assign \new_[6965]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][10] ;
  assign \new_[6966]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][35] ;
  assign \new_[6967]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][10] ;
  assign \new_[6968]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][19] ;
  assign \new_[6969]_  = ~\new_[9137]_  | ~\new_[8572]_  | ~\new_[8573]_  | ~\new_[9136]_ ;
  assign \new_[6970]_  = ~\new_[9140]_  | ~\new_[8576]_  | ~\new_[8117]_  | ~\new_[9139]_ ;
  assign \new_[6971]_  = ~\new_[8120]_  | ~\new_[9143]_  | ~\new_[8579]_  | ~\new_[9142]_ ;
  assign \new_[6972]_  = ~\new_[8583]_  | ~\new_[9145]_  | ~\new_[8584]_  | ~\new_[9144]_ ;
  assign \new_[6973]_  = ~\new_[9147]_  | ~\new_[8589]_  | ~\new_[8126]_  | ~\new_[9146]_ ;
  assign \new_[6974]_  = ~\new_[8593]_  | ~\new_[9149]_  | ~\new_[9148]_  | ~\new_[8592]_ ;
  assign \new_[6975]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][29] ;
  assign \new_[6976]_  = ~\new_[8597]_  | ~\new_[9151]_  | ~\new_[9150]_  | ~\new_[8596]_ ;
  assign \new_[6977]_  = ~\new_[9153]_  | ~\new_[8602]_  | ~\new_[8601]_  | ~\new_[9152]_ ;
  assign \new_[6978]_  = ~\new_[9155]_  | ~\new_[8607]_  | ~\new_[9154]_  | ~\new_[8606]_ ;
  assign \new_[6979]_  = ~\new_[9158]_  | ~\new_[8614]_  | ~\new_[8612]_  | ~\new_[9159]_ ;
  assign \new_[6980]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][3] ;
  assign \new_[6981]_  = ~\new_[9161]_  | ~\new_[8618]_  | ~\new_[8617]_  | ~\new_[9160]_ ;
  assign \new_[6982]_  = ~\new_[9162]_  | ~\new_[8620]_  | ~\new_[8139]_  | ~\new_[9163]_ ;
  assign \new_[6983]_  = ~\new_[9166]_  | ~\new_[9167]_  | ~\new_[8145]_  | ~\new_[8629]_ ;
  assign \new_[6984]_  = ~\new_[8630]_  | ~\new_[9169]_  | ~\new_[8147]_  | ~\new_[9168]_ ;
  assign \new_[6985]_  = ~\new_[8632]_  | ~\new_[8633]_  | ~\new_[9170]_  | ~\new_[9171]_ ;
  assign \pci_ad_oe_o[30]  = pci_io_mux_ad_iob30_en_out_reg;
  assign \new_[6987]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][29] ;
  assign \pci_ad_oe_o[0]  = pci_io_mux_ad_iob0_en_out_reg;
  assign \new_[6989]_  = ~\new_[9176]_  | ~\new_[8640]_  | ~\new_[8639]_  | ~\new_[9177]_ ;
  assign \new_[6990]_  = ~\new_[9179]_  | ~\new_[8641]_  | ~\new_[9178]_  | ~\new_[8337]_ ;
  assign \new_[6991]_  = ~\new_[8645]_  | ~\new_[9181]_  | ~\new_[8644]_  | ~\new_[9180]_ ;
  assign \new_[6992]_  = ~\new_[9182]_  | ~\new_[9183]_  | ~\new_[8648]_  | ~\new_[8647]_ ;
  assign \new_[6993]_  = ~\new_[8347]_  | ~\new_[8655]_  | ~\new_[9186]_  | ~\new_[8654]_ ;
  assign \new_[6994]_  = ~\new_[8657]_  | ~\new_[8351]_  | ~\new_[8656]_  | ~\new_[8350]_ ;
  assign \pci_ad_oe_o[6]  = pci_io_mux_ad_iob6_en_out_reg;
  assign \new_[6996]_  = ~\new_[8353]_  | ~\new_[8659]_  | ~\new_[8352]_  | ~\new_[8658]_ ;
  assign \new_[6997]_  = ~\new_[8355]_  | ~\new_[8660]_  | ~\new_[8356]_  | ~\new_[8661]_ ;
  assign \new_[6998]_  = ~\new_[8663]_  | ~\new_[8662]_  | ~\new_[8358]_  | ~\new_[8357]_ ;
  assign \new_[6999]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][18] ;
  assign \pci_ad_oe_o[12]  = pci_io_mux_ad_iob12_en_out_reg;
  assign \new_[7001]_  = ~\new_[8664]_  | ~\new_[8361]_  | ~\new_[8360]_  | ~\new_[8665]_ ;
  assign \pci_ad_oe_o[10]  = pci_io_mux_ad_iob10_en_out_reg;
  assign \new_[7003]_  = ~\new_[8667]_  | ~\new_[8364]_  | ~\new_[8666]_  | ~\new_[8363]_ ;
  assign \new_[7004]_  = ~\new_[8668]_  | ~\new_[8669]_  | ~\new_[8367]_  | ~\new_[8366]_ ;
  assign \new_[7005]_  = ~\new_[8671]_  | ~\new_[8369]_  | ~\new_[8670]_  | ~\new_[8186]_ ;
  assign \new_[7006]_  = ~\new_[8372]_  | ~\new_[8673]_  | ~\new_[8371]_  | ~\new_[8672]_ ;
  assign \pci_ad_oe_o[16]  = pci_io_mux_ad_iob16_en_out_reg;
  assign \new_[7008]_  = ~\new_[8674]_  | ~\new_[8375]_  | ~\new_[8374]_  | ~\new_[8675]_ ;
  assign \new_[7009]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][10] ;
  assign \new_[7010]_  = ~\new_[8676]_  | ~\new_[8379]_  | ~\new_[8378]_  | ~\new_[8677]_ ;
  assign \new_[7011]_  = ~\new_[8382]_  | ~\new_[8383]_  | ~\new_[8678]_  | ~\new_[8679]_ ;
  assign \new_[7012]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][3] ;
  assign \pci_ad_oe_o[20]  = pci_io_mux_ad_iob20_en_out_reg;
  assign \pci_ad_oe_o[24]  = pci_io_mux_ad_iob24_en_out_reg;
  assign \new_[7015]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][18] ;
  assign \new_[7016]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][10] ;
  assign \new_[7017]_  = ~\new_[19877]_  | ~\new_[18165]_ ;
  assign \new_[7018]_  = ~\new_[19877]_  | ~\new_[18226]_ ;
  assign \new_[7019]_  = ~\new_[19877]_  | ~\new_[18180]_ ;
  assign \new_[7020]_  = ~\new_[19877]_  | ~\new_[19541]_ ;
  assign \new_[7021]_  = ~\new_[19877]_  | ~\new_[17883]_ ;
  assign \new_[7022]_  = ~\new_[19876]_  | ~\new_[18236]_ ;
  assign \new_[7023]_  = ~\new_[19877]_  | ~\new_[18754]_ ;
  assign \new_[7024]_  = ~\new_[19877]_  | ~\new_[19690]_ ;
  assign \new_[7025]_  = ~\new_[19877]_  | ~\new_[18246]_ ;
  assign \new_[7026]_  = ~\new_[19877]_  | ~\new_[18864]_ ;
  assign \new_[7027]_  = ~\new_[19876]_  | ~\new_[17874]_ ;
  assign \new_[7028]_  = ~\new_[19876]_  | ~\new_[18139]_ ;
  assign \new_[7029]_  = ~\new_[19877]_  | ~\new_[19413]_ ;
  assign \new_[7030]_  = ~\new_[8092]_  | ~\new_[18217]_ ;
  assign \new_[7031]_  = ~\new_[8103]_  | ~\new_[18519]_ ;
  assign \new_[7032]_  = ~\new_[8092]_  | ~\new_[18882]_ ;
  assign \new_[7033]_  = ~\new_[8092]_  | ~\new_[18468]_ ;
  assign \new_[7034]_  = ~\new_[8103]_  | ~\new_[17808]_ ;
  assign \new_[7035]_  = ~\new_[8092]_  | ~\new_[17938]_ ;
  assign \new_[7036]_  = ~\new_[8103]_  | ~\new_[19488]_ ;
  assign \new_[7037]_  = ~\new_[8087]_  | ~\new_[18795]_ ;
  assign \new_[7038]_  = ~\new_[8087]_  | ~\new_[18698]_ ;
  assign \new_[7039]_  = ~\new_[8092]_  | ~\new_[19502]_ ;
  assign \new_[7040]_  = ~\new_[8092]_  | ~\new_[18865]_ ;
  assign \new_[7041]_  = ~\new_[8103]_  | ~\new_[18531]_ ;
  assign \new_[7042]_  = ~\new_[8092]_  | ~\new_[18812]_ ;
  assign \new_[7043]_  = ~\new_[8092]_  | ~\new_[19307]_ ;
  assign \new_[7044]_  = ~\new_[8092]_  | ~\new_[18768]_ ;
  assign \new_[7045]_  = ~\new_[8087]_  | ~\new_[18740]_ ;
  assign \new_[7046]_  = ~\new_[8092]_  | ~\new_[18714]_ ;
  assign \new_[7047]_  = ~\new_[8087]_  | ~\new_[18836]_ ;
  assign \new_[7048]_  = ~\new_[8092]_  | ~\new_[18780]_ ;
  assign \new_[7049]_  = ~\new_[8103]_  | ~\new_[19485]_ ;
  assign \new_[7050]_  = ~\new_[8087]_  | ~\new_[18118]_ ;
  assign \new_[7051]_  = ~\new_[8092]_  | ~\new_[17940]_ ;
  assign \new_[7052]_  = ~\new_[8103]_  | ~\new_[17845]_ ;
  assign \new_[7053]_  = ~\new_[8087]_  | ~\new_[19461]_ ;
  assign \new_[7054]_  = ~\new_[8092]_  | ~\new_[19500]_ ;
  assign \new_[7055]_  = ~\new_[8092]_  | ~\new_[17941]_ ;
  assign \new_[7056]_  = ~\new_[8092]_  | ~\new_[19142]_ ;
  assign \new_[7057]_  = ~\new_[8087]_  | ~\new_[18558]_ ;
  assign \new_[7058]_  = ~\new_[8087]_  | ~\new_[19329]_ ;
  assign \new_[7059]_  = ~\new_[8091]_  & ~\new_[11430]_ ;
  assign \new_[7060]_  = ~\new_[8087]_  | ~\new_[19330]_ ;
  assign \new_[7061]_  = ~\new_[8092]_  | ~\new_[18902]_ ;
  assign \new_[7062]_  = ~\new_[8092]_  | ~\new_[18591]_ ;
  assign \new_[7063]_  = ~\new_[8092]_  | ~\new_[18345]_ ;
  assign \new_[7064]_  = ~\new_[8087]_  | ~\new_[18000]_ ;
  assign \new_[7065]_  = ~\new_[8092]_  | ~\new_[18525]_ ;
  assign \new_[7066]_  = ~\new_[8087]_  | ~\new_[18656]_ ;
  assign \new_[7067]_  = ~\new_[8092]_  | ~\new_[19504]_ ;
  assign \new_[7068]_  = ~\new_[8092]_  | ~\new_[18566]_ ;
  assign \new_[7069]_  = ~\new_[8092]_  | ~\new_[19303]_ ;
  assign \new_[7070]_  = ~\new_[8092]_  | ~\new_[18281]_ ;
  assign \new_[7071]_  = ~\new_[8103]_  | ~\new_[17966]_ ;
  assign \new_[7072]_  = ~\new_[8103]_  | ~\new_[18632]_ ;
  assign \new_[7073]_  = ~\new_[8092]_  | ~\new_[19304]_ ;
  assign \new_[7074]_  = ~\new_[8087]_  | ~\new_[18114]_ ;
  assign \new_[7075]_  = ~\new_[8093]_  | ~\new_[19478]_ ;
  assign \new_[7076]_  = ~\new_[8107]_  | ~\new_[18679]_ ;
  assign \new_[7077]_  = ~\new_[8111]_  | ~\new_[17881]_ ;
  assign \new_[7078]_  = ~\new_[8100]_  | ~\new_[18683]_ ;
  assign \new_[7079]_  = ~\new_[8113]_  | ~\new_[17849]_ ;
  assign \new_[7080]_  = ~\new_[8101]_  | ~\new_[18489]_ ;
  assign \new_[7081]_  = ~\new_[8084]_  | ~\new_[19147]_ ;
  assign \new_[7082]_  = ~\new_[8083]_  | ~\new_[19367]_ ;
  assign \new_[7083]_  = ~\new_[8100]_  | ~\new_[18207]_ ;
  assign \new_[7084]_  = ~\new_[8094]_  | ~\new_[18937]_ ;
  assign \new_[7085]_  = ~\new_[8082]_  | ~\new_[18751]_ ;
  assign \new_[7086]_  = ~\new_[8094]_  | ~\new_[18282]_ ;
  assign \new_[7087]_  = ~\new_[8109]_  & ~\new_[11390]_ ;
  assign \new_[7088]_  = ~\new_[8101]_  | ~\new_[18291]_ ;
  assign \new_[7089]_  = ~\new_[8100]_  | ~\new_[19262]_ ;
  assign \new_[7090]_  = ~\new_[8083]_  | ~\new_[19632]_ ;
  assign \new_[7091]_  = ~\new_[8094]_  | ~\new_[19476]_ ;
  assign \new_[7092]_  = ~\new_[8110]_  | ~\new_[18611]_ ;
  assign \new_[7093]_  = ~\new_[8096]_  | ~\new_[18564]_ ;
  assign \new_[7094]_  = ~\new_[8108]_  | ~\new_[18650]_ ;
  assign \new_[7095]_  = ~\new_[8093]_  | ~\new_[19119]_ ;
  assign \new_[7096]_  = ~\new_[8100]_  | ~\new_[18663]_ ;
  assign \new_[7097]_  = ~\new_[8111]_  | ~\new_[19146]_ ;
  assign \new_[7098]_  = ~\new_[8113]_  | ~\new_[18012]_ ;
  assign \new_[7099]_  = ~\new_[8101]_  | ~\new_[18305]_ ;
  assign \new_[7100]_  = ~\new_[8084]_  | ~\new_[19150]_ ;
  assign \new_[7101]_  = ~\new_[8082]_  | ~\new_[19072]_ ;
  assign \new_[7102]_  = ~\new_[8113]_  | ~\new_[18129]_ ;
  assign \new_[7103]_  = ~\new_[8101]_  | ~\new_[19315]_ ;
  assign \new_[7104]_  = ~\new_[8107]_  | ~\new_[18446]_ ;
  assign \new_[7105]_  = ~\new_[8101]_  | ~\new_[18327]_ ;
  assign \new_[7106]_  = ~\new_[8082]_  | ~\new_[19548]_ ;
  assign \new_[7107]_  = ~\new_[8111]_  | ~\new_[18042]_ ;
  assign \new_[7108]_  = ~\new_[8100]_  | ~\new_[18240]_ ;
  assign \new_[7109]_  = ~\new_[8107]_  | ~\new_[19350]_ ;
  assign \new_[7110]_  = ~\new_[8093]_  | ~\new_[19681]_ ;
  assign \new_[7111]_  = ~\new_[8105]_  | ~\new_[19225]_ ;
  assign \new_[7112]_  = ~\new_[8107]_  | ~\new_[17905]_ ;
  assign \new_[7113]_  = ~\new_[8085]_  | ~\new_[18737]_ ;
  assign \new_[7114]_  = ~\new_[8098]_  | ~\new_[17847]_ ;
  assign \new_[7115]_  = ~\new_[8094]_  | ~\new_[18355]_ ;
  assign \new_[7116]_  = ~\new_[8107]_  | ~\new_[18613]_ ;
  assign \new_[7117]_  = ~\new_[8096]_  | ~\new_[19675]_ ;
  assign \new_[7118]_  = ~\new_[8112]_  & ~\new_[11446]_ ;
  assign \new_[7119]_  = ~\new_[8110]_  | ~\new_[18887]_ ;
  assign \new_[7120]_  = ~\new_[8094]_  | ~\new_[19474]_ ;
  assign \new_[7121]_  = ~\new_[8111]_  | ~\new_[18044]_ ;
  assign \new_[7122]_  = ~\new_[8105]_  | ~\new_[19637]_ ;
  assign \new_[7123]_  = ~\new_[8093]_  | ~\new_[17931]_ ;
  assign \new_[7124]_  = ~\new_[8107]_  | ~\new_[17906]_ ;
  assign \new_[7125]_  = ~\new_[8086]_  | ~\new_[19778]_ ;
  assign \new_[7126]_  = ~\new_[8099]_  | ~\new_[18333]_ ;
  assign \new_[7127]_  = ~\new_[8100]_  | ~\new_[18556]_ ;
  assign \new_[7128]_  = ~\new_[8082]_  | ~\new_[19207]_ ;
  assign \new_[7129]_  = ~\new_[8098]_  | ~\new_[18991]_ ;
  assign \new_[7130]_  = ~\new_[8110]_  | ~\new_[19283]_ ;
  assign \new_[7131]_  = ~\new_[8094]_  | ~\new_[18304]_ ;
  assign \new_[7132]_  = ~\new_[8099]_  | ~\new_[18919]_ ;
  assign \new_[7133]_  = ~\new_[8086]_  | ~\new_[19122]_ ;
  assign \new_[7134]_  = ~\new_[8094]_  | ~\new_[19473]_ ;
  assign \new_[7135]_  = ~\new_[8107]_  | ~\new_[19526]_ ;
  assign \new_[7136]_  = ~\new_[8096]_  | ~\new_[17937]_ ;
  assign \new_[7137]_  = ~\new_[8111]_  | ~\new_[18050]_ ;
  assign \new_[7138]_  = ~\new_[8108]_  | ~\new_[19527]_ ;
  assign \new_[7139]_  = ~\new_[8094]_  | ~\new_[19131]_ ;
  assign \new_[7140]_  = ~\new_[8083]_  | ~\new_[18805]_ ;
  assign \new_[7141]_  = ~\new_[8111]_  | ~\new_[18060]_ ;
  assign \new_[7142]_  = ~\new_[8100]_  | ~\new_[19316]_ ;
  assign \new_[7143]_  = ~\new_[8107]_  | ~\new_[19515]_ ;
  assign \new_[7144]_  = ~\new_[8094]_  | ~\new_[19471]_ ;
  assign \new_[7145]_  = ~\new_[8093]_  | ~\new_[19472]_ ;
  assign \new_[7146]_  = ~\new_[8096]_  | ~\new_[19068]_ ;
  assign \new_[7147]_  = ~\new_[8107]_  | ~\new_[19522]_ ;
  assign \new_[7148]_  = ~\new_[8086]_  | ~\new_[18374]_ ;
  assign \new_[7149]_  = ~\new_[8099]_  | ~\new_[18605]_ ;
  assign \new_[7150]_  = ~\new_[8101]_  | ~\new_[18361]_ ;
  assign \new_[7151]_  = ~\new_[8112]_  & ~\new_[11793]_ ;
  assign \new_[7152]_  = ~\new_[8082]_  | ~\new_[19190]_ ;
  assign \new_[7153]_  = ~\new_[8098]_  | ~\new_[18629]_ ;
  assign \new_[7154]_  = ~\new_[8111]_  | ~\new_[18832]_ ;
  assign \new_[7155]_  = ~\new_[8105]_  | ~\new_[18265]_ ;
  assign \new_[7156]_  = ~\new_[8094]_  | ~\new_[18268]_ ;
  assign \new_[7157]_  = ~\new_[8096]_  | ~\new_[18616]_ ;
  assign \new_[7158]_  = ~\new_[8110]_  | ~\new_[19506]_ ;
  assign \new_[7159]_  = ~\new_[8105]_  | ~\new_[19671]_ ;
  assign \new_[7160]_  = ~\new_[8093]_  | ~\new_[17951]_ ;
  assign \new_[7161]_  = ~\new_[8108]_  | ~\new_[17908]_ ;
  assign \new_[7162]_  = ~\new_[8084]_  | ~\new_[17921]_ ;
  assign \new_[7163]_  = ~\new_[8093]_  | ~\new_[17948]_ ;
  assign \new_[7164]_  = ~\new_[8107]_  | ~\new_[19525]_ ;
  assign \new_[7165]_  = ~\new_[8084]_  | ~\new_[17907]_ ;
  assign \new_[7166]_  = ~\new_[8110]_  | ~\new_[19713]_ ;
  assign \new_[7167]_  = ~\new_[8094]_  | ~\new_[19310]_ ;
  assign \new_[7168]_  = ~\new_[8113]_  | ~\new_[18142]_ ;
  assign \new_[7169]_  = ~\new_[8101]_  | ~\new_[19439]_ ;
  assign \new_[7170]_  = ~\new_[8085]_  | ~\new_[18535]_ ;
  assign \new_[7171]_  = ~\new_[8098]_  | ~\new_[18091]_ ;
  assign \new_[7172]_  = ~\new_[8100]_  | ~\new_[19565]_ ;
  assign \new_[7173]_  = ~\new_[8113]_  | ~\new_[19228]_ ;
  assign \new_[7174]_  = ~\new_[8085]_  | ~\new_[18170]_ ;
  assign \new_[7175]_  = ~\new_[8105]_  | ~\new_[18395]_ ;
  assign \new_[7176]_  = ~\new_[8094]_  | ~\new_[19491]_ ;
  assign \new_[7177]_  = ~\new_[8101]_  | ~\new_[19532]_ ;
  assign \new_[7178]_  = ~\new_[8100]_  | ~\new_[17835]_ ;
  assign \new_[7179]_  = ~\new_[8085]_  | ~\new_[19365]_ ;
  assign \new_[7180]_  = ~\new_[8105]_  | ~\new_[19004]_ ;
  assign \new_[7181]_  = ~\new_[8094]_  | ~\new_[19520]_ ;
  assign \new_[7182]_  = ~\new_[8107]_  | ~\new_[19523]_ ;
  assign \new_[7183]_  = ~\new_[8093]_  | ~\new_[18674]_ ;
  assign \new_[7184]_  = ~\new_[8107]_  | ~\new_[19524]_ ;
  assign \new_[7185]_  = ~\new_[8085]_  | ~\new_[18340]_ ;
  assign \new_[7186]_  = ~\new_[8098]_  | ~\new_[18450]_ ;
  assign \new_[7187]_  = ~\new_[8105]_  | ~\new_[17963]_ ;
  assign \new_[7188]_  = ~\new_[8093]_  | ~\new_[18241]_ ;
  assign \new_[7189]_  = ~\new_[8108]_  | ~\new_[19133]_ ;
  assign \new_[7190]_  = ~\new_[8098]_  | ~\new_[17809]_ ;
  assign \new_[7191]_  = ~\new_[8085]_  | ~\new_[18933]_ ;
  assign \new_[7192]_  = ~\new_[8108]_  | ~\new_[17917]_ ;
  assign \new_[7193]_  = ~\new_[8094]_  | ~\new_[19469]_ ;
  assign \new_[7194]_  = ~\new_[8098]_  | ~\new_[18068]_ ;
  assign \new_[7195]_  = ~\new_[8083]_  | ~\new_[18746]_ ;
  assign \new_[7196]_  = ~\new_[8094]_  | ~\new_[19319]_ ;
  assign \new_[7197]_  = ~\new_[8107]_  | ~\new_[18363]_ ;
  assign \new_[7198]_  = ~\new_[8111]_  | ~\new_[19324]_ ;
  assign \new_[7199]_  = ~\new_[8100]_  | ~\new_[18653]_ ;
  assign \new_[7200]_  = ~\new_[8113]_  | ~\new_[18895]_ ;
  assign \new_[7201]_  = ~\new_[8101]_  | ~\new_[18259]_ ;
  assign \new_[7202]_  = ~\new_[8101]_  | ~\new_[18276]_ ;
  assign \new_[7203]_  = ~\new_[8100]_  | ~\new_[18533]_ ;
  assign \new_[7204]_  = ~\new_[8082]_  | ~\new_[18943]_ ;
  assign \new_[7205]_  = ~\new_[8094]_  | ~\new_[18958]_ ;
  assign \new_[7206]_  = ~\new_[8101]_  | ~\new_[18719]_ ;
  assign \new_[7207]_  = ~\new_[8082]_  | ~\new_[19786]_ ;
  assign \new_[7208]_  = ~\new_[8111]_  | ~\new_[19571]_ ;
  assign \new_[7209]_  = ~\new_[8100]_  | ~\new_[18830]_ ;
  assign \new_[7210]_  = ~\new_[8094]_  | ~\new_[18659]_ ;
  assign \new_[7211]_  = ~\new_[8105]_  | ~\new_[19499]_ ;
  assign \new_[7212]_  = ~\new_[8093]_  | ~\new_[19479]_ ;
  assign \new_[7213]_  = ~\new_[8108]_  | ~\new_[18763]_ ;
  assign \new_[7214]_  = ~\new_[8086]_  | ~\new_[18407]_ ;
  assign \new_[7215]_  = ~\new_[8099]_  | ~\new_[17987]_ ;
  assign \new_[7216]_  = ~\new_[8093]_  | ~\new_[19480]_ ;
  assign \new_[7217]_  = ~\new_[8107]_  | ~\new_[18704]_ ;
  assign \new_[7218]_  = ~\new_[8084]_  | ~\new_[17885]_ ;
  assign \new_[7219]_  = ~\new_[8093]_  | ~\new_[18744]_ ;
  assign \new_[7220]_  = ~\new_[8108]_  | ~\new_[18755]_ ;
  assign \new_[7221]_  = ~\new_[8086]_  | ~\new_[19269]_ ;
  assign \new_[7222]_  = ~\new_[8112]_  & ~\new_[11724]_ ;
  assign \new_[7223]_  = ~\new_[8093]_  | ~\new_[18782]_ ;
  assign \new_[7224]_  = ~\new_[8107]_  | ~\new_[18371]_ ;
  assign \new_[7225]_  = ~\new_[8083]_  | ~\new_[18801]_ ;
  assign \new_[7226]_  = ~\new_[8105]_  | ~\new_[18742]_ ;
  assign \new_[7227]_  = ~\new_[8094]_  | ~\new_[19475]_ ;
  assign \new_[7228]_  = ~\new_[8109]_  & ~\new_[11308]_ ;
  assign \new_[7229]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][20] ;
  assign \new_[7230]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][0] ;
  assign \new_[7231]_  = ~\new_[7368]_ ;
  assign \new_[7232]_  = ~\new_[7395]_ ;
  assign \new_[7233]_  = ~\new_[7398]_ ;
  assign \new_[7234]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][1] ;
  assign \new_[7235]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][16] ;
  assign \new_[7236]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][9] ;
  assign \new_[7237]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][29] ;
  assign \new_[7238]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][21] ;
  assign \new_[7239]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][18] ;
  assign \new_[7240]_  = ~\new_[7419]_ ;
  assign \new_[7241]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][33] ;
  assign \new_[7242]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][32] ;
  assign \new_[7243]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][33] ;
  assign \new_[7244]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][33] ;
  assign \new_[7245]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][32] ;
  assign \new_[7246]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][32] ;
  assign \new_[7247]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][33] ;
  assign \new_[7248]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][32] ;
  assign \new_[7249]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][32] ;
  assign \new_[7250]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][33] ;
  assign \new_[7251]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][33] ;
  assign \new_[7252]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][32] ;
  assign \new_[7253]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][32] ;
  assign \new_[7254]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][32] ;
  assign \new_[7255]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][32] ;
  assign \new_[7256]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][32] ;
  assign \new_[7257]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][32] ;
  assign \new_[7258]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][32] ;
  assign \new_[7259]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][33] ;
  assign \new_[7260]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][32] ;
  assign \new_[7261]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][33] ;
  assign \new_[7262]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][32] ;
  assign \new_[7263]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][33] ;
  assign \new_[7264]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][32] ;
  assign \new_[7265]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][32] ;
  assign \new_[7266]_  = pci_target_unit_wishbone_master_first_data_is_burst_reg_reg;
  assign n3165 = \wbs_adr_i[11]  ? \new_[15279]_  : \new_[8551]_ ;
  assign n3170 = \wbs_adr_i[10]  ? \new_[15279]_  : \new_[8550]_ ;
  assign n3235 = \wbs_adr_i[12]  ? \new_[15279]_  : \new_[8552]_ ;
  assign n3175 = \wbs_adr_i[13]  ? \new_[15279]_  : \new_[8553]_ ;
  assign n3185 = \wbs_adr_i[15]  ? \new_[15279]_  : \new_[8555]_ ;
  assign n3180 = \wbs_adr_i[14]  ? \new_[15279]_  : \new_[8554]_ ;
  assign n3190 = \wbs_adr_i[16]  ? \new_[15279]_  : \new_[8558]_ ;
  assign n3195 = \wbs_adr_i[17]  ? \new_[15279]_  : \new_[8561]_ ;
  assign \new_[7275]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][33] ;
  assign n3295 = \wbs_adr_i[18]  ? \new_[15279]_  : \new_[8564]_ ;
  assign n3200 = \wbs_adr_i[19]  ? \new_[15279]_  : \new_[8568]_ ;
  assign n3205 = \wbs_adr_i[20]  ? \new_[15279]_  : \new_[8570]_ ;
  assign n3210 = \wbs_adr_i[21]  ? \new_[15279]_  : \new_[8574]_ ;
  assign n3290 = \wbs_adr_i[22]  ? \new_[15279]_  : \new_[8575]_ ;
  assign \new_[7281]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][33] ;
  assign n3215 = \wbs_adr_i[23]  ? \new_[15279]_  : \new_[8578]_ ;
  assign \new_[7283]_  = ~\new_[20026]_ ;
  assign n3220 = \wbs_adr_i[24]  ? \new_[15279]_  : \new_[8582]_ ;
  assign n3225 = \wbs_adr_i[25]  ? \new_[15279]_  : \new_[8585]_ ;
  assign n3305 = \wbs_adr_i[26]  ? \new_[15279]_  : \new_[8588]_ ;
  assign n3230 = \wbs_adr_i[27]  ? \new_[15279]_  : \new_[8591]_ ;
  assign \new_[7288]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][33] ;
  assign n3280 = \wbs_adr_i[28]  ? \new_[15279]_  : \new_[8594]_ ;
  assign n3315 = \wbs_adr_i[2]  ? \new_[15279]_  : \new_[8627]_ ;
  assign n3245 = \wbs_adr_i[30]  ? \new_[15279]_  : \new_[8600]_ ;
  assign n3240 = \wbs_adr_i[29]  ? \new_[15279]_  : \new_[8598]_ ;
  assign \new_[7293]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][33] ;
  assign n3250 = \wbs_adr_i[31]  ? \new_[15279]_  : \new_[8605]_ ;
  assign n3255 = \wbs_adr_i[3]  ? \new_[15279]_  : \new_[8608]_ ;
  assign n3310 = \wbs_adr_i[4]  ? \new_[15279]_  : \new_[8611]_ ;
  assign n3260 = \wbs_adr_i[5]  ? \new_[15279]_  : \new_[8613]_ ;
  assign n3265 = \wbs_adr_i[6]  ? \new_[15279]_  : \new_[8616]_ ;
  assign n3270 = \wbs_adr_i[7]  ? \new_[15279]_  : \new_[8619]_ ;
  assign n3275 = \wbs_adr_i[9]  ? \new_[15279]_  : \new_[8624]_ ;
  assign n3300 = \wbs_adr_i[8]  ? \new_[15279]_  : \new_[8621]_ ;
  assign \new_[7302]_  = ~\new_[9164]_  | ~\new_[9165]_  | ~\new_[8623]_  | ~\new_[8625]_ ;
  assign \new_[7303]_  = ~\new_[9172]_  | ~\new_[9173]_  | ~\new_[8635]_  | ~\new_[8636]_ ;
  assign \new_[7304]_  = ~\new_[9184]_  | ~\new_[9185]_  | ~\new_[8651]_  | ~\new_[8652]_ ;
  assign n3285 = ~\new_[8263]_  | (~\new_[14967]_  & ~\new_[17510]_ );
  assign \new_[7306]_  = ~\new_[8279]_  | ~\new_[18766]_ ;
  assign \new_[7307]_  = ~\new_[8284]_  | ~\new_[18772]_ ;
  assign \new_[7308]_  = ~\new_[8279]_  | ~\new_[18196]_ ;
  assign \new_[7309]_  = ~\new_[8279]_  | ~\new_[18538]_ ;
  assign \new_[7310]_  = ~\new_[8279]_  | ~\new_[17986]_ ;
  assign \new_[7311]_  = ~\new_[8284]_  | ~\new_[18645]_ ;
  assign \new_[7312]_  = ~\new_[8279]_  | ~\new_[19746]_ ;
  assign \new_[7313]_  = ~\new_[8279]_  | ~\new_[17857]_ ;
  assign \new_[7314]_  = ~\new_[8277]_  | ~\new_[17859]_ ;
  assign \new_[7315]_  = ~\new_[8284]_  | ~\new_[18797]_ ;
  assign \new_[7316]_  = ~\new_[8277]_  | ~\new_[19424]_ ;
  assign \new_[7317]_  = ~\new_[8279]_  | ~\new_[18439]_ ;
  assign \new_[7318]_  = ~\new_[8284]_  | ~\new_[19745]_ ;
  assign \new_[7319]_  = ~\new_[8279]_  | ~\new_[19860]_ ;
  assign \new_[7320]_  = ~\new_[8278]_  | ~\new_[19868]_ ;
  assign \new_[7321]_  = ~\new_[8277]_  | ~\new_[18955]_ ;
  assign \new_[7322]_  = ~\new_[8284]_  | ~\new_[19698]_ ;
  assign \new_[7323]_  = ~\new_[8278]_  | ~\new_[19161]_ ;
  assign \new_[7324]_  = ~\new_[8284]_  | ~\new_[18990]_ ;
  assign \new_[7325]_  = ~\new_[8278]_  | ~\new_[19589]_ ;
  assign \new_[7326]_  = ~\new_[8278]_  | ~\new_[18208]_ ;
  assign \new_[7327]_  = ~\new_[8285]_  | ~\new_[18787]_ ;
  assign \new_[7328]_  = ~\new_[8278]_  | ~\new_[19575]_ ;
  assign \new_[7329]_  = ~\new_[8279]_  | ~\new_[19346]_ ;
  assign \new_[7330]_  = ~\new_[8279]_  | ~\new_[19813]_ ;
  assign \new_[7331]_  = ~\new_[8277]_  | ~\new_[19837]_ ;
  assign \new_[7332]_  = ~\new_[8279]_  | ~\new_[18379]_ ;
  assign \new_[7333]_  = ~\new_[8279]_  | ~\new_[18420]_ ;
  assign \new_[7334]_  = ~\new_[8278]_  | ~\new_[19431]_ ;
  assign \new_[7335]_  = ~\new_[8285]_  | ~\new_[18697]_ ;
  assign \new_[7336]_  = ~\new_[8277]_  | ~\new_[17836]_ ;
  assign \new_[7337]_  = ~\new_[8285]_  | ~\new_[18424]_ ;
  assign \new_[7338]_  = ~\new_[8279]_  | ~\new_[17988]_ ;
  assign \new_[7339]_  = ~\new_[8278]_  | ~\new_[19127]_ ;
  assign \new_[7340]_  = ~\new_[8279]_  | ~\new_[17999]_ ;
  assign \new_[7341]_  = ~\new_[8279]_  | ~\new_[19419]_ ;
  assign \new_[7342]_  = ~\new_[8277]_  | ~\new_[19451]_ ;
  assign \new_[7343]_  = ~\new_[8284]_  | ~\new_[17995]_ ;
  assign \new_[7344]_  = ~\new_[8277]_  | ~\new_[19708]_ ;
  assign \new_[7345]_  = ~\new_[8279]_  | ~\new_[18097]_ ;
  assign \new_[7346]_  = ~\new_[8279]_  | ~\new_[19417]_ ;
  assign \new_[7347]_  = ~\new_[8284]_  | ~\new_[18551]_ ;
  assign \new_[7348]_  = ~\new_[8279]_  | ~\new_[19067]_ ;
  assign \new_[7349]_  = (~\new_[9190]_  | ~\new_[18293]_ ) & (~\new_[9239]_  | ~\new_[19678]_ );
  assign \new_[7350]_  = (~\new_[9190]_  | ~\new_[18083]_ ) & (~\new_[9239]_  | ~\new_[18788]_ );
  assign \new_[7351]_  = (~\new_[9190]_  | ~\new_[18061]_ ) & (~\new_[9239]_  | ~\new_[19865]_ );
  assign \new_[7352]_  = (~\new_[20501]_  | ~\new_[19785]_ ) & (~\new_[8388]_  | ~\new_[18110]_ );
  assign \new_[7353]_  = (~\new_[9190]_  | ~\new_[18262]_ ) & (~\new_[9239]_  | ~\new_[18920]_ );
  assign \new_[7354]_  = (~\new_[20504]_  | ~\new_[18202]_ ) & (~\new_[8388]_  | ~\new_[19863]_ );
  assign \new_[7355]_  = (~\new_[20504]_  | ~\new_[17933]_ ) & (~\new_[8388]_  | ~\new_[19784]_ );
  assign \new_[7356]_  = (~\new_[9190]_  | ~\new_[18175]_ ) & (~\new_[9239]_  | ~\new_[18542]_ );
  assign \new_[7357]_  = (~\new_[20504]_  | ~\new_[19759]_ ) & (~\new_[8388]_  | ~\new_[18120]_ );
  assign \new_[7358]_  = (~\new_[9190]_  | ~\new_[18161]_ ) & (~\new_[9239]_  | ~\new_[18944]_ );
  assign \new_[7359]_  = (~\new_[20501]_  | ~\new_[19271]_ ) & (~\new_[8388]_  | ~\new_[19232]_ );
  assign \new_[7360]_  = (~\new_[20504]_  | ~\new_[19538]_ ) & (~\new_[8388]_  | ~\new_[18306]_ );
  assign \new_[7361]_  = (~\new_[20504]_  | ~\new_[18222]_ ) & (~\new_[8388]_  | ~\new_[19577]_ );
  assign \new_[7362]_  = (~\new_[9190]_  | ~\new_[19737]_ ) & (~\new_[9239]_  | ~\new_[19121]_ );
  assign \new_[7363]_  = (~\new_[9190]_  | ~\new_[18908]_ ) & (~\new_[9239]_  | ~\new_[18514]_ );
  assign \new_[7364]_  = (~\new_[20504]_  | ~\new_[18258]_ ) & (~\new_[8388]_  | ~\new_[18166]_ );
  assign \new_[7365]_  = (~\new_[20504]_  | ~\new_[19764]_ ) & (~\new_[8388]_  | ~\new_[19792]_ );
  assign \new_[7366]_  = (~\new_[9190]_  | ~\new_[19820]_ ) & (~\new_[9239]_  | ~\new_[19258]_ );
  assign \new_[7367]_  = (~\new_[20504]_  | ~\new_[17838]_ ) & (~\new_[8388]_  | ~\new_[19246]_ );
  assign \new_[7368]_  = \new_[8088]_ ;
  assign \new_[7369]_  = ~\new_[8088]_ ;
  assign \new_[7370]_  = ~\new_[8088]_ ;
  assign \new_[7371]_  = ~\new_[8088]_ ;
  assign \new_[7372]_  = ~\new_[8089]_ ;
  assign \new_[7373]_  = ~\new_[8090]_ ;
  assign \new_[7374]_  = ~\new_[8090]_ ;
  assign \new_[7375]_  = ~\new_[8090]_ ;
  assign \new_[7376]_  = ~\new_[8091]_ ;
  assign \new_[7377]_  = ~\new_[8095]_ ;
  assign \new_[7378]_  = ~\new_[8095]_ ;
  assign \new_[7379]_  = ~\new_[8095]_ ;
  assign \new_[7380]_  = ~\new_[8095]_ ;
  assign \new_[7381]_  = ~\new_[8097]_ ;
  assign \new_[7382]_  = ~\new_[8098]_ ;
  assign \new_[7383]_  = ~\new_[8099]_ ;
  assign \new_[7384]_  = ~\new_[8099]_ ;
  assign \new_[7385]_  = \new_[8099]_ ;
  assign \new_[7386]_  = ~\new_[8102]_ ;
  assign \new_[7387]_  = ~\new_[8104]_ ;
  assign \new_[7388]_  = ~\new_[8105]_ ;
  assign \new_[7389]_  = ~\new_[8106]_ ;
  assign \new_[7390]_  = ~\new_[8106]_ ;
  assign \new_[7391]_  = ~\new_[8106]_ ;
  assign \new_[7392]_  = ~\new_[8106]_ ;
  assign \new_[7393]_  = ~\new_[8109]_ ;
  assign \new_[7394]_  = ~\new_[8112]_ ;
  assign \new_[7395]_  = ~\new_[8112]_ ;
  assign \new_[7396]_  = ~\new_[8113]_ ;
  assign \new_[7397]_  = ~\new_[8114]_ ;
  assign \new_[7398]_  = ~\new_[8114]_ ;
  assign \new_[7399]_  = ~\new_[8114]_ ;
  assign \new_[7400]_  = ~\new_[8114]_ ;
  assign \new_[7401]_  = ~\new_[8118]_ ;
  assign \new_[7402]_  = ~\new_[8122]_ ;
  assign \new_[7403]_  = ~\new_[8135]_ ;
  assign \new_[7404]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][33] ;
  assign \new_[7405]_  = ~\new_[8143]_ ;
  assign \new_[7406]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][33] ;
  assign \new_[7407]_  = ~\new_[8148]_ ;
  assign \new_[7408]_  = ~\new_[8156]_ ;
  assign \new_[7409]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][33] ;
  assign \new_[7410]_  = (~\new_[9290]_  | ~\new_[18973]_ ) & (~\new_[9509]_  | ~\new_[19834]_ );
  assign \new_[7411]_  = ~\new_[8168]_ ;
  assign \new_[7412]_  = (~\new_[9297]_  | ~\new_[19254]_ ) & (~\new_[9503]_  | ~\new_[19822]_ );
  assign \new_[7413]_  = (~\new_[19986]_  | ~\new_[18540]_ ) & (~\new_[20551]_  | ~\new_[18640]_ );
  assign \new_[7414]_  = ~\new_[8174]_ ;
  assign \new_[7415]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][34] ;
  assign \new_[7416]_  = (~\new_[9297]_  | ~\new_[18081]_ ) & (~\new_[9503]_  | ~\new_[18507]_ );
  assign \new_[7417]_  = ~\new_[8177]_ ;
  assign \new_[7418]_  = (~\new_[9297]_  | ~\new_[18947]_ ) & (~\new_[9206]_  | ~\new_[18339]_ );
  assign \new_[7419]_  = (~\new_[9297]_  | ~\new_[19692]_ ) & (~\new_[9503]_  | ~\new_[19763]_ );
  assign \new_[7420]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][5] ;
  assign \new_[7421]_  = ~\new_[8181]_ ;
  assign \new_[7422]_  = (~\new_[9297]_  | ~\new_[18636]_ ) & (~\new_[9206]_  | ~\new_[18559]_ );
  assign \new_[7423]_  = (~\new_[9297]_  | ~\new_[18245]_ ) & (~\new_[9206]_  | ~\new_[18666]_ );
  assign \new_[7424]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][4] ;
  assign \new_[7425]_  = (~\new_[9297]_  | ~\new_[19181]_ ) & (~\new_[9503]_  | ~\new_[18554]_ );
  assign \new_[7426]_  = ~\new_[8194]_ ;
  assign \new_[7427]_  = (~\new_[9297]_  | ~\new_[18329]_ ) & (~\new_[9206]_  | ~\new_[19391]_ );
  assign \new_[7428]_  = (~\new_[9297]_  | ~\new_[19607]_ ) & (~\new_[9206]_  | ~\new_[19370]_ );
  assign \new_[7429]_  = (~\new_[19986]_  | ~\new_[18881]_ ) & (~\new_[20551]_  | ~\new_[17982]_ );
  assign n3480 = ~\new_[9481]_  | (~\new_[9694]_  & ~\new_[8708]_ );
  assign \new_[7431]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][2] ;
  assign \new_[7432]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][25] ;
  assign \new_[7433]_  = i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg;
  assign \new_[7434]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][14] ;
  assign \new_[7435]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][22] ;
  assign \new_[7436]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][25] ;
  assign \new_[7437]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][4] ;
  assign \new_[7438]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][5] ;
  assign \new_[7439]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][14] ;
  assign \new_[7440]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][22] ;
  assign \new_[7441]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][2] ;
  assign \new_[7442]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][5] ;
  assign \new_[7443]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][4] ;
  assign \new_[7444]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][12] ;
  assign \new_[7445]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][22] ;
  assign \new_[7446]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][2] ;
  assign \new_[7447]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][34] ;
  assign \new_[7448]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][5] ;
  assign \new_[7449]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][12] ;
  assign \new_[7450]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][34] ;
  assign \new_[7451]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][4] ;
  assign \new_[7452]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][6] ;
  assign \new_[7453]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][12] ;
  assign \new_[7454]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][14] ;
  assign \new_[7455]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][4] ;
  assign \new_[7456]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][5] ;
  assign \new_[7457]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][22] ;
  assign \new_[7458]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][25] ;
  assign \new_[7459]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][4] ;
  assign \new_[7460]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][5] ;
  assign \new_[7461]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][12] ;
  assign \new_[7462]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][14] ;
  assign \new_[7463]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][22] ;
  assign \new_[7464]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][2] ;
  assign \new_[7465]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][4] ;
  assign \new_[7466]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][6] ;
  assign \new_[7467]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][5] ;
  assign \new_[7468]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][12] ;
  assign \new_[7469]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][22] ;
  assign \new_[7470]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][2] ;
  assign \new_[7471]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][4] ;
  assign \new_[7472]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][5] ;
  assign \new_[7473]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][12] ;
  assign \new_[7474]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][5] ;
  assign \new_[7475]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][12] ;
  assign \new_[7476]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][22] ;
  assign \new_[7477]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][2] ;
  assign \new_[7478]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][4] ;
  assign \new_[7479]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][5] ;
  assign \new_[7480]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][12] ;
  assign \new_[7481]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][22] ;
  assign \new_[7482]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][2] ;
  assign \new_[7483]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][4] ;
  assign \new_[7484]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][5] ;
  assign n3455 = ~\new_[9479]_  | (~\new_[9694]_  & ~\new_[8703]_ );
  assign \new_[7486]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][12] ;
  assign n3460 = ~\new_[9480]_  | (~\new_[9694]_  & ~\new_[8704]_ );
  assign \new_[7488]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][5] ;
  assign \new_[7489]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][12] ;
  assign n3465 = ~\new_[9532]_  | (~\new_[9694]_  & ~\new_[8705]_ );
  assign \new_[7491]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][34] ;
  assign \new_[7492]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][6] ;
  assign n3470 = ~\new_[9533]_  | (~\new_[9694]_  & ~\new_[8706]_ );
  assign \new_[7494]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][12] ;
  assign n3475 = ~\new_[9534]_  | (~\new_[9694]_  & ~\new_[8707]_ );
  assign \new_[7496]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][5] ;
  assign \new_[7497]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][6] ;
  assign \new_[7498]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][12] ;
  assign \new_[7499]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][22] ;
  assign \new_[7500]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][34] ;
  assign \new_[7501]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][6] ;
  assign n5355 = ~\new_[9482]_  | (~\new_[9694]_  & ~\new_[8709]_ );
  assign \new_[7503]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][34] ;
  assign \new_[7504]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][12] ;
  assign \new_[7505]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][22] ;
  assign n3485 = ~\new_[9483]_  | (~\new_[9694]_  & ~\new_[8710]_ );
  assign \new_[7507]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][34] ;
  assign \new_[7508]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][4] ;
  assign \new_[7509]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][5] ;
  assign \new_[7510]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][34] ;
  assign n3490 = ~\new_[9484]_  | (~\new_[9694]_  & ~\new_[8711]_ );
  assign n3495 = ~\new_[9485]_  | (~\new_[9694]_  & ~\new_[8712]_ );
  assign n5340 = ~\new_[9535]_  | (~\new_[9694]_  & ~\new_[8713]_ );
  assign n3500 = \new_[8719]_  ? \new_[9749]_  : \new_[17925]_ ;
  assign n3505 = \new_[8720]_  ? \new_[9718]_  : \new_[19369]_ ;
  assign n3510 = \new_[8721]_  ? \new_[9713]_  : \new_[19664]_ ;
  assign n3515 = \new_[8722]_  ? \new_[9716]_  : \new_[19825]_ ;
  assign n3520 = \new_[8723]_  ? \new_[9669]_  : \new_[18876]_ ;
  assign n3525 = \new_[8724]_  ? \new_[9738]_  : \new_[18654]_ ;
  assign n3530 = \new_[8725]_  ? \new_[9745]_  : \new_[18930]_ ;
  assign n3535 = \new_[8726]_  ? \new_[9735]_  : \new_[18573]_ ;
  assign n3540 = \new_[8727]_  ? \new_[9754]_  : \new_[18720]_ ;
  assign n5320 = \new_[8728]_  ? \new_[9740]_  : \new_[18443]_ ;
  assign n3545 = \new_[8729]_  ? \new_[9609]_  : \new_[18633]_ ;
  assign n3550 = \new_[8731]_  ? \new_[9722]_  : \new_[18366]_ ;
  assign n3555 = \new_[8732]_  ? \new_[9661]_  : \new_[18537]_ ;
  assign n3560 = \new_[8733]_  ? \new_[9669]_  : \new_[19107]_ ;
  assign n3565 = \new_[8734]_  ? \new_[9706]_  : \new_[19113]_ ;
  assign n5305 = \new_[8735]_  ? \new_[9701]_  : \new_[19858]_ ;
  assign n3570 = \new_[8736]_  ? \new_[9704]_  : \new_[18668]_ ;
  assign n3575 = \new_[8737]_  ? \new_[9668]_  : \new_[18292]_ ;
  assign n3580 = \new_[8738]_  ? \new_[9747]_  : \new_[17952]_ ;
  assign n3585 = \new_[8739]_  ? \new_[9733]_  : \new_[18973]_ ;
  assign n3590 = \new_[8740]_  ? \new_[9732]_  : \new_[19089]_ ;
  assign n3595 = \new_[8741]_  ? \new_[9669]_  : \new_[18777]_ ;
  assign n3600 = \new_[8742]_  ? \new_[9700]_  : \new_[18529]_ ;
  assign n3605 = \new_[8743]_  ? \new_[9740]_  : \new_[18820]_ ;
  assign n5285 = \new_[8744]_  ? \new_[9698]_  : \new_[19537]_ ;
  assign n3610 = \new_[8745]_  ? \new_[9723]_  : \new_[18752]_ ;
  assign n3615 = \new_[8746]_  ? \new_[9741]_  : \new_[19118]_ ;
  assign n3620 = \new_[8747]_  ? \new_[9733]_  : \new_[18627]_ ;
  assign n3625 = \new_[8748]_  ? \new_[9725]_  : \new_[18324]_ ;
  assign n3630 = \new_[8749]_  ? \new_[9733]_  : \new_[18342]_ ;
  assign n5275 = \new_[8750]_  ? \new_[9661]_  : \new_[19036]_ ;
  assign n3635 = \new_[8751]_  ? \new_[9669]_  : \new_[19251]_ ;
  assign n3640 = \new_[8752]_  ? \new_[9758]_  : \new_[18135]_ ;
  assign n3670 = \new_[8753]_  ? \new_[9699]_  : \new_[18557]_ ;
  assign n5270 = \new_[8755]_  ? \new_[9733]_  : \new_[18723]_ ;
  assign n3645 = \new_[8754]_  ? \new_[9698]_  : \new_[19372]_ ;
  assign n3650 = \new_[8756]_  ? \new_[9701]_  : \new_[18351]_ ;
  assign n3655 = \new_[8757]_  ? \new_[9722]_  : \new_[19854]_ ;
  assign n3660 = \new_[8758]_  ? \new_[9704]_  : \new_[18707]_ ;
  assign n3665 = \new_[8759]_  ? \new_[9694]_  : \new_[18846]_ ;
  assign n5260 = \new_[8760]_  ? \new_[9698]_  : \new_[17895]_ ;
  assign n5265 = \new_[8761]_  ? \new_[9698]_  : \new_[18869]_ ;
  assign n3675 = \new_[8762]_  ? \new_[9747]_  : \new_[19796]_ ;
  assign n3680 = \new_[8763]_  ? \new_[9753]_  : \new_[19797]_ ;
  assign n3685 = \new_[8764]_  ? \new_[9661]_  : \new_[17823]_ ;
  assign n3690 = \new_[8789]_  ? \new_[9661]_  : \new_[18528]_ ;
  assign n3695 = \new_[8765]_  ? \new_[9732]_  : \new_[18945]_ ;
  assign n3700 = \new_[8766]_  ? \new_[9742]_  : \new_[18826]_ ;
  assign n3705 = \new_[8767]_  ? \new_[9703]_  : \new_[19625]_ ;
  assign n5225 = \new_[8768]_  ? \new_[9746]_  : \new_[18993]_ ;
  assign n3710 = \new_[8769]_  ? \new_[9699]_  : \new_[19561]_ ;
  assign n3715 = \new_[8770]_  ? \new_[9669]_  : \new_[19157]_ ;
  assign n3720 = \new_[8771]_  ? \new_[9669]_  : \new_[17850]_ ;
  assign n3725 = \new_[8772]_  ? \new_[9730]_  : \new_[18191]_ ;
  assign n3730 = \new_[8774]_  ? \new_[9730]_  : \new_[19263]_ ;
  assign n3740 = \new_[8775]_  ? \new_[9757]_  : \new_[19144]_ ;
  assign n3745 = \new_[8776]_  ? \new_[9719]_  : \new_[19260]_ ;
  assign n3735 = \new_[8773]_  ? \new_[9730]_  : \new_[18631]_ ;
  assign n3750 = \new_[8777]_  ? \new_[9698]_  : \new_[18315]_ ;
  assign n5245 = \new_[8778]_  ? \new_[9723]_  : \new_[17942]_ ;
  assign n3755 = \new_[8779]_  ? \new_[9665]_  : \new_[18018]_ ;
  assign n3760 = \new_[8780]_  ? \new_[9729]_  : \new_[19055]_ ;
  assign n3765 = \new_[8781]_  ? \new_[9722]_  : \new_[18641]_ ;
  assign n3770 = \new_[8858]_  ? \new_[9748]_  : \new_[18394]_ ;
  assign n3775 = \new_[8782]_  ? \new_[9733]_  : \new_[18899]_ ;
  assign n5240 = \new_[8783]_  ? \new_[9748]_  : \new_[18225]_ ;
  assign n3780 = \new_[8784]_  ? \new_[9661]_  : \new_[18845]_ ;
  assign n3785 = \new_[8785]_  ? \new_[9702]_  : \new_[19265]_ ;
  assign n3790 = \new_[8786]_  ? \new_[9718]_  : \new_[18287]_ ;
  assign n3795 = \new_[8787]_  ? \new_[9733]_  : \new_[18299]_ ;
  assign n3800 = \new_[8857]_  ? \new_[9661]_  : \new_[19188]_ ;
  assign n3805 = \new_[8788]_  ? \new_[9752]_  : \new_[18501]_ ;
  assign n3810 = \new_[8790]_  ? \new_[9699]_  : \new_[18526]_ ;
  assign n3815 = \new_[8791]_  ? \new_[9733]_  : \new_[19855]_ ;
  assign n5235 = \new_[8792]_  ? \new_[9667]_  : \new_[18844]_ ;
  assign n3820 = \new_[8793]_  ? \new_[9698]_  : \new_[18483]_ ;
  assign n3825 = \new_[8794]_  ? \new_[9701]_  : \new_[19657]_ ;
  assign n3830 = \new_[8795]_  ? \new_[9733]_  : \new_[19648]_ ;
  assign n3835 = \new_[8796]_  ? \new_[9606]_  : \new_[17886]_ ;
  assign n3840 = \new_[8797]_  ? \new_[9722]_  : \new_[19156]_ ;
  assign n3325 = \new_[8798]_  ? \new_[9699]_  : \new_[19388]_ ;
  assign n3845 = \new_[8799]_  ? \new_[9660]_  : \new_[18140]_ ;
  assign n3850 = \new_[8800]_  ? \new_[9608]_  : \new_[19444]_ ;
  assign n3855 = \new_[8801]_  ? \new_[9724]_  : \new_[19279]_ ;
  assign n3860 = \new_[8716]_  ? \new_[9694]_  : \new_[18771]_ ;
  assign n3865 = \new_[8802]_  ? \new_[9698]_  : \new_[18856]_ ;
  assign n3870 = \new_[8803]_  ? \new_[9610]_  : \new_[18730]_ ;
  assign n3875 = \new_[8804]_  ? \new_[9698]_  : \new_[19364]_ ;
  assign n3880 = \new_[8805]_  ? \new_[9745]_  : \new_[18972]_ ;
  assign n3885 = \new_[8806]_  ? \new_[9666]_  : \new_[19320]_ ;
  assign n3890 = \new_[8807]_  ? \new_[9663]_  : \new_[19754]_ ;
  assign n3895 = \new_[8808]_  ? \new_[9721]_  : \new_[19019]_ ;
  assign n3900 = \new_[8809]_  ? \new_[9707]_  : \new_[18695]_ ;
  assign n3905 = \new_[8810]_  ? \new_[9733]_  : \new_[18889]_ ;
  assign n3910 = \new_[8811]_  ? \new_[9714]_  : \new_[19165]_ ;
  assign n5470 = \new_[8812]_  ? \new_[9698]_  : \new_[18749]_ ;
  assign n3915 = \new_[8813]_  ? \new_[9669]_  : \new_[19061]_ ;
  assign n3920 = \new_[8814]_  ? \new_[9730]_  : \new_[18811]_ ;
  assign n3925 = \new_[8815]_  ? \new_[9754]_  : \new_[18857]_ ;
  assign n3930 = \new_[8816]_  ? \new_[9719]_  : \new_[19179]_ ;
  assign n3935 = \new_[8817]_  ? \new_[9661]_  : \new_[19053]_ ;
  assign n5465 = \new_[8714]_  ? \new_[9733]_  : \new_[18891]_ ;
  assign n3940 = \new_[8818]_  ? \new_[9756]_  : \new_[18682]_ ;
  assign n3945 = \new_[8819]_  ? \new_[9734]_  : \new_[20002]_ ;
  assign n3950 = \new_[8820]_  ? \new_[9742]_  : \new_[19611]_ ;
  assign n5460 = \new_[8821]_  ? \new_[9724]_  : \new_[18736]_ ;
  assign n3955 = \new_[8822]_  ? \new_[9715]_  : \new_[18794]_ ;
  assign n3960 = \new_[8823]_  ? \new_[9732]_  : \new_[19602]_ ;
  assign n3965 = \new_[8834]_  ? \new_[9746]_  : \new_[19066]_ ;
  assign n3970 = \new_[8824]_  ? \new_[9712]_  : \new_[18385]_ ;
  assign n3975 = \new_[8825]_  ? \new_[9667]_  : \new_[19200]_ ;
  assign n3980 = \new_[8718]_  ? \new_[9660]_  : \new_[18341]_ ;
  assign n3985 = \new_[8826]_  ? \new_[9669]_  : \new_[18230]_ ;
  assign n3990 = \new_[8827]_  ? \new_[9661]_  : \new_[18776]_ ;
  assign n3995 = \new_[8828]_  ? \new_[9754]_  : \new_[18675]_ ;
  assign n4000 = \new_[8829]_  ? \new_[9721]_  : \new_[19007]_ ;
  assign n4005 = \new_[8830]_  ? \new_[9730]_  : \new_[18148]_ ;
  assign \new_[7631]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][34] ;
  assign n4010 = \new_[8831]_  ? \new_[9738]_  : \new_[17962]_ ;
  assign n4015 = \new_[8832]_  ? \new_[9745]_  : \new_[17910]_ ;
  assign n4020 = \new_[8833]_  ? \new_[9612]_  : \new_[19549]_ ;
  assign n5455 = \new_[8835]_  ? \new_[9664]_  : \new_[18705]_ ;
  assign n4025 = \new_[8836]_  ? \new_[9662]_  : \new_[17980]_ ;
  assign n4030 = \new_[8837]_  ? \new_[9710]_  : \new_[18960]_ ;
  assign n4035 = \new_[8838]_  ? \new_[9660]_  : \new_[19361]_ ;
  assign n4040 = \new_[8839]_  ? \new_[9733]_  : \new_[18359]_ ;
  assign n4045 = \new_[8840]_  ? \new_[9699]_  : \new_[17806]_ ;
  assign \new_[7641]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][4] ;
  assign \new_[7642]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][14] ;
  assign n4050 = \new_[8841]_  ? \new_[9698]_  : \new_[19230]_ ;
  assign n4055 = \new_[8842]_  ? \new_[9729]_  : \new_[19203]_ ;
  assign n4060 = \new_[8843]_  ? \new_[9744]_  : \new_[18195]_ ;
  assign n4065 = \new_[8715]_  ? \new_[9667]_  : \new_[18029]_ ;
  assign n5450 = \new_[8844]_  ? \new_[9663]_  : \new_[17877]_ ;
  assign \new_[7648]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][6] ;
  assign n4070 = \new_[8845]_  ? \new_[9730]_  : \new_[19767]_ ;
  assign n4075 = \new_[8846]_  ? \new_[9717]_  : \new_[18614]_ ;
  assign n4080 = \new_[8847]_  ? \new_[9727]_  : \new_[18532]_ ;
  assign n4085 = \new_[8848]_  ? \new_[9713]_  : \new_[18667]_ ;
  assign n4090 = \new_[8849]_  ? \new_[9665]_  : \new_[18986]_ ;
  assign n5300 = \new_[8850]_  ? \new_[9758]_  : \new_[19787]_ ;
  assign n4095 = \new_[8851]_  ? \new_[9698]_  : \new_[19714]_ ;
  assign n4105 = \new_[8853]_  ? \new_[9607]_  : \new_[19834]_ ;
  assign n4100 = \new_[8852]_  ? \new_[9725]_  : \new_[19800]_ ;
  assign \new_[7658]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][2] ;
  assign n4110 = \new_[8854]_  ? \new_[9733]_  : \new_[18637]_ ;
  assign n4115 = \new_[8855]_  ? \new_[9613]_  : \new_[18691]_ ;
  assign n4120 = \new_[8717]_  ? \new_[9667]_  : \new_[19794]_ ;
  assign n4125 = \new_[8856]_  ? \new_[9667]_  : \new_[17945]_ ;
  assign n4130 = \new_[8863]_  ? \new_[9669]_  : \new_[19853]_ ;
  assign n5445 = \new_[8864]_  ? \new_[9730]_  : \new_[19425]_ ;
  assign \new_[7665]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][25] ;
  assign n4135 = \new_[8865]_  ? \new_[9730]_  : \new_[18354]_ ;
  assign n4140 = \new_[8866]_  ? \new_[9730]_  : \new_[19332]_ ;
  assign n4145 = \new_[8867]_  ? \new_[9717]_  : \new_[17976]_ ;
  assign \new_[7669]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][4] ;
  assign n4150 = \new_[8868]_  ? \new_[9699]_  : \new_[17977]_ ;
  assign n4155 = \new_[8869]_  ? \new_[9699]_  : \new_[19832]_ ;
  assign n5440 = \new_[8870]_  ? \new_[9661]_  : \new_[18117]_ ;
  assign n4160 = \new_[8871]_  ? \new_[9708]_  : \new_[18030]_ ;
  assign \new_[7674]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][22] ;
  assign n4165 = \new_[8872]_  ? \new_[9699]_  : \new_[18569]_ ;
  assign n4170 = \new_[8873]_  ? \new_[9694]_  : \new_[17897]_ ;
  assign n4175 = \new_[8874]_  ? \new_[9699]_  : \new_[19109]_ ;
  assign n4180 = \new_[8875]_  ? \new_[9667]_  : \new_[18963]_ ;
  assign \new_[7679]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][4] ;
  assign n4185 = \new_[8876]_  ? \new_[9720]_  : \new_[19547]_ ;
  assign n4190 = \new_[8877]_  ? \new_[9698]_  : \new_[19645]_ ;
  assign n4195 = \new_[8878]_  ? \new_[9698]_  : \new_[19236]_ ;
  assign n4200 = \new_[8879]_  ? \new_[9710]_  : \new_[18238]_ ;
  assign n5370 = \new_[8880]_  ? \new_[9660]_  : \new_[17864]_ ;
  assign n4205 = \new_[8881]_  ? \new_[9701]_  : \new_[19276]_ ;
  assign n4210 = \new_[8882]_  ? \new_[9660]_  : \new_[19353]_ ;
  assign n5425 = \new_[8883]_  ? \new_[9730]_  : \new_[18101]_ ;
  assign \new_[7688]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][14] ;
  assign n4215 = \new_[8884]_  ? \new_[9733]_  : \new_[18670]_ ;
  assign n4220 = \new_[8885]_  ? \new_[9667]_  : \new_[18969]_ ;
  assign n4225 = \new_[8886]_  ? \new_[9660]_  : \new_[18311]_ ;
  assign n4230 = \new_[8887]_  ? \new_[9660]_  : \new_[18192]_ ;
  assign n5420 = \new_[8888]_  ? \new_[9699]_  : \new_[19305]_ ;
  assign n4235 = \new_[8889]_  ? \new_[9608]_  : \new_[19592]_ ;
  assign n4240 = \new_[8890]_  ? \new_[9730]_  : \new_[18216]_ ;
  assign n4245 = \new_[8891]_  ? \new_[9730]_  : \new_[19405]_ ;
  assign n4250 = \new_[8892]_  ? \new_[9712]_  : \new_[18071]_ ;
  assign n4255 = \new_[8893]_  ? \new_[9715]_  : \new_[19014]_ ;
  assign n5400 = \new_[8894]_  ? \new_[9611]_  : \new_[19700]_ ;
  assign n4260 = \new_[8895]_  ? \new_[9669]_  : \new_[18214]_ ;
  assign n4265 = \new_[8896]_  ? \new_[9730]_  : \new_[19753]_ ;
  assign n4270 = \new_[8897]_  ? \new_[9733]_  : \new_[18692]_ ;
  assign n4275 = \new_[8898]_  ? \new_[9661]_  : \new_[19624]_ ;
  assign \new_[7704]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][25] ;
  assign \new_[7705]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][5] ;
  assign n4280 = \new_[8899]_  ? \new_[9669]_  : \new_[19247]_ ;
  assign \new_[7707]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][22] ;
  assign n4285 = \new_[8900]_  ? \new_[9610]_  : \new_[19149]_ ;
  assign n4290 = \new_[8901]_  ? \new_[9733]_  : \new_[18906]_ ;
  assign n4295 = \new_[8903]_  ? \new_[9745]_  : \new_[19824]_ ;
  assign n4300 = \new_[8904]_  ? \new_[9745]_  : \new_[19394]_ ;
  assign n5385 = \new_[8905]_  ? \new_[9733]_  : \new_[19047]_ ;
  assign n4310 = \new_[8907]_  ? \new_[9745]_  : \new_[19668]_ ;
  assign n4305 = \new_[8906]_  ? \new_[9699]_  : \new_[19718]_ ;
  assign n5125 = ~\new_[20077]_  & ~\new_[20073]_ ;
  assign n5375 = \new_[8908]_  ? \new_[9670]_  : \new_[18416]_ ;
  assign n5220 = ~\new_[20073]_  & ~\new_[20083]_ ;
  assign n4315 = \new_[8909]_  ? \new_[9747]_  : \new_[18694]_ ;
  assign n4320 = \new_[8859]_  ? \new_[9733]_  : \new_[19344]_ ;
  assign n4325 = \new_[8910]_  ? \new_[9743]_  : \new_[19395]_ ;
  assign n4330 = \new_[8911]_  ? \new_[9711]_  : \new_[18718]_ ;
  assign n5350 = \new_[8912]_  ? \new_[9745]_  : \new_[19707]_ ;
  assign n4335 = \new_[8913]_  ? \new_[9743]_  : \new_[18052]_ ;
  assign n4340 = \new_[8914]_  ? \new_[9669]_  : \new_[19368]_ ;
  assign n4345 = \new_[8915]_  ? \new_[9699]_  : \new_[19428]_ ;
  assign n4350 = \new_[8861]_  ? \new_[9612]_  : \new_[18388]_ ;
  assign n4430 = \new_[8916]_  ? \new_[9660]_  : \new_[19383]_ ;
  assign n5365 = \new_[8918]_  ? \new_[9698]_  : \new_[17930]_ ;
  assign n4360 = \new_[8919]_  ? \new_[9669]_  : \new_[18401]_ ;
  assign \new_[7730]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][2] ;
  assign n4365 = \new_[8920]_  ? \new_[9755]_  : \new_[18399]_ ;
  assign n4355 = \new_[8917]_  ? \new_[9733]_  : \new_[19358]_ ;
  assign n4370 = \new_[8921]_  ? \new_[9612]_  : \new_[17929]_ ;
  assign \new_[7734]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][14] ;
  assign n4375 = \new_[8979]_  ? \new_[9698]_  : \new_[17927]_ ;
  assign n4380 = \new_[8922]_  ? \new_[9698]_  : \new_[19414]_ ;
  assign n4385 = \new_[8923]_  ? \new_[9730]_  : \new_[17926]_ ;
  assign \new_[7738]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][25] ;
  assign n4390 = \new_[8924]_  ? \new_[9730]_  : \new_[18455]_ ;
  assign n4395 = \new_[8925]_  ? \new_[9698]_  : \new_[19373]_ ;
  assign \new_[7741]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][25] ;
  assign n4400 = \new_[8926]_  ? \new_[9669]_  : \new_[19198]_ ;
  assign n4405 = \new_[8927]_  ? \new_[9737]_  : \new_[19408]_ ;
  assign n4410 = \new_[8928]_  ? \new_[9726]_  : \new_[17922]_ ;
  assign n4415 = \new_[8929]_  ? \new_[9726]_  : \new_[18453]_ ;
  assign \new_[7746]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][6] ;
  assign \new_[7747]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][6] ;
  assign n4420 = \new_[8930]_  ? \new_[9704]_  : \new_[17916]_ ;
  assign n4425 = \new_[8931]_  ? \new_[9733]_  : \new_[17915]_ ;
  assign n4435 = \new_[8932]_  ? \new_[9734]_  : \new_[19396]_ ;
  assign \new_[7751]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][2] ;
  assign n4440 = \new_[8933]_  ? \new_[9734]_  : \new_[17913]_ ;
  assign n5360 = \new_[8934]_  ? \new_[9745]_  : \new_[17911]_ ;
  assign n4445 = \new_[8935]_  ? \new_[9756]_  : \new_[19106]_ ;
  assign n4450 = \new_[8936]_  ? \new_[9734]_  : \new_[18604]_ ;
  assign n4455 = \new_[8937]_  ? \new_[9708]_  : \new_[19249]_ ;
  assign n4460 = \new_[8860]_  ? \new_[9724]_  : \new_[18952]_ ;
  assign n4465 = \new_[8938]_  ? \new_[9742]_  : \new_[18181]_ ;
  assign n5345 = \new_[8939]_  ? \new_[9716]_  : \new_[20016]_ ;
  assign n4470 = \new_[8940]_  ? \new_[9715]_  : \new_[18513]_ ;
  assign n4475 = \new_[8941]_  ? \new_[9703]_  : \new_[19253]_ ;
  assign n4480 = \new_[8942]_  ? \new_[9660]_  : \new_[19338]_ ;
  assign n5330 = \new_[8943]_  ? \new_[9732]_  : \new_[19335]_ ;
  assign \new_[7764]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][14] ;
  assign n4485 = \new_[8944]_  ? \new_[9735]_  : \new_[18019]_ ;
  assign n4490 = \new_[8945]_  ? \new_[9705]_  : \new_[17992]_ ;
  assign n4495 = \new_[8946]_  ? \new_[9699]_  : \new_[17949]_ ;
  assign n4500 = \new_[8947]_  ? \new_[9667]_  : \new_[17939]_ ;
  assign n4505 = \new_[8948]_  ? \new_[9660]_  : \new_[19514]_ ;
  assign n5335 = \new_[8949]_  ? \new_[9660]_  : \new_[17888]_ ;
  assign \new_[7771]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][34] ;
  assign n4510 = \new_[8950]_  ? \new_[9669]_  : \new_[19268]_ ;
  assign n4515 = \new_[8951]_  ? \new_[9708]_  : \new_[18783]_ ;
  assign n5325 = \new_[8952]_  ? \new_[9699]_  : \new_[17956]_ ;
  assign n4520 = \new_[8953]_  ? \new_[9745]_  : \new_[18796]_ ;
  assign n4525 = \new_[8954]_  ? \new_[9669]_  : \new_[18472]_ ;
  assign \new_[7777]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][25] ;
  assign n4530 = \new_[8955]_  ? \new_[9714]_  : \new_[19406]_ ;
  assign n4535 = \new_[8957]_  ? \new_[9660]_  : \new_[18781]_ ;
  assign n5310 = \new_[8962]_  ? \new_[9606]_  : \new_[18164]_ ;
  assign n4540 = \new_[8956]_  ? \new_[9750]_  : \new_[19223]_ ;
  assign n4545 = \new_[8958]_  ? \new_[9669]_  : \new_[19665]_ ;
  assign \new_[7783]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][34] ;
  assign n4550 = \new_[8959]_  ? \new_[9728]_  : \new_[19545]_ ;
  assign n4555 = \new_[8960]_  ? \new_[9660]_  : \new_[19658]_ ;
  assign n4560 = \new_[8961]_  ? \new_[9700]_  : \new_[18959]_ ;
  assign n5315 = \new_[8963]_  ? \new_[9730]_  : \new_[18516]_ ;
  assign \new_[7788]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][4] ;
  assign n4565 = \new_[8964]_  ? \new_[9731]_  : \new_[18571]_ ;
  assign n4570 = \new_[8965]_  ? \new_[9719]_  : \new_[18790]_ ;
  assign n4575 = \new_[8966]_  ? \new_[9750]_  : \new_[19006]_ ;
  assign n4580 = \new_[8967]_  ? \new_[9662]_  : \new_[18469]_ ;
  assign n4585 = \new_[8968]_  ? \new_[9757]_  : \new_[19788]_ ;
  assign n4590 = \new_[8969]_  ? \new_[9745]_  : \new_[19722]_ ;
  assign n4595 = \new_[8970]_  ? \new_[9738]_  : \new_[19022]_ ;
  assign n4600 = \new_[8971]_  ? \new_[9664]_  : \new_[19727]_ ;
  assign n4605 = \new_[8972]_  ? \new_[9669]_  : \new_[18563]_ ;
  assign n5290 = \new_[8973]_  ? \new_[9730]_  : \new_[19092]_ ;
  assign n4610 = \new_[8862]_  ? \new_[9660]_  : \new_[19612]_ ;
  assign n4615 = \new_[8974]_  ? \new_[9664]_  : \new_[18231]_ ;
  assign n5295 = \new_[8975]_  ? \new_[9698]_  : \new_[18559]_ ;
  assign \new_[7802]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][25] ;
  assign \new_[7803]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][2] ;
  assign n4620 = \new_[8976]_  ? \new_[9660]_  : \new_[19391]_ ;
  assign n4625 = \new_[8977]_  ? \new_[9660]_  : \new_[19370]_ ;
  assign \new_[7806]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][34] ;
  assign n4630 = \new_[8978]_  ? \new_[9723]_  : \new_[19059]_ ;
  assign n5190 = \new_[9094]_  ? \new_[9723]_  : \new_[18093]_ ;
  assign n4635 = \new_[8983]_  ? \new_[9660]_  : \new_[17983]_ ;
  assign n4640 = \new_[8984]_  ? \new_[9609]_  : \new_[19103]_ ;
  assign n4645 = \new_[8985]_  ? \new_[9741]_  : \new_[19079]_ ;
  assign n4650 = \new_[8986]_  ? \new_[9744]_  : \new_[18257]_ ;
  assign n4655 = \new_[8987]_  ? \new_[9729]_  : \new_[18655]_ ;
  assign n4660 = \new_[8988]_  ? \new_[9660]_  : \new_[18818]_ ;
  assign n4670 = \new_[8990]_  ? \new_[9733]_  : \new_[18504]_ ;
  assign n4665 = \new_[8989]_  ? \new_[9733]_  : \new_[19659]_ ;
  assign n5430 = ~\new_[8242]_ ;
  assign n5280 = \new_[8991]_  ? \new_[9667]_  : \new_[17879]_ ;
  assign \new_[7819]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][22] ;
  assign n4675 = \new_[8992]_  ? \new_[9717]_  : \new_[18444]_ ;
  assign n3450 = ~\new_[8242]_ ;
  assign \new_[7822]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][12] ;
  assign n4680 = \new_[8993]_  ? \new_[9663]_  : \new_[19495]_ ;
  assign n4685 = \new_[8994]_  ? \new_[9661]_  : \new_[19206]_ ;
  assign n3425 = ~\new_[8242]_ ;
  assign n4690 = \new_[8995]_  ? \new_[9730]_  : \new_[18106]_ ;
  assign n5435 = ~\new_[8242]_ ;
  assign n4695 = \new_[8996]_  ? \new_[9667]_  : \new_[18997]_ ;
  assign n3375 = ~\new_[8242]_ ;
  assign n5395 = ~\new_[8242]_ ;
  assign n4700 = \new_[8997]_  ? \new_[9727]_  : \new_[19581]_ ;
  assign n3410 = ~\new_[8242]_ ;
  assign n4705 = \new_[8998]_  ? \new_[9733]_  : \new_[18285]_ ;
  assign n5405 = ~\new_[8242]_ ;
  assign n4710 = \new_[8999]_  ? \new_[9727]_  : \new_[18121]_ ;
  assign n3360 = ~\new_[8242]_ ;
  assign n4715 = \new_[9000]_  ? \new_[9698]_  : \new_[19352]_ ;
  assign n5410 = ~\new_[8242]_ ;
  assign n3435 = ~\new_[8242]_ ;
  assign n5390 = ~\new_[8242]_ ;
  assign n4720 = \new_[9001]_  ? \new_[9712]_  : \new_[18578]_ ;
  assign n4725 = \new_[9002]_  ? \new_[9698]_  : \new_[17904]_ ;
  assign n4730 = \new_[9003]_  ? \new_[9698]_  : \new_[18947]_ ;
  assign \new_[7844]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][14] ;
  assign n4735 = \new_[9004]_  ? \new_[9698]_  : \new_[18636]_ ;
  assign n4740 = \new_[9005]_  ? \new_[9663]_  : \new_[18329]_ ;
  assign n4750 = \new_[9006]_  ? \new_[9660]_  : \new_[19607]_ ;
  assign n4745 = \new_[9007]_  ? \new_[9725]_  : \new_[18931]_ ;
  assign n4755 = \new_[9008]_  ? \new_[9702]_  : \new_[18484]_ ;
  assign n4760 = \new_[9009]_  ? \new_[9718]_  : \new_[18242]_ ;
  assign n5255 = \new_[9010]_  ? \new_[9713]_  : \new_[19446]_ ;
  assign n4765 = \new_[9011]_  ? \new_[9751]_  : \new_[19421]_ ;
  assign n4770 = \new_[9079]_  ? \new_[9739]_  : \new_[18077]_ ;
  assign n4775 = \new_[9012]_  ? \new_[9733]_  : \new_[18905]_ ;
  assign n4780 = \new_[9013]_  ? \new_[9733]_  : \new_[18064]_ ;
  assign n4785 = \new_[9014]_  ? \new_[9661]_  : \new_[18981]_ ;
  assign n5250 = \new_[9015]_  ? \new_[9718]_  : \new_[19697]_ ;
  assign n4790 = \new_[9016]_  ? \new_[9613]_  : \new_[19566]_ ;
  assign n4795 = \new_[9017]_  ? \new_[9702]_  : \new_[19087]_ ;
  assign n4800 = \new_[9018]_  ? \new_[9739]_  : \new_[18878]_ ;
  assign \new_[7861]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][6] ;
  assign n4805 = \new_[9019]_  ? \new_[9709]_  : \new_[17973]_ ;
  assign n4810 = \new_[9020]_  ? \new_[9607]_  : \new_[19988]_ ;
  assign n4815 = \new_[9021]_  ? \new_[9660]_  : \new_[18621]_ ;
  assign n4820 = \new_[9022]_  ? \new_[9709]_  : \new_[19057]_ ;
  assign \new_[7866]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][6] ;
  assign n4825 = \new_[9023]_  ? \new_[9663]_  : \new_[18326]_ ;
  assign n4830 = \new_[9024]_  ? \new_[9736]_  : \new_[19693]_ ;
  assign \new_[7869]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][34] ;
  assign n4835 = \new_[9025]_  ? \new_[9758]_  : \new_[19073]_ ;
  assign n4840 = \new_[9026]_  ? \new_[9661]_  : \new_[19680]_ ;
  assign n4845 = \new_[9027]_  ? \new_[9730]_  : \new_[19267]_ ;
  assign n4850 = \new_[9028]_  ? \new_[9698]_  : \new_[18863]_ ;
  assign n4855 = \new_[9029]_  ? \new_[9748]_  : \new_[19243]_ ;
  assign n4860 = \new_[9030]_  ? \new_[9733]_  : \new_[18898]_ ;
  assign n4865 = \new_[9031]_  ? \new_[9730]_  : \new_[18881]_ ;
  assign n4870 = \new_[9032]_  ? \new_[9605]_  : \new_[18070]_ ;
  assign n4875 = \new_[9033]_  ? \new_[9730]_  : \new_[18979]_ ;
  assign n4880 = \new_[9034]_  ? \new_[9752]_  : \new_[19035]_ ;
  assign n4885 = \new_[9035]_  ? \new_[9752]_  : \new_[19085]_ ;
  assign n4890 = \new_[9036]_  ? \new_[9752]_  : \new_[19300]_ ;
  assign n4895 = \new_[9037]_  ? \new_[9744]_  : \new_[19460]_ ;
  assign n4900 = \new_[9038]_  ? \new_[9661]_  : \new_[17901]_ ;
  assign n4905 = \new_[9039]_  ? \new_[9729]_  : \new_[18687]_ ;
  assign n5230 = \new_[9127]_  ? \new_[9699]_  : \new_[18964]_ ;
  assign n4910 = \new_[9040]_  ? \new_[9744]_  : \new_[18601]_ ;
  assign n4915 = \new_[9041]_  ? \new_[9698]_  : \new_[18983]_ ;
  assign n4920 = \new_[9042]_  ? \new_[9741]_  : \new_[18975]_ ;
  assign n4925 = \new_[9043]_  ? \new_[9665]_  : \new_[18567]_ ;
  assign n4930 = \new_[9044]_  ? \new_[9609]_  : \new_[18630]_ ;
  assign n4935 = \new_[9045]_  ? \new_[9667]_  : \new_[18381]_ ;
  assign n4940 = \new_[9046]_  ? \new_[9609]_  : \new_[19635]_ ;
  assign n4945 = \new_[9047]_  ? \new_[9749]_  : \new_[19101]_ ;
  assign n4950 = \new_[9048]_  ? \new_[9749]_  : \new_[18530]_ ;
  assign \new_[7895]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][14] ;
  assign n4955 = \new_[9049]_  ? \new_[9698]_  : \new_[19176]_ ;
  assign n4960 = \new_[9050]_  ? \new_[9731]_  : \new_[18218]_ ;
  assign n4965 = \new_[9051]_  ? \new_[9706]_  : \new_[18544]_ ;
  assign n4970 = \new_[9052]_  ? \new_[9612]_  : \new_[18186]_ ;
  assign \new_[7900]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][6] ;
  assign n4975 = \new_[9053]_  ? \new_[9710]_  : \new_[18112]_ ;
  assign n4980 = \new_[9054]_  ? \new_[9730]_  : \new_[19441]_ ;
  assign n4985 = \new_[9055]_  ? \new_[9745]_  : \new_[19443]_ ;
  assign n4990 = \new_[9056]_  ? \new_[9745]_  : \new_[18034]_ ;
  assign n4995 = \new_[9057]_  ? \new_[9661]_  : \new_[19450]_ ;
  assign n3320 = \new_[9058]_  ? \new_[9705]_  : \new_[18004]_ ;
  assign n5000 = \new_[9059]_  ? \new_[9606]_  : \new_[17990]_ ;
  assign n5005 = \new_[9060]_  ? \new_[9700]_  : \new_[19490]_ ;
  assign n5010 = \new_[9061]_  ? \new_[9730]_  : \new_[19749]_ ;
  assign \new_[7910]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][14] ;
  assign n5015 = \new_[9062]_  ? \new_[9700]_  : \new_[19518]_ ;
  assign n5020 = \new_[9063]_  ? \new_[9662]_  : \new_[19065]_ ;
  assign n3330 = \new_[9064]_  ? \new_[9706]_  : \new_[19699]_ ;
  assign n5025 = \new_[9065]_  ? \new_[9669]_  : \new_[19543]_ ;
  assign n5030 = \new_[9066]_  ? \new_[9667]_  : \new_[18722]_ ;
  assign n5035 = \new_[9067]_  ? \new_[9721]_  : \new_[17834]_ ;
  assign n5040 = \new_[9068]_  ? \new_[9661]_  : \new_[19086]_ ;
  assign n5045 = \new_[9069]_  ? \new_[9606]_  : \new_[19984]_ ;
  assign n5050 = \new_[8982]_  ? \new_[9705]_  : \new_[19757]_ ;
  assign n5055 = \new_[9070]_  ? \new_[9708]_  : \new_[19214]_ ;
  assign \new_[7921]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][12] ;
  assign n5060 = \new_[9071]_  ? \new_[9714]_  : \new_[18753]_ ;
  assign n5065 = \new_[9072]_  ? \new_[9669]_  : \new_[18103]_ ;
  assign n5070 = \new_[9073]_  ? \new_[9703]_  : \new_[17848]_ ;
  assign n5075 = \new_[9074]_  ? \new_[9661]_  : \new_[19386]_ ;
  assign \new_[7926]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][25] ;
  assign n5080 = \new_[9075]_  ? \new_[9730]_  : \new_[18014]_ ;
  assign n5085 = \new_[9076]_  ? \new_[9755]_  : \new_[19010]_ ;
  assign n5090 = \new_[8980]_  ? \new_[9668]_  : \new_[19097]_ ;
  assign n5095 = \new_[9077]_  ? \new_[9669]_  : \new_[19689]_ ;
  assign n5100 = \new_[9078]_  ? \new_[9694]_  : \new_[17982]_ ;
  assign n5105 = \new_[9080]_  ? \new_[9608]_  : \new_[18198]_ ;
  assign n5110 = \new_[9081]_  ? \new_[9745]_  : \new_[19600]_ ;
  assign n5115 = \new_[9082]_  ? \new_[9745]_  : \new_[18929]_ ;
  assign \new_[7935]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][14] ;
  assign n5120 = \new_[9083]_  ? \new_[9661]_  : \new_[17807]_ ;
  assign n5130 = \new_[9084]_  ? \new_[9711]_  : \new_[18581]_ ;
  assign n5135 = \new_[9102]_  ? \new_[9745]_  : \new_[18961]_ ;
  assign n5140 = \new_[9085]_  ? \new_[9745]_  : \new_[19238]_ ;
  assign n5485 = \new_[9086]_  ? \new_[9733]_  : \new_[20000]_ ;
  assign n5145 = \new_[9087]_  ? \new_[9733]_  : \new_[19867]_ ;
  assign n5150 = \new_[9128]_  ? \new_[9733]_  : \new_[19652]_ ;
  assign n5155 = \new_[9088]_  ? \new_[9711]_  : \new_[18384]_ ;
  assign \new_[7944]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][4] ;
  assign n5480 = \new_[9089]_  ? \new_[9666]_  : \new_[19840]_ ;
  assign n5160 = \new_[9100]_  ? \new_[9745]_  : \new_[18585]_ ;
  assign n5165 = \new_[9090]_  ? \new_[9660]_  : \new_[19677]_ ;
  assign n5170 = \new_[9091]_  ? \new_[9699]_  : \new_[18314]_ ;
  assign n5175 = \new_[9099]_  ? \new_[9720]_  : \new_[19205]_ ;
  assign n5180 = \new_[9092]_  ? \new_[9670]_  : \new_[19110]_ ;
  assign n5475 = \new_[9093]_  ? \new_[9660]_  : \new_[19241]_ ;
  assign n5185 = \new_[8981]_  ? \new_[9670]_  : \new_[18536]_ ;
  assign \new_[7953]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][6] ;
  assign \new_[7954]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][2] ;
  assign n5195 = \new_[9095]_  ? \new_[9753]_  : \new_[18436]_ ;
  assign n5200 = \new_[9096]_  ? \new_[9753]_  : \new_[19252]_ ;
  assign n5205 = \new_[9097]_  ? \new_[9728]_  : \new_[18219]_ ;
  assign n5210 = \new_[9101]_  ? \new_[9745]_  : \new_[19798]_ ;
  assign n5215 = \new_[9098]_  ? \new_[9660]_  : \new_[19033]_ ;
  assign \new_[7960]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][25] ;
  assign \new_[7961]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][22] ;
  assign \new_[7962]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][14] ;
  assign \new_[7963]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][6] ;
  assign \new_[7964]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][25] ;
  assign \new_[7965]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][14] ;
  assign \new_[7966]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][25] ;
  assign \new_[7967]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][6] ;
  assign \new_[7968]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][34] ;
  assign \new_[7969]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][2] ;
  assign \new_[7970]_  = (~\new_[20493]_  | ~\new_[19743]_ ) & (~\new_[8682]_  | ~\new_[19679]_ );
  assign \new_[7971]_  = (~\new_[20501]_  | ~\new_[19235]_ ) & (~\new_[8730]_  | ~\new_[18871]_ );
  assign \new_[7972]_  = (~\new_[20493]_  | ~\new_[17964]_ ) & (~\new_[8682]_  | ~\new_[19739]_ );
  assign \new_[7973]_  = (~\new_[20480]_  | ~\new_[18373]_ ) & (~\new_[8697]_  | ~\new_[19776]_ );
  assign \new_[7974]_  = (~\new_[20481]_  | ~\new_[18419]_ ) & (~\new_[8697]_  | ~\new_[19779]_ );
  assign \new_[7975]_  = (~\new_[20504]_  | ~\new_[19562]_ ) & (~\new_[9132]_  | ~\new_[19795]_ );
  assign \new_[7976]_  = (~\new_[20493]_  | ~\new_[19291]_ ) & (~\new_[8682]_  | ~\new_[19043]_ );
  assign \new_[7977]_  = (~\new_[20501]_  | ~\new_[19208]_ ) & (~\new_[8730]_  | ~\new_[19016]_ );
  assign \new_[7978]_  = (~\new_[20481]_  | ~\new_[19686]_ ) & (~\new_[8697]_  | ~\new_[19780]_ );
  assign \new_[7979]_  = (~\new_[9190]_  | ~\new_[18510]_ ) & (~\new_[8686]_  | ~\new_[18840]_ );
  assign \new_[7980]_  = (~\new_[20484]_  | ~\new_[19709]_ ) & (~\new_[8684]_  | ~\new_[18588]_ );
  assign \new_[7981]_  = (~\new_[20493]_  | ~\new_[19292]_ ) & (~\new_[8682]_  | ~\new_[17912]_ );
  assign \new_[7982]_  = (~\new_[20501]_  | ~\new_[18086]_ ) & (~\new_[8730]_  | ~\new_[19210]_ );
  assign \new_[7983]_  = (~\new_[20481]_  | ~\new_[19354]_ ) & (~\new_[8697]_  | ~\new_[19768]_ );
  assign \new_[7984]_  = (~\new_[9190]_  | ~\new_[19017]_ ) & (~\new_[8686]_  | ~\new_[18617]_ );
  assign \new_[7985]_  = (~\new_[20493]_  | ~\new_[18562]_ ) & (~\new_[8682]_  | ~\new_[19821]_ );
  assign \new_[7986]_  = (~\new_[20501]_  | ~\new_[19015]_ ) & (~\new_[8730]_  | ~\new_[18868]_ );
  assign \new_[7987]_  = (~\new_[20481]_  | ~\new_[17896]_ ) & (~\new_[8697]_  | ~\new_[18579]_ );
  assign \new_[7988]_  = (~\new_[20493]_  | ~\new_[19810]_ ) & (~\new_[8682]_  | ~\new_[17909]_ );
  assign \new_[7989]_  = (~\new_[9190]_  | ~\new_[18076]_ ) & (~\new_[8685]_  | ~\new_[18774]_ );
  assign \new_[7990]_  = (~\new_[20504]_  | ~\new_[19082]_ ) & (~\new_[8730]_  | ~\new_[19752]_ );
  assign \new_[7991]_  = (~\new_[20480]_  | ~\new_[19801]_ ) & (~\new_[8697]_  | ~\new_[18253]_ );
  assign \new_[7992]_  = (~\new_[9190]_  | ~\new_[18597]_ ) & (~\new_[8686]_  | ~\new_[18900]_ );
  assign \new_[7993]_  = (~\new_[20482]_  | ~\new_[19168]_ ) & (~\new_[8684]_  | ~\new_[18619]_ );
  assign \new_[7994]_  = (~\new_[20504]_  | ~\new_[19137]_ ) & (~\new_[9132]_  | ~\new_[19211]_ );
  assign \new_[7995]_  = (~\new_[9190]_  | ~\new_[18932]_ ) & (~\new_[8686]_  | ~\new_[18069]_ );
  assign \new_[7996]_  = (~\new_[20503]_  | ~\new_[19256]_ ) & (~\new_[9132]_  | ~\new_[19217]_ );
  assign \new_[7997]_  = (~\new_[20484]_  | ~\new_[18038]_ ) & (~\new_[8683]_  | ~\new_[19302]_ );
  assign \new_[7998]_  = (~\new_[9190]_  | ~\new_[19000]_ ) & (~\new_[9133]_  | ~\new_[18940]_ );
  assign \new_[7999]_  = (~\new_[20493]_  | ~\new_[19808]_ ) & (~\new_[8682]_  | ~\new_[19463]_ );
  assign \new_[8000]_  = (~\new_[20503]_  | ~\new_[18200]_ ) & (~\new_[9132]_  | ~\new_[18113]_ );
  assign \new_[8001]_  = (~\new_[20484]_  | ~\new_[17985]_ ) & (~\new_[8684]_  | ~\new_[19710]_ );
  assign \new_[8002]_  = (~\new_[9190]_  | ~\new_[18107]_ ) & (~\new_[9133]_  | ~\new_[18941]_ );
  assign \new_[8003]_  = (~\new_[20493]_  | ~\new_[18162]_ ) & (~\new_[8682]_  | ~\new_[19124]_ );
  assign \new_[8004]_  = (~\new_[20480]_  | ~\new_[19643]_ ) & (~\new_[8684]_  | ~\new_[18263]_ );
  assign \new_[8005]_  = (~\new_[20501]_  | ~\new_[19790]_ ) & (~\new_[8730]_  | ~\new_[18111]_ );
  assign \new_[8006]_  = (~\new_[20482]_  | ~\new_[19169]_ ) & (~\new_[8697]_  | ~\new_[19777]_ );
  assign \new_[8007]_  = (~\new_[9190]_  | ~\new_[19826]_ ) & (~\new_[9133]_  | ~\new_[19487]_ );
  assign \new_[8008]_  = (~\new_[20503]_  | ~\new_[18201]_ ) & (~\new_[9132]_  | ~\new_[19212]_ );
  assign \new_[8009]_  = (~\new_[20493]_  | ~\new_[17994]_ ) & (~\new_[8682]_  | ~\new_[19342]_ );
  assign \new_[8010]_  = (~\new_[9190]_  | ~\new_[19407]_ ) & (~\new_[8686]_  | ~\new_[19183]_ );
  assign \new_[8011]_  = (~\new_[20493]_  | ~\new_[19148]_ ) & (~\new_[8682]_  | ~\new_[19741]_ );
  assign \new_[8012]_  = (~\new_[20484]_  | ~\new_[17978]_ ) & (~\new_[8683]_  | ~\new_[19297]_ );
  assign \new_[8013]_  = (~\new_[20482]_  | ~\new_[19802]_ ) & (~\new_[8697]_  | ~\new_[19774]_ );
  assign \new_[8014]_  = (~\new_[20504]_  | ~\new_[19673]_ ) & (~\new_[8730]_  | ~\new_[19682]_ );
  assign \new_[8015]_  = (~\new_[20493]_  | ~\new_[17998]_ ) & (~\new_[8682]_  | ~\new_[19819]_ );
  assign \new_[8016]_  = (~\new_[9190]_  | ~\new_[18835]_ ) & (~\new_[8685]_  | ~\new_[19595]_ );
  assign \new_[8017]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][22] ;
  assign \new_[8018]_  = (~\new_[20484]_  | ~\new_[19747]_ ) & (~\new_[8697]_  | ~\new_[19400]_ );
  assign \new_[8019]_  = (~\new_[9190]_  | ~\new_[18179]_ ) & (~\new_[8685]_  | ~\new_[18522]_ );
  assign \new_[8020]_  = (~\new_[20493]_  | ~\new_[17997]_ ) & (~\new_[8682]_  | ~\new_[19459]_ );
  assign \new_[8021]_  = (~\new_[9190]_  | ~\new_[18178]_ ) & (~\new_[9133]_  | ~\new_[19399]_ );
  assign \new_[8022]_  = (~\new_[20493]_  | ~\new_[19725]_ ) & (~\new_[8682]_  | ~\new_[18331]_ );
  assign \new_[8023]_  = (~\new_[20503]_  | ~\new_[18213]_ ) & (~\new_[8730]_  | ~\new_[19598]_ );
  assign \new_[8024]_  = (~\new_[20484]_  | ~\new_[18067]_ ) & (~\new_[8683]_  | ~\new_[18422]_ );
  assign \new_[8025]_  = (~\new_[9190]_  | ~\new_[18174]_ ) & (~\new_[8686]_  | ~\new_[18476]_ );
  assign \new_[8026]_  = (~\new_[20503]_  | ~\new_[19120]_ ) & (~\new_[9132]_  | ~\new_[19218]_ );
  assign \new_[8027]_  = (~\new_[20484]_  | ~\new_[19799]_ ) & (~\new_[8683]_  | ~\new_[18380]_ );
  assign \new_[8028]_  = (~\new_[20482]_  | ~\new_[18055]_ ) & (~\new_[8697]_  | ~\new_[18938]_ );
  assign \new_[8029]_  = (~\new_[20504]_  | ~\new_[19789]_ ) & (~\new_[8730]_  | ~\new_[18126]_ );
  assign \new_[8030]_  = (~\new_[9190]_  | ~\new_[18169]_ ) & (~\new_[8686]_  | ~\new_[18935]_ );
  assign \new_[8031]_  = (~\new_[20484]_  | ~\new_[19174]_ ) & (~\new_[8697]_  | ~\new_[18036]_ );
  assign \new_[8032]_  = (~\new_[20493]_  | ~\new_[19512]_ ) & (~\new_[8682]_  | ~\new_[19816]_ );
  assign \new_[8033]_  = (~\new_[9190]_  | ~\new_[18168]_ ) & (~\new_[9133]_  | ~\new_[18353]_ );
  assign \new_[8034]_  = (~\new_[20480]_  | ~\new_[19672]_ ) & (~\new_[8684]_  | ~\new_[19008]_ );
  assign \new_[8035]_  = (~\new_[20504]_  | ~\new_[19117]_ ) & (~\new_[8730]_  | ~\new_[19584]_ );
  assign \new_[8036]_  = (~\new_[9190]_  | ~\new_[18160]_ ) & (~\new_[9133]_  | ~\new_[18539]_ );
  assign \new_[8037]_  = (~\new_[20481]_  | ~\new_[19748]_ ) & (~\new_[8697]_  | ~\new_[18350]_ );
  assign \new_[8038]_  = (~\new_[20503]_  | ~\new_[19013]_ ) & (~\new_[9132]_  | ~\new_[18159]_ );
  assign \new_[8039]_  = (~\new_[20493]_  | ~\new_[19582]_ ) & (~\new_[8682]_  | ~\new_[19807]_ );
  assign \new_[8040]_  = (~\new_[20480]_  | ~\new_[18062]_ ) & (~\new_[8684]_  | ~\new_[19773]_ );
  assign \new_[8041]_  = (~\new_[20493]_  | ~\new_[18989]_ ) & (~\new_[8682]_  | ~\new_[19812]_ );
  assign \new_[8042]_  = (~\new_[20482]_  | ~\new_[19653]_ ) & (~\new_[8697]_  | ~\new_[19685]_ );
  assign \new_[8043]_  = (~\new_[9190]_  | ~\new_[19114]_ ) & (~\new_[8685]_  | ~\new_[17839]_ );
  assign \new_[8044]_  = (~\new_[20493]_  | ~\new_[19151]_ ) & (~\new_[8682]_  | ~\new_[19108]_ );
  assign \new_[8045]_  = (~\new_[9190]_  | ~\new_[18580]_ ) & (~\new_[9133]_  | ~\new_[18312]_ );
  assign \new_[8046]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][25] ;
  assign \new_[8047]_  = (~\new_[20503]_  | ~\new_[18223]_ ) & (~\new_[9132]_  | ~\new_[19838]_ );
  assign \new_[8048]_  = (~\new_[20484]_  | ~\new_[19182]_ ) & (~\new_[8683]_  | ~\new_[18356]_ );
  assign \new_[8049]_  = (~\new_[20480]_  | ~\new_[19186]_ ) & (~\new_[8697]_  | ~\new_[19732]_ );
  assign \new_[8050]_  = (~\new_[20493]_  | ~\new_[19669]_ ) & (~\new_[8682]_  | ~\new_[19726]_ );
  assign \new_[8051]_  = (~\new_[20481]_  | ~\new_[18079]_ ) & (~\new_[8697]_  | ~\new_[19434]_ );
  assign \new_[8052]_  = (~\new_[20493]_  | ~\new_[18021]_ ) & (~\new_[9270]_  | ~\new_[19704]_ );
  assign \new_[8053]_  = (~\new_[20504]_  | ~\new_[19054]_ ) & (~\new_[9132]_  | ~\new_[19233]_ );
  assign \new_[8054]_  = (~\new_[20493]_  | ~\new_[19158]_ ) & (~\new_[8682]_  | ~\new_[18302]_ );
  assign \new_[8055]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][14] ;
  assign \new_[8056]_  = (~\new_[9190]_  | ~\new_[17892]_ ) & (~\new_[8685]_  | ~\new_[18874]_ );
  assign \new_[8057]_  = (~\new_[20484]_  | ~\new_[19623]_ ) & (~\new_[8683]_  | ~\new_[19438]_ );
  assign \new_[8058]_  = (~\new_[20482]_  | ~\new_[19202]_ ) & (~\new_[8697]_  | ~\new_[19771]_ );
  assign \new_[8059]_  = (~\new_[20504]_  | ~\new_[19782]_ ) & (~\new_[8730]_  | ~\new_[19716]_ );
  assign \new_[8060]_  = (~\new_[9190]_  | ~\new_[18096]_ ) & (~\new_[8685]_  | ~\new_[18925]_ );
  assign \new_[8061]_  = (~\new_[20493]_  | ~\new_[19164]_ ) & (~\new_[8682]_  | ~\new_[19317]_ );
  assign \new_[8062]_  = (~\new_[20504]_  | ~\new_[19783]_ ) & (~\new_[8730]_  | ~\new_[19756]_ );
  assign \new_[8063]_  = (~\new_[20493]_  | ~\new_[19160]_ ) & (~\new_[8682]_  | ~\new_[19833]_ );
  assign \new_[8064]_  = (~\new_[20480]_  | ~\new_[17889]_ ) & (~\new_[8697]_  | ~\new_[19772]_ );
  assign \new_[8065]_  = (~\new_[9190]_  | ~\new_[19309]_ ) & (~\new_[8685]_  | ~\new_[18194]_ );
  assign \new_[8066]_  = (~\new_[9190]_  | ~\new_[19021]_ ) & (~\new_[8686]_  | ~\new_[17919]_ );
  assign \new_[8067]_  = (~\new_[20493]_  | ~\new_[19803]_ ) & (~\new_[8682]_  | ~\new_[19670]_ );
  assign \new_[8068]_  = (~\new_[20482]_  | ~\new_[19617]_ ) & (~\new_[8697]_  | ~\new_[18367]_ );
  assign \new_[8069]_  = (~\new_[20481]_  | ~\new_[18092]_ ) & (~\new_[8697]_  | ~\new_[19347]_ );
  assign \new_[8070]_  = (~\new_[20503]_  | ~\new_[19765]_ ) & (~\new_[8730]_  | ~\new_[18212]_ );
  assign \new_[8071]_  = (~\new_[20493]_  | ~\new_[19650]_ ) & (~\new_[8682]_  | ~\new_[17955]_ );
  assign \new_[8072]_  = (~\new_[9190]_  | ~\new_[18924]_ ) & (~\new_[8685]_  | ~\new_[18197]_ );
  assign \new_[8073]_  = (~\new_[20482]_  | ~\new_[19363]_ ) & (~\new_[8697]_  | ~\new_[18370]_ );
  assign \new_[8074]_  = (~\new_[20481]_  | ~\new_[18147]_ ) & (~\new_[8697]_  | ~\new_[19435]_ );
  assign \new_[8075]_  = (~\new_[20504]_  | ~\new_[19864]_ ) & (~\new_[8730]_  | ~\new_[19791]_ );
  assign \new_[8076]_  = (~\new_[20493]_  | ~\new_[18024]_ ) & (~\new_[8682]_  | ~\new_[17853]_ );
  assign \new_[8077]_  = (~\new_[9190]_  | ~\new_[17900]_ ) & (~\new_[8685]_  | ~\new_[18547]_ );
  assign \new_[8078]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][12] ;
  assign \new_[8079]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][34] ;
  assign \new_[8080]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][6] ;
  assign \new_[8081]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][2] ;
  assign \new_[8082]_  = ~\new_[8275]_ ;
  assign \new_[8083]_  = ~\new_[8275]_ ;
  assign \new_[8084]_  = ~\new_[8275]_ ;
  assign \new_[8085]_  = ~\new_[8275]_ ;
  assign \new_[8086]_  = ~\new_[8275]_ ;
  assign \new_[8087]_  = \new_[8276]_ ;
  assign \new_[8088]_  = ~\new_[8276]_ ;
  assign \new_[8089]_  = ~\new_[8280]_ ;
  assign \new_[8090]_  = ~\new_[8280]_ ;
  assign \new_[8091]_  = \new_[20334]_ ;
  assign \new_[8092]_  = ~\new_[20334]_ ;
  assign \new_[8093]_  = ~\new_[8281]_ ;
  assign \new_[8094]_  = ~\new_[8281]_ ;
  assign \new_[8095]_  = ~\new_[8282]_ ;
  assign \new_[8096]_  = \new_[8282]_ ;
  assign \new_[8097]_  = ~\new_[8283]_ ;
  assign \new_[8098]_  = \new_[8283]_ ;
  assign \new_[8099]_  = \new_[8283]_ ;
  assign \new_[8100]_  = ~\new_[8286]_ ;
  assign \new_[8101]_  = \new_[8287]_ ;
  assign \new_[8102]_  = ~\new_[8287]_ ;
  assign \new_[8103]_  = \new_[8288]_ ;
  assign \new_[8104]_  = ~\new_[8288]_ ;
  assign \new_[8105]_  = \new_[8289]_ ;
  assign \new_[8106]_  = ~\new_[8289]_ ;
  assign \new_[8107]_  = ~\new_[8569]_ ;
  assign \new_[8108]_  = ~\new_[8569]_ ;
  assign \new_[8109]_  = \new_[8569]_ ;
  assign \new_[8110]_  = ~\new_[8569]_ ;
  assign \new_[8111]_  = \new_[8290]_ ;
  assign \new_[8112]_  = ~\new_[8290]_ ;
  assign \new_[8113]_  = \new_[8291]_ ;
  assign \new_[8114]_  = ~\new_[8291]_ ;
  assign \new_[8115]_  = ~\new_[8292]_ ;
  assign \new_[8116]_  = (~\new_[9297]_  | ~\new_[17983]_ ) & (~\new_[9206]_  | ~\new_[18781]_ );
  assign \new_[8117]_  = (~\new_[8700]_  | ~\new_[18979]_ ) & (~\new_[9510]_  | ~\new_[18752]_ );
  assign \new_[8118]_  = (~\new_[19986]_  | ~\new_[18242]_ ) & (~\new_[20552]_  | ~\new_[19450]_ );
  assign \new_[8119]_  = (~\new_[9290]_  | ~\new_[19369]_ ) & (~\new_[9298]_  | ~\new_[17980]_ );
  assign \new_[8120]_  = (~\new_[9295]_  | ~\new_[19035]_ ) & (~\new_[9510]_  | ~\new_[19118]_ );
  assign \new_[8121]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][22] ;
  assign \new_[8122]_  = (~\new_[19986]_  | ~\new_[19446]_ ) & (~\new_[20552]_  | ~\new_[18004]_ );
  assign \new_[8123]_  = (~\new_[9290]_  | ~\new_[19664]_ ) & (~\new_[9298]_  | ~\new_[18960]_ );
  assign \new_[8124]_  = ~\new_[8296]_ ;
  assign \new_[8125]_  = (~\new_[9297]_  | ~\new_[17981]_ ) & (~\new_[9206]_  | ~\new_[18115]_ );
  assign \new_[8126]_  = (~\new_[8700]_  | ~\new_[19085]_ ) & (~\new_[9510]_  | ~\new_[18627]_ );
  assign \new_[8127]_  = (~\new_[9290]_  | ~\new_[19825]_ ) & (~\new_[9298]_  | ~\new_[19361]_ );
  assign \new_[8128]_  = ~\new_[8300]_ ;
  assign \new_[8129]_  = (~\new_[9290]_  | ~\new_[19546]_ ) & (~\new_[9298]_  | ~\new_[19580]_ );
  assign \new_[8130]_  = ~\new_[8302]_ ;
  assign \new_[8131]_  = ~\new_[8306]_ ;
  assign \new_[8132]_  = (~\new_[9297]_  | ~\new_[18818]_ ) & (~\new_[9206]_  | ~\new_[19658]_ );
  assign \new_[8133]_  = ~\new_[8308]_ ;
  assign \new_[8134]_  = (~\new_[9297]_  | ~\new_[19659]_ ) & (~\new_[9206]_  | ~\new_[18959]_ );
  assign \new_[8135]_  = (~\new_[19986]_  | ~\new_[18981]_ ) & (~\new_[20552]_  | ~\new_[19065]_ );
  assign \new_[8136]_  = ~\new_[8311]_ ;
  assign \new_[8137]_  = ~\new_[8314]_ ;
  assign \new_[8138]_  = (~\new_[9297]_  | ~\new_[18444]_ ) & (~\new_[9206]_  | ~\new_[18790]_ );
  assign \new_[8139]_  = (~\new_[9295]_  | ~\new_[18983]_ ) & (~\new_[9510]_  | ~\new_[19372]_ );
  assign \new_[8140]_  = ~\new_[8317]_ ;
  assign \new_[8141]_  = (~\new_[9290]_  | ~\new_[18633]_ ) & (~\new_[9509]_  | ~\new_[17877]_ );
  assign \new_[8142]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][2] ;
  assign \new_[8143]_  = (~\new_[9297]_  | ~\new_[19206]_ ) & (~\new_[9503]_  | ~\new_[18469]_ );
  assign \new_[8144]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][6] ;
  assign \new_[8145]_  = (~\new_[8700]_  | ~\new_[19371]_ ) & (~\new_[9510]_  | ~\new_[18404]_ );
  assign \new_[8146]_  = ~\new_[8321]_ ;
  assign \new_[8147]_  = (~\new_[8700]_  | ~\new_[18567]_ ) & (~\new_[9510]_  | ~\new_[18351]_ );
  assign \new_[8148]_  = (~\new_[9290]_  | ~\new_[18537]_ ) & (~\new_[9509]_  | ~\new_[18614]_ );
  assign \new_[8149]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][5] ;
  assign \new_[8150]_  = ~\new_[16229]_  | ~\new_[20479]_  | ~\new_[8549]_  | ~\new_[9829]_ ;
  assign \new_[8151]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][34] ;
  assign \new_[8152]_  = ~\new_[8328]_ ;
  assign \new_[8153]_  = (~\new_[9297]_  | ~\new_[19189]_ ) & (~\new_[9503]_  | ~\new_[19018]_ );
  assign \new_[8154]_  = (~\new_[9295]_  | ~\new_[18381]_ ) & (~\new_[9510]_  | ~\new_[18707]_ );
  assign \new_[8155]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][25] ;
  assign \new_[8156]_  = (~\new_[9290]_  | ~\new_[19113]_ ) & (~\new_[9509]_  | ~\new_[18667]_ );
  assign \new_[8157]_  = ~\new_[8333]_ ;
  assign \new_[8158]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][14] ;
  assign \new_[8159]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][25] ;
  assign \new_[8160]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][2] ;
  assign \new_[8161]_  = (~\new_[19986]_  | ~\new_[19693]_ ) & (~\new_[20552]_  | ~\new_[18103]_ );
  assign \new_[8162]_  = ~\new_[8344]_ ;
  assign \new_[8163]_  = (~\new_[9297]_  | ~\new_[19337]_ ) & (~\new_[9206]_  | ~\new_[19056]_ );
  assign \new_[8164]_  = ~\new_[8345]_ ;
  assign \new_[8165]_  = (~\new_[9297]_  | ~\new_[18578]_ ) & (~\new_[9206]_  | ~\new_[19612]_ );
  assign \new_[8166]_  = ~\new_[8348]_ ;
  assign \new_[8167]_  = (~\new_[9292]_  | ~\new_[19680]_ ) & (~\new_[20551]_  | ~\new_[19386]_ );
  assign \new_[8168]_  = (~\new_[9204]_  | ~\new_[19594]_ ) & (~\new_[9510]_  | ~\new_[17815]_ );
  assign \new_[8169]_  = (~\new_[9500]_  | ~\new_[19180]_ ) & (~\new_[9203]_  | ~\new_[18657]_ );
  assign \new_[8170]_  = (~\new_[9502]_  | ~\new_[18108]_ ) & (~\new_[9208]_  | ~\new_[19687]_ );
  assign \new_[8171]_  = ~\new_[8354]_ ;
  assign \new_[8172]_  = (~\new_[9290]_  | ~\new_[19870]_ ) & (~\new_[9298]_  | ~\new_[18412]_ );
  assign \new_[8173]_  = (~\new_[20012]_  | ~\new_[19063]_ ) & (~\new_[20518]_  | ~\new_[18332]_ );
  assign \new_[8174]_  = (~\new_[9500]_  | ~\new_[19336]_ ) & (~\new_[9203]_  | ~\new_[18976]_ );
  assign \new_[8175]_  = (~\new_[9204]_  | ~\new_[18676]_ ) & (~\new_[9303]_  | ~\new_[18665]_ );
  assign \new_[8176]_  = (~\new_[9502]_  | ~\new_[17967]_ ) & (~\new_[9208]_  | ~\new_[17852]_ );
  assign \new_[8177]_  = (~\new_[9500]_  | ~\new_[18701]_ ) & (~\new_[9203]_  | ~\new_[19626]_ );
  assign \new_[8178]_  = (~\new_[9204]_  | ~\new_[18544]_ ) & (~\new_[9303]_  | ~\new_[18499]_ );
  assign \new_[8179]_  = (~\new_[9204]_  | ~\new_[18886]_ ) & (~\new_[9303]_  | ~\new_[18475]_ );
  assign \new_[8180]_  = (~\new_[9502]_  | ~\new_[17943]_ ) & (~\new_[9208]_  | ~\new_[18492]_ );
  assign \new_[8181]_  = (~\new_[9204]_  | ~\new_[18186]_ ) & (~\new_[9302]_  | ~\new_[17823]_ );
  assign \new_[8182]_  = (~\new_[9502]_  | ~\new_[18695]_ ) & (~\new_[9208]_  | ~\new_[18287]_ );
  assign \new_[8183]_  = ~\new_[8368]_ ;
  assign \new_[8184]_  = (~\new_[9204]_  | ~\new_[18297]_ ) & (~\new_[9303]_  | ~\new_[18459]_ );
  assign \new_[8185]_  = (~\new_[9500]_  | ~\new_[18124]_ ) & (~\new_[9203]_  | ~\new_[18421]_ );
  assign \new_[8186]_  = (~\new_[9295]_  | ~\new_[18153]_ ) & (~\new_[9510]_  | ~\new_[18335]_ );
  assign \new_[8187]_  = ~\new_[8370]_ ;
  assign \new_[8188]_  = (~\new_[9290]_  | ~\new_[18089]_ ) & (~\new_[9299]_  | ~\new_[18184]_ );
  assign \new_[8189]_  = (~\new_[9292]_  | ~\new_[18758]_ ) & (~\new_[20551]_  | ~\new_[19025]_ );
  assign \new_[8190]_  = (~\new_[20012]_  | ~\new_[19454]_ ) & (~\new_[20518]_  | ~\new_[19655]_ );
  assign \new_[8191]_  = ~\new_[8373]_ ;
  assign \new_[8192]_  = (~\new_[9204]_  | ~\new_[19404]_ ) & (~\new_[9510]_  | ~\new_[18322]_ );
  assign \new_[8193]_  = (~\new_[9500]_  | ~\new_[18457]_ ) & (~\new_[9203]_  | ~\new_[19846]_ );
  assign \new_[8194]_  = (~\new_[9204]_  | ~\new_[18112]_ ) & (~\new_[9302]_  | ~\new_[18528]_ );
  assign \new_[8195]_  = ~\new_[8380]_ ;
  assign \new_[8196]_  = (~\new_[9204]_  | ~\new_[19441]_ ) & (~\new_[9303]_  | ~\new_[18945]_ );
  assign \new_[8197]_  = ~\new_[8384]_ ;
  assign \new_[8198]_  = (~\new_[9290]_  | ~\new_[18820]_ ) & (~\new_[9299]_  | ~\new_[17945]_ );
  assign \new_[8199]_  = (~\new_[20012]_  | ~\new_[19406]_ ) & (~\new_[20518]_  | ~\new_[18311]_ );
  assign \new_[8200]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0] ;
  assign \new_[8201]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0] ;
  assign \new_[8202]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1] ;
  assign \new_[8203]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2] ;
  assign \new_[8204]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[0] ;
  assign \new_[8205]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[10] ;
  assign \new_[8206]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[11] ;
  assign \new_[8207]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[13] ;
  assign \new_[8208]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[15] ;
  assign \new_[8209]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[16] ;
  assign \new_[8210]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[17] ;
  assign \new_[8211]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[19] ;
  assign \new_[8212]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[1] ;
  assign \new_[8213]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[20] ;
  assign \new_[8214]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[23] ;
  assign \new_[8215]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[24] ;
  assign \new_[8216]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[26] ;
  assign \new_[8217]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[27] ;
  assign \new_[8218]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[28] ;
  assign \new_[8219]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[30] ;
  assign \new_[8220]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[31] ;
  assign \new_[8221]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[7] ;
  assign \new_[8222]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[8] ;
  assign \new_[8223]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[9] ;
  assign \new_[8224]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1] ;
  assign n17435 = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[0] ;
  assign \new_[8226]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0] ;
  assign n5495 = \new_[9217]_  ? \new_[9698]_  : \new_[18879]_ ;
  assign n5500 = \new_[9218]_  ? \new_[9730]_  : \new_[19870]_ ;
  assign n5510 = \new_[9219]_  ? \new_[9660]_  : \new_[17815]_ ;
  assign n5505 = \new_[9220]_  ? \new_[9699]_  : \new_[19852]_ ;
  assign n5515 = \new_[9221]_  ? \new_[9663]_  : \new_[19687]_ ;
  assign n5520 = \new_[9222]_  ? \new_[9669]_  : \new_[19002]_ ;
  assign n5525 = \new_[9223]_  ? \new_[9661]_  : \new_[18108]_ ;
  assign n5650 = \new_[9224]_  ? \new_[9743]_  : \new_[19380]_ ;
  assign n5530 = \new_[9225]_  ? \new_[9750]_  : \new_[18982]_ ;
  assign n5535 = \new_[9226]_  ? \new_[9660]_  : \new_[18151]_ ;
  assign n5545 = \new_[9227]_  ? \new_[9739]_  : \new_[19052]_ ;
  assign n5540 = \new_[9228]_  ? \new_[9751]_  : \new_[18412]_ ;
  assign n5550 = \new_[9233]_  ? \new_[9749]_  : \new_[19032]_ ;
  assign n5635 = \new_[9234]_  ? \new_[9707]_  : \new_[18332]_ ;
  assign \new_[8241]_  = ~\new_[19914]_ ;
  assign \new_[8242]_  = ~\new_[20074]_ ;
  assign n5555 = \new_[9235]_  ? \new_[9698]_  : \new_[19254]_ ;
  assign n5630 = \new_[9236]_  ? \new_[9665]_  : \new_[18040]_ ;
  assign n5560 = \new_[9237]_  ? \new_[9748]_  : \new_[19615]_ ;
  assign n5625 = \new_[9238]_  ? \new_[9730]_  : \new_[18540]_ ;
  assign n5565 = \new_[9240]_  ? \new_[9660]_  : \new_[19594]_ ;
  assign n5620 = \new_[9253]_  ? \new_[9669]_  : \new_[18553]_ ;
  assign n5570 = \new_[9241]_  ? \new_[9724]_  : \new_[18954]_ ;
  assign n5490 = \new_[9242]_  ? \new_[9730]_  : \new_[18640]_ ;
  assign n5575 = \new_[9243]_  ? \new_[9733]_  : \new_[18657]_ ;
  assign n5580 = \new_[9244]_  ? \new_[9698]_  : \new_[18988]_ ;
  assign n5585 = \new_[9245]_  ? \new_[9733]_  : \new_[19180]_ ;
  assign n5590 = \new_[9246]_  ? \new_[9698]_  : \new_[19449]_ ;
  assign n5595 = \new_[9247]_  ? \new_[9669]_  : \new_[18264]_ ;
  assign n5600 = \new_[9248]_  ? \new_[9661]_  : \new_[19063]_ ;
  assign n5605 = \new_[9249]_  ? \new_[9721]_  : \new_[19227]_ ;
  assign n5645 = \new_[9250]_  ? \new_[9663]_  : \new_[18548]_ ;
  assign n5610 = \new_[9251]_  ? \new_[9699]_  : \new_[19822]_ ;
  assign n5640 = \new_[9252]_  ? \new_[9666]_  : \new_[19080]_ ;
  assign \new_[8261]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[3] ;
  assign \new_[8262]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[29] ;
  assign \new_[8263]_  = ~\new_[9829]_  | ~\new_[17510]_  | ~\new_[10328]_  | ~\new_[9493]_ ;
  assign \new_[8264]_  = (~\new_[20493]_  | ~\new_[19811]_ ) & (~\new_[9187]_  | ~\new_[17924]_ );
  assign \new_[8265]_  = (~\new_[20493]_  | ~\new_[19138]_ ) & (~\new_[9187]_  | ~\new_[18203]_ );
  assign \new_[8266]_  = (~\new_[20493]_  | ~\new_[19266]_ ) & (~\new_[9187]_  | ~\new_[19026]_ );
  assign n5615 = \new_[19874]_  & \new_[10949]_ ;
  assign \new_[8268]_  = (~\new_[20493]_  | ~\new_[19560]_ ) & (~\new_[9187]_  | ~\new_[19818]_ );
  assign \new_[8269]_  = (~\new_[20493]_  | ~\new_[19806]_ ) & (~\new_[9187]_  | ~\new_[18323]_ );
  assign \new_[8270]_  = (~\new_[20493]_  | ~\new_[18157]_ ) & (~\new_[9187]_  | ~\new_[19334]_ );
  assign \new_[8271]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[18] ;
  assign \new_[8272]_  = (~\new_[20493]_  | ~\new_[19724]_ ) & (~\new_[9187]_  | ~\new_[19815]_ );
  assign \new_[8273]_  = (~\new_[20493]_  | ~\new_[19162]_ ) & (~\new_[9187]_  | ~\new_[18284]_ );
  assign \new_[8274]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[21] ;
  assign \new_[8275]_  = ~\new_[8556]_ ;
  assign \new_[8276]_  = ~\new_[8559]_ ;
  assign \new_[8277]_  = ~\new_[20457]_ ;
  assign \new_[8278]_  = ~\new_[20457]_ ;
  assign \new_[8279]_  = ~\new_[20457]_ ;
  assign \new_[8280]_  = ~\new_[8560]_ ;
  assign \new_[8281]_  = ~\new_[20322]_ ;
  assign \new_[8282]_  = ~\new_[8562]_ ;
  assign \new_[8283]_  = ~\new_[8563]_ ;
  assign \new_[8284]_  = \new_[8565]_ ;
  assign \new_[8285]_  = \new_[8565]_ ;
  assign \new_[8286]_  = ~\new_[8565]_ ;
  assign \new_[8287]_  = ~\new_[20144]_ ;
  assign \new_[8288]_  = ~\new_[8566]_ ;
  assign \new_[8289]_  = ~\new_[8567]_ ;
  assign \new_[8290]_  = ~\new_[20343]_ ;
  assign \new_[8291]_  = ~\new_[8571]_ ;
  assign \new_[8292]_  = (~\new_[9500]_  | ~\new_[18718]_ ) & (~\new_[9203]_  | ~\new_[18192]_ );
  assign \new_[8293]_  = (~\new_[9204]_  | ~\new_[18070]_ ) & (~\new_[9303]_  | ~\new_[19537]_ );
  assign \new_[8294]_  = (~\new_[9502]_  | ~\new_[18526]_ ) & (~\new_[9208]_  | ~\new_[19625]_ );
  assign \new_[8295]_  = (~\new_[9202]_  | ~\new_[17911]_ ) & (~\new_[20518]_  | ~\new_[19425]_ );
  assign \new_[8296]_  = (~\new_[9204]_  | ~\new_[18738]_ ) & (~\new_[9302]_  | ~\new_[18893]_ );
  assign \new_[8297]_  = ~\new_[8590]_ ;
  assign \new_[8298]_  = (~\new_[9202]_  | ~\new_[18604]_ ) & (~\new_[20518]_  | ~\new_[19332]_ );
  assign \new_[8299]_  = (~\new_[9292]_  | ~\new_[19421]_ ) & (~\new_[20551]_  | ~\new_[17990]_ );
  assign \new_[8300]_  = (~\new_[19986]_  | ~\new_[18303]_ ) & (~\new_[20552]_  | ~\new_[18301]_ );
  assign \new_[8301]_  = (~\new_[9202]_  | ~\new_[19288]_ ) & (~\new_[20518]_  | ~\new_[19519]_ );
  assign \new_[8302]_  = (~\new_[9497]_  | ~\new_[18581]_ ) & (~\new_[9207]_  | ~\new_[19053]_ );
  assign \new_[8303]_  = (~\new_[9290]_  | ~\new_[18876]_ ) & (~\new_[9299]_  | ~\new_[18359]_ );
  assign \new_[8304]_  = (~\new_[9292]_  | ~\new_[18077]_ ) & (~\new_[20551]_  | ~\new_[19490]_ );
  assign \new_[8305]_  = (~\new_[20012]_  | ~\new_[19249]_ ) & (~\new_[20518]_  | ~\new_[17976]_ );
  assign \new_[8306]_  = (~\new_[9500]_  | ~\new_[18388]_ ) & (~\new_[9203]_  | ~\new_[18071]_ );
  assign \new_[8307]_  = (~\new_[9204]_  | ~\new_[19460]_ ) & (~\new_[9510]_  | ~\new_[18342]_ );
  assign \new_[8308]_  = (~\new_[9204]_  | ~\new_[17901]_ ) & (~\new_[9302]_  | ~\new_[19036]_ );
  assign \new_[8309]_  = (~\new_[9500]_  | ~\new_[19383]_ ) & (~\new_[9203]_  | ~\new_[19014]_ );
  assign \new_[8310]_  = (~\new_[9295]_  | ~\new_[18687]_ ) & (~\new_[9510]_  | ~\new_[19251]_ );
  assign \new_[8311]_  = (~\new_[19986]_  | ~\new_[19697]_ ) & (~\new_[20552]_  | ~\new_[19699]_ );
  assign \new_[8312]_  = (~\new_[9290]_  | ~\new_[18720]_ ) & (~\new_[9299]_  | ~\new_[18195]_ );
  assign \new_[8313]_  = (~\new_[20012]_  | ~\new_[18513]_ ) & (~\new_[20518]_  | ~\new_[18030]_ );
  assign \new_[8314]_  = (~\new_[9502]_  | ~\new_[18140]_ ) & (~\new_[9511]_  | ~\new_[19260]_ );
  assign \new_[8315]_  = (~\new_[9500]_  | ~\new_[18401]_ ) & (~\new_[9203]_  | ~\new_[19753]_ );
  assign \new_[8316]_  = (~\new_[9204]_  | ~\new_[18601]_ ) & (~\new_[9303]_  | ~\new_[18557]_ );
  assign \new_[8317]_  = (~\new_[9497]_  | ~\new_[18384]_ ) & (~\new_[9207]_  | ~\new_[18794]_ );
  assign \new_[8318]_  = (~\new_[9292]_  | ~\new_[19087]_ ) & (~\new_[20551]_  | ~\new_[18722]_ );
  assign \new_[8319]_  = (~\new_[20012]_  | ~\new_[19338]_ ) & (~\new_[20518]_  | ~\new_[17897]_ );
  assign \new_[8320]_  = (~\new_[9204]_  | ~\new_[18975]_ ) & (~\new_[9510]_  | ~\new_[18723]_ );
  assign \new_[8321]_  = (~\new_[19986]_  | ~\new_[18234]_ ) & (~\new_[20552]_  | ~\new_[17833]_ );
  assign \new_[8322]_  = (~\new_[9202]_  | ~\new_[18007]_ ) & (~\new_[20518]_  | ~\new_[18608]_ );
  assign \new_[8323]_  = (~\new_[19999]_  | ~\new_[18769]_ ) & (~\new_[20001]_  | ~\new_[19529]_ );
  assign \new_[8324]_  = (~\new_[9290]_  | ~\new_[19775]_ ) & (~\new_[9299]_  | ~\new_[19418]_ );
  assign \new_[8325]_  = (~\new_[19999]_  | ~\new_[18585]_ ) & (~\new_[20001]_  | ~\new_[19066]_ );
  assign \new_[8326]_  = (~\new_[9292]_  | ~\new_[17973]_ ) & (~\new_[20552]_  | ~\new_[19086]_ );
  assign \new_[8327]_  = ~\new_[8634]_ ;
  assign \new_[8328]_  = (~\new_[9204]_  | ~\new_[18434]_ ) & (~\new_[9510]_  | ~\new_[19630]_ );
  assign \new_[8329]_  = (~\new_[9502]_  | ~\new_[18295]_ ) & (~\new_[9208]_  | ~\new_[17903]_ );
  assign \new_[8330]_  = (~\new_[9500]_  | ~\new_[19755]_ ) & (~\new_[9203]_  | ~\new_[18978]_ );
  assign \new_[8331]_  = (~\new_[9202]_  | ~\new_[17949]_ ) & (~\new_[20518]_  | ~\new_[19645]_ );
  assign \new_[8332]_  = (~\new_[9292]_  | ~\new_[18621]_ ) & (~\new_[20552]_  | ~\new_[19757]_ );
  assign \new_[8333]_  = (~\new_[19986]_  | ~\new_[19057]_ ) & (~\new_[20552]_  | ~\new_[19214]_ );
  assign \new_[8334]_  = (~\new_[9290]_  | ~\new_[19858]_ ) & (~\new_[9298]_  | ~\new_[18986]_ );
  assign \new_[8335]_  = (~\new_[9202]_  | ~\new_[17939]_ ) & (~\new_[20518]_  | ~\new_[19236]_ );
  assign \new_[8336]_  = (~\new_[19999]_  | ~\new_[19205]_ ) & (~\new_[20001]_  | ~\new_[18341]_ );
  assign \new_[8337]_  = (~\new_[9295]_  | ~\new_[19101]_ ) & (~\new_[9510]_  | ~\new_[17895]_ );
  assign \new_[8338]_  = ~\new_[8642]_ ;
  assign \new_[8339]_  = (~\new_[9290]_  | ~\new_[18668]_ ) & (~\new_[9299]_  | ~\new_[19787]_ );
  assign \new_[8340]_  = (~\new_[9292]_  | ~\new_[18326]_ ) & (~\new_[20552]_  | ~\new_[18753]_ );
  assign \new_[8341]_  = ~\new_[8646]_ ;
  assign \new_[8342]_  = (~\new_[9290]_  | ~\new_[18292]_ ) & (~\new_[9298]_  | ~\new_[19714]_ );
  assign \new_[8343]_  = (~\new_[19999]_  | ~\new_[19241]_ ) & (~\new_[20001]_  | ~\new_[18776]_ );
  assign \new_[8344]_  = (~\new_[9204]_  | ~\new_[18204]_ ) & (~\new_[9510]_  | ~\new_[18390]_ );
  assign \new_[8345]_  = (~\new_[9502]_  | ~\new_[19754]_ ) & (~\new_[9511]_  | ~\new_[18845]_ );
  assign \new_[8346]_  = (~\new_[9204]_  | ~\new_[19176]_ ) & (~\new_[9510]_  | ~\new_[19796]_ );
  assign \new_[8347]_  = (~\new_[9295]_  | ~\new_[18218]_ ) & (~\new_[9510]_  | ~\new_[19797]_ );
  assign \new_[8348]_  = (~\new_[9291]_  | ~\new_[18783]_ ) & (~\new_[20518]_  | ~\new_[19353]_ );
  assign \new_[8349]_  = (~\new_[19999]_  | ~\new_[18093]_ ) & (~\new_[9300]_  | ~\new_[19007]_ );
  assign \new_[8350]_  = (~\new_[9290]_  | ~\new_[18879]_ ) & (~\new_[9509]_  | ~\new_[19052]_ );
  assign \new_[8351]_  = (~\new_[19986]_  | ~\new_[19615]_ ) & (~\new_[20551]_  | ~\new_[18954]_ );
  assign \new_[8352]_  = (~\new_[9297]_  | ~\new_[18040]_ ) & (~\new_[9504]_  | ~\new_[19080]_ );
  assign \new_[8353]_  = (~\new_[9295]_  | ~\new_[18553]_ ) & (~\new_[9510]_  | ~\new_[19852]_ );
  assign \new_[8354]_  = (~\new_[9497]_  | ~\new_[18548]_ ) & (~\new_[9301]_  | ~\new_[18151]_ );
  assign \new_[8355]_  = (~\new_[9290]_  | ~\new_[18503]_ ) & (~\new_[9509]_  | ~\new_[19696]_ );
  assign \new_[8356]_  = (~\new_[19987]_  | ~\new_[18762]_ ) & (~\new_[20552]_  | ~\new_[19760]_ );
  assign \new_[8357]_  = (~\new_[9290]_  | ~\new_[18747]_ ) & (~\new_[9509]_  | ~\new_[19152]_ );
  assign \new_[8358]_  = (~\new_[19986]_  | ~\new_[19267]_ ) & (~\new_[20552]_  | ~\new_[18014]_ );
  assign \new_[8359]_  = (~\new_[9502]_  | ~\new_[17969]_ ) & (~\new_[9304]_  | ~\new_[19172]_ );
  assign \new_[8360]_  = (~\new_[19986]_  | ~\new_[19640]_ ) & (~\new_[20552]_  | ~\new_[18518]_ );
  assign \new_[8361]_  = (~\new_[9290]_  | ~\new_[18967]_ ) & (~\new_[9509]_  | ~\new_[19590]_ );
  assign \new_[8362]_  = (~\new_[9500]_  | ~\new_[18427]_ ) & (~\new_[9294]_  | ~\new_[18409]_ );
  assign \new_[8363]_  = (~\new_[9292]_  | ~\new_[18863]_ ) & (~\new_[20551]_  | ~\new_[19010]_ );
  assign \new_[8364]_  = (~\new_[9290]_  | ~\new_[19089]_ ) & (~\new_[9509]_  | ~\new_[18637]_ );
  assign \new_[8365]_  = (~\new_[9500]_  | ~\new_[18453]_ ) & (~\new_[9294]_  | ~\new_[18416]_ );
  assign \new_[8366]_  = (~\new_[9290]_  | ~\new_[18693]_ ) & (~\new_[9509]_  | ~\new_[17893]_ );
  assign \new_[8367]_  = (~\new_[19986]_  | ~\new_[18272]_ ) & (~\new_[20552]_  | ~\new_[19719]_ );
  assign \new_[8368]_  = (~\new_[9502]_  | ~\new_[18684]_ ) & (~\new_[9511]_  | ~\new_[18487]_ );
  assign \new_[8369]_  = (~\new_[9297]_  | ~\new_[18828]_ ) & (~\new_[9506]_  | ~\new_[19027]_ );
  assign \new_[8370]_  = (~\new_[9497]_  | ~\new_[19649]_ ) & (~\new_[9301]_  | ~\new_[18022]_ );
  assign \new_[8371]_  = (~\new_[9292]_  | ~\new_[18977]_ ) & (~\new_[20552]_  | ~\new_[18966]_ );
  assign \new_[8372]_  = (~\new_[9290]_  | ~\new_[18923]_ ) & (~\new_[9509]_  | ~\new_[18775]_ );
  assign \new_[8373]_  = (~\new_[9502]_  | ~\new_[19828]_ ) & (~\new_[9511]_  | ~\new_[19591]_ );
  assign \new_[8374]_  = (~\new_[19986]_  | ~\new_[19243]_ ) & (~\new_[20552]_  | ~\new_[19097]_ );
  assign \new_[8375]_  = (~\new_[9290]_  | ~\new_[18777]_ ) & (~\new_[9509]_  | ~\new_[18691]_ );
  assign \new_[8376]_  = (~\new_[9500]_  | ~\new_[17916]_ ) & (~\new_[9294]_  | ~\new_[18694]_ );
  assign \new_[8377]_  = (~\new_[9502]_  | ~\new_[18889]_ ) & (~\new_[9304]_  | ~\new_[18299]_ );
  assign \new_[8378]_  = (~\new_[9292]_  | ~\new_[18898]_ ) & (~\new_[20552]_  | ~\new_[19689]_ );
  assign \new_[8379]_  = (~\new_[9290]_  | ~\new_[18529]_ ) & (~\new_[9509]_  | ~\new_[19794]_ );
  assign \new_[8380]_  = (~\new_[9502]_  | ~\new_[19165]_ ) & (~\new_[9511]_  | ~\new_[19188]_ );
  assign \new_[8381]_  = (~\new_[9500]_  | ~\new_[17915]_ ) & (~\new_[9294]_  | ~\new_[19344]_ );
  assign \new_[8382]_  = (~\new_[9295]_  | ~\new_[19443]_ ) & (~\new_[9510]_  | ~\new_[18826]_ );
  assign \new_[8383]_  = (~\new_[9297]_  | ~\new_[18931]_ ) & (~\new_[9507]_  | ~\new_[19059]_ );
  assign \new_[8384]_  = (~\new_[9497]_  | ~\new_[19033]_ ) & (~\new_[9301]_  | ~\new_[19549]_ );
  assign \new_[8385]_  = \\pci_target_unit_pci_target_sm_c_state_reg[0] ;
  assign \new_[8386]_  = \\pci_target_unit_pci_target_sm_c_state_reg[1] ;
  assign \new_[8387]_  = \\pci_target_unit_pci_target_sm_c_state_reg[2] ;
  assign \new_[8388]_  = ~\new_[9307]_ ;
  assign \new_[8389]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2] ;
  assign \new_[8390]_  = \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0] ;
  assign \new_[8391]_  = \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1] ;
  assign \new_[8392]_  = \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3] ;
  assign n17450 = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[1] ;
  assign \new_[8394]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3] ;
  assign \new_[8395]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[0] ;
  assign \new_[8396]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[1] ;
  assign \new_[8397]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[2] ;
  assign \new_[8398]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[3] ;
  assign n17285 = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[2] ;
  assign \new_[8400]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][36] ;
  assign \new_[8401]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][36] ;
  assign n6220 = \new_[9316]_  ? \new_[9605]_  : \new_[18994]_ ;
  assign n6215 = \new_[9317]_  ? \new_[9660]_  : \new_[19546]_ ;
  assign n5690 = \new_[9318]_  ? \new_[9709]_  : \new_[19775]_ ;
  assign n5695 = \new_[9319]_  ? \new_[9699]_  : \new_[19809]_ ;
  assign n6130 = \new_[9320]_  ? \new_[9669]_  : \new_[18511]_ ;
  assign n6200 = \new_[9311]_  ? \new_[9737]_  : \new_[18503]_ ;
  assign n5700 = \new_[9321]_  ? \new_[9742]_  : \new_[18693]_ ;
  assign n5705 = \new_[9322]_  ? \new_[9735]_  : \new_[18089]_ ;
  assign n6190 = \new_[9323]_  ? \new_[9699]_  : \new_[18923]_ ;
  assign n6180 = \new_[9324]_  ? \new_[9661]_  : \new_[18893]_ ;
  assign n5710 = \new_[9325]_  ? \new_[9736]_  : \new_[18939]_ ;
  assign n5715 = \new_[9326]_  ? \new_[9669]_  : \new_[18404]_ ;
  assign n6160 = \new_[9327]_  ? \new_[9661]_  : \new_[19630]_ ;
  assign n5720 = \new_[9328]_  ? \new_[9660]_  : \new_[18390]_ ;
  assign n6140 = \new_[9312]_  ? \new_[9669]_  : \new_[18665]_ ;
  assign n5730 = \new_[9329]_  ? \new_[9610]_  : \new_[18459]_ ;
  assign n5725 = \new_[9330]_  ? \new_[9738]_  : \new_[18335]_ ;
  assign n6120 = \new_[9331]_  ? \new_[9730]_  : \new_[18322]_ ;
  assign n5735 = \new_[9332]_  ? \new_[9667]_  : \new_[19125]_ ;
  assign n6105 = \new_[9333]_  ? \new_[9745]_  : \new_[19257]_ ;
  assign n5740 = \new_[9334]_  ? \new_[9726]_  : \new_[18851]_ ;
  assign n6085 = \new_[9335]_  ? \new_[9663]_  : \new_[17903]_ ;
  assign n5745 = \new_[9336]_  ? \new_[9725]_  : \new_[18696]_ ;
  assign n5750 = \new_[9313]_  ? \new_[9669]_  : \new_[17852]_ ;
  assign n5755 = \new_[9338]_  ? \new_[9613]_  : \new_[18685]_ ;
  assign n6065 = \new_[9337]_  ? \new_[9661]_  : \new_[18487]_ ;
  assign n6050 = \new_[9339]_  ? \new_[9714]_  : \new_[19591]_ ;
  assign n5760 = \new_[9340]_  ? \new_[9698]_  : \new_[19331]_ ;
  assign n6045 = \new_[9341]_  ? \new_[9730]_  : \new_[18090]_ ;
  assign n6300 = \new_[9342]_  ? \new_[9755]_  : \new_[18907]_ ;
  assign n6370 = \new_[9343]_  ? \new_[9740]_  : \new_[18295]_ ;
  assign n6375 = \new_[9344]_  ? \new_[9699]_  : \new_[18158]_ ;
  assign n5765 = \new_[9314]_  ? \new_[9733]_  : \new_[17967]_ ;
  assign n5770 = \new_[9345]_  ? \new_[9711]_  : \new_[18684]_ ;
  assign n6350 = \new_[9346]_  ? \new_[9611]_  : \new_[18847]_ ;
  assign n5775 = \new_[9347]_  ? \new_[9660]_  : \new_[19828]_ ;
  assign n5780 = \new_[9348]_  ? \new_[9737]_  : \new_[18058]_ ;
  assign n5785 = \new_[9349]_  ? \new_[9737]_  : \new_[19440]_ ;
  assign n6335 = \new_[9350]_  ? \new_[9746]_  : \new_[19529]_ ;
  assign n6305 = \new_[9351]_  ? \new_[9667]_  : \new_[18724]_ ;
  assign n6330 = \new_[9352]_  ? \new_[9669]_  : \new_[19245]_ ;
  assign n6320 = \new_[9315]_  ? \new_[9728]_  : \new_[19378]_ ;
  assign n5790 = \new_[9353]_  ? \new_[9731]_  : \new_[18054]_ ;
  assign n5795 = \new_[9354]_  ? \new_[9663]_  : \new_[18022]_ ;
  assign n5680 = ~\new_[9493]_  | (~wbs_stb_i & ~\new_[17473]_ );
  assign n6325 = \new_[9355]_  ? \new_[9757]_  : \new_[19477]_ ;
  assign n6315 = \new_[9356]_  ? \new_[9726]_  : \new_[18205]_ ;
  assign n6310 = \new_[9357]_  ? \new_[9660]_  : \new_[19580]_ ;
  assign n5800 = \new_[9358]_  ? \new_[9715]_  : \new_[19418]_ ;
  assign n5805 = \new_[9359]_  ? \new_[9751]_  : \new_[18639]_ ;
  assign n6295 = \new_[9360]_  ? \new_[9736]_  : \new_[19793]_ ;
  assign n6290 = \new_[9310]_  ? \new_[9739]_  : \new_[19696]_ ;
  assign n5810 = \new_[9361]_  ? \new_[9669]_  : \new_[17893]_ ;
  assign n5815 = \new_[9362]_  ? \new_[9613]_  : \new_[18184]_ ;
  assign n6285 = \new_[9363]_  ? \new_[9669]_  : \new_[18775]_ ;
  assign n5820 = \new_[9365]_  ? \new_[9730]_  : \new_[18343]_ ;
  assign n5825 = \new_[9366]_  ? \new_[9758]_  : \new_[19519]_ ;
  assign n5830 = \new_[9367]_  ? \new_[9667]_  : \new_[18608]_ ;
  assign n6280 = \new_[9368]_  ? \new_[9605]_  : \new_[18460]_ ;
  assign n5835 = \new_[9369]_  ? \new_[9730]_  : \new_[18877]_ ;
  assign n5840 = \new_[9370]_  ? \new_[9733]_  : \new_[18921]_ ;
  assign n5850 = \new_[9371]_  ? \new_[9660]_  : \new_[19655]_ ;
  assign n5845 = \new_[9372]_  ? \new_[9733]_  : \new_[19817]_ ;
  assign n5855 = \new_[9373]_  ? \new_[9669]_  : \new_[18741]_ ;
  assign n6275 = \new_[9374]_  ? \new_[9703]_  : \new_[19191]_ ;
  assign n5860 = \new_[9375]_  ? \new_[9740]_  : \new_[19656]_ ;
  assign n6270 = \new_[9376]_  ? \new_[9661]_  : \new_[18978]_ ;
  assign n5865 = \new_[9377]_  ? \new_[9666]_  : \new_[18506]_ ;
  assign n5870 = \new_[9378]_  ? \new_[9663]_  : \new_[18421]_ ;
  assign n5875 = \new_[9379]_  ? \new_[9753]_  : \new_[19094]_ ;
  assign n6265 = \new_[9380]_  ? \new_[9663]_  : \new_[19846]_ ;
  assign n5880 = \new_[9381]_  ? \new_[9743]_  : \new_[18541]_ ;
  assign n6260 = \new_[9382]_  ? \new_[9745]_  : \new_[19494]_ ;
  assign n6255 = \new_[9383]_  ? \new_[9610]_  : \new_[17928]_ ;
  assign n6250 = \new_[9384]_  ? \new_[9661]_  : \new_[19755]_ ;
  assign n6245 = \new_[9385]_  ? \new_[9669]_  : \new_[18440]_ ;
  assign n6235 = \new_[9364]_  ? \new_[9719]_  : \new_[18124]_ ;
  assign n5885 = \new_[9386]_  ? \new_[9704]_  : \new_[17918]_ ;
  assign n6240 = \new_[9387]_  ? \new_[9661]_  : \new_[18457]_ ;
  assign n5890 = \new_[9388]_  ? \new_[9756]_  : \new_[19390]_ ;
  assign n6230 = \new_[9389]_  ? \new_[9756]_  : \new_[19288]_ ;
  assign n5895 = \new_[9390]_  ? \new_[9735]_  : \new_[18007]_ ;
  assign n6225 = \new_[9391]_  ? \new_[9746]_  : \new_[17944]_ ;
  assign n5900 = \new_[9392]_  ? \new_[9669]_  : \new_[19270]_ ;
  assign n5905 = \new_[9393]_  ? \new_[9669]_  : \new_[18171]_ ;
  assign n5910 = \new_[9394]_  ? \new_[9661]_  : \new_[19454]_ ;
  assign n6210 = \new_[9395]_  ? \new_[9669]_  : \new_[19569]_ ;
  assign n5915 = \new_[9396]_  ? \new_[9661]_  : \new_[18115]_ ;
  assign n6205 = \new_[9397]_  ? \new_[9730]_  : \new_[19313]_ ;
  assign n5920 = \new_[9398]_  ? \new_[9757]_  : \new_[19712]_ ;
  assign n6115 = \new_[9399]_  ? \new_[9745]_  : \new_[19018]_ ;
  assign n5925 = \new_[9400]_  ? \new_[9710]_  : \new_[19056]_ ;
  assign n5930 = \new_[9401]_  ? \new_[9730]_  : \new_[18666]_ ;
  assign n5935 = \new_[9402]_  ? \new_[9730]_  : \new_[19027]_ ;
  assign n6195 = \new_[9403]_  ? \new_[9731]_  : \new_[18554]_ ;
  assign n6170 = \new_[9407]_  ? \new_[9733]_  : \new_[18296]_ ;
  assign n5940 = \new_[9408]_  ? \new_[9660]_  : \new_[17981]_ ;
  assign n6185 = \new_[9409]_  ? \new_[9741]_  : \new_[19289]_ ;
  assign n6175 = \new_[9410]_  ? \new_[9605]_  : \new_[18057]_ ;
  assign n6145 = \new_[9411]_  ? \new_[9667]_  : \new_[19189]_ ;
  assign n6165 = \new_[9412]_  ? \new_[9713]_  : \new_[19337]_ ;
  assign n6150 = \new_[9413]_  ? \new_[9712]_  : \new_[18081]_ ;
  assign n6155 = \new_[9414]_  ? \new_[9698]_  : \new_[18245]_ ;
  assign n5945 = \new_[9415]_  ? \new_[9736]_  : \new_[18828]_ ;
  assign n6125 = \new_[9416]_  ? \new_[9607]_  : \new_[19181]_ ;
  assign n5950 = \new_[9417]_  ? \new_[9702]_  : \new_[19842]_ ;
  assign n6135 = \new_[9418]_  ? \new_[9709]_  : \new_[18303]_ ;
  assign n6095 = \new_[9419]_  ? \new_[9661]_  : \new_[18234]_ ;
  assign n6110 = \new_[9420]_  ? \new_[9607]_  : \new_[18072]_ ;
  assign n6100 = \new_[9445]_  ? \new_[9669]_  : \new_[19091]_ ;
  assign n5955 = \new_[9421]_  ? \new_[9751]_  : \new_[18762]_ ;
  assign n6075 = \new_[9422]_  ? \new_[9730]_  : \new_[18272]_ ;
  assign n6090 = \new_[9423]_  ? \new_[9733]_  : \new_[18758]_ ;
  assign n5960 = \new_[9424]_  ? \new_[9727]_  : \new_[18977]_ ;
  assign n5965 = \new_[9425]_  ? \new_[9707]_  : \new_[18738]_ ;
  assign n6080 = \new_[9426]_  ? \new_[9663]_  : \new_[19823]_ ;
  assign n6070 = \new_[9427]_  ? \new_[9699]_  : \new_[19371]_ ;
  assign n6060 = \new_[9428]_  ? \new_[9720]_  : \new_[18434]_ ;
  assign n6055 = \new_[9429]_  ? \new_[9705]_  : \new_[18204]_ ;
  assign n6035 = \new_[9430]_  ? \new_[9698]_  : \new_[18676]_ ;
  assign n6040 = \new_[9431]_  ? \new_[9669]_  : \new_[18297]_ ;
  assign n5970 = \new_[9432]_  ? \new_[9745]_  : \new_[18153]_ ;
  assign n5975 = \new_[9433]_  ? \new_[9664]_  : \new_[19404]_ ;
  assign n5980 = \new_[9434]_  ? \new_[9750]_  : \new_[19242]_ ;
  assign n5685 = \new_[9435]_  ? \new_[9662]_  : \new_[18301]_ ;
  assign n5985 = \new_[9436]_  ? \new_[9706]_  : \new_[17833]_ ;
  assign n5675 = \new_[9437]_  ? \new_[9754]_  : \new_[17832]_ ;
  assign n5670 = \new_[9438]_  ? \new_[9730]_  : \new_[18759]_ ;
  assign n5990 = \new_[9439]_  ? \new_[9730]_  : \new_[19760]_ ;
  assign n5665 = \new_[9440]_  ? \new_[9668]_  : \new_[19719]_ ;
  assign n5660 = \new_[9441]_  ? \new_[9668]_  : \new_[19025]_ ;
  assign n5995 = \new_[9442]_  ? \new_[9611]_  : \new_[18966]_ ;
  assign n5655 = \new_[9404]_  ? \new_[9661]_  : \new_[18976]_ ;
  assign n6355 = \new_[9443]_  ? \new_[9720]_  : \new_[19336]_ ;
  assign n6000 = \new_[9444]_  ? \new_[9608]_  : \new_[18286]_ ;
  assign n6005 = \new_[9452]_  ? \new_[9669]_  : \new_[19662]_ ;
  assign n6365 = \new_[9446]_  ? \new_[9733]_  : \new_[19132]_ ;
  assign n6010 = \new_[9447]_  ? \new_[9699]_  : \new_[18769]_ ;
  assign n6360 = \new_[9448]_  ? \new_[9728]_  : \new_[19733]_ ;
  assign n6340 = \new_[9449]_  ? \new_[9670]_  : \new_[18618]_ ;
  assign n6015 = \new_[9406]_  ? \new_[9747]_  : \new_[19558]_ ;
  assign n6020 = \new_[9453]_  ? \new_[9733]_  : \new_[18873]_ ;
  assign n6025 = \new_[9450]_  ? \new_[9717]_  : \new_[19649]_ ;
  assign n6345 = \new_[9451]_  ? \new_[9699]_  : \new_[18402]_ ;
  assign n6030 = \new_[9405]_  ? \new_[9707]_  : \new_[18507]_ ;
  assign n17250 = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[3] ;
  assign \new_[8548]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2] ;
  assign \new_[8549]_  = ~\new_[10459]_  & (~\new_[16993]_  | ~\new_[9286]_ );
  assign \new_[8550]_  = \new_[6304]_  ? \new_[9286]_  : \new_[15380]_ ;
  assign \new_[8551]_  = \new_[6303]_  ? \new_[9286]_  : \new_[15628]_ ;
  assign \new_[8552]_  = \new_[6317]_  ? \new_[9286]_  : \new_[15610]_ ;
  assign \new_[8553]_  = \new_[6305]_  ? \new_[9567]_  : \new_[15157]_ ;
  assign \new_[8554]_  = \new_[6306]_  ? \new_[9286]_  : \new_[14974]_ ;
  assign \new_[8555]_  = \new_[6307]_  ? \new_[9286]_  : \new_[15250]_ ;
  assign \new_[8556]_  = ~\new_[9134]_ ;
  assign \new_[8557]_  = ~\new_[20335]_  | ~\new_[20390]_ ;
  assign \new_[8558]_  = \new_[6308]_  ? \new_[9567]_  : \new_[15238]_ ;
  assign \new_[8559]_  = ~\new_[9216]_  | ~\new_[20335]_ ;
  assign \new_[8560]_  = ~\new_[20459]_  | ~\new_[20390]_ ;
  assign \new_[8561]_  = \new_[6309]_  ? \new_[9286]_  : \new_[14986]_ ;
  assign \new_[8562]_  = ~\new_[20345]_  | ~\new_[20458]_ ;
  assign \new_[8563]_  = ~\new_[9216]_  | ~\new_[20323]_ ;
  assign \new_[8564]_  = \new_[6329]_  ? \new_[9286]_  : \new_[14193]_ ;
  assign \new_[8565]_  = ~\new_[9135]_ ;
  assign \new_[8566]_  = ~\new_[20345]_  | ~\new_[20390]_ ;
  assign \new_[8567]_  = ~\new_[20344]_  | ~\new_[20459]_ ;
  assign \new_[8568]_  = \new_[6310]_  ? \new_[9286]_  : \new_[15242]_ ;
  assign \new_[8569]_  = ~\new_[20345]_  | ~\new_[9216]_ ;
  assign \new_[8570]_  = \new_[6311]_  ? \new_[9286]_  : \new_[15243]_ ;
  assign \new_[8571]_  = ~\new_[9216]_  | ~\new_[20459]_ ;
  assign \new_[8572]_  = (~\new_[9290]_  | ~\new_[17925]_ ) & (~\new_[9509]_  | ~\new_[18705]_ );
  assign \new_[8573]_  = (~\new_[19986]_  | ~\new_[18484]_ ) & (~\new_[20552]_  | ~\new_[18034]_ );
  assign \new_[8574]_  = \new_[6312]_  ? \new_[9286]_  : \new_[15159]_ ;
  assign \new_[8575]_  = \new_[6328]_  ? \new_[9567]_  : \new_[14851]_ ;
  assign \new_[8576]_  = (~\new_[9297]_  | ~\new_[19103]_ ) & (~\new_[9506]_  | ~\new_[18164]_ );
  assign \new_[8577]_  = (~\new_[19999]_  | ~\new_[19600]_ ) & (~\new_[9300]_  | ~\new_[18811]_ );
  assign \new_[8578]_  = \new_[6313]_  ? \new_[9286]_  : \new_[15244]_ ;
  assign \new_[8579]_  = (~\new_[9297]_  | ~\new_[19079]_ ) & (~\new_[9505]_  | ~\new_[19223]_ );
  assign \new_[8580]_  = (~\new_[9291]_  | ~\new_[19106]_ ) & (~\new_[20518]_  | ~\new_[18354]_ );
  assign \new_[8581]_  = (~\new_[19999]_  | ~\new_[18929]_ ) & (~\new_[9300]_  | ~\new_[18857]_ );
  assign \new_[8582]_  = \new_[6314]_  ? \new_[9286]_  : \new_[15005]_ ;
  assign \new_[8583]_  = (~\new_[9290]_  | ~\new_[18994]_ ) & (~\new_[9509]_  | ~\new_[18205]_ );
  assign \new_[8584]_  = (~\new_[19986]_  | ~\new_[19842]_ ) & (~\new_[20552]_  | ~\new_[19242]_ );
  assign \new_[8585]_  = \new_[6315]_  ? \new_[9286]_  : \new_[14981]_ ;
  assign \new_[8586]_  = (~\new_[9500]_  | ~\new_[18541]_ ) & (~\new_[9294]_  | ~\new_[18741]_ );
  assign \new_[8587]_  = (~\new_[9502]_  | ~\new_[19331]_ ) & (~\new_[9304]_  | ~\new_[19125]_ );
  assign \new_[8588]_  = \new_[6552]_  ? \new_[9286]_  : \new_[13788]_ ;
  assign \new_[8589]_  = (~\new_[9297]_  | ~\new_[18257]_ ) & (~\new_[9507]_  | ~\new_[19665]_ );
  assign \new_[8590]_  = (~\new_[9497]_  | ~\new_[17807]_ ) & (~\new_[9301]_  | ~\new_[19179]_ );
  assign \new_[8591]_  = \new_[6316]_  ? \new_[9286]_  : \new_[14877]_ ;
  assign \new_[8592]_  = (~\new_[9297]_  | ~\new_[19289]_ ) & (~\new_[9504]_  | ~\new_[19313]_ );
  assign \new_[8593]_  = (~\new_[9295]_  | ~\new_[19823]_ ) & (~\new_[9510]_  | ~\new_[18939]_ );
  assign \new_[8594]_  = \new_[6326]_  ? \new_[9286]_  : \new_[14869]_ ;
  assign \new_[8595]_  = (~\new_[19999]_  | ~\new_[19132]_ ) & (~\new_[9300]_  | ~\new_[19440]_ );
  assign \new_[8596]_  = (~\new_[9297]_  | ~\new_[18655]_ ) & (~\new_[9504]_  | ~\new_[19545]_ );
  assign \new_[8597]_  = (~\new_[9295]_  | ~\new_[19300]_ ) & (~\new_[9510]_  | ~\new_[18324]_ );
  assign \new_[8598]_  = (~\new_[9286]_  & ~\new_[6318]_ ) | (~\new_[9493]_  & ~\new_[14195]_ );
  assign \new_[8599]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1] ;
  assign \new_[8600]_  = \new_[6319]_  ? \new_[9567]_  : \new_[13606]_ ;
  assign \new_[8601]_  = (~\new_[9292]_  | ~\new_[18905]_ ) & (~\new_[20552]_  | ~\new_[19749]_ );
  assign \new_[8602]_  = (~\new_[9290]_  | ~\new_[18654]_ ) & (~\new_[9509]_  | ~\new_[17806]_ );
  assign \new_[8603]_  = \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2] ;
  assign \new_[8604]_  = (~\new_[9502]_  | ~\new_[19648]_ ) & (~\new_[9304]_  | ~\new_[18191]_ );
  assign \new_[8605]_  = (~\new_[9286]_  & ~\new_[6320]_ ) | (~\new_[9493]_  & ~\new_[14210]_ );
  assign \new_[8606]_  = (~\new_[9292]_  | ~\new_[18064]_ ) & (~\new_[20551]_  | ~\new_[19518]_ );
  assign \new_[8607]_  = (~\new_[9290]_  | ~\new_[18930]_ ) & (~\new_[9509]_  | ~\new_[19230]_ );
  assign \new_[8608]_  = \new_[6321]_  ? \new_[9286]_  : \new_[17286]_ ;
  assign \new_[8609]_  = (~\new_[9502]_  | ~\new_[17886]_ ) & (~\new_[9304]_  | ~\new_[19263]_ );
  assign \new_[8610]_  = (~\new_[9297]_  | ~\new_[18504]_ ) & (~\new_[9505]_  | ~\new_[18516]_ );
  assign \new_[8611]_  = \new_[6553]_  ? \new_[9286]_  : \new_[16469]_ ;
  assign \new_[8612]_  = (~\new_[9297]_  | ~\new_[17879]_ ) & (~\new_[9503]_  | ~\new_[18571]_ );
  assign \new_[8613]_  = \new_[6322]_  ? \new_[9286]_  : \new_[15945]_ ;
  assign \new_[8614]_  = (~\new_[9295]_  | ~\new_[18964]_ ) & (~\new_[9510]_  | ~\new_[18135]_ );
  assign \new_[8615]_  = (~\new_[19999]_  | ~\new_[19867]_ ) & (~\new_[9300]_  | ~\new_[19611]_ );
  assign \new_[8616]_  = \new_[6323]_  ? \new_[9286]_  : \new_[15789]_ ;
  assign \new_[8617]_  = (~\new_[9290]_  | ~\new_[18443]_ ) & (~\new_[9509]_  | ~\new_[18029]_ );
  assign \new_[8618]_  = (~\new_[19986]_  | ~\new_[19566]_ ) & (~\new_[20551]_  | ~\new_[19543]_ );
  assign \new_[8619]_  = \new_[6324]_  ? \new_[9286]_  : \new_[15987]_ ;
  assign \new_[8620]_  = (~\new_[9297]_  | ~\new_[19495]_ ) & (~\new_[9506]_  | ~\new_[19006]_ );
  assign \new_[8621]_  = \new_[6551]_  ? \new_[9286]_  : \new_[15958]_ ;
  assign \new_[8622]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3] ;
  assign \new_[8623]_  = (~\new_[9290]_  | ~\new_[18366]_ ) & (~\new_[9509]_  | ~\new_[19767]_ );
  assign \new_[8624]_  = \new_[6325]_  ? \new_[9286]_  : \new_[15595]_ ;
  assign \new_[8625]_  = (~\new_[9292]_  | ~\new_[18878]_ ) & (~\new_[20551]_  | ~\new_[17834]_ );
  assign \new_[8626]_  = (~\new_[9502]_  | ~\new_[19279]_ ) & (~\new_[9304]_  | ~\new_[17942]_ );
  assign \new_[8627]_  = \new_[6554]_  ^ \new_[9286]_ ;
  assign \new_[8628]_  = (~\new_[9500]_  | ~\new_[17929]_ ) & (~\new_[9294]_  | ~\new_[19624]_ );
  assign \new_[8629]_  = (~\new_[9297]_  | ~\new_[18057]_ ) & (~\new_[9504]_  | ~\new_[19712]_ );
  assign \new_[8630]_  = (~\new_[9297]_  | ~\new_[18106]_ ) & (~\new_[9505]_  | ~\new_[19788]_ );
  assign \new_[8631]_  = (~\new_[9291]_  | ~\new_[18019]_ ) & (~\new_[20518]_  | ~\new_[18963]_ );
  assign \new_[8632]_  = (~\new_[9295]_  | ~\new_[18630]_ ) & (~\new_[9510]_  | ~\new_[19854]_ );
  assign \new_[8633]_  = (~\new_[9297]_  | ~\new_[18997]_ ) & (~\new_[9507]_  | ~\new_[19722]_ );
  assign \new_[8634]_  = (~\new_[9291]_  | ~\new_[17992]_ ) & (~\new_[20518]_  | ~\new_[19547]_ );
  assign \new_[8635]_  = (~\new_[9290]_  | ~\new_[19809]_ ) & (~\new_[9509]_  | ~\new_[18639]_ );
  assign \new_[8636]_  = (~\new_[9292]_  | ~\new_[18072]_ ) & (~\new_[20551]_  | ~\new_[17832]_ );
  assign \new_[8637]_  = (~\new_[9297]_  | ~\new_[19581]_ ) & (~\new_[9507]_  | ~\new_[19022]_ );
  assign \new_[8638]_  = (~\new_[19999]_  | ~\new_[18314]_ ) & (~\new_[9300]_  | ~\new_[19200]_ );
  assign \new_[8639]_  = (~\new_[9297]_  | ~\new_[18285]_ ) & (~\new_[9505]_  | ~\new_[19727]_ );
  assign \new_[8640]_  = (~\new_[9295]_  | ~\new_[19635]_ ) & (~\new_[9510]_  | ~\new_[18846]_ );
  assign \new_[8641]_  = (~\new_[9297]_  | ~\new_[18121]_ ) & (~\new_[9506]_  | ~\new_[18563]_ );
  assign \new_[8642]_  = (~\new_[9291]_  | ~\new_[19514]_ ) & (~\new_[20518]_  | ~\new_[18238]_ );
  assign \new_[8643]_  = (~\new_[19999]_  | ~\new_[19110]_ ) & (~\new_[9300]_  | ~\new_[18230]_ );
  assign \new_[8644]_  = (~\new_[9297]_  | ~\new_[19352]_ ) & (~\new_[9504]_  | ~\new_[19092]_ );
  assign \new_[8645]_  = (~\new_[9295]_  | ~\new_[18530]_ ) & (~\new_[9510]_  | ~\new_[18869]_ );
  assign \new_[8646]_  = (~\new_[9291]_  | ~\new_[17888]_ ) & (~\new_[20518]_  | ~\new_[17864]_ );
  assign \new_[8647]_  = (~\new_[9290]_  | ~\new_[18511]_ ) & (~\new_[9509]_  | ~\new_[19793]_ );
  assign \new_[8648]_  = (~\new_[19987]_  | ~\new_[19091]_ ) & (~\new_[20552]_  | ~\new_[18759]_ );
  assign \new_[8649]_  = (~\new_[9502]_  | ~\new_[18158]_ ) & (~\new_[9304]_  | ~\new_[18696]_ );
  assign \new_[8650]_  = (~\new_[9500]_  | ~\new_[18440]_ ) & (~\new_[9294]_  | ~\new_[18506]_ );
  assign \new_[8651]_  = (~\new_[9290]_  | ~\new_[17952]_ ) & (~\new_[9509]_  | ~\new_[19800]_ );
  assign \new_[8652]_  = (~\new_[9292]_  | ~\new_[19073]_ ) & (~\new_[20551]_  | ~\new_[17848]_ );
  assign \new_[8653]_  = (~\new_[9500]_  | ~\new_[19408]_ ) & (~\new_[9294]_  | ~\new_[19718]_ );
  assign \new_[8654]_  = (~\new_[9297]_  | ~\new_[17904]_ ) & (~\new_[9504]_  | ~\new_[18231]_ );
  assign \new_[8655]_  = (~\new_[9500]_  | ~\new_[17922]_ ) & (~\new_[9499]_  | ~\new_[19668]_ );
  assign \new_[8656]_  = (~\new_[20012]_  | ~\new_[18264]_ ) & (~\new_[20518]_  | ~\new_[19032]_ );
  assign \new_[8657]_  = (~\new_[9497]_  | ~\new_[19227]_ ) & (~\new_[19997]_  | ~\new_[18982]_ );
  assign \new_[8658]_  = (~\new_[9500]_  | ~\new_[19449]_ ) & (~\new_[9499]_  | ~\new_[18988]_ );
  assign \new_[8659]_  = (~\new_[9502]_  | ~\new_[19380]_ ) & (~\new_[9511]_  | ~\new_[19002]_ );
  assign \new_[8660]_  = (~\new_[20012]_  | ~\new_[18286]_ ) & (~\new_[20518]_  | ~\new_[18296]_ );
  assign \new_[8661]_  = (~\new_[19999]_  | ~\new_[19558]_ ) & (~\new_[19997]_  | ~\new_[19378]_ );
  assign \new_[8662]_  = (~\new_[20012]_  | ~\new_[17813]_ ) & (~\new_[20518]_  | ~\new_[18220]_ );
  assign \new_[8663]_  = (~\new_[19999]_  | ~\new_[18436]_ ) & (~\new_[19997]_  | ~\new_[18956]_ );
  assign \new_[8664]_  = (~\new_[20012]_  | ~\new_[18382]_ ) & (~\new_[20518]_  | ~\new_[19285]_ );
  assign \new_[8665]_  = (~\new_[9497]_  | ~\new_[19154]_ ) & (~\new_[19997]_  | ~\new_[19750]_ );
  assign \new_[8666]_  = (~\new_[9497]_  | ~\new_[19252]_ ) & (~\new_[19997]_  | ~\new_[18148]_ );
  assign \new_[8667]_  = (~\new_[20012]_  | ~\new_[17956]_ ) & (~\new_[20518]_  | ~\new_[18101]_ );
  assign \new_[8668]_  = (~\new_[9497]_  | ~\new_[18873]_ ) & (~\new_[19997]_  | ~\new_[18054]_ );
  assign \new_[8669]_  = (~\new_[20012]_  | ~\new_[18171]_ ) & (~\new_[20518]_  | ~\new_[18921]_ );
  assign \new_[8670]_  = (~\new_[9500]_  | ~\new_[17918]_ ) & (~\new_[9499]_  | ~\new_[19094]_ );
  assign \new_[8671]_  = (~\new_[9502]_  | ~\new_[18847]_ ) & (~\new_[9511]_  | ~\new_[18685]_ );
  assign \new_[8672]_  = (~\new_[20012]_  | ~\new_[19569]_ ) & (~\new_[20518]_  | ~\new_[19817]_ );
  assign \new_[8673]_  = (~\new_[19999]_  | ~\new_[18402]_ ) & (~\new_[19997]_  | ~\new_[19477]_ );
  assign \new_[8674]_  = (~\new_[9497]_  | ~\new_[18219]_ ) & (~\new_[19997]_  | ~\new_[17962]_ );
  assign \new_[8675]_  = (~\new_[20012]_  | ~\new_[18796]_ ) & (~\new_[20518]_  | ~\new_[18670]_ );
  assign \new_[8676]_  = (~\new_[9497]_  | ~\new_[19798]_ ) & (~\new_[19997]_  | ~\new_[17910]_ );
  assign \new_[8677]_  = (~\new_[20012]_  | ~\new_[18472]_ ) & (~\new_[20518]_  | ~\new_[18969]_ );
  assign \new_[8678]_  = (~\new_[9502]_  | ~\new_[18749]_ ) & (~\new_[9511]_  | ~\new_[18501]_ );
  assign \new_[8679]_  = (~\new_[9500]_  | ~\new_[19396]_ ) & (~\new_[9499]_  | ~\new_[19395]_ );
  assign n6380 = \new_[11344]_  ? \new_[16604]_  : \new_[9512]_ ;
  assign \new_[8681]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[0] ;
  assign \new_[8682]_  = ~\new_[9188]_ ;
  assign \new_[8683]_  = ~\new_[9189]_ ;
  assign \new_[8684]_  = ~\new_[9189]_ ;
  assign \new_[8685]_  = \new_[9239]_ ;
  assign \new_[8686]_  = \new_[9239]_ ;
  assign \new_[8687]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3] ;
  assign \new_[8688]_  = ~\\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[1] ;
  assign \new_[8689]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[12] ;
  assign \new_[8690]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[22] ;
  assign \new_[8691]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[2] ;
  assign \new_[8692]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[5] ;
  assign \new_[8693]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[4] ;
  assign \new_[8694]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][36] ;
  assign \new_[8695]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][36] ;
  assign \new_[8696]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][36] ;
  assign \new_[8697]_  = ~\new_[9189]_ ;
  assign \new_[8698]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[25] ;
  assign n6385 = ~\new_[9288]_  | (~\new_[16604]_  & ~\new_[11344]_ );
  assign \new_[8700]_  = ~\new_[9205]_ ;
  assign n6390 = \new_[10876]_  ? \new_[16604]_  : \new_[9529]_ ;
  assign n6395 = \new_[11345]_  ? \new_[16604]_  : \new_[9530]_ ;
  assign \new_[8703]_  = ~\new_[9462]_  & (~\new_[18220]_  | ~\new_[16662]_ );
  assign \new_[8704]_  = ~\new_[9463]_  & (~\new_[18747]_  | ~\new_[17003]_ );
  assign \new_[8705]_  = ~\new_[9464]_  & (~\new_[18499]_  | ~\new_[16804]_ );
  assign \new_[8706]_  = ~\new_[9465]_  & (~\new_[19626]_  | ~\new_[16790]_ );
  assign \new_[8707]_  = ~\new_[9466]_  & (~\new_[18701]_  | ~\new_[16896]_ );
  assign \new_[8708]_  = ~\new_[9467]_  & (~\new_[19172]_  | ~\new_[17001]_ );
  assign \new_[8709]_  = ~\new_[9468]_  & (~\new_[17813]_  | ~\new_[16679]_ );
  assign \new_[8710]_  = ~\new_[9469]_  & (~\new_[17969]_  | ~\new_[16805]_ );
  assign \new_[8711]_  = ~\new_[9470]_  & (~\new_[18956]_  | ~\new_[17131]_ );
  assign \new_[8712]_  = ~\new_[9471]_  & (~\new_[18339]_  | ~\new_[16796]_ );
  assign \new_[8713]_  = ~\new_[9472]_  & (~\new_[19152]_  | ~\new_[16797]_ );
  assign \new_[8714]_  = \new_[9541]_  ? \new_[17131]_  : \new_[18891]_ ;
  assign \new_[8715]_  = \new_[9545]_  ? \new_[16797]_  : \new_[18029]_ ;
  assign \new_[8716]_  = \new_[9548]_  ? \new_[16805]_  : \new_[18771]_ ;
  assign \new_[8717]_  = \new_[9558]_  ? \new_[16797]_  : \new_[19794]_ ;
  assign \new_[8718]_  = \new_[9551]_  ? \new_[17131]_  : \new_[18341]_ ;
  assign \new_[8719]_  = \new_[9536]_  ? \new_[17003]_  : \new_[17925]_ ;
  assign \new_[8720]_  = \new_[9537]_  ? \new_[17003]_  : \new_[19369]_ ;
  assign \new_[8721]_  = \new_[9538]_  ? \new_[17003]_  : \new_[19664]_ ;
  assign \new_[8722]_  = \new_[9539]_  ? \new_[17003]_  : \new_[19825]_ ;
  assign \new_[8723]_  = \new_[9540]_  ? \new_[17003]_  : \new_[18876]_ ;
  assign \new_[8724]_  = \new_[9541]_  ? \new_[17003]_  : \new_[18654]_ ;
  assign \new_[8725]_  = \new_[9542]_  ? \new_[17003]_  : \new_[18930]_ ;
  assign \new_[8726]_  = \new_[9543]_  ? \new_[17003]_  : \new_[18573]_ ;
  assign \new_[8727]_  = \new_[9544]_  ? \new_[17003]_  : \new_[18720]_ ;
  assign \new_[8728]_  = \new_[9545]_  ? \new_[17003]_  : \new_[18443]_ ;
  assign \new_[8729]_  = \new_[9546]_  ? \new_[17003]_  : \new_[18633]_ ;
  assign \new_[8730]_  = \new_[8388]_ ;
  assign \new_[8731]_  = \new_[9547]_  ? \new_[17003]_  : \new_[18366]_ ;
  assign \new_[8732]_  = \new_[9548]_  ? \new_[17003]_  : \new_[18537]_ ;
  assign \new_[8733]_  = \new_[9549]_  ? \new_[17003]_  : \new_[19107]_ ;
  assign \new_[8734]_  = \new_[9550]_  ? \new_[17003]_  : \new_[19113]_ ;
  assign \new_[8735]_  = \new_[9551]_  ? \new_[17003]_  : \new_[19858]_ ;
  assign \new_[8736]_  = \new_[9552]_  ? \new_[17003]_  : \new_[18668]_ ;
  assign \new_[8737]_  = \new_[9553]_  ? \new_[17003]_  : \new_[18292]_ ;
  assign \new_[8738]_  = \new_[9554]_  ? \new_[17003]_  : \new_[17952]_ ;
  assign \new_[8739]_  = \new_[9555]_  ? \new_[17003]_  : \new_[18973]_ ;
  assign \new_[8740]_  = \new_[9556]_  ? \new_[17003]_  : \new_[19089]_ ;
  assign \new_[8741]_  = \new_[9557]_  ? \new_[17003]_  : \new_[18777]_ ;
  assign \new_[8742]_  = \new_[9558]_  ? \new_[17003]_  : \new_[18529]_ ;
  assign \new_[8743]_  = \new_[9559]_  ? \new_[17003]_  : \new_[18820]_ ;
  assign \new_[8744]_  = \new_[9536]_  ? \new_[16804]_  : \new_[19537]_ ;
  assign \new_[8745]_  = \new_[9537]_  ? \new_[16804]_  : \new_[18752]_ ;
  assign \new_[8746]_  = \new_[9538]_  ? \new_[16804]_  : \new_[19118]_ ;
  assign \new_[8747]_  = \new_[9539]_  ? \new_[16804]_  : \new_[18627]_ ;
  assign \new_[8748]_  = \new_[9540]_  ? \new_[16804]_  : \new_[18324]_ ;
  assign \new_[8749]_  = \new_[9541]_  ? \new_[16804]_  : \new_[18342]_ ;
  assign \new_[8750]_  = \new_[9542]_  ? \new_[16804]_  : \new_[19036]_ ;
  assign \new_[8751]_  = \new_[9543]_  ? \new_[16804]_  : \new_[19251]_ ;
  assign \new_[8752]_  = \new_[9544]_  ? \new_[16804]_  : \new_[18135]_ ;
  assign \new_[8753]_  = \new_[9545]_  ? \new_[16804]_  : \new_[18557]_ ;
  assign \new_[8754]_  = \new_[9546]_  ? \new_[16804]_  : \new_[19372]_ ;
  assign \new_[8755]_  = \new_[9547]_  ? \new_[16804]_  : \new_[18723]_ ;
  assign \new_[8756]_  = \new_[9548]_  ? \new_[16804]_  : \new_[18351]_ ;
  assign \new_[8757]_  = \new_[9549]_  ? \new_[16804]_  : \new_[19854]_ ;
  assign \new_[8758]_  = \new_[9550]_  ? \new_[16804]_  : \new_[18707]_ ;
  assign \new_[8759]_  = \new_[9551]_  ? \new_[16804]_  : \new_[18846]_ ;
  assign \new_[8760]_  = \new_[9552]_  ? \new_[16804]_  : \new_[17895]_ ;
  assign \new_[8761]_  = \new_[9553]_  ? \new_[16804]_  : \new_[18869]_ ;
  assign \new_[8762]_  = \new_[9554]_  ? \new_[16804]_  : \new_[19796]_ ;
  assign \new_[8763]_  = \new_[9555]_  ? \new_[16804]_  : \new_[19797]_ ;
  assign \new_[8764]_  = \new_[9556]_  ? \new_[16804]_  : \new_[17823]_ ;
  assign \new_[8765]_  = \new_[9558]_  ? \new_[16804]_  : \new_[18945]_ ;
  assign \new_[8766]_  = \new_[9559]_  ? \new_[16804]_  : \new_[18826]_ ;
  assign \new_[8767]_  = \new_[9536]_  ? \new_[17001]_  : \new_[19625]_ ;
  assign \new_[8768]_  = \new_[9537]_  ? \new_[17001]_  : \new_[18993]_ ;
  assign \new_[8769]_  = \new_[9538]_  ? \new_[17001]_  : \new_[19561]_ ;
  assign \new_[8770]_  = \new_[9539]_  ? \new_[17001]_  : \new_[19157]_ ;
  assign \new_[8771]_  = \new_[9540]_  ? \new_[17001]_  : \new_[17850]_ ;
  assign \new_[8772]_  = \new_[9541]_  ? \new_[17001]_  : \new_[18191]_ ;
  assign \new_[8773]_  = \new_[9543]_  ? \new_[17001]_  : \new_[18631]_ ;
  assign \new_[8774]_  = \new_[9542]_  ? \new_[17001]_  : \new_[19263]_ ;
  assign \new_[8775]_  = \new_[9544]_  ? \new_[17001]_  : \new_[19144]_ ;
  assign \new_[8776]_  = \new_[9545]_  ? \new_[17001]_  : \new_[19260]_ ;
  assign \new_[8777]_  = \new_[9546]_  ? \new_[17001]_  : \new_[18315]_ ;
  assign \new_[8778]_  = \new_[9547]_  ? \new_[17001]_  : \new_[17942]_ ;
  assign \new_[8779]_  = \new_[9548]_  ? \new_[17001]_  : \new_[18018]_ ;
  assign \new_[8780]_  = \new_[9549]_  ? \new_[17001]_  : \new_[19055]_ ;
  assign \new_[8781]_  = \new_[9550]_  ? \new_[17001]_  : \new_[18641]_ ;
  assign \new_[8782]_  = \new_[9552]_  ? \new_[17001]_  : \new_[18899]_ ;
  assign \new_[8783]_  = \new_[9553]_  ? \new_[17001]_  : \new_[18225]_ ;
  assign \new_[8784]_  = \new_[9554]_  ? \new_[17001]_  : \new_[18845]_ ;
  assign \new_[8785]_  = \new_[9555]_  ? \new_[17001]_  : \new_[19265]_ ;
  assign \new_[8786]_  = \new_[9556]_  ? \new_[17001]_  : \new_[18287]_ ;
  assign \new_[8787]_  = \new_[9557]_  ? \new_[17001]_  : \new_[18299]_ ;
  assign \new_[8788]_  = \new_[9559]_  ? \new_[17001]_  : \new_[18501]_ ;
  assign \new_[8789]_  = \new_[9557]_  ? \new_[16804]_  : \new_[18528]_ ;
  assign \new_[8790]_  = \new_[9536]_  ? \new_[16805]_  : \new_[18526]_ ;
  assign \new_[8791]_  = \new_[9537]_  ? \new_[16805]_  : \new_[19855]_ ;
  assign \new_[8792]_  = \new_[9538]_  ? \new_[16805]_  : \new_[18844]_ ;
  assign \new_[8793]_  = \new_[9539]_  ? \new_[16805]_  : \new_[18483]_ ;
  assign \new_[8794]_  = \new_[9540]_  ? \new_[16805]_  : \new_[19657]_ ;
  assign \new_[8795]_  = \new_[9541]_  ? \new_[16805]_  : \new_[19648]_ ;
  assign \new_[8796]_  = \new_[9542]_  ? \new_[16805]_  : \new_[17886]_ ;
  assign \new_[8797]_  = \new_[9543]_  ? \new_[16805]_  : \new_[19156]_ ;
  assign \new_[8798]_  = \new_[9544]_  ? \new_[16805]_  : \new_[19388]_ ;
  assign \new_[8799]_  = \new_[9545]_  ? \new_[16805]_  : \new_[18140]_ ;
  assign \new_[8800]_  = \new_[9546]_  ? \new_[16805]_  : \new_[19444]_ ;
  assign \new_[8801]_  = \new_[9547]_  ? \new_[16805]_  : \new_[19279]_ ;
  assign \new_[8802]_  = \new_[9549]_  ? \new_[16805]_  : \new_[18856]_ ;
  assign \new_[8803]_  = \new_[9550]_  ? \new_[16805]_  : \new_[18730]_ ;
  assign \new_[8804]_  = \new_[9551]_  ? \new_[16805]_  : \new_[19364]_ ;
  assign \new_[8805]_  = \new_[9552]_  ? \new_[16805]_  : \new_[18972]_ ;
  assign \new_[8806]_  = \new_[9553]_  ? \new_[16805]_  : \new_[19320]_ ;
  assign \new_[8807]_  = \new_[9554]_  ? \new_[16805]_  : \new_[19754]_ ;
  assign \new_[8808]_  = \new_[9555]_  ? \new_[16805]_  : \new_[19019]_ ;
  assign \new_[8809]_  = \new_[9556]_  ? \new_[16805]_  : \new_[18695]_ ;
  assign \new_[8810]_  = \new_[9557]_  ? \new_[16805]_  : \new_[18889]_ ;
  assign \new_[8811]_  = \new_[9558]_  ? \new_[16805]_  : \new_[19165]_ ;
  assign \new_[8812]_  = \new_[9559]_  ? \new_[16805]_  : \new_[18749]_ ;
  assign \new_[8813]_  = \new_[9536]_  ? \new_[17131]_  : \new_[19061]_ ;
  assign \new_[8814]_  = \new_[9537]_  ? \new_[17131]_  : \new_[18811]_ ;
  assign \new_[8815]_  = \new_[9538]_  ? \new_[17131]_  : \new_[18857]_ ;
  assign \new_[8816]_  = \new_[9539]_  ? \new_[17131]_  : \new_[19179]_ ;
  assign \new_[8817]_  = \new_[9540]_  ? \new_[17131]_  : \new_[19053]_ ;
  assign \new_[8818]_  = \new_[9542]_  ? \new_[17131]_  : \new_[18682]_ ;
  assign \new_[8819]_  = \new_[9543]_  ? \new_[17131]_  : \new_[20002]_ ;
  assign \new_[8820]_  = \new_[9544]_  ? \new_[17131]_  : \new_[19611]_ ;
  assign \new_[8821]_  = \new_[9545]_  ? \new_[17131]_  : \new_[18736]_ ;
  assign \new_[8822]_  = \new_[9546]_  ? \new_[17131]_  : \new_[18794]_ ;
  assign \new_[8823]_  = \new_[9547]_  ? \new_[17131]_  : \new_[19602]_ ;
  assign \new_[8824]_  = \new_[9549]_  ? \new_[17131]_  : \new_[18385]_ ;
  assign \new_[8825]_  = \new_[9550]_  ? \new_[17131]_  : \new_[19200]_ ;
  assign \new_[8826]_  = \new_[9552]_  ? \new_[17131]_  : \new_[18230]_ ;
  assign \new_[8827]_  = \new_[9553]_  ? \new_[17131]_  : \new_[18776]_ ;
  assign \new_[8828]_  = \new_[9554]_  ? \new_[17131]_  : \new_[18675]_ ;
  assign \new_[8829]_  = \new_[9555]_  ? \new_[17131]_  : \new_[19007]_ ;
  assign \new_[8830]_  = \new_[9556]_  ? \new_[17131]_  : \new_[18148]_ ;
  assign \new_[8831]_  = \new_[9557]_  ? \new_[17131]_  : \new_[17962]_ ;
  assign \new_[8832]_  = \new_[9558]_  ? \new_[17131]_  : \new_[17910]_ ;
  assign \new_[8833]_  = \new_[9559]_  ? \new_[17131]_  : \new_[19549]_ ;
  assign \new_[8834]_  = \new_[9548]_  ? \new_[17131]_  : \new_[19066]_ ;
  assign \new_[8835]_  = \new_[9536]_  ? \new_[16797]_  : \new_[18705]_ ;
  assign \new_[8836]_  = \new_[9537]_  ? \new_[16797]_  : \new_[17980]_ ;
  assign \new_[8837]_  = \new_[9538]_  ? \new_[16797]_  : \new_[18960]_ ;
  assign \new_[8838]_  = \new_[9539]_  ? \new_[16797]_  : \new_[19361]_ ;
  assign \new_[8839]_  = \new_[9540]_  ? \new_[16797]_  : \new_[18359]_ ;
  assign \new_[8840]_  = \new_[9541]_  ? \new_[16797]_  : \new_[17806]_ ;
  assign \new_[8841]_  = \new_[9542]_  ? \new_[16797]_  : \new_[19230]_ ;
  assign \new_[8842]_  = \new_[9543]_  ? \new_[16797]_  : \new_[19203]_ ;
  assign \new_[8843]_  = \new_[9544]_  ? \new_[16797]_  : \new_[18195]_ ;
  assign \new_[8844]_  = \new_[9546]_  ? \new_[16797]_  : \new_[17877]_ ;
  assign \new_[8845]_  = \new_[9547]_  ? \new_[16797]_  : \new_[19767]_ ;
  assign \new_[8846]_  = \new_[9548]_  ? \new_[16797]_  : \new_[18614]_ ;
  assign \new_[8847]_  = \new_[9549]_  ? \new_[16797]_  : \new_[18532]_ ;
  assign \new_[8848]_  = \new_[9550]_  ? \new_[16797]_  : \new_[18667]_ ;
  assign \new_[8849]_  = \new_[9551]_  ? \new_[16797]_  : \new_[18986]_ ;
  assign \new_[8850]_  = \new_[9552]_  ? \new_[16797]_  : \new_[19787]_ ;
  assign \new_[8851]_  = \new_[9553]_  ? \new_[16797]_  : \new_[19714]_ ;
  assign \new_[8852]_  = \new_[9554]_  ? \new_[16797]_  : \new_[19800]_ ;
  assign \new_[8853]_  = \new_[9555]_  ? \new_[16797]_  : \new_[19834]_ ;
  assign \new_[8854]_  = \new_[9556]_  ? \new_[16797]_  : \new_[18637]_ ;
  assign \new_[8855]_  = \new_[9557]_  ? \new_[16797]_  : \new_[18691]_ ;
  assign \new_[8856]_  = \new_[9559]_  ? \new_[16797]_  : \new_[17945]_ ;
  assign \new_[8857]_  = \new_[9558]_  ? \new_[17001]_  : \new_[19188]_ ;
  assign \new_[8858]_  = \new_[9551]_  ? \new_[17001]_  : \new_[18394]_ ;
  assign \new_[8859]_  = \new_[9558]_  ? \new_[16790]_  : \new_[19344]_ ;
  assign \new_[8860]_  = \new_[9541]_  ? \new_[16679]_  : \new_[18952]_ ;
  assign \new_[8861]_  = \new_[9541]_  ? \new_[16896]_  : \new_[18388]_ ;
  assign \new_[8862]_  = \new_[9554]_  ? \new_[16796]_  : \new_[19612]_ ;
  assign \new_[8863]_  = \new_[9536]_  ? \new_[16662]_  : \new_[19853]_ ;
  assign \new_[8864]_  = \new_[9537]_  ? \new_[16662]_  : \new_[19425]_ ;
  assign \new_[8865]_  = \new_[9538]_  ? \new_[16662]_  : \new_[18354]_ ;
  assign \new_[8866]_  = \new_[9539]_  ? \new_[16662]_  : \new_[19332]_ ;
  assign \new_[8867]_  = \new_[9540]_  ? \new_[16662]_  : \new_[17976]_ ;
  assign \new_[8868]_  = \new_[9541]_  ? \new_[16662]_  : \new_[17977]_ ;
  assign \new_[8869]_  = \new_[9542]_  ? \new_[16662]_  : \new_[19832]_ ;
  assign \new_[8870]_  = \new_[9543]_  ? \new_[16662]_  : \new_[18117]_ ;
  assign \new_[8871]_  = \new_[9544]_  ? \new_[16662]_  : \new_[18030]_ ;
  assign \new_[8872]_  = \new_[9545]_  ? \new_[16662]_  : \new_[18569]_ ;
  assign \new_[8873]_  = \new_[9546]_  ? \new_[16662]_  : \new_[17897]_ ;
  assign \new_[8874]_  = \new_[9547]_  ? \new_[16662]_  : \new_[19109]_ ;
  assign \new_[8875]_  = \new_[9548]_  ? \new_[16662]_  : \new_[18963]_ ;
  assign \new_[8876]_  = \new_[9549]_  ? \new_[16662]_  : \new_[19547]_ ;
  assign \new_[8877]_  = \new_[9550]_  ? \new_[16662]_  : \new_[19645]_ ;
  assign \new_[8878]_  = \new_[9551]_  ? \new_[16662]_  : \new_[19236]_ ;
  assign \new_[8879]_  = \new_[9552]_  ? \new_[16662]_  : \new_[18238]_ ;
  assign \new_[8880]_  = \new_[9553]_  ? \new_[16662]_  : \new_[17864]_ ;
  assign \new_[8881]_  = \new_[9554]_  ? \new_[16662]_  : \new_[19276]_ ;
  assign \new_[8882]_  = \new_[9555]_  ? \new_[16662]_  : \new_[19353]_ ;
  assign \new_[8883]_  = \new_[9556]_  ? \new_[16662]_  : \new_[18101]_ ;
  assign \new_[8884]_  = \new_[9557]_  ? \new_[16662]_  : \new_[18670]_ ;
  assign \new_[8885]_  = \new_[9558]_  ? \new_[16662]_  : \new_[18969]_ ;
  assign \new_[8886]_  = \new_[9559]_  ? \new_[16662]_  : \new_[18311]_ ;
  assign \new_[8887]_  = \new_[9536]_  ? \new_[16790]_  : \new_[18192]_ ;
  assign \new_[8888]_  = \new_[9537]_  ? \new_[16790]_  : \new_[19305]_ ;
  assign \new_[8889]_  = \new_[9538]_  ? \new_[16790]_  : \new_[19592]_ ;
  assign \new_[8890]_  = \new_[9539]_  ? \new_[16790]_  : \new_[18216]_ ;
  assign \new_[8891]_  = \new_[9540]_  ? \new_[16790]_  : \new_[19405]_ ;
  assign \new_[8892]_  = \new_[9541]_  ? \new_[16790]_  : \new_[18071]_ ;
  assign \new_[8893]_  = \new_[9542]_  ? \new_[16790]_  : \new_[19014]_ ;
  assign \new_[8894]_  = \new_[9543]_  ? \new_[16790]_  : \new_[19700]_ ;
  assign \new_[8895]_  = \new_[9544]_  ? \new_[16790]_  : \new_[18214]_ ;
  assign \new_[8896]_  = \new_[9545]_  ? \new_[16790]_  : \new_[19753]_ ;
  assign \new_[8897]_  = \new_[9546]_  ? \new_[16790]_  : \new_[18692]_ ;
  assign \new_[8898]_  = \new_[9547]_  ? \new_[16790]_  : \new_[19624]_ ;
  assign \new_[8899]_  = \new_[9548]_  ? \new_[16790]_  : \new_[19247]_ ;
  assign \new_[8900]_  = \new_[9549]_  ? \new_[16790]_  : \new_[19149]_ ;
  assign \new_[8901]_  = \new_[9550]_  ? \new_[16790]_  : \new_[18906]_ ;
  assign \new_[8902]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[6] ;
  assign \new_[8903]_  = \new_[9551]_  ? \new_[16790]_  : \new_[19824]_ ;
  assign \new_[8904]_  = \new_[9552]_  ? \new_[16790]_  : \new_[19394]_ ;
  assign \new_[8905]_  = \new_[9553]_  ? \new_[16790]_  : \new_[19047]_ ;
  assign \new_[8906]_  = \new_[9554]_  ? \new_[16790]_  : \new_[19718]_ ;
  assign \new_[8907]_  = \new_[9555]_  ? \new_[16790]_  : \new_[19668]_ ;
  assign \new_[8908]_  = \new_[9556]_  ? \new_[16790]_  : \new_[18416]_ ;
  assign \new_[8909]_  = \new_[9557]_  ? \new_[16790]_  : \new_[18694]_ ;
  assign \new_[8910]_  = \new_[9559]_  ? \new_[16790]_  : \new_[19395]_ ;
  assign \new_[8911]_  = \new_[9536]_  ? \new_[16896]_  : \new_[18718]_ ;
  assign \new_[8912]_  = \new_[9537]_  ? \new_[16896]_  : \new_[19707]_ ;
  assign \new_[8913]_  = \new_[9538]_  ? \new_[16896]_  : \new_[18052]_ ;
  assign \new_[8914]_  = \new_[9539]_  ? \new_[16896]_  : \new_[19368]_ ;
  assign \new_[8915]_  = \new_[9540]_  ? \new_[16896]_  : \new_[19428]_ ;
  assign \new_[8916]_  = \new_[9542]_  ? \new_[16896]_  : \new_[19383]_ ;
  assign \new_[8917]_  = \new_[9543]_  ? \new_[16896]_  : \new_[19358]_ ;
  assign \new_[8918]_  = \new_[9544]_  ? \new_[16896]_  : \new_[17930]_ ;
  assign \new_[8919]_  = \new_[9545]_  ? \new_[16896]_  : \new_[18401]_ ;
  assign \new_[8920]_  = \new_[9546]_  ? \new_[16896]_  : \new_[18399]_ ;
  assign \new_[8921]_  = \new_[9547]_  ? \new_[16896]_  : \new_[17929]_ ;
  assign \new_[8922]_  = \new_[9549]_  ? \new_[16896]_  : \new_[19414]_ ;
  assign \new_[8923]_  = \new_[9550]_  ? \new_[16896]_  : \new_[17926]_ ;
  assign \new_[8924]_  = \new_[9551]_  ? \new_[16896]_  : \new_[18455]_ ;
  assign \new_[8925]_  = \new_[9552]_  ? \new_[16896]_  : \new_[19373]_ ;
  assign \new_[8926]_  = \new_[9553]_  ? \new_[16896]_  : \new_[19198]_ ;
  assign \new_[8927]_  = \new_[9554]_  ? \new_[16896]_  : \new_[19408]_ ;
  assign \new_[8928]_  = \new_[9555]_  ? \new_[16896]_  : \new_[17922]_ ;
  assign \new_[8929]_  = \new_[9556]_  ? \new_[16896]_  : \new_[18453]_ ;
  assign \new_[8930]_  = \new_[9557]_  ? \new_[16896]_  : \new_[17916]_ ;
  assign \new_[8931]_  = \new_[9558]_  ? \new_[16896]_  : \new_[17915]_ ;
  assign \new_[8932]_  = \new_[9559]_  ? \new_[16896]_  : \new_[19396]_ ;
  assign \new_[8933]_  = \new_[9536]_  ? \new_[16679]_  : \new_[17913]_ ;
  assign \new_[8934]_  = \new_[9537]_  ? \new_[16679]_  : \new_[17911]_ ;
  assign \new_[8935]_  = \new_[9538]_  ? \new_[16679]_  : \new_[19106]_ ;
  assign \new_[8936]_  = \new_[9539]_  ? \new_[16679]_  : \new_[18604]_ ;
  assign \new_[8937]_  = \new_[9540]_  ? \new_[16679]_  : \new_[19249]_ ;
  assign \new_[8938]_  = \new_[9542]_  ? \new_[16679]_  : \new_[18181]_ ;
  assign \new_[8939]_  = \new_[9543]_  ? \new_[16679]_  : \new_[20016]_ ;
  assign \new_[8940]_  = \new_[9544]_  ? \new_[16679]_  : \new_[18513]_ ;
  assign \new_[8941]_  = \new_[9545]_  ? \new_[16679]_  : \new_[19253]_ ;
  assign \new_[8942]_  = \new_[9546]_  ? \new_[16679]_  : \new_[19338]_ ;
  assign \new_[8943]_  = \new_[9547]_  ? \new_[16679]_  : \new_[19335]_ ;
  assign \new_[8944]_  = \new_[9548]_  ? \new_[16679]_  : \new_[18019]_ ;
  assign \new_[8945]_  = \new_[9549]_  ? \new_[16679]_  : \new_[17992]_ ;
  assign \new_[8946]_  = \new_[9550]_  ? \new_[16679]_  : \new_[17949]_ ;
  assign \new_[8947]_  = \new_[9551]_  ? \new_[16679]_  : \new_[17939]_ ;
  assign \new_[8948]_  = \new_[9552]_  ? \new_[16679]_  : \new_[19514]_ ;
  assign \new_[8949]_  = \new_[9553]_  ? \new_[16679]_  : \new_[17888]_ ;
  assign \new_[8950]_  = \new_[9554]_  ? \new_[16679]_  : \new_[19268]_ ;
  assign \new_[8951]_  = \new_[9555]_  ? \new_[16679]_  : \new_[18783]_ ;
  assign \new_[8952]_  = \new_[9556]_  ? \new_[16679]_  : \new_[17956]_ ;
  assign \new_[8953]_  = \new_[9557]_  ? \new_[16679]_  : \new_[18796]_ ;
  assign \new_[8954]_  = \new_[9558]_  ? \new_[16679]_  : \new_[18472]_ ;
  assign \new_[8955]_  = \new_[9559]_  ? \new_[16679]_  : \new_[19406]_ ;
  assign \new_[8956]_  = \new_[9538]_  ? \new_[16796]_  : \new_[19223]_ ;
  assign \new_[8957]_  = \new_[9536]_  ? \new_[16796]_  : \new_[18781]_ ;
  assign \new_[8958]_  = \new_[9539]_  ? \new_[16796]_  : \new_[19665]_ ;
  assign \new_[8959]_  = \new_[9540]_  ? \new_[16796]_  : \new_[19545]_ ;
  assign \new_[8960]_  = \new_[9541]_  ? \new_[16796]_  : \new_[19658]_ ;
  assign \new_[8961]_  = \new_[9542]_  ? \new_[16796]_  : \new_[18959]_ ;
  assign \new_[8962]_  = \new_[9537]_  ? \new_[16796]_  : \new_[18164]_ ;
  assign \new_[8963]_  = \new_[9543]_  ? \new_[16796]_  : \new_[18516]_ ;
  assign \new_[8964]_  = \new_[9544]_  ? \new_[16796]_  : \new_[18571]_ ;
  assign \new_[8965]_  = \new_[9545]_  ? \new_[16796]_  : \new_[18790]_ ;
  assign \new_[8966]_  = \new_[9546]_  ? \new_[16796]_  : \new_[19006]_ ;
  assign \new_[8967]_  = \new_[9547]_  ? \new_[16796]_  : \new_[18469]_ ;
  assign \new_[8968]_  = \new_[9548]_  ? \new_[16796]_  : \new_[19788]_ ;
  assign \new_[8969]_  = \new_[9549]_  ? \new_[16796]_  : \new_[19722]_ ;
  assign \new_[8970]_  = \new_[9550]_  ? \new_[16796]_  : \new_[19022]_ ;
  assign \new_[8971]_  = \new_[9551]_  ? \new_[16796]_  : \new_[19727]_ ;
  assign \new_[8972]_  = \new_[9552]_  ? \new_[16796]_  : \new_[18563]_ ;
  assign \new_[8973]_  = \new_[9553]_  ? \new_[16796]_  : \new_[19092]_ ;
  assign \new_[8974]_  = \new_[9555]_  ? \new_[16796]_  : \new_[18231]_ ;
  assign \new_[8975]_  = \new_[9556]_  ? \new_[16796]_  : \new_[18559]_ ;
  assign \new_[8976]_  = \new_[9557]_  ? \new_[16796]_  : \new_[19391]_ ;
  assign \new_[8977]_  = \new_[9558]_  ? \new_[16796]_  : \new_[19370]_ ;
  assign \new_[8978]_  = \new_[9559]_  ? \new_[16796]_  : \new_[19059]_ ;
  assign \new_[8979]_  = \new_[9548]_  ? \new_[16896]_  : \new_[17927]_ ;
  assign \new_[8980]_  = \new_[19097]_  ? \new_[17191]_  : \new_[9557]_ ;
  assign \new_[8981]_  = \new_[18536]_  ? \new_[16911]_  : \new_[9554]_ ;
  assign \new_[8982]_  = \new_[19757]_  ? \new_[17191]_  : \new_[9550]_ ;
  assign \new_[8983]_  = \new_[17983]_  ? \new_[16975]_  : \new_[9536]_ ;
  assign \new_[8984]_  = \new_[19103]_  ? \new_[16975]_  : \new_[9537]_ ;
  assign \new_[8985]_  = \new_[19079]_  ? \new_[16975]_  : \new_[9538]_ ;
  assign \new_[8986]_  = \new_[18257]_  ? \new_[16975]_  : \new_[9539]_ ;
  assign \new_[8987]_  = \new_[18655]_  ? \new_[16975]_  : \new_[9540]_ ;
  assign \new_[8988]_  = \new_[18818]_  ? \new_[16975]_  : \new_[9541]_ ;
  assign \new_[8989]_  = \new_[19659]_  ? \new_[16975]_  : \new_[9542]_ ;
  assign \new_[8990]_  = \new_[18504]_  ? \new_[16975]_  : \new_[9543]_ ;
  assign \new_[8991]_  = \new_[17879]_  ? \new_[16975]_  : \new_[9544]_ ;
  assign \new_[8992]_  = \new_[18444]_  ? \new_[16975]_  : \new_[9545]_ ;
  assign \new_[8993]_  = \new_[19495]_  ? \new_[16975]_  : \new_[9546]_ ;
  assign \new_[8994]_  = \new_[19206]_  ? \new_[16975]_  : \new_[9547]_ ;
  assign \new_[8995]_  = \new_[18106]_  ? \new_[16975]_  : \new_[9548]_ ;
  assign \new_[8996]_  = \new_[18997]_  ? \new_[16975]_  : \new_[9549]_ ;
  assign \new_[8997]_  = \new_[19581]_  ? \new_[16975]_  : \new_[9550]_ ;
  assign \new_[8998]_  = \new_[18285]_  ? \new_[16975]_  : \new_[9551]_ ;
  assign \new_[8999]_  = \new_[18121]_  ? \new_[16975]_  : \new_[9552]_ ;
  assign \new_[9000]_  = \new_[19352]_  ? \new_[16975]_  : \new_[9553]_ ;
  assign \new_[9001]_  = \new_[18578]_  ? \new_[16975]_  : \new_[9554]_ ;
  assign \new_[9002]_  = \new_[17904]_  ? \new_[16975]_  : \new_[9555]_ ;
  assign \new_[9003]_  = \new_[18947]_  ? \new_[16975]_  : \new_[9531]_ ;
  assign \new_[9004]_  = \new_[18636]_  ? \new_[16975]_  : \new_[9556]_ ;
  assign \new_[9005]_  = \new_[18329]_  ? \new_[16975]_  : \new_[9557]_ ;
  assign \new_[9006]_  = \new_[19607]_  ? \new_[16975]_  : \new_[9558]_ ;
  assign \new_[9007]_  = \new_[18931]_  ? \new_[16975]_  : \new_[9559]_ ;
  assign \new_[9008]_  = \new_[18484]_  ? \new_[16976]_  : \new_[9536]_ ;
  assign \new_[9009]_  = \new_[18242]_  ? \new_[16976]_  : \new_[9537]_ ;
  assign \new_[9010]_  = \new_[19446]_  ? \new_[16976]_  : \new_[9538]_ ;
  assign \new_[9011]_  = \new_[19421]_  ? \new_[16976]_  : \new_[9539]_ ;
  assign \new_[9012]_  = \new_[18905]_  ? \new_[16976]_  : \new_[9541]_ ;
  assign \new_[9013]_  = \new_[18064]_  ? \new_[16976]_  : \new_[9542]_ ;
  assign \new_[9014]_  = \new_[18981]_  ? \new_[16976]_  : \new_[9543]_ ;
  assign \new_[9015]_  = \new_[19697]_  ? \new_[16976]_  : \new_[9544]_ ;
  assign \new_[9016]_  = \new_[19566]_  ? \new_[16976]_  : \new_[9545]_ ;
  assign \new_[9017]_  = \new_[19087]_  ? \new_[16976]_  : \new_[9546]_ ;
  assign \new_[9018]_  = \new_[18878]_  ? \new_[16976]_  : \new_[9547]_ ;
  assign \new_[9019]_  = \new_[17973]_  ? \new_[16976]_  : \new_[9548]_ ;
  assign \new_[9020]_  = \new_[19988]_  ? \new_[16976]_  : \new_[9549]_ ;
  assign \new_[9021]_  = \new_[18621]_  ? \new_[16976]_  : \new_[9550]_ ;
  assign \new_[9022]_  = \new_[19057]_  ? \new_[16976]_  : \new_[9551]_ ;
  assign \new_[9023]_  = \new_[18326]_  ? \new_[16976]_  : \new_[9552]_ ;
  assign \new_[9024]_  = \new_[19693]_  ? \new_[16976]_  : \new_[9553]_ ;
  assign \new_[9025]_  = \new_[19073]_  ? \new_[16976]_  : \new_[9554]_ ;
  assign \new_[9026]_  = \new_[19680]_  ? \new_[16976]_  : \new_[9555]_ ;
  assign \new_[9027]_  = \new_[19267]_  ? \new_[16976]_  : \new_[9531]_ ;
  assign \new_[9028]_  = \new_[18863]_  ? \new_[16976]_  : \new_[9556]_ ;
  assign \new_[9029]_  = \new_[19243]_  ? \new_[16976]_  : \new_[9557]_ ;
  assign \new_[9030]_  = \new_[18898]_  ? \new_[16976]_  : \new_[9558]_ ;
  assign \new_[9031]_  = \new_[18881]_  ? \new_[16976]_  : \new_[9559]_ ;
  assign \new_[9032]_  = \new_[18070]_  ? \new_[16900]_  : \new_[9536]_ ;
  assign \new_[9033]_  = \new_[18979]_  ? \new_[16900]_  : \new_[9537]_ ;
  assign \new_[9034]_  = \new_[19035]_  ? \new_[16900]_  : \new_[9538]_ ;
  assign \new_[9035]_  = \new_[19085]_  ? \new_[16900]_  : \new_[9539]_ ;
  assign \new_[9036]_  = \new_[19300]_  ? \new_[16900]_  : \new_[9540]_ ;
  assign \new_[9037]_  = \new_[19460]_  ? \new_[16900]_  : \new_[9541]_ ;
  assign \new_[9038]_  = \new_[17901]_  ? \new_[16900]_  : \new_[9542]_ ;
  assign \new_[9039]_  = \new_[18687]_  ? \new_[16900]_  : \new_[9543]_ ;
  assign \new_[9040]_  = \new_[18601]_  ? \new_[16900]_  : \new_[9545]_ ;
  assign \new_[9041]_  = \new_[18983]_  ? \new_[16900]_  : \new_[9546]_ ;
  assign \new_[9042]_  = \new_[18975]_  ? \new_[16900]_  : \new_[9547]_ ;
  assign \new_[9043]_  = \new_[18567]_  ? \new_[16900]_  : \new_[9548]_ ;
  assign \new_[9044]_  = \new_[18630]_  ? \new_[16900]_  : \new_[9549]_ ;
  assign \new_[9045]_  = \new_[18381]_  ? \new_[16900]_  : \new_[9550]_ ;
  assign \new_[9046]_  = \new_[19635]_  ? \new_[16900]_  : \new_[9551]_ ;
  assign \new_[9047]_  = \new_[19101]_  ? \new_[16900]_  : \new_[9552]_ ;
  assign \new_[9048]_  = \new_[18530]_  ? \new_[16900]_  : \new_[9553]_ ;
  assign \new_[9049]_  = \new_[19176]_  ? \new_[16900]_  : \new_[9554]_ ;
  assign \new_[9050]_  = \new_[18218]_  ? \new_[16900]_  : \new_[9555]_ ;
  assign \new_[9051]_  = \new_[18544]_  ? \new_[16900]_  : \new_[9531]_ ;
  assign \new_[9052]_  = \new_[18186]_  ? \new_[16900]_  : \new_[9556]_ ;
  assign \new_[9053]_  = \new_[18112]_  ? \new_[16900]_  : \new_[9557]_ ;
  assign \new_[9054]_  = \new_[19441]_  ? \new_[16900]_  : \new_[9558]_ ;
  assign \new_[9055]_  = \new_[19443]_  ? \new_[16900]_  : \new_[9559]_ ;
  assign \new_[9056]_  = \new_[18034]_  ? \new_[17191]_  : \new_[9536]_ ;
  assign \new_[9057]_  = \new_[19450]_  ? \new_[17191]_  : \new_[9537]_ ;
  assign \new_[9058]_  = \new_[18004]_  ? \new_[17191]_  : \new_[9538]_ ;
  assign \new_[9059]_  = \new_[17990]_  ? \new_[17191]_  : \new_[9539]_ ;
  assign \new_[9060]_  = \new_[19490]_  ? \new_[17191]_  : \new_[9540]_ ;
  assign \new_[9061]_  = \new_[19749]_  ? \new_[17191]_  : \new_[9541]_ ;
  assign \new_[9062]_  = \new_[19518]_  ? \new_[17191]_  : \new_[9542]_ ;
  assign \new_[9063]_  = \new_[19065]_  ? \new_[17191]_  : \new_[9543]_ ;
  assign \new_[9064]_  = \new_[19699]_  ? \new_[17191]_  : \new_[9544]_ ;
  assign \new_[9065]_  = \new_[19543]_  ? \new_[17191]_  : \new_[9545]_ ;
  assign \new_[9066]_  = \new_[18722]_  ? \new_[17191]_  : \new_[9546]_ ;
  assign \new_[9067]_  = \new_[17834]_  ? \new_[17191]_  : \new_[9547]_ ;
  assign \new_[9068]_  = \new_[19086]_  ? \new_[17191]_  : \new_[9548]_ ;
  assign \new_[9069]_  = \new_[19984]_  ? \new_[17191]_  : \new_[9549]_ ;
  assign \new_[9070]_  = \new_[19214]_  ? \new_[17191]_  : \new_[9551]_ ;
  assign \new_[9071]_  = \new_[18753]_  ? \new_[17191]_  : \new_[9552]_ ;
  assign \new_[9072]_  = \new_[18103]_  ? \new_[17191]_  : \new_[9553]_ ;
  assign \new_[9073]_  = \new_[17848]_  ? \new_[17191]_  : \new_[9554]_ ;
  assign \new_[9074]_  = \new_[19386]_  ? \new_[17191]_  : \new_[9555]_ ;
  assign \new_[9075]_  = \new_[18014]_  ? \new_[17191]_  : \new_[9531]_ ;
  assign \new_[9076]_  = \new_[19010]_  ? \new_[17191]_  : \new_[9556]_ ;
  assign \new_[9077]_  = \new_[19689]_  ? \new_[17191]_  : \new_[9558]_ ;
  assign \new_[9078]_  = \new_[17982]_  ? \new_[17191]_  : \new_[9559]_ ;
  assign \new_[9079]_  = \new_[18077]_  ? \new_[16976]_  : \new_[9540]_ ;
  assign \new_[9080]_  = \new_[18198]_  ? \new_[16911]_  : \new_[9536]_ ;
  assign \new_[9081]_  = \new_[19600]_  ? \new_[16911]_  : \new_[9537]_ ;
  assign \new_[9082]_  = \new_[18929]_  ? \new_[16911]_  : \new_[9538]_ ;
  assign \new_[9083]_  = \new_[17807]_  ? \new_[16911]_  : \new_[9539]_ ;
  assign \new_[9084]_  = \new_[18581]_  ? \new_[16911]_  : \new_[9540]_ ;
  assign \new_[9085]_  = \new_[19238]_  ? \new_[16911]_  : \new_[9542]_ ;
  assign \new_[9086]_  = \new_[20000]_  ? \new_[16911]_  : \new_[9543]_ ;
  assign \new_[9087]_  = \new_[19867]_  ? \new_[16911]_  : \new_[9544]_ ;
  assign \new_[9088]_  = \new_[18384]_  ? \new_[16911]_  : \new_[9546]_ ;
  assign \new_[9089]_  = \new_[19840]_  ? \new_[16911]_  : \new_[9547]_ ;
  assign \new_[9090]_  = \new_[19677]_  ? \new_[16911]_  : \new_[9549]_ ;
  assign \new_[9091]_  = \new_[18314]_  ? \new_[16911]_  : \new_[9550]_ ;
  assign \new_[9092]_  = \new_[19110]_  ? \new_[16911]_  : \new_[9552]_ ;
  assign \new_[9093]_  = \new_[19241]_  ? \new_[16911]_  : \new_[9553]_ ;
  assign \new_[9094]_  = \new_[18093]_  ? \new_[16911]_  : \new_[9555]_ ;
  assign \new_[9095]_  = \new_[18436]_  ? \new_[16911]_  : \new_[9531]_ ;
  assign \new_[9096]_  = \new_[19252]_  ? \new_[16911]_  : \new_[9556]_ ;
  assign \new_[9097]_  = \new_[18219]_  ? \new_[16911]_  : \new_[9557]_ ;
  assign \new_[9098]_  = \new_[19033]_  ? \new_[16911]_  : \new_[9559]_ ;
  assign \new_[9099]_  = \new_[19205]_  ? \new_[16911]_  : \new_[9551]_ ;
  assign \new_[9100]_  = \new_[18585]_  ? \new_[16911]_  : \new_[9548]_ ;
  assign \new_[9101]_  = \new_[19798]_  ? \new_[16911]_  : \new_[9558]_ ;
  assign \new_[9102]_  = \new_[18961]_  ? \new_[16911]_  : \new_[9541]_ ;
  assign n6400 = \new_[18020]_  ? \new_[10324]_  : \new_[9536]_ ;
  assign n6405 = \new_[17876]_  ? \new_[10324]_  : \new_[9537]_ ;
  assign n6410 = \new_[17821]_  ? \new_[10324]_  : \new_[9538]_ ;
  assign n6415 = \new_[19563]_  ? \new_[10324]_  : \new_[9539]_ ;
  assign n6420 = \new_[17816]_  ? \new_[10324]_  : \new_[9540]_ ;
  assign n6425 = \new_[17891]_  ? \new_[10324]_  : \new_[9541]_ ;
  assign n6430 = \new_[18779]_  ? \new_[10324]_  : \new_[9542]_ ;
  assign n6525 = \new_[19578]_  ? \new_[10324]_  : \new_[9543]_ ;
  assign n6435 = \new_[18987]_  ? \new_[10324]_  : \new_[9544]_ ;
  assign n6440 = \new_[18917]_  ? \new_[10324]_  : \new_[9545]_ ;
  assign n6445 = \new_[18568]_  ? \new_[10324]_  : \new_[9546]_ ;
  assign n6530 = \new_[17863]_  ? \new_[10324]_  : \new_[9547]_ ;
  assign n6450 = \new_[19576]_  ? \new_[10324]_  : \new_[9548]_ ;
  assign n6455 = \new_[18150]_  ? \new_[10324]_  : \new_[9549]_ ;
  assign n6460 = \new_[19366]_  ? \new_[10324]_  : \new_[9550]_ ;
  assign n6465 = \new_[19349]_  ? \new_[10324]_  : \new_[9551]_ ;
  assign n6470 = \new_[18357]_  ? \new_[10324]_  : \new_[9552]_ ;
  assign n6520 = \new_[19282]_  ? \new_[10324]_  : \new_[9553]_ ;
  assign n6475 = \new_[19610]_  ? \new_[10324]_  : \new_[9554]_ ;
  assign n6480 = \new_[17854]_  ? \new_[10324]_  : \new_[9555]_ ;
  assign n6515 = \new_[18116]_  ? \new_[10324]_  : \new_[9556]_ ;
  assign n6485 = \new_[19604]_  ? \new_[10324]_  : \new_[9557]_ ;
  assign n6490 = \new_[17841]_  ? \new_[10324]_  : \new_[9558]_ ;
  assign n6495 = \new_[18047]_  ? \new_[10324]_  : \new_[9559]_ ;
  assign \new_[9127]_  = \new_[18964]_  ? \new_[16900]_  : \new_[9544]_ ;
  assign \new_[9128]_  = \new_[19652]_  ? \new_[16911]_  : \new_[9545]_ ;
  assign n6500 = ~\new_[9477]_  | ~\new_[9604]_ ;
  assign n6505 = ~\new_[9478]_  | ~\new_[9604]_ ;
  assign n6510 = ~\new_[9476]_  | (~\new_[9613]_  & ~\new_[17640]_ );
  assign \new_[9132]_  = \new_[8388]_ ;
  assign \new_[9133]_  = \new_[9239]_ ;
  assign \new_[9134]_  = ~\new_[20458]_  | ~\new_[20323]_ ;
  assign \new_[9135]_  = ~\new_[20323]_  | ~\new_[20344]_ ;
  assign \new_[9136]_  = (~\new_[20012]_  | ~\new_[17913]_ ) & (~\new_[20518]_  | ~\new_[19853]_ );
  assign \new_[9137]_  = (~\new_[9497]_  | ~\new_[18198]_ ) & (~\new_[19997]_  | ~\new_[19061]_ );
  assign \new_[9138]_  = ~\\wishbone_slave_unit_del_sync_addr_out_reg[14] ;
  assign \new_[9139]_  = (~\new_[9502]_  | ~\new_[19855]_ ) & (~\new_[9511]_  | ~\new_[18993]_ );
  assign \new_[9140]_  = (~\new_[9500]_  | ~\new_[19707]_ ) & (~\new_[9499]_  | ~\new_[19305]_ );
  assign \new_[9141]_  = ~\\wishbone_slave_unit_fifos_inGreyCount_reg[0] ;
  assign \new_[9142]_  = (~\new_[9500]_  | ~\new_[18052]_ ) & (~\new_[9499]_  | ~\new_[19592]_ );
  assign \new_[9143]_  = (~\new_[9502]_  | ~\new_[18844]_ ) & (~\new_[9511]_  | ~\new_[19561]_ );
  assign \new_[9144]_  = (~\new_[19999]_  | ~\new_[19662]_ ) & (~\new_[19997]_  | ~\new_[18058]_ );
  assign \new_[9145]_  = (~\new_[20012]_  | ~\new_[19390]_ ) & (~\new_[20518]_  | ~\new_[18343]_ );
  assign \new_[9146]_  = (~\new_[9502]_  | ~\new_[18483]_ ) & (~\new_[9511]_  | ~\new_[19157]_ );
  assign \new_[9147]_  = (~\new_[9500]_  | ~\new_[19368]_ ) & (~\new_[9499]_  | ~\new_[18216]_ );
  assign \new_[9148]_  = (~\new_[9500]_  | ~\new_[19494]_ ) & (~\new_[9499]_  | ~\new_[19191]_ );
  assign \new_[9149]_  = (~\new_[9502]_  | ~\new_[18090]_ ) & (~\new_[9511]_  | ~\new_[19257]_ );
  assign \new_[9150]_  = (~\new_[9502]_  | ~\new_[19657]_ ) & (~\new_[9511]_  | ~\new_[17850]_ );
  assign \new_[9151]_  = (~\new_[9500]_  | ~\new_[19428]_ ) & (~\new_[9499]_  | ~\new_[19405]_ );
  assign \new_[9152]_  = (~\new_[20012]_  | ~\new_[18952]_ ) & (~\new_[20518]_  | ~\new_[17977]_ );
  assign \new_[9153]_  = (~\new_[9497]_  | ~\new_[18961]_ ) & (~\new_[19997]_  | ~\new_[18891]_ );
  assign \new_[9154]_  = (~\new_[20012]_  | ~\new_[18181]_ ) & (~\new_[20518]_  | ~\new_[19832]_ );
  assign \new_[9155]_  = (~\new_[19999]_  | ~\new_[19238]_ ) & (~\new_[19997]_  | ~\new_[18682]_ );
  assign \new_[9156]_  = (~\new_[9500]_  | ~\new_[19358]_ ) & (~\new_[9499]_  | ~\new_[19700]_ );
  assign \new_[9157]_  = (~\new_[9502]_  | ~\new_[19156]_ ) & (~\new_[9511]_  | ~\new_[18631]_ );
  assign \new_[9158]_  = (~\new_[9502]_  | ~\new_[19388]_ ) & (~\new_[9511]_  | ~\new_[19144]_ );
  assign \new_[9159]_  = (~\new_[9500]_  | ~\new_[17930]_ ) & (~\new_[9499]_  | ~\new_[18214]_ );
  assign \new_[9160]_  = (~\new_[19999]_  | ~\new_[19652]_ ) & (~\new_[19997]_  | ~\new_[18736]_ );
  assign \new_[9161]_  = (~\new_[20012]_  | ~\new_[19253]_ ) & (~\new_[20518]_  | ~\new_[18569]_ );
  assign \new_[9162]_  = (~\new_[9500]_  | ~\new_[18399]_ ) & (~\new_[9499]_  | ~\new_[18692]_ );
  assign \new_[9163]_  = (~\new_[9502]_  | ~\new_[19444]_ ) & (~\new_[9511]_  | ~\new_[18315]_ );
  assign \new_[9164]_  = (~\new_[9497]_  | ~\new_[19840]_ ) & (~\new_[19997]_  | ~\new_[19602]_ );
  assign \new_[9165]_  = (~\new_[20012]_  | ~\new_[19335]_ ) & (~\new_[20518]_  | ~\new_[19109]_ );
  assign \new_[9166]_  = (~\new_[9502]_  | ~\new_[18907]_ ) & (~\new_[9511]_  | ~\new_[18851]_ );
  assign \new_[9167]_  = (~\new_[9500]_  | ~\new_[17928]_ ) & (~\new_[9499]_  | ~\new_[19656]_ );
  assign \new_[9168]_  = (~\new_[9500]_  | ~\new_[17927]_ ) & (~\new_[9499]_  | ~\new_[19247]_ );
  assign \new_[9169]_  = (~\new_[9502]_  | ~\new_[18771]_ ) & (~\new_[9511]_  | ~\new_[18018]_ );
  assign \new_[9170]_  = (~\new_[9502]_  | ~\new_[18856]_ ) & (~\new_[9511]_  | ~\new_[19055]_ );
  assign \new_[9171]_  = (~\new_[9500]_  | ~\new_[19414]_ ) & (~\new_[9499]_  | ~\new_[19149]_ );
  assign \new_[9172]_  = (~\new_[20012]_  | ~\new_[17944]_ ) & (~\new_[20518]_  | ~\new_[18460]_ );
  assign \new_[9173]_  = (~\new_[19999]_  | ~\new_[19733]_ ) & (~\new_[19997]_  | ~\new_[18724]_ );
  assign \new_[9174]_  = (~\new_[9500]_  | ~\new_[17926]_ ) & (~\new_[9499]_  | ~\new_[18906]_ );
  assign \new_[9175]_  = (~\new_[9502]_  | ~\new_[18730]_ ) & (~\new_[9511]_  | ~\new_[18641]_ );
  assign \new_[9176]_  = (~\new_[9502]_  | ~\new_[19364]_ ) & (~\new_[9511]_  | ~\new_[18394]_ );
  assign \new_[9177]_  = (~\new_[9500]_  | ~\new_[18455]_ ) & (~\new_[9499]_  | ~\new_[19824]_ );
  assign \new_[9178]_  = (~\new_[9500]_  | ~\new_[19373]_ ) & (~\new_[9499]_  | ~\new_[19394]_ );
  assign \new_[9179]_  = (~\new_[9502]_  | ~\new_[18972]_ ) & (~\new_[9511]_  | ~\new_[18899]_ );
  assign \new_[9180]_  = (~\new_[9500]_  | ~\new_[19198]_ ) & (~\new_[9499]_  | ~\new_[19047]_ );
  assign \new_[9181]_  = (~\new_[9502]_  | ~\new_[19320]_ ) & (~\new_[9511]_  | ~\new_[18225]_ );
  assign \new_[9182]_  = (~\new_[20012]_  | ~\new_[19270]_ ) & (~\new_[20518]_  | ~\new_[18877]_ );
  assign \new_[9183]_  = (~\new_[19999]_  | ~\new_[18618]_ ) & (~\new_[19997]_  | ~\new_[19245]_ );
  assign \new_[9184]_  = (~\new_[19999]_  | ~\new_[18536]_ ) & (~\new_[19997]_  | ~\new_[18675]_ );
  assign \new_[9185]_  = (~\new_[20012]_  | ~\new_[19268]_ ) & (~\new_[20518]_  | ~\new_[19276]_ );
  assign \new_[9186]_  = (~\new_[9502]_  | ~\new_[19019]_ ) & (~\new_[9511]_  | ~\new_[19265]_ );
  assign \new_[9187]_  = \new_[9270]_ ;
  assign \new_[9188]_  = ~\new_[9270]_ ;
  assign \new_[9189]_  = ~\new_[9285]_ ;
  assign \new_[9190]_  = ~\new_[9271]_ ;
  assign \new_[9191]_  = ~\\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2] ;
  assign \new_[9192]_  = ~\\wishbone_slave_unit_fifos_inGreyCount_reg[1] ;
  assign \new_[9193]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][36] ;
  assign \new_[9194]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][36] ;
  assign \new_[9195]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][36] ;
  assign \new_[9196]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][36] ;
  assign \new_[9197]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][36] ;
  assign \new_[9198]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][36] ;
  assign \new_[9199]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][36] ;
  assign \new_[9200]_  = ~\new_[9513]_  | ~\new_[9820]_ ;
  assign \new_[9201]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][36] ;
  assign \new_[9202]_  = ~\new_[20011]_ ;
  assign \new_[9203]_  = ~\new_[9293]_ ;
  assign \new_[9204]_  = \new_[9295]_ ;
  assign \new_[9205]_  = ~\new_[9295]_ ;
  assign \new_[9206]_  = ~\new_[9296]_ ;
  assign \new_[9207]_  = ~\new_[19996]_ ;
  assign \new_[9208]_  = ~\new_[9305]_ ;
  assign n6635 = \new_[16543]_  ? \new_[16604]_  : \new_[9595]_ ;
  assign n6550 = \new_[15939]_  ? \new_[16604]_  : \new_[9594]_ ;
  assign n6625 = \new_[16887]_  ? \new_[16604]_  : \new_[9596]_ ;
  assign n6555 = n16725 ? \new_[16604]_  : \new_[9597]_ ;
  assign n6560 = n17050 ? \new_[16604]_  : \new_[9598]_ ;
  assign n6630 = n17080 ? \new_[16604]_  : \new_[9599]_ ;
  assign n6565 = n17040 ? \new_[16604]_  : \new_[9600]_ ;
  assign \new_[9216]_  = ~\new_[20003]_ ;
  assign \new_[9217]_  = \new_[9601]_  ? \new_[17003]_  : \new_[18879]_ ;
  assign \new_[9218]_  = \new_[9602]_  ? \new_[17003]_  : \new_[19870]_ ;
  assign \new_[9219]_  = \new_[9601]_  ? \new_[16804]_  : \new_[17815]_ ;
  assign \new_[9220]_  = \new_[9602]_  ? \new_[16804]_  : \new_[19852]_ ;
  assign \new_[9221]_  = \new_[9601]_  ? \new_[17001]_  : \new_[19687]_ ;
  assign \new_[9222]_  = \new_[9602]_  ? \new_[17001]_  : \new_[19002]_ ;
  assign \new_[9223]_  = \new_[9601]_  ? \new_[16805]_  : \new_[18108]_ ;
  assign \new_[9224]_  = \new_[9602]_  ? \new_[16805]_  : \new_[19380]_ ;
  assign \new_[9225]_  = \new_[9601]_  ? \new_[17131]_  : \new_[18982]_ ;
  assign \new_[9226]_  = \new_[9602]_  ? \new_[17131]_  : \new_[18151]_ ;
  assign \new_[9227]_  = \new_[9601]_  ? \new_[16797]_  : \new_[19052]_ ;
  assign \new_[9228]_  = \new_[9602]_  ? \new_[16797]_  : \new_[18412]_ ;
  assign \new_[9229]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][36] ;
  assign \new_[9230]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][36] ;
  assign \new_[9231]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][36] ;
  assign \new_[9232]_  = ~\\wishbone_slave_unit_fifos_inGreyCount_reg[2] ;
  assign \new_[9233]_  = \new_[9601]_  ? \new_[16662]_  : \new_[19032]_ ;
  assign \new_[9234]_  = \new_[9602]_  ? \new_[16662]_  : \new_[18332]_ ;
  assign \new_[9235]_  = \new_[19254]_  ? \new_[16975]_  : \new_[9601]_ ;
  assign \new_[9236]_  = \new_[18040]_  ? \new_[16975]_  : \new_[9602]_ ;
  assign \new_[9237]_  = \new_[19615]_  ? \new_[16976]_  : \new_[9601]_ ;
  assign \new_[9238]_  = \new_[18540]_  ? \new_[16976]_  : \new_[9602]_ ;
  assign \new_[9239]_  = ~\new_[9272]_ ;
  assign \new_[9240]_  = \new_[19594]_  ? \new_[16900]_  : \new_[9601]_ ;
  assign \new_[9241]_  = \new_[18954]_  ? \new_[17191]_  : \new_[9601]_ ;
  assign \new_[9242]_  = \new_[18640]_  ? \new_[17191]_  : \new_[9602]_ ;
  assign \new_[9243]_  = \new_[9601]_  ? \new_[16790]_  : \new_[18657]_ ;
  assign \new_[9244]_  = \new_[9602]_  ? \new_[16790]_  : \new_[18988]_ ;
  assign \new_[9245]_  = \new_[9601]_  ? \new_[16896]_  : \new_[19180]_ ;
  assign \new_[9246]_  = \new_[9602]_  ? \new_[16896]_  : \new_[19449]_ ;
  assign \new_[9247]_  = \new_[9601]_  ? \new_[16679]_  : \new_[18264]_ ;
  assign \new_[9248]_  = \new_[9602]_  ? \new_[16679]_  : \new_[19063]_ ;
  assign \new_[9249]_  = \new_[19227]_  ? \new_[16911]_  : \new_[9601]_ ;
  assign \new_[9250]_  = \new_[18548]_  ? \new_[16911]_  : \new_[9602]_ ;
  assign \new_[9251]_  = \new_[9601]_  ? \new_[16796]_  : \new_[19822]_ ;
  assign \new_[9252]_  = \new_[9602]_  ? \new_[16796]_  : \new_[19080]_ ;
  assign \new_[9253]_  = \new_[18553]_  ? \new_[16900]_  : \new_[9602]_ ;
  assign n6620 = \new_[16189]_  ? \new_[9613]_  : \new_[8548]_ ;
  assign n6570 = \new_[16806]_  ? \new_[9613]_  : n17450;
  assign n6605 = \new_[10036]_  ? \new_[9611]_  : \new_[19590]_ ;
  assign n6575 = \new_[16523]_  ? \new_[9613]_  : \new_[8394]_ ;
  assign n6610 = \new_[10037]_  ? \new_[9694]_  : \new_[19154]_ ;
  assign n6580 = n17435 ? \new_[9613]_  : \new_[8395]_ ;
  assign n6585 = n17450 ? \new_[9613]_  : \new_[8396]_ ;
  assign n6590 = n17285 ? \new_[9613]_  : \new_[8397]_ ;
  assign n6595 = n17250 ? \new_[9613]_  : \new_[8398]_ ;
  assign n6600 = \new_[16660]_  ? \new_[9613]_  : n17285;
  assign n6615 = \new_[8394]_  ? \new_[9613]_  : n17250;
  assign n6535 = \new_[8385]_  ? \new_[9590]_  : \new_[16735]_ ;
  assign n6540 = \new_[8386]_  ? \new_[9590]_  : \new_[16800]_ ;
  assign n6545 = \new_[8387]_  ? \new_[9590]_  : \new_[16904]_ ;
  assign \new_[9268]_  = ~\\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0] ;
  assign \new_[9269]_  = i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg;
  assign \new_[9270]_  = ~\new_[9490]_ ;
  assign \new_[9271]_  = ~\new_[9820]_  | ~\new_[9588]_ ;
  assign \new_[9272]_  = ~\new_[9819]_  | ~\new_[9588]_ ;
  assign \new_[9273]_  = ~\new_[9820]_  | ~\new_[19968]_ ;
  assign n6640 = ~\new_[9568]_  | (~\new_[13215]_  & ~\new_[17656]_ );
  assign \new_[9275]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2] ;
  assign \new_[9276]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1] ;
  assign \new_[9277]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2] ;
  assign n17160 = \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0] ;
  assign n17360 = \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1] ;
  assign \new_[9280]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[0] ;
  assign \new_[9281]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[1] ;
  assign \new_[9282]_  = wishbone_slave_unit_del_sync_burst_out_reg;
  assign \new_[9283]_  = pci_target_unit_wishbone_master_addr_into_cnt_reg_reg;
  assign \new_[9284]_  = ~\new_[9492]_ ;
  assign \new_[9285]_  = ~\new_[9881]_  & ~\new_[9587]_ ;
  assign \new_[9286]_  = ~\new_[9493]_ ;
  assign \new_[9287]_  = output_backup_trdy_en_out_reg;
  assign \new_[9288]_  = ~\new_[9593]_  | ~\new_[16604]_ ;
  assign \new_[9289]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0] ;
  assign \new_[9290]_  = ~\new_[9496]_ ;
  assign \new_[9291]_  = \new_[20012]_ ;
  assign \new_[9292]_  = ~\new_[9498]_ ;
  assign \new_[9293]_  = ~\new_[9499]_ ;
  assign \new_[9294]_  = \new_[9499]_ ;
  assign \new_[9295]_  = ~\new_[9501]_ ;
  assign \new_[9296]_  = ~\new_[9503]_ ;
  assign \new_[9297]_  = ~\new_[9508]_ ;
  assign \new_[9298]_  = \new_[9509]_ ;
  assign \new_[9299]_  = \new_[9509]_ ;
  assign \new_[9300]_  = \new_[19997]_ ;
  assign \new_[9301]_  = \new_[19997]_ ;
  assign \new_[9302]_  = \new_[9510]_ ;
  assign \new_[9303]_  = \new_[9510]_ ;
  assign \new_[9304]_  = \new_[9511]_ ;
  assign \new_[9305]_  = ~\new_[9511]_ ;
  assign n6645 = \new_[11343]_  ? \new_[16604]_  : \new_[20392]_ ;
  assign \new_[9307]_  = ~\new_[9819]_  | ~\new_[19968]_ ;
  assign n6650 = ~\new_[9592]_  | (~\new_[8688]_  & ~\new_[9689]_ );
  assign n6710 = ~\new_[9592]_  | (~\new_[9141]_  & ~\new_[9689]_ );
  assign \new_[9310]_  = \new_[9650]_  ? \new_[16797]_  : \new_[19696]_ ;
  assign \new_[9311]_  = \new_[9650]_  ? \new_[17003]_  : \new_[18503]_ ;
  assign \new_[9312]_  = \new_[9650]_  ? \new_[16804]_  : \new_[18665]_ ;
  assign \new_[9313]_  = \new_[9650]_  ? \new_[17001]_  : \new_[17852]_ ;
  assign \new_[9314]_  = \new_[9650]_  ? \new_[16805]_  : \new_[17967]_ ;
  assign \new_[9315]_  = \new_[9650]_  ? \new_[17131]_  : \new_[19378]_ ;
  assign \new_[9316]_  = \new_[9651]_  ? \new_[17003]_  : \new_[18994]_ ;
  assign \new_[9317]_  = \new_[9652]_  ? \new_[17003]_  : \new_[19546]_ ;
  assign \new_[9318]_  = \new_[9653]_  ? \new_[17003]_  : \new_[19775]_ ;
  assign \new_[9319]_  = \new_[9654]_  ? \new_[17003]_  : \new_[19809]_ ;
  assign \new_[9320]_  = \new_[9655]_  ? \new_[17003]_  : \new_[18511]_ ;
  assign \new_[9321]_  = \new_[9656]_  ? \new_[17003]_  : \new_[18693]_ ;
  assign \new_[9322]_  = \new_[9657]_  ? \new_[17003]_  : \new_[18089]_ ;
  assign \new_[9323]_  = \new_[9658]_  ? \new_[17003]_  : \new_[18923]_ ;
  assign \new_[9324]_  = \new_[9651]_  ? \new_[16804]_  : \new_[18893]_ ;
  assign \new_[9325]_  = \new_[9652]_  ? \new_[16804]_  : \new_[18939]_ ;
  assign \new_[9326]_  = \new_[9653]_  ? \new_[16804]_  : \new_[18404]_ ;
  assign \new_[9327]_  = \new_[9654]_  ? \new_[16804]_  : \new_[19630]_ ;
  assign \new_[9328]_  = \new_[9655]_  ? \new_[16804]_  : \new_[18390]_ ;
  assign \new_[9329]_  = \new_[9656]_  ? \new_[16804]_  : \new_[18459]_ ;
  assign \new_[9330]_  = \new_[9657]_  ? \new_[16804]_  : \new_[18335]_ ;
  assign \new_[9331]_  = \new_[9658]_  ? \new_[16804]_  : \new_[18322]_ ;
  assign \new_[9332]_  = \new_[9651]_  ? \new_[17001]_  : \new_[19125]_ ;
  assign \new_[9333]_  = \new_[9652]_  ? \new_[17001]_  : \new_[19257]_ ;
  assign \new_[9334]_  = \new_[9653]_  ? \new_[17001]_  : \new_[18851]_ ;
  assign \new_[9335]_  = \new_[9654]_  ? \new_[17001]_  : \new_[17903]_ ;
  assign \new_[9336]_  = \new_[9655]_  ? \new_[17001]_  : \new_[18696]_ ;
  assign \new_[9337]_  = \new_[9656]_  ? \new_[17001]_  : \new_[18487]_ ;
  assign \new_[9338]_  = \new_[9657]_  ? \new_[17001]_  : \new_[18685]_ ;
  assign \new_[9339]_  = \new_[9658]_  ? \new_[17001]_  : \new_[19591]_ ;
  assign \new_[9340]_  = \new_[9651]_  ? \new_[16805]_  : \new_[19331]_ ;
  assign \new_[9341]_  = \new_[9652]_  ? \new_[16805]_  : \new_[18090]_ ;
  assign \new_[9342]_  = \new_[9653]_  ? \new_[16805]_  : \new_[18907]_ ;
  assign \new_[9343]_  = \new_[9654]_  ? \new_[16805]_  : \new_[18295]_ ;
  assign \new_[9344]_  = \new_[9655]_  ? \new_[16805]_  : \new_[18158]_ ;
  assign \new_[9345]_  = \new_[9656]_  ? \new_[16805]_  : \new_[18684]_ ;
  assign \new_[9346]_  = \new_[9657]_  ? \new_[16805]_  : \new_[18847]_ ;
  assign \new_[9347]_  = \new_[9658]_  ? \new_[16805]_  : \new_[19828]_ ;
  assign \new_[9348]_  = \new_[9651]_  ? \new_[17131]_  : \new_[18058]_ ;
  assign \new_[9349]_  = \new_[9652]_  ? \new_[17131]_  : \new_[19440]_ ;
  assign \new_[9350]_  = \new_[9653]_  ? \new_[17131]_  : \new_[19529]_ ;
  assign \new_[9351]_  = \new_[9654]_  ? \new_[17131]_  : \new_[18724]_ ;
  assign \new_[9352]_  = \new_[9655]_  ? \new_[17131]_  : \new_[19245]_ ;
  assign \new_[9353]_  = \new_[9656]_  ? \new_[17131]_  : \new_[18054]_ ;
  assign \new_[9354]_  = \new_[9657]_  ? \new_[17131]_  : \new_[18022]_ ;
  assign \new_[9355]_  = \new_[9658]_  ? \new_[17131]_  : \new_[19477]_ ;
  assign \new_[9356]_  = \new_[9651]_  ? \new_[16797]_  : \new_[18205]_ ;
  assign \new_[9357]_  = \new_[9652]_  ? \new_[16797]_  : \new_[19580]_ ;
  assign \new_[9358]_  = \new_[9653]_  ? \new_[16797]_  : \new_[19418]_ ;
  assign \new_[9359]_  = \new_[9654]_  ? \new_[16797]_  : \new_[18639]_ ;
  assign \new_[9360]_  = \new_[9655]_  ? \new_[16797]_  : \new_[19793]_ ;
  assign \new_[9361]_  = \new_[9656]_  ? \new_[16797]_  : \new_[17893]_ ;
  assign \new_[9362]_  = \new_[9657]_  ? \new_[16797]_  : \new_[18184]_ ;
  assign \new_[9363]_  = \new_[9658]_  ? \new_[16797]_  : \new_[18775]_ ;
  assign \new_[9364]_  = \new_[9656]_  ? \new_[16896]_  : \new_[18124]_ ;
  assign \new_[9365]_  = \new_[9651]_  ? \new_[16662]_  : \new_[18343]_ ;
  assign \new_[9366]_  = \new_[9652]_  ? \new_[16662]_  : \new_[19519]_ ;
  assign \new_[9367]_  = \new_[9653]_  ? \new_[16662]_  : \new_[18608]_ ;
  assign \new_[9368]_  = \new_[9654]_  ? \new_[16662]_  : \new_[18460]_ ;
  assign \new_[9369]_  = \new_[9655]_  ? \new_[16662]_  : \new_[18877]_ ;
  assign \new_[9370]_  = \new_[9656]_  ? \new_[16662]_  : \new_[18921]_ ;
  assign \new_[9371]_  = \new_[9657]_  ? \new_[16662]_  : \new_[19655]_ ;
  assign \new_[9372]_  = \new_[9658]_  ? \new_[16662]_  : \new_[19817]_ ;
  assign \new_[9373]_  = \new_[9651]_  ? \new_[16790]_  : \new_[18741]_ ;
  assign \new_[9374]_  = \new_[9652]_  ? \new_[16790]_  : \new_[19191]_ ;
  assign \new_[9375]_  = \new_[9653]_  ? \new_[16790]_  : \new_[19656]_ ;
  assign \new_[9376]_  = \new_[9654]_  ? \new_[16790]_  : \new_[18978]_ ;
  assign \new_[9377]_  = \new_[9655]_  ? \new_[16790]_  : \new_[18506]_ ;
  assign \new_[9378]_  = \new_[9656]_  ? \new_[16790]_  : \new_[18421]_ ;
  assign \new_[9379]_  = \new_[9657]_  ? \new_[16790]_  : \new_[19094]_ ;
  assign \new_[9380]_  = \new_[9658]_  ? \new_[16790]_  : \new_[19846]_ ;
  assign \new_[9381]_  = \new_[9651]_  ? \new_[16896]_  : \new_[18541]_ ;
  assign \new_[9382]_  = \new_[9652]_  ? \new_[16896]_  : \new_[19494]_ ;
  assign \new_[9383]_  = \new_[9653]_  ? \new_[16896]_  : \new_[17928]_ ;
  assign \new_[9384]_  = \new_[9654]_  ? \new_[16896]_  : \new_[19755]_ ;
  assign \new_[9385]_  = \new_[9655]_  ? \new_[16896]_  : \new_[18440]_ ;
  assign \new_[9386]_  = \new_[9657]_  ? \new_[16896]_  : \new_[17918]_ ;
  assign \new_[9387]_  = \new_[9658]_  ? \new_[16896]_  : \new_[18457]_ ;
  assign \new_[9388]_  = \new_[9651]_  ? \new_[16679]_  : \new_[19390]_ ;
  assign \new_[9389]_  = \new_[9652]_  ? \new_[16679]_  : \new_[19288]_ ;
  assign \new_[9390]_  = \new_[9653]_  ? \new_[16679]_  : \new_[18007]_ ;
  assign \new_[9391]_  = \new_[9654]_  ? \new_[16679]_  : \new_[17944]_ ;
  assign \new_[9392]_  = \new_[9655]_  ? \new_[16679]_  : \new_[19270]_ ;
  assign \new_[9393]_  = \new_[9656]_  ? \new_[16679]_  : \new_[18171]_ ;
  assign \new_[9394]_  = \new_[9657]_  ? \new_[16679]_  : \new_[19454]_ ;
  assign \new_[9395]_  = \new_[9658]_  ? \new_[16679]_  : \new_[19569]_ ;
  assign \new_[9396]_  = \new_[9651]_  ? \new_[16796]_  : \new_[18115]_ ;
  assign \new_[9397]_  = \new_[9652]_  ? \new_[16796]_  : \new_[19313]_ ;
  assign \new_[9398]_  = \new_[9653]_  ? \new_[16796]_  : \new_[19712]_ ;
  assign \new_[9399]_  = \new_[9654]_  ? \new_[16796]_  : \new_[19018]_ ;
  assign \new_[9400]_  = \new_[9655]_  ? \new_[16796]_  : \new_[19056]_ ;
  assign \new_[9401]_  = \new_[9656]_  ? \new_[16796]_  : \new_[18666]_ ;
  assign \new_[9402]_  = \new_[9657]_  ? \new_[16796]_  : \new_[19027]_ ;
  assign \new_[9403]_  = \new_[9658]_  ? \new_[16796]_  : \new_[18554]_ ;
  assign \new_[9404]_  = \new_[9650]_  ? \new_[16790]_  : \new_[18976]_ ;
  assign \new_[9405]_  = \new_[9650]_  ? \new_[16796]_  : \new_[18507]_ ;
  assign \new_[9406]_  = \new_[19558]_  ? \new_[16911]_  : \new_[9650]_ ;
  assign \new_[9407]_  = \new_[9650]_  ? \new_[16662]_  : \new_[18296]_ ;
  assign \new_[9408]_  = \new_[17981]_  ? \new_[16975]_  : \new_[9651]_ ;
  assign \new_[9409]_  = \new_[19289]_  ? \new_[16975]_  : \new_[9652]_ ;
  assign \new_[9410]_  = \new_[18057]_  ? \new_[16975]_  : \new_[9653]_ ;
  assign \new_[9411]_  = \new_[19189]_  ? \new_[16975]_  : \new_[9654]_ ;
  assign \new_[9412]_  = \new_[19337]_  ? \new_[16975]_  : \new_[9655]_ ;
  assign \new_[9413]_  = \new_[18081]_  ? \new_[16975]_  : \new_[9650]_ ;
  assign \new_[9414]_  = \new_[18245]_  ? \new_[16975]_  : \new_[9656]_ ;
  assign \new_[9415]_  = \new_[18828]_  ? \new_[16975]_  : \new_[9657]_ ;
  assign \new_[9416]_  = \new_[19181]_  ? \new_[16975]_  : \new_[9658]_ ;
  assign \new_[9417]_  = \new_[19842]_  ? \new_[16976]_  : \new_[9651]_ ;
  assign \new_[9418]_  = \new_[18303]_  ? \new_[16976]_  : \new_[9652]_ ;
  assign \new_[9419]_  = \new_[18234]_  ? \new_[16976]_  : \new_[9653]_ ;
  assign \new_[9420]_  = \new_[18072]_  ? \new_[16976]_  : \new_[9654]_ ;
  assign \new_[9421]_  = \new_[18762]_  ? \new_[16976]_  : \new_[9650]_ ;
  assign \new_[9422]_  = \new_[18272]_  ? \new_[16976]_  : \new_[9656]_ ;
  assign \new_[9423]_  = \new_[18758]_  ? \new_[16976]_  : \new_[9657]_ ;
  assign \new_[9424]_  = \new_[18977]_  ? \new_[16976]_  : \new_[9658]_ ;
  assign \new_[9425]_  = \new_[18738]_  ? \new_[16900]_  : \new_[9651]_ ;
  assign \new_[9426]_  = \new_[19823]_  ? \new_[16900]_  : \new_[9652]_ ;
  assign \new_[9427]_  = \new_[19371]_  ? \new_[16900]_  : \new_[9653]_ ;
  assign \new_[9428]_  = \new_[18434]_  ? \new_[16900]_  : \new_[9654]_ ;
  assign \new_[9429]_  = \new_[18204]_  ? \new_[16900]_  : \new_[9655]_ ;
  assign \new_[9430]_  = \new_[18676]_  ? \new_[16900]_  : \new_[9650]_ ;
  assign \new_[9431]_  = \new_[18297]_  ? \new_[16900]_  : \new_[9656]_ ;
  assign \new_[9432]_  = \new_[18153]_  ? \new_[16900]_  : \new_[9657]_ ;
  assign \new_[9433]_  = \new_[19404]_  ? \new_[16900]_  : \new_[9658]_ ;
  assign \new_[9434]_  = \new_[19242]_  ? \new_[17191]_  : \new_[9651]_ ;
  assign \new_[9435]_  = \new_[18301]_  ? \new_[17191]_  : \new_[9652]_ ;
  assign \new_[9436]_  = \new_[17833]_  ? \new_[17191]_  : \new_[9653]_ ;
  assign \new_[9437]_  = \new_[17832]_  ? \new_[17191]_  : \new_[9654]_ ;
  assign \new_[9438]_  = \new_[18759]_  ? \new_[17191]_  : \new_[9655]_ ;
  assign \new_[9439]_  = \new_[19760]_  ? \new_[17191]_  : \new_[9650]_ ;
  assign \new_[9440]_  = \new_[19719]_  ? \new_[17191]_  : \new_[9656]_ ;
  assign \new_[9441]_  = \new_[19025]_  ? \new_[17191]_  : \new_[9657]_ ;
  assign \new_[9442]_  = \new_[18966]_  ? \new_[17191]_  : \new_[9658]_ ;
  assign \new_[9443]_  = \new_[9650]_  ? \new_[16896]_  : \new_[19336]_ ;
  assign \new_[9444]_  = \new_[9650]_  ? \new_[16679]_  : \new_[18286]_ ;
  assign \new_[9445]_  = \new_[19091]_  ? \new_[16976]_  : \new_[9655]_ ;
  assign \new_[9446]_  = \new_[19132]_  ? \new_[16911]_  : \new_[9652]_ ;
  assign \new_[9447]_  = \new_[18769]_  ? \new_[16911]_  : \new_[9653]_ ;
  assign \new_[9448]_  = \new_[19733]_  ? \new_[16911]_  : \new_[9654]_ ;
  assign \new_[9449]_  = \new_[18618]_  ? \new_[16911]_  : \new_[9655]_ ;
  assign \new_[9450]_  = \new_[19649]_  ? \new_[16911]_  : \new_[9657]_ ;
  assign \new_[9451]_  = \new_[18402]_  ? \new_[16911]_  : \new_[9658]_ ;
  assign \new_[9452]_  = \new_[19662]_  ? \new_[16911]_  : \new_[9651]_ ;
  assign \new_[9453]_  = \new_[18873]_  ? \new_[16911]_  : \new_[9656]_ ;
  assign n6655 = \new_[17810]_  ? \new_[10324]_  : \new_[9651]_ ;
  assign n6705 = \new_[19564]_  ? \new_[10324]_  : \new_[9652]_ ;
  assign n6660 = \new_[19572]_  ? \new_[10324]_  : \new_[9653]_ ;
  assign n6695 = \new_[19409]_  ? \new_[10324]_  : \new_[9654]_ ;
  assign n6665 = \new_[19296]_  ? \new_[10324]_  : \new_[9655]_ ;
  assign n6675 = \new_[19614]_  ? \new_[10324]_  : \new_[9656]_ ;
  assign n6670 = \new_[17844]_  ? \new_[10324]_  : \new_[9657]_ ;
  assign n6700 = \new_[18748]_  ? \new_[10324]_  : \new_[9658]_ ;
  assign \new_[9462]_  = ~\new_[9603]_  & ~\new_[16662]_ ;
  assign \new_[9463]_  = ~\new_[9603]_  & ~\new_[17003]_ ;
  assign \new_[9464]_  = ~\new_[9603]_  & ~\new_[16804]_ ;
  assign \new_[9465]_  = ~\new_[9603]_  & ~\new_[16790]_ ;
  assign \new_[9466]_  = ~\new_[9603]_  & ~\new_[16896]_ ;
  assign \new_[9467]_  = ~\new_[9603]_  & ~\new_[17001]_ ;
  assign \new_[9468]_  = ~\new_[9603]_  & ~\new_[16679]_ ;
  assign \new_[9469]_  = ~\new_[9603]_  & ~\new_[16805]_ ;
  assign \new_[9470]_  = ~\new_[9603]_  & ~\new_[17131]_ ;
  assign \new_[9471]_  = ~\new_[9603]_  & ~\new_[16796]_ ;
  assign \new_[9472]_  = ~\new_[9603]_  & ~\new_[16797]_ ;
  assign n6680 = \new_[10027]_  ? \new_[9669]_  : \new_[19285]_ ;
  assign n6685 = \new_[10035]_  ? \new_[9661]_  : \new_[19763]_ ;
  assign n6690 = \new_[10038]_  ? \new_[9661]_  : \new_[19692]_ ;
  assign \new_[9476]_  = ~\new_[9613]_  | ~\new_[17640]_ ;
  assign \new_[9477]_  = ~\new_[9612]_  | ~\new_[8224]_ ;
  assign \new_[9478]_  = ~\new_[9613]_  | ~n17435;
  assign \new_[9479]_  = ~\new_[9612]_  | ~\new_[18220]_ ;
  assign \new_[9480]_  = ~\new_[9612]_  | ~\new_[18747]_ ;
  assign \new_[9481]_  = ~\new_[9612]_  | ~\new_[19172]_ ;
  assign \new_[9482]_  = ~\new_[9612]_  | ~\new_[17813]_ ;
  assign \new_[9483]_  = ~\new_[9612]_  | ~\new_[17969]_ ;
  assign \new_[9484]_  = ~\new_[9612]_  | ~\new_[18956]_ ;
  assign \new_[9485]_  = ~\new_[9612]_  | ~\new_[18339]_ ;
  assign n17185 = \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2] ;
  assign \new_[9487]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[2] ;
  assign \new_[9488]_  = \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1] ;
  assign pci_trdy_oe_o = pci_io_mux_trdy_iob_en_out_reg;
  assign \new_[9490]_  = ~\new_[9819]_  | ~\new_[9646]_ ;
  assign \new_[9491]_  = ~\new_[9820]_  | ~\new_[9646]_ ;
  assign \new_[9492]_  = \new_[9642]_  | \new_[20531]_ ;
  assign \new_[9493]_  = ~\new_[9567]_ ;
  assign pci_stop_oe_o = pci_io_mux_stop_iob_en_out_reg;
  assign pci_devsel_oe_o = pci_io_mux_devsel_iob_en_out_reg;
  assign \new_[9496]_  = ~\new_[20193]_  | ~\new_[20445]_ ;
  assign \new_[9497]_  = ~\new_[20468]_ ;
  assign \new_[9498]_  = ~\new_[19987]_ ;
  assign \new_[9499]_  = ~\new_[9570]_ ;
  assign \new_[9500]_  = ~\new_[9571]_ ;
  assign \new_[9501]_  = ~\new_[9683]_  | ~\new_[19960]_ ;
  assign \new_[9502]_  = ~\new_[9572]_ ;
  assign \new_[9503]_  = ~\new_[9573]_ ;
  assign \new_[9504]_  = ~\new_[9573]_ ;
  assign \new_[9505]_  = ~\new_[9573]_ ;
  assign \new_[9506]_  = ~\new_[9573]_ ;
  assign \new_[9507]_  = ~\new_[9573]_ ;
  assign \new_[9508]_  = ~\new_[19960]_  | ~\new_[9682]_ ;
  assign \new_[9509]_  = ~\new_[9574]_ ;
  assign \new_[9510]_  = ~\new_[9575]_ ;
  assign \new_[9511]_  = ~\new_[9576]_ ;
  assign \new_[9512]_  = ~\new_[20346]_ ;
  assign \new_[9513]_  = ~\new_[9587]_ ;
  assign n6715 = \new_[19273]_  ? \new_[9689]_  : \new_[16145]_ ;
  assign n6720 = n17015 ? \new_[9689]_  : \new_[17034]_ ;
  assign n6780 = n17005 ? \new_[9689]_  : \new_[19273]_ ;
  assign n6785 = \new_[18890]_  ^ \new_[9689]_ ;
  assign n6725 = \new_[10026]_  ? \new_[9745]_  : \new_[18967]_ ;
  assign n6760 = \new_[10028]_  ? \new_[9745]_  : \new_[18475]_ ;
  assign n6730 = \new_[10029]_  ? \new_[9733]_  : \new_[18409]_ ;
  assign n6735 = \new_[10030]_  ? \new_[9733]_  : \new_[18427]_ ;
  assign n6740 = \new_[10031]_  ? \new_[9716]_  : \new_[18492]_ ;
  assign n6775 = \new_[10032]_  ? \new_[9730]_  : \new_[18382]_ ;
  assign n6770 = \new_[10033]_  ? \new_[9716]_  : \new_[17943]_ ;
  assign n6745 = \new_[10034]_  ? \new_[9730]_  : \new_[19750]_ ;
  assign n6750 = \new_[10039]_  ? \new_[9755]_  : \new_[19640]_ ;
  assign n6755 = \new_[10040]_  ? \new_[9733]_  : \new_[18886]_ ;
  assign n6765 = \new_[10041]_  ? \new_[9730]_  : \new_[18518]_ ;
  assign \new_[9529]_  = ~\new_[20190]_ ;
  assign \new_[9530]_  = ~\new_[20462]_ ;
  assign \new_[9531]_  = ~\new_[9603]_ ;
  assign \new_[9532]_  = ~\new_[9663]_  | ~\new_[18499]_ ;
  assign \new_[9533]_  = ~\new_[9663]_  | ~\new_[19626]_ ;
  assign \new_[9534]_  = ~\new_[9663]_  | ~\new_[18701]_ ;
  assign \new_[9535]_  = ~\new_[9663]_  | ~\new_[19152]_ ;
  assign \new_[9536]_  = \new_[13679]_  ? \new_[9979]_  : \new_[18041]_ ;
  assign \new_[9537]_  = \new_[6304]_  ? \new_[9760]_  : \new_[19197]_ ;
  assign \new_[9538]_  = \new_[6303]_  ? \new_[9760]_  : \new_[18063]_ ;
  assign \new_[9539]_  = \new_[6305]_  ? \new_[9979]_  : \new_[17858]_ ;
  assign \new_[9540]_  = \new_[6307]_  ? \new_[9979]_  : \new_[17814]_ ;
  assign \new_[9541]_  = \new_[6308]_  ? \new_[9979]_  : \new_[18075]_ ;
  assign \new_[9542]_  = \new_[6309]_  ? \new_[9979]_  : \new_[19038]_ ;
  assign \new_[9543]_  = \new_[6329]_  ? \new_[9760]_  : \new_[18678]_ ;
  assign \new_[9544]_  = \new_[6310]_  ? \new_[9760]_  : \new_[19143]_ ;
  assign \new_[9545]_  = \new_[13686]_  ? \new_[9760]_  : \new_[18102]_ ;
  assign \new_[9546]_  = \new_[6311]_  ? \new_[9979]_  : \new_[18156]_ ;
  assign \new_[9547]_  = \new_[6312]_  ? \new_[9979]_  : \new_[18099]_ ;
  assign \new_[9548]_  = \new_[6313]_  ? \new_[9760]_  : \new_[18227]_ ;
  assign \new_[9549]_  = \new_[6314]_  ? \new_[9979]_  : \new_[18839]_ ;
  assign \new_[9550]_  = \new_[6552]_  ? \new_[9979]_  : \new_[18628]_ ;
  assign \new_[9551]_  = \new_[6316]_  ? \new_[9979]_  : \new_[17824]_ ;
  assign \new_[9552]_  = \new_[6326]_  ? \new_[9760]_  : \new_[17884]_ ;
  assign \new_[9553]_  = \new_[18545]_  ? \new_[9979]_  : \new_[17860]_ ;
  assign \new_[9554]_  = \new_[6319]_  ? \new_[9979]_  : \new_[18406]_ ;
  assign \new_[9555]_  = \new_[17959]_  ? \new_[9979]_  : \new_[18290]_ ;
  assign \new_[9556]_  = \new_[6321]_  ? \new_[9760]_  : \new_[18520]_ ;
  assign \new_[9557]_  = \new_[6324]_  ? \new_[9979]_  : \new_[18733]_ ;
  assign \new_[9558]_  = \new_[6551]_  ? \new_[9979]_  : \new_[18814]_ ;
  assign \new_[9559]_  = \new_[6325]_  ? \new_[9979]_  : \new_[18260]_ ;
  assign \new_[9560]_  = ~\new_[9901]_  | ~\wbm_adr_o[0] ;
  assign \new_[9561]_  = ~\new_[9901]_  | ~\wbm_adr_o[1] ;
  assign \new_[9562]_  = \\pci_target_unit_wishbone_master_rty_counter_reg[0] ;
  assign n6845 = \new_[17656]_  ? \new_[13215]_  : \new_[9820]_ ;
  assign n6840 = ~n6875;
  assign \new_[9565]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0] ;
  assign n6790 = (~\new_[9829]_  & ~wbs_err_o) | (~wbs_stb_i & ~\new_[17475]_ );
  assign \new_[9567]_  = ~\new_[9642]_ ;
  assign \new_[9568]_  = ~\new_[9686]_  | ~\new_[13215]_ ;
  assign \new_[9569]_  = ~\new_[20445]_  | ~\new_[9690]_ ;
  assign \new_[9570]_  = ~\new_[9682]_  | ~\new_[9690]_ ;
  assign \new_[9571]_  = ~\new_[20445]_  | ~\new_[20471]_ ;
  assign \new_[9572]_  = ~\new_[20470]_  | ~\new_[9690]_ ;
  assign \new_[9573]_  = ~\new_[9691]_  | ~\new_[20445]_ ;
  assign \new_[9574]_  = ~\new_[9691]_  | ~\new_[9682]_ ;
  assign \new_[9575]_  = ~\new_[9683]_  | ~\new_[9691]_ ;
  assign \new_[9576]_  = ~\new_[20471]_  | ~\new_[9682]_ ;
  assign n6795 = \new_[15967]_  ? \new_[13215]_  : \new_[9833]_ ;
  assign n6860 = \new_[17002]_  ? \new_[13215]_  : \new_[9836]_ ;
  assign n6800 = \new_[10004]_  ? \new_[13215]_  : \new_[19973]_ ;
  assign n6805 = \new_[10074]_  ? \new_[13215]_  : \new_[19972]_ ;
  assign n6810 = n17065 ? \new_[13215]_  : \new_[9837]_ ;
  assign n6815 = n17035 ? \new_[13215]_  : \new_[9838]_ ;
  assign n6850 = n17020 ? \new_[13215]_  : \new_[9839]_ ;
  assign n6820 = \new_[10012]_  ? \new_[13215]_  : \new_[9840]_ ;
  assign n6825 = \new_[10006]_  ? \new_[13215]_  : \new_[9842]_ ;
  assign n6855 = \new_[10077]_  ? \new_[13215]_  : \new_[9841]_ ;
  assign \new_[9587]_  = ~\new_[9688]_  | ~\new_[9687]_ ;
  assign \new_[9588]_  = ~\new_[9688]_  & ~\new_[19973]_ ;
  assign n6830 = ~\new_[10019]_  | ~\new_[9685]_ ;
  assign \new_[9590]_  = ~\new_[16510]_  | ~\new_[17257]_  | ~\new_[9681]_  | ~\new_[16584]_ ;
  assign \new_[9591]_  = ~\\wishbone_slave_unit_del_sync_bc_out_reg[3] ;
  assign \new_[9592]_  = ~\new_[17009]_  | ~\new_[9689]_ ;
  assign \new_[9593]_  = \new_[19683]_  ^ \new_[20100]_ ;
  assign \new_[9594]_  = \new_[20288]_  ? \new_[20100]_  : \new_[16696]_ ;
  assign \new_[9595]_  = \new_[18185]_  ? \new_[20100]_  : \new_[16175]_ ;
  assign \new_[9596]_  = \new_[20188]_  ? \new_[20100]_  : \new_[17014]_ ;
  assign \new_[9597]_  = \new_[8390]_  ? \new_[20100]_  : \new_[17107]_ ;
  assign \new_[9598]_  = \new_[8391]_  ? \new_[20100]_  : \new_[17431]_ ;
  assign \new_[9599]_  = \new_[8603]_  ? \new_[20100]_  : \new_[17105]_ ;
  assign \new_[9600]_  = \new_[8392]_  ? \new_[20100]_  : \new_[18680]_ ;
  assign \new_[9601]_  = ~\new_[18589]_  | ~\new_[9692]_  | ~\new_[9979]_ ;
  assign \new_[9602]_  = ~\new_[18288]_  | ~\new_[9692]_  | ~\new_[9979]_ ;
  assign \new_[9603]_  = ~\new_[9693]_  | ~\new_[9692]_ ;
  assign \new_[9604]_  = \new_[16981]_  | \new_[9694]_ ;
  assign \new_[9605]_  = ~\new_[9659]_ ;
  assign \new_[9606]_  = ~\new_[9659]_ ;
  assign \new_[9607]_  = ~\new_[9659]_ ;
  assign \new_[9608]_  = ~\new_[9659]_ ;
  assign \new_[9609]_  = ~\new_[9659]_ ;
  assign \new_[9610]_  = ~\new_[9659]_ ;
  assign \new_[9611]_  = ~\new_[9659]_ ;
  assign \new_[9612]_  = ~\new_[9854]_ ;
  assign \new_[9613]_  = ~\new_[9854]_ ;
  assign \new_[9614]_  = ~\new_[9761]_  & ~\new_[20499]_ ;
  assign \new_[9615]_  = ~\new_[9813]_  | (~\new_[15688]_  & ~\new_[16436]_ );
  assign \new_[9616]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0] ;
  assign \new_[9617]_  = output_backup_frame_out_reg;
  assign \new_[9618]_  = \\pci_target_unit_wishbone_master_rty_counter_reg[5] ;
  assign \new_[9619]_  = \\pci_target_unit_wishbone_master_rty_counter_reg[6] ;
  assign \new_[9620]_  = ~\\wishbone_slave_unit_del_sync_bc_out_reg[2] ;
  assign \new_[9621]_  = \\pci_target_unit_wishbone_master_rty_counter_reg[1] ;
  assign \new_[9622]_  = \\pci_target_unit_wishbone_master_rty_counter_reg[2] ;
  assign \new_[9623]_  = \\pci_target_unit_wishbone_master_rty_counter_reg[4] ;
  assign \new_[9624]_  = \\wishbone_slave_unit_fifos_outGreyCount_reg[0] ;
  assign \new_[9625]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2] ;
  assign \new_[9626]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3] ;
  assign \new_[9627]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1] ;
  assign \new_[9628]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2] ;
  assign \new_[9629]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[0] ;
  assign \new_[9630]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[1] ;
  assign \new_[9631]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[2] ;
  assign \new_[9632]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[0] ;
  assign \new_[9633]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[1] ;
  assign \new_[9634]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[2] ;
  assign \new_[9635]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[0] ;
  assign \new_[9636]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[2] ;
  assign \new_[9637]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[3] ;
  assign \new_[9638]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[3] ;
  assign \new_[9639]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[1] ;
  assign \new_[9640]_  = ~\\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[3] ;
  assign \new_[9641]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3] ;
  assign \new_[9642]_  = ~\new_[10973]_  & ~\new_[9830]_ ;
  assign \new_[9643]_  = ~\new_[17914]_  | ~\new_[16214]_  | ~\new_[9918]_  | ~\new_[15849]_ ;
  assign \new_[9644]_  = \\pci_target_unit_wishbone_master_rty_counter_reg[3] ;
  assign n6880 = ~\new_[9888]_  | ~\new_[9834]_ ;
  assign \new_[9646]_  = \new_[19972]_  & \new_[19973]_ ;
  assign \new_[9647]_  = \\pci_target_unit_wishbone_master_rty_counter_reg[7] ;
  assign pci_frame_o = pci_io_mux_frame_iob_dat_out_reg;
  assign n6875 = ~\new_[15499]_  & ~\new_[9814]_ ;
  assign \new_[9650]_  = ~\new_[9853]_  & (~\new_[9979]_  | ~\new_[18596]_ );
  assign \new_[9651]_  = \new_[6317]_  ? \new_[9979]_  : \new_[19123]_ ;
  assign \new_[9652]_  = \new_[6306]_  ? \new_[9979]_  : \new_[17894]_ ;
  assign \new_[9653]_  = \new_[6328]_  ? \new_[9979]_  : \new_[18035]_ ;
  assign \new_[9654]_  = \new_[6315]_  ? \new_[9979]_  : \new_[19250]_ ;
  assign \new_[9655]_  = \new_[6554]_  ? \new_[9979]_  : \new_[18441]_ ;
  assign \new_[9656]_  = \new_[6553]_  ? \new_[9979]_  : \new_[18843]_ ;
  assign \new_[9657]_  = \new_[6322]_  ? \new_[9979]_  : \new_[18277]_ ;
  assign \new_[9658]_  = \new_[6323]_  ? \new_[9979]_  : \new_[19069]_ ;
  assign \new_[9659]_  = ~\new_[9694]_ ;
  assign \new_[9660]_  = ~\new_[9695]_ ;
  assign \new_[9661]_  = ~\new_[9695]_ ;
  assign \new_[9662]_  = ~\new_[9696]_ ;
  assign \new_[9663]_  = ~\new_[9696]_ ;
  assign \new_[9664]_  = ~\new_[9696]_ ;
  assign \new_[9665]_  = ~\new_[9696]_ ;
  assign \new_[9666]_  = ~\new_[9696]_ ;
  assign \new_[9667]_  = ~\new_[9697]_ ;
  assign \new_[9668]_  = ~\new_[9697]_ ;
  assign \new_[9669]_  = ~\new_[9697]_ ;
  assign \new_[9670]_  = ~\new_[9697]_ ;
  assign \new_[9671]_  = ~pci_target_unit_pci_target_sm_rd_request_reg;
  assign \new_[9672]_  = pci_target_unit_pci_target_sm_rd_progress_reg;
  assign \new_[9673]_  = \\wishbone_slave_unit_del_sync_be_out_reg[0] ;
  assign \new_[9674]_  = \\wishbone_slave_unit_del_sync_be_out_reg[1] ;
  assign \new_[9675]_  = \\wishbone_slave_unit_del_sync_be_out_reg[2] ;
  assign \new_[9676]_  = ~wishbone_slave_unit_del_sync_we_out_reg;
  assign \new_[9677]_  = ~\\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[1] ;
  assign \new_[9678]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1] ;
  assign \new_[9679]_  = \\wishbone_slave_unit_del_sync_be_out_reg[3] ;
  assign \new_[9680]_  = ~\\wishbone_slave_unit_del_sync_bc_out_reg[1] ;
  assign \new_[9681]_  = ~\new_[9814]_ ;
  assign \new_[9682]_  = \new_[20449]_  & \new_[20447]_ ;
  assign \new_[9683]_  = \new_[9885]_  & \new_[20446]_ ;
  assign n6890 = ~\new_[9887]_  | (~\new_[10324]_  & ~\new_[9591]_ );
  assign \new_[9685]_  = ~\new_[10021]_  | ~\new_[15612]_  | ~\new_[20509]_  | ~\new_[20532]_ ;
  assign \new_[9686]_  = ~\new_[9886]_  | (~\new_[10020]_  & ~\new_[18056]_ );
  assign \new_[9687]_  = ~\new_[19973]_ ;
  assign \new_[9688]_  = ~\new_[19972]_ ;
  assign \new_[9689]_  = ~\new_[9895]_  & ~\new_[11150]_ ;
  assign \new_[9690]_  = \new_[20472]_  & \new_[20474]_ ;
  assign \new_[9691]_  = ~\new_[20472]_  & ~n7075;
  assign \new_[9692]_  = ~\new_[9853]_ ;
  assign \new_[9693]_  = ~\new_[9899]_  & ~\new_[18594]_ ;
  assign \new_[9694]_  = ~\new_[9854]_ ;
  assign \new_[9695]_  = \new_[9854]_ ;
  assign \new_[9696]_  = \new_[9854]_ ;
  assign \new_[9697]_  = \new_[9854]_ ;
  assign \new_[9698]_  = ~\new_[9896]_ ;
  assign \new_[9699]_  = ~\new_[9856]_ ;
  assign \new_[9700]_  = ~\new_[9856]_ ;
  assign \new_[9701]_  = ~\new_[9856]_ ;
  assign \new_[9702]_  = ~\new_[9856]_ ;
  assign \new_[9703]_  = ~\new_[9856]_ ;
  assign \new_[9704]_  = ~\new_[9856]_ ;
  assign \new_[9705]_  = ~\new_[9855]_ ;
  assign \new_[9706]_  = ~\new_[9855]_ ;
  assign \new_[9707]_  = ~\new_[9855]_ ;
  assign \new_[9708]_  = ~\new_[9855]_ ;
  assign \new_[9709]_  = ~\new_[9855]_ ;
  assign \new_[9710]_  = ~\new_[9855]_ ;
  assign \new_[9711]_  = ~\new_[9855]_ ;
  assign \new_[9712]_  = ~\new_[9855]_ ;
  assign \new_[9713]_  = ~\new_[9856]_ ;
  assign \new_[9714]_  = ~\new_[9856]_ ;
  assign \new_[9715]_  = ~\new_[9856]_ ;
  assign \new_[9716]_  = ~\new_[9856]_ ;
  assign \new_[9717]_  = ~\new_[9856]_ ;
  assign \new_[9718]_  = ~\new_[9856]_ ;
  assign \new_[9719]_  = ~\new_[9856]_ ;
  assign \new_[9720]_  = ~\new_[9856]_ ;
  assign \new_[9721]_  = ~\new_[9855]_ ;
  assign \new_[9722]_  = ~\new_[9855]_ ;
  assign \new_[9723]_  = ~\new_[9855]_ ;
  assign \new_[9724]_  = ~\new_[9855]_ ;
  assign \new_[9725]_  = ~\new_[9855]_ ;
  assign \new_[9726]_  = ~\new_[9855]_ ;
  assign \new_[9727]_  = ~\new_[9855]_ ;
  assign \new_[9728]_  = ~\new_[9855]_ ;
  assign \new_[9729]_  = ~\new_[9857]_ ;
  assign \new_[9730]_  = ~\new_[9857]_ ;
  assign \new_[9731]_  = ~\new_[9857]_ ;
  assign \new_[9732]_  = ~\new_[9857]_ ;
  assign \new_[9733]_  = ~\new_[9857]_ ;
  assign \new_[9734]_  = ~\new_[9857]_ ;
  assign \new_[9735]_  = ~\new_[9855]_ ;
  assign \new_[9736]_  = ~\new_[9855]_ ;
  assign \new_[9737]_  = ~\new_[9855]_ ;
  assign \new_[9738]_  = ~\new_[9855]_ ;
  assign \new_[9739]_  = ~\new_[9855]_ ;
  assign \new_[9740]_  = ~\new_[9856]_ ;
  assign \new_[9741]_  = ~\new_[9856]_ ;
  assign \new_[9742]_  = ~\new_[9856]_ ;
  assign \new_[9743]_  = ~\new_[9856]_ ;
  assign \new_[9744]_  = ~\new_[9856]_ ;
  assign \new_[9745]_  = ~\new_[9855]_ ;
  assign \new_[9746]_  = ~\new_[9855]_ ;
  assign \new_[9747]_  = ~\new_[9855]_ ;
  assign \new_[9748]_  = ~\new_[9855]_ ;
  assign \new_[9749]_  = ~\new_[9855]_ ;
  assign \new_[9750]_  = ~\new_[9855]_ ;
  assign \new_[9751]_  = ~\new_[9856]_ ;
  assign \new_[9752]_  = ~\new_[9856]_ ;
  assign \new_[9753]_  = ~\new_[9856]_ ;
  assign \new_[9754]_  = ~\new_[9856]_ ;
  assign \new_[9755]_  = ~\new_[9856]_ ;
  assign \new_[9756]_  = ~\new_[9856]_ ;
  assign \new_[9757]_  = ~\new_[9856]_ ;
  assign \new_[9758]_  = ~\new_[9856]_ ;
  assign n6885 = ~\new_[9900]_  | (~\new_[9565]_  & ~\new_[19875]_ );
  assign \new_[9760]_  = ~\new_[9899]_ ;
  assign \new_[9761]_  = \new_[9901]_  | \new_[15361]_ ;
  assign \new_[9762]_  = ~\new_[20497]_  & ~\new_[9901]_ ;
  assign \new_[9763]_  = ~\new_[9901]_ ;
  assign \new_[9764]_  = ~\\wishbone_slave_unit_del_sync_comp_cycle_count_reg[12] ;
  assign \new_[9765]_  = pci_target_unit_pci_target_if_norm_prf_en_reg;
  assign \new_[9766]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[0] ;
  assign \new_[9767]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[10] ;
  assign \new_[9768]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[11] ;
  assign \new_[9769]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[13] ;
  assign \new_[9770]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[14] ;
  assign \new_[9771]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[15] ;
  assign \new_[9772]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[17] ;
  assign \new_[9773]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[18] ;
  assign \new_[9774]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[1] ;
  assign \new_[9775]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[21] ;
  assign \new_[9776]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[23] ;
  assign \new_[9777]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[25] ;
  assign \new_[9778]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[26] ;
  assign \new_[9779]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[27] ;
  assign \new_[9780]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[29] ;
  assign \new_[9781]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[2] ;
  assign \new_[9782]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[30] ;
  assign \new_[9783]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[32] ;
  assign \new_[9784]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[33] ;
  assign \new_[9785]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[34] ;
  assign \new_[9786]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[3] ;
  assign \new_[9787]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[5] ;
  assign \new_[9788]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[8] ;
  assign \new_[9789]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[7] ;
  assign \new_[9790]_  = \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[0] ;
  assign \new_[9791]_  = ~\\wishbone_slave_unit_del_sync_comp_cycle_count_reg[10] ;
  assign \new_[9792]_  = ~\\wishbone_slave_unit_del_sync_comp_cycle_count_reg[11] ;
  assign \new_[9793]_  = ~\\wishbone_slave_unit_del_sync_comp_cycle_count_reg[14] ;
  assign \new_[9794]_  = \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[1] ;
  assign \new_[9795]_  = \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[3] ;
  assign \new_[9796]_  = \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[5] ;
  assign \new_[9797]_  = ~\\wishbone_slave_unit_del_sync_comp_cycle_count_reg[9] ;
  assign \new_[9798]_  = \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[7] ;
  assign \new_[9799]_  = ~\\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0] ;
  assign \new_[9800]_  = pci_target_unit_pci_target_if_pciw_fifo_wenable_out_reg;
  assign \new_[9801]_  = \\wishbone_slave_unit_fifos_outGreyCount_reg[2] ;
  assign \new_[9802]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[6] ;
  assign \new_[9803]_  = \\wishbone_slave_unit_fifos_outGreyCount_reg[1] ;
  assign \new_[9804]_  = ~\\wishbone_slave_unit_del_sync_bc_out_reg[0] ;
  assign \new_[9805]_  = ~\\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2] ;
  assign \new_[9806]_  = i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg;
  assign \new_[9807]_  = \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[6] ;
  assign \new_[9808]_  = \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[4] ;
  assign \new_[9809]_  = ~\\wishbone_slave_unit_del_sync_comp_cycle_count_reg[13] ;
  assign \new_[9810]_  = \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[2] ;
  assign \new_[9811]_  = ~\\wishbone_slave_unit_del_sync_comp_cycle_count_reg[15] ;
  assign \new_[9812]_  = ~\\wishbone_slave_unit_del_sync_comp_cycle_count_reg[16] ;
  assign \new_[9813]_  = ~\new_[20325]_  | ~\new_[20340]_ ;
  assign \new_[9814]_  = \new_[20325]_  | \new_[16904]_ ;
  assign \new_[9815]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[9] ;
  assign \new_[9816]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[4] ;
  assign \new_[9817]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[35] ;
  assign \new_[9818]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[31] ;
  assign \new_[9819]_  = ~\new_[9881]_ ;
  assign \new_[9820]_  = \new_[9881]_ ;
  assign \new_[9821]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[22] ;
  assign \new_[9822]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[28] ;
  assign \new_[9823]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[24] ;
  assign \new_[9824]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[16] ;
  assign \new_[9825]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[20] ;
  assign \new_[9826]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[12] ;
  assign \new_[9827]_  = ~\\wishbone_slave_unit_wishbone_slave_d_incoming_reg[19] ;
  assign \new_[9828]_  = ~\\wishbone_slave_unit_del_sync_comp_cycle_count_reg[8] ;
  assign \new_[9829]_  = ~\new_[9972]_  & (~\new_[16208]_  | ~\new_[12545]_ );
  assign \new_[9830]_  = ~\new_[20394]_  | ~\new_[16594]_  | ~\new_[11115]_ ;
  assign n6900 = ~\new_[9931]_  | (~\new_[14942]_  & ~\new_[17971]_ );
  assign n7035 = ~\new_[9931]_  | (~\new_[14942]_  & ~\new_[18999]_ );
  assign \new_[9833]_  = \new_[16694]_  ? \new_[10020]_  : \new_[19647]_ ;
  assign \new_[9834]_  = ~\new_[17878]_  | ~wbm_rty_i | ~\new_[19940]_  | ~\new_[10017]_ ;
  assign n6895 = ~\new_[20448]_ ;
  assign \new_[9836]_  = \new_[17017]_  ? \new_[10020]_  : \new_[9488]_ ;
  assign \new_[9837]_  = \new_[19145]_  ? \new_[10020]_  : n17160;
  assign \new_[9838]_  = \new_[18347]_  ? \new_[10020]_  : n17360;
  assign \new_[9839]_  = \new_[19684]_  ? \new_[10020]_  : n17185;
  assign \new_[9840]_  = \new_[17093]_  ? \new_[10020]_  : \new_[19145]_ ;
  assign \new_[9841]_  = \new_[18085]_  ? \new_[10020]_  : \new_[19684]_ ;
  assign \new_[9842]_  = \new_[17244]_  ? \new_[10020]_  : \new_[18347]_ ;
  assign n6905 = ~\new_[9968]_  & (~\new_[15228]_  | ~\new_[17021]_ );
  assign n6910 = ~\new_[9968]_  & (~\new_[15229]_  | ~\new_[16824]_ );
  assign n7030 = ~\new_[9968]_  & (~\new_[15407]_  | ~\new_[16823]_ );
  assign \new_[9846]_  = ~n7270 | ~\new_[17914]_ ;
  assign \new_[9847]_  = n7270 | \new_[17914]_ ;
  assign n6925 = ~\new_[9968]_  & (~\new_[16822]_  | ~\new_[15227]_ );
  assign n7025 = ~\new_[9968]_  & (~\new_[16825]_  | ~\new_[15286]_ );
  assign n6930 = ~\new_[9968]_  & (~\new_[16650]_  | ~\new_[15391]_ );
  assign n6915 = ~\new_[9970]_  | (~\new_[10324]_  & ~\new_[9620]_ );
  assign n6920 = ~\new_[9968]_  & (~\new_[15990]_  | ~\new_[15433]_ );
  assign \new_[9853]_  = ~\new_[9979]_  & ~\new_[18458]_ ;
  assign \new_[9854]_  = ~\new_[9895]_ ;
  assign \new_[9855]_  = \new_[9896]_ ;
  assign \new_[9856]_  = \new_[9896]_ ;
  assign \new_[9857]_  = \new_[9896]_ ;
  assign n6935 = ~\new_[9980]_  | ~\new_[10025]_ ;
  assign n6940 = \new_[16470]_  ? \new_[19875]_  : \new_[9625]_ ;
  assign n6945 = \new_[15944]_  ? \new_[19875]_  : \new_[9626]_ ;
  assign n6950 = \new_[17282]_  ? \new_[19875]_  : \new_[9627]_ ;
  assign n6955 = ~\new_[20449]_ ;
  assign n7020 = ~\new_[20472]_ ;
  assign n6960 = \new_[9635]_  ? \new_[19875]_  : \new_[18031]_ ;
  assign n6965 = \new_[9639]_  ? \new_[19875]_  : \new_[19167]_ ;
  assign n6970 = \new_[9636]_  ? \new_[19875]_  : \new_[19166]_ ;
  assign n7015 = \new_[9637]_  ? \new_[19875]_  : \new_[17989]_ ;
  assign n6975 = \new_[18031]_  ? \new_[19875]_  : n17090;
  assign n6980 = \new_[19167]_  ? \new_[19875]_  : n17025;
  assign n6985 = \new_[19166]_  ? \new_[19875]_  : n17075;
  assign n7005 = \new_[17989]_  ? \new_[19875]_  : n17045;
  assign n6990 = \new_[17414]_  ? \new_[19875]_  : \new_[9635]_ ;
  assign n7010 = \new_[17363]_  ? \new_[19875]_  : \new_[9639]_ ;
  assign n6995 = \new_[17350]_  ? \new_[19875]_  : \new_[9636]_ ;
  assign n7000 = \new_[9641]_  ? \new_[19875]_  : \new_[9637]_ ;
  assign n6835 = ~\new_[9901]_ ;
  assign \new_[9877]_  = pci_target_unit_pci_target_sm_wr_progress_reg;
  assign \new_[9878]_  = pci_target_unit_wishbone_master_w_attempt_reg;
  assign \new_[9879]_  = \\configuration_wb_am2_reg[31] ;
  assign \new_[9880]_  = \\configuration_wb_am1_reg[31] ;
  assign \new_[9881]_  = \new_[18056]_  ? \new_[19974]_  : \new_[19392]_ ;
  assign n7045 = ~\new_[10016]_  | ~\new_[15225]_ ;
  assign n7040 = ~\new_[10013]_  | (~\new_[9671]_  & ~\new_[16572]_ );
  assign \new_[9884]_  = pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg;
  assign \new_[9885]_  = ~\new_[20447]_ ;
  assign \new_[9886]_  = ~\new_[10020]_  | ~\new_[18056]_ ;
  assign \new_[9887]_  = ~\new_[20509]_  | ~\new_[10018]_  | ~\new_[19194]_ ;
  assign \new_[9888]_  = ~\new_[18523]_  | ~\new_[10017]_  | ~\new_[9562]_ ;
  assign n7085 = \new_[18515]_  ? \new_[10324]_  : \new_[16438]_ ;
  assign n7050 = \new_[9673]_  ? \new_[10324]_  : \new_[13794]_ ;
  assign n7055 = \new_[9674]_  ? \new_[10324]_  : \new_[13802]_ ;
  assign n7060 = \new_[9675]_  ? \new_[10324]_  : \new_[13763]_ ;
  assign n7080 = \new_[9679]_  ? \new_[10324]_  : \new_[13809]_ ;
  assign n7065 = \new_[19139]_  ? \new_[10324]_  : \new_[20531]_ ;
  assign \new_[9895]_  = ~\new_[9971]_ ;
  assign \new_[9896]_  = \new_[9971]_ ;
  assign n7070 = ~\new_[10025]_  | (~\new_[9677]_  & ~\new_[10465]_ );
  assign n7075 = ~\new_[20474]_ ;
  assign \new_[9899]_  = ~\new_[9979]_ ;
  assign \new_[9900]_  = ~\new_[9565]_  | ~\new_[19875]_ ;
  assign \new_[9901]_  = ~\new_[9982]_ ;
  assign \new_[9902]_  = \\output_backup_cbe_out_reg[1] ;
  assign \new_[9903]_  = wishbone_slave_unit_pci_initiator_if_del_read_req_reg;
  assign \new_[9904]_  = \\configuration_pci_img_ctrl1_bit2_1_reg[1] ;
  assign \new_[9905]_  = \\configuration_pci_img_ctrl1_bit2_1_reg[2] ;
  assign \new_[9906]_  = \\configuration_wb_ta1_reg[31] ;
  assign \new_[9907]_  = configuration_wb_err_cs_bit0_reg;
  assign \new_[9908]_  = \\configuration_wb_ta2_reg[31] ;
  assign \pci_cbe_o[1]  = pci_io_mux_cbe_iob1_dat_out_reg;
  assign \new_[9910]_  = pci_target_unit_pci_target_sm_master_will_request_read_reg;
  assign n7090 = ~\new_[15009]_  & ~\new_[10315]_ ;
  assign n7390 = ~\new_[15679]_  & ~\new_[10315]_ ;
  assign n7095 = ~\new_[15882]_  | ~\new_[10293]_ ;
  assign n7240 = ~\new_[17092]_  & ~\new_[10315]_ ;
  assign \new_[9915]_  = \new_[10312]_  | \new_[9275]_ ;
  assign n7225 = ~\new_[15427]_  & ~\new_[10315]_ ;
  assign n7255 = ~\new_[15827]_  & ~\new_[10315]_ ;
  assign \new_[9918]_  = ~\new_[10321]_  | ~\new_[16213]_ ;
  assign \new_[9919]_  = ~\new_[19974]_  | ~\new_[18085]_ ;
  assign n7220 = ~\new_[10315]_  & ~\new_[9790]_ ;
  assign n7230 = ~\new_[15395]_  & ~\new_[10315]_ ;
  assign n7315 = ~\new_[15598]_  & ~\new_[10315]_ ;
  assign n7235 = ~\new_[15146]_  & ~\new_[10315]_ ;
  assign n7325 = ~\new_[15113]_  & ~\new_[10315]_ ;
  assign n7320 = ~\new_[16695]_  & ~\new_[10315]_ ;
  assign n7245 = ~\new_[16174]_  & ~\new_[10315]_ ;
  assign n7310 = ~\new_[15896]_  & ~\new_[10315]_ ;
  assign n7250 = ~\new_[16487]_  & ~\new_[10315]_ ;
  assign n7305 = ~\new_[16187]_  & ~\new_[10315]_ ;
  assign n7260 = ~\new_[15913]_  & ~\new_[10315]_ ;
  assign \new_[9931]_  = ~\new_[16706]_  | ~\new_[10320]_  | ~\new_[14942]_ ;
  assign n7100 = \new_[18041]_  ? \new_[20384]_  : \new_[18396]_ ;
  assign n7105 = \new_[19197]_  ? \new_[20384]_  : \new_[18173]_ ;
  assign n7110 = \new_[18063]_  ? \new_[20384]_  : \new_[18033]_ ;
  assign n7380 = \new_[19123]_  ? \new_[20384]_  : \new_[18073]_ ;
  assign n7115 = \new_[17858]_  ? \new_[20384]_  : \new_[18001]_ ;
  assign n7120 = \new_[17894]_  ? \new_[20384]_  : \new_[18586]_ ;
  assign n7125 = \new_[17814]_  ? \new_[20384]_  : \new_[18176]_ ;
  assign n7370 = \new_[18075]_  ? \new_[20384]_  : \new_[18574]_ ;
  assign n7130 = \new_[19038]_  ? \new_[20384]_  : \new_[19322]_ ;
  assign n7135 = \new_[18678]_  ? \new_[20384]_  : \new_[19501]_ ;
  assign n7385 = \new_[19143]_  ? \new_[20384]_  : \new_[17920]_ ;
  assign n7140 = \new_[18102]_  ? \new_[20384]_  : \new_[17887]_ ;
  assign n7375 = \new_[18156]_  ? \new_[20384]_  : \new_[19544]_ ;
  assign n7145 = \new_[18099]_  ? \new_[20384]_  : \new_[18049]_ ;
  assign n7355 = \new_[18035]_  ? \new_[20384]_  : \new_[18310]_ ;
  assign n7150 = \new_[18227]_  ? \new_[20384]_  : \new_[19616]_ ;
  assign n7365 = \new_[18839]_  ? \new_[20384]_  : \new_[18852]_ ;
  assign n7155 = \new_[19250]_  ? \new_[20384]_  : \new_[18389]_ ;
  assign n7160 = \new_[18628]_  ? \new_[20384]_  : \new_[18770]_ ;
  assign n7165 = \new_[17824]_  ? \new_[20384]_  : \new_[18187]_ ;
  assign n7360 = \new_[17884]_  ? \new_[20384]_  : \new_[18560]_ ;
  assign n7170 = \new_[17860]_  ? \new_[20384]_  : \new_[19333]_ ;
  assign n7175 = \new_[18441]_  ? \new_[20384]_  : \new_[19711]_ ;
  assign n7180 = \new_[18406]_  ? \new_[20384]_  : \new_[19674]_ ;
  assign n7350 = \new_[18290]_  ? \new_[20384]_  : \new_[19389]_ ;
  assign n7185 = \new_[18589]_  ? \new_[20384]_  : \new_[13794]_ ;
  assign n7190 = \new_[18288]_  ? \new_[20384]_  : \new_[13802]_ ;
  assign n7195 = \new_[18596]_  ? \new_[20384]_  : \new_[13763]_ ;
  assign n7345 = \new_[18594]_  ? \new_[20384]_  : \new_[13809]_ ;
  assign n7200 = \new_[18520]_  ? \new_[20384]_  : \new_[19738]_ ;
  assign n7340 = \new_[18843]_  ? \new_[20384]_  : \new_[18897]_ ;
  assign n7205 = \new_[18277]_  ? \new_[20384]_  : \new_[18555]_ ;
  assign n7280 = \new_[19069]_  ? \new_[20384]_  : \new_[18149]_ ;
  assign n7215 = \new_[18733]_  ? \new_[20384]_  : \new_[19720]_ ;
  assign n7210 = \new_[18814]_  ? \new_[20384]_  : \new_[17822]_ ;
  assign n7335 = \new_[18260]_  ? \new_[20384]_  : \new_[19835]_ ;
  assign \new_[9968]_  = ~\new_[10017]_ ;
  assign n7290 = ~\new_[10324]_  & ~\new_[9804]_ ;
  assign \new_[9970]_  = ~\new_[10018]_ ;
  assign \new_[9971]_  = ~\new_[10022]_ ;
  assign \new_[9972]_  = \new_[15812]_  | \new_[10332]_ ;
  assign n7270 = ~\new_[10023]_ ;
  assign n7295 = \new_[19224]_  ? \new_[10465]_  : \new_[16225]_ ;
  assign n7285 = \new_[9803]_  ? \new_[10465]_  : \new_[17005]_ ;
  assign n7265 = \new_[18199]_  ^ \new_[10465]_ ;
  assign n7275 = \new_[9801]_  ? \new_[10465]_  : \new_[19224]_ ;
  assign n7300 = \new_[10459]_  ? wbs_rty_o : \new_[19918]_ ;
  assign \new_[9979]_  = ~wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg;
  assign \new_[9980]_  = ~\new_[10329]_  | ~\new_[9624]_ ;
  assign n7330 = ~\new_[13709]_  & ~\new_[10315]_ ;
  assign \new_[9982]_  = ~\new_[20406]_ ;
  assign \new_[9983]_  = ~output_backup_par_out_reg;
  assign pci_par_o = pci_io_mux_par_iob_dat_out_reg;
  assign \new_[9985]_  = configuration_pci_err_cs_bit0_reg;
  assign \new_[9986]_  = \\configuration_wb_img_ctrl1_bit2_0_reg[2] ;
  assign \new_[9987]_  = \\configuration_interrupt_line_reg[6] ;
  assign \new_[9988]_  = \\configuration_wb_img_ctrl2_bit2_0_reg[1] ;
  assign \new_[9989]_  = \\configuration_interrupt_line_reg[2] ;
  assign n16740 = wishbone_slave_unit_del_sync_req_req_pending_reg;
  assign \new_[9991]_  = \\configuration_wb_img_ctrl1_bit2_0_reg[0] ;
  assign \new_[9992]_  = \\configuration_wb_img_ctrl1_bit2_0_reg[1] ;
  assign \new_[9993]_  = \\configuration_interrupt_line_reg[0] ;
  assign \new_[9994]_  = \\configuration_interrupt_line_reg[1] ;
  assign \new_[9995]_  = \\configuration_wb_img_ctrl2_bit2_0_reg[0] ;
  assign \new_[9996]_  = \\configuration_wb_img_ctrl2_bit2_0_reg[2] ;
  assign \new_[9997]_  = \\configuration_command_bit2_0_reg[0] ;
  assign \new_[9998]_  = \\configuration_command_bit2_0_reg[1] ;
  assign n17430 = \\configuration_command_bit2_0_reg[2] ;
  assign \new_[10000]_  = configuration_wb_ba1_bit0_reg;
  assign \new_[10001]_  = configuration_wb_ba2_bit0_reg;
  assign \new_[10002]_  = configuration_command_bit8_reg;
  assign \new_[10003]_  = configuration_wb_err_cs_bit8_reg;
  assign \new_[10004]_  = \\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1] ;
  assign \new_[10005]_  = \\configuration_status_bit15_11_reg[11] ;
  assign \new_[10006]_  = \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1] ;
  assign \new_[10007]_  = \\configuration_status_bit15_11_reg[12] ;
  assign \new_[10008]_  = \\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0] ;
  assign \new_[10009]_  = \\configuration_status_bit15_11_reg[13] ;
  assign \new_[10010]_  = \\configuration_isr_bit2_0_reg[1] ;
  assign \new_[10011]_  = ~wishbone_slave_unit_del_sync_comp_comp_pending_reg;
  assign \new_[10012]_  = \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[0] ;
  assign \new_[10013]_  = ~\new_[17254]_  | ~\new_[15879]_  | ~\new_[10825]_ ;
  assign n7415 = ~\new_[15881]_  | ~\new_[10449]_ ;
  assign n7395 = ~\new_[15002]_  | ~\new_[10449]_  | ~\new_[15869]_ ;
  assign \new_[10016]_  = \new_[16363]_  & \new_[10450]_ ;
  assign \new_[10017]_  = ~pci_target_unit_wishbone_master_reset_rty_cnt_reg;
  assign \new_[10018]_  = ~\new_[10453]_  & ~\new_[10497]_ ;
  assign \new_[10019]_  = ~\new_[10453]_  | ~\new_[9282]_ ;
  assign \new_[10020]_  = \new_[19974]_ ;
  assign \new_[10021]_  = ~\new_[17354]_  & ~\new_[10453]_ ;
  assign \new_[10022]_  = ~\new_[10456]_  | ~\new_[16227]_ ;
  assign \new_[10023]_  = ~\new_[10321]_ ;
  assign n7400 = ~\new_[10455]_  | (~\new_[20517]_  & ~\new_[15841]_ );
  assign \new_[10025]_  = ~\new_[17004]_  | ~\new_[10465]_ ;
  assign \new_[10026]_  = ~\new_[16637]_  | (~\new_[17003]_  & ~\new_[10830]_ );
  assign \new_[10027]_  = ~\new_[16375]_  | (~\new_[16662]_  & ~\new_[10830]_ );
  assign \new_[10028]_  = ~\new_[16380]_  | (~\new_[16804]_  & ~\new_[10830]_ );
  assign \new_[10029]_  = ~\new_[16365]_  | (~\new_[16790]_  & ~\new_[10830]_ );
  assign \new_[10030]_  = ~\new_[16592]_  | (~\new_[16896]_  & ~\new_[10830]_ );
  assign \new_[10031]_  = ~\new_[16590]_  | (~\new_[17001]_  & ~\new_[10830]_ );
  assign \new_[10032]_  = ~\new_[16371]_  | (~\new_[16679]_  & ~\new_[10830]_ );
  assign \new_[10033]_  = ~\new_[16366]_  | (~\new_[16805]_  & ~\new_[10830]_ );
  assign \new_[10034]_  = ~\new_[16841]_  | (~\new_[17131]_  & ~\new_[10830]_ );
  assign \new_[10035]_  = ~\new_[16364]_  | (~\new_[16796]_  & ~\new_[10830]_ );
  assign \new_[10036]_  = ~\new_[16373]_  | (~\new_[16797]_  & ~\new_[10830]_ );
  assign \new_[10037]_  = ~\new_[10464]_  | (~\new_[8401]_  & ~\new_[16911]_ );
  assign \new_[10038]_  = ~\new_[10460]_  | (~\new_[8696]_  & ~\new_[16975]_ );
  assign \new_[10039]_  = ~\new_[10461]_  | (~\new_[9198]_  & ~\new_[16976]_ );
  assign \new_[10040]_  = ~\new_[10462]_  | (~\new_[9199]_  & ~\new_[16900]_ );
  assign \new_[10041]_  = ~\new_[10463]_  | (~\new_[9229]_  & ~\new_[17191]_ );
  assign \new_[10042]_  = \\configuration_wb_ba2_bit31_12_reg[31] ;
  assign \new_[10043]_  = \\configuration_wb_ba1_bit31_12_reg[31] ;
  assign n7410 = ~\new_[10414]_  | (~\new_[11123]_  & ~\new_[16418]_ );
  assign n7405 = ~\new_[10415]_  | (~\new_[11124]_  & ~\new_[16418]_ );
  assign \new_[10046]_  = configuration_command_bit6_reg;
  assign \new_[10047]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][1] ;
  assign \new_[10048]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][6] ;
  assign \new_[10049]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][3] ;
  assign \new_[10050]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[1] ;
  assign \new_[10051]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][26] ;
  assign \new_[10052]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][31] ;
  assign \new_[10053]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][2] ;
  assign \new_[10054]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][22] ;
  assign \new_[10055]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][24] ;
  assign \new_[10056]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][19] ;
  assign \new_[10057]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][20] ;
  assign \new_[10058]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][11] ;
  assign \new_[10059]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][0] ;
  assign \new_[10060]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][8] ;
  assign \new_[10061]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][15] ;
  assign \new_[10062]_  = \\configuration_icr_bit2_0_reg[0] ;
  assign \new_[10063]_  = \\configuration_icr_bit2_0_reg[1] ;
  assign \new_[10064]_  = \\configuration_icr_bit2_0_reg[2] ;
  assign \new_[10065]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][4] ;
  assign \new_[10066]_  = \\configuration_interrupt_line_reg[3] ;
  assign n16995 = \\configuration_cache_line_size_reg_reg[3] ;
  assign \new_[10068]_  = \\configuration_interrupt_line_reg[5] ;
  assign \new_[10069]_  = \\configuration_interrupt_line_reg[4] ;
  assign n17500 = \\configuration_cache_line_size_reg_reg[5] ;
  assign n17350 = \\configuration_cache_line_size_reg_reg[4] ;
  assign \new_[10072]_  = ~configuration_sync_isr_2_del_bit_reg;
  assign \new_[10073]_  = ~configuration_sync_pci_err_cs_8_del_bit_reg;
  assign \new_[10074]_  = \\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2] ;
  assign \new_[10075]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[0] ;
  assign \new_[10076]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[2] ;
  assign \new_[10077]_  = \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2] ;
  assign \new_[10078]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][0] ;
  assign \new_[10079]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][10] ;
  assign \new_[10080]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][12] ;
  assign \new_[10081]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][14] ;
  assign \new_[10082]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][16] ;
  assign \new_[10083]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][18] ;
  assign \new_[10084]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][1] ;
  assign \new_[10085]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][20] ;
  assign \new_[10086]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][21] ;
  assign \new_[10087]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][23] ;
  assign \new_[10088]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][25] ;
  assign \new_[10089]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][27] ;
  assign \new_[10090]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][29] ;
  assign \new_[10091]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][30] ;
  assign \new_[10092]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][37] ;
  assign \new_[10093]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][4] ;
  assign \new_[10094]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][5] ;
  assign \new_[10095]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][6] ;
  assign \new_[10096]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][8] ;
  assign \new_[10097]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][0] ;
  assign \new_[10098]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][11] ;
  assign \new_[10099]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][12] ;
  assign \new_[10100]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][13] ;
  assign \new_[10101]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][15] ;
  assign \new_[10102]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][16] ;
  assign \new_[10103]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][17] ;
  assign \new_[10104]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][19] ;
  assign \new_[10105]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][1] ;
  assign \new_[10106]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][20] ;
  assign \new_[10107]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][22] ;
  assign \new_[10108]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][24] ;
  assign \new_[10109]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][26] ;
  assign \new_[10110]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][28] ;
  assign \new_[10111]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][2] ;
  assign \new_[10112]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][31] ;
  assign \new_[10113]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][3] ;
  assign \new_[10114]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][4] ;
  assign \new_[10115]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][5] ;
  assign \new_[10116]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][7] ;
  assign \new_[10117]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][8] ;
  assign \new_[10118]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][9] ;
  assign \new_[10119]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][10] ;
  assign \new_[10120]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][11] ;
  assign \new_[10121]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][12] ;
  assign \new_[10122]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][14] ;
  assign \new_[10123]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][16] ;
  assign \new_[10124]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][18] ;
  assign \new_[10125]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][19] ;
  assign \new_[10126]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][1] ;
  assign \new_[10127]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][21] ;
  assign \new_[10128]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][23] ;
  assign \new_[10129]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][25] ;
  assign \new_[10130]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][26] ;
  assign \new_[10131]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][27] ;
  assign \new_[10132]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][29] ;
  assign \new_[10133]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][30] ;
  assign \new_[10134]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][37] ;
  assign \new_[10135]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][3] ;
  assign \new_[10136]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][4] ;
  assign \new_[10137]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][6] ;
  assign \new_[10138]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][7] ;
  assign \new_[10139]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][8] ;
  assign \new_[10140]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][0] ;
  assign \new_[10141]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][10] ;
  assign \new_[10142]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][11] ;
  assign \new_[10143]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][13] ;
  assign \new_[10144]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][15] ;
  assign \new_[10145]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][17] ;
  assign \new_[10146]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][18] ;
  assign \new_[10147]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][19] ;
  assign \new_[10148]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][20] ;
  assign \new_[10149]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][22] ;
  assign \new_[10150]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][24] ;
  assign \new_[10151]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][25] ;
  assign \new_[10152]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][26] ;
  assign \new_[10153]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][28] ;
  assign \new_[10154]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][29] ;
  assign \new_[10155]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][2] ;
  assign \new_[10156]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][31] ;
  assign \new_[10157]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][37] ;
  assign \new_[10158]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][3] ;
  assign \new_[10159]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][5] ;
  assign \new_[10160]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][7] ;
  assign \new_[10161]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][9] ;
  assign \new_[10162]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][14] ;
  assign \new_[10163]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][15] ;
  assign \new_[10164]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][16] ;
  assign \new_[10165]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][18] ;
  assign \new_[10166]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][1] ;
  assign \new_[10167]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][21] ;
  assign \new_[10168]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][22] ;
  assign \new_[10169]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][23] ;
  assign \new_[10170]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][25] ;
  assign \new_[10171]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][27] ;
  assign \new_[10172]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][29] ;
  assign \new_[10173]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][2] ;
  assign \new_[10174]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][30] ;
  assign \new_[10175]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][37] ;
  assign \new_[10176]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][4] ;
  assign \new_[10177]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][6] ;
  assign \new_[10178]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][7] ;
  assign \new_[10179]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][8] ;
  assign \new_[10180]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][0] ;
  assign \new_[10181]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][11] ;
  assign \new_[10182]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][13] ;
  assign \new_[10183]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][14] ;
  assign \new_[10184]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][15] ;
  assign \new_[10185]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][17] ;
  assign \new_[10186]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][18] ;
  assign \new_[10187]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][19] ;
  assign \new_[10188]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][20] ;
  assign \new_[10189]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][22] ;
  assign \new_[10190]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][24] ;
  assign \new_[10191]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][26] ;
  assign \new_[10192]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][28] ;
  assign \new_[10193]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][29] ;
  assign \new_[10194]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][2] ;
  assign \new_[10195]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][31] ;
  assign \new_[10196]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][3] ;
  assign \new_[10197]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][5] ;
  assign \new_[10198]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][7] ;
  assign \new_[10199]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][9] ;
  assign \new_[10200]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][10] ;
  assign \new_[10201]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][12] ;
  assign \new_[10202]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][13] ;
  assign \new_[10203]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][14] ;
  assign \new_[10204]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][16] ;
  assign \new_[10205]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][17] ;
  assign \new_[10206]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][18] ;
  assign \new_[10207]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][1] ;
  assign \new_[10208]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][21] ;
  assign \new_[10209]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][23] ;
  assign \new_[10210]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][25] ;
  assign \new_[10211]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][27] ;
  assign \new_[10212]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][28] ;
  assign \new_[10213]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][29] ;
  assign \new_[10214]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][30] ;
  assign \new_[10215]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][37] ;
  assign \new_[10216]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][4] ;
  assign \new_[10217]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][5] ;
  assign \new_[10218]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][6] ;
  assign \new_[10219]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][8] ;
  assign \new_[10220]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][9] ;
  assign \new_[10221]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][0] ;
  assign \new_[10222]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][11] ;
  assign \new_[10223]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][13] ;
  assign \new_[10224]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][15] ;
  assign \new_[10225]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][17] ;
  assign \new_[10226]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][19] ;
  assign \new_[10227]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][1] ;
  assign \new_[10228]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][20] ;
  assign \new_[10229]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][22] ;
  assign \new_[10230]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][24] ;
  assign \new_[10231]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][26] ;
  assign \new_[10232]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][27] ;
  assign \new_[10233]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][28] ;
  assign \new_[10234]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][2] ;
  assign \new_[10235]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][31] ;
  assign \new_[10236]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][3] ;
  assign \new_[10237]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][4] ;
  assign \new_[10238]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][5] ;
  assign \new_[10239]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][7] ;
  assign \new_[10240]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][9] ;
  assign \new_[10241]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][10] ;
  assign \new_[10242]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][12] ;
  assign \new_[10243]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][30] ;
  assign \new_[10244]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][37] ;
  assign \new_[10245]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][25] ;
  assign \new_[10246]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][27] ;
  assign \new_[10247]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][23] ;
  assign n7475 = \new_[12358]_  ? \new_[11095]_  : \new_[10937]_ ;
  assign \new_[10249]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][21] ;
  assign \new_[10250]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][1] ;
  assign \new_[10251]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][16] ;
  assign \new_[10252]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][9] ;
  assign \new_[10253]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][10] ;
  assign \new_[10254]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][12] ;
  assign \new_[10255]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][26] ;
  assign \new_[10256]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][21] ;
  assign n17335 = \\configuration_cache_line_size_reg_reg[7] ;
  assign \new_[10258]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][3] ;
  assign \new_[10259]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][5] ;
  assign \new_[10260]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][31] ;
  assign \new_[10261]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][28] ;
  assign \new_[10262]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][24] ;
  assign \new_[10263]_  = \\configuration_interrupt_line_reg[7] ;
  assign \new_[10264]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][19] ;
  assign \new_[10265]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][20] ;
  assign \new_[10266]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][17] ;
  assign \new_[10267]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][4] ;
  assign \new_[10268]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][8] ;
  assign \new_[10269]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][6] ;
  assign \new_[10270]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][30] ;
  assign \new_[10271]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][27] ;
  assign \new_[10272]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][23] ;
  assign \new_[10273]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][8] ;
  assign \new_[10274]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][9] ;
  assign \new_[10275]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][28] ;
  assign \new_[10276]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][14] ;
  assign \new_[10277]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][16] ;
  assign \new_[10278]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][12] ;
  assign \new_[10279]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][5] ;
  assign \new_[10280]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][2] ;
  assign \new_[10281]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][31] ;
  assign \new_[10282]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][24] ;
  assign \new_[10283]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][22] ;
  assign \new_[10284]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][0] ;
  assign \new_[10285]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][0] ;
  assign \new_[10286]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][20] ;
  assign \new_[10287]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][11] ;
  assign \new_[10288]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][13] ;
  assign \new_[10289]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][17] ;
  assign \new_[10290]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][13] ;
  assign \new_[10291]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][15] ;
  assign \new_[10292]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][29] ;
  assign \new_[10293]_  = ~\new_[16572]_  | ~\new_[10825]_  | ~\new_[9904]_ ;
  assign \new_[10294]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][6] ;
  assign \new_[10295]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][6] ;
  assign \new_[10296]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][37] ;
  assign \new_[10297]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][21] ;
  assign \new_[10298]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][30] ;
  assign \new_[10299]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][29] ;
  assign \new_[10300]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][30] ;
  assign \new_[10301]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][37] ;
  assign \new_[10302]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][25] ;
  assign \new_[10303]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][23] ;
  assign \new_[10304]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][25] ;
  assign \new_[10305]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][10] ;
  assign \new_[10306]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][18] ;
  assign \new_[10307]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][27] ;
  assign \new_[10308]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][16] ;
  assign \new_[10309]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][18] ;
  assign \new_[10310]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][23] ;
  assign \new_[10311]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][12] ;
  assign \new_[10312]_  = ~\new_[19975]_ ;
  assign \new_[10313]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][14] ;
  assign n7425 = ~\new_[10948]_  | ~\new_[13823]_  | ~\new_[15277]_ ;
  assign \new_[10315]_  = ~\new_[19933]_  | ~\new_[16802]_  | ~\new_[20443]_ ;
  assign \new_[10316]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][21] ;
  assign \new_[10317]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][14] ;
  assign \new_[10318]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][10] ;
  assign \new_[10319]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][9] ;
  assign \new_[10320]_  = ~\new_[11145]_  | ~\new_[19742]_  | ~\new_[19360]_  | ~\new_[15632]_ ;
  assign \new_[10321]_  = ~\new_[10826]_  | ~\new_[13126]_ ;
  assign n7420 = \new_[10958]_  ? \new_[12484]_  : \new_[9902]_ ;
  assign n7455 = \pci_cbe_o[1]  ? \new_[15613]_  : \new_[10958]_ ;
  assign \new_[10324]_  = ~\new_[10453]_ ;
  assign \new_[10325]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][7] ;
  assign n7460 = ~\new_[10458]_ ;
  assign \new_[10327]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][7] ;
  assign \new_[10328]_  = ~\new_[10459]_ ;
  assign \new_[10329]_  = ~\new_[10465]_ ;
  assign n7465 = ~\new_[10835]_  | (~\new_[16687]_  & ~\new_[20398]_ );
  assign \new_[10331]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][28] ;
  assign \new_[10332]_  = ~\new_[16791]_  & (~\new_[12469]_  | ~\new_[10935]_ );
  assign n7430 = ~\new_[10836]_  | (~\new_[12238]_  & ~\new_[15934]_ );
  assign n7435 = ~\new_[10837]_  | (~\new_[12238]_  & ~\new_[16122]_ );
  assign \new_[10335]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][2] ;
  assign \new_[10336]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][3] ;
  assign \new_[10337]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][31] ;
  assign \new_[10338]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][26] ;
  assign \new_[10339]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][22] ;
  assign \new_[10340]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][24] ;
  assign \new_[10341]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][13] ;
  assign \new_[10342]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][19] ;
  assign \new_[10343]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][17] ;
  assign \new_[10344]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][15] ;
  assign n7440 = ~\new_[10531]_  | (~\new_[11667]_  & ~\new_[16418]_ );
  assign n7480 = ~\new_[10533]_  | (~\new_[11669]_  & ~\new_[15899]_ );
  assign n7445 = ~\new_[10535]_  | (~\new_[11671]_  & ~\new_[15899]_ );
  assign n7450 = ~\new_[10532]_  | (~\new_[16418]_  & ~\new_[11672]_ );
  assign \new_[10349]_  = ~\\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][11] ;
  assign \new_[10350]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[5] ;
  assign \new_[10351]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[7] ;
  assign \new_[10352]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[8] ;
  assign \new_[10353]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[23] ;
  assign \new_[10354]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[4] ;
  assign \new_[10355]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[31] ;
  assign \new_[10356]_  = \\configuration_pci_ba0_bit31_8_reg[12] ;
  assign \new_[10357]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[27] ;
  assign \new_[10358]_  = \\configuration_latency_timer_reg[1] ;
  assign \new_[10359]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[12] ;
  assign \new_[10360]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[1] ;
  assign \new_[10361]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[21] ;
  assign \new_[10362]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[14] ;
  assign \new_[10363]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[16] ;
  assign \new_[10364]_  = \\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1] ;
  assign \new_[10365]_  = configuration_icr_bit31_reg;
  assign \new_[10366]_  = wishbone_slave_unit_wishbone_slave_img_wallow_reg;
  assign \new_[10367]_  = wishbone_slave_unit_wishbone_slave_do_del_request_reg;
  assign \new_[10368]_  = ~wishbone_slave_unit_wishbone_slave_mrl_en_reg;
  assign \new_[10369]_  = ~wishbone_slave_unit_wishbone_slave_pref_en_reg;
  assign \new_[10370]_  = wishbone_slave_unit_wishbone_slave_del_addr_hit_reg;
  assign \new_[10371]_  = \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[1] ;
  assign \new_[10372]_  = wishbone_slave_unit_wishbone_slave_del_completion_allow_reg;
  assign n16895 = pci_target_unit_del_sync_comp_comp_pending_reg;
  assign \new_[10374]_  = pci_target_unit_del_sync_comp_req_pending_reg;
  assign \new_[10375]_  = \\pci_target_unit_wishbone_master_c_state_reg[2] ;
  assign \new_[10376]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][37] ;
  assign \new_[10377]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][37] ;
  assign \new_[10378]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][37] ;
  assign \new_[10379]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][37] ;
  assign \new_[10380]_  = wishbone_slave_unit_pci_initiator_if_intermediate_last_reg;
  assign \new_[10381]_  = ~\\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[1] ;
  assign \new_[10382]_  = \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1] ;
  assign \new_[10383]_  = \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0] ;
  assign \new_[10384]_  = \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2] ;
  assign \new_[10385]_  = \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3] ;
  assign \new_[10386]_  = \\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0] ;
  assign \new_[10387]_  = \\configuration_latency_timer_reg[0] ;
  assign \new_[10388]_  = \\configuration_latency_timer_reg[2] ;
  assign \new_[10389]_  = \\configuration_latency_timer_reg[3] ;
  assign \new_[10390]_  = \\configuration_latency_timer_reg[4] ;
  assign \new_[10391]_  = \\configuration_latency_timer_reg[5] ;
  assign \new_[10392]_  = \\configuration_latency_timer_reg[6] ;
  assign \new_[10393]_  = \\configuration_latency_timer_reg[7] ;
  assign \new_[10394]_  = \\configuration_cache_line_size_reg_reg[0] ;
  assign \new_[10395]_  = \\configuration_pci_ba0_bit31_8_reg[14] ;
  assign \new_[10396]_  = \\configuration_cache_line_size_reg_reg[1] ;
  assign n17220 = \\configuration_cache_line_size_reg_reg[2] ;
  assign \new_[10398]_  = \\configuration_pci_ba0_bit31_8_reg[13] ;
  assign \new_[10399]_  = \\configuration_pci_ba0_bit31_8_reg[17] ;
  assign n17280 = \\configuration_cache_line_size_reg_reg[6] ;
  assign \new_[10401]_  = \\configuration_pci_ba0_bit31_8_reg[16] ;
  assign \new_[10402]_  = \\configuration_pci_ba0_bit31_8_reg[20] ;
  assign \new_[10403]_  = \\configuration_pci_ba0_bit31_8_reg[23] ;
  assign \new_[10404]_  = \\configuration_pci_ba0_bit31_8_reg[18] ;
  assign \new_[10405]_  = \\configuration_pci_ba0_bit31_8_reg[15] ;
  assign \new_[10406]_  = \\configuration_pci_ba0_bit31_8_reg[19] ;
  assign \new_[10407]_  = \\configuration_pci_ba0_bit31_8_reg[25] ;
  assign \new_[10408]_  = \\configuration_pci_ba0_bit31_8_reg[27] ;
  assign \new_[10409]_  = \\configuration_pci_ba0_bit31_8_reg[28] ;
  assign \new_[10410]_  = \\configuration_pci_ba0_bit31_8_reg[30] ;
  assign \new_[10411]_  = \\configuration_pci_ba0_bit31_8_reg[29] ;
  assign \new_[10412]_  = \\pci_target_unit_wishbone_master_read_count_reg[1] ;
  assign \new_[10413]_  = ~\\pci_target_unit_wishbone_master_read_count_reg[2] ;
  assign \new_[10414]_  = ~\new_[9880]_  | (~\new_[11123]_  & ~\new_[17476]_ );
  assign \new_[10415]_  = ~\new_[9879]_  | (~\new_[11124]_  & ~\new_[17476]_ );
  assign \new_[10416]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[0] ;
  assign \new_[10417]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[10] ;
  assign \new_[10418]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[11] ;
  assign \new_[10419]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[13] ;
  assign \new_[10420]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[15] ;
  assign \new_[10421]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[17] ;
  assign \new_[10422]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[18] ;
  assign \new_[10423]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[19] ;
  assign \new_[10424]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[20] ;
  assign \new_[10425]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[22] ;
  assign \new_[10426]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[24] ;
  assign \new_[10427]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[25] ;
  assign \new_[10428]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[26] ;
  assign \new_[10429]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[28] ;
  assign \new_[10430]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[29] ;
  assign \new_[10431]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[2] ;
  assign \new_[10432]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[3] ;
  assign \new_[10433]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[6] ;
  assign \new_[10434]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[9] ;
  assign \new_[10435]_  = \\wishbone_slave_unit_pci_initiator_if_data_out_reg[30] ;
  assign n7570 = ~\new_[10921]_  | (~\new_[14242]_  & ~\new_[19466]_ );
  assign n7590 = ~\new_[10928]_  | ~\new_[15252]_ ;
  assign n7605 = ~\new_[10922]_  | (~\new_[17578]_  & ~\new_[14242]_ );
  assign n7600 = ~\new_[10926]_  | ~\new_[16103]_ ;
  assign n7575 = ~\new_[10931]_  | ~\new_[11104]_ ;
  assign n7615 = ~\new_[10932]_  | ~\new_[11104]_ ;
  assign n7585 = ~\new_[10930]_  | (~\new_[16408]_  & ~\new_[11675]_ );
  assign n7595 = ~\new_[10929]_  | (~\new_[11675]_  & ~\new_[17656]_ );
  assign \new_[10444]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][37] ;
  assign \new_[10445]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][37] ;
  assign \new_[10446]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][37] ;
  assign \new_[10447]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][37] ;
  assign \new_[10448]_  = ~wishbone_slave_unit_del_sync_comp_req_pending_reg;
  assign \new_[10449]_  = ~\new_[20332]_  | ~\new_[16572]_ ;
  assign \new_[10450]_  = ~\new_[16572]_  | ~\new_[20332]_  | ~\new_[17254]_ ;
  assign n7610 = ~\new_[10942]_  & (~\new_[17743]_  | ~n17480);
  assign n7505 = ~\new_[15500]_  & (~\new_[11138]_  | ~\new_[19012]_ );
  assign \new_[10453]_  = ~\new_[19012]_  | ~\new_[10954]_  | ~\new_[17308]_ ;
  assign n7620 = ~\new_[17029]_  | ~\new_[10949]_ ;
  assign \new_[10455]_  = ~\new_[10949]_  | ~\new_[17752]_ ;
  assign \new_[10456]_  = ~\new_[20388]_  | ~\new_[20389]_  | ~\new_[11150]_ ;
  assign \new_[10457]_  = ~\new_[14966]_  | ~\new_[10961]_  | ~\new_[15315]_ ;
  assign \new_[10458]_  = ~\new_[19201]_  | ~\new_[17843]_  | ~\new_[11016]_  | ~\new_[15908]_ ;
  assign \new_[10459]_  = ~\new_[12482]_  | ~\new_[11018]_ ;
  assign \new_[10460]_  = ~\new_[16975]_  | ~\new_[10974]_ ;
  assign \new_[10461]_  = ~\new_[16976]_  | ~\new_[10974]_ ;
  assign \new_[10462]_  = ~\new_[16900]_  | ~\new_[10974]_ ;
  assign \new_[10463]_  = ~\new_[17191]_  | ~\new_[10974]_ ;
  assign \new_[10464]_  = ~\new_[16911]_  | ~\new_[10974]_ ;
  assign \new_[10465]_  = \new_[20185]_  & \new_[19308]_ ;
  assign n7510 = ~\new_[11026]_  | (~\new_[12576]_  & ~\new_[15899]_ );
  assign n7485 = ~\new_[11028]_  | (~\new_[12576]_  & ~\new_[16122]_ );
  assign n7515 = ~\new_[11027]_  | (~\new_[12576]_  & ~\new_[15934]_ );
  assign n7580 = ~\new_[10925]_  | ~\new_[16406]_ ;
  assign n7555 = ~\new_[10872]_  | (~\new_[12290]_  & ~\new_[15899]_ );
  assign n7630 = ~\new_[10871]_  | (~\new_[12290]_  & ~\new_[16418]_ );
  assign n7560 = ~\new_[10873]_  | (~\new_[12289]_  & ~\new_[15899]_ );
  assign n7625 = ~\new_[10874]_  | (~\new_[12289]_  & ~\new_[16418]_ );
  assign n7565 = ~\new_[10875]_  | (~\new_[12295]_  & ~\new_[16677]_ );
  assign n7520 = ~\new_[10838]_ ;
  assign n7525 = ~\new_[10839]_ ;
  assign n7500 = ~\new_[10840]_ ;
  assign n7530 = ~\new_[10841]_ ;
  assign n7495 = ~\new_[10842]_ ;
  assign n7535 = ~\new_[10843]_ ;
  assign \new_[10481]_  = \\configuration_pci_ba0_bit31_8_reg[31] ;
  assign n7490 = ~\new_[10844]_ ;
  assign \new_[10483]_  = \\configuration_pci_ba0_bit31_8_reg[26] ;
  assign \new_[10484]_  = \\configuration_pci_ba0_bit31_8_reg[24] ;
  assign \new_[10485]_  = \\configuration_pci_ba0_bit31_8_reg[21] ;
  assign \new_[10486]_  = \\configuration_pci_ba0_bit31_8_reg[22] ;
  assign n7540 = ~\new_[10849]_ ;
  assign n7545 = ~\new_[10850]_ ;
  assign n7550 = ~\new_[10851]_ ;
  assign n7635 = ~\new_[10852]_ ;
  assign \new_[10491]_  = \\configuration_pci_am1_reg[16] ;
  assign \new_[10492]_  = \\configuration_pci_am1_reg[15] ;
  assign \new_[10493]_  = \\configuration_pci_am1_reg[24] ;
  assign \new_[10494]_  = \\configuration_pci_ba1_bit31_8_reg[11] ;
  assign \new_[10495]_  = \\configuration_pci_ba1_bit31_8_reg[15] ;
  assign \new_[10496]_  = ~\\wishbone_slave_unit_pci_initiator_if_read_count_reg[3] ;
  assign \new_[10497]_  = wishbone_slave_unit_wishbone_slave_map_reg;
  assign \new_[10498]_  = \\configuration_pci_ba1_bit31_8_reg[18] ;
  assign \new_[10499]_  = \\configuration_pci_ba1_bit31_8_reg[19] ;
  assign \new_[10500]_  = \\configuration_pci_ba1_bit31_8_reg[20] ;
  assign \new_[10501]_  = \\configuration_pci_ba1_bit31_8_reg[21] ;
  assign \new_[10502]_  = \\configuration_pci_ba1_bit31_8_reg[23] ;
  assign \new_[10503]_  = \\configuration_pci_ba1_bit31_8_reg[25] ;
  assign \new_[10504]_  = \\configuration_pci_ba1_bit31_8_reg[26] ;
  assign \new_[10505]_  = \\configuration_pci_ba1_bit31_8_reg[27] ;
  assign \new_[10506]_  = \\configuration_pci_ba1_bit31_8_reg[29] ;
  assign \new_[10507]_  = \\configuration_pci_ba1_bit31_8_reg[30] ;
  assign \new_[10508]_  = \\configuration_pci_ba1_bit31_8_reg[10] ;
  assign \new_[10509]_  = \\configuration_pci_ba1_bit31_8_reg[12] ;
  assign \new_[10510]_  = \\configuration_pci_ba1_bit31_8_reg[13] ;
  assign \new_[10511]_  = \\configuration_pci_ba1_bit31_8_reg[14] ;
  assign \new_[10512]_  = \\configuration_pci_ba1_bit31_8_reg[16] ;
  assign \new_[10513]_  = \\pci_target_unit_wishbone_master_c_state_reg[1] ;
  assign \new_[10514]_  = \\configuration_pci_am1_reg[21] ;
  assign \new_[10515]_  = \\configuration_pci_am1_reg[10] ;
  assign \new_[10516]_  = \\configuration_pci_am1_reg[12] ;
  assign \new_[10517]_  = \\configuration_pci_am1_reg[11] ;
  assign \new_[10518]_  = \\configuration_pci_am1_reg[13] ;
  assign \new_[10519]_  = \\configuration_pci_am1_reg[18] ;
  assign \new_[10520]_  = \\configuration_pci_am1_reg[17] ;
  assign \new_[10521]_  = \\configuration_pci_am1_reg[20] ;
  assign \new_[10522]_  = \\configuration_pci_am1_reg[14] ;
  assign \new_[10523]_  = \\configuration_pci_am1_reg[22] ;
  assign \new_[10524]_  = \\configuration_pci_am1_reg[23] ;
  assign \new_[10525]_  = \\configuration_pci_am1_reg[25] ;
  assign \new_[10526]_  = \\configuration_pci_am1_reg[19] ;
  assign \new_[10527]_  = \\configuration_pci_am1_reg[29] ;
  assign \new_[10528]_  = \\configuration_pci_am1_reg[31] ;
  assign \new_[10529]_  = \\configuration_pci_am1_reg[30] ;
  assign \new_[10530]_  = \\configuration_pci_am1_reg[28] ;
  assign \new_[10531]_  = ~\new_[9906]_  | (~\new_[11667]_  & ~\new_[17476]_ );
  assign \new_[10532]_  = ~\new_[9908]_  | (~\new_[11672]_  & ~\new_[17476]_ );
  assign \new_[10533]_  = ~\new_[9985]_  | (~\new_[11669]_  & ~\new_[17258]_ );
  assign \new_[10534]_  = \\pci_target_unit_wishbone_master_read_count_reg[0] ;
  assign \new_[10535]_  = ~\new_[9907]_  | (~\new_[11671]_  & ~\new_[17258]_ );
  assign n7735 = ~\new_[11118]_  | (~\new_[14229]_  & ~\new_[13723]_ );
  assign n7750 = ~\new_[11119]_  | (~\new_[14229]_  & ~\new_[13722]_ );
  assign n7745 = ~\new_[11120]_  | (~\new_[14229]_  & ~\new_[13724]_ );
  assign n8715 = ~\new_[11121]_  | (~\new_[14229]_  & ~\new_[13725]_ );
  assign n7740 = ~\new_[11125]_  | (~\new_[14229]_  & ~\new_[13863]_ );
  assign n7760 = ~\new_[11122]_  | (~\new_[14229]_  & ~\new_[13862]_ );
  assign n7755 = ~\new_[11127]_  | (~\new_[14229]_  & ~\new_[13860]_ );
  assign n8685 = ~\new_[11129]_  | (~\new_[14229]_  & ~\new_[13864]_ );
  assign n7765 = ~\new_[11103]_  & (~\new_[16725]_  | ~n16670);
  assign n7770 = ~\new_[11102]_  & (~\new_[16724]_  | ~n16665);
  assign n7795 = \new_[16011]_  ? \new_[11680]_  : \new_[19678]_ ;
  assign n7800 = \new_[16018]_  ? \new_[11679]_  : \new_[18788]_ ;
  assign n9045 = \new_[15929]_  ? \new_[11680]_  : \new_[19865]_ ;
  assign n7805 = \new_[16128]_  ? \new_[11679]_  : \new_[18840]_ ;
  assign n9025 = \new_[16019]_  ? \new_[11681]_  : \new_[18617]_ ;
  assign n7810 = \new_[15996]_  ? \new_[11679]_  : \new_[18774]_ ;
  assign n9040 = \new_[16014]_  ? \new_[13577]_  : \new_[18920]_ ;
  assign n7815 = \new_[15998]_  ? \new_[11678]_  : \new_[18900]_ ;
  assign n9035 = \new_[16005]_  ? \new_[11673]_  : \new_[18069]_ ;
  assign n7820 = \new_[16001]_  ? \new_[11675]_  : \new_[18940]_ ;
  assign n9030 = \new_[16022]_  ? \new_[11681]_  : \new_[18941]_ ;
  assign n7825 = \new_[16007]_  ? \new_[11678]_  : \new_[19487]_ ;
  assign n7830 = \new_[16000]_  ? \new_[11674]_  : \new_[19183]_ ;
  assign n7835 = \new_[15999]_  ? \new_[11676]_  : \new_[19595]_ ;
  assign n9015 = \new_[16020]_  ? \new_[13577]_  : \new_[18522]_ ;
  assign n7840 = \new_[16010]_  ? \new_[11674]_  : \new_[19399]_ ;
  assign n9020 = \new_[16015]_  ? \new_[11677]_  : \new_[18476]_ ;
  assign n7845 = \new_[15997]_  ? \new_[11680]_  : \new_[18542]_ ;
  assign n9010 = \new_[16012]_  ? \new_[11677]_  : \new_[18935]_ ;
  assign n7850 = \new_[16131]_  ? \new_[11679]_  : \new_[18353]_ ;
  assign n8990 = \new_[16009]_  ? \new_[11675]_  : \new_[18539]_ ;
  assign n7855 = \new_[16133]_  ? \new_[11681]_  : \new_[18944]_ ;
  assign n8995 = \new_[16008]_  ? \new_[11679]_  : \new_[17839]_ ;
  assign n7860 = \new_[16006]_  ? \new_[11679]_  : \new_[18312]_ ;
  assign n9005 = \new_[16004]_  ? \new_[11678]_  : \new_[19121]_ ;
  assign n7865 = \new_[13920]_  ? \new_[11679]_  : \new_[18514]_ ;
  assign n9000 = \new_[16003]_  ? \new_[11674]_  : \new_[18874]_ ;
  assign n7870 = \new_[16136]_  ? \new_[11675]_  : \new_[18925]_ ;
  assign n7875 = \new_[16002]_  ? \new_[11680]_  : \new_[18194]_ ;
  assign n7880 = \new_[16023]_  ? \new_[11678]_  : \new_[17919]_ ;
  assign n8985 = \new_[16021]_  ? \new_[11678]_  : \new_[19258]_ ;
  assign n7885 = \new_[16017]_  ? \new_[11680]_  : \new_[18197]_ ;
  assign n8975 = \new_[16016]_  ? \new_[11674]_  : \new_[18547]_ ;
  assign n7890 = \new_[16248]_  ? \new_[11676]_  : \new_[18293]_ ;
  assign n8970 = \new_[16238]_  ? \new_[11681]_  : \new_[18083]_ ;
  assign n7895 = \new_[16149]_  ? \new_[11675]_  : \new_[18061]_ ;
  assign n7900 = \new_[16235]_  ? \new_[11677]_  : \new_[18510]_ ;
  assign n7905 = \new_[16269]_  ? \new_[11675]_  : \new_[19017]_ ;
  assign n8965 = \new_[16167]_  ? \new_[11680]_  : \new_[18076]_ ;
  assign n7910 = \new_[16188]_  ? \new_[11673]_  : \new_[18262]_ ;
  assign n7915 = \new_[16282]_  ? \new_[11678]_  : \new_[18597]_ ;
  assign n7920 = \new_[16278]_  ? \new_[11675]_  : \new_[18932]_ ;
  assign n8940 = \new_[16257]_  ? \new_[11677]_  : \new_[19000]_ ;
  assign n7925 = \new_[16277]_  ? \new_[11676]_  : \new_[18107]_ ;
  assign n7930 = \new_[16237]_  ? \new_[11681]_  : \new_[19826]_ ;
  assign n7935 = \new_[16437]_  ? \new_[11680]_  : \new_[19407]_ ;
  assign n8960 = \new_[16284]_  ? \new_[11679]_  : \new_[18835]_ ;
  assign n7940 = \new_[16275]_  ? \new_[11677]_  : \new_[18179]_ ;
  assign n8945 = \new_[16286]_  ? \new_[11678]_  : \new_[18178]_ ;
  assign n7945 = \new_[16283]_  ? \new_[11677]_  : \new_[18174]_ ;
  assign n8915 = \new_[16273]_  ? \new_[11675]_  : \new_[18175]_ ;
  assign n7950 = \new_[16274]_  ? \new_[11679]_  : \new_[18169]_ ;
  assign n8930 = \new_[16268]_  ? \new_[11679]_  : \new_[18168]_ ;
  assign n7955 = \new_[16266]_  ? \new_[11673]_  : \new_[18160]_ ;
  assign n8860 = \new_[16239]_  ? \new_[11680]_  : \new_[18161]_ ;
  assign n7960 = \new_[16249]_  ? \new_[11675]_  : \new_[19114]_ ;
  assign n8895 = \new_[16242]_  ? \new_[11675]_  : \new_[18580]_ ;
  assign n7965 = \new_[16162]_  ? \new_[11680]_  : \new_[19737]_ ;
  assign n8900 = \new_[13923]_  ? \new_[11680]_  : \new_[18908]_ ;
  assign n7970 = \new_[16279]_  ? \new_[11681]_  : \new_[17892]_ ;
  assign n7975 = \new_[16258]_  ? \new_[11679]_  : \new_[18096]_ ;
  assign n7980 = \new_[16256]_  ? \new_[11681]_  : \new_[19309]_ ;
  assign n8870 = \new_[16245]_  ? \new_[11678]_  : \new_[19021]_ ;
  assign n7985 = \new_[16246]_  ? \new_[11680]_  : \new_[19820]_ ;
  assign n7990 = \new_[16272]_  ? \new_[11680]_  : \new_[18924]_ ;
  assign n7995 = \new_[16247]_  ? \new_[11678]_  : \new_[17900]_ ;
  assign n8820 = \new_[16241]_  ? \new_[11676]_  : \new_[19679]_ ;
  assign n8000 = \new_[16255]_  ? \new_[11680]_  : \new_[19739]_ ;
  assign n8005 = \new_[16280]_  ? \new_[11676]_  : \new_[19043]_ ;
  assign n8010 = \new_[16270]_  ? \new_[11673]_  : \new_[17912]_ ;
  assign n8840 = \new_[16264]_  ? \new_[11678]_  : \new_[19821]_ ;
  assign n8015 = \new_[16260]_  ? \new_[11676]_  : \new_[17909]_ ;
  assign n8855 = \new_[16252]_  ? \new_[11676]_  : \new_[17924]_ ;
  assign n8020 = \new_[16243]_  ? \new_[11677]_  : \new_[18203]_ ;
  assign n8845 = \new_[16263]_  ? \new_[11674]_  : \new_[19026]_ ;
  assign n8025 = \new_[16271]_  ? \new_[11674]_  : \new_[19463]_ ;
  assign n8030 = \new_[16240]_  ? \new_[11681]_  : \new_[19124]_ ;
  assign n8035 = \new_[16281]_  ? \new_[13577]_  : \new_[19342]_ ;
  assign n8830 = \new_[16267]_  ? \new_[11677]_  : \new_[19741]_ ;
  assign n8040 = \new_[16190]_  ? \new_[11680]_  : \new_[19819]_ ;
  assign n8815 = \new_[16198]_  ? \new_[11676]_  : \new_[19459]_ ;
  assign n8045 = \new_[16154]_  ? \new_[11681]_  : \new_[18331]_ ;
  assign n8810 = \new_[16261]_  ? \new_[11673]_  : \new_[19818]_ ;
  assign n8050 = \new_[16413]_  ? \new_[11680]_  : \new_[18323]_ ;
  assign n8055 = \new_[16276]_  ? \new_[11677]_  : \new_[19816]_ ;
  assign n8060 = \new_[16244]_  ? \new_[11678]_  : \new_[19334]_ ;
  assign n8775 = \new_[16285]_  ? \new_[11677]_  : \new_[19807]_ ;
  assign n8065 = \new_[16236]_  ? \new_[11679]_  : \new_[19812]_ ;
  assign n8800 = \new_[16254]_  ? \new_[11676]_  : \new_[19108]_ ;
  assign n8070 = \new_[16262]_  ? \new_[11681]_  : \new_[19815]_ ;
  assign n8805 = \new_[16259]_  ? \new_[11676]_  : \new_[19726]_ ;
  assign n8075 = \new_[13922]_  ? \new_[11676]_  : \new_[19704]_ ;
  assign n8080 = \new_[16234]_  ? \new_[11680]_  : \new_[18302]_ ;
  assign n8085 = \new_[16250]_  ? \new_[11679]_  : \new_[19317]_ ;
  assign n8795 = \new_[16139]_  ? \new_[11679]_  : \new_[19833]_ ;
  assign n8090 = \new_[16206]_  ? \new_[11679]_  : \new_[19670]_ ;
  assign n8095 = \new_[16251]_  ? \new_[11677]_  : \new_[18284]_ ;
  assign n8100 = \new_[16265]_  ? \new_[11679]_  : \new_[17955]_ ;
  assign n8770 = \new_[16253]_  ? \new_[11678]_  : \new_[17853]_ ;
  assign n8105 = \new_[16526]_  ? \new_[11677]_  : \new_[19743]_ ;
  assign n8110 = \new_[16527]_  ? \new_[11674]_  : \new_[17964]_ ;
  assign n8115 = \new_[16498]_  ? \new_[11674]_  : \new_[19291]_ ;
  assign n8790 = \new_[16521]_  ? \new_[11675]_  : \new_[19292]_ ;
  assign n8120 = \new_[16525]_  ? \new_[11679]_  : \new_[18562]_ ;
  assign n8780 = \new_[16542]_  ? \new_[11678]_  : \new_[19810]_ ;
  assign n8125 = \new_[16540]_  ? \new_[11678]_  : \new_[19811]_ ;
  assign n8785 = \new_[16539]_  ? \new_[11678]_  : \new_[19138]_ ;
  assign n8130 = \new_[16537]_  ? \new_[11678]_  : \new_[19266]_ ;
  assign n8135 = \new_[16535]_  ? \new_[11673]_  : \new_[19808]_ ;
  assign n8140 = \new_[16492]_  ? \new_[11679]_  : \new_[18162]_ ;
  assign n7640 = \new_[16531]_  ? \new_[11680]_  : \new_[17994]_ ;
  assign n8145 = \new_[16496]_  ? \new_[11675]_  : \new_[19148]_ ;
  assign n8680 = \new_[16522]_  ? \new_[11679]_  : \new_[17998]_ ;
  assign n8150 = \new_[16529]_  ? \new_[11679]_  : \new_[17997]_ ;
  assign n8760 = \new_[16480]_  ? \new_[11677]_  : \new_[19725]_ ;
  assign n8155 = \new_[16538]_  ? \new_[11677]_  : \new_[19560]_ ;
  assign n8160 = \new_[16519]_  ? \new_[11680]_  : \new_[19806]_ ;
  assign n8165 = \new_[16532]_  ? \new_[11676]_  : \new_[19512]_ ;
  assign n8755 = \new_[16524]_  ? \new_[11674]_  : \new_[18157]_ ;
  assign n8170 = \new_[16541]_  ? \new_[11674]_  : \new_[19582]_ ;
  assign n8175 = \new_[16528]_  ? \new_[11681]_  : \new_[18989]_ ;
  assign n8180 = \new_[16520]_  ? \new_[11678]_  : \new_[19151]_ ;
  assign n8750 = \new_[16544]_  ? \new_[11679]_  : \new_[19724]_ ;
  assign n8185 = \new_[16534]_  ? \new_[11681]_  : \new_[19669]_ ;
  assign n8190 = \new_[13925]_  ? \new_[11678]_  : \new_[18021]_ ;
  assign n8195 = \new_[16533]_  ? \new_[11678]_  : \new_[19158]_ ;
  assign n8735 = \new_[16482]_  ? \new_[11681]_  : \new_[19164]_ ;
  assign n8200 = \new_[16536]_  ? \new_[11681]_  : \new_[19160]_ ;
  assign n8745 = \new_[16481]_  ? \new_[11680]_  : \new_[19803]_ ;
  assign n8205 = \new_[16530]_  ? \new_[11674]_  : \new_[19162]_ ;
  assign n8740 = \new_[16456]_  ? \new_[11680]_  : \new_[19650]_ ;
  assign n8210 = \new_[16478]_  ? \new_[11674]_  : \new_[18024]_ ;
  assign n8220 = \new_[16287]_  ? \new_[11678]_  : \new_[19801]_ ;
  assign n8225 = \new_[16334]_  ? \new_[11676]_  : \new_[19168]_ ;
  assign n8730 = \new_[16342]_  ? \new_[11680]_  : \new_[18038]_ ;
  assign n8230 = \new_[16340]_  ? \new_[11674]_  : \new_[17985]_ ;
  assign n8720 = \new_[16288]_  ? \new_[11674]_  : \new_[19643]_ ;
  assign n8235 = \new_[16289]_  ? \new_[11676]_  : \new_[19169]_ ;
  assign n8725 = \new_[16347]_  ? \new_[11676]_  : \new_[17978]_ ;
  assign n8240 = \new_[16348]_  ? \new_[11673]_  : \new_[19802]_ ;
  assign n8245 = \new_[16168]_  ? \new_[11681]_  : \new_[19747]_ ;
  assign n8250 = \new_[16290]_  ? \new_[11678]_  : \new_[18067]_ ;
  assign n8710 = \new_[16291]_  ? \new_[11675]_  : \new_[19799]_ ;
  assign n8255 = \new_[16292]_  ? \new_[11678]_  : \new_[18055]_ ;
  assign n8675 = \new_[16339]_  ? \new_[11681]_  : \new_[19174]_ ;
  assign n8260 = \new_[16293]_  ? \new_[11678]_  : \new_[19672]_ ;
  assign n8705 = \new_[16338]_  ? \new_[11679]_  : \new_[19748]_ ;
  assign n8265 = \new_[16337]_  ? \new_[11674]_  : \new_[18062]_ ;
  assign n8270 = \new_[16294]_  ? \new_[11679]_  : \new_[19653]_ ;
  assign n8275 = \new_[16295]_  ? \new_[11676]_  : \new_[19182]_ ;
  assign n8700 = \new_[16296]_  ? \new_[11677]_  : \new_[19186]_ ;
  assign n8280 = \new_[13927]_  ? \new_[11673]_  : \new_[18079]_ ;
  assign n8690 = \new_[16328]_  ? \new_[11674]_  : \new_[19623]_ ;
  assign n8285 = \new_[16297]_  ? \new_[11675]_  : \new_[19202]_ ;
  assign n8695 = \new_[16327]_  ? \new_[11676]_  : \new_[17889]_ ;
  assign n8290 = \new_[16298]_  ? \new_[11676]_  : \new_[19617]_ ;
  assign n8295 = \new_[16326]_  ? \new_[11677]_  : \new_[18092]_ ;
  assign n8300 = \new_[16325]_  ? \new_[11680]_  : \new_[19363]_ ;
  assign n8660 = \new_[16324]_  ? \new_[11677]_  : \new_[18147]_ ;
  assign n8305 = \new_[16299]_  ? \new_[11681]_  : \new_[18871]_ ;
  assign n8665 = \new_[16319]_  ? \new_[11678]_  : \new_[19016]_ ;
  assign n8310 = \new_[16346]_  ? \new_[11679]_  : \new_[19795]_ ;
  assign n8670 = \new_[16300]_  ? \new_[11674]_  : \new_[19210]_ ;
  assign n8315 = \new_[16301]_  ? \new_[11676]_  : \new_[18868]_ ;
  assign n8320 = \new_[16302]_  ? \new_[11677]_  : \new_[19752]_ ;
  assign n8325 = \new_[16303]_  ? \new_[11673]_  : \new_[18110]_ ;
  assign n8655 = \new_[16304]_  ? \new_[11681]_  : \new_[19211]_ ;
  assign n8330 = \new_[16178]_  ? \new_[11676]_  : \new_[19217]_ ;
  assign n8335 = \new_[16305]_  ? \new_[11676]_  : \new_[18113]_ ;
  assign n8340 = \new_[16163]_  ? \new_[11679]_  : \new_[18111]_ ;
  assign n8650 = \new_[16306]_  ? \new_[11681]_  : \new_[19212]_ ;
  assign n8345 = \new_[16307]_  ? \new_[11681]_  : \new_[19863]_ ;
  assign n8645 = \new_[16407]_  ? \new_[11674]_  : \new_[19682]_ ;
  assign n8350 = \new_[16335]_  ? \new_[11680]_  : \new_[19784]_ ;
  assign n8640 = \new_[16308]_  ? \new_[11674]_  : \new_[19598]_ ;
  assign n8355 = \new_[16441]_  ? \new_[11673]_  : \new_[19218]_ ;
  assign n8630 = \new_[16309]_  ? \new_[11677]_  : \new_[18126]_ ;
  assign n8360 = \new_[16310]_  ? \new_[11676]_  : \new_[18120]_ ;
  assign n8635 = \new_[16311]_  ? \new_[11676]_  : \new_[19584]_ ;
  assign n8365 = \new_[16330]_  ? \new_[11681]_  : \new_[18159]_ ;
  assign n8370 = \new_[16177]_  ? \new_[11677]_  : \new_[19232]_ ;
  assign n8375 = \new_[16312]_  ? \new_[11673]_  : \new_[18306]_ ;
  assign n8620 = \new_[16444]_  ? \new_[11679]_  : \new_[19838]_ ;
  assign n8380 = \new_[16313]_  ? \new_[11674]_  : \new_[19577]_ ;
  assign n8625 = \new_[13929]_  ? \new_[11680]_  : \new_[19233]_ ;
  assign n8385 = \new_[16333]_  ? \new_[11677]_  : \new_[18166]_ ;
  assign n7730 = \new_[16314]_  ? \new_[11677]_  : \new_[19716]_ ;
  assign n8390 = \new_[16321]_  ? \new_[11675]_  : \new_[19756]_ ;
  assign n7645 = \new_[16315]_  ? \new_[11675]_  : \new_[19792]_ ;
  assign n8395 = \new_[16316]_  ? \new_[11674]_  : \new_[18212]_ ;
  assign n7705 = \new_[16317]_  ? \new_[11681]_  : \new_[19246]_ ;
  assign n8400 = \new_[16322]_  ? \new_[11678]_  : \new_[19791]_ ;
  assign n7700 = \new_[16488]_  ? \new_[11681]_  : \new_[19235]_ ;
  assign n8405 = \new_[16546]_  ? \new_[11679]_  : \new_[19208]_ ;
  assign n7695 = \new_[16447]_  ? \new_[11677]_  : \new_[19562]_ ;
  assign n8410 = \new_[16448]_  ? \new_[11675]_  : \new_[18086]_ ;
  assign n8415 = \new_[16547]_  ? \new_[11676]_  : \new_[19015]_ ;
  assign n8420 = \new_[16555]_  ? \new_[11676]_  : \new_[19082]_ ;
  assign \new_[10744]_  = \\configuration_pci_ba1_bit31_8_reg[31] ;
  assign n7710 = \new_[16548]_  ? \new_[11680]_  : \new_[19785]_ ;
  assign n8425 = \new_[16559]_  ? \new_[11681]_  : \new_[19137]_ ;
  assign n8430 = \new_[16556]_  ? \new_[11673]_  : \new_[19256]_ ;
  assign n8435 = \new_[16549]_  ? \new_[11673]_  : \new_[18200]_ ;
  assign n7685 = \new_[16564]_  ? \new_[11678]_  : \new_[19790]_ ;
  assign n8440 = \new_[16550]_  ? \new_[11679]_  : \new_[18201]_ ;
  assign n7690 = \new_[16560]_  ? \new_[11677]_  : \new_[18202]_ ;
  assign n8445 = \new_[16486]_  ? \new_[11676]_  : \new_[19673]_ ;
  assign n7675 = \new_[16490]_  ? \new_[11681]_  : \new_[17933]_ ;
  assign n8450 = \new_[16571]_  ? \new_[11674]_  : \new_[18213]_ ;
  assign n7680 = \new_[16570]_  ? \new_[11679]_  : \new_[19120]_ ;
  assign n8455 = \new_[16568]_  ? \new_[11676]_  : \new_[19789]_ ;
  assign n7660 = \new_[16566]_  ? \new_[11673]_  : \new_[19759]_ ;
  assign n8460 = \new_[16565]_  ? \new_[11678]_  : \new_[19117]_ ;
  assign \new_[10759]_  = \\wishbone_slave_unit_wishbone_slave_img_hit_reg[1] ;
  assign n8465 = \new_[16562]_  ? \new_[11681]_  : \new_[19013]_ ;
  assign n8470 = \new_[16567]_  ? \new_[11680]_  : \new_[19271]_ ;
  assign n7670 = \new_[16454]_  ? \new_[11677]_  : \new_[19538]_ ;
  assign n8475 = \new_[16551]_  ? \new_[11680]_  : \new_[18223]_ ;
  assign n7665 = \new_[16552]_  ? \new_[11677]_  : \new_[18222]_ ;
  assign n8480 = \new_[13928]_  ? \new_[11680]_  : \new_[19054]_ ;
  assign n7650 = \new_[16553]_  ? \new_[11677]_  : \new_[18258]_ ;
  assign n8485 = \new_[16554]_  ? \new_[11673]_  : \new_[19782]_ ;
  assign n8490 = \new_[16569]_  ? \new_[11679]_  : \new_[19783]_ ;
  assign n8495 = \new_[16494]_  ? \new_[11677]_  : \new_[19764]_ ;
  assign n8980 = \new_[16449]_  ? \new_[11676]_  : \new_[19765]_ ;
  assign n8500 = \new_[16563]_  ? \new_[13577]_  : \new_[17838]_ ;
  assign n8505 = \new_[16561]_  ? \new_[11676]_  : \new_[19864]_ ;
  assign \new_[10773]_  = \\configuration_pci_ba1_bit31_8_reg[8] ;
  assign \new_[10774]_  = \\configuration_pci_ba1_bit31_8_reg[9] ;
  assign \new_[10775]_  = \\configuration_pci_ba1_bit31_8_reg[22] ;
  assign n8510 = \new_[16028]_  ? \new_[11675]_  : \new_[18588]_ ;
  assign n8920 = \new_[16026]_  ? \new_[11681]_  : \new_[19776]_ ;
  assign n8515 = \new_[16043]_  ? \new_[11675]_  : \new_[19779]_ ;
  assign n8950 = \new_[16025]_  ? \new_[11674]_  : \new_[19780]_ ;
  assign n8520 = \new_[16044]_  ? \new_[11673]_  : \new_[19768]_ ;
  assign n8955 = \new_[16045]_  ? \new_[11674]_  : \new_[18579]_ ;
  assign n8525 = \new_[16036]_  ? \new_[11677]_  : \new_[18253]_ ;
  assign n8935 = \new_[16046]_  ? \new_[11676]_  : \new_[18619]_ ;
  assign n8530 = \new_[16047]_  ? \new_[11674]_  : \new_[19302]_ ;
  assign n8925 = \new_[16048]_  ? \new_[11677]_  : \new_[19710]_ ;
  assign n8535 = \new_[16049]_  ? \new_[11680]_  : \new_[18263]_ ;
  assign n8540 = \new_[16135]_  ? \new_[11679]_  : \new_[19777]_ ;
  assign n8545 = \new_[16024]_  ? \new_[11674]_  : \new_[19297]_ ;
  assign n8880 = \new_[15916]_  ? \new_[11677]_  : \new_[19774]_ ;
  assign n8550 = \new_[16050]_  ? \new_[11679]_  : \new_[19400]_ ;
  assign n8910 = \new_[16051]_  ? \new_[11678]_  : \new_[18422]_ ;
  assign n8555 = \new_[16039]_  ? \new_[11676]_  : \new_[18380]_ ;
  assign n8905 = \new_[16041]_  ? \new_[11675]_  : \new_[18938]_ ;
  assign \new_[10794]_  = \\configuration_pci_ba1_bit31_8_reg[28] ;
  assign n8560 = \new_[16029]_  ? \new_[11681]_  : \new_[18036]_ ;
  assign n8565 = \new_[16052]_  ? \new_[11678]_  : \new_[19008]_ ;
  assign n8570 = \new_[16042]_  ? \new_[11676]_  : \new_[18350]_ ;
  assign n8890 = \new_[16053]_  ? \new_[11675]_  : \new_[19773]_ ;
  assign n8575 = \new_[16040]_  ? \new_[11678]_  : \new_[19685]_ ;
  assign n8885 = \new_[16054]_  ? \new_[11678]_  : \new_[18356]_ ;
  assign n8580 = \new_[16055]_  ? \new_[11681]_  : \new_[19732]_ ;
  assign n8875 = \new_[13930]_  ? \new_[11677]_  : \new_[19434]_ ;
  assign n8585 = \new_[16037]_  ? \new_[11678]_  : \new_[19438]_ ;
  assign n8590 = \new_[16034]_  ? \new_[11681]_  : \new_[19771]_ ;
  assign n8595 = \new_[16033]_  ? \new_[11681]_  : \new_[19772]_ ;
  assign n8865 = \new_[16056]_  ? \new_[11681]_  : \new_[18367]_ ;
  assign n8600 = \new_[16057]_  ? \new_[11674]_  : \new_[19347]_ ;
  assign n8765 = \new_[16058]_  ? \new_[11674]_  : \new_[18370]_ ;
  assign n8605 = \new_[16059]_  ? \new_[11680]_  : \new_[19435]_ ;
  assign n8825 = \new_[16323]_  ? \new_[11680]_  : \new_[19709]_ ;
  assign n8610 = \new_[16140]_  ? \new_[11674]_  : \new_[18373]_ ;
  assign n8835 = \new_[16318]_  ? \new_[11680]_  : \new_[18419]_ ;
  assign n8615 = \new_[16349]_  ? \new_[11674]_  : \new_[19686]_ ;
  assign n8850 = \new_[16350]_  ? \new_[11674]_  : \new_[19354]_ ;
  assign n8215 = \new_[16351]_  ? \new_[11674]_  : \new_[17896]_ ;
  assign \new_[10816]_  = \\configuration_pci_ba1_bit31_8_reg[24] ;
  assign n7775 = \new_[15967]_  ? \new_[11675]_  : \new_[10074]_ ;
  assign n7655 = \new_[10006]_  ? \new_[11675]_  : n17035;
  assign n7780 = \new_[10012]_  ? \new_[11675]_  : n17065;
  assign n7785 = \new_[10077]_  ? \new_[11675]_  : n17020;
  assign n7790 = \new_[10074]_  ? \new_[11675]_  : \new_[10077]_ ;
  assign \new_[10822]_  = \\configuration_pci_ba1_bit31_8_reg[17] ;
  assign \new_[10823]_  = wishbone_slave_unit_pci_initiator_if_current_last_reg;
  assign \new_[10824]_  = \\wishbone_slave_unit_wishbone_slave_img_hit_reg[0] ;
  assign \new_[10825]_  = ~\new_[20332]_ ;
  assign \new_[10826]_  = ~\new_[18729]_  | ~\new_[17096]_  | ~\new_[11865]_ ;
  assign \new_[10827]_  = ~\new_[16517]_  | ~\new_[15891]_  | ~\new_[11874]_ ;
  assign \new_[10828]_  = ~\new_[16655]_  & (~\new_[11887]_  | ~\new_[15324]_ );
  assign \new_[10829]_  = ~\new_[16434]_  & (~\new_[11888]_  | ~\new_[15747]_ );
  assign \new_[10830]_  = ~\new_[10974]_ ;
  assign \new_[10831]_  = \new_[11206]_  | \new_[16655]_ ;
  assign n7715 = ~\new_[11203]_  | (~\new_[13298]_  & ~\new_[15899]_ );
  assign n7720 = ~\new_[11204]_  | (~\new_[13298]_  & ~\new_[15934]_ );
  assign n7725 = ~\new_[11205]_  | (~\new_[13298]_  & ~\new_[16122]_ );
  assign \new_[10835]_  = ~\new_[20398]_  | (~\new_[13130]_  & ~\new_[11328]_ );
  assign \new_[10836]_  = ~\new_[11135]_  | ~\new_[9904]_ ;
  assign \new_[10837]_  = ~\new_[11135]_  | ~\new_[9905]_ ;
  assign \new_[10838]_  = (~\new_[11612]_  | ~\new_[9993]_ ) & (~\new_[13117]_  | ~\new_[15931]_ );
  assign \new_[10839]_  = (~\new_[11612]_  | ~\new_[9994]_ ) & (~\new_[13117]_  | ~\new_[15801]_ );
  assign \new_[10840]_  = (~\new_[11612]_  | ~\new_[9989]_ ) & (~\new_[13117]_  | ~\new_[15901]_ );
  assign \new_[10841]_  = (~\new_[11613]_  | ~\new_[9995]_ ) & (~\new_[13118]_  | ~\new_[15931]_ );
  assign \new_[10842]_  = (~\new_[11613]_  | ~\new_[9988]_ ) & (~\new_[13118]_  | ~\new_[15801]_ );
  assign \new_[10843]_  = (~\new_[11613]_  | ~\new_[9996]_ ) & (~\new_[13118]_  | ~\new_[15901]_ );
  assign \new_[10844]_  = (~\new_[11612]_  | ~\new_[9987]_ ) & (~\new_[16120]_  | ~\new_[13117]_ );
  assign \new_[10845]_  = \\configuration_pci_am1_reg[26] ;
  assign \new_[10846]_  = \\configuration_pci_am1_reg[8] ;
  assign \new_[10847]_  = \\configuration_pci_am1_reg[9] ;
  assign \new_[10848]_  = \\configuration_pci_am1_reg[27] ;
  assign \new_[10849]_  = (~\new_[11614]_  | ~\new_[9997]_ ) & (~\new_[13121]_  | ~\new_[15931]_ );
  assign \new_[10850]_  = (~\new_[11614]_  | ~\new_[9998]_ ) & (~\new_[13121]_  | ~\new_[15801]_ );
  assign \new_[10851]_  = (~\new_[11614]_  | ~n17430) & (~\new_[13121]_  | ~\new_[15901]_ );
  assign \new_[10852]_  = (~\new_[11614]_  | ~\new_[10046]_ ) & (~\new_[13121]_  | ~\new_[16120]_ );
  assign \new_[10853]_  = \\wishbone_slave_unit_wishbone_slave_c_state_reg[1] ;
  assign \new_[10854]_  = \\configuration_pci_ta1_reg[10] ;
  assign \new_[10855]_  = pci_target_unit_wishbone_master_read_bound_reg;
  assign n9365 = ~\new_[11636]_  | (~\new_[15022]_  & ~\new_[12575]_ );
  assign \new_[10857]_  = \\configuration_pci_ta1_reg[29] ;
  assign \new_[10858]_  = \\configuration_pci_ta1_reg[16] ;
  assign \new_[10859]_  = \\wishbone_slave_unit_pci_initiator_if_read_count_reg[2] ;
  assign \new_[10860]_  = \\configuration_pci_ta1_reg[17] ;
  assign \new_[10861]_  = \\configuration_pci_ta1_reg[18] ;
  assign \new_[10862]_  = \\configuration_pci_ta1_reg[20] ;
  assign \new_[10863]_  = \\configuration_pci_ta1_reg[21] ;
  assign \new_[10864]_  = \\configuration_pci_ta1_reg[24] ;
  assign \new_[10865]_  = \\configuration_pci_ta1_reg[23] ;
  assign \new_[10866]_  = \\configuration_pci_ta1_reg[30] ;
  assign \new_[10867]_  = \\configuration_pci_ta1_reg[28] ;
  assign \new_[10868]_  = \\configuration_pci_ta1_reg[31] ;
  assign \new_[10869]_  = \\configuration_pci_ta1_reg[14] ;
  assign \new_[10870]_  = wishbone_slave_unit_pci_initiator_if_err_recovery_reg;
  assign \new_[10871]_  = ~\new_[10043]_  | (~\new_[12290]_  & ~\new_[17476]_ );
  assign \new_[10872]_  = ~\new_[10000]_  | (~\new_[12290]_  & ~\new_[17258]_ );
  assign \new_[10873]_  = ~\new_[10001]_  | (~\new_[12289]_  & ~\new_[17258]_ );
  assign \new_[10874]_  = ~\new_[10042]_  | (~\new_[12289]_  & ~\new_[17476]_ );
  assign \new_[10875]_  = ~\new_[10002]_  | (~\new_[12295]_  & ~\new_[16838]_ );
  assign \new_[10876]_  = \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1] ;
  assign \new_[10877]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][37] ;
  assign \new_[10878]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][37] ;
  assign \new_[10879]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][37] ;
  assign \new_[10880]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][37] ;
  assign \new_[10881]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][37] ;
  assign \new_[10882]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][37] ;
  assign \new_[10883]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][37] ;
  assign \new_[10884]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][37] ;
  assign \new_[10885]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][37] ;
  assign \new_[10886]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][37] ;
  assign \new_[10887]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][37] ;
  assign \new_[10888]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][37] ;
  assign n9370 = \new_[19517]_  ? \new_[12293]_  : \new_[10416]_ ;
  assign n9375 = \new_[18261]_  ? \new_[12293]_  : \new_[10417]_ ;
  assign n9380 = \new_[18321]_  ? \new_[12292]_  : \new_[10418]_ ;
  assign n9095 = \new_[19530]_  ? \new_[12292]_  : \new_[10359]_ ;
  assign n9385 = \new_[18951]_  ? \new_[12293]_  : \new_[10419]_ ;
  assign n9110 = \new_[19318]_  ? \new_[12293]_  : \new_[10362]_ ;
  assign n9390 = \new_[19178]_  ? \new_[12292]_  : \new_[10420]_ ;
  assign n9115 = \new_[18308]_  ? \new_[12292]_  : \new_[10363]_ ;
  assign n9395 = \new_[19111]_  ? \new_[12293]_  : \new_[10421]_ ;
  assign n9400 = \new_[17867]_  ? \new_[12292]_  : \new_[10422]_ ;
  assign n9405 = \new_[17840]_  ? \new_[12293]_  : \new_[10423]_ ;
  assign n9100 = \new_[19083]_  ? \new_[12293]_  : \new_[10360]_ ;
  assign n9410 = \new_[18946]_  ? \new_[12293]_  : \new_[10424]_ ;
  assign n9105 = \new_[18534]_  ? \new_[12293]_  : \new_[10361]_ ;
  assign n9415 = \new_[18337]_  ? \new_[12293]_  : \new_[10425]_ ;
  assign n9065 = \new_[19845]_  ? \new_[12292]_  : \new_[10353]_ ;
  assign n9420 = \new_[19341]_  ? \new_[12292]_  : \new_[10426]_ ;
  assign n9425 = \new_[18934]_  ? \new_[12293]_  : \new_[10427]_ ;
  assign n9430 = \new_[18362]_  ? \new_[12292]_  : \new_[10428]_ ;
  assign n9085 = \new_[19381]_  ? \new_[12292]_  : \new_[10357]_ ;
  assign n9435 = \new_[19362]_  ? \new_[12293]_  : \new_[10429]_ ;
  assign n9440 = \new_[18425]_  ? \new_[12292]_  : \new_[10430]_ ;
  assign n9445 = \new_[18435]_  ? \new_[12293]_  : \new_[10431]_ ;
  assign n9465 = \new_[18462]_  ? \new_[12292]_  : \new_[10435]_ ;
  assign n9075 = \new_[18565]_  ? \new_[12293]_  : \new_[10355]_ ;
  assign n9450 = \new_[18664]_  ? \new_[12292]_  : \new_[10432]_ ;
  assign n9070 = \new_[18481]_  ? \new_[12292]_  : \new_[10354]_ ;
  assign n9050 = \new_[18926]_  ? \new_[12292]_  : \new_[10350]_ ;
  assign n9455 = \new_[19226]_  ? \new_[12292]_  : \new_[10433]_ ;
  assign n9055 = \new_[18517]_  ? \new_[12293]_  : \new_[10351]_ ;
  assign n9060 = \new_[19497]_  ? \new_[12292]_  : \new_[10352]_ ;
  assign n9460 = \new_[19608]_  ? \new_[12293]_  : \new_[10434]_ ;
  assign \new_[10921]_  = ~\new_[10003]_  | (~\new_[15051]_  & ~\new_[14229]_ );
  assign \new_[10922]_  = ~\new_[10010]_  | (~\new_[14567]_  & ~\new_[14229]_ );
  assign \new_[10923]_  = ~\new_[3738]_  | (~\new_[15064]_  & ~\new_[14229]_ );
  assign \new_[10924]_  = ~\new_[4136]_  | (~\new_[15065]_  & ~\new_[14229]_ );
  assign \new_[10925]_  = ~\new_[10005]_  | (~\new_[15066]_  & ~\new_[14229]_ );
  assign \new_[10926]_  = ~\new_[10009]_  | (~\new_[15063]_  & ~\new_[14229]_ );
  assign \new_[10927]_  = ~\new_[4267]_  | (~\new_[15060]_  & ~\new_[14229]_ );
  assign \new_[10928]_  = ~\new_[10007]_  | (~\new_[15067]_  & ~\new_[14229]_ );
  assign \new_[10929]_  = ~\new_[11675]_  | ~\new_[17656]_ ;
  assign \new_[10930]_  = ~\new_[11675]_  | ~\new_[10006]_ ;
  assign \new_[10931]_  = ~\new_[11675]_  | ~\new_[10004]_ ;
  assign \new_[10932]_  = ~\new_[11675]_  | ~\new_[10012]_ ;
  assign \new_[10933]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][37] ;
  assign \new_[10934]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][37] ;
  assign \new_[10935]_  = ~\new_[12571]_  | ~\new_[5297]_  | ~\new_[11974]_  | ~\new_[20397]_ ;
  assign \new_[10936]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][37] ;
  assign \new_[10937]_  = \new_[17342]_  ^ \new_[12359]_ ;
  assign \new_[10938]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][37] ;
  assign n9150 = ~\new_[11864]_  | ~\new_[11850]_ ;
  assign n9135 = ~\new_[11868]_  | ~\new_[11849]_ ;
  assign n9130 = ~\new_[11869]_  | ~\new_[11852]_ ;
  assign \new_[10942]_  = ~n16890 & (~\new_[12399]_  | ~\new_[17946]_ );
  assign n9140 = ~\new_[13141]_  | (~\new_[15627]_  & ~\new_[12386]_ );
  assign n9145 = ~\new_[13142]_  | (~\new_[15626]_  & ~\new_[12386]_ );
  assign n9490 = (~\new_[16923]_  & ~\new_[16664]_  & ~\new_[17946]_ ) | (~\new_[12399]_  & ~\new_[16459]_  & ~\new_[16506]_ );
  assign n9155 = \new_[10371]_  ? \new_[16782]_  : \new_[12403]_ ;
  assign \new_[10947]_  = ~\new_[9884]_  | ~\new_[15906]_  | ~\new_[12470]_ ;
  assign \new_[10948]_  = ~\new_[16782]_  | ~\new_[11875]_  | ~\new_[15226]_ ;
  assign \new_[10949]_  = ~\new_[11872]_  & ~\new_[16988]_ ;
  assign \new_[10950]_  = ~\new_[16434]_  & (~\new_[12476]_  | ~\new_[15326]_ );
  assign \new_[10951]_  = ~\new_[16434]_  & (~\new_[12477]_  | ~\new_[15305]_ );
  assign \new_[10952]_  = ~\new_[16434]_  & (~\new_[12479]_  | ~\new_[15289]_ );
  assign n9170 = ~\new_[15418]_  & (~\new_[12464]_  | ~\new_[17747]_ );
  assign \new_[10954]_  = ~\new_[11138]_ ;
  assign \new_[10955]_  = ~\new_[16434]_  & (~\new_[20017]_  | ~\new_[15352]_ );
  assign \new_[10956]_  = ~\new_[16658]_  & (~\new_[11970]_  | ~\new_[15310]_ );
  assign n9160 = \new_[12286]_  ? \new_[13804]_  : \new_[10372]_ ;
  assign \new_[10958]_  = ~\new_[11877]_  | ~\new_[16986]_ ;
  assign n9165 = ~\new_[11871]_  & (~\new_[16061]_  | ~n16480);
  assign \new_[10960]_  = ~\new_[13154]_  & (~\new_[17026]_  | ~\new_[12467]_ );
  assign \new_[10961]_  = ~\new_[14217]_  & ~\new_[11870]_ ;
  assign \new_[10962]_  = ~\new_[11876]_  & (~\new_[15388]_  | ~\new_[19948]_ );
  assign n9185 = \new_[11965]_  ? \new_[15274]_  : \new_[19062]_ ;
  assign n9180 = \new_[11969]_  ? \new_[15274]_  : \new_[18715]_ ;
  assign n9485 = \new_[11966]_  ? \new_[15485]_  : \new_[19028]_ ;
  assign n9480 = \new_[11968]_  ? \new_[15274]_  : \new_[19071]_ ;
  assign \new_[10967]_  = (~\new_[16904]_  | ~\new_[13154]_ ) & (~\new_[12470]_  | ~\new_[15907]_ );
  assign n9470 = \new_[11971]_  ? \new_[15484]_  : \new_[18904]_ ;
  assign n9190 = \new_[11972]_  ? \new_[15488]_  : \new_[18732]_ ;
  assign n9475 = \new_[11973]_  ? \new_[15592]_  : \new_[19187]_ ;
  assign n9195 = \new_[11975]_  ? \new_[15274]_  : \new_[18838]_ ;
  assign \new_[10972]_  = \\configuration_pci_ta1_reg[11] ;
  assign \new_[10973]_  = ~\new_[20386]_ ;
  assign \new_[10974]_  = ~\new_[11150]_ ;
  assign \new_[10975]_  = ~\new_[11893]_  | ~\new_[4212]_ ;
  assign \new_[10976]_  = ~\new_[12487]_  | ~\new_[4213]_ ;
  assign \new_[10977]_  = ~\new_[12487]_  | ~\new_[4214]_ ;
  assign \new_[10978]_  = ~\new_[11893]_  | ~\new_[4215]_ ;
  assign \new_[10979]_  = ~\new_[12487]_  | ~\new_[4260]_ ;
  assign \new_[10980]_  = ~\new_[11893]_  | ~\new_[4216]_ ;
  assign \new_[10981]_  = ~\new_[12487]_  | ~\pci_ad_o[29] ;
  assign \new_[10982]_  = ~\new_[12485]_  | ~\new_[4265]_ ;
  assign \new_[10983]_  = ~\new_[12487]_  | ~\new_[4217]_ ;
  assign \new_[10984]_  = ~\new_[12484]_  | ~\new_[4181]_ ;
  assign \new_[10985]_  = ~\new_[12484]_  | ~\new_[4182]_ ;
  assign \new_[10986]_  = ~\new_[12487]_  | ~\new_[4456]_ ;
  assign \new_[10987]_  = ~\new_[12487]_  | ~\new_[4268]_ ;
  assign \new_[10988]_  = ~\new_[12487]_  | ~\new_[4183]_ ;
  assign \new_[10989]_  = ~\new_[12484]_  | ~\new_[4184]_ ;
  assign \new_[10990]_  = ~\new_[12484]_  | ~\new_[4185]_ ;
  assign \new_[10991]_  = ~\new_[12484]_  | ~\new_[4186]_ ;
  assign \new_[10992]_  = ~\new_[12487]_  | ~\new_[4261]_ ;
  assign \new_[10993]_  = ~\new_[12487]_  | ~\new_[4187]_ ;
  assign \new_[10994]_  = ~\new_[12487]_  | ~\new_[4188]_ ;
  assign \new_[10995]_  = ~\new_[12487]_  | ~\new_[4189]_ ;
  assign \new_[10996]_  = ~\new_[12487]_  | ~\new_[4190]_ ;
  assign \new_[10997]_  = ~\new_[11893]_  | ~\new_[4191]_ ;
  assign \new_[10998]_  = ~\new_[12487]_  | ~\new_[4218]_ ;
  assign \new_[10999]_  = ~\new_[12487]_  | ~\pci_ad_o[18] ;
  assign \new_[11000]_  = ~\new_[12487]_  | ~\pci_ad_o[19] ;
  assign \new_[11001]_  = ~\new_[12485]_  | ~\pci_ad_o[25] ;
  assign \new_[11002]_  = ~\new_[12487]_  | ~\pci_ad_o[27] ;
  assign \new_[11003]_  = ~\new_[12487]_  | ~\pci_ad_o[28] ;
  assign \new_[11004]_  = ~\new_[12487]_  | ~\pci_ad_o[7] ;
  assign \new_[11005]_  = ~\new_[12485]_  | ~\pci_ad_o[9] ;
  assign \new_[11006]_  = ~\new_[12487]_  | ~\pci_ad_o[10] ;
  assign \new_[11007]_  = ~\new_[12485]_  | ~\new_[4345]_ ;
  assign \new_[11008]_  = ~\new_[12485]_  | ~\new_[4226]_ ;
  assign \new_[11009]_  = ~\new_[11893]_  | ~\new_[4228]_ ;
  assign \new_[11010]_  = ~\new_[11893]_  | ~\new_[4229]_ ;
  assign \new_[11011]_  = ~\new_[12484]_  | ~\new_[4210]_ ;
  assign \new_[11012]_  = ~\new_[12485]_  | ~\new_[4211]_ ;
  assign \new_[11013]_  = ~\new_[12487]_  | ~\pci_ad_o[16] ;
  assign \new_[11014]_  = ~\new_[12487]_  | ~\new_[4180]_ ;
  assign n9125 = ~\new_[11883]_  | (~\new_[13298]_  & ~\new_[16418]_ );
  assign \new_[11016]_  = ~\new_[11885]_  | (~\new_[16612]_  & ~\new_[16577]_ );
  assign n9200 = \new_[20500]_  ? \new_[12189]_  : \new_[15894]_ ;
  assign \new_[11018]_  = ~\new_[16400]_  | ~\new_[20525]_  | ~\new_[12542]_  | ~\new_[20397]_ ;
  assign n9205 = \new_[19872]_  ? \new_[12189]_  : \new_[16951]_ ;
  assign n9220 = \new_[20514]_  ? \new_[12338]_  : \new_[14291]_ ;
  assign n9225 = \new_[20512]_  ? \new_[12338]_  : \new_[15355]_ ;
  assign n9215 = \new_[17558]_  ? \new_[12338]_  : \new_[14971]_ ;
  assign n9210 = \new_[17592]_  ? \new_[12338]_  : \new_[14950]_ ;
  assign n9230 = \new_[10386]_  ? \new_[12338]_  : \new_[16102]_ ;
  assign n9120 = \new_[17279]_  ? \new_[12338]_  : \new_[15633]_ ;
  assign \new_[11026]_  = ~\new_[11273]_  | ~\new_[9991]_ ;
  assign \new_[11027]_  = ~\new_[11273]_  | ~\new_[9992]_ ;
  assign \new_[11028]_  = ~\new_[11273]_  | ~\new_[9986]_ ;
  assign \new_[11029]_  = \\configuration_pci_ta1_reg[13] ;
  assign n9360 = ~\new_[11841]_  | (~\new_[15069]_  & ~\new_[12575]_ );
  assign \new_[11031]_  = \\configuration_pci_ta1_reg[15] ;
  assign n9235 = ~\new_[11208]_ ;
  assign n9090 = ~\new_[11209]_ ;
  assign n9240 = ~\new_[11210]_ ;
  assign n9245 = ~\new_[11212]_ ;
  assign \new_[11036]_  = \\configuration_pci_ta1_reg[12] ;
  assign n9305 = ~\new_[11213]_ ;
  assign n9250 = ~\new_[11214]_ ;
  assign n9255 = ~\new_[11216]_ ;
  assign n9260 = ~\new_[11218]_ ;
  assign n9265 = ~\new_[11220]_ ;
  assign n9270 = ~\new_[11221]_ ;
  assign n9325 = ~\new_[11233]_ ;
  assign n9280 = ~\new_[11235]_ ;
  assign n9285 = ~\new_[11238]_ ;
  assign \new_[11046]_  = \\configuration_pci_ta1_reg[8] ;
  assign \new_[11047]_  = \\configuration_pci_ta1_reg[9] ;
  assign n9080 = ~\new_[11244]_ ;
  assign n9290 = ~\new_[11245]_ ;
  assign n9275 = ~\new_[11246]_ ;
  assign n9320 = ~\new_[11247]_ ;
  assign n9300 = ~\new_[11248]_ ;
  assign n9295 = ~\new_[11249]_ ;
  assign n9330 = ~\new_[11250]_ ;
  assign n9310 = ~\new_[11251]_ ;
  assign n9510 = ~\new_[11252]_ ;
  assign n9515 = ~\new_[11253]_ ;
  assign n9315 = ~\new_[11254]_ ;
  assign n9505 = ~\new_[11255]_ ;
  assign n9335 = ~\new_[11256]_ ;
  assign n9500 = ~\new_[11257]_ ;
  assign n9340 = ~\new_[11258]_ ;
  assign n9345 = ~\new_[11259]_ ;
  assign n9355 = ~\new_[11260]_ ;
  assign n9350 = ~\new_[11261]_ ;
  assign n9495 = ~\new_[11262]_ ;
  assign \new_[11067]_  = \\configuration_pci_ta1_reg[27] ;
  assign \new_[11068]_  = \\configuration_pci_ta1_reg[26] ;
  assign \new_[11069]_  = \\configuration_pci_ta1_reg[25] ;
  assign \new_[11070]_  = \\configuration_pci_ta1_reg[22] ;
  assign \new_[11071]_  = \\configuration_pci_ta1_reg[19] ;
  assign \new_[11072]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][32] ;
  assign n9720 = \new_[15093]_  ? \new_[12575]_  : \new_[14895]_ ;
  assign \new_[11074]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][32] ;
  assign \new_[11075]_  = wishbone_slave_unit_pci_initiator_if_posted_write_req_reg;
  assign pci_frame_oe_o = pci_io_mux_frame_iob_en_out_reg;
  assign \new_[11077]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[27] ;
  assign \new_[11078]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[17] ;
  assign \new_[11079]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[19] ;
  assign \new_[11080]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[20] ;
  assign \new_[11081]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[22] ;
  assign \new_[11082]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[23] ;
  assign \new_[11083]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[24] ;
  assign \new_[11084]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[28] ;
  assign \new_[11085]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[29] ;
  assign \new_[11086]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[2] ;
  assign \new_[11087]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[31] ;
  assign \new_[11088]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[3] ;
  assign \new_[11089]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[4] ;
  assign \new_[11090]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[6] ;
  assign \new_[11091]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[8] ;
  assign \new_[11092]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[16] ;
  assign \new_[11093]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[14] ;
  assign \new_[11094]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[0] ;
  assign \new_[11095]_  = output_backup_cbe_en_out_reg;
  assign \new_[11096]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][32] ;
  assign \new_[11097]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][32] ;
  assign \new_[11098]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][32] ;
  assign \new_[11099]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][32] ;
  assign \new_[11100]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][36] ;
  assign \new_[11101]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][32] ;
  assign \new_[11102]_  = ~n17085 & (~\new_[13778]_  | ~\new_[20129]_ );
  assign \new_[11103]_  = ~n16920 & (~\new_[14568]_  | ~\new_[20129]_ );
  assign \new_[11104]_  = ~\new_[13123]_  | ~\new_[17002]_ ;
  assign \new_[11105]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[13] ;
  assign \new_[11106]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[15] ;
  assign \new_[11107]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[9] ;
  assign \new_[11108]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[5] ;
  assign \new_[11109]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[7] ;
  assign \new_[11110]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][36] ;
  assign \new_[11111]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[26] ;
  assign \new_[11112]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[30] ;
  assign \new_[11113]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[18] ;
  assign \new_[11114]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[21] ;
  assign \new_[11115]_  = (~\new_[16497]_  | ~\new_[12545]_ ) & (~\new_[16788]_  | ~\new_[19909]_ );
  assign \new_[11116]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[1] ;
  assign \new_[11117]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[12] ;
  assign \new_[11118]_  = ~\new_[14229]_  | ~\new_[10066]_ ;
  assign \new_[11119]_  = ~\new_[14229]_  | ~\new_[10069]_ ;
  assign \new_[11120]_  = ~\new_[14229]_  | ~\new_[10068]_ ;
  assign \new_[11121]_  = ~\new_[14229]_  | ~\new_[10263]_ ;
  assign \new_[11122]_  = ~\new_[14229]_  | ~n17350;
  assign \new_[11123]_  = ~\new_[17033]_  | ~\new_[20129]_  | ~\new_[15271]_ ;
  assign \new_[11124]_  = ~\new_[17033]_  | ~\new_[20129]_  | ~\new_[15696]_ ;
  assign \new_[11125]_  = ~\new_[14229]_  | ~n16995;
  assign \new_[11126]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[25] ;
  assign \new_[11127]_  = ~\new_[14229]_  | ~n17500;
  assign \new_[11128]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[11] ;
  assign \new_[11129]_  = ~\new_[14229]_  | ~n17335;
  assign \new_[11130]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[0] ;
  assign \new_[11131]_  = ~\\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[10] ;
  assign \new_[11132]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][36] ;
  assign \new_[11133]_  = \\wishbone_slave_unit_pci_initiator_if_be_out_reg[1] ;
  assign \new_[11134]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][32] ;
  assign \new_[11135]_  = \new_[12238]_  | \new_[17258]_ ;
  assign \new_[11136]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][36] ;
  assign \new_[11137]_  = ~n9175;
  assign \new_[11138]_  = ~\new_[13697]_  | ~\new_[20525]_  | ~\new_[12471]_  | ~\new_[12542]_ ;
  assign \new_[11139]_  = \new_[12389]_  | \new_[16655]_ ;
  assign \new_[11140]_  = \new_[12390]_  | \new_[16655]_ ;
  assign \new_[11141]_  = \new_[12391]_  | \new_[16658]_ ;
  assign \new_[11142]_  = \new_[12392]_  | \new_[16655]_ ;
  assign \new_[11143]_  = \new_[12393]_  | \new_[16658]_ ;
  assign n9545 = ~\new_[12400]_  | (~\new_[14221]_  & ~\new_[10496]_ );
  assign \new_[11145]_  = ~\new_[17012]_  & (~\new_[13152]_  | ~\new_[15572]_ );
  assign n9550 = ~\new_[13144]_  | (~\new_[13804]_  & ~\new_[15625]_ );
  assign n9770 = \new_[16161]_  ? \new_[13804]_  : \new_[10824]_ ;
  assign n9730 = \new_[16215]_  ? \new_[13804]_  : \new_[10759]_ ;
  assign n9765 = \new_[13152]_  ? \new_[13572]_  : \new_[10823]_ ;
  assign \new_[11150]_  = ~\new_[20387]_  | ~\new_[16687]_ ;
  assign \new_[11151]_  = ~\new_[12487]_  | ~\pci_ad_o[5] ;
  assign \new_[11152]_  = ~\new_[12487]_  | ~\pci_ad_o[4] ;
  assign \new_[11153]_  = ~\new_[12487]_  | ~\pci_ad_o[2] ;
  assign \new_[11154]_  = \new_[17797]_  & \new_[12467]_ ;
  assign \new_[11155]_  = ~\new_[12485]_  | ~\new_[4192]_ ;
  assign \new_[11156]_  = ~\new_[12485]_  | ~\pci_ad_o[26] ;
  assign \new_[11157]_  = ~\new_[12487]_  | ~\pci_ad_o[23] ;
  assign \new_[11158]_  = ~\new_[12485]_  | ~\pci_ad_o[20] ;
  assign \new_[11159]_  = ~\new_[12485]_  | ~\pci_ad_o[0] ;
  assign \new_[11160]_  = ~\new_[12487]_  | ~\pci_ad_o[13] ;
  assign \new_[11161]_  = ~\new_[12487]_  | ~\pci_ad_o[14] ;
  assign \new_[11162]_  = ~\new_[12487]_  | ~\pci_ad_o[15] ;
  assign \new_[11163]_  = ~\new_[12487]_  | ~\pci_ad_o[17] ;
  assign \new_[11164]_  = ~\new_[12487]_  | ~\pci_ad_o[1] ;
  assign \new_[11165]_  = ~\new_[12487]_  | ~\pci_ad_o[21] ;
  assign \new_[11166]_  = ~\new_[12487]_  | ~\pci_ad_o[22] ;
  assign \new_[11167]_  = ~\new_[12487]_  | ~\pci_ad_o[24] ;
  assign \new_[11168]_  = ~\new_[12487]_  | ~\pci_ad_o[30] ;
  assign \new_[11169]_  = ~\new_[12487]_  | ~\pci_ad_o[3] ;
  assign \new_[11170]_  = ~\new_[12487]_  | ~\pci_ad_o[6] ;
  assign \new_[11171]_  = ~\new_[12485]_  | ~\pci_ad_o[8] ;
  assign \new_[11172]_  = ~\new_[12487]_  | ~\pci_ad_o[11] ;
  assign \new_[11173]_  = \new_[20387]_  | \new_[16609]_ ;
  assign n9630 = \new_[11867]_ ;
  assign \new_[11175]_  = ~\new_[11867]_ ;
  assign \new_[11176]_  = ~\new_[12485]_  | ~\pci_ad_o[12] ;
  assign \new_[11177]_  = ~\new_[15478]_  | ~\new_[15685]_  | ~\new_[12474]_  | ~\new_[15747]_ ;
  assign \new_[11178]_  = \new_[12472]_  | \new_[16658]_ ;
  assign n9555 = ~\new_[12439]_  | (~\new_[13820]_  & ~\new_[16118]_ );
  assign n9560 = ~\new_[12440]_  | (~\new_[13820]_  & ~\new_[16126]_ );
  assign n9565 = ~\new_[12441]_  | (~\new_[13820]_  & ~\new_[16116]_ );
  assign n9745 = ~\new_[12443]_  | (~\new_[13820]_  & ~\new_[16111]_ );
  assign n9570 = ~\new_[12442]_  | (~\new_[13820]_  & ~\new_[16124]_ );
  assign n9575 = ~\new_[12444]_  | (~\new_[13820]_  & ~\new_[16117]_ );
  assign n9755 = ~\new_[12445]_  | (~\new_[13820]_  & ~\new_[16146]_ );
  assign n9580 = ~\new_[12446]_  | (~\new_[13820]_  & ~\new_[16110]_ );
  assign n9585 = ~\new_[12447]_  | (~\new_[13820]_  & ~\new_[15933]_ );
  assign n9590 = ~\new_[12449]_  | (~\new_[13820]_  & ~\new_[16152]_ );
  assign n9750 = ~\new_[12450]_  | (~\new_[13820]_  & ~\new_[16151]_ );
  assign n9595 = ~\new_[12451]_  | (~\new_[13820]_  & ~\new_[16424]_ );
  assign n9600 = ~\new_[12452]_  | (~\new_[13820]_  & ~\new_[16147]_ );
  assign n9725 = ~\new_[12453]_  | (~\new_[13820]_  & ~\new_[16418]_ );
  assign n9740 = ~\new_[12455]_  | (~\new_[13820]_  & ~\new_[16431]_ );
  assign n9735 = ~\new_[12454]_  | (~\new_[13820]_  & ~\new_[16677]_ );
  assign n9605 = ~\new_[12456]_  | (~\new_[13820]_  & ~\new_[16425]_ );
  assign n9535 = ~\new_[12457]_  | (~\new_[13820]_  & ~\new_[16159]_ );
  assign n9610 = ~\new_[12458]_  | (~\new_[13820]_  & ~\new_[16160]_ );
  assign n9615 = ~\new_[12459]_  | (~\new_[13820]_  & ~\new_[16419]_ );
  assign n9620 = ~\new_[12460]_  | (~\new_[13820]_  & ~\new_[16141]_ );
  assign n9540 = ~\new_[12461]_  | (~\new_[13820]_  & ~\new_[16427]_ );
  assign n9625 = ~\new_[12462]_  | (~\new_[13820]_  & ~\new_[16119]_ );
  assign n9760 = ~\new_[12463]_  | (~\new_[13820]_  & ~\new_[16109]_ );
  assign \new_[11203]_  = ~\new_[12041]_  | ~\new_[10062]_ ;
  assign \new_[11204]_  = ~\new_[12041]_  | ~\new_[10063]_ ;
  assign \new_[11205]_  = ~\new_[12041]_  | ~\new_[10064]_ ;
  assign \new_[11206]_  = ~\new_[12002]_  & ~\new_[14246]_ ;
  assign n9700 = ~\new_[11900]_ ;
  assign \new_[11208]_  = (~\new_[12569]_  | ~\new_[10387]_ ) & (~\new_[13717]_  | ~\new_[16632]_ );
  assign \new_[11209]_  = (~\new_[12569]_  | ~\new_[10358]_ ) & (~\new_[13717]_  | ~\new_[16635]_ );
  assign \new_[11210]_  = (~\new_[12569]_  | ~\new_[10388]_ ) & (~\new_[13717]_  | ~\new_[16633]_ );
  assign n9710 = ~\new_[11902]_ ;
  assign \new_[11212]_  = (~\new_[12569]_  | ~\new_[10389]_ ) & (~\new_[13717]_  | ~\new_[16457]_ );
  assign \new_[11213]_  = (~\new_[12566]_  | ~\new_[10401]_ ) & (~\new_[20121]_  | ~\new_[16423]_ );
  assign \new_[11214]_  = (~\new_[12569]_  | ~\new_[10390]_ ) & (~\new_[13717]_  | ~\new_[16458]_ );
  assign n9780 = ~\new_[11903]_ ;
  assign \new_[11216]_  = (~\new_[12569]_  | ~\new_[10391]_ ) & (~\new_[13717]_  | ~\new_[16631]_ );
  assign n9680 = ~\new_[11904]_ ;
  assign \new_[11218]_  = (~\new_[12569]_  | ~\new_[10392]_ ) & (~\new_[13717]_  | ~\new_[16636]_ );
  assign n9775 = ~\new_[11905]_ ;
  assign \new_[11220]_  = (~\new_[12569]_  | ~\new_[10393]_ ) & (~\new_[13717]_  | ~\new_[16634]_ );
  assign \new_[11221]_  = (~\new_[12568]_  | ~\new_[10394]_ ) & (~\new_[13717]_  | ~\new_[15931]_ );
  assign n9640 = ~\new_[11906]_ ;
  assign n9650 = ~\new_[11908]_ ;
  assign n9645 = ~\new_[11909]_ ;
  assign n9655 = ~\new_[11911]_ ;
  assign n9675 = ~\new_[11912]_ ;
  assign n9525 = ~\new_[11913]_ ;
  assign n9520 = ~\new_[11914]_ ;
  assign n9665 = ~\new_[11916]_ ;
  assign n9660 = ~\new_[11917]_ ;
  assign n9670 = ~\new_[11918]_ ;
  assign n9635 = ~\new_[11923]_ ;
  assign \new_[11233]_  = (~\new_[12565]_  | ~\new_[10405]_ ) & (~\new_[20121]_  | ~\new_[16634]_ );
  assign n9685 = ~\new_[11927]_ ;
  assign \new_[11235]_  = (~\new_[12568]_  | ~\new_[10396]_ ) & (~\new_[13717]_  | ~\new_[15801]_ );
  assign n9530 = ~\new_[11931]_ ;
  assign n9690 = ~\new_[11936]_ ;
  assign \new_[11238]_  = (~\new_[12568]_  | ~n17220) & (~\new_[13717]_  | ~\new_[15901]_ );
  assign n9695 = ~\new_[11939]_ ;
  assign n9790 = ~\new_[11940]_ ;
  assign n9715 = ~\new_[11944]_ ;
  assign n9705 = ~\new_[11945]_ ;
  assign n9785 = ~\new_[11946]_ ;
  assign \new_[11244]_  = (~\new_[12565]_  | ~\new_[10356]_ ) & (~\new_[20121]_  | ~\new_[16458]_ );
  assign \new_[11245]_  = (~\new_[12565]_  | ~\new_[10398]_ ) & (~\new_[20121]_  | ~\new_[16631]_ );
  assign \new_[11246]_  = (~\new_[12565]_  | ~\new_[10395]_ ) & (~\new_[20121]_  | ~\new_[16636]_ );
  assign \new_[11247]_  = (~\new_[12566]_  | ~\new_[10404]_ ) & (~\new_[20121]_  | ~\new_[16422]_ );
  assign \new_[11248]_  = (~\new_[12568]_  | ~n17280) & (~\new_[16120]_  | ~\new_[13717]_ );
  assign \new_[11249]_  = (~\new_[12566]_  | ~\new_[10399]_ ) & (~\new_[20121]_  | ~\new_[16156]_ );
  assign \new_[11250]_  = (~\new_[12566]_  | ~\new_[10406]_ ) & (~\new_[20121]_  | ~\new_[16429]_ );
  assign \new_[11251]_  = (~\new_[12566]_  | ~\new_[10402]_ ) & (~\new_[20121]_  | ~\new_[16420]_ );
  assign \new_[11252]_  = (~\new_[12566]_  | ~\new_[10485]_ ) & (~\new_[20121]_  | ~\new_[16428]_ );
  assign \new_[11253]_  = (~\new_[12566]_  | ~\new_[10486]_ ) & (~\new_[20121]_  | ~\new_[16417]_ );
  assign \new_[11254]_  = (~\new_[12566]_  | ~\new_[10403]_ ) & (~\new_[20121]_  | ~\new_[16421]_ );
  assign \new_[11255]_  = (~\new_[12567]_  | ~\new_[10484]_ ) & (~\new_[20121]_  | ~\new_[16125]_ );
  assign \new_[11256]_  = (~\new_[12567]_  | ~\new_[10407]_ ) & (~\new_[20121]_  | ~\new_[16155]_ );
  assign \new_[11257]_  = (~\new_[12567]_  | ~\new_[10483]_ ) & (~\new_[20121]_  | ~\new_[16416]_ );
  assign \new_[11258]_  = (~\new_[12567]_  | ~\new_[10408]_ ) & (~\new_[20121]_  | ~\new_[16113]_ );
  assign \new_[11259]_  = (~\new_[12567]_  | ~\new_[10409]_ ) & (~\new_[20121]_  | ~\new_[16114]_ );
  assign \new_[11260]_  = (~\new_[12567]_  | ~\new_[10411]_ ) & (~\new_[20121]_  | ~\new_[16121]_ );
  assign \new_[11261]_  = (~\new_[12567]_  | ~\new_[10410]_ ) & (~\new_[20121]_  | ~\new_[16123]_ );
  assign \new_[11262]_  = (~\new_[12567]_  | ~\new_[10481]_ ) & (~\new_[20121]_  | ~\new_[16112]_ );
  assign \new_[11263]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][6] ;
  assign \new_[11264]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][4] ;
  assign \new_[11265]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][13] ;
  assign \new_[11266]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][3] ;
  assign \new_[11267]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][7] ;
  assign \new_[11268]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][9] ;
  assign \new_[11269]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][0] ;
  assign \new_[11270]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][19] ;
  assign \new_[11271]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][6] ;
  assign \new_[11272]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][15] ;
  assign \new_[11273]_  = \new_[12576]_  | \new_[17258]_ ;
  assign \new_[11274]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][7] ;
  assign \new_[11275]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][16] ;
  assign \new_[11276]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][8] ;
  assign \new_[11277]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][17] ;
  assign \new_[11278]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][7] ;
  assign \new_[11279]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][30] ;
  assign \new_[11280]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][25] ;
  assign \new_[11281]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][0] ;
  assign \new_[11282]_  = \\wishbone_slave_unit_wishbone_slave_img_hit_reg[4] ;
  assign \new_[11283]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][12] ;
  assign \new_[11284]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][3] ;
  assign \new_[11285]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][12] ;
  assign \new_[11286]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][10] ;
  assign \new_[11287]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][36] ;
  assign \new_[11288]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][11] ;
  assign \new_[11289]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][9] ;
  assign \new_[11290]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][2] ;
  assign \new_[11291]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][29] ;
  assign \new_[11292]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][8] ;
  assign \new_[11293]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][7] ;
  assign \new_[11294]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][8] ;
  assign \new_[11295]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][25] ;
  assign \new_[11296]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][23] ;
  assign \new_[11297]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][14] ;
  assign \new_[11298]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][6] ;
  assign \new_[11299]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][16] ;
  assign \new_[11300]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][27] ;
  assign \new_[11301]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][13] ;
  assign \new_[11302]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][28] ;
  assign \new_[11303]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][1] ;
  assign \new_[11304]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][25] ;
  assign \new_[11305]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][26] ;
  assign \new_[11306]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][23] ;
  assign \new_[11307]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][16] ;
  assign \new_[11308]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][16] ;
  assign \new_[11309]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][8] ;
  assign \new_[11310]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][12] ;
  assign \new_[11311]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][10] ;
  assign \new_[11312]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][9] ;
  assign \new_[11313]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][25] ;
  assign \new_[11314]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][31] ;
  assign \new_[11315]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][4] ;
  assign \new_[11316]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][22] ;
  assign \new_[11317]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][18] ;
  assign \new_[11318]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][27] ;
  assign \new_[11319]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][29] ;
  assign \new_[11320]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][21] ;
  assign \new_[11321]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][27] ;
  assign \new_[11322]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][23] ;
  assign \new_[11323]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][1] ;
  assign \new_[11324]_  = ~\\pci_target_unit_del_sync_comp_cycle_count_reg[16] ;
  assign \new_[11325]_  = ~configuration_set_isr_bit2_reg;
  assign \new_[11326]_  = \\wishbone_slave_unit_wishbone_slave_img_hit_reg[2] ;
  assign \new_[11327]_  = \\wishbone_slave_unit_wishbone_slave_img_hit_reg[3] ;
  assign \new_[11328]_  = wishbone_slave_unit_wishbone_slave_wb_conf_hit_reg;
  assign \new_[11329]_  = \\configuration_wb_err_addr_reg[0] ;
  assign \new_[11330]_  = \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6] ;
  assign \new_[11331]_  = \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2] ;
  assign \new_[11332]_  = output_backup_frame_en_out_reg;
  assign \new_[11333]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][0] ;
  assign \new_[11334]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][0] ;
  assign n9805 = ~\new_[12575]_  & (~\new_[15541]_  | ~\new_[15202]_ );
  assign \new_[11336]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][0] ;
  assign \new_[11337]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][0] ;
  assign \new_[11338]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][1] ;
  assign \new_[11339]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][0] ;
  assign \new_[11340]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][0] ;
  assign \pci_cbe_oe_o[3]  = pci_io_mux_cbe_iob3_en_out_reg;
  assign \pci_cbe_oe_o[2]  = pci_io_mux_cbe_iob2_en_out_reg;
  assign \new_[11343]_  = \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3] ;
  assign \new_[11344]_  = \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0] ;
  assign \new_[11345]_  = \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2] ;
  assign \new_[11346]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[3] ;
  assign \new_[11347]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][0] ;
  assign \new_[11348]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][10] ;
  assign \new_[11349]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][12] ;
  assign \new_[11350]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][14] ;
  assign \new_[11351]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][10] ;
  assign \new_[11352]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][16] ;
  assign \new_[11353]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][18] ;
  assign \new_[11354]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][1] ;
  assign \new_[11355]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][21] ;
  assign \new_[11356]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][23] ;
  assign \new_[11357]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][24] ;
  assign \new_[11358]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][25] ;
  assign \new_[11359]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][27] ;
  assign \new_[11360]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][28] ;
  assign \new_[11361]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][29] ;
  assign \new_[11362]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][30] ;
  assign \new_[11363]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][4] ;
  assign \new_[11364]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][6] ;
  assign \new_[11365]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][8] ;
  assign \new_[11366]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][0] ;
  assign \new_[11367]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][11] ;
  assign \new_[11368]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][13] ;
  assign \new_[11369]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][15] ;
  assign \new_[11370]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][17] ;
  assign \new_[11371]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][19] ;
  assign \new_[11372]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][20] ;
  assign \new_[11373]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][22] ;
  assign \new_[11374]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][24] ;
  assign \new_[11375]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][26] ;
  assign \new_[11376]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][28] ;
  assign \new_[11377]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][30] ;
  assign \new_[11378]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][2] ;
  assign \new_[11379]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][3] ;
  assign \new_[11380]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][5] ;
  assign \new_[11381]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][7] ;
  assign \new_[11382]_  = \new_[12570]_  | \new_[13716]_ ;
  assign \new_[11383]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][0] ;
  assign \new_[11384]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][11] ;
  assign \new_[11385]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][13] ;
  assign \new_[11386]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][14] ;
  assign \new_[11387]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][15] ;
  assign \new_[11388]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][17] ;
  assign \new_[11389]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][18] ;
  assign \new_[11390]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][19] ;
  assign \new_[11391]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][20] ;
  assign \new_[11392]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][21] ;
  assign \new_[11393]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][22] ;
  assign \new_[11394]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][24] ;
  assign \new_[11395]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][2] ;
  assign \new_[11396]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][3] ;
  assign \new_[11397]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][5] ;
  assign \new_[11398]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][7] ;
  assign \new_[11399]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][9] ;
  assign \new_[11400]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][0] ;
  assign \new_[11401]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][11] ;
  assign \new_[11402]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][13] ;
  assign \new_[11403]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][15] ;
  assign \new_[11404]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][17] ;
  assign \new_[11405]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][18] ;
  assign \new_[11406]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][19] ;
  assign \new_[11407]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][20] ;
  assign \new_[11408]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][22] ;
  assign \new_[11409]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][24] ;
  assign \new_[11410]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][25] ;
  assign \new_[11411]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][26] ;
  assign \new_[11412]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][28] ;
  assign \new_[11413]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][2] ;
  assign \new_[11414]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][31] ;
  assign \new_[11415]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][3] ;
  assign \new_[11416]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][5] ;
  assign \new_[11417]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][6] ;
  assign \new_[11418]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][7] ;
  assign \new_[11419]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][9] ;
  assign \new_[11420]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][10] ;
  assign \new_[11421]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][12] ;
  assign \new_[11422]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][13] ;
  assign \new_[11423]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][14] ;
  assign \new_[11424]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][16] ;
  assign \new_[11425]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][1] ;
  assign \new_[11426]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][27] ;
  assign \new_[11427]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][31] ;
  assign \new_[11428]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][30] ;
  assign \new_[11429]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][4] ;
  assign \new_[11430]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][6] ;
  assign \new_[11431]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][8] ;
  assign \new_[11432]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][9] ;
  assign \new_[11433]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][0] ;
  assign \new_[11434]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][15] ;
  assign \new_[11435]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][19] ;
  assign \new_[11436]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][20] ;
  assign \new_[11437]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][22] ;
  assign \new_[11438]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][23] ;
  assign \new_[11439]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][24] ;
  assign \new_[11440]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][26] ;
  assign \new_[11441]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][28] ;
  assign \new_[11442]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][30] ;
  assign \new_[11443]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][2] ;
  assign \new_[11444]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][3] ;
  assign \new_[11445]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][5] ;
  assign \new_[11446]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][24] ;
  assign \new_[11447]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][7] ;
  assign \new_[11448]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][9] ;
  assign \new_[11449]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][10] ;
  assign \new_[11450]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][12] ;
  assign \new_[11451]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][14] ;
  assign \new_[11452]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][15] ;
  assign \new_[11453]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][16] ;
  assign \new_[11454]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][18] ;
  assign \new_[11455]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][19] ;
  assign \new_[11456]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][1] ;
  assign \new_[11457]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][21] ;
  assign \new_[11458]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][22] ;
  assign \new_[11459]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][23] ;
  assign \new_[11460]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][25] ;
  assign \new_[11461]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][27] ;
  assign \new_[11462]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][29] ;
  assign \new_[11463]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][2] ;
  assign \new_[11464]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][30] ;
  assign \new_[11465]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][4] ;
  assign \new_[11466]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][6] ;
  assign \new_[11467]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][8] ;
  assign \new_[11468]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][0] ;
  assign \new_[11469]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][11] ;
  assign \new_[11470]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][13] ;
  assign \new_[11471]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][14] ;
  assign \new_[11472]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][15] ;
  assign \new_[11473]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][17] ;
  assign \new_[11474]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][18] ;
  assign \new_[11475]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][19] ;
  assign \new_[11476]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][20] ;
  assign \new_[11477]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][21] ;
  assign \new_[11478]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][22] ;
  assign \new_[11479]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][24] ;
  assign \new_[11480]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][26] ;
  assign \new_[11481]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][28] ;
  assign \new_[11482]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][29] ;
  assign \new_[11483]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][2] ;
  assign \new_[11484]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][23] ;
  assign \new_[11485]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][9] ;
  assign \new_[11486]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][10] ;
  assign \new_[11487]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][12] ;
  assign \new_[11488]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][1] ;
  assign \new_[11489]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][21] ;
  assign \new_[11490]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][17] ;
  assign \new_[11491]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][27] ;
  assign \new_[11492]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][30] ;
  assign \new_[11493]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][4] ;
  assign \new_[11494]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][10] ;
  assign \new_[11495]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][12] ;
  assign \new_[11496]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][14] ;
  assign \new_[11497]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][16] ;
  assign \new_[11498]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][18] ;
  assign \new_[11499]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][19] ;
  assign \new_[11500]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][1] ;
  assign \new_[11501]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][21] ;
  assign \new_[11502]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][23] ;
  assign \new_[11503]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][25] ;
  assign \new_[11504]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][29] ;
  assign \new_[11505]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][4] ;
  assign \new_[11506]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][0] ;
  assign \new_[11507]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][13] ;
  assign \new_[11508]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][24] ;
  assign \new_[11509]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][26] ;
  assign \new_[11510]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][28] ;
  assign \new_[11511]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][29] ;
  assign \new_[11512]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][2] ;
  assign \new_[11513]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][3] ;
  assign \new_[11514]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][5] ;
  assign \new_[11515]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][6] ;
  assign \new_[11516]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][7] ;
  assign \new_[11517]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][9] ;
  assign \new_[11518]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][36] ;
  assign \new_[11519]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][36] ;
  assign \new_[11520]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][36] ;
  assign \new_[11521]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][36] ;
  assign \new_[11522]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][36] ;
  assign \new_[11523]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][14] ;
  assign \new_[11524]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][36] ;
  assign \new_[11525]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][36] ;
  assign \new_[11526]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][36] ;
  assign \new_[11527]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][13] ;
  assign \new_[11528]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][15] ;
  assign \new_[11529]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][19] ;
  assign \new_[11530]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][20] ;
  assign \new_[11531]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][24] ;
  assign \new_[11532]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][28] ;
  assign \new_[11533]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][31] ;
  assign \new_[11534]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][5] ;
  assign \new_[11535]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][9] ;
  assign \new_[11536]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][10] ;
  assign \new_[11537]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][14] ;
  assign \new_[11538]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][1] ;
  assign \new_[11539]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][23] ;
  assign \new_[11540]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][4] ;
  assign \new_[11541]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][27] ;
  assign \new_[11542]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][29] ;
  assign \new_[11543]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][4] ;
  assign \new_[11544]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][6] ;
  assign \new_[11545]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][8] ;
  assign \new_[11546]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][0] ;
  assign \new_[11547]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][19] ;
  assign \new_[11548]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][20] ;
  assign \new_[11549]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][22] ;
  assign \new_[11550]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][2] ;
  assign \new_[11551]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][31] ;
  assign \new_[11552]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][3] ;
  assign \new_[11553]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][5] ;
  assign \new_[11554]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][14] ;
  assign \new_[11555]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][18] ;
  assign \new_[11556]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][1] ;
  assign \new_[11557]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][25] ;
  assign \new_[11558]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][27] ;
  assign \new_[11559]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][29] ;
  assign \new_[11560]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][29] ;
  assign \new_[11561]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][30] ;
  assign \new_[11562]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][36] ;
  assign \new_[11563]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][36] ;
  assign \new_[11564]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][36] ;
  assign \new_[11565]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][10] ;
  assign \new_[11566]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][14] ;
  assign \new_[11567]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][18] ;
  assign \new_[11568]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][1] ;
  assign \new_[11569]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][23] ;
  assign \new_[11570]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][29] ;
  assign \new_[11571]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][36] ;
  assign \new_[11572]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][6] ;
  assign \new_[11573]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][16] ;
  assign \new_[11574]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][18] ;
  assign \new_[11575]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][30] ;
  assign \new_[11576]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][22] ;
  assign \new_[11577]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][21] ;
  assign \new_[11578]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][36] ;
  assign \new_[11579]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][1] ;
  assign \new_[11580]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][1] ;
  assign \new_[11581]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][26] ;
  assign \new_[11582]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][14] ;
  assign \new_[11583]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][27] ;
  assign \new_[11584]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][28] ;
  assign \new_[11585]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][10] ;
  assign \new_[11586]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][12] ;
  assign \new_[11587]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][24] ;
  assign \new_[11588]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][25] ;
  assign \new_[11589]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][0] ;
  assign \new_[11590]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][11] ;
  assign \new_[11591]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][21] ;
  assign \new_[11592]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][10] ;
  assign \new_[11593]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][23] ;
  assign \new_[11594]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][11] ;
  assign \new_[11595]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][16] ;
  assign \new_[11596]_  = ~\new_[10002]_  | ~n16645 | ~\new_[13120]_  | ~\new_[17519]_ ;
  assign \new_[11597]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][17] ;
  assign \new_[11598]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][18] ;
  assign \new_[11599]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][14] ;
  assign \new_[11600]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][12] ;
  assign \new_[11601]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][15] ;
  assign \new_[11602]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][13] ;
  assign \new_[11603]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][3] ;
  assign \new_[11604]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][8] ;
  assign \new_[11605]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][9] ;
  assign \new_[11606]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][14] ;
  assign \new_[11607]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][20] ;
  assign \new_[11608]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][9] ;
  assign \new_[11609]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][22] ;
  assign \new_[11610]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][5] ;
  assign \new_[11611]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][5] ;
  assign \new_[11612]_  = ~\new_[13117]_  | ~\new_[20340]_ ;
  assign \new_[11613]_  = ~\new_[13118]_  | ~\new_[20340]_ ;
  assign \new_[11614]_  = ~\new_[13121]_  | ~\new_[20340]_ ;
  assign n9880 = ~\new_[13122]_  | ~\new_[13571]_ ;
  assign \new_[11616]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][5] ;
  assign \new_[11617]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][7] ;
  assign n9945 = \new_[19690]_  ? \new_[13896]_  : \new_[13597]_ ;
  assign n9885 = \new_[19277]_  ? \new_[13838]_  : \new_[13582]_ ;
  assign n9890 = \new_[19346]_  ? \new_[13839]_  : \new_[13589]_ ;
  assign n9900 = \new_[18815]_  ? \new_[14919]_  : \new_[13595]_ ;
  assign \new_[11622]_  = \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3] ;
  assign n9960 = \new_[17921]_  ? \new_[13838]_  : \new_[13594]_ ;
  assign \new_[11624]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][6] ;
  assign n9910 = \new_[17934]_  ? \new_[13839]_  : \new_[13596]_ ;
  assign n9915 = \new_[20336]_  ? \new_[13902]_  : \new_[13585]_ ;
  assign n9920 = \new_[19671]_  ? \new_[13902]_  : \new_[13593]_ ;
  assign n9925 = \new_[19484]_  ? \new_[13896]_  : \new_[13586]_ ;
  assign n9950 = \new_[17951]_  ? \new_[13908]_  : \new_[13592]_ ;
  assign \new_[11630]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][7] ;
  assign n9955 = \new_[19173]_  ? \new_[13907]_  : \new_[13587]_ ;
  assign n9930 = \new_[19462]_  ? \new_[13908]_  : \new_[13591]_ ;
  assign \new_[11633]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][27] ;
  assign \new_[11634]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][19] ;
  assign n9935 = \new_[18144]_  ? \new_[14920]_  : \new_[13588]_ ;
  assign \new_[11636]_  = ~\new_[13832]_  | ~\new_[12575]_ ;
  assign \new_[11637]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][8] ;
  assign \new_[11638]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][4] ;
  assign n9940 = \new_[19403]_  ? \new_[13900]_  : \new_[13590]_ ;
  assign \new_[11640]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][30] ;
  assign \new_[11641]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][31] ;
  assign n9895 = \new_[17908]_  ? \new_[14920]_  : \new_[13583]_ ;
  assign n9905 = \new_[18448]_  ? \new_[14920]_  : \new_[13584]_ ;
  assign \new_[11644]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][20] ;
  assign \new_[11645]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][1] ;
  assign \new_[11646]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][23] ;
  assign \new_[11647]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][25] ;
  assign \new_[11648]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][21] ;
  assign \new_[11649]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][22] ;
  assign \new_[11650]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][31] ;
  assign \new_[11651]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][3] ;
  assign \new_[11652]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][16] ;
  assign \new_[11653]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][10] ;
  assign \new_[11654]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][11] ;
  assign \new_[11655]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][12] ;
  assign \new_[11656]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][17] ;
  assign \new_[11657]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][24] ;
  assign \new_[11658]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][15] ;
  assign \new_[11659]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][31] ;
  assign \new_[11660]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][2] ;
  assign \new_[11661]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][5] ;
  assign \new_[11662]_  = ~\new_[13127]_  & (~\new_[5011]_  | ~\new_[19906]_ );
  assign \new_[11663]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][3] ;
  assign \new_[11664]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][18] ;
  assign \new_[11665]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][15] ;
  assign \new_[11666]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][17] ;
  assign \new_[11667]_  = ~\new_[15055]_  | ~\new_[20129]_ ;
  assign \new_[11668]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][4] ;
  assign \new_[11669]_  = \new_[14229]_  | \new_[14838]_ ;
  assign \new_[11670]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][1] ;
  assign \new_[11671]_  = \new_[14229]_  | \new_[15550]_ ;
  assign \new_[11672]_  = ~\new_[15397]_  | ~\new_[16608]_  | ~\new_[20129]_  | ~\new_[15893]_ ;
  assign \new_[11673]_  = ~\new_[13123]_ ;
  assign \new_[11674]_  = ~\new_[13123]_ ;
  assign \new_[11675]_  = ~\new_[13123]_ ;
  assign \new_[11676]_  = ~\new_[13123]_ ;
  assign \new_[11677]_  = ~\new_[13123]_ ;
  assign \new_[11678]_  = ~\new_[13123]_ ;
  assign \new_[11679]_  = ~\new_[13123]_ ;
  assign \new_[11680]_  = ~\new_[13123]_ ;
  assign \new_[11681]_  = ~\new_[13123]_ ;
  assign \new_[11682]_  = configuration_wb_err_cs_bit9_reg;
  assign \new_[11683]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][5] ;
  assign \new_[11684]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][23] ;
  assign \new_[11685]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][0] ;
  assign \new_[11686]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][0] ;
  assign \new_[11687]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][17] ;
  assign \new_[11688]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][26] ;
  assign \new_[11689]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][0] ;
  assign \new_[11690]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][1] ;
  assign \new_[11691]_  = \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[0] ;
  assign \new_[11692]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][1] ;
  assign \new_[11693]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][9] ;
  assign \new_[11694]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][36] ;
  assign \new_[11695]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][26] ;
  assign \new_[11696]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][25] ;
  assign \new_[11697]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][11] ;
  assign \new_[11698]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][17] ;
  assign \new_[11699]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][30] ;
  assign \new_[11700]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][7] ;
  assign \new_[11701]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][5] ;
  assign \new_[11702]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][24] ;
  assign \new_[11703]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][28] ;
  assign \new_[11704]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][18] ;
  assign \new_[11705]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][31] ;
  assign \new_[11706]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][26] ;
  assign \new_[11707]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][26] ;
  assign \new_[11708]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][7] ;
  assign \new_[11709]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][19] ;
  assign \new_[11710]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][20] ;
  assign \new_[11711]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][15] ;
  assign \new_[11712]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][2] ;
  assign \new_[11713]_  = \wbm_adr_o[30]  ? \new_[15502]_  : \new_[13607]_ ;
  assign \new_[11714]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][22] ;
  assign \new_[11715]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][28] ;
  assign \new_[11716]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][8] ;
  assign \new_[11717]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][19] ;
  assign \new_[11718]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][16] ;
  assign \new_[11719]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][24] ;
  assign \new_[11720]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][27] ;
  assign \new_[11721]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][3] ;
  assign \new_[11722]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][29] ;
  assign \new_[11723]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][13] ;
  assign \new_[11724]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][14] ;
  assign \new_[11725]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][2] ;
  assign \new_[11726]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][28] ;
  assign \new_[11727]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][20] ;
  assign \new_[11728]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][29] ;
  assign \new_[11729]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][7] ;
  assign \new_[11730]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][6] ;
  assign \new_[11731]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][10] ;
  assign \new_[11732]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][11] ;
  assign \new_[11733]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][20] ;
  assign \new_[11734]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][31] ;
  assign \new_[11735]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][1] ;
  assign \new_[11736]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][17] ;
  assign \new_[11737]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][27] ;
  assign \new_[11738]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][26] ;
  assign \new_[11739]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][26] ;
  assign \new_[11740]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][0] ;
  assign \new_[11741]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][9] ;
  assign \new_[11742]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][28] ;
  assign \new_[11743]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][18] ;
  assign \new_[11744]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][6] ;
  assign \new_[11745]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][20] ;
  assign \new_[11746]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][21] ;
  assign \new_[11747]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][13] ;
  assign \new_[11748]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][22] ;
  assign \new_[11749]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][5] ;
  assign \new_[11750]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][13] ;
  assign \new_[11751]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][3] ;
  assign \new_[11752]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][11] ;
  assign \new_[11753]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][17] ;
  assign \new_[11754]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][11] ;
  assign \new_[11755]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][4] ;
  assign \new_[11756]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[2] ;
  assign \new_[11757]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][18] ;
  assign \new_[11758]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][30] ;
  assign \new_[11759]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][6] ;
  assign \new_[11760]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][1] ;
  assign \new_[11761]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][7] ;
  assign \new_[11762]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][30] ;
  assign \new_[11763]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][13] ;
  assign \new_[11764]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][19] ;
  assign \new_[11765]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][8] ;
  assign \new_[11766]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][15] ;
  assign \new_[11767]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][4] ;
  assign \new_[11768]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][8] ;
  assign \new_[11769]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][17] ;
  assign \new_[11770]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][29] ;
  assign \new_[11771]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][27] ;
  assign \new_[11772]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][31] ;
  assign \new_[11773]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][11] ;
  assign \new_[11774]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][9] ;
  assign \new_[11775]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][31] ;
  assign \new_[11776]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][25] ;
  assign \new_[11777]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][15] ;
  assign \new_[11778]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][23] ;
  assign \new_[11779]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][0] ;
  assign \new_[11780]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][2] ;
  assign \new_[11781]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][31] ;
  assign \new_[11782]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[1] ;
  assign \new_[11783]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][5] ;
  assign \new_[11784]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][3] ;
  assign \new_[11785]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][16] ;
  assign \new_[11786]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][8] ;
  assign \new_[11787]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][10] ;
  assign \new_[11788]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][25] ;
  assign \new_[11789]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][29] ;
  assign \new_[11790]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][0] ;
  assign \new_[11791]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][36] ;
  assign \new_[11792]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][27] ;
  assign \new_[11793]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][31] ;
  assign \new_[11794]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][4] ;
  assign \new_[11795]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][20] ;
  assign \new_[11796]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][28] ;
  assign \new_[11797]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][25] ;
  assign \new_[11798]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][21] ;
  assign \new_[11799]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][3] ;
  assign \new_[11800]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][27] ;
  assign \new_[11801]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][12] ;
  assign \pci_cbe_oe_o[1]  = pci_io_mux_cbe_iob1_en_out_reg;
  assign \pci_cbe_oe_o[0]  = pci_io_mux_cbe_iob0_en_out_reg;
  assign \new_[11804]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][2] ;
  assign \new_[11805]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][29] ;
  assign \new_[11806]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][30] ;
  assign \new_[11807]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][30] ;
  assign \new_[11808]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][30] ;
  assign \new_[11809]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][31] ;
  assign \new_[11810]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][21] ;
  assign \new_[11811]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][2] ;
  assign \new_[11812]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][20] ;
  assign \new_[11813]_  = ~\new_[13131]_  & (~\new_[4972]_  | ~\new_[19906]_ );
  assign \new_[11814]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][25] ;
  assign \new_[11815]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][23] ;
  assign \new_[11816]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][12] ;
  assign \new_[11817]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][24] ;
  assign \new_[11818]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][12] ;
  assign \new_[11819]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][1] ;
  assign \new_[11820]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][21] ;
  assign \new_[11821]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][22] ;
  assign \new_[11822]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][14] ;
  assign \new_[11823]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][16] ;
  assign \new_[11824]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][26] ;
  assign \new_[11825]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][10] ;
  assign \new_[11826]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][13] ;
  assign \new_[11827]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][19] ;
  assign \new_[11828]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][8] ;
  assign \new_[11829]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][17] ;
  assign \new_[11830]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][4] ;
  assign \new_[11831]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][1] ;
  assign \new_[11832]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][6] ;
  assign \new_[11833]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][1] ;
  assign \new_[11834]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][15] ;
  assign \new_[11835]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][1] ;
  assign \new_[11836]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][16] ;
  assign \new_[11837]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][9] ;
  assign \new_[11838]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][11] ;
  assign \new_[11839]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][0] ;
  assign \new_[11840]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][36] ;
  assign \new_[11841]_  = ~\new_[12575]_  | ~\new_[20434]_ ;
  assign \new_[11842]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][31] ;
  assign \new_[11843]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][6] ;
  assign \new_[11844]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][7] ;
  assign \new_[11845]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][28] ;
  assign \new_[11846]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][26] ;
  assign \new_[11847]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][8] ;
  assign \new_[11848]_  = ~\new_[14837]_  | ~\new_[13674]_  | ~\new_[12547]_  | ~\new_[15529]_ ;
  assign \new_[11849]_  = ~\new_[19012]_  | ~\new_[16098]_  | ~\new_[13138]_  | ~\new_[17149]_ ;
  assign \new_[11850]_  = ~\new_[16920]_  | ~\new_[16921]_  | ~\new_[13136]_  | ~\new_[15029]_ ;
  assign \new_[11851]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][5] ;
  assign \new_[11852]_  = ~\new_[16098]_  | ~\new_[13146]_  | ~\new_[17149]_ ;
  assign \new_[11853]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][3] ;
  assign \new_[11854]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][2] ;
  assign \new_[11855]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][4] ;
  assign \new_[11856]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][28] ;
  assign \new_[11857]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][22] ;
  assign \new_[11858]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][26] ;
  assign \new_[11859]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][11] ;
  assign \new_[11860]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][24] ;
  assign \new_[11861]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][21] ;
  assign \new_[11862]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][21] ;
  assign n9820 = ~\new_[13643]_  | (~\new_[16484]_  & ~\new_[13436]_ );
  assign \new_[11864]_  = ~\new_[13804]_  | ~\new_[10370]_ ;
  assign \new_[11865]_  = ~\new_[15257]_  | ~\new_[13153]_ ;
  assign n9795 = ~\new_[13804]_  | ~\new_[13814]_ ;
  assign \new_[11867]_  = ~\new_[14925]_  | ~\new_[13157]_  | ~\new_[20216]_ ;
  assign \new_[11868]_  = ~\new_[13804]_  | ~\new_[10367]_ ;
  assign \new_[11869]_  = ~\new_[13804]_  | ~\new_[10366]_ ;
  assign \new_[11870]_  = ~\new_[16069]_  | ~\new_[12543]_  | ~\new_[15358]_ ;
  assign \new_[11871]_  = ~n16895 & (~\new_[13213]_  | ~\new_[17747]_ );
  assign \new_[11872]_  = ~\new_[13845]_  | ~\new_[15740]_  | ~\new_[16383]_  | ~\new_[13600]_ ;
  assign \new_[11873]_  = ~\new_[16434]_  & (~\new_[13599]_  | ~\new_[15318]_ );
  assign \new_[11874]_  = ~\new_[17365]_  | ~\new_[19947]_  | ~\new_[16684]_ ;
  assign \new_[11875]_  = ~\new_[12399]_ ;
  assign \new_[11876]_  = ~\new_[15693]_  | (~\new_[20505]_  & ~\new_[17181]_ );
  assign \new_[11877]_  = (~\new_[13223]_  | ~\new_[17279]_ ) & (~\new_[17038]_  | ~\new_[10371]_ );
  assign \new_[11878]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][11] ;
  assign \new_[11879]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][12] ;
  assign \new_[11880]_  = \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5] ;
  assign \new_[11881]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][12] ;
  assign \new_[11882]_  = \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1] ;
  assign \new_[11883]_  = ~\new_[10365]_  | (~\new_[13298]_  & ~\new_[17476]_ );
  assign \new_[11884]_  = ~\new_[14750]_  | ~\new_[15747]_  | ~\new_[13160]_  | ~\new_[14891]_ ;
  assign \new_[11885]_  = ~\new_[12468]_ ;
  assign \new_[11886]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][22] ;
  assign \new_[11887]_  = ~\new_[13151]_  & ~\new_[15574]_ ;
  assign \new_[11888]_  = ~\new_[13155]_  & (~\new_[20158]_  | ~\new_[17799]_ );
  assign \new_[11889]_  = \new_[12538]_  | \new_[16658]_ ;
  assign \new_[11890]_  = i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg;
  assign \new_[11891]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][18] ;
  assign \new_[11892]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][1] ;
  assign \new_[11893]_  = ~\new_[13635]_ ;
  assign \new_[11894]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][36] ;
  assign n9875 = ~\new_[13125]_  | (~\new_[19308]_  & ~\new_[20065]_ );
  assign \new_[11896]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][20] ;
  assign n10015 = ~\new_[12489]_ ;
  assign n9810 = ~\new_[12491]_ ;
  assign \new_[11899]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][23] ;
  assign \new_[11900]_  = (~\new_[13297]_  | ~\new_[10527]_ ) & (~\new_[13841]_  | ~\new_[16121]_ );
  assign \new_[11901]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][13] ;
  assign \new_[11902]_  = (~\new_[13297]_  | ~\new_[10529]_ ) & (~\new_[13841]_  | ~\new_[16123]_ );
  assign \new_[11903]_  = (~\new_[13295]_  | ~\new_[10846]_ ) & (~\new_[20526]_  | ~\new_[16632]_ );
  assign \new_[11904]_  = (~\new_[13296]_  | ~\new_[10523]_ ) & (~\new_[13841]_  | ~\new_[16417]_ );
  assign \new_[11905]_  = (~\new_[13297]_  | ~\new_[10845]_ ) & (~\new_[13841]_  | ~\new_[16416]_ );
  assign \new_[11906]_  = (~\new_[13295]_  | ~\new_[10515]_ ) & (~\new_[20526]_  | ~\new_[16633]_ );
  assign n9995 = ~\new_[12496]_ ;
  assign \new_[11908]_  = (~\new_[13295]_  | ~\new_[10517]_ ) & (~\new_[13841]_  | ~\new_[16457]_ );
  assign \new_[11909]_  = (~\new_[13295]_  | ~\new_[10516]_ ) & (~\new_[13841]_  | ~\new_[16458]_ );
  assign \new_[11910]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][19] ;
  assign \new_[11911]_  = (~\new_[13295]_  | ~\new_[10518]_ ) & (~\new_[13841]_  | ~\new_[16631]_ );
  assign \new_[11912]_  = (~\new_[13295]_  | ~\new_[10522]_ ) & (~\new_[20526]_  | ~\new_[16636]_ );
  assign \new_[11913]_  = (~\new_[13295]_  | ~\new_[10492]_ ) & (~\new_[20526]_  | ~\new_[16634]_ );
  assign \new_[11914]_  = (~\new_[13296]_  | ~\new_[10491]_ ) & (~\new_[20526]_  | ~\new_[16423]_ );
  assign n9800 = ~\new_[12497]_ ;
  assign \new_[11916]_  = (~\new_[13296]_  | ~\new_[10520]_ ) & (~\new_[13841]_  | ~\new_[16156]_ );
  assign \new_[11917]_  = (~\new_[13296]_  | ~\new_[10519]_ ) & (~\new_[13841]_  | ~\new_[16422]_ );
  assign \new_[11918]_  = (~\new_[13296]_  | ~\new_[10521]_ ) & (~\new_[13841]_  | ~\new_[16420]_ );
  assign n9965 = ~\new_[12499]_ ;
  assign n9980 = ~\new_[12500]_ ;
  assign n9970 = ~\new_[12501]_ ;
  assign n9870 = ~\new_[12502]_ ;
  assign \new_[11923]_  = (~\new_[13296]_  | ~\new_[10514]_ ) & (~\new_[13841]_  | ~\new_[16428]_ );
  assign n9815 = ~\new_[12504]_ ;
  assign n9825 = ~\new_[12505]_ ;
  assign n9830 = ~\new_[12506]_ ;
  assign \new_[11927]_  = (~\new_[13296]_  | ~\new_[10524]_ ) & (~\new_[13841]_  | ~\new_[16421]_ );
  assign n9835 = ~\new_[12507]_ ;
  assign n9840 = ~\new_[12510]_ ;
  assign n10010 = ~\new_[12511]_ ;
  assign \new_[11931]_  = (~\new_[13297]_  | ~\new_[10493]_ ) & (~\new_[13841]_  | ~\new_[16125]_ );
  assign n9850 = ~\new_[12512]_ ;
  assign n9845 = ~\new_[12513]_ ;
  assign \new_[11934]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][24] ;
  assign n10005 = ~\new_[12514]_ ;
  assign \new_[11936]_  = (~\new_[13297]_  | ~\new_[10525]_ ) & (~\new_[20526]_  | ~\new_[16155]_ );
  assign n10000 = ~\new_[12516]_ ;
  assign \new_[11938]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][36] ;
  assign \new_[11939]_  = (~\new_[13296]_  | ~\new_[10526]_ ) & (~\new_[20526]_  | ~\new_[16429]_ );
  assign \new_[11940]_  = (~\new_[13297]_  | ~\new_[10848]_ ) & (~\new_[13841]_  | ~\new_[16113]_ );
  assign n9865 = ~\new_[12519]_ ;
  assign n9985 = ~\new_[12520]_ ;
  assign n9990 = ~\new_[12521]_ ;
  assign \new_[11944]_  = (~\new_[13297]_  | ~\new_[10530]_ ) & (~\new_[20526]_  | ~\new_[16114]_ );
  assign \new_[11945]_  = (~\new_[13297]_  | ~\new_[10528]_ ) & (~\new_[13841]_  | ~\new_[16112]_ );
  assign \new_[11946]_  = (~\new_[13295]_  | ~\new_[10847]_ ) & (~\new_[13841]_  | ~\new_[16635]_ );
  assign \new_[11947]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][36] ;
  assign \new_[11948]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][17] ;
  assign \new_[11949]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][15] ;
  assign n9860 = ~\new_[12530]_ ;
  assign n9975 = ~\new_[12531]_ ;
  assign n9855 = ~\new_[12533]_ ;
  assign \new_[11953]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][16] ;
  assign \new_[11954]_  = \\configuration_wb_err_addr_reg[11] ;
  assign \new_[11955]_  = \\configuration_wb_err_data_reg[0] ;
  assign \new_[11956]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][20] ;
  assign \new_[11957]_  = \\configuration_wb_err_cs_bit31_24_reg[30] ;
  assign \new_[11958]_  = \\configuration_wb_err_addr_reg[19] ;
  assign \new_[11959]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][25] ;
  assign \new_[11960]_  = \\configuration_pci_err_data_reg[28] ;
  assign \new_[11961]_  = wishbone_slave_unit_pci_initiator_if_data_source_reg;
  assign \new_[11962]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][9] ;
  assign \new_[11963]_  = \\configuration_wb_err_cs_bit31_24_reg[28] ;
  assign \new_[11964]_  = \\configuration_wb_err_addr_reg[15] ;
  assign \new_[11965]_  = \new_[13692]_  ? \new_[16795]_  : \new_[19062]_ ;
  assign \new_[11966]_  = \new_[13692]_  ? \new_[16794]_  : \new_[19028]_ ;
  assign \new_[11967]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][16] ;
  assign \new_[11968]_  = \new_[13692]_  ? \new_[16783]_  : \new_[19071]_ ;
  assign \new_[11969]_  = \new_[13692]_  ? \new_[16803]_  : \new_[18715]_ ;
  assign \new_[11970]_  = ~\new_[13647]_  & (~\new_[20298]_  | ~\new_[12401]_ );
  assign \new_[11971]_  = \new_[18904]_  ? \new_[16883]_  : \new_[13692]_ ;
  assign \new_[11972]_  = \new_[18732]_  ? \new_[16784]_  : \new_[13692]_ ;
  assign \new_[11973]_  = \new_[19187]_  ? \new_[16984]_  : \new_[13692]_ ;
  assign \new_[11974]_  = ~\new_[12542]_ ;
  assign \new_[11975]_  = \new_[18838]_  ? \new_[16789]_  : \new_[13692]_ ;
  assign \new_[11976]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][4] ;
  assign \new_[11977]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][14] ;
  assign \new_[11978]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][22] ;
  assign \new_[11979]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][4] ;
  assign \new_[11980]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][30] ;
  assign \new_[11981]_  = \\configuration_wb_err_data_reg[6] ;
  assign \new_[11982]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][21] ;
  assign \new_[11983]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][24] ;
  assign \new_[11984]_  = \\configuration_wb_err_data_reg[8] ;
  assign \new_[11985]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][27] ;
  assign \new_[11986]_  = \\configuration_wb_err_data_reg[30] ;
  assign \new_[11987]_  = \\configuration_wb_err_data_reg[4] ;
  assign \new_[11988]_  = \\configuration_wb_err_data_reg[31] ;
  assign \new_[11989]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][15] ;
  assign \new_[11990]_  = \\configuration_wb_err_data_reg[28] ;
  assign \new_[11991]_  = \\configuration_wb_err_data_reg[27] ;
  assign \new_[11992]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][29] ;
  assign \new_[11993]_  = \\configuration_wb_err_data_reg[24] ;
  assign \new_[11994]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][23] ;
  assign \new_[11995]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][22] ;
  assign \new_[11996]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][18] ;
  assign \new_[11997]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][21] ;
  assign \new_[11998]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][21] ;
  assign \new_[11999]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][16] ;
  assign \new_[12000]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][12] ;
  assign \new_[12001]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][35] ;
  assign \new_[12002]_  = ~\new_[13870]_  | ~\new_[14962]_  | ~\new_[15037]_  | ~\new_[15694]_ ;
  assign \new_[12003]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][26] ;
  assign \new_[12004]_  = \\configuration_wb_err_data_reg[20] ;
  assign \new_[12005]_  = wishbone_slave_unit_pci_initiator_if_read_bound_reg;
  assign \new_[12006]_  = configuration_pci_err_cs_bit9_reg;
  assign \new_[12007]_  = configuration_pci_err_cs_bit10_reg;
  assign \new_[12008]_  = \\configuration_pci_err_cs_bit31_24_reg[30] ;
  assign \new_[12009]_  = \\configuration_pci_err_cs_bit31_24_reg[28] ;
  assign \new_[12010]_  = \\configuration_pci_err_cs_bit31_24_reg[29] ;
  assign \new_[12011]_  = \\wishbone_slave_unit_pci_initiator_if_read_count_reg[1] ;
  assign \new_[12012]_  = \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4] ;
  assign \new_[12013]_  = \\configuration_pci_err_addr_reg[0] ;
  assign \new_[12014]_  = \\configuration_pci_err_addr_reg[11] ;
  assign \new_[12015]_  = \\configuration_pci_err_addr_reg[12] ;
  assign \new_[12016]_  = \\configuration_pci_err_addr_reg[15] ;
  assign \new_[12017]_  = \\configuration_pci_err_addr_reg[19] ;
  assign \new_[12018]_  = \\configuration_pci_err_addr_reg[20] ;
  assign \new_[12019]_  = \\configuration_pci_err_addr_reg[22] ;
  assign \new_[12020]_  = \\configuration_pci_err_addr_reg[26] ;
  assign \new_[12021]_  = \\configuration_pci_err_addr_reg[28] ;
  assign \new_[12022]_  = \\configuration_pci_err_addr_reg[2] ;
  assign \new_[12023]_  = \\configuration_pci_err_addr_reg[31] ;
  assign \new_[12024]_  = \\configuration_pci_err_addr_reg[4] ;
  assign \new_[12025]_  = \\configuration_pci_err_addr_reg[6] ;
  assign \new_[12026]_  = \\configuration_pci_err_addr_reg[8] ;
  assign \new_[12027]_  = \\configuration_pci_err_data_reg[0] ;
  assign \new_[12028]_  = \\configuration_pci_err_data_reg[11] ;
  assign \new_[12029]_  = \\configuration_pci_err_data_reg[13] ;
  assign \new_[12030]_  = \\configuration_pci_err_data_reg[15] ;
  assign \new_[12031]_  = \\configuration_pci_err_data_reg[17] ;
  assign \new_[12032]_  = \\configuration_pci_err_data_reg[19] ;
  assign \new_[12033]_  = \\configuration_pci_err_data_reg[21] ;
  assign \new_[12034]_  = \\configuration_pci_err_data_reg[25] ;
  assign \new_[12035]_  = \\configuration_pci_err_data_reg[29] ;
  assign \new_[12036]_  = \\configuration_pci_err_data_reg[31] ;
  assign \new_[12037]_  = \\configuration_pci_err_data_reg[3] ;
  assign \new_[12038]_  = \\configuration_pci_err_data_reg[7] ;
  assign \new_[12039]_  = pci_target_unit_pci_target_sm_same_read_reg_reg;
  assign \new_[12040]_  = \\configuration_wb_err_cs_bit31_24_reg[25] ;
  assign \new_[12041]_  = \new_[13298]_  | \new_[17258]_ ;
  assign \new_[12042]_  = \\configuration_wb_err_cs_bit31_24_reg[31] ;
  assign \new_[12043]_  = \\configuration_wb_err_data_reg[10] ;
  assign \new_[12044]_  = \\configuration_wb_err_data_reg[11] ;
  assign \new_[12045]_  = \\configuration_wb_err_data_reg[12] ;
  assign \new_[12046]_  = \\configuration_wb_err_data_reg[14] ;
  assign \new_[12047]_  = \\configuration_wb_err_data_reg[15] ;
  assign \new_[12048]_  = \\configuration_wb_err_data_reg[16] ;
  assign \new_[12049]_  = \\configuration_wb_err_data_reg[18] ;
  assign \new_[12050]_  = \\configuration_wb_err_data_reg[19] ;
  assign \new_[12051]_  = \\configuration_wb_err_data_reg[1] ;
  assign \new_[12052]_  = \\configuration_wb_err_data_reg[21] ;
  assign \new_[12053]_  = \\configuration_wb_err_data_reg[22] ;
  assign \new_[12054]_  = \\configuration_wb_err_data_reg[23] ;
  assign \new_[12055]_  = \\configuration_wb_err_data_reg[25] ;
  assign \new_[12056]_  = \\configuration_wb_err_data_reg[26] ;
  assign \new_[12057]_  = ~\new_[13299]_  & ~\new_[14244]_ ;
  assign \new_[12058]_  = \\configuration_wb_err_data_reg[29] ;
  assign \new_[12059]_  = \\configuration_wb_err_data_reg[2] ;
  assign \new_[12060]_  = \\configuration_wb_err_data_reg[3] ;
  assign \new_[12061]_  = \\configuration_wb_err_data_reg[5] ;
  assign \new_[12062]_  = \\configuration_wb_err_data_reg[9] ;
  assign \new_[12063]_  = \\configuration_wb_err_data_reg[7] ;
  assign \new_[12064]_  = \\configuration_wb_err_addr_reg[10] ;
  assign \new_[12065]_  = \\configuration_wb_err_addr_reg[12] ;
  assign \new_[12066]_  = \\configuration_wb_err_addr_reg[13] ;
  assign \new_[12067]_  = \\configuration_wb_err_addr_reg[14] ;
  assign \new_[12068]_  = \\configuration_wb_err_addr_reg[16] ;
  assign \new_[12069]_  = \\configuration_wb_err_addr_reg[18] ;
  assign \new_[12070]_  = \\configuration_wb_err_addr_reg[20] ;
  assign \new_[12071]_  = \\configuration_wb_err_addr_reg[22] ;
  assign \new_[12072]_  = \\configuration_wb_err_addr_reg[24] ;
  assign \new_[12073]_  = \\configuration_wb_err_addr_reg[26] ;
  assign \new_[12074]_  = \\configuration_wb_err_addr_reg[28] ;
  assign \new_[12075]_  = \\configuration_wb_err_addr_reg[2] ;
  assign \new_[12076]_  = \\configuration_wb_err_addr_reg[31] ;
  assign \new_[12077]_  = \\configuration_wb_err_addr_reg[4] ;
  assign \new_[12078]_  = \\configuration_wb_err_addr_reg[6] ;
  assign \new_[12079]_  = \\configuration_wb_err_addr_reg[7] ;
  assign \new_[12080]_  = \\configuration_wb_err_addr_reg[8] ;
  assign \new_[12081]_  = ~\\pci_target_unit_fifos_pciw_inTransactionCount_reg[1] ;
  assign \new_[12082]_  = ~\\pci_target_unit_fifos_inGreyCount_reg[0] ;
  assign \new_[12083]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][17] ;
  assign \new_[12084]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][12] ;
  assign \new_[12085]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][11] ;
  assign \new_[12086]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][20] ;
  assign \new_[12087]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][7] ;
  assign \new_[12088]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][24] ;
  assign \new_[12089]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][3] ;
  assign \new_[12090]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][34] ;
  assign \new_[12091]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][33] ;
  assign \new_[12092]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][15] ;
  assign \new_[12093]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][29] ;
  assign \new_[12094]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][11] ;
  assign \new_[12095]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][13] ;
  assign \new_[12096]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][15] ;
  assign \new_[12097]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][17] ;
  assign \new_[12098]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][20] ;
  assign \new_[12099]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][23] ;
  assign \new_[12100]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][25] ;
  assign \new_[12101]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][28] ;
  assign \new_[12102]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][18] ;
  assign \new_[12103]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][30] ;
  assign \new_[12104]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][34] ;
  assign \new_[12105]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][35] ;
  assign \new_[12106]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][5] ;
  assign \new_[12107]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][7] ;
  assign \new_[12108]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][10] ;
  assign \new_[12109]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][12] ;
  assign \new_[12110]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][17] ;
  assign \new_[12111]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][22] ;
  assign \new_[12112]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][24] ;
  assign \new_[12113]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][31] ;
  assign \new_[12114]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][8] ;
  assign \new_[12115]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][16] ;
  assign \new_[12116]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][19] ;
  assign \new_[12117]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][22] ;
  assign \new_[12118]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][26] ;
  assign \new_[12119]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][2] ;
  assign \new_[12120]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][34] ;
  assign \new_[12121]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][33] ;
  assign \new_[12122]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][5] ;
  assign \new_[12123]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][7] ;
  assign \new_[12124]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][9] ;
  assign \new_[12125]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][14] ;
  assign \new_[12126]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][10] ;
  assign \new_[12127]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][17] ;
  assign \new_[12128]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][20] ;
  assign \new_[12129]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][22] ;
  assign \new_[12130]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][24] ;
  assign \new_[12131]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][23] ;
  assign \new_[12132]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][21] ;
  assign \new_[12133]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][25] ;
  assign \new_[12134]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][12] ;
  assign \new_[12135]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][34] ;
  assign \new_[12136]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][5] ;
  assign \new_[12137]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][7] ;
  assign \new_[12138]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][16] ;
  assign \new_[12139]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][23] ;
  assign \new_[12140]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][21] ;
  assign \new_[12141]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][14] ;
  assign \new_[12142]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][11] ;
  assign \new_[12143]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][13] ;
  assign \new_[12144]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][15] ;
  assign \new_[12145]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][17] ;
  assign \new_[12146]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][19] ;
  assign \new_[12147]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][27] ;
  assign \new_[12148]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][2] ;
  assign \new_[12149]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][3] ;
  assign \new_[12150]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][4] ;
  assign \new_[12151]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][6] ;
  assign \new_[12152]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][7] ;
  assign \new_[12153]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][16] ;
  assign \new_[12154]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][20] ;
  assign \new_[12155]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][22] ;
  assign \new_[12156]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][27] ;
  assign \new_[12157]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][29] ;
  assign \new_[12158]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][33] ;
  assign \new_[12159]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][6] ;
  assign \new_[12160]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][8] ;
  assign \new_[12161]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][10] ;
  assign \new_[12162]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][14] ;
  assign \new_[12163]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][9] ;
  assign \new_[12164]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][19] ;
  assign \new_[12165]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][23] ;
  assign \new_[12166]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][28] ;
  assign \new_[12167]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][8] ;
  assign \new_[12168]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][11] ;
  assign \new_[12169]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][21] ;
  assign \new_[12170]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][24] ;
  assign \new_[12171]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][27] ;
  assign \new_[12172]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][2] ;
  assign \new_[12173]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][18] ;
  assign \new_[12174]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][29] ;
  assign \new_[12175]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][35] ;
  assign \new_[12176]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][26] ;
  assign \new_[12177]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][38] ;
  assign \new_[12178]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][38] ;
  assign \new_[12179]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][38] ;
  assign \new_[12180]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][38] ;
  assign \new_[12181]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][13] ;
  assign \new_[12182]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][18] ;
  assign \new_[12183]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][13] ;
  assign \new_[12184]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][25] ;
  assign \new_[12185]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][19] ;
  assign \new_[12186]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][15] ;
  assign n10250 = \new_[16209]_  ? \new_[13718]_  : \new_[11133]_ ;
  assign n10035 = ~n10605;
  assign \new_[12189]_  = (~\new_[13719]_  & ~\new_[20500]_ ) | (~\new_[16599]_  & ~\new_[17062]_ );
  assign \new_[12190]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][20] ;
  assign n10105 = \new_[13727]_  ? \new_[17510]_  : \new_[18149]_ ;
  assign \new_[12192]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][28] ;
  assign n10075 = \new_[13740]_  ? \new_[17510]_  : \new_[18560]_ ;
  assign \new_[12194]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][12] ;
  assign \new_[12195]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][14] ;
  assign \new_[12196]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][9] ;
  assign \new_[12197]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][18] ;
  assign \new_[12198]_  = \\configuration_wb_err_cs_bit31_24_reg[29] ;
  assign \new_[12199]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][33] ;
  assign n10195 = \new_[13731]_  ? \new_[17510]_  : \new_[18770]_ ;
  assign \new_[12201]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][27] ;
  assign \new_[12202]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][6] ;
  assign n10225 = \new_[13729]_  ? \new_[17510]_  : \new_[18389]_ ;
  assign n10110 = \new_[13756]_  ? \new_[17510]_  : \new_[17822]_ ;
  assign \new_[12205]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][35] ;
  assign n10215 = \new_[13738]_  ? \new_[17510]_  : \new_[17887]_ ;
  assign n10065 = \new_[13734]_  ? \new_[17510]_  : \new_[19616]_ ;
  assign n10230 = \new_[13748]_  ? \new_[17510]_  : \new_[18033]_ ;
  assign n10220 = \new_[13736]_  ? \new_[17510]_  : \new_[18073]_ ;
  assign n10165 = \new_[13737]_  ? \new_[17510]_  : \new_[18001]_ ;
  assign n10045 = \new_[13749]_  ? \new_[17510]_  : \new_[19322]_ ;
  assign \new_[12212]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][5] ;
  assign n10210 = \new_[13739]_  ? \new_[17510]_  : \new_[18049]_ ;
  assign n10070 = \new_[13733]_  ? \new_[17510]_  : \new_[18852]_ ;
  assign n10040 = \new_[13728]_  ? \new_[17510]_  : \new_[18187]_ ;
  assign n10115 = \new_[13735]_  ? \new_[17510]_  : \new_[18574]_ ;
  assign n10080 = \new_[13758]_  ? \new_[17510]_  : \new_[19333]_ ;
  assign n10085 = \new_[13730]_  ? \new_[17510]_  : \new_[19711]_ ;
  assign n10200 = \new_[13741]_  ? \new_[17510]_  : \new_[19674]_ ;
  assign n10090 = \new_[13742]_  ? \new_[17510]_  : \new_[19389]_ ;
  assign n10095 = \new_[13743]_  ? \new_[17510]_  : \new_[19738]_ ;
  assign n10100 = \new_[13732]_  ? \new_[17510]_  : \new_[18897]_ ;
  assign \new_[12223]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][6] ;
  assign n10180 = \new_[13745]_  ? \new_[17510]_  : \new_[18555]_ ;
  assign n10050 = \new_[13754]_  ? \new_[17510]_  : \new_[17920]_ ;
  assign n10185 = \new_[13746]_  ? \new_[17510]_  : \new_[19720]_ ;
  assign n10175 = \new_[13753]_  ? \new_[17510]_  : \new_[19835]_ ;
  assign n10170 = \new_[13744]_  ? \new_[17510]_  : \new_[18176]_ ;
  assign n10205 = \new_[13747]_  ? \new_[17510]_  : \new_[19501]_ ;
  assign n10235 = \new_[13751]_  ? \new_[17510]_  : \new_[18396]_ ;
  assign n10240 = \new_[13752]_  ? \new_[17510]_  : \new_[18173]_ ;
  assign n10120 = \new_[13750]_  ? \new_[17510]_  : \new_[18586]_ ;
  assign n10055 = \new_[13755]_  ? \new_[17510]_  : \new_[19544]_ ;
  assign \new_[12234]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][6] ;
  assign \new_[12235]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][3] ;
  assign \new_[12236]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][8] ;
  assign n10060 = \new_[13757]_  ? \new_[17510]_  : \new_[18310]_ ;
  assign \new_[12238]_  = ~\new_[16372]_  | ~\new_[15578]_  | ~\new_[20129]_ ;
  assign n10125 = ~\new_[13571]_  | (~\new_[11094]_  & ~\new_[14878]_ );
  assign n10130 = ~n12765;
  assign \new_[12241]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][23] ;
  assign \new_[12242]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][22] ;
  assign \new_[12243]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][4] ;
  assign \new_[12244]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][9] ;
  assign \new_[12245]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][6] ;
  assign \new_[12246]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][15] ;
  assign \new_[12247]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][30] ;
  assign \new_[12248]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][8] ;
  assign \new_[12249]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][11] ;
  assign \new_[12250]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][13] ;
  assign \new_[12251]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][9] ;
  assign \new_[12252]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][14] ;
  assign \new_[12253]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][19] ;
  assign \new_[12254]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][4] ;
  assign \new_[12255]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][3] ;
  assign \new_[12256]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][33] ;
  assign \new_[12257]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][2] ;
  assign \new_[12258]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][31] ;
  assign \new_[12259]_  = \\configuration_wb_err_data_reg[13] ;
  assign \new_[12260]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][27] ;
  assign \new_[12261]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][29] ;
  assign n10135 = \new_[13765]_  ? \new_[15590]_  : \new_[18429]_ ;
  assign n10020 = \new_[13766]_  ? \new_[15493]_  : \new_[17856]_ ;
  assign n10025 = \new_[13764]_  ? \new_[15492]_  : \new_[18703]_ ;
  assign n10140 = \new_[13767]_  ? \new_[15494]_  : \new_[18606]_ ;
  assign \new_[12266]_  = \\configuration_wb_err_cs_bit31_24_reg[24] ;
  assign \new_[12267]_  = \\configuration_wb_err_cs_bit31_24_reg[27] ;
  assign \new_[12268]_  = \\configuration_wb_err_cs_bit31_24_reg[26] ;
  assign \new_[12269]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][12] ;
  assign \new_[12270]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][3] ;
  assign \new_[12271]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][10] ;
  assign \new_[12272]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][7] ;
  assign \new_[12273]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][4] ;
  assign \new_[12274]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][29] ;
  assign n10155 = \new_[13768]_  ? \new_[15275]_  : \new_[18661]_ ;
  assign n10145 = \new_[13772]_  ? \new_[15494]_  : \new_[19731]_ ;
  assign \new_[12277]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][11] ;
  assign \new_[12278]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][28] ;
  assign n10260 = \new_[13777]_  ? \new_[15495]_  : \new_[19193]_ ;
  assign n10245 = \new_[13773]_  ? \new_[15488]_  : \new_[19306]_ ;
  assign \new_[12281]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][5] ;
  assign \new_[12282]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][16] ;
  assign n10150 = \new_[13769]_  ? \new_[15486]_  : \new_[19751]_ ;
  assign n10190 = \new_[13770]_  ? \new_[15494]_  : \new_[18346]_ ;
  assign n10255 = \new_[13775]_  ? \new_[15488]_  : \new_[17991]_ ;
  assign \new_[12286]_  = (~\new_[9676]_  & ~\new_[17308]_  & ~\new_[20532]_ ) | (~\new_[16360]_  & ~\new_[20039]_  & ~\new_[17752]_ );
  assign \new_[12287]_  = \\configuration_wb_err_data_reg[17] ;
  assign n10160 = \new_[13776]_  ? \new_[15591]_  : \new_[19470]_ ;
  assign \new_[12289]_  = ~\new_[16837]_  | ~\new_[20129]_  | ~\new_[15696]_ ;
  assign \new_[12290]_  = ~\new_[16837]_  | ~\new_[20129]_  | ~\new_[15271]_ ;
  assign \new_[12291]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][4] ;
  assign \new_[12292]_  = ~\new_[13119]_ ;
  assign \new_[12293]_  = ~\new_[13119]_ ;
  assign \new_[12294]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][31] ;
  assign \new_[12295]_  = ~\new_[13121]_ ;
  assign \new_[12296]_  = \\configuration_pci_err_data_reg[2] ;
  assign \new_[12297]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][35] ;
  assign \new_[12298]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][31] ;
  assign \new_[12299]_  = \\configuration_wb_err_addr_reg[1] ;
  assign \new_[12300]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][22] ;
  assign \new_[12301]_  = \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[7] ;
  assign \new_[12302]_  = pci_target_unit_pci_target_if_same_read_reg_reg;
  assign \new_[12303]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][34] ;
  assign \new_[12304]_  = \\configuration_pci_err_data_reg[8] ;
  assign \new_[12305]_  = \\configuration_pci_err_data_reg[30] ;
  assign \new_[12306]_  = \\configuration_pci_err_data_reg[9] ;
  assign \new_[12307]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][13] ;
  assign \new_[12308]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][20] ;
  assign \new_[12309]_  = \\configuration_pci_err_data_reg[5] ;
  assign \new_[12310]_  = \\configuration_pci_err_data_reg[6] ;
  assign \new_[12311]_  = \\configuration_pci_err_data_reg[4] ;
  assign \new_[12312]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][6] ;
  assign \new_[12313]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][2] ;
  assign \new_[12314]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][30] ;
  assign \new_[12315]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][23] ;
  assign \new_[12316]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][4] ;
  assign \new_[12317]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][26] ;
  assign \new_[12318]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][7] ;
  assign \new_[12319]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][24] ;
  assign \new_[12320]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][26] ;
  assign \new_[12321]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][31] ;
  assign \new_[12322]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][29] ;
  assign \new_[12323]_  = \\configuration_pci_err_data_reg[23] ;
  assign \new_[12324]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][26] ;
  assign \new_[12325]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][25] ;
  assign \new_[12326]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][23] ;
  assign \new_[12327]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][5] ;
  assign \new_[12328]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][10] ;
  assign \new_[12329]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][31] ;
  assign \new_[12330]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][2] ;
  assign \new_[12331]_  = \\configuration_wb_err_addr_reg[17] ;
  assign \new_[12332]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][25] ;
  assign \new_[12333]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][9] ;
  assign \new_[12334]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][6] ;
  assign \new_[12335]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][24] ;
  assign \new_[12336]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][8] ;
  assign \new_[12337]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][17] ;
  assign \new_[12338]_  = ~\new_[14955]_  | ~\new_[13848]_  | ~\new_[16589]_  | ~\new_[16678]_ ;
  assign \new_[12339]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][31] ;
  assign \new_[12340]_  = \\configuration_pci_err_data_reg[24] ;
  assign \new_[12341]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][33] ;
  assign \new_[12342]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][9] ;
  assign \new_[12343]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][18] ;
  assign \new_[12344]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][21] ;
  assign \new_[12345]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][19] ;
  assign \new_[12346]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][33] ;
  assign \new_[12347]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][10] ;
  assign \new_[12348]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][15] ;
  assign \new_[12349]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][3] ;
  assign \new_[12350]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][15] ;
  assign \new_[12351]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][14] ;
  assign \new_[12352]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][34] ;
  assign \new_[12353]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][11] ;
  assign \new_[12354]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][12] ;
  assign \new_[12355]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][34] ;
  assign \new_[12356]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][13] ;
  assign \new_[12357]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][8] ;
  assign \new_[12358]_  = \new_[16709]_  ^ \new_[13792]_ ;
  assign \new_[12359]_  = \new_[4174]_  ^ \new_[13793]_ ;
  assign \new_[12360]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][19] ;
  assign \new_[12361]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][25] ;
  assign \new_[12362]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][17] ;
  assign \new_[12363]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][30] ;
  assign \new_[12364]_  = \new_[15429]_  ^ \new_[13797]_ ;
  assign \new_[12365]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][5] ;
  assign \new_[12366]_  = \\configuration_pci_err_data_reg[26] ;
  assign \new_[12367]_  = \\configuration_pci_err_data_reg[27] ;
  assign \new_[12368]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][34] ;
  assign \new_[12369]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][35] ;
  assign \new_[12370]_  = ~\new_[13135]_ ;
  assign \new_[12371]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][28] ;
  assign \new_[12372]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][35] ;
  assign \new_[12373]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][38] ;
  assign \new_[12374]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][28] ;
  assign \new_[12375]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][16] ;
  assign \new_[12376]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][26] ;
  assign \new_[12377]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][27] ;
  assign \new_[12378]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][10] ;
  assign \new_[12379]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][7] ;
  assign \new_[12380]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][8] ;
  assign \new_[12381]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][18] ;
  assign \new_[12382]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][18] ;
  assign \new_[12383]_  = \\configuration_pci_err_addr_reg[7] ;
  assign \new_[12384]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][20] ;
  assign \new_[12385]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][38] ;
  assign \new_[12386]_  = ~\new_[13630]_  | ~\new_[15612]_ ;
  assign \new_[12387]_  = ~\new_[16655]_  & (~\new_[13811]_  | ~\new_[15474]_ );
  assign \new_[12388]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][14] ;
  assign \new_[12389]_  = ~\new_[13623]_  & ~\new_[13843]_ ;
  assign \new_[12390]_  = ~\new_[13624]_  & ~\new_[13849]_ ;
  assign \new_[12391]_  = ~\new_[13625]_  & ~\new_[13844]_ ;
  assign \new_[12392]_  = ~\new_[13626]_  & ~\new_[13852]_ ;
  assign \new_[12393]_  = ~\new_[13627]_  & ~\new_[13846]_ ;
  assign \new_[12394]_  = ~\new_[16658]_  & (~\new_[13683]_  | ~\new_[15293]_ );
  assign \new_[12395]_  = ~\new_[16655]_  & (~\new_[13682]_  | ~\new_[15295]_ );
  assign \new_[12396]_  = ~\new_[16655]_  & (~\new_[13680]_  | ~\new_[15297]_ );
  assign \new_[12397]_  = ~\new_[16655]_  & (~\new_[13677]_  | ~\new_[15316]_ );
  assign \new_[12398]_  = ~\new_[16655]_  & (~\new_[13676]_  | ~\new_[15299]_ );
  assign \new_[12399]_  = ~\new_[14940]_  | (~\new_[13780]_  & ~\new_[15496]_ );
  assign \new_[12400]_  = (~\new_[15843]_  | ~\new_[14221]_ ) & (~\new_[16180]_  | ~\new_[13710]_ );
  assign \new_[12401]_  = \\configuration_pci_err_addr_reg[9] ;
  assign \new_[12402]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][12] ;
  assign \new_[12403]_  = \new_[19498]_  ? \new_[20186]_  : \new_[18515]_ ;
  assign \new_[12404]_  = \\configuration_pci_err_data_reg[18] ;
  assign \new_[12405]_  = \\configuration_pci_err_data_reg[1] ;
  assign \new_[12406]_  = \\configuration_pci_err_data_reg[20] ;
  assign \new_[12407]_  = \\configuration_pci_err_data_reg[22] ;
  assign \new_[12408]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][10] ;
  assign \new_[12409]_  = \\configuration_pci_err_data_reg[14] ;
  assign \new_[12410]_  = \\configuration_pci_err_cs_bit31_24_reg[24] ;
  assign \new_[12411]_  = \\configuration_pci_err_data_reg[16] ;
  assign \new_[12412]_  = \\configuration_pci_err_cs_bit31_24_reg[25] ;
  assign \new_[12413]_  = \\configuration_pci_err_data_reg[10] ;
  assign \new_[12414]_  = \\configuration_pci_err_data_reg[12] ;
  assign \new_[12415]_  = \\configuration_pci_err_cs_bit31_24_reg[26] ;
  assign \new_[12416]_  = \\configuration_pci_err_cs_bit31_24_reg[27] ;
  assign \new_[12417]_  = \\configuration_pci_err_addr_reg[3] ;
  assign \new_[12418]_  = \\configuration_pci_err_addr_reg[10] ;
  assign \new_[12419]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][5] ;
  assign \new_[12420]_  = \\configuration_wb_err_addr_reg[21] ;
  assign \new_[12421]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][38] ;
  assign \new_[12422]_  = \\configuration_pci_err_addr_reg[5] ;
  assign \new_[12423]_  = \\configuration_pci_err_addr_reg[30] ;
  assign \new_[12424]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][11] ;
  assign \new_[12425]_  = \\configuration_pci_err_addr_reg[27] ;
  assign \new_[12426]_  = \\configuration_pci_err_addr_reg[29] ;
  assign \new_[12427]_  = \\configuration_pci_err_addr_reg[25] ;
  assign \new_[12428]_  = \\configuration_pci_err_addr_reg[1] ;
  assign \new_[12429]_  = \\configuration_pci_err_addr_reg[23] ;
  assign \new_[12430]_  = \\configuration_pci_err_addr_reg[24] ;
  assign \new_[12431]_  = \\configuration_pci_err_addr_reg[21] ;
  assign \new_[12432]_  = \\configuration_pci_err_addr_reg[13] ;
  assign \new_[12433]_  = \\configuration_pci_err_addr_reg[18] ;
  assign \new_[12434]_  = \\configuration_pci_err_addr_reg[17] ;
  assign \new_[12435]_  = \\configuration_pci_err_addr_reg[14] ;
  assign \new_[12436]_  = \\configuration_pci_err_addr_reg[16] ;
  assign \new_[12437]_  = \\configuration_pci_err_cs_bit31_24_reg[31] ;
  assign \new_[12438]_  = ~\new_[16655]_  & (~\new_[13726]_  | ~\new_[14943]_ );
  assign \new_[12439]_  = ~\new_[13610]_  | ~\new_[10498]_ ;
  assign \new_[12440]_  = ~\new_[13610]_  | ~\new_[10499]_ ;
  assign \new_[12441]_  = ~\new_[13610]_  | ~\new_[10500]_ ;
  assign \new_[12442]_  = ~\new_[13610]_  | ~\new_[10501]_ ;
  assign \new_[12443]_  = ~\new_[13610]_  | ~\new_[10775]_ ;
  assign \new_[12444]_  = ~\new_[13610]_  | ~\new_[10502]_ ;
  assign \new_[12445]_  = ~\new_[13214]_  | ~\new_[10816]_ ;
  assign \new_[12446]_  = ~\new_[13214]_  | ~\new_[10503]_ ;
  assign \new_[12447]_  = ~\new_[13214]_  | ~\new_[10504]_ ;
  assign \new_[12448]_  = \\wishbone_slave_unit_pci_initiator_if_read_count_reg[0] ;
  assign \new_[12449]_  = ~\new_[13214]_  | ~\new_[10505]_ ;
  assign \new_[12450]_  = ~\new_[13214]_  | ~\new_[10794]_ ;
  assign \new_[12451]_  = ~\new_[13214]_  | ~\new_[10506]_ ;
  assign \new_[12452]_  = ~\new_[13214]_  | ~\new_[10507]_ ;
  assign \new_[12453]_  = ~\new_[13214]_  | ~\new_[10744]_ ;
  assign \new_[12454]_  = ~\new_[13611]_  | ~\new_[10773]_ ;
  assign \new_[12455]_  = ~\new_[13611]_  | ~\new_[10774]_ ;
  assign \new_[12456]_  = ~\new_[13611]_  | ~\new_[10508]_ ;
  assign \new_[12457]_  = ~\new_[13611]_  | ~\new_[10494]_ ;
  assign \new_[12458]_  = ~\new_[13611]_  | ~\new_[10509]_ ;
  assign \new_[12459]_  = ~\new_[13611]_  | ~\new_[10510]_ ;
  assign \new_[12460]_  = ~\new_[13611]_  | ~\new_[10511]_ ;
  assign \new_[12461]_  = ~\new_[13611]_  | ~\new_[10495]_ ;
  assign \new_[12462]_  = ~\new_[13610]_  | ~\new_[10512]_ ;
  assign \new_[12463]_  = ~\new_[13610]_  | ~\new_[10822]_ ;
  assign \new_[12464]_  = \new_[13213]_  | \new_[15010]_ ;
  assign \new_[12465]_  = ~\new_[16655]_  & (~\new_[13706]_  | ~\new_[15516]_ );
  assign \new_[12466]_  = ~\new_[16658]_  & (~\new_[13707]_  | ~\new_[15520]_ );
  assign \new_[12467]_  = \new_[20505]_  & \new_[17467]_ ;
  assign \new_[12468]_  = \new_[20505]_  & \new_[16904]_ ;
  assign \new_[12469]_  = ~\new_[15887]_  | ~\new_[20397]_ ;
  assign \new_[12470]_  = ~\new_[13153]_ ;
  assign \new_[12471]_  = ~\new_[19958]_ ;
  assign \new_[12472]_  = ~\new_[13649]_  & ~\new_[13847]_ ;
  assign \new_[12473]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][3] ;
  assign \new_[12474]_  = ~\new_[13212]_  & (~\new_[20158]_  | ~\new_[17686]_ );
  assign \new_[12475]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][25] ;
  assign \new_[12476]_  = ~\new_[13646]_  & ~\new_[15574]_ ;
  assign \new_[12477]_  = ~\new_[13645]_  & ~\new_[15574]_ ;
  assign \new_[12478]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][33] ;
  assign \new_[12479]_  = ~\new_[13644]_  & ~\new_[15574]_ ;
  assign n10030 = ~\new_[20186]_  | (~\new_[13779]_  & ~\new_[20151]_ );
  assign \new_[12481]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][31] ;
  assign \new_[12482]_  = ~\new_[16074]_  | (~\new_[13696]_  & ~\new_[13817]_ );
  assign \new_[12483]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][2] ;
  assign \new_[12484]_  = ~\new_[13635]_ ;
  assign \new_[12485]_  = ~\new_[13635]_ ;
  assign \new_[12486]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][24] ;
  assign \new_[12487]_  = ~\new_[13635]_ ;
  assign \new_[12488]_  = ~\new_[13635]_ ;
  assign \new_[12489]_  = (~\new_[13695]_  | ~\new_[11071]_ ) & (~\new_[19920]_  | ~\new_[16429]_ );
  assign \new_[12490]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][13] ;
  assign \new_[12491]_  = (~\new_[13693]_  | ~\new_[10857]_ ) & (~\new_[19920]_  | ~\new_[16121]_ );
  assign \new_[12492]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][21] ;
  assign \new_[12493]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][26] ;
  assign \new_[12494]_  = \\configuration_wb_err_addr_reg[9] ;
  assign \new_[12495]_  = \\configuration_wb_err_addr_reg[5] ;
  assign \new_[12496]_  = (~\new_[13693]_  | ~\new_[11067]_ ) & (~\new_[19920]_  | ~\new_[16113]_ );
  assign \new_[12497]_  = (~\new_[13694]_  | ~\new_[10854]_ ) & (~\new_[19920]_  | ~\new_[16633]_ );
  assign \new_[12498]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][30] ;
  assign \new_[12499]_  = (~\new_[13694]_  | ~\new_[10972]_ ) & (~\new_[19920]_  | ~\new_[16457]_ );
  assign \new_[12500]_  = (~\new_[13694]_  | ~\new_[11036]_ ) & (~\new_[19920]_  | ~\new_[16458]_ );
  assign \new_[12501]_  = (~\new_[13694]_  | ~\new_[11029]_ ) & (~\new_[19920]_  | ~\new_[16631]_ );
  assign \new_[12502]_  = (~\new_[13694]_  | ~\new_[10869]_ ) & (~\new_[19920]_  | ~\new_[16636]_ );
  assign \new_[12503]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][30] ;
  assign \new_[12504]_  = (~\new_[13695]_  | ~\new_[10858]_ ) & (~\new_[19920]_  | ~\new_[16423]_ );
  assign \new_[12505]_  = (~\new_[13695]_  | ~\new_[10860]_ ) & (~\new_[19920]_  | ~\new_[16156]_ );
  assign \new_[12506]_  = (~\new_[13695]_  | ~\new_[10861]_ ) & (~\new_[19920]_  | ~\new_[16422]_ );
  assign \new_[12507]_  = (~\new_[13695]_  | ~\new_[10862]_ ) & (~\new_[19920]_  | ~\new_[16420]_ );
  assign \new_[12508]_  = \\configuration_wb_err_addr_reg[3] ;
  assign \new_[12509]_  = \\configuration_wb_err_addr_reg[23] ;
  assign \new_[12510]_  = (~\new_[13695]_  | ~\new_[10863]_ ) & (~\new_[19920]_  | ~\new_[16428]_ );
  assign \new_[12511]_  = (~\new_[13695]_  | ~\new_[11070]_ ) & (~\new_[19920]_  | ~\new_[16417]_ );
  assign \new_[12512]_  = (~\new_[13695]_  | ~\new_[10865]_ ) & (~\new_[19920]_  | ~\new_[16421]_ );
  assign \new_[12513]_  = (~\new_[13693]_  | ~\new_[10864]_ ) & (~\new_[19920]_  | ~\new_[16125]_ );
  assign \new_[12514]_  = (~\new_[13693]_  | ~\new_[11069]_ ) & (~\new_[19920]_  | ~\new_[16155]_ );
  assign \new_[12515]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][27] ;
  assign \new_[12516]_  = (~\new_[13693]_  | ~\new_[11068]_ ) & (~\new_[19920]_  | ~\new_[16416]_ );
  assign \new_[12517]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][30] ;
  assign \new_[12518]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][28] ;
  assign \new_[12519]_  = (~\new_[13693]_  | ~\new_[10868]_ ) & (~\new_[19920]_  | ~\new_[16112]_ );
  assign \new_[12520]_  = (~\new_[13694]_  | ~\new_[11046]_ ) & (~\new_[19920]_  | ~\new_[16632]_ );
  assign \new_[12521]_  = (~\new_[13694]_  | ~\new_[11047]_ ) & (~\new_[19920]_  | ~\new_[16635]_ );
  assign \new_[12522]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][29] ;
  assign \new_[12523]_  = \\configuration_wb_err_addr_reg[30] ;
  assign \new_[12524]_  = \\configuration_wb_err_addr_reg[29] ;
  assign \new_[12525]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][19] ;
  assign \new_[12526]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][35] ;
  assign \new_[12527]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][16] ;
  assign \new_[12528]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][28] ;
  assign \new_[12529]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][17] ;
  assign \new_[12530]_  = (~\new_[13693]_  | ~\new_[10867]_ ) & (~\new_[19920]_  | ~\new_[16114]_ );
  assign \new_[12531]_  = (~\new_[13694]_  | ~\new_[11031]_ ) & (~\new_[19920]_  | ~\new_[16634]_ );
  assign \new_[12532]_  = \\configuration_wb_err_addr_reg[25] ;
  assign \new_[12533]_  = (~\new_[13693]_  | ~\new_[10866]_ ) & (~\new_[19920]_  | ~\new_[16123]_ );
  assign \new_[12534]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][2] ;
  assign \new_[12535]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][3] ;
  assign \new_[12536]_  = \\configuration_wb_err_addr_reg[27] ;
  assign \new_[12537]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][38] ;
  assign \new_[12538]_  = ~\new_[13703]_  & ~\new_[14245]_ ;
  assign n10600 = \new_[10388]_  ? \new_[15633]_  : \new_[13834]_ ;
  assign n13045 = \new_[10391]_  ? \new_[15633]_  : \new_[13835]_ ;
  assign n13055 = \new_[10358]_  ? \new_[15633]_  : \new_[13833]_ ;
  assign \new_[12542]_  = ~\new_[13208]_ ;
  assign \new_[12543]_  = ~\new_[13711]_  & (~\new_[11955]_  | ~\new_[20056]_ );
  assign n12210 = \new_[10387]_  ? \new_[15633]_  : \new_[13837]_ ;
  assign \new_[12545]_  = ~\new_[19935]_ ;
  assign n12200 = \new_[13876]_  ? \new_[15485]_  : \new_[18010]_ ;
  assign \new_[12547]_  = ~\new_[13702]_  & (~\new_[11069]_  | ~\new_[20506]_ );
  assign \new_[12548]_  = \\pci_target_unit_fifos_pciw_inTransactionCount_reg[0] ;
  assign \new_[12549]_  = ~\\pci_target_unit_fifos_inGreyCount_reg[1] ;
  assign n12185 = \new_[13877]_  ? \new_[15488]_  : \new_[18028]_ ;
  assign n12215 = \new_[13875]_  ? \new_[15491]_  : \new_[18025]_ ;
  assign n12205 = \new_[13871]_  ? \new_[15591]_  : \new_[17996]_ ;
  assign n10610 = \new_[13878]_  ? \new_[15488]_  : \new_[19064]_ ;
  assign n10615 = \new_[13879]_  ? \new_[15489]_  : \new_[19153]_ ;
  assign n12160 = \new_[13880]_  ? \new_[15592]_  : \new_[19805]_ ;
  assign n10605 = ~\new_[16678]_  | ~\new_[15098]_  | ~\new_[14290]_  | ~\new_[13848]_ ;
  assign n10620 = \new_[13885]_  ? \new_[15492]_  : \new_[17818]_ ;
  assign n12920 = \new_[13886]_  ? \new_[15591]_  : \new_[19766]_ ;
  assign n12910 = \new_[13887]_  ? \new_[15273]_  : \new_[18182]_ ;
  assign n10625 = \new_[13889]_  ? \new_[15493]_  : \new_[18017]_ ;
  assign n10630 = \new_[13890]_  ? \new_[15591]_  : \new_[19095]_ ;
  assign n10635 = \new_[13891]_  ? \new_[15488]_  : \new_[18016]_ ;
  assign n12900 = \new_[13888]_  ? \new_[15485]_  : \new_[18243]_ ;
  assign n10640 = \new_[13892]_  ? \new_[15488]_  : \new_[19096]_ ;
  assign \new_[12565]_  = ~\new_[20121]_  | ~\new_[17383]_ ;
  assign \new_[12566]_  = ~\new_[20121]_  | ~\new_[17080]_ ;
  assign \new_[12567]_  = ~\new_[20121]_  | ~\new_[20143]_ ;
  assign \new_[12568]_  = ~\new_[13717]_  | ~\new_[20340]_ ;
  assign \new_[12569]_  = ~\new_[13717]_  | ~\new_[17383]_ ;
  assign \new_[12570]_  = ~\new_[14250]_  | ~\new_[11328]_ ;
  assign \new_[12571]_  = ~\new_[13716]_  & ~\new_[11328]_ ;
  assign \new_[12572]_  = ~\new_[4458]_  | ~\new_[13718]_ ;
  assign \new_[12573]_  = ~\new_[4459]_  | ~\new_[13718]_ ;
  assign \new_[12574]_  = ~\new_[4460]_  | ~\new_[13718]_ ;
  assign \new_[12575]_  = ~\new_[14278]_  & ~\new_[20216]_ ;
  assign \new_[12576]_  = ~\new_[16073]_  | ~\new_[17033]_  | ~\new_[20129]_  | ~\new_[16829]_ ;
  assign n12660 = n17050 ? \new_[14878]_  : \new_[16614]_ ;
  assign n12765 = ~\new_[13715]_  & ~\new_[14562]_ ;
  assign n10530 = \new_[19327]_  ? \new_[13897]_  : \new_[13950]_ ;
  assign n10695 = \new_[18276]_  ? \new_[13897]_  : \new_[14582]_ ;
  assign n10470 = \new_[17906]_  ? \new_[13896]_  : \new_[13961]_ ;
  assign n10675 = \new_[19030]_  ? \new_[13898]_  : \new_[13947]_ ;
  assign n10680 = \new_[18136]_  ? \new_[13899]_  : \new_[14731]_ ;
  assign n12520 = \new_[17874]_  ? \new_[13899]_  : \new_[14729]_ ;
  assign n10685 = \new_[19585]_  ? \new_[13904]_  : \new_[14726]_ ;
  assign n12485 = \new_[18139]_  ? \new_[13896]_  : \new_[14079]_ ;
  assign n10690 = \new_[19412]_  ? \new_[13894]_  : \new_[14046]_ ;
  assign n12115 = \new_[19413]_  ? \new_[13898]_  : \new_[14661]_ ;
  assign n10700 = \new_[19415]_  ? \new_[13903]_  : \new_[14689]_ ;
  assign n12190 = \new_[19427]_  ? \new_[14917]_  : \new_[14019]_ ;
  assign n10705 = \new_[18141]_  ? \new_[13838]_  : \new_[14039]_ ;
  assign n12335 = \new_[18391]_  ? \new_[13899]_  : \new_[13992]_ ;
  assign n10710 = \new_[18143]_  ? \new_[13903]_  : \new_[14596]_ ;
  assign n12385 = \new_[18146]_  ? \new_[13910]_  : \new_[14727]_ ;
  assign n10715 = \new_[18221]_  ? \new_[13897]_  : \new_[14096]_ ;
  assign n12320 = \new_[19231]_  ? \new_[13895]_  : \new_[14732]_ ;
  assign n10720 = \new_[19234]_  ? \new_[13908]_  : \new_[14734]_ ;
  assign n10725 = \new_[18165]_  ? \new_[14881]_  : \new_[14038]_ ;
  assign n10730 = \new_[18226]_  ? \new_[14919]_  : \new_[14576]_ ;
  assign n12290 = \new_[19248]_  ? \new_[13898]_  : \new_[14092]_ ;
  assign n10735 = \new_[18180]_  ? \new_[13902]_  : \new_[14110]_ ;
  assign n10740 = \new_[19259]_  ? \new_[13903]_  : \new_[14022]_ ;
  assign n10745 = \new_[19541]_  ? \new_[13895]_  : \new_[13954]_ ;
  assign n12125 = \new_[17883]_  ? \new_[14917]_  : \new_[13946]_ ;
  assign n10840 = \new_[18792]_  ? \new_[14921]_  : \new_[14590]_ ;
  assign n10750 = \new_[18236]_  ? \new_[13895]_  : \new_[14574]_ ;
  assign n12075 = \new_[19694]_  ? \new_[13900]_  : \new_[14097]_ ;
  assign n12080 = \new_[18246]_  ? \new_[13839]_  : \new_[14747]_ ;
  assign n10755 = \new_[18700]_  ? \new_[13898]_  : \new_[13948]_ ;
  assign n10760 = \new_[18248]_  ? \new_[13899]_  : \new_[14581]_ ;
  assign n11995 = \new_[18403]_  ? \new_[14878]_  : \new_[14593]_ ;
  assign n10765 = \new_[19287]_  ? \new_[13902]_  : \new_[14090]_ ;
  assign n11970 = \new_[18864]_  ? \new_[13911]_  : \new_[14579]_ ;
  assign n10770 = \new_[18259]_  ? \new_[14944]_  : \new_[13945]_ ;
  assign n10775 = \new_[18719]_  ? \new_[13899]_  : \new_[14577]_ ;
  assign n10360 = \new_[18267]_  ? \new_[14878]_  : \new_[14583]_ ;
  assign n10780 = \new_[19540]_  ? \new_[14916]_  : \new_[13941]_ ;
  assign n10430 = \new_[18266]_  ? \new_[13894]_  : \new_[13949]_ ;
  assign n10785 = \new_[19509]_  ? \new_[13906]_  : \new_[14575]_ ;
  assign n10480 = \new_[19596]_  ? \new_[14918]_  : \new_[14584]_ ;
  assign n10790 = \new_[18489]_  ? \new_[14919]_  : \new_[13939]_ ;
  assign n10795 = \new_[19539]_  ? \new_[14919]_  : \new_[14071]_ ;
  assign n10560 = \new_[18291]_  ? \new_[13904]_  : \new_[14585]_ ;
  assign n10800 = \new_[18305]_  ? \new_[13904]_  : \new_[14601]_ ;
  assign n10805 = \new_[18327]_  ? \new_[13897]_  : \new_[14603]_ ;
  assign n10555 = \new_[19275]_  ? \new_[13902]_  : \new_[14586]_ ;
  assign n10810 = \new_[19536]_  ? \new_[13909]_  : \new_[13966]_ ;
  assign n10510 = \new_[19534]_  ? \new_[13903]_  : \new_[14587]_ ;
  assign n10815 = \new_[19535]_  ? \new_[13895]_  : \new_[13965]_ ;
  assign n10820 = \new_[19703]_  ? \new_[13895]_  : \new_[13962]_ ;
  assign n10540 = \new_[18942]_  ? \new_[14919]_  : \new_[13953]_ ;
  assign n10830 = \new_[19533]_  ? \new_[14917]_  : \new_[13937]_ ;
  assign n10825 = \new_[18330]_  ? \new_[14921]_  : \new_[14588]_ ;
  assign n10515 = \new_[18361]_  ? \new_[14921]_  : \new_[13955]_ ;
  assign n10835 = \new_[18358]_  ? \new_[13895]_  : \new_[14589]_ ;
  assign n10520 = \new_[19439]_  ? \new_[13895]_  : \new_[13957]_ ;
  assign n10435 = \new_[19532]_  ? \new_[13906]_  : \new_[14748]_ ;
  assign n10845 = \new_[18716]_  ? \new_[13900]_  : \new_[14591]_ ;
  assign n10490 = \new_[17898]_  ? \new_[13896]_  : \new_[14108]_ ;
  assign n10850 = \new_[18363]_  ? \new_[13905]_  : \new_[14056]_ ;
  assign n10500 = \new_[18365]_  ? \new_[13898]_  : \new_[14745]_ ;
  assign n10855 = \new_[18369]_  ? \new_[14878]_  : \new_[14594]_ ;
  assign n10495 = \new_[18763]_  ? \new_[13912]_  : \new_[14738]_ ;
  assign n10860 = \new_[18704]_  ? \new_[13838]_  : \new_[14089]_ ;
  assign n10865 = \new_[18755]_  ? \new_[13904]_  : \new_[13956]_ ;
  assign n10485 = \new_[18834]_  ? \new_[13904]_  : \new_[14730]_ ;
  assign n10880 = \new_[19348]_  ? \new_[13910]_  : \new_[13958]_ ;
  assign n10885 = \new_[19432]_  ? \new_[13903]_  : \new_[13959]_ ;
  assign n10460 = \new_[18611]_  ? \new_[13902]_  : \new_[14703]_ ;
  assign n10890 = \new_[18650]_  ? \new_[13838]_  : \new_[14698]_ ;
  assign n10895 = \new_[18446]_  ? \new_[13838]_  : \new_[13960]_ ;
  assign n10900 = \new_[19350]_  ? \new_[13899]_  : \new_[14595]_ ;
  assign n10475 = \new_[17905]_  ? \new_[14918]_  : \new_[14706]_ ;
  assign n10905 = \new_[18613]_  ? \new_[13896]_  : \new_[13999]_ ;
  assign n10465 = \new_[18887]_  ? \new_[13907]_  : \new_[14580]_ ;
  assign n10445 = \new_[18397]_  ? \new_[13898]_  : \new_[13943]_ ;
  assign n10455 = \new_[19283]_  ? \new_[13905]_  : \new_[14109]_ ;
  assign n12390 = \new_[19526]_  ? \new_[13903]_  : \new_[13963]_ ;
  assign n10910 = \new_[19527]_  ? \new_[13838]_  : \new_[14074]_ ;
  assign n12785 = \new_[19515]_  ? \new_[13898]_  : \new_[14692]_ ;
  assign n12795 = \new_[19522]_  ? \new_[13901]_  : \new_[14045]_ ;
  assign n10915 = \new_[19525]_  ? \new_[14920]_  : \new_[14691]_ ;
  assign n12895 = \new_[19713]_  ? \new_[14918]_  : \new_[14026]_ ;
  assign n10920 = \new_[19422]_  ? \new_[13909]_  : \new_[14639]_ ;
  assign n10925 = \new_[19524]_  ? \new_[13901]_  : \new_[14602]_ ;
  assign n10930 = \new_[17917]_  ? \new_[13904]_  : \new_[14598]_ ;
  assign n10535 = \new_[18320]_  ? \new_[13838]_  : \new_[13952]_ ;
  assign n12885 = \new_[19133]_  ? \new_[13904]_  : \new_[13964]_ ;
  assign n10935 = \new_[18449]_  ? \new_[13904]_  : \new_[14104]_ ;
  assign n12870 = \new_[19374]_  ? \new_[13903]_  : \new_[14604]_ ;
  assign n10940 = \new_[19521]_  ? \new_[13897]_  : \new_[14735]_ ;
  assign n12835 = \new_[19376]_  ? \new_[13902]_  : \new_[14605]_ ;
  assign n10945 = \new_[18244]_  ? \new_[13902]_  : \new_[14094]_ ;
  assign n12855 = \new_[19516]_  ? \new_[13838]_  : \new_[13968]_ ;
  assign n10950 = \new_[18995]_  ? \new_[13909]_  : \new_[14572]_ ;
  assign n12860 = \new_[18463]_  ? \new_[13912]_  : \new_[14606]_ ;
  assign n10955 = \new_[19382]_  ? \new_[13901]_  : \new_[14091]_ ;
  assign n10965 = \new_[18479]_  ? \new_[13895]_  : \new_[14035]_ ;
  assign n12840 = \new_[19513]_  ? \new_[13901]_  : \new_[14607]_ ;
  assign n10970 = \new_[18546]_  ? \new_[13838]_  : \new_[14740]_ ;
  assign n12800 = \new_[18470]_  ? \new_[13895]_  : \new_[13970]_ ;
  assign n12820 = \new_[18883]_  ? \new_[13899]_  : \new_[14608]_ ;
  assign n10985 = \new_[17932]_  ? \new_[14919]_  : \new_[14737]_ ;
  assign n10545 = \new_[19315]_  ? \new_[13900]_  : \new_[13951]_ ;
  assign n12750 = \new_[19510]_  ? \new_[13908]_  : \new_[13971]_ ;
  assign n10995 = \new_[19511]_  ? \new_[13905]_  : \new_[14101]_ ;
  assign n12780 = \new_[18985]_  ? \new_[13838]_  : \new_[14610]_ ;
  assign n11010 = \new_[18646]_  ? \new_[14921]_  : \new_[14611]_ ;
  assign n12720 = \new_[19339]_  ? \new_[13894]_  : \new_[14037]_ ;
  assign n11020 = \new_[19503]_  ? \new_[13904]_  : \new_[14573]_ ;
  assign n11025 = \new_[18495]_  ? \new_[13838]_  : \new_[14613]_ ;
  assign n12680 = \new_[19024]_  ? \new_[13895]_  : \new_[14112]_ ;
  assign n11030 = \new_[18550]_  ? \new_[13908]_  : \new_[14615]_ ;
  assign n12700 = \new_[18525]_  ? \new_[13906]_  : \new_[13973]_ ;
  assign n11035 = \new_[19505]_  ? \new_[13902]_  : \new_[14663]_ ;
  assign n12410 = \new_[17842]_  ? \new_[14878]_  : \new_[14616]_ ;
  assign n11040 = \new_[19504]_  ? \new_[13902]_  : \new_[14741]_ ;
  assign n11045 = \new_[18566]_  ? \new_[13905]_  : \new_[13974]_ ;
  assign n11050 = \new_[19303]_  ? \new_[13895]_  : \new_[14098]_ ;
  assign n12635 = \new_[18281]_  ? \new_[13904]_  : \new_[14617]_ ;
  assign n11055 = \new_[19304]_  ? \new_[13899]_  : \new_[14733]_ ;
  assign n12595 = \new_[18217]_  ? \new_[14922]_  : \new_[13975]_ ;
  assign n12535 = \new_[18882]_  ? \new_[14944]_  : \new_[13976]_ ;
  assign n12570 = \new_[18468]_  ? \new_[13905]_  : \new_[13977]_ ;
  assign n11060 = \new_[18880]_  ? \new_[13899]_  : \new_[14722]_ ;
  assign n12415 = \new_[17938]_  ? \new_[13903]_  : \new_[14618]_ ;
  assign n12480 = \new_[18643]_  ? \new_[13898]_  : \new_[13978]_ ;
  assign n12490 = \new_[18602]_  ? \new_[14878]_  : \new_[14619]_ ;
  assign n12175 = \new_[19502]_  ? \new_[13899]_  : \new_[14723]_ ;
  assign n12110 = \new_[18865]_  ? \new_[13906]_  : \new_[13979]_ ;
  assign n12235 = \new_[18812]_  ? \new_[13898]_  : \new_[14620]_ ;
  assign n12195 = \new_[19307]_  ? \new_[13912]_  : \new_[14077]_ ;
  assign n11065 = \new_[18768]_  ? \new_[13904]_  : \new_[14083]_ ;
  assign n12325 = \new_[18714]_  ? \new_[13896]_  : \new_[13980]_ ;
  assign n12360 = \new_[18780]_  ? \new_[13910]_  : \new_[14081]_ ;
  assign n12375 = \new_[17940]_  ? \new_[13906]_  : \new_[13981]_ ;
  assign n11075 = \new_[18793]_  ? \new_[13838]_  : \new_[14719]_ ;
  assign n11070 = \new_[19500]_  ? \new_[13913]_  : \new_[14078]_ ;
  assign n12355 = \new_[17941]_  ? \new_[13904]_  : \new_[14717]_ ;
  assign n11080 = \new_[19142]_  ? \new_[13838]_  : \new_[14073]_ ;
  assign n12260 = \new_[18593]_  ? \new_[13894]_  : \new_[14716]_ ;
  assign n11085 = \new_[18914]_  ? \new_[13894]_  : \new_[14621]_ ;
  assign n12295 = \new_[18902]_  ? \new_[13838]_  : \new_[14714]_ ;
  assign n11090 = \new_[18591]_  ? \new_[14919]_  : \new_[13982]_ ;
  assign n11095 = \new_[18345]_  ? \new_[13838]_  : \new_[14712]_ ;
  assign n11100 = \new_[19453]_  ? \new_[14918]_  : \new_[13983]_ ;
  assign n12090 = \new_[18183]_  ? \new_[13894]_  : \new_[14622]_ ;
  assign n12095 = \new_[19398]_  ? \new_[14878]_  : \new_[14711]_ ;
  assign n12100 = \new_[19499]_  ? \new_[13900]_  : \new_[14623]_ ;
  assign n10450 = \new_[17890]_  ? \new_[13913]_  : \new_[13984]_ ;
  assign n11960 = \new_[17827]_  ? \new_[13901]_  : \new_[13985]_ ;
  assign n11105 = \new_[17869]_  ? \new_[13909]_  : \new_[14709]_ ;
  assign n10440 = \new_[18742]_  ? \new_[13896]_  : \new_[14624]_ ;
  assign n12515 = \new_[18862]_  ? \new_[13911]_  : \new_[14065]_ ;
  assign n12465 = \new_[19375]_  ? \new_[13900]_  : \new_[13986]_ ;
  assign n11110 = \new_[18336]_  ? \new_[13900]_  : \new_[14063]_ ;
  assign n12425 = \new_[19871]_  ? \new_[13838]_  : \new_[14707]_ ;
  assign n11115 = \new_[18474]_  ? \new_[13898]_  : \new_[14625]_ ;
  assign n12740 = \new_[19579]_  ? \new_[13896]_  : \new_[13987]_ ;
  assign n11120 = \new_[19437]_  ? \new_[13838]_  : \new_[14704]_ ;
  assign n11125 = \new_[19225]_  ? \new_[13894]_  : \new_[14702]_ ;
  assign n11130 = \new_[19629]_  ? \new_[13900]_  : \new_[14058]_ ;
  assign n12690 = \new_[19654]_  ? \new_[13908]_  : \new_[14626]_ ;
  assign n11135 = \new_[19637]_  ? \new_[13897]_  : \new_[14057]_ ;
  assign n12435 = \new_[19729]_  ? \new_[13901]_  : \new_[13988]_ ;
  assign n11140 = \new_[17960]_  ? \new_[13904]_  : \new_[14055]_ ;
  assign n12600 = \new_[17961]_  ? \new_[14920]_  : \new_[13989]_ ;
  assign n11150 = \new_[19666]_  ? \new_[13901]_  : \new_[14054]_ ;
  assign n11145 = \new_[18998]_  ? \new_[14918]_  : \new_[14699]_ ;
  assign n12625 = \new_[18911]_  ? \new_[13909]_  : \new_[13990]_ ;
  assign n11155 = \new_[19311]_  ? \new_[13902]_  : \new_[14627]_ ;
  assign n12585 = \new_[18872]_  ? \new_[13901]_  : \new_[14051]_ ;
  assign n11160 = \new_[18395]_  ? \new_[13904]_  : \new_[14697]_ ;
  assign n12545 = \new_[19004]_  ? \new_[13902]_  : \new_[14695]_ ;
  assign n11170 = \new_[19850]_  ? \new_[13902]_  : \new_[14628]_ ;
  assign n12575 = \new_[17963]_  ? \new_[13838]_  : \new_[14049]_ ;
  assign n11175 = \new_[19848]_  ? \new_[13838]_  : \new_[14629]_ ;
  assign n12450 = \new_[19695]_  ? \new_[13838]_  : \new_[14048]_ ;
  assign n11180 = \new_[19430]_  ? \new_[13898]_  : \new_[14694]_ ;
  assign n12510 = \new_[19045]_  ? \new_[13898]_  : \new_[14630]_ ;
  assign n11185 = \new_[18349]_  ? \new_[13838]_  : \new_[14631]_ ;
  assign n12500 = \new_[17965]_  ? \new_[13900]_  : \new_[14042]_ ;
  assign n11190 = \new_[19489]_  ? \new_[13900]_  : \new_[14041]_ ;
  assign n11195 = \new_[17966]_  ? \new_[14916]_  : \new_[14632]_ ;
  assign n11200 = \new_[18632]_  ? \new_[14916]_  : \new_[14633]_ ;
  assign n12105 = \new_[18294]_  ? \new_[13903]_  : \new_[13993]_ ;
  assign n11205 = \new_[18519]_  ? \new_[13902]_  : \new_[14040]_ ;
  assign n12905 = \new_[19523]_  ? \new_[14881]_  : \new_[14597]_ ;
  assign n11215 = \new_[17808]_  ? \new_[14881]_  : \new_[14690]_ ;
  assign n12305 = \new_[19314]_  ? \new_[13902]_  : \new_[14635]_ ;
  assign n11225 = \new_[17968]_  ? \new_[13902]_  : \new_[14636]_ ;
  assign n11230 = \new_[19481]_  ? \new_[13902]_  : \new_[14634]_ ;
  assign n12345 = \new_[18531]_  ? \new_[13838]_  : \new_[13995]_ ;
  assign n11235 = \new_[19099]_  ? \new_[13898]_  : \new_[14578]_ ;
  assign n12285 = \new_[19093]_  ? \new_[13898]_  : \new_[13944]_ ;
  assign n11240 = \new_[19631]_  ? \new_[13895]_  : \new_[13996]_ ;
  assign n12270 = \new_[17846]_  ? \new_[13895]_  : \new_[13997]_ ;
  assign n11245 = \new_[19485]_  ? \new_[13912]_  : \new_[13967]_ ;
  assign n11250 = \new_[17845]_  ? \new_[13903]_  : \new_[13940]_ ;
  assign n11255 = \new_[17870]_  ? \new_[13901]_  : \new_[14637]_ ;
  assign n12120 = \new_[19196]_  ? \new_[13895]_  : \new_[13998]_ ;
  assign n11945 = \new_[17974]_  ? \new_[13896]_  : \new_[14638]_ ;
  assign n11260 = \new_[17837]_  ? \new_[13901]_  : \new_[14000]_ ;
  assign n11985 = \new_[17975]_  ? \new_[13838]_  : \new_[14693]_ ;
  assign n11265 = \new_[18078]_  ? \new_[13901]_  : \new_[14688]_ ;
  assign n10410 = \new_[19483]_  ? \new_[13901]_  : \new_[14686]_ ;
  assign n11270 = \new_[18039]_  ? \new_[13902]_  : \new_[14001]_ ;
  assign n12455 = \new_[19482]_  ? \new_[13902]_  : \new_[14687]_ ;
  assign n11275 = \new_[19319]_  ? \new_[13899]_  : \new_[14113]_ ;
  assign n12685 = \new_[18958]_  ? \new_[13899]_  : \new_[14640]_ ;
  assign n12755 = \new_[19479]_  ? \new_[13897]_  : \new_[14642]_ ;
  assign n11285 = \new_[19480]_  ? \new_[13897]_  : \new_[14060]_ ;
  assign n11290 = \new_[18744]_  ? \new_[13900]_  : \new_[14002]_ ;
  assign n11295 = \new_[18782]_  ? \new_[14917]_  : \new_[14713]_ ;
  assign n12675 = \new_[19475]_  ? \new_[13908]_  : \new_[14643]_ ;
  assign n11300 = \new_[19478]_  ? \new_[13905]_  : \new_[14111]_ ;
  assign n11305 = \new_[18937]_  ? \new_[13908]_  : \new_[14003]_ ;
  assign n11310 = \new_[18282]_  ? \new_[13908]_  : \new_[14004]_ ;
  assign n12550 = \new_[19476]_  ? \new_[13838]_  : \new_[14644]_ ;
  assign n11315 = \new_[19119]_  ? \new_[13839]_  : \new_[14724]_ ;
  assign n11320 = \new_[17902]_  ? \new_[14878]_  : \new_[14088]_ ;
  assign n11325 = \new_[17899]_  ? \new_[14878]_  : \new_[14645]_ ;
  assign n12640 = \new_[19681]_  ? \new_[13895]_  : \new_[14646]_ ;
  assign n11330 = \new_[18355]_  ? \new_[13895]_  : \new_[14080]_ ;
  assign n12630 = \new_[19474]_  ? \new_[13894]_  : \new_[14647]_ ;
  assign n11335 = \new_[17931]_  ? \new_[13838]_  : \new_[14076]_ ;
  assign n12605 = \new_[19323]_  ? \new_[13904]_  : \new_[14005]_ ;
  assign n11340 = \new_[18304]_  ? \new_[13838]_  : \new_[14075]_ ;
  assign n11345 = \new_[19473]_  ? \new_[13907]_  : \new_[14006]_ ;
  assign n11350 = \new_[19131]_  ? \new_[13907]_  : \new_[14007]_ ;
  assign n12540 = \new_[19471]_  ? \new_[14878]_  : \new_[14648]_ ;
  assign n12420 = \new_[19472]_  ? \new_[14878]_  : \new_[14070]_ ;
  assign n12505 = \new_[17948]_  ? \new_[13900]_  : \new_[14649]_ ;
  assign n12525 = \new_[19310]_  ? \new_[13906]_  : \new_[14053]_ ;
  assign n12495 = \new_[19491]_  ? \new_[13906]_  : \new_[14650]_ ;
  assign n12470 = \new_[19520]_  ? \new_[13902]_  : \new_[14651]_ ;
  assign n12395 = \new_[18674]_  ? \new_[13900]_  : \new_[14652]_ ;
  assign n10415 = \new_[18241]_  ? \new_[14878]_  : \new_[14047]_ ;
  assign n11360 = \new_[19469]_  ? \new_[13902]_  : \new_[14653]_ ;
  assign n12180 = \new_[19324]_  ? \new_[13894]_  : \new_[14044]_ ;
  assign n11365 = \new_[18405]_  ? \new_[13894]_  : \new_[14654]_ ;
  assign n12240 = \new_[19571]_  ? \new_[13905]_  : \new_[14655]_ ;
  assign n11370 = \new_[18209]_  ? \new_[14922]_  : \new_[14746]_ ;
  assign n12365 = \new_[19325]_  ? \new_[13839]_  : \new_[14008]_ ;
  assign n12370 = \new_[19862]_  ? \new_[14878]_  : \new_[14009]_ ;
  assign n12310 = \new_[18229]_  ? \new_[13906]_  : \new_[14656]_ ;
  assign n12340 = \new_[19586]_  ? \new_[13901]_  : \new_[14742]_ ;
  assign n12245 = \new_[17881]_  ? \new_[13895]_  : \new_[14010]_ ;
  assign n12275 = \new_[18026]_  ? \new_[13838]_  : \new_[14103]_ ;
  assign n12300 = \new_[19177]_  ? \new_[14922]_  : \new_[14011]_ ;
  assign n11375 = \new_[19170]_  ? \new_[14944]_  : \new_[14728]_ ;
  assign n11965 = \new_[19146]_  ? \new_[13906]_  : \new_[14657]_ ;
  assign n11380 = \new_[19644]_  ? \new_[13906]_  : \new_[14086]_ ;
  assign n11975 = \new_[18042]_  ? \new_[13838]_  : \new_[14658]_ ;
  assign n10425 = \new_[18043]_  ? \new_[13838]_  : \new_[14721]_ ;
  assign n11165 = \new_[18045]_  ? \new_[13899]_  : \new_[14012]_ ;
  assign n10420 = \new_[18044]_  ? \new_[13903]_  : \new_[14720]_ ;
  assign n12445 = \new_[19326]_  ? \new_[13903]_  : \new_[14013]_ ;
  assign n11390 = \new_[18048]_  ? \new_[13898]_  : \new_[14082]_ ;
  assign n12460 = \new_[19135]_  ? \new_[13899]_  : \new_[14014]_ ;
  assign n12695 = \new_[18050]_  ? \new_[13899]_  : \new_[14015]_ ;
  assign n12650 = \new_[19467]_  ? \new_[13894]_  : \new_[14016]_ ;
  assign n11395 = \new_[18060]_  ? \new_[13894]_  : \new_[14715]_ ;
  assign n12715 = \new_[19129]_  ? \new_[13901]_  : \new_[14017]_ ;
  assign n12670 = \new_[18059]_  ? \new_[13904]_  : \new_[14609]_ ;
  assign n11400 = \new_[19702]_  ? \new_[13838]_  : \new_[14018]_ ;
  assign n12665 = \new_[18280]_  ? \new_[13907]_  : \new_[14659]_ ;
  assign n12400 = \new_[18145]_  ? \new_[13902]_  : \new_[14660]_ ;
  assign n12555 = \new_[18109]_  ? \new_[13896]_  : \new_[14710]_ ;
  assign n12590 = \new_[18672]_  ? \new_[13905]_  : \new_[14067]_ ;
  assign n12620 = \new_[18686]_  ? \new_[13907]_  : \new_[14708]_ ;
  assign n12645 = \new_[18000]_  ? \new_[13910]_  : \new_[14107]_ ;
  assign n11405 = \new_[18867]_  ? \new_[13896]_  : \new_[14739]_ ;
  assign n12615 = \new_[18859]_  ? \new_[13894]_  : \new_[14662]_ ;
  assign n11410 = \new_[18656]_  ? \new_[13838]_  : \new_[14664]_ ;
  assign n12565 = \new_[18750]_  ? \new_[13902]_  : \new_[14020]_ ;
  assign n11415 = \new_[18855]_  ? \new_[13903]_  : \new_[14100]_ ;
  assign n12580 = \new_[19464]_  ? \new_[13904]_  : \new_[14665]_ ;
  assign n11420 = \new_[18114]_  ? \new_[13899]_  : \new_[14744]_ ;
  assign n12430 = \new_[19213]_  ? \new_[13899]_  : \new_[14021]_ ;
  assign n11425 = \new_[19455]_  ? \new_[13895]_  : \new_[14106]_ ;
  assign n11430 = \new_[18765]_  ? \new_[13905]_  : \new_[14023]_ ;
  assign n11435 = \new_[18842]_  ? \new_[13913]_  : \new_[14666]_ ;
  assign n12475 = \new_[19215]_  ? \new_[13898]_  : \new_[14667]_ ;
  assign n11440 = \new_[18795]_  ? \new_[13911]_  : \new_[14095]_ ;
  assign n10525 = \new_[18698]_  ? \new_[13908]_  : \new_[14668]_ ;
  assign n11445 = \new_[19220]_  ? \new_[13904]_  : \new_[14669]_ ;
  assign n12265 = \new_[19599]_  ? \new_[13838]_  : \new_[14024]_ ;
  assign n11450 = \new_[18721]_  ? \new_[13908]_  : \new_[14718]_ ;
  assign n12350 = \new_[18740]_  ? \new_[14944]_  : \new_[14066]_ ;
  assign n12380 = \new_[18817]_  ? \new_[13900]_  : \new_[14027]_ ;
  assign n11455 = \new_[18836]_  ? \new_[13894]_  : \new_[14062]_ ;
  assign n12315 = \new_[18118]_  ? \new_[13902]_  : \new_[14061]_ ;
  assign n12250 = \new_[18831]_  ? \new_[13896]_  : \new_[14705]_ ;
  assign n12280 = \new_[19461]_  ? \new_[14920]_  : \new_[14028]_ ;
  assign n12135 = \new_[19328]_  ? \new_[13899]_  : \new_[14670]_ ;
  assign n11460 = \new_[19221]_  ? \new_[13895]_  : \new_[14029]_ ;
  assign n11980 = \new_[18558]_  ? \new_[13902]_  : \new_[14701]_ ;
  assign n12005 = \new_[19329]_  ? \new_[13839]_  : \new_[14671]_ ;
  assign n12010 = \new_[19330]_  ? \new_[13904]_  : \new_[14672]_ ;
  assign n11950 = \new_[18319]_  ? \new_[13899]_  : \new_[14030]_ ;
  assign n11955 = \new_[18620]_  ? \new_[13896]_  : \new_[14700]_ ;
  assign n11465 = \new_[18895]_  ? \new_[13907]_  : \new_[14052]_ ;
  assign n12405 = \new_[18916]_  ? \new_[13901]_  : \new_[14673]_ ;
  assign n13035 = \new_[19458]_  ? \new_[14878]_  : \new_[14696]_ ;
  assign n13040 = \new_[18008]_  ? \new_[13912]_  : \new_[14674]_ ;
  assign n11470 = \new_[18587]_  ? \new_[13913]_  : \new_[14050]_ ;
  assign n11550 = \new_[18125]_  ? \new_[13899]_  : \new_[13991]_ ;
  assign n12145 = \new_[18009]_  ? \new_[13900]_  : \new_[14675]_ ;
  assign n12085 = \new_[19457]_  ? \new_[14881]_  : \new_[14676]_ ;
  assign n12150 = \new_[17849]_  ? \new_[13905]_  : \new_[14085]_ ;
  assign n12140 = \new_[18128]_  ? \new_[13838]_  : \new_[14084]_ ;
  assign n12020 = \new_[18011]_  ? \new_[14916]_  : \new_[14031]_ ;
  assign n12165 = ~\new_[13698]_  | (~\new_[14242]_  & ~\new_[16103]_ );
  assign n12050 = \new_[19456]_  ? \new_[13899]_  : \new_[14677]_ ;
  assign n12045 = \new_[18012]_  ? \new_[13838]_  : \new_[14600]_ ;
  assign n12065 = \new_[18129]_  ? \new_[13911]_  : \new_[14032]_ ;
  assign n12070 = \new_[18013]_  ? \new_[13897]_  : \new_[14678]_ ;
  assign n12055 = \new_[19037]_  ? \new_[13838]_  : \new_[14679]_ ;
  assign n11475 = \new_[18130]_  ? \new_[13894]_  : \new_[14069]_ ;
  assign n12060 = \new_[18131]_  ? \new_[14916]_  : \new_[14680]_ ;
  assign n11480 = \new_[18132]_  ? \new_[13907]_  : \new_[14059]_ ;
  assign n12015 = \new_[19588]_  ? \new_[13900]_  : \new_[14033]_ ;
  assign n11485 = \new_[18456]_  ? \new_[13897]_  : \new_[14068]_ ;
  assign n11490 = \new_[18927]_  ? \new_[13898]_  : \new_[14034]_ ;
  assign n11495 = \new_[19587]_  ? \new_[13838]_  : \new_[14064]_ ;
  assign n12035 = \new_[18965]_  ? \new_[13900]_  : \new_[14681]_ ;
  assign n12040 = \new_[18137]_  ? \new_[13907]_  : \new_[14043]_ ;
  assign n11500 = \new_[19831]_  ? \new_[13909]_  : \new_[14682]_ ;
  assign n12030 = \new_[18142]_  ? \new_[13897]_  : \new_[13942]_ ;
  assign n11505 = \new_[19228]_  ? \new_[13902]_  : \new_[14683]_ ;
  assign n11510 = \new_[18138]_  ? \new_[13897]_  : \new_[14725]_ ;
  assign n11515 = \new_[19229]_  ? \new_[13897]_  : \new_[14684]_ ;
  assign n12025 = \new_[19423]_  ? \new_[13906]_  : \new_[14087]_ ;
  assign n11520 = \new_[18383]_  ? \new_[14881]_  : \new_[14685]_ ;
  assign n11015 = \new_[19340]_  ? \new_[13897]_  : \new_[14612]_ ;
  assign n11220 = \new_[19488]_  ? \new_[13897]_  : \new_[14036]_ ;
  assign n11210 = \new_[19084]_  ? \new_[13902]_  : \new_[13994]_ ;
  assign n12230 = \new_[18743]_  ? \new_[13901]_  : \new_[14025]_ ;
  assign n10960 = \new_[18467]_  ? \new_[14918]_  : \new_[13969]_ ;
  assign n11280 = \new_[18659]_  ? \new_[13902]_  : \new_[14641]_ ;
  assign n10875 = \new_[18679]_  ? \new_[13897]_  : \new_[14072]_ ;
  assign n10870 = \new_[18371]_  ? \new_[13904]_  : \new_[14736]_ ;
  assign n10990 = \new_[18478]_  ? \new_[13897]_  : \new_[14099]_ ;
  assign n10980 = \new_[18473]_  ? \new_[14881]_  : \new_[14114]_ ;
  assign n10505 = \new_[18368]_  ? \new_[13901]_  : \new_[14592]_ ;
  assign n11005 = \new_[19155]_  ? \new_[13901]_  : \new_[14102]_ ;
  assign n11000 = \new_[19507]_  ? \new_[13906]_  : \new_[14105]_ ;
  assign n12775 = \new_[18734]_  ? \new_[14881]_  : \new_[13972]_ ;
  assign n10975 = \new_[19295]_  ? \new_[13894]_  : \new_[14743]_ ;
  assign n11990 = \new_[18250]_  ? \new_[13906]_  : \new_[14599]_ ;
  assign n10655 = \new_[11343]_  ? \new_[14878]_  : \new_[16543]_ ;
  assign n11555 = \new_[13918]_  ? \new_[15486]_  : \new_[18561]_ ;
  assign n11530 = \new_[13919]_  ? \new_[15488]_  : \new_[18249]_ ;
  assign n13110 = \new_[18689]_  ? \new_[13897]_  : \new_[16231]_ ;
  assign n13080 = \new_[19506]_  ? \new_[13902]_  : \new_[15860]_ ;
  assign n11525 = \new_[13921]_  ? \new_[15486]_  : \new_[19284]_ ;
  assign n11535 = \new_[18265]_  ? \new_[13908]_  : \new_[16169]_ ;
  assign n11540 = \new_[18268]_  ? \new_[13898]_  : \new_[15809]_ ;
  assign n13115 = \new_[18832]_  ? \new_[13897]_  : \new_[16233]_ ;
  assign n11545 = \new_[18739]_  ? \new_[13909]_  : \new_[16232]_ ;
  assign n11560 = \new_[13924]_  ? \new_[15489]_  : \new_[19436]_ ;
  assign n10660 = \new_[11344]_  ^ \new_[14878]_ ;
  assign n10345 = \new_[18439]_  ? \new_[13907]_  : \new_[14760]_ ;
  assign n11605 = \new_[18379]_  ? \new_[13894]_  : \new_[14763]_ ;
  assign n11830 = \new_[18538]_  ? \new_[13838]_  : \new_[14758]_ ;
  assign n11675 = \new_[17828]_  ? \new_[13894]_  : \new_[14778]_ ;
  assign n11805 = \new_[18688]_  ? \new_[13900]_  : \new_[14121]_ ;
  assign n11610 = \new_[17988]_  ? \new_[13898]_  : \new_[14230]_ ;
  assign n11575 = \new_[19417]_  ? \new_[13898]_  : \new_[14793]_ ;
  assign n11565 = \new_[18754]_  ? \new_[13897]_  : \new_[16557]_ ;
  assign n11880 = \new_[19127]_  ? \new_[13896]_  : \new_[14178]_ ;
  assign n11885 = \new_[19419]_  ? \new_[13903]_  : \new_[14826]_ ;
  assign n11865 = \new_[19451]_  ? \new_[13900]_  : \new_[14756]_ ;
  assign n11845 = \new_[18097]_  ? \new_[13907]_  : \new_[14120]_ ;
  assign n11800 = \new_[19067]_  ? \new_[13898]_  : \new_[14757]_ ;
  assign n11385 = \new_[18766]_  ? \new_[14916]_  : \new_[14119]_ ;
  assign n11580 = \new_[18196]_  ? \new_[13894]_  : \new_[14117]_ ;
  assign n11585 = \new_[17986]_  ? \new_[13838]_  : \new_[14822]_ ;
  assign n11355 = \new_[17859]_  ? \new_[13905]_  : \new_[14759]_ ;
  assign n11590 = \new_[19424]_  ? \new_[14916]_  : \new_[14164]_ ;
  assign n12865 = \new_[19860]_  ? \new_[13908]_  : \new_[14125]_ ;
  assign n10395 = \new_[19589]_  ? \new_[13838]_  : \new_[13826]_ ;
  assign n11600 = \new_[18208]_  ? \new_[13897]_  : \new_[14126]_ ;
  assign n10270 = \new_[19837]_  ? \new_[13900]_  : \new_[14116]_ ;
  assign n10305 = \new_[18420]_  ? \new_[13911]_  : \new_[14827]_ ;
  assign n10315 = \new_[19431]_  ? \new_[13838]_  : \new_[14764]_ ;
  assign n10325 = \new_[17836]_  ? \new_[13900]_  : \new_[14131]_ ;
  assign n10295 = \new_[18727]_  ? \new_[13898]_  : \new_[14127]_ ;
  assign n11615 = \new_[19130]_  ? \new_[13899]_  : \new_[14765]_ ;
  assign n13015 = \new_[19001]_  ? \new_[14916]_  : \new_[14813]_ ;
  assign n13050 = \new_[17987]_  ? \new_[13911]_  : \new_[14766]_ ;
  assign n13125 = \new_[19638]_  ? \new_[13838]_  : \new_[14831]_ ;
  assign n13120 = \new_[18850]_  ? \new_[13905]_  : \new_[14168]_ ;
  assign n13100 = \new_[18447]_  ? \new_[13896]_  : \new_[14145]_ ;
  assign n13085 = \new_[18454]_  ? \new_[13907]_  : \new_[14819]_ ;
  assign n13030 = \new_[19429]_  ? \new_[14878]_  : \new_[14130]_ ;
  assign n12970 = \new_[18333]_  ? \new_[14881]_  : \new_[14177]_ ;
  assign n12965 = \new_[18919]_  ? \new_[13900]_  : \new_[14162]_ ;
  assign n11645 = \new_[19184]_  ? \new_[13909]_  : \new_[14133]_ ;
  assign n12990 = \new_[19621]_  ? \new_[13899]_  : \new_[14157]_ ;
  assign n12655 = \new_[18605]_  ? \new_[13913]_  : \new_[13829]_ ;
  assign n11650 = \new_[18091]_  ? \new_[13901]_  : \new_[14134]_ ;
  assign n11655 = \new_[19628]_  ? \new_[13896]_  : \new_[14824]_ ;
  assign n11660 = \new_[17809]_  ? \new_[13912]_  : \new_[14171]_ ;
  assign n11665 = \new_[18813]_  ? \new_[14878]_  : \new_[14144]_ ;
  assign n11860 = \new_[19866]_  ? \new_[13913]_  : \new_[14815]_ ;
  assign n11930 = \new_[19701]_  ? \new_[13901]_  : \new_[14212]_ ;
  assign n11940 = \new_[18154]_  ? \new_[13907]_  : \new_[14153]_ ;
  assign n11925 = \new_[19633]_  ? \new_[13900]_  : \new_[14167]_ ;
  assign n11910 = \new_[19040]_  ? \new_[14918]_  : \new_[14776]_ ;
  assign n11915 = \new_[18829]_  ? \new_[13899]_  : \new_[14135]_ ;
  assign n11920 = \new_[19676]_  ? \new_[13895]_  : \new_[14154]_ ;
  assign n11670 = \new_[19651]_  ? \new_[13896]_  : \new_[14118]_ ;
  assign n11835 = \new_[18564]_  ? \new_[13896]_  : \new_[14777]_ ;
  assign n11890 = \new_[19836]_  ? \new_[13896]_  : \new_[14174]_ ;
  assign n11680 = \new_[17923]_  ? \new_[13899]_  : \new_[14829]_ ;
  assign n11900 = \new_[18728]_  ? \new_[14878]_  : \new_[14779]_ ;
  assign n11875 = \new_[19128]_  ? \new_[13904]_  : \new_[14798]_ ;
  assign n11840 = \new_[18003]_  ? \new_[13839]_  : \new_[14169]_ ;
  assign n11850 = \new_[18824]_  ? \new_[13894]_  : \new_[14170]_ ;
  assign n11730 = \new_[17937]_  ? \new_[13899]_  : \new_[14176]_ ;
  assign n11685 = \new_[18658]_  ? \new_[13902]_  : \new_[13828]_ ;
  assign n11810 = \new_[18690]_  ? \new_[13895]_  : \new_[14781]_ ;
  assign n11690 = \new_[19068]_  ? \new_[14918]_  : \new_[14137]_ ;
  assign n11825 = \new_[18616]_  ? \new_[13899]_  : \new_[16341]_ ;
  assign n11695 = \new_[17970]_  ? \new_[14920]_  : \new_[14782]_ ;
  assign n11635 = \new_[19851]_  ? \new_[13838]_  : \new_[13926]_ ;
  assign n11700 = \new_[19351]_  ? \new_[13838]_  : \new_[14810]_ ;
  assign n10335 = \new_[19239]_  ? \new_[14944]_  : \new_[14784]_ ;
  assign n10365 = \new_[19813]_  ? \new_[14920]_  : \new_[14762]_ ;
  assign n10390 = \new_[18087]_  ? \new_[13896]_  : \new_[14811]_ ;
  assign n10385 = \new_[19786]_  ? \new_[14919]_  : \new_[14830]_ ;
  assign n10370 = \new_[18407]_  ? \new_[13902]_  : \new_[14787]_ ;
  assign n10275 = \new_[17885]_  ? \new_[13894]_  : \new_[14156]_ ;
  assign n10310 = \new_[18950]_  ? \new_[13838]_  : \new_[14825]_ ;
  assign n10330 = \new_[19147]_  ? \new_[13838]_  : \new_[14184]_ ;
  assign n13020 = \new_[19574]_  ? \new_[13900]_  : \new_[14186]_ ;
  assign n10300 = \new_[18751]_  ? \new_[14944]_  : \new_[14182]_ ;
  assign n11715 = \new_[19632]_  ? \new_[13894]_  : \new_[14789]_ ;
  assign n12725 = \new_[19150]_  ? \new_[13908]_  : \new_[14834]_ ;
  assign n13060 = \new_[19548]_  ? \new_[13838]_  : \new_[14833]_ ;
  assign n13105 = \new_[19104]_  ? \new_[13894]_  : \new_[14181]_ ;
  assign n13010 = \new_[19778]_  ? \new_[13902]_  : \new_[14180]_ ;
  assign n11725 = \new_[19207]_  ? \new_[13911]_  : \new_[14142]_ ;
  assign n13000 = \new_[19122]_  ? \new_[13897]_  : \new_[14179]_ ;
  assign n12805 = \new_[18318]_  ? \new_[13904]_  : \new_[14175]_ ;
  assign n12950 = \new_[18374]_  ? \new_[13908]_  : \new_[14183]_ ;
  assign n12995 = \new_[18535]_  ? \new_[13838]_  : \new_[14159]_ ;
  assign n12975 = \new_[18933]_  ? \new_[13911]_  : \new_[14115]_ ;
  assign n12930 = \new_[18746]_  ? \new_[13898]_  : \new_[14797]_ ;
  assign n12945 = \new_[18918]_  ? \new_[13904]_  : \new_[16332]_ ;
  assign n11755 = \new_[18970]_  ? \new_[13903]_  : \new_[16344]_ ;
  assign n12790 = \new_[18417]_  ? \new_[13913]_  : \new_[14770]_ ;
  assign n11760 = \new_[18533]_  ? \new_[13905]_  : \new_[14799]_ ;
  assign n12935 = \new_[18830]_  ? \new_[13902]_  : \new_[14821]_ ;
  assign n12825 = \new_[17995]_  ? \new_[13895]_  : \new_[14800]_ ;
  assign n12875 = \new_[18095]_  ? \new_[13899]_  : \new_[14166]_ ;
  assign n11765 = \new_[18015]_  ? \new_[13913]_  : \new_[14165]_ ;
  assign n12915 = \new_[19827]_  ? \new_[13910]_  : \new_[14237]_ ;
  assign n12925 = \new_[18551]_  ? \new_[13902]_  : \new_[14820]_ ;
  assign n12890 = \new_[18683]_  ? \new_[13899]_  : \new_[14147]_ ;
  assign n11770 = \new_[18207]_  ? \new_[13904]_  : \new_[14148]_ ;
  assign n12880 = \new_[18772]_  ? \new_[13838]_  : \new_[14161]_ ;
  assign n11775 = \new_[19262]_  ? \new_[13903]_  : \new_[14801]_ ;
  assign n12810 = \new_[18663]_  ? \new_[13902]_  : \new_[14802]_ ;
  assign n12845 = \new_[18645]_  ? \new_[13906]_  : \new_[14163]_ ;
  assign n12850 = \new_[18240]_  ? \new_[13904]_  : \new_[14817]_ ;
  assign n11780 = \new_[18797]_  ? \new_[13838]_  : \new_[14803]_ ;
  assign n12815 = \new_[19745]_  ? \new_[13894]_  : \new_[14804]_ ;
  assign n12440 = \new_[18211]_  ? \new_[13910]_  : \new_[13840]_ ;
  assign n12710 = \new_[18556]_  ? \new_[13896]_  : \new_[14149]_ ;
  assign n12730 = \new_[19698]_  ? \new_[13910]_  : \new_[14150]_ ;
  assign n11785 = \new_[18990]_  ? \new_[13896]_  : \new_[14151]_ ;
  assign n12770 = \new_[19050]_  ? \new_[13904]_  : \new_[14160]_ ;
  assign n12560 = \new_[19316]_  ? \new_[14878]_  : \new_[14816]_ ;
  assign n12610 = \new_[18206]_  ? \new_[13910]_  : \new_[13850]_ ;
  assign n11790 = \new_[18787]_  ? \new_[13904]_  : \new_[16442]_ ;
  assign n10280 = \new_[19856]_  ? \new_[13908]_  : \new_[14805]_ ;
  assign n12155 = \new_[19620]_  ? \new_[13907]_  : \new_[14152]_ ;
  assign n12170 = \new_[19565]_  ? \new_[13904]_  : \new_[14806]_ ;
  assign n11795 = \new_[17835]_  ? \new_[13905]_  : \new_[14823]_ ;
  assign n12255 = \new_[18697]_  ? \new_[13896]_  : \new_[14807]_ ;
  assign n12330 = \new_[18424]_  ? \new_[13912]_  : \new_[13936]_ ;
  assign n12220 = \new_[18352]_  ? \new_[13838]_  : \new_[14808]_ ;
  assign n12225 = \new_[18414]_  ? \new_[13902]_  : \new_[16343]_ ;
  assign n12745 = \new_[18648]_  ? \new_[13907]_  : \new_[14771]_ ;
  assign n10405 = \new_[18426]_  ? \new_[13898]_  : \new_[14138]_ ;
  assign n11710 = \new_[19367]_  ? \new_[13838]_  : \new_[14140]_ ;
  assign n11705 = \new_[19269]_  ? \new_[13904]_  : \new_[14139]_ ;
  assign n11905 = \new_[18875]_  ? \new_[13906]_  : \new_[14775]_ ;
  assign n12980 = \new_[18170]_  ? \new_[13912]_  : \new_[14795]_ ;
  assign n11630 = \new_[17847]_  ? \new_[13899]_  : \new_[14768]_ ;
  assign n10350 = \new_[18767]_  ? \new_[13907]_  : \new_[14158]_ ;
  assign n13005 = \new_[19847]_  ? \new_[13901]_  : \new_[14812]_ ;
  assign n12830 = \new_[18576]_  ? \new_[13899]_  : \new_[14093]_ ;
  assign n12735 = \new_[19613]_  ? \new_[14922]_  : \new_[14769]_ ;
  assign n11815 = \new_[17857]_  ? \new_[14922]_  : \new_[14809]_ ;
  assign n12940 = \new_[18653]_  ? \new_[13905]_  : \new_[14146]_ ;
  assign n11625 = \new_[18644]_  ? \new_[13897]_  : \new_[14216]_ ;
  assign n10375 = \new_[18943]_  ? \new_[14922]_  : \new_[14786]_ ;
  assign n11820 = \new_[19746]_  ? \new_[14921]_  : \new_[14122]_ ;
  assign n13070 = \new_[19468]_  ? \new_[14917]_  : \new_[14129]_ ;
  assign n11750 = \new_[19553]_  ? \new_[14921]_  : \new_[16331]_ ;
  assign n10290 = \new_[18068]_  ? \new_[14878]_  : \new_[14774]_ ;
  assign n11870 = \new_[19675]_  ? \new_[13904]_  : \new_[14136]_ ;
  assign n10265 = \new_[19486]_  ? \new_[14917]_  : \new_[14783]_ ;
  assign n10320 = \new_[18801]_  ? \new_[14944]_  : \new_[14788]_ ;
  assign n10400 = \new_[19161]_  ? \new_[13901]_  : \new_[14124]_ ;
  assign n12985 = \new_[17907]_  ? \new_[13838]_  : \new_[14794]_ ;
  assign n11570 = \new_[19708]_  ? \new_[13838]_  : \new_[14173]_ ;
  assign n10285 = \new_[18450]_  ? \new_[13838]_  : \new_[14773]_ ;
  assign n11895 = \new_[17999]_  ? \new_[13901]_  : \new_[14755]_ ;
  assign n10550 = \new_[19868]_  ? \new_[13895]_  : \new_[14123]_ ;
  assign n11745 = \new_[19190]_  ? \new_[13899]_  : \new_[16558]_ ;
  assign n11595 = \new_[18955]_  ? \new_[14944]_  : \new_[14155]_ ;
  assign n13130 = \new_[19770]_  ? \new_[14917]_  : \new_[14767]_ ;
  assign n11740 = \new_[18805]_  ? \new_[13901]_  : \new_[14792]_ ;
  assign n12705 = \new_[18629]_  ? \new_[13904]_  : \new_[16030]_ ;
  assign n11855 = \new_[19619]_  ? \new_[14878]_  : \new_[14172]_ ;
  assign n11935 = \new_[18451]_  ? \new_[13906]_  : \new_[14828]_ ;
  assign n11640 = \new_[18991]_  ? \new_[13904]_  : \new_[14132]_ ;
  assign n10340 = \new_[18582]_  ? \new_[13838]_  : \new_[14761]_ ;
  assign n10380 = \new_[19575]_  ? \new_[14921]_  : \new_[16320]_ ;
  assign n11735 = \new_[18127]_  ? \new_[14917]_  : \new_[14143]_ ;
  assign n11720 = \new_[18486]_  ? \new_[14878]_  : \new_[14791]_ ;
  assign n13090 = \new_[18737]_  ? \new_[14921]_  : \new_[14790]_ ;
  assign n13025 = \new_[19072]_  ? \new_[14922]_  : \new_[14141]_ ;
  assign n12955 = \new_[19365]_  ? \new_[13839]_  : \new_[14835]_ ;
  assign n12960 = \new_[18340]_  ? \new_[13895]_  : \new_[14796]_ ;
  assign n12130 = \new_[19609]_  ? \new_[13897]_  : \new_[14772]_ ;
  assign n11620 = \new_[18892]_  ? \new_[13905]_  : \new_[14128]_ ;
  assign n13095 = \new_[19705]_  ? \new_[14922]_  : \new_[14185]_ ;
  assign n10665 = \new_[11345]_  ? \new_[14878]_  : \new_[15939]_ ;
  assign n12530 = n17080 ? \new_[14878]_  : \new_[16884]_ ;
  assign n10670 = n17040 ? \new_[14878]_  : \new_[11343]_ ;
  assign \new_[13117]_  = ~\new_[14229]_  & ~\new_[15359]_ ;
  assign \new_[13118]_  = ~\new_[15276]_  & ~\new_[14229]_ ;
  assign \new_[13119]_  = ~\new_[13719]_ ;
  assign \new_[13120]_  = ~\new_[15784]_  | ~\new_[13759]_ ;
  assign \new_[13121]_  = ~\new_[14229]_  & ~\new_[15563]_ ;
  assign \new_[13122]_  = ~\new_[10876]_  | ~\new_[14287]_ ;
  assign \new_[13123]_  = ~\new_[13577]_ ;
  assign n16910 = pci_target_unit_del_sync_comp_rty_exp_reg_reg;
  assign \new_[13125]_  = ~\new_[20065]_  | ~\new_[13701]_  | ~\new_[19742]_ ;
  assign \new_[13126]_  = ~\new_[17025]_  | ~\new_[14292]_  | ~\new_[17028]_  | ~\new_[18729]_ ;
  assign \new_[13127]_  = ~\new_[13784]_  & ~\new_[19906]_ ;
  assign \new_[13128]_  = ~\new_[13782]_  & (~\new_[4896]_  | ~\new_[19906]_ );
  assign \new_[13129]_  = \wbm_adr_o[26]  ? \new_[15502]_  : \new_[14194]_ ;
  assign \new_[13130]_  = ~\new_[20397]_ ;
  assign \new_[13131]_  = ~\new_[13789]_  & ~\new_[19906]_ ;
  assign \new_[13132]_  = \wbm_adr_o[29]  ? \new_[15502]_  : \new_[14198]_ ;
  assign n12000 = \new_[10389]_  ? \new_[15633]_  : \new_[14201]_ ;
  assign \new_[13134]_  = \\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2] ;
  assign \new_[13135]_  = ~\new_[17318]_  | ~\new_[17101]_  | ~\new_[14780]_  | ~\new_[17031]_ ;
  assign \new_[13136]_  = ~\new_[13804]_  & ~\new_[15451]_ ;
  assign n10565 = ~\new_[13800]_  & ~\new_[15836]_ ;
  assign \new_[13138]_  = ~\new_[13804]_  & ~\new_[17019]_ ;
  assign n10575 = \new_[13804]_  & \new_[11326]_ ;
  assign n10580 = \new_[13804]_  & \new_[11327]_ ;
  assign \new_[13141]_  = ~\new_[13804]_  | ~\new_[19194]_ ;
  assign \new_[13142]_  = ~\new_[13804]_  | ~\new_[19410]_ ;
  assign n10585 = \new_[13804]_  & \new_[11328]_ ;
  assign \new_[13144]_  = ~\new_[13804]_  | ~\new_[10497]_ ;
  assign n10355 = \new_[13804]_  & \new_[11282]_ ;
  assign \new_[13146]_  = ~\new_[13804]_  & ~\new_[15619]_ ;
  assign \new_[13147]_  = ~\new_[13803]_  & (~\new_[18791]_  | ~\new_[19906]_ );
  assign n10570 = ~\new_[13620]_ ;
  assign \new_[13149]_  = \wbm_adr_o[31]  ? \new_[15502]_  : \new_[13815]_ ;
  assign \new_[13150]_  = ~configuration_set_pci_err_cs_bit8_reg;
  assign \new_[13151]_  = ~\new_[15050]_  | ~\new_[15323]_  | ~\new_[15475]_  | ~\new_[13853]_ ;
  assign \new_[13152]_  = ~\new_[20105]_  | ~\new_[13690]_  | ~\new_[17312]_ ;
  assign \new_[13153]_  = ~\new_[19887]_  | ~\new_[19948]_ ;
  assign \new_[13154]_  = \new_[20505]_  & \new_[15015]_ ;
  assign \new_[13155]_  = ~\new_[15042]_  | ~\new_[15291]_  | ~\new_[15455]_  | ~\new_[13842]_ ;
  assign n13065 = ~\new_[14924]_  | ~\new_[13781]_ ;
  assign \new_[13157]_  = ~\new_[13762]_  & (~\new_[14908]_  | ~\new_[16603]_ );
  assign \new_[13158]_  = wishbone_slave_unit_pci_initiator_if_del_write_req_reg;
  assign n10590 = ~\new_[13700]_  | (~\new_[15003]_  & ~\new_[14242]_ );
  assign \new_[13160]_  = ~\new_[13721]_  & ~\new_[13699]_ ;
  assign n13075 = \new_[13872]_  ? \new_[15484]_  : \new_[18279]_ ;
  assign n10595 = \new_[10392]_  ? \new_[15633]_  : \new_[13836]_ ;
  assign n13420 = \wbm_adr_o[2]  ? \new_[14219]_  : \new_[12022]_ ;
  assign n15035 = \wbm_adr_o[30]  ? \new_[14218]_  : \new_[12423]_ ;
  assign n13425 = \wbm_adr_o[31]  ? \new_[14218]_  : \new_[12023]_ ;
  assign n15005 = \wbm_adr_o[3]  ? \new_[14996]_  : \new_[12417]_ ;
  assign n13430 = \wbm_adr_o[4]  ? \new_[14996]_  : \new_[12024]_ ;
  assign n15030 = \wbm_adr_o[5]  ? \new_[14219]_  : \new_[12422]_ ;
  assign n13435 = \wbm_adr_o[6]  ? \new_[14219]_  : \new_[12025]_ ;
  assign n14910 = \wbm_adr_o[7]  ? \new_[14219]_  : \new_[12383]_ ;
  assign n13440 = \wbm_adr_o[8]  ? \new_[14219]_  : \new_[12026]_ ;
  assign n14930 = \wbm_adr_o[9]  ? \new_[14219]_  : \new_[12401]_ ;
  assign n14970 = \new_[18909]_  ? \new_[14219]_  : \new_[12410]_ ;
  assign n14980 = \new_[19219]_  ? \new_[14219]_  : \new_[12412]_ ;
  assign n14995 = \new_[19116]_  ? \new_[14219]_  : \new_[12415]_ ;
  assign n15000 = \new_[19573]_  ? \new_[14996]_  : \new_[12416]_ ;
  assign n13445 = \wbm_dat_o[0]  ? \new_[14218]_  : \new_[12027]_ ;
  assign n14985 = \wbm_dat_o[10]  ? \new_[14219]_  : \new_[12413]_ ;
  assign n13450 = \wbm_dat_o[11]  ? \new_[14218]_  : \new_[12028]_ ;
  assign n14990 = \wbm_dat_o[12]  ? \new_[14218]_  : \new_[12414]_ ;
  assign n13455 = \wbm_dat_o[13]  ? \new_[14218]_  : \new_[12029]_ ;
  assign n14965 = \wbm_dat_o[14]  ? \new_[14219]_  : \new_[12409]_ ;
  assign n13460 = \wbm_dat_o[15]  ? \new_[14219]_  : \new_[12030]_ ;
  assign n14975 = \wbm_dat_o[16]  ? \new_[14219]_  : \new_[12411]_ ;
  assign n13465 = \wbm_dat_o[17]  ? \new_[14219]_  : \new_[12031]_ ;
  assign n14940 = \wbm_dat_o[18]  ? \new_[14219]_  : \new_[12404]_ ;
  assign n13470 = \wbm_dat_o[19]  ? \new_[14219]_  : \new_[12032]_ ;
  assign n14945 = \wbm_dat_o[1]  ? \new_[14219]_  : \new_[12405]_ ;
  assign n14950 = \wbm_dat_o[20]  ? \new_[14219]_  : \new_[12406]_ ;
  assign n13475 = \wbm_dat_o[21]  ? \new_[14219]_  : \new_[12033]_ ;
  assign n14955 = \wbm_dat_o[22]  ? \new_[14219]_  : \new_[12407]_ ;
  assign n14635 = \wbm_dat_o[23]  ? \new_[14219]_  : \new_[12323]_ ;
  assign n14715 = \wbm_dat_o[24]  ? \new_[14219]_  : \new_[12340]_ ;
  assign n13480 = \wbm_dat_o[25]  ? \new_[14218]_  : \new_[12034]_ ;
  assign n14830 = \wbm_dat_o[26]  ? \new_[14218]_  : \new_[12366]_ ;
  assign n14835 = \wbm_dat_o[27]  ? \new_[14218]_  : \new_[12367]_ ;
  assign n13165 = \wbm_dat_o[28]  ? \new_[14218]_  : \new_[11960]_ ;
  assign n13485 = \wbm_dat_o[29]  ? \new_[14218]_  : \new_[12035]_ ;
  assign n14545 = \wbm_dat_o[30]  ? \new_[14219]_  : \new_[12305]_ ;
  assign n13490 = \wbm_dat_o[31]  ? \new_[14996]_  : \new_[12036]_ ;
  assign n13495 = \wbm_dat_o[3]  ? \new_[14996]_  : \new_[12037]_ ;
  assign n14575 = \wbm_dat_o[4]  ? \new_[14219]_  : \new_[12311]_ ;
  assign n14565 = \wbm_dat_o[5]  ? \new_[14996]_  : \new_[12309]_ ;
  assign n13500 = \wbm_dat_o[7]  ? \new_[14219]_  : \new_[12038]_ ;
  assign n14540 = \wbm_dat_o[8]  ? \new_[14219]_  : \new_[12304]_ ;
  assign n14550 = \wbm_dat_o[9]  ? \new_[14219]_  : \new_[12306]_ ;
  assign n14500 = \wbm_dat_o[2]  ? \new_[14219]_  : \new_[12296]_ ;
  assign \new_[13208]_  = ~\new_[19965]_ ;
  assign n14570 = \wbm_dat_o[6]  ? \new_[14219]_  : \new_[12310]_ ;
  assign \new_[13210]_  = \wbm_adr_o[27]  ? \new_[15502]_  : \new_[14233]_ ;
  assign n13370 = \new_[10390]_  ? \new_[15633]_  : \new_[14234]_ ;
  assign \new_[13212]_  = ~\new_[14923]_  | ~\new_[15086]_  | ~\new_[15530]_  | ~\new_[15514]_ ;
  assign \new_[13213]_  = pci_target_unit_wishbone_master_wb_read_done_out_reg;
  assign \new_[13214]_  = \new_[13820]_  | \new_[17476]_ ;
  assign \new_[13215]_  = ~pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg;
  assign \new_[13216]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[0] ;
  assign \new_[13217]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1] ;
  assign \new_[13218]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[0] ;
  assign \new_[13219]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0] ;
  assign n16930 = pci_target_unit_del_sync_req_done_reg_reg;
  assign \new_[13221]_  = \\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1] ;
  assign \new_[13222]_  = \\pci_target_unit_pci_target_if_strd_address_reg[2] ;
  assign \new_[13223]_  = \new_[14261]_  ? \new_[17323]_  : \new_[16951]_ ;
  assign n14530 = ~\new_[15866]_  | ~\new_[13822]_ ;
  assign n13510 = \new_[10371]_  ? \new_[14243]_  : \new_[12040]_ ;
  assign n14430 = \new_[5045]_  ? \new_[14242]_  : \new_[12268]_ ;
  assign n14425 = \new_[5046]_  ? \new_[14242]_  : \new_[12267]_ ;
  assign n13180 = \new_[4174]_  ? \new_[14258]_  : \new_[11963]_ ;
  assign n14265 = \new_[9902]_  ? \new_[14242]_  : \new_[12198]_ ;
  assign n13150 = \new_[4178]_  ? \new_[14243]_  : \new_[11957]_ ;
  assign n13515 = \new_[4175]_  ? \new_[14243]_  : \new_[12042]_ ;
  assign n13140 = \new_[4345]_  ? \new_[14258]_  : \new_[11955]_ ;
  assign n13520 = \new_[4226]_  ? \new_[14242]_  : \new_[12043]_ ;
  assign n13525 = \new_[4228]_  ? \new_[14242]_  : \new_[12044]_ ;
  assign n13530 = \new_[4229]_  ? \new_[14242]_  : \new_[12045]_ ;
  assign n14405 = \new_[4210]_  ? \new_[14242]_  : \new_[12259]_ ;
  assign n13535 = \new_[4211]_  ? \new_[14258]_  : \new_[12046]_ ;
  assign n13540 = \new_[4180]_  ? \new_[14242]_  : \new_[12047]_ ;
  assign n13545 = \new_[4212]_  ? \new_[14242]_  : \new_[12048]_ ;
  assign n14485 = \new_[4213]_  ? \new_[14242]_  : \new_[12287]_ ;
  assign n13550 = \new_[4214]_  ? \new_[14242]_  : \new_[12049]_ ;
  assign n13555 = \new_[4215]_  ? \new_[14258]_  : \new_[12050]_ ;
  assign n13560 = \new_[4260]_  ? \new_[14243]_  : \new_[12051]_ ;
  assign n13330 = \new_[4216]_  ? \new_[14258]_  : \new_[12004]_ ;
  assign n13565 = \new_[4265]_  ? \new_[14242]_  : \new_[12052]_ ;
  assign n13570 = \new_[4217]_  ? \new_[14242]_  : \new_[12053]_ ;
  assign n13575 = \new_[4181]_  ? \new_[14243]_  : \new_[12054]_ ;
  assign n13280 = \new_[4182]_  ? \new_[14243]_  : \new_[11993]_ ;
  assign n13580 = \new_[4456]_  ? \new_[14242]_  : \new_[12055]_ ;
  assign n13585 = \new_[4268]_  ? \new_[14242]_  : \new_[12056]_ ;
  assign n13270 = \new_[4183]_  ? \new_[14242]_  : \new_[11991]_ ;
  assign n13265 = \new_[4184]_  ? \new_[14258]_  : \new_[11990]_ ;
  assign n13590 = \new_[4185]_  ? \new_[14242]_  : \new_[12058]_ ;
  assign n13595 = \new_[4186]_  ? \new_[14243]_  : \new_[12059]_ ;
  assign n13245 = \new_[4261]_  ? \new_[14258]_  : \new_[11986]_ ;
  assign n13255 = \new_[4130]_  ? \new_[14258]_  : \new_[11988]_ ;
  assign n13600 = \new_[4187]_  ? \new_[14258]_  : \new_[12060]_ ;
  assign n13250 = \new_[4188]_  ? \new_[14242]_  : \new_[11987]_ ;
  assign n13605 = \new_[4189]_  ? \new_[14243]_  : \new_[12061]_ ;
  assign n13220 = \new_[4190]_  ? \new_[14242]_  : \new_[11981]_ ;
  assign n13615 = \new_[4191]_  ? \new_[14242]_  : \new_[12063]_ ;
  assign n13235 = \new_[4192]_  ? \new_[14242]_  : \new_[11984]_ ;
  assign n13610 = \new_[4218]_  ? \new_[14258]_  : \new_[12062]_ ;
  assign n13620 = \new_[5043]_  ? \new_[14243]_  : \new_[12064]_ ;
  assign n13135 = \new_[5090]_  ? \new_[14242]_  : \new_[11954]_ ;
  assign n13625 = \new_[5044]_  ? \new_[14242]_  : \new_[12065]_ ;
  assign n13630 = \new_[5038]_  ? \new_[14243]_  : \new_[12066]_ ;
  assign n13635 = \new_[4963]_  ? \new_[14258]_  : \new_[12067]_ ;
  assign n13185 = \new_[5039]_  ? \new_[14243]_  : \new_[11964]_ ;
  assign n13640 = \new_[4964]_  ? \new_[14258]_  : \new_[12068]_ ;
  assign n14675 = \new_[5040]_  ? \new_[14242]_  : \new_[12331]_ ;
  assign n13645 = \new_[5012]_  ? \new_[14243]_  : \new_[12069]_ ;
  assign n13155 = \new_[4965]_  ? \new_[14242]_  : \new_[11958]_ ;
  assign n13650 = \new_[4966]_  ? \new_[14242]_  : \new_[12070]_ ;
  assign n15020 = \new_[5009]_  ? \new_[14242]_  : \new_[12420]_ ;
  assign n13655 = \new_[4967]_  ? \new_[14242]_  : \new_[12071]_ ;
  assign n15185 = \new_[4968]_  ? \new_[14243]_  : \new_[12509]_ ;
  assign n13660 = \new_[4969]_  ? \new_[14242]_  : \new_[12072]_ ;
  assign n15245 = \new_[5010]_  ? \new_[14242]_  : \new_[12532]_ ;
  assign n13665 = \new_[4896]_  ? \new_[14242]_  : \new_[12073]_ ;
  assign n15260 = \new_[4970]_  ? \new_[14242]_  : \new_[12536]_ ;
  assign n13670 = \new_[4971]_  ? \new_[14258]_  : \new_[12074]_ ;
  assign n15215 = \new_[4972]_  ? \new_[14242]_  : \new_[12524]_ ;
  assign n13675 = \new_[5008]_  ? \new_[14242]_  : \new_[12075]_ ;
  assign n15210 = \new_[5011]_  ? \new_[14243]_  : \new_[12523]_ ;
  assign n13680 = \new_[18791]_  ? \new_[14243]_  : \new_[12076]_ ;
  assign n15180 = \new_[5041]_  ? \new_[14243]_  : \new_[12508]_ ;
  assign n13685 = \new_[4974]_  ? \new_[14258]_  : \new_[12077]_ ;
  assign n15165 = \new_[4962]_  ? \new_[14242]_  : \new_[12495]_ ;
  assign n13690 = \new_[4975]_  ? \new_[14242]_  : \new_[12078]_ ;
  assign n13695 = \new_[4976]_  ? \new_[14242]_  : \new_[12079]_ ;
  assign n13700 = \new_[5042]_  ? \new_[14242]_  : \new_[12080]_ ;
  assign n15160 = \new_[4977]_  ? \new_[14258]_  : \new_[12494]_ ;
  assign n14420 = \new_[5047]_  ? \new_[14242]_  : \new_[12266]_ ;
  assign \new_[13295]_  = ~\new_[13841]_  | ~\new_[17383]_ ;
  assign \new_[13296]_  = ~\new_[13841]_  | ~\new_[17080]_ ;
  assign \new_[13297]_  = ~\new_[13841]_  | ~\new_[20143]_ ;
  assign \new_[13298]_  = ~\new_[15791]_  | ~\new_[17033]_  | ~\new_[20129]_  | ~\new_[16078]_ ;
  assign \new_[13299]_  = ~\new_[14941]_  | ~\new_[14960]_  | ~\new_[15035]_  | ~\new_[15689]_ ;
  assign n13705 = ~\new_[13851]_  | (~\new_[14932]_  & ~\new_[12081]_ );
  assign n13710 = ~\new_[13851]_  | (~\new_[12082]_  & ~\new_[14932]_ );
  assign n13920 = \new_[14408]_  ? \new_[15484]_  : \new_[18708]_ ;
  assign n14665 = \new_[14419]_  ? \new_[15273]_  : \new_[18922]_ ;
  assign n13720 = \new_[14297]_  ? \new_[15488]_  : \new_[18163]_ ;
  assign n13900 = \new_[14335]_  ? \new_[15488]_  : \new_[18543]_ ;
  assign n14215 = \new_[14295]_  ? \new_[15590]_  : \new_[19730]_ ;
  assign n13875 = \new_[14326]_  ? \new_[15486]_  : \new_[19397]_ ;
  assign n14315 = \new_[14319]_  ? \new_[15486]_  : \new_[18461]_ ;
  assign n13965 = \new_[14350]_  ? \new_[15592]_  : \new_[19496]_ ;
  assign n13915 = \new_[14346]_  ? \new_[15590]_  : \new_[18626]_ ;
  assign n13300 = \new_[14301]_  ? \new_[15488]_  : \new_[18433]_ ;
  assign n15140 = \new_[14304]_  ? \new_[15275]_  : \new_[18497]_ ;
  assign n13910 = \new_[14329]_  ? \new_[15273]_  : \new_[19402]_ ;
  assign n15225 = \new_[14334]_  ? \new_[15590]_  : \new_[18706]_ ;
  assign n14335 = \new_[14372]_  ? \new_[15489]_  : \new_[17953]_ ;
  assign n14365 = \new_[14328]_  ? \new_[15494]_  : \new_[19280]_ ;
  assign n13870 = \new_[14307]_  ? \new_[15493]_  : \new_[19134]_ ;
  assign n14670 = \new_[14422]_  ? \new_[15493]_  : \new_[18549]_ ;
  assign n14295 = \new_[14296]_  ? \new_[15273]_  : \new_[19717]_ ;
  assign n13745 = \new_[14311]_  ? \new_[15491]_  : \new_[19861]_ ;
  assign n14290 = \new_[14314]_  ? \new_[15488]_  : \new_[18398]_ ;
  assign n13740 = \new_[14305]_  ? \new_[15485]_  : \new_[18235]_ ;
  assign n14325 = \new_[14315]_  ? \new_[15488]_  : \new_[19281]_ ;
  assign n13945 = \new_[14313]_  ? \new_[15590]_  : \new_[18493]_ ;
  assign n14305 = \new_[14316]_  ? \new_[15275]_  : \new_[19359]_ ;
  assign n13320 = \new_[14321]_  ? \new_[15273]_  : \new_[18307]_ ;
  assign n14285 = \new_[14356]_  ? \new_[15485]_  : \new_[18252]_ ;
  assign n15150 = \new_[14318]_  ? \new_[15273]_  : \new_[18849]_ ;
  assign n13295 = \new_[14327]_  ? \new_[15494]_  : \new_[19706]_ ;
  assign n13750 = \new_[14323]_  ? \new_[15484]_  : \new_[19286]_ ;
  assign n13755 = \new_[14325]_  ? \new_[15491]_  : \new_[19290]_ ;
  assign n14345 = \new_[14320]_  ? \new_[15590]_  : \new_[19278]_ ;
  assign n14280 = \new_[14333]_  ? \new_[15486]_  : \new_[18577]_ ;
  assign n13195 = \new_[14302]_  ? \new_[15491]_  : \new_[18912]_ ;
  assign n13930 = \new_[14303]_  ? \new_[15491]_  : \new_[18400]_ ;
  assign n15130 = \new_[14299]_  ? \new_[15493]_  : \new_[18255]_ ;
  assign n13975 = \new_[14399]_  ? \new_[15488]_  : \new_[18527]_ ;
  assign n13865 = \new_[14322]_  ? \new_[15592]_  : \new_[19618]_ ;
  assign n15170 = \new_[14337]_  ? \new_[15590]_  : \new_[19298]_ ;
  assign n15135 = \new_[14341]_  ? \new_[15484]_  : \new_[19508]_ ;
  assign n14630 = \new_[14331]_  ? \new_[15590]_  : \new_[18984]_ ;
  assign n13760 = \new_[14336]_  ? \new_[15489]_  : \new_[18710]_ ;
  assign n14880 = \new_[14338]_  ? \new_[15489]_  : \new_[19076]_ ;
  assign n13765 = \new_[14385]_  ? \new_[15592]_  : \new_[19299]_ ;
  assign n14330 = \new_[14371]_  ? \new_[15495]_  : \new_[18372]_ ;
  assign n13215 = \new_[14364]_  ? \new_[15495]_  : \new_[18466]_ ;
  assign n14390 = \new_[14355]_  ? \new_[15590]_  : \new_[18572]_ ;
  assign n14865 = \new_[14389]_  ? \new_[15273]_  : \new_[18757]_ ;
  assign n15145 = \new_[14348]_  ? \new_[15489]_  : \new_[19401]_ ;
  assign n14875 = \new_[14376]_  ? \new_[15274]_  : \new_[19734]_ ;
  assign n14275 = \new_[14380]_  ? \new_[15590]_  : \new_[19355]_ ;
  assign n13925 = \new_[14345]_  ? \new_[15274]_  : \new_[19387]_ ;
  assign n14640 = \new_[14344]_  ? \new_[15489]_  : \new_[18821]_ ;
  assign n13895 = \new_[14349]_  ? \new_[15489]_  : \new_[18477]_ ;
  assign n14645 = \new_[14343]_  ? \new_[15491]_  : \new_[18761]_ ;
  assign n13815 = \new_[14340]_  ? \new_[15273]_  : \new_[18784]_ ;
  assign n14395 = \new_[14351]_  ? \new_[15488]_  : \new_[18713]_ ;
  assign n14895 = \new_[14342]_  ? \new_[15275]_  : \new_[18269]_ ;
  assign n14660 = \new_[14384]_  ? \new_[15488]_  : \new_[18270]_ ;
  assign n14300 = \new_[14363]_  ? \new_[15488]_  : \new_[18635]_ ;
  assign n14375 = \new_[14386]_  ? \new_[15275]_  : \new_[18853]_ ;
  assign n13795 = \new_[14378]_  ? \new_[15484]_  : \new_[18275]_ ;
  assign n13950 = \new_[14330]_  ? \new_[15495]_  : \new_[18496]_ ;
  assign n13890 = \new_[14370]_  ? \new_[15495]_  : \new_[19379]_ ;
  assign n13805 = \new_[14369]_  ? \new_[15590]_  : \new_[18896]_ ;
  assign n14400 = \new_[14387]_  ? \new_[15488]_  : \new_[18360]_ ;
  assign n14270 = \new_[14391]_  ? \new_[15592]_  : \new_[18652]_ ;
  assign n13820 = \new_[14382]_  ? \new_[15488]_  : \new_[18699]_ ;
  assign n13810 = \new_[14362]_  ? \new_[15486]_  : \new_[18378]_ ;
  assign n13785 = \new_[14353]_  ? \new_[15275]_  : \new_[18625]_ ;
  assign n13840 = \new_[14411]_  ? \new_[15491]_  : \new_[18377]_ ;
  assign n14480 = \new_[14357]_  ? \new_[15488]_  : \new_[18638]_ ;
  assign n13845 = \new_[14407]_  ? \new_[15273]_  : \new_[18051]_ ;
  assign n14250 = \new_[14403]_  ? \new_[15273]_  : \new_[19005]_ ;
  assign n14210 = \new_[14392]_  ? \new_[15489]_  : \new_[19660]_ ;
  assign n13780 = \new_[14359]_  ? \new_[15491]_  : \new_[18273]_ ;
  assign n14000 = \new_[14420]_  ? \new_[15494]_  : \new_[17811]_ ;
  assign n14370 = \new_[14361]_  ? \new_[15485]_  : \new_[18623]_ ;
  assign n13775 = \new_[14358]_  ? \new_[15485]_  : \new_[18702]_ ;
  assign n13315 = \new_[14365]_  ? \new_[15493]_  : \new_[18271]_ ;
  assign n13735 = \new_[14310]_  ? \new_[15493]_  : \new_[18237]_ ;
  assign n13725 = \new_[14300]_  ? \new_[15484]_  : \new_[19550]_ ;
  assign n14415 = \new_[14366]_  ? \new_[15592]_  : \new_[18949]_ ;
  assign n14230 = \new_[14417]_  ? \new_[15491]_  : \new_[18418]_ ;
  assign n13715 = \new_[14324]_  ? \new_[15590]_  : \new_[19356]_ ;
  assign n13880 = \new_[14317]_  ? \new_[15493]_  : \new_[18432]_ ;
  assign n13730 = \new_[14306]_  ? \new_[15493]_  : \new_[19448]_ ;
  assign n13885 = \new_[14414]_  ? \new_[15591]_  : \new_[18431]_ ;
  assign n13325 = \new_[14424]_  ? \new_[15591]_  : \new_[18452]_ ;
  assign n14410 = \new_[14368]_  ? \new_[15486]_  : \new_[18423]_ ;
  assign n13905 = \new_[14377]_  ? \new_[15492]_  : \new_[18465]_ ;
  assign n14380 = \new_[14352]_  ? \new_[15491]_  : \new_[19301]_ ;
  assign n13210 = \new_[14309]_  ? \new_[15486]_  : \new_[19385]_ ;
  assign n14350 = \new_[14298]_  ? \new_[15491]_  : \new_[18283]_ ;
  assign n14245 = \new_[14395]_  ? \new_[15493]_  : \new_[18764]_ ;
  assign n14385 = \new_[14373]_  ? \new_[15484]_  : \new_[18745]_ ;
  assign n15230 = \new_[14410]_  ? \new_[15484]_  : \new_[18482]_ ;
  assign n13800 = \new_[14375]_  ? \new_[15488]_  : \new_[18622]_ ;
  assign n13830 = \new_[14360]_  ? \new_[15488]_  : \new_[18773]_ ;
  assign n13955 = \new_[14383]_  ? \new_[15494]_  : \new_[18494]_ ;
  assign n15200 = \new_[14354]_  ? \new_[15275]_  : \new_[18785]_ ;
  assign n13770 = \new_[14367]_  ? \new_[15488]_  : \new_[18032]_ ;
  assign n13825 = \new_[14381]_  ? \new_[15273]_  : \new_[18364]_ ;
  assign n13960 = \new_[14390]_  ? \new_[15484]_  : \new_[19433]_ ;
  assign n13205 = \new_[14388]_  ? \new_[15484]_  : \new_[18612]_ ;
  assign n14225 = \new_[14426]_  ? \new_[15591]_  : \new_[18500]_ ;
  assign n13850 = \new_[14396]_  ? \new_[15273]_  : \new_[18053]_ ;
  assign n14260 = \new_[14394]_  ? \new_[15275]_  : \new_[18155]_ ;
  assign n13790 = \new_[14401]_  ? \new_[15489]_  : \new_[18274]_ ;
  assign n13990 = \new_[14398]_  ? \new_[15494]_  : \new_[19031]_ ;
  assign n15040 = \new_[14400]_  ? \new_[15484]_  : \new_[18485]_ ;
  assign n14255 = \new_[14402]_  ? \new_[15492]_  : \new_[19556]_ ;
  assign n14340 = \new_[14397]_  ? \new_[15591]_  : \new_[18376]_ ;
  assign n14310 = \new_[14404]_  ? \new_[15273]_  : \new_[17861]_ ;
  assign n14885 = \new_[14405]_  ? \new_[15492]_  : \new_[19384]_ ;
  assign n14360 = \new_[14308]_  ? \new_[15495]_  : \new_[18375]_ ;
  assign n13935 = \new_[14393]_  ? \new_[15492]_  : \new_[19020]_ ;
  assign n13985 = \new_[14406]_  ? \new_[15492]_  : \new_[18974]_ ;
  assign n13835 = \new_[14339]_  ? \new_[15273]_  : \new_[18837]_ ;
  assign n14355 = \new_[14409]_  ? \new_[15273]_  : \new_[18660]_ ;
  assign n13980 = \new_[14332]_  ? \new_[15494]_  : \new_[18344]_ ;
  assign n14220 = \new_[14425]_  ? \new_[15494]_  : \new_[18816]_ ;
  assign n13860 = \new_[14347]_  ? \new_[15274]_  : \new_[19357]_ ;
  assign n13995 = \new_[14413]_  ? \new_[15494]_  : \new_[19554]_ ;
  assign n13275 = \new_[14412]_  ? \new_[15590]_  : \new_[18464]_ ;
  assign n15255 = \new_[14379]_  ? \new_[15274]_  : \new_[18800]_ ;
  assign n14005 = \new_[14423]_  ? \new_[15274]_  : \new_[18712]_ ;
  assign n13940 = \new_[14312]_  ? \new_[15274]_  : \new_[18870]_ ;
  assign n13855 = \new_[14416]_  ? \new_[15489]_  : \new_[19603]_ ;
  assign n14240 = \new_[14415]_  ? \new_[15489]_  : \new_[19605]_ ;
  assign n13240 = \new_[14421]_  ? \new_[15492]_  : \new_[19377]_ ;
  assign n14235 = \new_[14418]_  ? \new_[15492]_  : \new_[19081]_ ;
  assign n15220 = \new_[14374]_  ? \new_[15591]_  : \new_[18866]_ ;
  assign \new_[13434]_  = ~\new_[14964]_  | ~\new_[15357]_  | ~\new_[15463]_  | ~\new_[15522]_ ;
  assign \new_[13435]_  = ~\new_[14963]_  | ~\new_[15357]_  | ~\new_[15462]_  | ~\new_[15519]_ ;
  assign \new_[13436]_  = ~\new_[13710]_ ;
  assign \new_[13437]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1] ;
  assign n14180 = \new_[14559]_  ? \new_[15591]_  : \new_[18316]_ ;
  assign n14445 = \new_[14428]_  ? \new_[15491]_  : \new_[17993]_ ;
  assign n14010 = \new_[14542]_  ? \new_[15591]_  : \new_[17954]_ ;
  assign n14435 = \new_[14429]_  ? \new_[15488]_  : \new_[19661]_ ;
  assign n14015 = \new_[14430]_  ? \new_[15488]_  : \new_[19622]_ ;
  assign n13200 = \new_[14432]_  ? \new_[15488]_  : \new_[19804]_ ;
  assign n14020 = \new_[14433]_  ? \new_[15491]_  : \new_[19244]_ ;
  assign n13190 = \new_[14434]_  ? \new_[15275]_  : \new_[18006]_ ;
  assign n14520 = \new_[14538]_  ? \new_[15488]_  : \new_[18172]_ ;
  assign n14025 = \new_[14437]_  ? \new_[15488]_  : \new_[19642]_ ;
  assign n14490 = \new_[14436]_  ? \new_[15488]_  : \new_[19736]_ ;
  assign n14165 = \new_[14438]_  ? \new_[15485]_  : \new_[18570]_ ;
  assign n14030 = \new_[14440]_  ? \new_[15485]_  : \new_[18662]_ ;
  assign n13145 = \new_[14536]_  ? \new_[15275]_  : \new_[19442]_ ;
  assign n13225 = \new_[14442]_  ? \new_[15485]_  : \new_[18819]_ ;
  assign n14320 = \new_[14443]_  ? \new_[15484]_  : \new_[18005]_ ;
  assign n13285 = \new_[14444]_  ? \new_[15495]_  : \new_[18508]_ ;
  assign n13230 = \new_[14535]_  ? \new_[15488]_  : \new_[18647]_ ;
  assign n13160 = \new_[14445]_  ? \new_[15488]_  : \new_[18524]_ ;
  assign n14620 = \new_[14446]_  ? \new_[15486]_  : \new_[18410]_ ;
  assign n14035 = \new_[14448]_  ? \new_[15493]_  : \new_[18233]_ ;
  assign n15235 = \new_[14449]_  ? \new_[15488]_  : \new_[17862]_ ;
  assign n14170 = \new_[14450]_  ? \new_[15488]_  : \new_[19447]_ ;
  assign n15195 = \new_[14533]_  ? \new_[15488]_  : \new_[19839]_ ;
  assign n14625 = \new_[14532]_  ? \new_[15274]_  : \new_[19060]_ ;
  assign n14805 = \new_[14453]_  ? \new_[15273]_  : \new_[19769]_ ;
  assign n14720 = \new_[14454]_  ? \new_[15488]_  : \new_[18387]_ ;
  assign n14840 = \new_[14455]_  ? \new_[15486]_  : \new_[18841]_ ;
  assign n14855 = \new_[14456]_  ? \new_[15488]_  : \new_[19034]_ ;
  assign n14045 = \new_[14458]_  ? \new_[15488]_  : \new_[19112]_ ;
  assign n14050 = \new_[14459]_  ? \new_[15273]_  : \new_[18957]_ ;
  assign n14825 = \new_[14460]_  ? \new_[15592]_  : \new_[18278]_ ;
  assign n14055 = \new_[14461]_  ? \new_[15486]_  : \new_[18717]_ ;
  assign n14060 = \new_[14462]_  ? \new_[15492]_  : \new_[18442]_ ;
  assign n14800 = \new_[14463]_  ? \new_[15493]_  : \new_[18610]_ ;
  assign n14140 = \new_[14539]_  ? \new_[15493]_  : \new_[18408]_ ;
  assign n14725 = \new_[14464]_  ? \new_[15488]_  : \new_[18858]_ ;
  assign n14815 = \new_[14527]_  ? \new_[15495]_  : \new_[19841]_ ;
  assign n14750 = \new_[14467]_  ? \new_[15591]_  : \new_[19761]_ ;
  assign n14780 = \new_[14468]_  ? \new_[15491]_  : \new_[19646]_ ;
  assign n14795 = \new_[14470]_  ? \new_[15488]_  : \new_[18094]_ ;
  assign n14770 = \new_[14472]_  ? \new_[15489]_  : \new_[18104]_ ;
  assign n14765 = \new_[14473]_  ? \new_[15495]_  : \new_[19426]_ ;
  assign n14705 = \new_[14475]_  ? \new_[15488]_  : \new_[18592]_ ;
  assign n14730 = \new_[14476]_  ? \new_[15273]_  : \new_[19465]_ ;
  assign n14740 = \new_[14478]_  ? \new_[15485]_  : \new_[19492]_ ;
  assign n14070 = \new_[14479]_  ? \new_[15493]_  : \new_[17935]_ ;
  assign n14755 = \new_[14525]_  ? \new_[15493]_  : \new_[18669]_ ;
  assign n14735 = \new_[14480]_  ? \new_[15273]_  : \new_[17950]_ ;
  assign n14075 = \new_[14481]_  ? \new_[15492]_  : \new_[19688]_ ;
  assign n14650 = \new_[14483]_  ? \new_[15486]_  : \new_[18505]_ ;
  assign n14695 = \new_[14484]_  ? \new_[15488]_  : \new_[18348]_ ;
  assign \new_[13490]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0] ;
  assign n14680 = \new_[14485]_  ? \new_[15273]_  : \new_[19606]_ ;
  assign n14605 = \new_[14544]_  ? \new_[15484]_  : \new_[19601]_ ;
  assign n14080 = \new_[14486]_  ? \new_[15592]_  : \new_[19641]_ ;
  assign n14470 = \new_[14488]_  ? \new_[15273]_  : \new_[18599]_ ;
  assign n14085 = \new_[14541]_  ? \new_[15491]_  : \new_[18415]_ ;
  assign n14585 = \new_[14489]_  ? \new_[15488]_  : \new_[19843]_ ;
  assign n14590 = \new_[14490]_  ? \new_[15495]_  : \new_[19098]_ ;
  assign n14495 = \new_[14491]_  ? \new_[15275]_  : \new_[18177]_ ;
  assign n14090 = \new_[14492]_  ? \new_[15488]_  : \new_[19814]_ ;
  assign n14535 = \new_[14493]_  ? \new_[15486]_  : \new_[19105]_ ;
  assign n14505 = \new_[14496]_  ? \new_[15486]_  : \new_[18411]_ ;
  assign n14935 = \new_[14494]_  ? \new_[15488]_  : \new_[18778]_ ;
  assign n14440 = \new_[14498]_  ? \new_[15488]_  : \new_[18634]_ ;
  assign n14455 = \new_[14513]_  ? \new_[15275]_  : \new_[19597]_ ;
  assign n14475 = \new_[14499]_  ? \new_[15488]_  : \new_[17936]_ ;
  assign n14095 = \new_[14500]_  ? \new_[15491]_  : \new_[18334]_ ;
  assign n14450 = \new_[14501]_  ? \new_[15488]_  : \new_[17820]_ ;
  assign n14100 = \new_[14502]_  ? \new_[15485]_  : \new_[19195]_ ;
  assign n13175 = \new_[14503]_  ? \new_[15273]_  : \new_[18232]_ ;
  assign n14105 = \new_[14495]_  ? \new_[15274]_  : \new_[18996]_ ;
  assign n14465 = \new_[14504]_  ? \new_[15592]_  : \new_[17872]_ ;
  assign n13970 = \new_[14505]_  ? \new_[15488]_  : \new_[17829]_ ;
  assign n15115 = \new_[14497]_  ? \new_[15275]_  : \new_[19723]_ ;
  assign n14205 = \new_[14482]_  ? \new_[15488]_  : \new_[19691]_ ;
  assign n14115 = \new_[14452]_  ? \new_[15590]_  : \new_[18309]_ ;
  assign n14110 = \new_[14506]_  ? \new_[15488]_  : \new_[19551]_ ;
  assign n13260 = \new_[14471]_  ? \new_[15488]_  : \new_[19568]_ ;
  assign n13310 = \new_[14465]_  ? \new_[15590]_  : \new_[18575]_ ;
  assign n15240 = \new_[14507]_  ? \new_[15493]_  : \new_[17871]_ ;
  assign n14905 = \new_[14508]_  ? \new_[15486]_  : \new_[19046]_ ;
  assign n14120 = \new_[14457]_  ? \new_[15495]_  : \new_[19240]_ ;
  assign n14560 = \new_[14509]_  ? \new_[15488]_  : \new_[19293]_ ;
  assign n13305 = \new_[14447]_  ? \new_[15485]_  : \new_[18735]_ ;
  assign n13290 = \new_[14510]_  ? \new_[15488]_  : \new_[19049]_ ;
  assign n14125 = \new_[14439]_  ? \new_[15488]_  : \new_[19090]_ ;
  assign n14615 = \new_[14511]_  ? \new_[15488]_  : \new_[17972]_ ;
  assign n15120 = \new_[14431]_  ? \new_[15592]_  : \new_[19003]_ ;
  assign n15155 = \new_[14512]_  ? \new_[15494]_  : \new_[19559]_ ;
  assign n15190 = \new_[14514]_  ? \new_[15275]_  : \new_[19452]_ ;
  assign n14130 = \new_[14515]_  ? \new_[15494]_  : \new_[18894]_ ;
  assign n15205 = \new_[14516]_  ? \new_[15494]_  : \new_[18552]_ ;
  assign n15250 = \new_[14518]_  ? \new_[15488]_  : \new_[19115]_ ;
  assign n15175 = \new_[14487]_  ? \new_[15273]_  : \new_[19528]_ ;
  assign n14510 = \new_[14519]_  ? \new_[15488]_  : \new_[18827]_ ;
  assign n15125 = \new_[14520]_  ? \new_[15488]_  : \new_[17875]_ ;
  assign n14790 = \new_[14466]_  ? \new_[15488]_  : \new_[19237]_ ;
  assign n14845 = \new_[14521]_  ? \new_[15273]_  : \new_[18809]_ ;
  assign n14580 = \new_[14522]_  ? \new_[15488]_  : \new_[19531]_ ;
  assign n14135 = \new_[14435]_  ? \new_[15489]_  : \new_[18980]_ ;
  assign n14960 = \new_[14523]_  ? \new_[15591]_  : \new_[18913]_ ;
  assign n14555 = \new_[14524]_  ? \new_[15592]_  : \new_[18651]_ ;
  assign n14925 = \new_[14477]_  ? \new_[15592]_  : \new_[18498]_ ;
  assign n14870 = \new_[14526]_  ? \new_[15274]_  : \new_[19744]_ ;
  assign n14900 = \new_[14545]_  ? \new_[15485]_  : \new_[18413]_ ;
  assign n14915 = \new_[14528]_  ? \new_[15488]_  : \new_[19039]_ ;
  assign n14145 = \new_[14441]_  ? \new_[15592]_  : \new_[19102]_ ;
  assign n14595 = \new_[14543]_  ? \new_[15492]_  : \new_[18210]_ ;
  assign n14150 = \new_[14529]_  ? \new_[15492]_  : \new_[18430]_ ;
  assign n14810 = \new_[14427]_  ? \new_[15494]_  : \new_[18760]_ ;
  assign n14155 = \new_[14530]_  ? \new_[15592]_  : \new_[19100]_ ;
  assign n14460 = \new_[14537]_  ? \new_[15484]_  : \new_[17979]_ ;
  assign n14820 = \new_[14555]_  ? \new_[15492]_  : \new_[18731]_ ;
  assign n14785 = \new_[14469]_  ? \new_[15273]_  : \new_[19667]_ ;
  assign n14760 = \new_[14552]_  ? \new_[15591]_  : \new_[19740]_ ;
  assign n14655 = \new_[14548]_  ? \new_[15273]_  : \new_[19411]_ ;
  assign n14690 = \new_[14557]_  ? \new_[15274]_  : \new_[19185]_ ;
  assign n14610 = \new_[14554]_  ? \new_[15495]_  : \new_[19445]_ ;
  assign n14685 = \new_[14546]_  ? \new_[15495]_  : \new_[18490]_ ;
  assign n14040 = \new_[14451]_  ? \new_[15492]_  : \new_[19557]_ ;
  assign n14890 = \new_[14517]_  ? \new_[15495]_  : \new_[17865]_ ;
  assign n14065 = \new_[14474]_  ? \new_[15495]_  : \new_[19570]_ ;
  assign n15015 = \new_[14558]_  ? \new_[15273]_  : \new_[18854]_ ;
  assign n14775 = \new_[14549]_  ? \new_[15274]_  : \new_[18833]_ ;
  assign n14175 = \new_[14534]_  ? \new_[15273]_  : \new_[18313]_ ;
  assign n14700 = \new_[14547]_  ? \new_[15591]_  : \new_[18074]_ ;
  assign n14745 = \new_[14550]_  ? \new_[15495]_  : \new_[18393]_ ;
  assign n14600 = \new_[14551]_  ? \new_[15273]_  : \new_[19078]_ ;
  assign n14710 = \new_[14553]_  ? \new_[15485]_  : \new_[19715]_ ;
  assign n14160 = \new_[14556]_  ? \new_[15591]_  : \new_[18193]_ ;
  assign n14850 = \new_[14531]_  ? \new_[15273]_  : \new_[19294]_ ;
  assign \new_[13571]_  = ~\new_[16887]_  | ~\new_[14878]_ ;
  assign \new_[13572]_  = ~\new_[13915]_  & (~\new_[15867]_  | ~\new_[15994]_ );
  assign n15025 = \new_[14753]_  ? \new_[15275]_  : \new_[18709]_ ;
  assign n14185 = \new_[14752]_  ? \new_[15488]_  : \new_[19209]_ ;
  assign n15265 = \new_[14751]_  ? \new_[15275]_  : \new_[18167]_ ;
  assign n14190 = \new_[14754]_  ? \new_[15273]_  : \new_[18803]_ ;
  assign \new_[13577]_  = (~\new_[17036]_  | ~\new_[14560]_ ) & (~\new_[17360]_  | ~\new_[14560]_ );
  assign n14195 = \new_[14814]_  ? \new_[15494]_  : \new_[18806]_ ;
  assign n14200 = \new_[14818]_  ? \new_[15488]_  : \new_[18804]_ ;
  assign n14860 = \new_[14836]_  ? \new_[15488]_  : \new_[18799]_ ;
  assign n14920 = \new_[14832]_  ? \new_[15484]_  : \new_[18802]_ ;
  assign \new_[13582]_  = ~\new_[16639]_  | (~\new_[14749]_  & ~\new_[16998]_ );
  assign \new_[13583]_  = ~\new_[16070]_  | (~\new_[14749]_  & ~\new_[16615]_ );
  assign \new_[13584]_  = ~\new_[13934]_  | (~\new_[10881]_  & ~\new_[16983]_ );
  assign \new_[13585]_  = ~\new_[16500]_  | (~\new_[14749]_  & ~\new_[16881]_ );
  assign \new_[13586]_  = ~\new_[16579]_  | (~\new_[14749]_  & ~\new_[17013]_ );
  assign \new_[13587]_  = ~\new_[16582]_  | (~\new_[14749]_  & ~\new_[16985]_ );
  assign \new_[13588]_  = ~\new_[16587]_  | (~\new_[14749]_  & ~\new_[16888]_ );
  assign \new_[13589]_  = ~\new_[13932]_  | (~\new_[10878]_  & ~\new_[16987]_ );
  assign \new_[13590]_  = ~\new_[16583]_  | (~\new_[14749]_  & ~\new_[16864]_ );
  assign \new_[13591]_  = ~\new_[13933]_  | (~\new_[10886]_  & ~\new_[16977]_ );
  assign \new_[13592]_  = ~\new_[16075]_  | (~\new_[14749]_  & ~\new_[16613]_ );
  assign \new_[13593]_  = ~\new_[16586]_  | (~\new_[14749]_  & ~\new_[16997]_ );
  assign \new_[13594]_  = ~\new_[13935]_  | (~\new_[10938]_  & ~\new_[17103]_ );
  assign \new_[13595]_  = ~\new_[13931]_  | (~\new_[10880]_  & ~\new_[16792]_ );
  assign \new_[13596]_  = ~\new_[16595]_  | (~\new_[14749]_  & ~\new_[16991]_ );
  assign \new_[13597]_  = ~\new_[16740]_  | (~\new_[14749]_  & ~\new_[17067]_ );
  assign \new_[13598]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1] ;
  assign \new_[13599]_  = ~\new_[13819]_  & (~\new_[20298]_  | ~\new_[12418]_ );
  assign \new_[13600]_  = ~n15300 & (~\new_[17460]_  | ~\new_[10375]_ );
  assign \new_[13601]_  = wishbone_slave_unit_pci_initiator_sm_timeout_reg;
  assign n13505 = ~\new_[15875]_  | ~\new_[13822]_ ;
  assign \new_[13603]_  = \new_[14846]_  ? \new_[19906]_  : \new_[5012]_ ;
  assign n14525 = \new_[10393]_  ? \new_[15633]_  : \new_[14844]_ ;
  assign n14515 = \new_[15432]_  ? \new_[14258]_  : \new_[12299]_ ;
  assign \new_[13606]_  = \new_[6319]_  ^ \new_[14849]_ ;
  assign \new_[13607]_  = \wbm_adr_o[30]  ^ \new_[14850]_ ;
  assign \new_[13608]_  = \wbm_adr_o[18]  ? \new_[15502]_  : \new_[14852]_ ;
  assign \new_[13609]_  = \wbm_adr_o[22]  ? \new_[15502]_  : \new_[14853]_ ;
  assign \new_[13610]_  = \new_[13820]_  | \new_[17318]_ ;
  assign \new_[13611]_  = \new_[13820]_  | \new_[16838]_ ;
  assign \new_[13612]_  = \\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0] ;
  assign \new_[13613]_  = ~\new_[14196]_  & (~\new_[5010]_  | ~\new_[19906]_ );
  assign \new_[13614]_  = \wbm_adr_o[25]  ? \new_[15502]_  : \new_[14859]_ ;
  assign \new_[13615]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][39] ;
  assign \new_[13616]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][39] ;
  assign \new_[13617]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][39] ;
  assign \new_[13618]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][39] ;
  assign n13170 = \new_[11961]_  ? \new_[16782]_  : \new_[14540]_ ;
  assign \new_[13620]_  = (~\new_[17158]_  | ~\new_[18953]_ ) & (~\new_[14204]_  | ~\new_[10064]_ );
  assign \new_[13621]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][39] ;
  assign \new_[13622]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][39] ;
  assign \new_[13623]_  = ~\new_[15076]_  | ~\new_[15747]_  | ~\new_[15075]_  | ~\new_[14903]_ ;
  assign \new_[13624]_  = ~\new_[15087]_  | ~\new_[15352]_  | ~\new_[15077]_  | ~\new_[14907]_ ;
  assign \new_[13625]_  = ~\new_[14904]_  | ~\new_[15352]_  | ~\new_[15078]_  | ~\new_[15085]_ ;
  assign \new_[13626]_  = ~\new_[15080]_  | ~\new_[15747]_  | ~\new_[15079]_  | ~\new_[14909]_ ;
  assign \new_[13627]_  = ~\new_[14905]_  | ~\new_[15747]_  | ~\new_[15082]_  | ~\new_[15081]_ ;
  assign \new_[13628]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][39] ;
  assign \new_[13629]_  = ~\new_[13827]_  | ~\new_[16603]_ ;
  assign \new_[13630]_  = ~\new_[13804]_ ;
  assign n13345 = ~\new_[14200]_  | ~\new_[14862]_ ;
  assign n13340 = ~\new_[14187]_  | ~\new_[14862]_ ;
  assign \new_[13633]_  = ~\\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][39] ;
  assign n13335 = ~\new_[13893]_  | (~\new_[14906]_  & ~\new_[17312]_ );
  assign \new_[13635]_  = ~\new_[13807]_ ;
  assign n13355 = ~\new_[14192]_  | (~\new_[14996]_  & ~\wbm_sel_o[0] );
  assign n13360 = ~\new_[14191]_  | (~\new_[14996]_  & ~\wbm_sel_o[1] );
  assign n13350 = ~\new_[14190]_  | (~\new_[14996]_  & ~\wbm_sel_o[2] );
  assign n15105 = ~\new_[14188]_  | (~\new_[14996]_  & ~\wbm_sel_o[3] );
  assign \new_[13640]_  = ~\new_[13938]_  & (~\new_[4970]_  | ~\new_[19906]_ );
  assign n15110 = \new_[12448]_  ? \new_[14221]_  : \new_[15842]_ ;
  assign n13365 = \new_[12011]_  ? \new_[14221]_  : \new_[15832]_ ;
  assign \new_[13643]_  = \new_[19663]_  ? \new_[14221]_  : \new_[15979]_ ;
  assign \new_[13644]_  = ~\new_[15312]_  | ~\new_[15479]_  | ~\new_[19989]_ ;
  assign \new_[13645]_  = ~\new_[15327]_  | ~\new_[20045]_  | ~\new_[15477]_ ;
  assign \new_[13646]_  = ~\new_[15325]_  | ~\new_[15476]_  | ~\new_[14262]_ ;
  assign \new_[13647]_  = ~\new_[15527]_  | ~\new_[15423]_  | ~\new_[14259]_ ;
  assign \new_[13648]_  = ~\new_[19909]_  & ~\new_[13817]_ ;
  assign \new_[13649]_  = ~\new_[15523]_  | ~\new_[15468]_  | ~\new_[20032]_ ;
  assign n13375 = \wbm_adr_o[0]  ? \new_[14219]_  : \new_[12013]_ ;
  assign n15010 = \wbm_adr_o[10]  ? \new_[14219]_  : \new_[12418]_ ;
  assign n13380 = \wbm_adr_o[11]  ? \new_[14219]_  : \new_[12014]_ ;
  assign n13385 = \wbm_adr_o[12]  ? \new_[14219]_  : \new_[12015]_ ;
  assign n15080 = \wbm_adr_o[13]  ? \new_[14219]_  : \new_[12432]_ ;
  assign n15095 = \wbm_adr_o[14]  ? \new_[14219]_  : \new_[12435]_ ;
  assign n13390 = \wbm_adr_o[15]  ? \new_[14218]_  : \new_[12016]_ ;
  assign n15100 = \wbm_adr_o[16]  ? \new_[14219]_  : \new_[12436]_ ;
  assign n15090 = \wbm_adr_o[17]  ? \new_[14219]_  : \new_[12434]_ ;
  assign n15085 = \wbm_adr_o[18]  ? \new_[14218]_  : \new_[12433]_ ;
  assign n13395 = \wbm_adr_o[19]  ? \new_[14218]_  : \new_[12017]_ ;
  assign n15060 = \wbm_adr_o[1]  ? \new_[14219]_  : \new_[12428]_ ;
  assign n13400 = \wbm_adr_o[20]  ? \new_[14996]_  : \new_[12018]_ ;
  assign n15075 = \wbm_adr_o[21]  ? \new_[14219]_  : \new_[12431]_ ;
  assign n13405 = \wbm_adr_o[22]  ? \new_[14219]_  : \new_[12019]_ ;
  assign n15065 = \wbm_adr_o[23]  ? \new_[14996]_  : \new_[12429]_ ;
  assign n15070 = \wbm_adr_o[24]  ? \new_[14218]_  : \new_[12430]_ ;
  assign n15055 = \wbm_adr_o[25]  ? \new_[14218]_  : \new_[12427]_ ;
  assign n15045 = \wbm_adr_o[27]  ? \new_[14219]_  : \new_[12425]_ ;
  assign n13410 = \wbm_adr_o[26]  ? \new_[14219]_  : \new_[12020]_ ;
  assign n13415 = \wbm_adr_o[28]  ? \new_[14219]_  : \new_[12021]_ ;
  assign n15050 = \wbm_adr_o[29]  ? \new_[14219]_  : \new_[12426]_ ;
  assign \new_[13672]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[2] ;
  assign n17395 = \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[0] ;
  assign \new_[13674]_  = \new_[14238]_  & \new_[15747]_ ;
  assign n17165 = \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[2] ;
  assign \new_[13676]_  = ~\new_[14226]_  & ~\new_[15574]_ ;
  assign \new_[13677]_  = ~\new_[14225]_  & ~\new_[15574]_ ;
  assign \new_[13678]_  = pci_target_unit_pci_target_sm_wr_to_fifo_reg;
  assign \new_[13679]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0] ;
  assign \new_[13680]_  = ~\new_[14224]_  & ~\new_[15574]_ ;
  assign \new_[13681]_  = \new_[20044]_  & \new_[16400]_ ;
  assign \new_[13682]_  = ~\new_[14223]_  & ~\new_[15574]_ ;
  assign \new_[13683]_  = ~\new_[14222]_  & ~\new_[15574]_ ;
  assign \new_[13684]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[15] ;
  assign \new_[13685]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[2] ;
  assign \new_[13686]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1] ;
  assign \new_[13687]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[2] ;
  assign \new_[13688]_  = pci_target_unit_del_sync_req_comp_pending_reg;
  assign \new_[13689]_  = wishbone_slave_unit_pci_initiator_sm_transfer_reg;
  assign \new_[13690]_  = (~\new_[14910]_  | ~\new_[20153]_ ) & (~\new_[19555]_  | ~\new_[9903]_ );
  assign n17355 = \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[1] ;
  assign \new_[13692]_  = \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[1] ;
  assign \new_[13693]_  = ~\new_[19920]_  | ~\new_[20143]_ ;
  assign \new_[13694]_  = ~\new_[19920]_  | ~\new_[17383]_ ;
  assign \new_[13695]_  = ~\new_[19920]_  | ~\new_[17080]_ ;
  assign \new_[13696]_  = ~\new_[13818]_ ;
  assign \new_[13697]_  = \new_[10367]_  & \new_[14250]_ ;
  assign \new_[13698]_  = ~\new_[14242]_  | ~\new_[11682]_ ;
  assign \new_[13699]_  = ~\new_[14260]_  | (~\new_[15420]_  & ~\new_[16607]_ );
  assign \new_[13700]_  = ~\new_[14242]_  | ~\new_[11329]_ ;
  assign \new_[13701]_  = ~\new_[14242]_  & ~\new_[20500]_ ;
  assign \new_[13702]_  = ~\new_[15083]_  | ~\new_[15545]_  | ~\new_[15524]_  | ~\new_[16076]_ ;
  assign \new_[13703]_  = ~\new_[15045]_  | ~\new_[15322]_  | ~\new_[14939]_  | ~\new_[16076]_ ;
  assign \new_[13704]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[14] ;
  assign \new_[13705]_  = (~\new_[20212]_  | ~\new_[14933]_ ) & (~\new_[16882]_  | ~\new_[17747]_ );
  assign \new_[13706]_  = ~\new_[14253]_  & (~\new_[20092]_  | ~\new_[12037]_ );
  assign \new_[13707]_  = ~\new_[14254]_  & (~\new_[20092]_  | ~\new_[12309]_ );
  assign n17365 = wishbone_slave_unit_del_sync_comp_rty_exp_reg_reg;
  assign \new_[13709]_  = n16770 ^ \new_[14880]_ ;
  assign \new_[13710]_  = \new_[14221]_  & \new_[17323]_ ;
  assign \new_[13711]_  = ~\new_[15089]_  | ~\new_[14965]_  | ~\new_[14912]_ ;
  assign n15275 = n17055 ? \new_[14932]_  : \new_[17868]_ ;
  assign n15270 = \new_[12548]_  ^ \new_[14932]_ ;
  assign \new_[13714]_  = ~\new_[14293]_  | ~\new_[16672]_ ;
  assign \new_[13715]_  = ~\new_[14290]_  | ~\new_[15814]_ ;
  assign \new_[13716]_  = ~\new_[14890]_ ;
  assign \new_[13717]_  = ~\new_[14229]_  & ~\new_[15564]_ ;
  assign \new_[13718]_  = \new_[19906]_  & \new_[14289]_ ;
  assign \new_[13719]_  = \new_[19884]_  | \new_[17062]_ ;
  assign \new_[13720]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2] ;
  assign \new_[13721]_  = ~\new_[15088]_  | ~\new_[15308]_  | ~\new_[15062]_  | ~\new_[14946]_ ;
  assign \new_[13722]_  = ~\new_[14951]_  & (~\new_[14953]_  | ~\new_[10069]_ );
  assign \new_[13723]_  = ~\new_[14952]_  & (~\new_[14953]_  | ~\new_[10066]_ );
  assign \new_[13724]_  = ~\new_[14947]_  & (~\new_[14953]_  | ~\new_[10068]_ );
  assign \new_[13725]_  = ~\new_[14948]_  & (~\new_[14953]_  | ~\new_[10263]_ );
  assign \new_[13726]_  = ~\new_[14288]_  & (~\new_[16077]_  | ~n17280);
  assign \new_[13727]_  = \wbs_dat_i[6]  ? \new_[14967]_  : \new_[18149]_ ;
  assign \new_[13728]_  = \wbs_dat_i[27]  ? \new_[14967]_  : \new_[18187]_ ;
  assign \new_[13729]_  = \wbs_dat_i[25]  ? \new_[14967]_  : \new_[18389]_ ;
  assign \new_[13730]_  = \wbs_dat_i[2]  ? \new_[14967]_  : \new_[19711]_ ;
  assign \new_[13731]_  = \wbs_dat_i[26]  ? \new_[14967]_  : \new_[18770]_ ;
  assign \new_[13732]_  = \wbs_dat_i[4]  ? \new_[14967]_  : \new_[18897]_ ;
  assign \new_[13733]_  = \wbs_dat_i[24]  ? \new_[14967]_  : \new_[18852]_ ;
  assign \new_[13734]_  = \wbs_dat_i[23]  ? \new_[14967]_  : \new_[19616]_ ;
  assign \new_[13735]_  = \wbs_dat_i[16]  ? \new_[14967]_  : \new_[18574]_ ;
  assign \new_[13736]_  = \wbs_dat_i[12]  ? \new_[14967]_  : \new_[18073]_ ;
  assign \new_[13737]_  = \wbs_dat_i[13]  ? \new_[14967]_  : \new_[18001]_ ;
  assign \new_[13738]_  = \wbs_dat_i[1]  ? \new_[14967]_  : \new_[17887]_ ;
  assign \new_[13739]_  = \wbs_dat_i[21]  ? \new_[14967]_  : \new_[18049]_ ;
  assign \new_[13740]_  = \wbs_dat_i[28]  ? \new_[14967]_  : \new_[18560]_ ;
  assign \new_[13741]_  = \wbs_dat_i[30]  ? \new_[14967]_  : \new_[19674]_ ;
  assign \new_[13742]_  = \wbs_dat_i[31]  ? \new_[14967]_  : \new_[19389]_ ;
  assign \new_[13743]_  = \wbs_dat_i[3]  ? \new_[14967]_  : \new_[19738]_ ;
  assign \new_[13744]_  = \wbs_dat_i[15]  ? \new_[14967]_  : \new_[18176]_ ;
  assign \new_[13745]_  = \wbs_dat_i[5]  ? \new_[14967]_  : \new_[18555]_ ;
  assign \new_[13746]_  = \wbs_dat_i[7]  ? \new_[14967]_  : \new_[19720]_ ;
  assign \new_[13747]_  = \wbs_dat_i[18]  ? \new_[14967]_  : \new_[19501]_ ;
  assign \new_[13748]_  = \wbs_dat_i[11]  ? \new_[14967]_  : \new_[18033]_ ;
  assign \new_[13749]_  = \wbs_dat_i[17]  ? \new_[14967]_  : \new_[19322]_ ;
  assign \new_[13750]_  = \wbs_dat_i[14]  ? \new_[14967]_  : \new_[18586]_ ;
  assign \new_[13751]_  = \wbs_dat_i[0]  ? \new_[14967]_  : \new_[18396]_ ;
  assign \new_[13752]_  = \wbs_dat_i[10]  ? \new_[14967]_  : \new_[18173]_ ;
  assign \new_[13753]_  = \wbs_dat_i[9]  ? \new_[14967]_  : \new_[19835]_ ;
  assign \new_[13754]_  = \wbs_dat_i[19]  ? \new_[14967]_  : \new_[17920]_ ;
  assign \new_[13755]_  = \wbs_dat_i[20]  ? \new_[14967]_  : \new_[19544]_ ;
  assign \new_[13756]_  = \wbs_dat_i[8]  ? \new_[14967]_  : \new_[17822]_ ;
  assign \new_[13757]_  = \wbs_dat_i[22]  ? \new_[14967]_  : \new_[18310]_ ;
  assign \new_[13758]_  = \wbs_dat_i[29]  ? \new_[14967]_  : \new_[19333]_ ;
  assign \new_[13759]_  = ~parity_checker_check_for_serr_on_second_reg;
  assign n15285 = ~\new_[16654]_  | ~\new_[14563]_ ;
  assign \new_[13761]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[1] ;
  assign \new_[13762]_  = ~\new_[14228]_  & ~\new_[20218]_ ;
  assign \new_[13763]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[2] ;
  assign \new_[13764]_  = \new_[14970]_  ? \new_[16795]_  : \new_[18703]_ ;
  assign \new_[13765]_  = \new_[14970]_  ? \new_[16794]_  : \new_[18429]_ ;
  assign \new_[13766]_  = \new_[14970]_  ? \new_[16783]_  : \new_[17856]_ ;
  assign \new_[13767]_  = \new_[14970]_  ? \new_[16803]_  : \new_[18606]_ ;
  assign \new_[13768]_  = ~\new_[14566]_  | (~\new_[11100]_  & ~\new_[16883]_ );
  assign \new_[13769]_  = \new_[19751]_  ? \new_[16984]_  : \new_[14970]_ ;
  assign \new_[13770]_  = ~\new_[14565]_  | (~\new_[11110]_  & ~\new_[16984]_ );
  assign \new_[13771]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2] ;
  assign \new_[13772]_  = \new_[19731]_  ? \new_[16784]_  : \new_[14970]_ ;
  assign \new_[13773]_  = ~\new_[14569]_  | (~\new_[11132]_  & ~\new_[16789]_ );
  assign \new_[13774]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[1] ;
  assign \new_[13775]_  = \new_[17991]_  ? \new_[16883]_  : \new_[14970]_ ;
  assign \new_[13776]_  = \new_[19470]_  ? \new_[16789]_  : \new_[14970]_ ;
  assign \new_[13777]_  = ~\new_[14564]_  | (~\new_[11136]_  & ~\new_[16784]_ );
  assign \new_[13778]_  = ~\new_[14838]_  & ~\new_[16677]_ ;
  assign \new_[13779]_  = \new_[14857]_  & \new_[15994]_ ;
  assign \new_[13780]_  = ~\new_[15994]_  | (~\new_[14901]_  & ~\new_[16992]_ );
  assign \new_[13781]_  = ~\new_[20554]_  | ~\new_[17726]_  | ~\new_[14892]_ ;
  assign \new_[13782]_  = ~\new_[14843]_  & ~\new_[19906]_ ;
  assign \new_[13783]_  = ~\new_[14840]_  & (~\new_[4967]_  | ~\new_[19906]_ );
  assign \new_[13784]_  = \new_[5011]_  ^ \new_[14973]_ ;
  assign \new_[13785]_  = ~\new_[14839]_  & (~\new_[4963]_  | ~\new_[19906]_ );
  assign n15280 = ~\new_[15950]_  | ~\new_[14220]_ ;
  assign \new_[13787]_  = \wbm_adr_o[14]  ? \new_[15502]_  : \new_[14975]_ ;
  assign \new_[13788]_  = ~\new_[14847]_  | (~\new_[15127]_  & ~\new_[6552]_ );
  assign \new_[13789]_  = \new_[4972]_  ^ \new_[14979]_ ;
  assign \new_[13790]_  = \wbm_adr_o[17]  ? \new_[15502]_  : \new_[14982]_ ;
  assign \new_[13791]_  = \new_[14985]_  ? \new_[19906]_  : \new_[5040]_ ;
  assign \new_[13792]_  = \new_[16710]_  ^ \new_[14865]_ ;
  assign \new_[13793]_  = \new_[4175]_  ^ \new_[14865]_ ;
  assign \new_[13794]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[0] ;
  assign \new_[13795]_  = ~\new_[16935]_  | ~\new_[16940]_  | ~\new_[14785]_  | ~\new_[16944]_ ;
  assign \new_[13796]_  = ~\new_[14863]_  & (~\new_[4971]_  | ~\new_[19906]_ );
  assign \new_[13797]_  = \new_[15964]_  ^ \new_[14876]_ ;
  assign \new_[13798]_  = \wbm_adr_o[28]  ? \new_[15502]_  : \new_[14868]_ ;
  assign \new_[13799]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[0] ;
  assign \new_[13800]_  = n16755 ^ \new_[14879]_ ;
  assign \new_[13801]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[12] ;
  assign \new_[13802]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[1] ;
  assign \new_[13803]_  = ~\new_[14231]_  & ~\new_[19906]_ ;
  assign \new_[13804]_  = ~\new_[17264]_  | ~\new_[18502]_  | ~\new_[16098]_  | ~\new_[19882]_ ;
  assign n15290 = \new_[16891]_  | \new_[14204]_ ;
  assign n15295 = ~\new_[14294]_  | (~\new_[15044]_  & ~\new_[20105]_ );
  assign \new_[13807]_  = ~\new_[15438]_  & (~\new_[14936]_  | ~\new_[17113]_ );
  assign \new_[13808]_  = ~\new_[14207]_  & (~\new_[17454]_  | ~\new_[10416]_ );
  assign \new_[13809]_  = \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[3] ;
  assign \new_[13810]_  = i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg;
  assign \new_[13811]_  = ~\new_[14227]_  & ~\new_[15090]_ ;
  assign \new_[13812]_  = \wbm_adr_o[24]  ? \new_[15502]_  : \new_[15006]_ ;
  assign \new_[13813]_  = pci_target_unit_pci_target_if_target_rd_reg;
  assign \new_[13814]_  = ~\new_[20398]_  | ~\new_[19882]_  | ~\new_[11328]_ ;
  assign \new_[13815]_  = \wbm_adr_o[31]  ^ \new_[15020]_ ;
  assign \new_[13816]_  = \wbm_adr_o[19]  ? \new_[15502]_  : \new_[15021]_ ;
  assign \new_[13817]_  = ~\new_[16227]_  & ~\new_[14890]_ ;
  assign \new_[13818]_  = \new_[16224]_  | \new_[14890]_ ;
  assign \new_[13819]_  = ~\new_[15695]_  | ~\new_[15317]_  | ~\new_[15533]_  | ~\new_[15534]_ ;
  assign \new_[13820]_  = ~\new_[16170]_  | ~\new_[16828]_  | ~\new_[20129]_  | ~\new_[20126]_ ;
  assign \new_[13821]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[11] ;
  assign \new_[13822]_  = ~\new_[15351]_  | ~\new_[16572]_  | ~\new_[14931]_  | ~\new_[15618]_ ;
  assign \new_[13823]_  = \new_[16581]_  | \new_[14901]_ ;
  assign n15360 = \new_[14894]_  & \new_[15994]_ ;
  assign n15300 = ~\new_[16839]_  & (~\new_[15853]_  | ~\new_[15030]_ );
  assign \new_[13826]_  = \new_[19589]_  ? \new_[16987]_  : \new_[15130]_ ;
  assign \new_[13827]_  = ~\new_[15434]_  | ~\new_[15853]_  | ~\new_[15030]_ ;
  assign \new_[13828]_  = \new_[18658]_  ? \new_[16983]_  : \new_[15130]_ ;
  assign \new_[13829]_  = \new_[18605]_  ? \new_[16792]_  : \new_[15137]_ ;
  assign \new_[13830]_  = ~\new_[14873]_  & (~\new_[4968]_  | ~\new_[19906]_ );
  assign n15305 = ~\new_[16873]_  | (~\new_[15736]_  & ~\new_[19941]_ );
  assign \new_[13832]_  = ~\new_[20085]_ ;
  assign \new_[13833]_  = ~\new_[14897]_  | (~\new_[16996]_  & ~\new_[15255]_ );
  assign \new_[13834]_  = ~\new_[14899]_  | (~\new_[16485]_  & ~\new_[15255]_ );
  assign \new_[13835]_  = ~\new_[14898]_  | (~\new_[16464]_  & ~\new_[15255]_ );
  assign \new_[13836]_  = ~\new_[14900]_  | (~\new_[15955]_  & ~\new_[15255]_ );
  assign \new_[13837]_  = ~\new_[14896]_  | (~\new_[11691]_  & ~\new_[15255]_ );
  assign \new_[13838]_  = ~\new_[14287]_ ;
  assign \new_[13839]_  = ~\new_[14287]_ ;
  assign \new_[13840]_  = \new_[18211]_  ? \new_[16977]_  : \new_[15148]_ ;
  assign \new_[13841]_  = \new_[15483]_  & \new_[20129]_ ;
  assign \new_[13842]_  = \new_[14938]_  & \new_[15357]_ ;
  assign \new_[13843]_  = ~\new_[15294]_  | ~\new_[15538]_  | ~\new_[15043]_ ;
  assign \new_[13844]_  = ~\new_[15321]_  | ~\new_[15532]_  | ~\new_[15046]_ ;
  assign \new_[13845]_  = ~\new_[14935]_  | ~\new_[20212]_ ;
  assign \new_[13846]_  = ~\new_[15302]_  | ~\new_[15517]_  | ~\new_[15048]_ ;
  assign \new_[13847]_  = ~\new_[15383]_  | ~\new_[15304]_  | ~\new_[15068]_ ;
  assign \new_[13848]_  = ~\new_[16196]_  | ~\new_[16610]_  | ~\new_[15041]_ ;
  assign \new_[13849]_  = ~\new_[15311]_  | ~\new_[15525]_  | ~\new_[15049]_ ;
  assign \new_[13850]_  = \new_[18206]_  ? \new_[16977]_  : \new_[15137]_ ;
  assign \new_[13851]_  = ~\new_[17221]_  | ~\new_[14932]_ ;
  assign \new_[13852]_  = ~\new_[15301]_  | ~\new_[15515]_  | ~\new_[15047]_ ;
  assign \new_[13853]_  = \new_[20052]_  & \new_[15357]_ ;
  assign \new_[13854]_  = ~\new_[14250]_ ;
  assign n15315 = ~\new_[14930]_  | ~\new_[15253]_ ;
  assign n15320 = ~\new_[14928]_  | ~\new_[15253]_ ;
  assign n15310 = ~\new_[14252]_ ;
  assign \new_[13858]_  = ~\new_[16201]_  & (~\new_[15061]_  | ~\new_[5047]_ );
  assign n15355 = ~\new_[14256]_ ;
  assign \new_[13860]_  = ~\new_[15053]_  & (~\new_[15056]_  | ~n17500);
  assign n15345 = ~\new_[14927]_  | (~\new_[16410]_  & ~\new_[15488]_ );
  assign \new_[13862]_  = ~\new_[15054]_  & (~\new_[15056]_  | ~n17350);
  assign \new_[13863]_  = ~\new_[15052]_  & (~\new_[15056]_  | ~n16995);
  assign \new_[13864]_  = ~\new_[15059]_  & (~\new_[15056]_  | ~n17335);
  assign n15395 = \new_[15106]_  ? \new_[15592]_  : \new_[18228]_ ;
  assign n15400 = \new_[15104]_  ? \new_[15485]_  : \new_[19274]_ ;
  assign n15405 = \new_[15108]_  ? \new_[15274]_  : \new_[18725]_ ;
  assign n15380 = \new_[15109]_  ? \new_[15489]_  : \new_[18807]_ ;
  assign \new_[13869]_  = pci_target_unit_pci_target_sm_rd_from_fifo_reg;
  assign \new_[13870]_  = ~\new_[14937]_  & (~\new_[20092]_  | ~\new_[12296]_ );
  assign \new_[13871]_  = \new_[15040]_  ? \new_[16783]_  : \new_[17996]_ ;
  assign \new_[13872]_  = \new_[15040]_  ? \new_[16795]_  : \new_[18279]_ ;
  assign n15325 = ~\new_[14926]_  | (~\new_[13219]_  & ~\new_[15488]_ );
  assign n15350 = ~\new_[14929]_  | (~\new_[17654]_  & ~\new_[15488]_ );
  assign \new_[13875]_  = \new_[15040]_  ? \new_[16803]_  : \new_[18025]_ ;
  assign \new_[13876]_  = \new_[15039]_  ? \new_[16795]_  : \new_[18010]_ ;
  assign \new_[13877]_  = \new_[15039]_  ? \new_[16803]_  : \new_[18028]_ ;
  assign \new_[13878]_  = \new_[15039]_  ? \new_[16794]_  : \new_[19064]_ ;
  assign \new_[13879]_  = \new_[15039]_  ? \new_[16783]_  : \new_[19153]_ ;
  assign \new_[13880]_  = \new_[15040]_  ? \new_[16794]_  : \new_[19805]_ ;
  assign n15385 = \new_[15151]_  ? \new_[15489]_  : \new_[18711]_ ;
  assign n15390 = \new_[15115]_  ? \new_[15590]_  : \new_[18215]_ ;
  assign n15375 = \new_[15117]_  ? \new_[15492]_  : \new_[18188]_ ;
  assign n15370 = \new_[15119]_  ? \new_[15273]_  : \new_[19261]_ ;
  assign \new_[13885]_  = \new_[17818]_  ? \new_[16784]_  : \new_[15039]_ ;
  assign \new_[13886]_  = \new_[19766]_  ? \new_[16784]_  : \new_[15040]_ ;
  assign \new_[13887]_  = \new_[18182]_  ? \new_[16789]_  : \new_[15040]_ ;
  assign \new_[13888]_  = \new_[18243]_  ? \new_[16883]_  : \new_[15040]_ ;
  assign \new_[13889]_  = \new_[18017]_  ? \new_[16984]_  : \new_[15039]_ ;
  assign \new_[13890]_  = \new_[19095]_  ? \new_[16984]_  : \new_[15040]_ ;
  assign \new_[13891]_  = \new_[18016]_  ? \new_[16883]_  : \new_[15039]_ ;
  assign \new_[13892]_  = \new_[19096]_  ? \new_[16789]_  : \new_[15039]_ ;
  assign \new_[13893]_  = ~\new_[10496]_  | ~\new_[17323]_  | ~\new_[14906]_  | ~\new_[19663]_ ;
  assign \new_[13894]_  = ~\new_[14279]_ ;
  assign \new_[13895]_  = ~\new_[14280]_ ;
  assign \new_[13896]_  = ~\new_[14281]_ ;
  assign \new_[13897]_  = ~\new_[14282]_ ;
  assign \new_[13898]_  = ~\new_[14247]_ ;
  assign \new_[13899]_  = ~\new_[14284]_ ;
  assign \new_[13900]_  = ~\new_[14241]_ ;
  assign \new_[13901]_  = ~\new_[14283]_ ;
  assign \new_[13902]_  = ~\new_[15025]_ ;
  assign \new_[13903]_  = ~\new_[15025]_ ;
  assign \new_[13904]_  = ~\new_[14284]_ ;
  assign \new_[13905]_  = ~\new_[14285]_ ;
  assign \new_[13906]_  = ~\new_[15025]_ ;
  assign \new_[13907]_  = ~\new_[14286]_ ;
  assign \new_[13908]_  = ~\new_[14287]_ ;
  assign \new_[13909]_  = ~\new_[14287]_ ;
  assign \new_[13910]_  = ~\new_[14287]_ ;
  assign \new_[13911]_  = ~\new_[14287]_ ;
  assign \new_[13912]_  = ~\new_[14287]_ ;
  assign \new_[13913]_  = ~\new_[14287]_ ;
  assign n15365 = ~\new_[14949]_  & ~\new_[13612]_ ;
  assign \new_[13915]_  = ~\new_[14289]_ ;
  assign n15335 = ~\new_[16874]_  & ~\new_[14949]_ ;
  assign n15330 = ~\new_[16780]_  & (~\new_[15096]_  | ~\new_[18860]_ );
  assign \new_[13918]_  = ~\new_[16370]_  | (~\new_[16795]_  & ~\new_[15330]_ );
  assign \new_[13919]_  = ~\new_[16385]_  | (~\new_[16794]_  & ~\new_[15330]_ );
  assign \new_[13920]_  = \new_[15095]_  ? \new_[16787]_  : \new_[18514]_ ;
  assign \new_[13921]_  = ~\new_[16377]_  | (~\new_[16783]_  & ~\new_[15330]_ );
  assign \new_[13922]_  = \new_[15095]_  ? \new_[16989]_  : \new_[19704]_ ;
  assign \new_[13923]_  = \new_[15095]_  ? \new_[16973]_  : \new_[18908]_ ;
  assign \new_[13924]_  = ~\new_[16378]_  | (~\new_[16803]_  & ~\new_[15330]_ );
  assign \new_[13925]_  = \new_[15095]_  ? \new_[17150]_  : \new_[18021]_ ;
  assign \new_[13926]_  = \new_[19851]_  ? \new_[16983]_  : \new_[15129]_ ;
  assign \new_[13927]_  = \new_[18079]_  ? \new_[16971]_  : \new_[15095]_ ;
  assign \new_[13928]_  = \new_[19054]_  ? \new_[17169]_  : \new_[15095]_ ;
  assign \new_[13929]_  = \new_[19233]_  ? \new_[16910]_  : \new_[15095]_ ;
  assign \new_[13930]_  = \new_[19434]_  ? \new_[16785]_  : \new_[15095]_ ;
  assign \new_[13931]_  = ~\new_[14961]_  | ~\new_[16792]_ ;
  assign \new_[13932]_  = ~\new_[14961]_  | ~\new_[16987]_ ;
  assign \new_[13933]_  = ~\new_[14961]_  | ~\new_[16977]_ ;
  assign \new_[13934]_  = ~\new_[14961]_  | ~\new_[16983]_ ;
  assign \new_[13935]_  = ~\new_[14961]_  | ~\new_[17103]_ ;
  assign \new_[13936]_  = \new_[18424]_  ? \new_[16977]_  : \new_[15134]_ ;
  assign \new_[13937]_  = \new_[15130]_  ? \new_[16998]_  : \new_[19533]_ ;
  assign \new_[13938]_  = ~\new_[14875]_  & ~\new_[19906]_ ;
  assign \new_[13939]_  = \new_[15141]_  ? \new_[16998]_  : \new_[18489]_ ;
  assign \new_[13940]_  = \new_[15130]_  ? \new_[17013]_  : \new_[17845]_ ;
  assign \new_[13941]_  = \new_[15140]_  ? \new_[16998]_  : \new_[19540]_ ;
  assign \new_[13942]_  = \new_[15129]_  ? \new_[16864]_  : \new_[18142]_ ;
  assign \new_[13943]_  = \new_[15145]_  ? \new_[16615]_  : \new_[18397]_ ;
  assign \new_[13944]_  = \new_[15148]_  ? \new_[17013]_  : \new_[19093]_ ;
  assign \new_[13945]_  = \new_[15132]_  ? \new_[16998]_  : \new_[18259]_ ;
  assign \new_[13946]_  = \new_[15130]_  ? \new_[17067]_  : \new_[17883]_ ;
  assign \new_[13947]_  = \new_[15132]_  ? \new_[17067]_  : \new_[19030]_ ;
  assign \new_[13948]_  = \new_[15129]_  ? \new_[17067]_  : \new_[18700]_ ;
  assign \new_[13949]_  = \new_[15143]_  ? \new_[16998]_  : \new_[18266]_ ;
  assign \new_[13950]_  = \new_[15147]_  ? \new_[16998]_  : \new_[19327]_ ;
  assign \new_[13951]_  = \new_[15139]_  ? \new_[16998]_  : \new_[19315]_ ;
  assign \new_[13952]_  = \new_[15145]_  ? \new_[16998]_  : \new_[18320]_ ;
  assign \new_[13953]_  = \new_[15131]_  ? \new_[16998]_  : \new_[18942]_ ;
  assign \new_[13954]_  = \new_[15131]_  ? \new_[17067]_  : \new_[19541]_ ;
  assign \new_[13955]_  = \new_[15137]_  ? \new_[16998]_  : \new_[18361]_ ;
  assign \new_[13956]_  = \new_[15143]_  ? \new_[16615]_  : \new_[18755]_ ;
  assign \new_[13957]_  = \new_[15129]_  ? \new_[16998]_  : \new_[19439]_ ;
  assign \new_[13958]_  = \new_[15147]_  ? \new_[16615]_  : \new_[19348]_ ;
  assign \new_[13959]_  = \new_[15138]_  ? \new_[16615]_  : \new_[19432]_ ;
  assign \new_[13960]_  = \new_[15139]_  ? \new_[16615]_  : \new_[18446]_ ;
  assign \new_[13961]_  = \new_[15148]_  ? \new_[16615]_  : \new_[17906]_ ;
  assign \new_[13962]_  = \new_[15142]_  ? \new_[16998]_  : \new_[19703]_ ;
  assign \new_[13963]_  = \new_[15131]_  ? \new_[16615]_  : \new_[19526]_ ;
  assign \new_[13964]_  = \new_[15134]_  ? \new_[16615]_  : \new_[19133]_ ;
  assign \new_[13965]_  = \new_[15148]_  ? \new_[16998]_  : \new_[19535]_ ;
  assign \new_[13966]_  = \new_[15136]_  ? \new_[16998]_  : \new_[19536]_ ;
  assign \new_[13967]_  = \new_[15131]_  ? \new_[17013]_  : \new_[19485]_ ;
  assign \new_[13968]_  = \new_[15143]_  ? \new_[16991]_  : \new_[19516]_ ;
  assign \new_[13969]_  = \new_[15147]_  ? \new_[16991]_  : \new_[18467]_ ;
  assign \new_[13970]_  = \new_[15139]_  ? \new_[16991]_  : \new_[18470]_ ;
  assign \new_[13971]_  = \new_[15145]_  ? \new_[16991]_  : \new_[19510]_ ;
  assign \new_[13972]_  = \new_[15131]_  ? \new_[16991]_  : \new_[18734]_ ;
  assign \new_[13973]_  = \new_[15132]_  ? \new_[16881]_  : \new_[18525]_ ;
  assign \new_[13974]_  = \new_[15140]_  ? \new_[16881]_  : \new_[18566]_ ;
  assign \new_[13975]_  = \new_[15141]_  ? \new_[16881]_  : \new_[18217]_ ;
  assign \new_[13976]_  = \new_[15147]_  ? \new_[16881]_  : \new_[18882]_ ;
  assign \new_[13977]_  = \new_[15138]_  ? \new_[16881]_  : \new_[18468]_ ;
  assign \new_[13978]_  = \new_[15139]_  ? \new_[16881]_  : \new_[18643]_ ;
  assign \new_[13979]_  = \new_[15136]_  ? \new_[16881]_  : \new_[18865]_ ;
  assign \new_[13980]_  = \new_[15142]_  ? \new_[16881]_  : \new_[18714]_ ;
  assign \new_[13981]_  = \new_[15130]_  ? \new_[16881]_  : \new_[17940]_ ;
  assign \new_[13982]_  = \new_[15134]_  ? \new_[16881]_  : \new_[18591]_ ;
  assign \new_[13983]_  = \new_[15132]_  ? \new_[16997]_  : \new_[19453]_ ;
  assign \new_[13984]_  = \new_[15140]_  ? \new_[16997]_  : \new_[17890]_ ;
  assign \new_[13985]_  = \new_[15143]_  ? \new_[16997]_  : \new_[17827]_ ;
  assign \new_[13986]_  = \new_[15147]_  ? \new_[16997]_  : \new_[19375]_ ;
  assign \new_[13987]_  = \new_[15139]_  ? \new_[16997]_  : \new_[19579]_ ;
  assign \new_[13988]_  = \new_[15145]_  ? \new_[16997]_  : \new_[19729]_ ;
  assign \new_[13989]_  = \new_[15131]_  ? \new_[16997]_  : \new_[17961]_ ;
  assign \new_[13990]_  = \new_[15137]_  ? \new_[16997]_  : \new_[18911]_ ;
  assign \new_[13991]_  = \new_[15143]_  ? \new_[16864]_  : \new_[18125]_ ;
  assign \new_[13992]_  = \new_[15138]_  ? \new_[17067]_  : \new_[18391]_ ;
  assign \new_[13993]_  = \new_[15141]_  ? \new_[17013]_  : \new_[18294]_ ;
  assign \new_[13994]_  = \new_[15138]_  ? \new_[17013]_  : \new_[19084]_ ;
  assign \new_[13995]_  = \new_[15136]_  ? \new_[17013]_  : \new_[18531]_ ;
  assign \new_[13996]_  = \new_[15145]_  ? \new_[17013]_  : \new_[19631]_ ;
  assign \new_[13997]_  = \new_[15142]_  ? \new_[17013]_  : \new_[17846]_ ;
  assign \new_[13998]_  = \new_[15137]_  ? \new_[17013]_  : \new_[19196]_ ;
  assign \new_[13999]_  = \new_[15136]_  ? \new_[16615]_  : \new_[18613]_ ;
  assign \new_[14000]_  = \new_[15129]_  ? \new_[17013]_  : \new_[17837]_ ;
  assign \new_[14001]_  = \new_[15134]_  ? \new_[17013]_  : \new_[18039]_ ;
  assign \new_[14002]_  = \new_[15143]_  ? \new_[16613]_  : \new_[18744]_ ;
  assign \new_[14003]_  = \new_[15147]_  ? \new_[16613]_  : \new_[18937]_ ;
  assign \new_[14004]_  = \new_[15138]_  ? \new_[16613]_  : \new_[18282]_ ;
  assign \new_[14005]_  = \new_[15145]_  ? \new_[16613]_  : \new_[19323]_ ;
  assign \new_[14006]_  = \new_[15131]_  ? \new_[16613]_  : \new_[19473]_ ;
  assign \new_[14007]_  = \new_[15130]_  ? \new_[16613]_  : \new_[19131]_ ;
  assign \new_[14008]_  = \new_[15140]_  ? \new_[16985]_  : \new_[19325]_ ;
  assign \new_[14009]_  = \new_[15143]_  ? \new_[16985]_  : \new_[19862]_ ;
  assign \new_[14010]_  = \new_[15141]_  ? \new_[16985]_  : \new_[17881]_ ;
  assign \new_[14011]_  = \new_[15138]_  ? \new_[16985]_  : \new_[19177]_ ;
  assign \new_[14012]_  = \new_[15136]_  ? \new_[16985]_  : \new_[18045]_ ;
  assign \new_[14013]_  = \new_[15148]_  ? \new_[16985]_  : \new_[19326]_ ;
  assign \new_[14014]_  = \new_[15142]_  ? \new_[16985]_  : \new_[19135]_ ;
  assign \new_[14015]_  = \new_[15131]_  ? \new_[16985]_  : \new_[18050]_ ;
  assign \new_[14016]_  = \new_[15130]_  ? \new_[16985]_  : \new_[19467]_ ;
  assign \new_[14017]_  = \new_[15137]_  ? \new_[16985]_  : \new_[19129]_ ;
  assign \new_[14018]_  = \new_[15129]_  ? \new_[16985]_  : \new_[19702]_ ;
  assign \new_[14019]_  = \new_[15141]_  ? \new_[17067]_  : \new_[19427]_ ;
  assign \new_[14020]_  = \new_[15140]_  ? \new_[16888]_  : \new_[18750]_ ;
  assign \new_[14021]_  = \new_[15141]_  ? \new_[16888]_  : \new_[19213]_ ;
  assign \new_[14022]_  = \new_[15142]_  ? \new_[17067]_  : \new_[19259]_ ;
  assign \new_[14023]_  = \new_[15138]_  ? \new_[16888]_  : \new_[18765]_ ;
  assign \new_[14024]_  = \new_[15136]_  ? \new_[16888]_  : \new_[19599]_ ;
  assign \new_[14025]_  = \new_[15148]_  ? \new_[16888]_  : \new_[18743]_ ;
  assign \new_[14026]_  = \new_[15129]_  ? \new_[16615]_  : \new_[19713]_ ;
  assign \new_[14027]_  = \new_[15142]_  ? \new_[16888]_  : \new_[18817]_ ;
  assign \new_[14028]_  = \new_[15137]_  ? \new_[16888]_  : \new_[19461]_ ;
  assign \new_[14029]_  = \new_[15129]_  ? \new_[16888]_  : \new_[19221]_ ;
  assign \new_[14030]_  = \new_[15134]_  ? \new_[16888]_  : \new_[18319]_ ;
  assign \new_[14031]_  = \new_[15138]_  ? \new_[16864]_  : \new_[18011]_ ;
  assign \new_[14032]_  = \new_[15139]_  ? \new_[16864]_  : \new_[18129]_ ;
  assign \new_[14033]_  = \new_[15145]_  ? \new_[16864]_  : \new_[19588]_ ;
  assign \new_[14034]_  = \new_[15131]_  ? \new_[16864]_  : \new_[18927]_ ;
  assign \new_[14035]_  = \new_[15138]_  ? \new_[16991]_  : \new_[18479]_ ;
  assign \new_[14036]_  = \new_[15139]_  ? \new_[17013]_  : \new_[19488]_ ;
  assign \new_[14037]_  = \new_[15129]_  ? \new_[16991]_  : \new_[19339]_ ;
  assign \new_[14038]_  = \new_[15136]_  ? \new_[17067]_  : \new_[18165]_ ;
  assign \new_[14039]_  = \new_[15147]_  ? \new_[17067]_  : \new_[18141]_ ;
  assign \new_[14040]_  = \new_[15147]_  ? \new_[17013]_  : \new_[18519]_ ;
  assign \new_[14041]_  = \new_[15143]_  ? \new_[17013]_  : \new_[19489]_ ;
  assign \new_[14042]_  = \new_[15140]_  ? \new_[17013]_  : \new_[17965]_ ;
  assign \new_[14043]_  = \new_[15137]_  ? \new_[16864]_  : \new_[18137]_ ;
  assign \new_[14044]_  = \new_[15132]_  ? \new_[16985]_  : \new_[19324]_ ;
  assign \new_[14045]_  = \new_[15137]_  ? \new_[16615]_  : \new_[19522]_ ;
  assign \new_[14046]_  = \new_[15143]_  ? \new_[17067]_  : \new_[19412]_ ;
  assign \new_[14047]_  = \new_[15134]_  ? \new_[16613]_  : \new_[18241]_ ;
  assign \new_[14048]_  = \new_[15132]_  ? \new_[17013]_  : \new_[19695]_ ;
  assign \new_[14049]_  = \new_[15134]_  ? \new_[16997]_  : \new_[17963]_ ;
  assign \new_[14050]_  = \new_[15140]_  ? \new_[16864]_  : \new_[18587]_ ;
  assign \new_[14051]_  = \new_[15129]_  ? \new_[16997]_  : \new_[18872]_ ;
  assign \new_[14052]_  = \new_[15132]_  ? \new_[16864]_  : \new_[18895]_ ;
  assign \new_[14053]_  = \new_[15129]_  ? \new_[16613]_  : \new_[19310]_ ;
  assign \new_[14054]_  = \new_[15130]_  ? \new_[16997]_  : \new_[19666]_ ;
  assign \new_[14055]_  = \new_[15142]_  ? \new_[16997]_  : \new_[17960]_ ;
  assign \new_[14056]_  = \new_[15132]_  ? \new_[16615]_  : \new_[18363]_ ;
  assign \new_[14057]_  = \new_[15148]_  ? \new_[16997]_  : \new_[19637]_ ;
  assign \new_[14058]_  = \new_[15136]_  ? \new_[16997]_  : \new_[19629]_ ;
  assign \new_[14059]_  = \new_[15148]_  ? \new_[16864]_  : \new_[18132]_ ;
  assign \new_[14060]_  = \new_[15140]_  ? \new_[16613]_  : \new_[19480]_ ;
  assign \new_[14061]_  = \new_[15130]_  ? \new_[16888]_  : \new_[18118]_ ;
  assign \new_[14062]_  = \new_[15131]_  ? \new_[16888]_  : \new_[18836]_ ;
  assign \new_[14063]_  = \new_[15138]_  ? \new_[16997]_  : \new_[18336]_ ;
  assign \new_[14064]_  = \new_[15130]_  ? \new_[16864]_  : \new_[19587]_ ;
  assign \new_[14065]_  = \new_[15141]_  ? \new_[16997]_  : \new_[18862]_ ;
  assign \new_[14066]_  = \new_[15145]_  ? \new_[16888]_  : \new_[18740]_ ;
  assign \new_[14067]_  = \new_[15134]_  ? \new_[16985]_  : \new_[18672]_ ;
  assign \new_[14068]_  = \new_[15142]_  ? \new_[16864]_  : \new_[18456]_ ;
  assign \new_[14069]_  = \new_[15136]_  ? \new_[16864]_  : \new_[18130]_ ;
  assign \new_[14070]_  = \new_[15137]_  ? \new_[16613]_  : \new_[19472]_ ;
  assign \new_[14071]_  = \new_[15138]_  ? \new_[16998]_  : \new_[19539]_ ;
  assign \new_[14072]_  = \new_[15141]_  ? \new_[16615]_  : \new_[18679]_ ;
  assign \new_[14073]_  = \new_[15129]_  ? \new_[16881]_  : \new_[19142]_ ;
  assign \new_[14074]_  = \new_[15130]_  ? \new_[16615]_  : \new_[19527]_ ;
  assign \new_[14075]_  = \new_[15142]_  ? \new_[16613]_  : \new_[18304]_ ;
  assign \new_[14076]_  = \new_[15148]_  ? \new_[16613]_  : \new_[17931]_ ;
  assign \new_[14077]_  = \new_[15148]_  ? \new_[16881]_  : \new_[19307]_ ;
  assign \new_[14078]_  = \new_[15137]_  ? \new_[16881]_  : \new_[19500]_ ;
  assign \new_[14079]_  = \new_[15140]_  ? \new_[17067]_  : \new_[18139]_ ;
  assign \new_[14080]_  = \new_[15136]_  ? \new_[16613]_  : \new_[18355]_ ;
  assign \new_[14081]_  = \new_[15131]_  ? \new_[16881]_  : \new_[18780]_ ;
  assign \new_[14082]_  = \new_[15145]_  ? \new_[16985]_  : \new_[18048]_ ;
  assign \new_[14083]_  = \new_[15145]_  ? \new_[16881]_  : \new_[18768]_ ;
  assign \new_[14084]_  = \new_[15147]_  ? \new_[16864]_  : \new_[18128]_ ;
  assign \new_[14085]_  = \new_[15141]_  ? \new_[16864]_  : \new_[17849]_ ;
  assign \new_[14086]_  = \new_[15139]_  ? \new_[16985]_  : \new_[19644]_ ;
  assign \new_[14087]_  = \new_[15134]_  ? \new_[16864]_  : \new_[19423]_ ;
  assign \new_[14088]_  = \new_[15139]_  ? \new_[16613]_  : \new_[17902]_ ;
  assign \new_[14089]_  = \new_[15140]_  ? \new_[16615]_  : \new_[18704]_ ;
  assign \new_[14090]_  = \new_[15134]_  ? \new_[17067]_  : \new_[19287]_ ;
  assign \new_[14091]_  = \new_[15141]_  ? \new_[16991]_  : \new_[19382]_ ;
  assign \new_[14092]_  = \new_[15148]_  ? \new_[17067]_  : \new_[19248]_ ;
  assign \new_[14093]_  = \new_[18576]_  ? \new_[16977]_  : \new_[15136]_ ;
  assign \new_[14094]_  = \new_[15140]_  ? \new_[16991]_  : \new_[18244]_ ;
  assign \new_[14095]_  = \new_[15139]_  ? \new_[16888]_  : \new_[18795]_ ;
  assign \new_[14096]_  = \new_[15139]_  ? \new_[17067]_  : \new_[18221]_ ;
  assign \new_[14097]_  = \new_[15137]_  ? \new_[17067]_  : \new_[19694]_ ;
  assign \new_[14098]_  = \new_[15143]_  ? \new_[16881]_  : \new_[19303]_ ;
  assign \new_[14099]_  = \new_[15148]_  ? \new_[16991]_  : \new_[18478]_ ;
  assign \new_[14100]_  = \new_[15143]_  ? \new_[16888]_  : \new_[18855]_ ;
  assign \new_[14101]_  = \new_[15142]_  ? \new_[16991]_  : \new_[19511]_ ;
  assign \new_[14102]_  = \new_[15137]_  ? \new_[16991]_  : \new_[19155]_ ;
  assign \new_[14103]_  = \new_[15147]_  ? \new_[16985]_  : \new_[18026]_ ;
  assign \new_[14104]_  = \new_[15132]_  ? \new_[16991]_  : \new_[18449]_ ;
  assign \new_[14105]_  = \new_[15130]_  ? \new_[16991]_  : \new_[19507]_ ;
  assign \new_[14106]_  = \new_[15147]_  ? \new_[16888]_  : \new_[19455]_ ;
  assign \new_[14107]_  = \new_[15132]_  ? \new_[16888]_  : \new_[18000]_ ;
  assign \new_[14108]_  = \new_[15134]_  ? \new_[16998]_  : \new_[17898]_ ;
  assign \new_[14109]_  = \new_[15142]_  ? \new_[16615]_  : \new_[19283]_ ;
  assign \new_[14110]_  = \new_[15145]_  ? \new_[17067]_  : \new_[18180]_ ;
  assign \new_[14111]_  = \new_[15141]_  ? \new_[16613]_  : \new_[19478]_ ;
  assign \new_[14112]_  = \new_[15134]_  ? \new_[16991]_  : \new_[19024]_ ;
  assign \new_[14113]_  = \new_[15132]_  ? \new_[16613]_  : \new_[19319]_ ;
  assign \new_[14114]_  = \new_[15136]_  ? \new_[16991]_  : \new_[18473]_ ;
  assign \new_[14115]_  = \new_[18933]_  ? \new_[17103]_  : \new_[15134]_ ;
  assign \new_[14116]_  = \new_[19837]_  ? \new_[16987]_  : \new_[15129]_ ;
  assign \new_[14117]_  = \new_[18196]_  ? \new_[16987]_  : \new_[15138]_ ;
  assign \new_[14118]_  = \new_[19651]_  ? \new_[16983]_  : \new_[15138]_ ;
  assign \new_[14119]_  = \new_[18766]_  ? \new_[16987]_  : \new_[15141]_ ;
  assign \new_[14120]_  = \new_[18097]_  ? \new_[16987]_  : \new_[15143]_ ;
  assign \new_[14121]_  = \new_[18688]_  ? \new_[16987]_  : \new_[15147]_ ;
  assign \new_[14122]_  = \new_[19746]_  ? \new_[16987]_  : \new_[15139]_ ;
  assign \new_[14123]_  = \new_[19868]_  ? \new_[16987]_  : \new_[15145]_ ;
  assign \new_[14124]_  = \new_[19161]_  ? \new_[16987]_  : \new_[15131]_ ;
  assign \new_[14125]_  = \new_[19860]_  ? \new_[16987]_  : \new_[15148]_ ;
  assign \new_[14126]_  = \new_[18208]_  ? \new_[16987]_  : \new_[15137]_ ;
  assign \new_[14127]_  = \new_[18727]_  ? \new_[16792]_  : \new_[15132]_ ;
  assign \new_[14128]_  = \new_[18892]_  ? \new_[16792]_  : \new_[15143]_ ;
  assign \new_[14129]_  = \new_[19468]_  ? \new_[16792]_  : \new_[15147]_ ;
  assign \new_[14130]_  = \new_[19429]_  ? \new_[16792]_  : \new_[15139]_ ;
  assign \new_[14131]_  = \new_[17836]_  ? \new_[16987]_  : \new_[15134]_ ;
  assign \new_[14132]_  = \new_[18991]_  ? \new_[16792]_  : \new_[15145]_ ;
  assign \new_[14133]_  = \new_[19184]_  ? \new_[16792]_  : \new_[15131]_ ;
  assign \new_[14134]_  = \new_[18091]_  ? \new_[16792]_  : \new_[15129]_ ;
  assign \new_[14135]_  = \new_[18829]_  ? \new_[16983]_  : \new_[15141]_ ;
  assign \new_[14136]_  = \new_[19675]_  ? \new_[16983]_  : \new_[15136]_ ;
  assign \new_[14137]_  = \new_[19068]_  ? \new_[16983]_  : \new_[15137]_ ;
  assign \new_[14138]_  = \new_[18426]_  ? \new_[16983]_  : \new_[15134]_ ;
  assign \new_[14139]_  = \new_[19269]_  ? \new_[17103]_  : \new_[15143]_ ;
  assign \new_[14140]_  = \new_[19367]_  ? \new_[17103]_  : \new_[15147]_ ;
  assign \new_[14141]_  = \new_[19072]_  ? \new_[17103]_  : \new_[15139]_ ;
  assign \new_[14142]_  = \new_[19207]_  ? \new_[17103]_  : \new_[15145]_ ;
  assign \new_[14143]_  = \new_[18127]_  ? \new_[17103]_  : \new_[15131]_ ;
  assign \new_[14144]_  = \new_[18813]_  ? \new_[16983]_  : \new_[15132]_ ;
  assign \new_[14145]_  = \new_[18447]_  ? \new_[16792]_  : \new_[15138]_ ;
  assign \new_[14146]_  = \new_[18653]_  ? \new_[16977]_  : \new_[15132]_ ;
  assign \new_[14147]_  = \new_[18683]_  ? \new_[16977]_  : \new_[15141]_ ;
  assign \new_[14148]_  = \new_[18207]_  ? \new_[16977]_  : \new_[15147]_ ;
  assign \new_[14149]_  = \new_[18556]_  ? \new_[16977]_  : \new_[15145]_ ;
  assign \new_[14150]_  = \new_[19698]_  ? \new_[16977]_  : \new_[15142]_ ;
  assign \new_[14151]_  = \new_[18990]_  ? \new_[16977]_  : \new_[15131]_ ;
  assign \new_[14152]_  = \new_[19620]_  ? \new_[16977]_  : \new_[15129]_ ;
  assign \new_[14153]_  = \new_[18154]_  ? \new_[16983]_  : \new_[15140]_ ;
  assign \new_[14154]_  = \new_[19676]_  ? \new_[16983]_  : \new_[15147]_ ;
  assign \new_[14155]_  = \new_[18955]_  ? \new_[16987]_  : \new_[15142]_ ;
  assign \new_[14156]_  = \new_[17885]_  ? \new_[17103]_  : \new_[15140]_ ;
  assign \new_[14157]_  = \new_[19621]_  ? \new_[16792]_  : \new_[15130]_ ;
  assign \new_[14158]_  = \new_[18767]_  ? \new_[17103]_  : \new_[15132]_ ;
  assign \new_[14159]_  = \new_[18535]_  ? \new_[17103]_  : \new_[15129]_ ;
  assign \new_[14160]_  = \new_[19050]_  ? \new_[16977]_  : \new_[15130]_ ;
  assign \new_[14161]_  = \new_[18772]_  ? \new_[16977]_  : \new_[15138]_ ;
  assign \new_[14162]_  = \new_[18919]_  ? \new_[16792]_  : \new_[15142]_ ;
  assign \new_[14163]_  = \new_[18645]_  ? \new_[16977]_  : \new_[15139]_ ;
  assign \new_[14164]_  = \new_[19424]_  ? \new_[16987]_  : \new_[15136]_ ;
  assign \new_[14165]_  = \new_[18015]_  ? \new_[16977]_  : \new_[15143]_ ;
  assign \new_[14166]_  = \new_[18095]_  ? \new_[16977]_  : \new_[15140]_ ;
  assign \new_[14167]_  = \new_[19633]_  ? \new_[16983]_  : \new_[15143]_ ;
  assign \new_[14168]_  = \new_[18850]_  ? \new_[16792]_  : \new_[15141]_ ;
  assign \new_[14169]_  = \new_[18003]_  ? \new_[16983]_  : \new_[15148]_ ;
  assign \new_[14170]_  = \new_[18824]_  ? \new_[16983]_  : \new_[15145]_ ;
  assign \new_[14171]_  = \new_[17809]_  ? \new_[16792]_  : \new_[15134]_ ;
  assign \new_[14172]_  = \new_[19619]_  ? \new_[16983]_  : \new_[15142]_ ;
  assign \new_[14173]_  = \new_[19708]_  ? \new_[16987]_  : \new_[15140]_ ;
  assign \new_[14174]_  = \new_[19836]_  ? \new_[16983]_  : \new_[15139]_ ;
  assign \new_[14175]_  = \new_[18318]_  ? \new_[17103]_  : \new_[15130]_ ;
  assign \new_[14176]_  = \new_[17937]_  ? \new_[16983]_  : \new_[15131]_ ;
  assign \new_[14177]_  = \new_[18333]_  ? \new_[16792]_  : \new_[15148]_ ;
  assign \new_[14178]_  = \new_[19127]_  ? \new_[16987]_  : \new_[15132]_ ;
  assign \new_[14179]_  = \new_[19122]_  ? \new_[17103]_  : \new_[15142]_ ;
  assign \new_[14180]_  = \new_[19778]_  ? \new_[17103]_  : \new_[15148]_ ;
  assign \new_[14181]_  = \new_[19104]_  ? \new_[17103]_  : \new_[15136]_ ;
  assign \new_[14182]_  = \new_[18751]_  ? \new_[17103]_  : \new_[15138]_ ;
  assign \new_[14183]_  = \new_[18374]_  ? \new_[17103]_  : \new_[15137]_ ;
  assign \new_[14184]_  = \new_[19147]_  ? \new_[17103]_  : \new_[15141]_ ;
  assign \new_[14185]_  = \new_[19705]_  ? \new_[16792]_  : \new_[15140]_ ;
  assign \new_[14186]_  = \new_[19574]_  ? \new_[16792]_  : \new_[15136]_ ;
  assign \new_[14187]_  = ~\new_[14996]_  | ~\new_[12006]_ ;
  assign \new_[14188]_  = ~\new_[14996]_  | ~\new_[12437]_ ;
  assign n15340 = ~\new_[16065]_  | (~\new_[16837]_  & ~\new_[16572]_ );
  assign \new_[14190]_  = ~\new_[14996]_  | ~\new_[12008]_ ;
  assign \new_[14191]_  = ~\new_[14996]_  | ~\new_[12010]_ ;
  assign \new_[14192]_  = ~\new_[14996]_  | ~\new_[12009]_ ;
  assign \new_[14193]_  = \new_[6329]_  ^ \new_[15121]_ ;
  assign \new_[14194]_  = \wbm_adr_o[26]  ^ \new_[15133]_ ;
  assign \new_[14195]_  = \new_[18545]_  ^ \new_[15150]_ ;
  assign \new_[14196]_  = ~\new_[14980]_  & ~\new_[19906]_ ;
  assign \new_[14197]_  = ~\new_[14978]_  & (~\new_[5009]_  | ~\new_[19906]_ );
  assign \new_[14198]_  = \wbm_adr_o[29]  ^ \new_[15156]_ ;
  assign \new_[14199]_  = \new_[14987]_  ? \new_[19906]_  : \new_[5038]_ ;
  assign \new_[14200]_  = ~\new_[14996]_  | ~\new_[12007]_ ;
  assign \new_[14201]_  = ~\new_[14889]_  | (~\new_[16166]_  & ~\new_[15255]_ );
  assign \new_[14202]_  = ~\new_[14958]_  & (~\new_[4969]_  | ~\new_[19906]_ );
  assign \new_[14203]_  = ~\new_[14959]_  & (~\new_[4964]_  | ~\new_[19906]_ );
  assign \new_[14204]_  = ~\new_[14996]_  & ~\new_[19175]_ ;
  assign \new_[14205]_  = \wbm_adr_o[16]  ? \new_[15502]_  : \new_[15237]_ ;
  assign pci_inta_oe_o = pci_resets_and_interrupts_inta_en_out_reg;
  assign \new_[14207]_  = ~\new_[15003]_  & ~\new_[17027]_ ;
  assign \new_[14208]_  = \\pci_target_unit_pci_target_if_norm_bc_reg[0] ;
  assign \new_[14209]_  = \\pci_target_unit_pci_target_if_strd_address_reg[3] ;
  assign \new_[14210]_  = \new_[17959]_  ^ \new_[15240]_ ;
  assign \new_[14211]_  = \wbm_adr_o[20]  ? \new_[15502]_  : \new_[15245]_ ;
  assign \new_[14212]_  = \new_[19701]_  ? \new_[16983]_  : \new_[15162]_ ;
  assign \new_[14213]_  = \wbm_adr_o[23]  ? \new_[15502]_  : \new_[15248]_ ;
  assign \new_[14214]_  = \new_[15251]_  ? \new_[19906]_  : \new_[5039]_ ;
  assign \new_[14215]_  = \wbm_adr_o[15]  ? \new_[15502]_  : \new_[15249]_ ;
  assign \new_[14216]_  = \new_[18644]_  ? \new_[16792]_  : \new_[15370]_ ;
  assign \new_[14217]_  = ~\new_[15070]_  | ~\new_[15472]_  | ~\new_[15482]_ ;
  assign \new_[14218]_  = ~\new_[14872]_ ;
  assign \new_[14219]_  = ~\new_[14872]_ ;
  assign \new_[14220]_  = ~\new_[17747]_  | ~\new_[15010]_  | ~\new_[18251]_ ;
  assign \new_[14221]_  = ~\new_[15018]_  | ~\new_[9903]_ ;
  assign \new_[14222]_  = ~\new_[15513]_  | ~\new_[15506]_  | ~\new_[15457]_  | ~\new_[15292]_ ;
  assign \new_[14223]_  = ~\new_[15507]_  | ~\new_[15508]_  | ~\new_[15458]_  | ~\new_[15306]_ ;
  assign \new_[14224]_  = ~\new_[15566]_  | ~\new_[15528]_  | ~\new_[15467]_  | ~\new_[15296]_ ;
  assign \new_[14225]_  = ~\new_[15511]_  | ~\new_[15531]_  | ~\new_[15464]_  | ~\new_[15313]_ ;
  assign \new_[14226]_  = ~\new_[15512]_  | ~\new_[15509]_  | ~\new_[15456]_  | ~\new_[15298]_ ;
  assign \new_[14227]_  = ~\new_[15536]_  | ~\new_[15549]_  | ~\new_[15537]_  | ~\new_[15357]_ ;
  assign \new_[14228]_  = ~\new_[15604]_  & (~\new_[16990]_  | ~\new_[20528]_ );
  assign \new_[14229]_  = ~\new_[20129]_ ;
  assign \new_[14230]_  = \new_[17988]_  ? \new_[16987]_  : \new_[15368]_ ;
  assign \new_[14231]_  = \new_[18791]_  ^ \new_[15241]_ ;
  assign \new_[14232]_  = ~\new_[14998]_  & (~\new_[4965]_  | ~\new_[19906]_ );
  assign \new_[14233]_  = ~\new_[15013]_  | (~\new_[15453]_  & ~\wbm_adr_o[27] );
  assign \new_[14234]_  = \new_[16412]_  ? \new_[15255]_  : \new_[12012]_ ;
  assign \new_[14235]_  = ~\new_[15012]_  & (~\new_[4974]_  | ~\new_[19906]_ );
  assign \new_[14236]_  = ~\new_[15014]_  & (~\new_[4976]_  | ~\new_[19906]_ );
  assign \new_[14237]_  = \new_[19827]_  ? \new_[16977]_  : \new_[15377]_ ;
  assign \new_[14238]_  = ~\new_[15017]_  & (~\new_[20158]_  | ~\new_[17766]_ );
  assign \new_[14239]_  = ~\new_[15011]_  | (~\new_[5008]_  & ~\new_[19906]_ );
  assign n15525 = ~\new_[15008]_  & ~\new_[15836]_ ;
  assign \new_[14241]_  = ~\new_[14881]_ ;
  assign \new_[14242]_  = ~\new_[14888]_ ;
  assign \new_[14243]_  = ~\new_[14888]_ ;
  assign \new_[14244]_  = ~\new_[15261]_  | ~\new_[15074]_ ;
  assign \new_[14245]_  = ~\new_[15573]_  | ~\new_[15459]_  | ~\new_[15282]_ ;
  assign \new_[14246]_  = ~\new_[15269]_  | ~\new_[15071]_ ;
  assign \new_[14247]_  = ~\new_[14919]_ ;
  assign n15470 = \new_[15938]_  & \new_[15033]_ ;
  assign n15480 = \new_[15024]_  & n17365;
  assign \new_[14250]_  = ~\new_[14902]_ ;
  assign n15495 = \new_[16808]_  ? \new_[15488]_  : \new_[13761]_ ;
  assign \new_[14252]_  = ~\new_[15258]_  & (~\new_[15488]_  | ~\new_[13216]_ );
  assign \new_[14253]_  = ~\new_[15034]_  | ~\new_[15687]_ ;
  assign \new_[14254]_  = ~\new_[15036]_  | ~\new_[15691]_ ;
  assign n15485 = \new_[15968]_  ? \new_[15488]_  : \new_[13720]_ ;
  assign \new_[14256]_  = ~\new_[15258]_  & (~\new_[13598]_  | ~\new_[15488]_ );
  assign n15505 = \new_[16137]_  ? \new_[15488]_  : \new_[13771]_ ;
  assign \new_[14258]_  = ~\new_[14888]_ ;
  assign \new_[14259]_  = ~\new_[15032]_  & (~\new_[20450]_  | ~\new_[11682]_ );
  assign \new_[14260]_  = ~\new_[15031]_  & (~\new_[20375]_  | ~\new_[17690]_ );
  assign \new_[14261]_  = \new_[19498]_  ? \new_[15498]_  : \new_[19872]_ ;
  assign \new_[14262]_  = ~\new_[15028]_  & (~\new_[20049]_  | ~\new_[10398]_ );
  assign n15415 = \new_[13216]_  ? \new_[15488]_  : n17395;
  assign n15420 = \new_[13685]_  ? \new_[15488]_  : n17165;
  assign n15520 = n17395 ? \new_[15488]_  : \new_[13799]_ ;
  assign n15410 = n17165 ? \new_[15488]_  : \new_[13672]_ ;
  assign n15440 = \new_[13720]_  ? \new_[15488]_  : \new_[13685]_ ;
  assign n15450 = \new_[13771]_  ? \new_[15488]_  : \new_[13687]_ ;
  assign n15510 = n17355 ? \new_[15488]_  : \new_[13774]_ ;
  assign n15465 = \new_[13437]_  ? \new_[15488]_  : n17355;
  assign n15430 = \wbs_adr_i[0]  ? \new_[15279]_  : \new_[13679]_ ;
  assign n15445 = \wbs_adr_i[1]  ? \new_[15279]_  : \new_[13686]_ ;
  assign n15515 = \wbs_sel_i[0]  ? \new_[15279]_  : \new_[13794]_ ;
  assign n15530 = \wbs_sel_i[1]  ? \new_[15279]_  : \new_[13802]_ ;
  assign n15500 = \wbs_sel_i[2]  ? \new_[15279]_  : \new_[13763]_ ;
  assign n15535 = \wbs_sel_i[3]  ? \new_[15279]_  : \new_[13809]_ ;
  assign n15540 = wbs_we_i ? \new_[15279]_  : \new_[20531]_ ;
  assign \new_[14278]_  = pci_target_unit_wishbone_master_retried_reg;
  assign \new_[14279]_  = ~\new_[14944]_ ;
  assign \new_[14280]_  = ~\new_[14916]_ ;
  assign \new_[14281]_  = ~\new_[14917]_ ;
  assign \new_[14282]_  = ~\new_[14918]_ ;
  assign \new_[14283]_  = ~\new_[14920]_ ;
  assign \new_[14284]_  = ~\new_[13902]_ ;
  assign \new_[14285]_  = ~\new_[14921]_ ;
  assign \new_[14286]_  = ~\new_[14922]_ ;
  assign \new_[14287]_  = ~\new_[14878]_ ;
  assign \new_[14288]_  = ~\new_[15084]_  | ~\new_[15521]_ ;
  assign \new_[14289]_  = \new_[15041]_  | \new_[16782]_ ;
  assign \new_[14290]_  = ~\new_[16665]_  | ~\new_[19360]_  | ~\new_[20081]_  | ~\new_[15355]_ ;
  assign \new_[14291]_  = ~\new_[15098]_  | (~\new_[15572]_  & ~\new_[16678]_ );
  assign \new_[14292]_  = ~n16380 & (~\new_[15331]_  | ~\new_[16577]_ );
  assign \new_[14293]_  = ~\new_[20039]_ ;
  assign \new_[14294]_  = ~\new_[20105]_  | ~\new_[19139]_  | ~\new_[15000]_  | ~\new_[20151]_ ;
  assign \new_[14295]_  = \new_[15203]_  ? \new_[16795]_  : \new_[19730]_ ;
  assign \new_[14296]_  = \new_[15213]_  ? \new_[20485]_  : \new_[19717]_ ;
  assign \new_[14297]_  = \new_[15221]_  ? \new_[16795]_  : \new_[18163]_ ;
  assign \new_[14298]_  = \new_[15211]_  ? \new_[16795]_  : \new_[18283]_ ;
  assign \new_[14299]_  = \new_[15344]_  ? \new_[16795]_  : \new_[18255]_ ;
  assign \new_[14300]_  = \new_[15333]_  ? \new_[16795]_  : \new_[19550]_ ;
  assign \new_[14301]_  = \new_[15206]_  ? \new_[16795]_  : \new_[18433]_ ;
  assign \new_[14302]_  = \new_[15212]_  ? \new_[16783]_  : \new_[18912]_ ;
  assign \new_[14303]_  = \new_[15332]_  ? \new_[16795]_  : \new_[18400]_ ;
  assign \new_[14304]_  = \new_[15345]_  ? \new_[16783]_  : \new_[18497]_ ;
  assign \new_[14305]_  = \new_[15345]_  ? \new_[16795]_  : \new_[18235]_ ;
  assign \new_[14306]_  = \new_[15208]_  ? \new_[16795]_  : \new_[19448]_ ;
  assign \new_[14307]_  = \new_[15211]_  ? \new_[16794]_  : \new_[19134]_ ;
  assign \new_[14308]_  = \new_[15203]_  ? \new_[16794]_  : \new_[18375]_ ;
  assign \new_[14309]_  = \new_[15212]_  ? \new_[16795]_  : \new_[19385]_ ;
  assign \new_[14310]_  = \new_[15342]_  ? \new_[16794]_  : \new_[18237]_ ;
  assign \new_[14311]_  = \new_[15340]_  ? \new_[16795]_  : \new_[19861]_ ;
  assign \new_[14312]_  = \new_[15208]_  ? \new_[16783]_  : \new_[18870]_ ;
  assign \new_[14313]_  = \new_[15219]_  ? \new_[16783]_  : \new_[18493]_ ;
  assign \new_[14314]_  = \new_[15341]_  ? \new_[16794]_  : \new_[18398]_ ;
  assign \new_[14315]_  = \new_[15212]_  ? \new_[16794]_  : \new_[19281]_ ;
  assign \new_[14316]_  = \new_[15340]_  ? \new_[16794]_  : \new_[19359]_ ;
  assign \new_[14317]_  = \new_[15335]_  ? \new_[16795]_  : \new_[18432]_ ;
  assign \new_[14318]_  = \new_[15206]_  ? \new_[16783]_  : \new_[18849]_ ;
  assign \new_[14319]_  = \new_[15336]_  ? \new_[16795]_  : \new_[18461]_ ;
  assign \new_[14320]_  = \new_[15217]_  ? \new_[16783]_  : \new_[19278]_ ;
  assign \new_[14321]_  = \new_[15207]_  ? \new_[16794]_  : \new_[18307]_ ;
  assign \new_[14322]_  = \new_[15344]_  ? \new_[16794]_  : \new_[19618]_ ;
  assign \new_[14323]_  = \new_[15339]_  ? \new_[16794]_  : \new_[19286]_ ;
  assign \new_[14324]_  = \new_[15349]_  ? \new_[16795]_  : \new_[19356]_ ;
  assign \new_[14325]_  = \new_[15214]_  ? \new_[16794]_  : \new_[19290]_ ;
  assign \new_[14326]_  = \new_[15334]_  ? \new_[16795]_  : \new_[19397]_ ;
  assign \new_[14327]_  = \new_[15220]_  ? \new_[16795]_  : \new_[19706]_ ;
  assign \new_[14328]_  = \new_[15343]_  ? \new_[20485]_  : \new_[19280]_ ;
  assign \new_[14329]_  = \new_[15341]_  ? \new_[16795]_  : \new_[19402]_ ;
  assign \new_[14330]_  = \new_[15345]_  ? \new_[16803]_  : \new_[18496]_ ;
  assign \new_[14331]_  = \new_[15215]_  ? \new_[16783]_  : \new_[18984]_ ;
  assign \new_[14332]_  = \new_[15341]_  ? \new_[16783]_  : \new_[18344]_ ;
  assign \new_[14333]_  = \new_[15213]_  ? \new_[16783]_  : \new_[18577]_ ;
  assign \new_[14334]_  = \new_[15207]_  ? \new_[16783]_  : \new_[18706]_ ;
  assign \new_[14335]_  = \new_[15339]_  ? \new_[16795]_  : \new_[18543]_ ;
  assign \new_[14336]_  = \new_[15347]_  ? \new_[16783]_  : \new_[18710]_ ;
  assign \new_[14337]_  = \new_[15217]_  ? \new_[16794]_  : \new_[19298]_ ;
  assign \new_[14338]_  = \new_[15209]_  ? \new_[16783]_  : \new_[19076]_ ;
  assign \new_[14339]_  = \new_[15342]_  ? \new_[16803]_  : \new_[18837]_ ;
  assign \new_[14340]_  = \new_[15217]_  ? \new_[16803]_  : \new_[18784]_ ;
  assign \new_[14341]_  = \new_[15338]_  ? \new_[16794]_  : \new_[19508]_ ;
  assign \new_[14342]_  = \new_[15211]_  ? \new_[16803]_  : \new_[18269]_ ;
  assign \new_[14343]_  = \new_[15348]_  ? \new_[16794]_  : \new_[18761]_ ;
  assign \new_[14344]_  = \new_[15218]_  ? \new_[16794]_  : \new_[18821]_ ;
  assign \new_[14345]_  = \new_[15346]_  ? \new_[16783]_  : \new_[19387]_ ;
  assign \new_[14346]_  = \new_[15342]_  ? \new_[16795]_  : \new_[18626]_ ;
  assign \new_[14347]_  = \new_[15345]_  ? \new_[16794]_  : \new_[19357]_ ;
  assign \new_[14348]_  = \new_[15203]_  ? \new_[16783]_  : \new_[19401]_ ;
  assign \new_[14349]_  = \new_[15338]_  ? \new_[16795]_  : \new_[18477]_ ;
  assign \new_[14350]_  = \new_[15348]_  ? \new_[16783]_  : \new_[19496]_ ;
  assign \new_[14351]_  = \new_[15338]_  ? \new_[16803]_  : \new_[18713]_ ;
  assign \new_[14352]_  = \new_[15212]_  ? \new_[16803]_  : \new_[19301]_ ;
  assign \new_[14353]_  = \new_[15349]_  ? \new_[16803]_  : \new_[18625]_ ;
  assign \new_[14354]_  = \new_[15337]_  ? \new_[16783]_  : \new_[18785]_ ;
  assign \new_[14355]_  = \new_[15214]_  ? \new_[16783]_  : \new_[18572]_ ;
  assign \new_[14356]_  = \new_[15207]_  ? \new_[16795]_  : \new_[18252]_ ;
  assign \new_[14357]_  = \new_[15334]_  ? \new_[16803]_  : \new_[18638]_ ;
  assign \new_[14358]_  = \new_[15203]_  ? \new_[16803]_  : \new_[18702]_ ;
  assign \new_[14359]_  = \new_[15347]_  ? \new_[16803]_  : \new_[18273]_ ;
  assign \new_[14360]_  = \new_[15341]_  ? \new_[16803]_  : \new_[18773]_ ;
  assign \new_[14361]_  = \new_[15346]_  ? \new_[16803]_  : \new_[18623]_ ;
  assign \new_[14362]_  = \new_[15220]_  ? \new_[16803]_  : \new_[18378]_ ;
  assign \new_[14363]_  = \new_[15213]_  ? \new_[16803]_  : \new_[18635]_ ;
  assign \new_[14364]_  = \new_[15217]_  ? \new_[16795]_  : \new_[18466]_ ;
  assign \new_[14365]_  = \new_[15221]_  ? \new_[16803]_  : \new_[18271]_ ;
  assign \new_[14366]_  = \new_[15215]_  ? \new_[16803]_  : \new_[18949]_ ;
  assign \new_[14367]_  = \new_[15333]_  ? \new_[16803]_  : \new_[18032]_ ;
  assign \new_[14368]_  = \new_[15209]_  ? \new_[16803]_  : \new_[18423]_ ;
  assign \new_[14369]_  = \new_[15337]_  ? \new_[16803]_  : \new_[18896]_ ;
  assign \new_[14370]_  = \new_[15218]_  ? \new_[16803]_  : \new_[19379]_ ;
  assign \new_[14371]_  = \new_[15343]_  ? \new_[16803]_  : \new_[18372]_ ;
  assign \new_[14372]_  = \new_[15213]_  ? \new_[16795]_  : \new_[17953]_ ;
  assign \new_[14373]_  = \new_[15340]_  ? \new_[16803]_  : \new_[18745]_ ;
  assign \new_[14374]_  = \new_[15335]_  ? \new_[16783]_  : \new_[18866]_ ;
  assign \new_[14375]_  = \new_[15348]_  ? \new_[16803]_  : \new_[18622]_ ;
  assign \new_[14376]_  = \new_[15218]_  ? \new_[16783]_  : \new_[19734]_ ;
  assign \new_[14377]_  = \new_[15214]_  ? \new_[16795]_  : \new_[18465]_ ;
  assign \new_[14378]_  = \new_[15336]_  ? \new_[16803]_  : \new_[18275]_ ;
  assign \new_[14379]_  = \new_[15340]_  ? \new_[16783]_  : \new_[18800]_ ;
  assign \new_[14380]_  = \new_[15209]_  ? \new_[20485]_  : \new_[19355]_ ;
  assign \new_[14381]_  = \new_[15207]_  ? \new_[16803]_  : \new_[18364]_ ;
  assign \new_[14382]_  = \new_[15339]_  ? \new_[16803]_  : \new_[18699]_ ;
  assign \new_[14383]_  = \new_[15336]_  ? \new_[16783]_  : \new_[18494]_ ;
  assign \new_[14384]_  = \new_[15332]_  ? \new_[16803]_  : \new_[18270]_ ;
  assign \new_[14385]_  = \new_[15215]_  ? \new_[16794]_  : \new_[19299]_ ;
  assign \new_[14386]_  = \new_[15335]_  ? \new_[16803]_  : \new_[18853]_ ;
  assign \new_[14387]_  = \new_[15344]_  ? \new_[16803]_  : \new_[18360]_ ;
  assign \new_[14388]_  = \new_[15219]_  ? \new_[16803]_  : \new_[18612]_ ;
  assign \new_[14389]_  = \new_[15337]_  ? \new_[20485]_  : \new_[18757]_ ;
  assign \new_[14390]_  = \new_[15206]_  ? \new_[16803]_  : \new_[19433]_ ;
  assign \new_[14391]_  = \new_[15214]_  ? \new_[16803]_  : \new_[18652]_ ;
  assign \new_[14392]_  = \new_[15220]_  ? \new_[16794]_  : \new_[19660]_ ;
  assign \new_[14393]_  = \new_[15349]_  ? \new_[16783]_  : \new_[19020]_ ;
  assign \new_[14394]_  = \new_[15220]_  ? \new_[16783]_  : \new_[18155]_ ;
  assign \new_[14395]_  = \new_[15221]_  ? \new_[16783]_  : \new_[18764]_ ;
  assign \new_[14396]_  = \new_[15349]_  ? \new_[20485]_  : \new_[18053]_ ;
  assign \new_[14397]_  = \new_[15347]_  ? \new_[16794]_  : \new_[18376]_ ;
  assign \new_[14398]_  = \new_[15334]_  ? \new_[16794]_  : \new_[19031]_ ;
  assign \new_[14399]_  = \new_[15339]_  ? \new_[16783]_  : \new_[18527]_ ;
  assign \new_[14400]_  = \new_[15333]_  ? \new_[16783]_  : \new_[18485]_ ;
  assign \new_[14401]_  = \new_[15208]_  ? \new_[16803]_  : \new_[18274]_ ;
  assign \new_[14402]_  = \new_[15343]_  ? \new_[16783]_  : \new_[19556]_ ;
  assign \new_[14403]_  = \new_[15346]_  ? \new_[16794]_  : \new_[19005]_ ;
  assign \new_[14404]_  = \new_[15211]_  ? \new_[16783]_  : \new_[17861]_ ;
  assign \new_[14405]_  = \new_[15332]_  ? \new_[16783]_  : \new_[19384]_ ;
  assign \new_[14406]_  = \new_[15342]_  ? \new_[16783]_  : \new_[18974]_ ;
  assign \new_[14407]_  = \new_[15221]_  ? \new_[16794]_  : \new_[18051]_ ;
  assign \new_[14408]_  = \new_[15343]_  ? \new_[16795]_  : \new_[18708]_ ;
  assign \new_[14409]_  = \new_[15333]_  ? \new_[20485]_  : \new_[18660]_ ;
  assign \new_[14410]_  = \new_[15334]_  ? \new_[16783]_  : \new_[18482]_ ;
  assign \new_[14411]_  = \new_[15332]_  ? \new_[16794]_  : \new_[18377]_ ;
  assign \new_[14412]_  = \new_[15215]_  ? \new_[16795]_  : \new_[18464]_ ;
  assign \new_[14413]_  = \new_[15336]_  ? \new_[20485]_  : \new_[19554]_ ;
  assign \new_[14414]_  = \new_[15219]_  ? \new_[16795]_  : \new_[18431]_ ;
  assign \new_[14415]_  = \new_[15337]_  ? \new_[16795]_  : \new_[19605]_ ;
  assign \new_[14416]_  = \new_[15219]_  ? \new_[16794]_  : \new_[19603]_ ;
  assign \new_[14417]_  = \new_[15347]_  ? \new_[16795]_  : \new_[18418]_ ;
  assign \new_[14418]_  = \new_[15208]_  ? \new_[16794]_  : \new_[19081]_ ;
  assign \new_[14419]_  = \new_[15344]_  ? \new_[16783]_  : \new_[18922]_ ;
  assign \new_[14420]_  = \new_[15206]_  ? \new_[20485]_  : \new_[17811]_ ;
  assign \new_[14421]_  = \new_[15209]_  ? \new_[16795]_  : \new_[19377]_ ;
  assign \new_[14422]_  = \new_[15338]_  ? \new_[16783]_  : \new_[18549]_ ;
  assign \new_[14423]_  = \new_[15346]_  ? \new_[16795]_  : \new_[18712]_ ;
  assign \new_[14424]_  = \new_[15218]_  ? \new_[16795]_  : \new_[18452]_ ;
  assign \new_[14425]_  = \new_[15348]_  ? \new_[16795]_  : \new_[18816]_ ;
  assign \new_[14426]_  = \new_[15335]_  ? \new_[16794]_  : \new_[18500]_ ;
  assign \new_[14427]_  = \new_[18760]_  ? \new_[16789]_  : \new_[15348]_ ;
  assign \new_[14428]_  = \new_[17993]_  ? \new_[16784]_  : \new_[15332]_ ;
  assign \new_[14429]_  = \new_[19661]_  ? \new_[16784]_  : \new_[15221]_ ;
  assign \new_[14430]_  = \new_[19622]_  ? \new_[16784]_  : \new_[15203]_ ;
  assign \new_[14431]_  = \new_[19003]_  ? \new_[16883]_  : \new_[15348]_ ;
  assign \new_[14432]_  = \new_[19804]_  ? \new_[16784]_  : \new_[15346]_ ;
  assign \new_[14433]_  = \new_[19244]_  ? \new_[16784]_  : \new_[15347]_ ;
  assign \new_[14434]_  = \new_[18006]_  ? \new_[16784]_  : \new_[15334]_ ;
  assign \new_[14435]_  = \new_[18980]_  ? \new_[16883]_  : \new_[15211]_ ;
  assign \new_[14436]_  = \new_[19736]_  ? \new_[16883]_  : \new_[15212]_ ;
  assign \new_[14437]_  = \new_[19642]_  ? \new_[16784]_  : \new_[15349]_ ;
  assign \new_[14438]_  = \new_[18570]_  ? \new_[16784]_  : \new_[15220]_ ;
  assign \new_[14439]_  = \new_[19090]_  ? \new_[16883]_  : \new_[15336]_ ;
  assign \new_[14440]_  = \new_[18662]_  ? \new_[16784]_  : \new_[15335]_ ;
  assign \new_[14441]_  = \new_[19102]_  ? \new_[16789]_  : \new_[15206]_ ;
  assign \new_[14442]_  = \new_[18819]_  ? \new_[16784]_  : \new_[15206]_ ;
  assign \new_[14443]_  = \new_[18005]_  ? \new_[16784]_  : \new_[15219]_ ;
  assign \new_[14444]_  = \new_[18508]_  ? \new_[16784]_  : \new_[15336]_ ;
  assign \new_[14445]_  = \new_[18524]_  ? \new_[16784]_  : \new_[15348]_ ;
  assign \new_[14446]_  = \new_[18410]_  ? \new_[16784]_  : \new_[15218]_ ;
  assign \new_[14447]_  = \new_[18735]_  ? \new_[16883]_  : \new_[15206]_ ;
  assign \new_[14448]_  = \new_[18233]_  ? \new_[16784]_  : \new_[15209]_ ;
  assign \new_[14449]_  = \new_[17862]_  ? \new_[16784]_  : \new_[15337]_ ;
  assign \new_[14450]_  = \new_[19447]_  ? \new_[16784]_  : \new_[15215]_ ;
  assign \new_[14451]_  = \new_[19557]_  ? \new_[16784]_  : \new_[15338]_ ;
  assign \new_[14452]_  = \new_[18309]_  ? \new_[16883]_  : \new_[15343]_ ;
  assign \new_[14453]_  = \new_[19769]_  ? \new_[16789]_  : \new_[15335]_ ;
  assign \new_[14454]_  = \new_[18387]_  ? \new_[16784]_  : \new_[15214]_ ;
  assign \new_[14455]_  = \new_[18841]_  ? \new_[16784]_  : \new_[15339]_ ;
  assign \new_[14456]_  = \new_[19034]_  ? \new_[16784]_  : \new_[15207]_ ;
  assign \new_[14457]_  = \new_[19240]_  ? \new_[16883]_  : \new_[15335]_ ;
  assign \new_[14458]_  = \new_[19112]_  ? \new_[16784]_  : \new_[15340]_ ;
  assign \new_[14459]_  = \new_[18957]_  ? \new_[16784]_  : \new_[15212]_ ;
  assign \new_[14460]_  = \new_[18278]_  ? \new_[16784]_  : \new_[15341]_ ;
  assign \new_[14461]_  = \new_[18717]_  ? \new_[16784]_  : \new_[15213]_ ;
  assign \new_[14462]_  = \new_[18442]_  ? \new_[16784]_  : \new_[15342]_ ;
  assign \new_[14463]_  = \new_[18610]_  ? \new_[16784]_  : \new_[15211]_ ;
  assign \new_[14464]_  = \new_[18858]_  ? \new_[16784]_  : \new_[15343]_ ;
  assign \new_[14465]_  = \new_[18575]_  ? \new_[16883]_  : \new_[15334]_ ;
  assign \new_[14466]_  = \new_[19237]_  ? \new_[16883]_  : \new_[15339]_ ;
  assign \new_[14467]_  = \new_[19761]_  ? \new_[16984]_  : \new_[15332]_ ;
  assign \new_[14468]_  = \new_[19646]_  ? \new_[16984]_  : \new_[15333]_ ;
  assign \new_[14469]_  = \new_[19667]_  ? \new_[16984]_  : \new_[15221]_ ;
  assign \new_[14470]_  = \new_[18094]_  ? \new_[16984]_  : \new_[15203]_ ;
  assign \new_[14471]_  = \new_[19568]_  ? \new_[16883]_  : \new_[15347]_ ;
  assign \new_[14472]_  = \new_[18104]_  ? \new_[16984]_  : \new_[15346]_ ;
  assign \new_[14473]_  = \new_[19426]_  ? \new_[16984]_  : \new_[15347]_ ;
  assign \new_[14474]_  = \new_[19570]_  ? \new_[16984]_  : \new_[15334]_ ;
  assign \new_[14475]_  = \new_[18592]_  ? \new_[16984]_  : \new_[15349]_ ;
  assign \new_[14476]_  = \new_[19465]_  ? \new_[16984]_  : \new_[15220]_ ;
  assign \new_[14477]_  = \new_[18498]_  ? \new_[16789]_  : \new_[15346]_ ;
  assign \new_[14478]_  = \new_[19492]_  ? \new_[16984]_  : \new_[15335]_ ;
  assign \new_[14479]_  = \new_[17935]_  ? \new_[16984]_  : \new_[15208]_ ;
  assign \new_[14480]_  = \new_[17950]_  ? \new_[16984]_  : \new_[15206]_ ;
  assign \new_[14481]_  = \new_[19688]_  ? \new_[16984]_  : \new_[15219]_ ;
  assign \new_[14482]_  = \new_[19691]_  ? \new_[16883]_  : \new_[15203]_ ;
  assign \new_[14483]_  = \new_[18505]_  ? \new_[16984]_  : \new_[15336]_ ;
  assign \new_[14484]_  = \new_[18348]_  ? \new_[16984]_  : \new_[15345]_ ;
  assign \new_[14485]_  = \new_[19606]_  ? \new_[16984]_  : \new_[15348]_ ;
  assign \new_[14486]_  = \new_[19641]_  ? \new_[16984]_  : \new_[15209]_ ;
  assign \new_[14487]_  = \new_[19528]_  ? \new_[16883]_  : \new_[15217]_ ;
  assign \new_[14488]_  = \new_[18599]_  ? \new_[16984]_  : \new_[15337]_ ;
  assign \new_[14489]_  = \new_[19843]_  ? \new_[16984]_  : \new_[15338]_ ;
  assign \new_[14490]_  = \new_[19098]_  ? \new_[16984]_  : \new_[15217]_ ;
  assign \new_[14491]_  = \new_[18177]_  ? \new_[16984]_  : \new_[15344]_ ;
  assign \new_[14492]_  = \new_[19814]_  ? \new_[16984]_  : \new_[15214]_ ;
  assign \new_[14493]_  = \new_[19105]_  ? \new_[16984]_  : \new_[15339]_ ;
  assign \new_[14494]_  = \new_[18778]_  ? \new_[16789]_  : \new_[15221]_ ;
  assign \new_[14495]_  = \new_[18996]_  ? \new_[16883]_  : \new_[15332]_ ;
  assign \new_[14496]_  = \new_[18411]_  ? \new_[16984]_  : \new_[15207]_ ;
  assign \new_[14497]_  = \new_[19723]_  ? \new_[16883]_  : \new_[15340]_ ;
  assign \new_[14498]_  = \new_[18634]_  ? \new_[16984]_  : \new_[15340]_ ;
  assign \new_[14499]_  = \new_[17936]_  ? \new_[16984]_  : \new_[15341]_ ;
  assign \new_[14500]_  = \new_[18334]_  ? \new_[16984]_  : \new_[15213]_ ;
  assign \new_[14501]_  = \new_[17820]_  ? \new_[16984]_  : \new_[15342]_ ;
  assign \new_[14502]_  = \new_[19195]_  ? \new_[16984]_  : \new_[15211]_ ;
  assign \new_[14503]_  = \new_[18232]_  ? \new_[16984]_  : \new_[15343]_ ;
  assign \new_[14504]_  = \new_[17872]_  ? \new_[16883]_  : \new_[15333]_ ;
  assign \new_[14505]_  = \new_[17829]_  ? \new_[16883]_  : \new_[15221]_ ;
  assign \new_[14506]_  = \new_[19551]_  ? \new_[16883]_  : \new_[15346]_ ;
  assign \new_[14507]_  = \new_[17871]_  ? \new_[16883]_  : \new_[15349]_ ;
  assign \new_[14508]_  = \new_[19046]_  ? \new_[16883]_  : \new_[15220]_ ;
  assign \new_[14509]_  = \new_[19293]_  ? \new_[16883]_  : \new_[15208]_ ;
  assign \new_[14510]_  = \new_[19049]_  ? \new_[16883]_  : \new_[15219]_ ;
  assign \new_[14511]_  = \new_[17972]_  ? \new_[16883]_  : \new_[15345]_ ;
  assign \new_[14512]_  = \new_[19559]_  ? \new_[16883]_  : \new_[15218]_ ;
  assign \new_[14513]_  = \new_[19597]_  ? \new_[16984]_  : \new_[15212]_ ;
  assign \new_[14514]_  = \new_[19452]_  ? \new_[16883]_  : \new_[15209]_ ;
  assign \new_[14515]_  = \new_[18894]_  ? \new_[16883]_  : \new_[15337]_ ;
  assign \new_[14516]_  = \new_[18552]_  ? \new_[16883]_  : \new_[15215]_ ;
  assign \new_[14517]_  = \new_[17865]_  ? \new_[16883]_  : \new_[15342]_ ;
  assign \new_[14518]_  = \new_[19115]_  ? \new_[16883]_  : \new_[15338]_ ;
  assign \new_[14519]_  = \new_[18827]_  ? \new_[16883]_  : \new_[15344]_ ;
  assign \new_[14520]_  = \new_[17875]_  ? \new_[16883]_  : \new_[15214]_ ;
  assign \new_[14521]_  = \new_[18809]_  ? \new_[16883]_  : \new_[15207]_ ;
  assign \new_[14522]_  = \new_[19531]_  ? \new_[16883]_  : \new_[15213]_ ;
  assign \new_[14523]_  = \new_[18913]_  ? \new_[16789]_  : \new_[15332]_ ;
  assign \new_[14524]_  = \new_[18651]_  ? \new_[16789]_  : \new_[15203]_ ;
  assign \new_[14525]_  = \new_[18669]_  ? \new_[16789]_  : \new_[15347]_ ;
  assign \new_[14526]_  = \new_[19744]_  ? \new_[16789]_  : \new_[15334]_ ;
  assign \new_[14527]_  = \new_[19841]_  ? \new_[16789]_  : \new_[15349]_ ;
  assign \new_[14528]_  = \new_[19039]_  ? \new_[16789]_  : \new_[15208]_ ;
  assign \new_[14529]_  = \new_[18430]_  ? \new_[16789]_  : \new_[15345]_ ;
  assign \new_[14530]_  = \new_[19100]_  ? \new_[16789]_  : \new_[15209]_ ;
  assign \new_[14531]_  = \new_[19294]_  ? \new_[16789]_  : \new_[15337]_ ;
  assign \new_[14532]_  = \new_[19060]_  ? \new_[16784]_  : \new_[15344]_ ;
  assign \new_[14533]_  = \new_[19839]_  ? \new_[16784]_  : \new_[15217]_ ;
  assign \new_[14534]_  = \new_[18313]_  ? \new_[16789]_  : \new_[15207]_ ;
  assign \new_[14535]_  = \new_[18647]_  ? \new_[16784]_  : \new_[15345]_ ;
  assign \new_[14536]_  = \new_[19442]_  ? \new_[16784]_  : \new_[15208]_ ;
  assign \new_[14537]_  = \new_[17979]_  ? \new_[16789]_  : \new_[15215]_ ;
  assign \new_[14538]_  = \new_[18172]_  ? \new_[16789]_  : \new_[15219]_ ;
  assign \new_[14539]_  = \new_[18408]_  ? \new_[16789]_  : \new_[15333]_ ;
  assign \new_[14540]_  = ~\new_[14945]_ ;
  assign \new_[14541]_  = \new_[18415]_  ? \new_[16984]_  : \new_[15215]_ ;
  assign \new_[14542]_  = \new_[17954]_  ? \new_[16784]_  : \new_[15333]_ ;
  assign \new_[14543]_  = \new_[18210]_  ? \new_[16789]_  : \new_[15336]_ ;
  assign \new_[14544]_  = \new_[19601]_  ? \new_[16984]_  : \new_[15218]_ ;
  assign \new_[14545]_  = \new_[18413]_  ? \new_[16789]_  : \new_[15220]_ ;
  assign \new_[14546]_  = \new_[18490]_  ? \new_[16789]_  : \new_[15343]_ ;
  assign \new_[14547]_  = \new_[18074]_  ? \new_[16789]_  : \new_[15211]_ ;
  assign \new_[14548]_  = \new_[19411]_  ? \new_[16789]_  : \new_[15341]_ ;
  assign \new_[14549]_  = \new_[18833]_  ? \new_[16789]_  : \new_[15339]_ ;
  assign \new_[14550]_  = \new_[18393]_  ? \new_[16789]_  : \new_[15214]_ ;
  assign \new_[14551]_  = \new_[19078]_  ? \new_[16789]_  : \new_[15212]_ ;
  assign \new_[14552]_  = \new_[19740]_  ? \new_[16789]_  : \new_[15340]_ ;
  assign \new_[14553]_  = \new_[19715]_  ? \new_[16789]_  : \new_[15344]_ ;
  assign \new_[14554]_  = \new_[19445]_  ? \new_[16789]_  : \new_[15342]_ ;
  assign \new_[14555]_  = \new_[18731]_  ? \new_[16789]_  : \new_[15217]_ ;
  assign \new_[14556]_  = \new_[18193]_  ? \new_[16789]_  : \new_[15338]_ ;
  assign \new_[14557]_  = \new_[19185]_  ? \new_[16789]_  : \new_[15213]_ ;
  assign \new_[14558]_  = \new_[18854]_  ? \new_[16883]_  : \new_[15341]_ ;
  assign \new_[14559]_  = \new_[18316]_  ? \new_[16789]_  : \new_[15218]_ ;
  assign \new_[14560]_  = pci_target_unit_wishbone_master_pcir_fifo_wenable_out_reg;
  assign n15460 = ~\new_[15602]_  & ~\new_[15743]_ ;
  assign \new_[14562]_  = ~\new_[15921]_  | ~\new_[15098]_ ;
  assign \new_[14563]_  = ~\new_[14949]_ ;
  assign \new_[14564]_  = ~\new_[16784]_  | ~\new_[15094]_ ;
  assign \new_[14565]_  = ~\new_[16984]_  | ~\new_[15094]_ ;
  assign \new_[14566]_  = ~\new_[16883]_  | ~\new_[15094]_ ;
  assign \new_[14567]_  = \new_[15100]_  | \new_[15934]_ ;
  assign \new_[14568]_  = ~\new_[15100]_  & ~\new_[16122]_ ;
  assign \new_[14569]_  = ~\new_[16789]_  | ~\new_[15094]_ ;
  assign n15455 = \new_[16597]_  & \new_[15096]_ ;
  assign n15490 = ~\new_[14956]_ ;
  assign \new_[14572]_  = \new_[15377]_  ? \new_[16991]_  : \new_[18995]_ ;
  assign \new_[14573]_  = \new_[15372]_  ? \new_[16991]_  : \new_[19503]_ ;
  assign \new_[14574]_  = \new_[15367]_  ? \new_[17067]_  : \new_[18236]_ ;
  assign \new_[14575]_  = \new_[15377]_  ? \new_[16998]_  : \new_[19509]_ ;
  assign \new_[14576]_  = \new_[15369]_  ? \new_[17067]_  : \new_[18226]_ ;
  assign \new_[14577]_  = \new_[15374]_  ? \new_[16998]_  : \new_[18719]_ ;
  assign \new_[14578]_  = \new_[15369]_  ? \new_[17013]_  : \new_[19099]_ ;
  assign \new_[14579]_  = \new_[15368]_  ? \new_[17067]_  : \new_[18864]_ ;
  assign \new_[14580]_  = \new_[15369]_  ? \new_[16615]_  : \new_[18887]_ ;
  assign \new_[14581]_  = \new_[15372]_  ? \new_[17067]_  : \new_[18248]_ ;
  assign \new_[14582]_  = \new_[15365]_  ? \new_[16998]_  : \new_[18276]_ ;
  assign \new_[14583]_  = \new_[15162]_  ? \new_[16998]_  : \new_[18267]_ ;
  assign \new_[14584]_  = \new_[15371]_  ? \new_[16998]_  : \new_[19596]_ ;
  assign \new_[14585]_  = \new_[15370]_  ? \new_[16998]_  : \new_[18291]_ ;
  assign \new_[14586]_  = \new_[15410]_  ? \new_[16998]_  : \new_[19275]_ ;
  assign \new_[14587]_  = \new_[15369]_  ? \new_[16998]_  : \new_[19534]_ ;
  assign \new_[14588]_  = \new_[15367]_  ? \new_[16998]_  : \new_[18330]_ ;
  assign \new_[14589]_  = \new_[15373]_  ? \new_[16998]_  : \new_[18358]_ ;
  assign \new_[14590]_  = \new_[15378]_  ? \new_[16998]_  : \new_[18792]_ ;
  assign \new_[14591]_  = \new_[15366]_  ? \new_[16998]_  : \new_[18716]_ ;
  assign \new_[14592]_  = \new_[15368]_  ? \new_[16998]_  : \new_[18368]_ ;
  assign \new_[14593]_  = \new_[15366]_  ? \new_[17067]_  : \new_[18403]_ ;
  assign \new_[14594]_  = \new_[15374]_  ? \new_[16615]_  : \new_[18369]_ ;
  assign \new_[14595]_  = \new_[15375]_  ? \new_[16615]_  : \new_[19350]_ ;
  assign \new_[14596]_  = \new_[15370]_  ? \new_[17067]_  : \new_[18143]_ ;
  assign \new_[14597]_  = \new_[15372]_  ? \new_[16615]_  : \new_[19523]_ ;
  assign \new_[14598]_  = \new_[15368]_  ? \new_[16615]_  : \new_[17917]_ ;
  assign \new_[14599]_  = \new_[15378]_  ? \new_[17067]_  : \new_[18250]_ ;
  assign \new_[14600]_  = \new_[15376]_  ? \new_[16864]_  : \new_[18012]_ ;
  assign \new_[14601]_  = \new_[15376]_  ? \new_[16998]_  : \new_[18305]_ ;
  assign \new_[14602]_  = \new_[15366]_  ? \new_[16615]_  : \new_[19524]_ ;
  assign \new_[14603]_  = \new_[15375]_  ? \new_[16998]_  : \new_[18327]_ ;
  assign \new_[14604]_  = \new_[15365]_  ? \new_[16991]_  : \new_[19374]_ ;
  assign \new_[14605]_  = \new_[15162]_  ? \new_[16991]_  : \new_[19376]_ ;
  assign \new_[14606]_  = \new_[15371]_  ? \new_[16991]_  : \new_[18463]_ ;
  assign \new_[14607]_  = \new_[15370]_  ? \new_[16991]_  : \new_[19513]_ ;
  assign \new_[14608]_  = \new_[15410]_  ? \new_[16991]_  : \new_[18883]_ ;
  assign \new_[14609]_  = \new_[15373]_  ? \new_[16985]_  : \new_[18059]_ ;
  assign \new_[14610]_  = \new_[15367]_  ? \new_[16991]_  : \new_[18985]_ ;
  assign \new_[14611]_  = \new_[15373]_  ? \new_[16991]_  : \new_[18646]_ ;
  assign \new_[14612]_  = \new_[15378]_  ? \new_[16991]_  : \new_[19340]_ ;
  assign \new_[14613]_  = \new_[15366]_  ? \new_[16991]_  : \new_[18495]_ ;
  assign \new_[14614]_  = pci_target_unit_pci_target_sm_rw_cbe0_reg;
  assign \new_[14615]_  = \new_[15368]_  ? \new_[16991]_  : \new_[18550]_ ;
  assign \new_[14616]_  = \new_[15374]_  ? \new_[16881]_  : \new_[17842]_ ;
  assign \new_[14617]_  = \new_[15377]_  ? \new_[16881]_  : \new_[18281]_ ;
  assign \new_[14618]_  = \new_[15376]_  ? \new_[16881]_  : \new_[17938]_ ;
  assign \new_[14619]_  = \new_[15375]_  ? \new_[16881]_  : \new_[18602]_ ;
  assign \new_[14620]_  = \new_[15369]_  ? \new_[16881]_  : \new_[18812]_ ;
  assign \new_[14621]_  = \new_[15372]_  ? \new_[16881]_  : \new_[18914]_ ;
  assign \new_[14622]_  = \new_[15365]_  ? \new_[16997]_  : \new_[18183]_ ;
  assign \new_[14623]_  = \new_[15162]_  ? \new_[16997]_  : \new_[19499]_ ;
  assign \new_[14624]_  = \new_[15371]_  ? \new_[16997]_  : \new_[18742]_ ;
  assign \new_[14625]_  = \new_[15376]_  ? \new_[16997]_  : \new_[18474]_ ;
  assign \new_[14626]_  = \new_[15369]_  ? \new_[16997]_  : \new_[19654]_ ;
  assign \new_[14627]_  = \new_[15373]_  ? \new_[16997]_  : \new_[19311]_ ;
  assign \new_[14628]_  = \new_[15366]_  ? \new_[16997]_  : \new_[19850]_ ;
  assign \new_[14629]_  = \new_[15368]_  ? \new_[16997]_  : \new_[19848]_ ;
  assign \new_[14630]_  = \new_[15374]_  ? \new_[17013]_  : \new_[19045]_ ;
  assign \new_[14631]_  = \new_[15162]_  ? \new_[17013]_  : \new_[18349]_ ;
  assign \new_[14632]_  = \new_[15377]_  ? \new_[17013]_  : \new_[17966]_ ;
  assign \new_[14633]_  = \new_[15371]_  ? \new_[17013]_  : \new_[18632]_ ;
  assign \new_[14634]_  = \new_[15410]_  ? \new_[17013]_  : \new_[19481]_ ;
  assign \new_[14635]_  = \new_[15376]_  ? \new_[17013]_  : \new_[19314]_ ;
  assign \new_[14636]_  = \new_[15375]_  ? \new_[17013]_  : \new_[17968]_ ;
  assign \new_[14637]_  = \new_[15367]_  ? \new_[17013]_  : \new_[17870]_ ;
  assign \new_[14638]_  = \new_[15373]_  ? \new_[17013]_  : \new_[17974]_ ;
  assign \new_[14639]_  = \new_[15378]_  ? \new_[16615]_  : \new_[19422]_ ;
  assign \new_[14640]_  = \new_[15365]_  ? \new_[16613]_  : \new_[18958]_ ;
  assign \new_[14641]_  = \new_[15374]_  ? \new_[16613]_  : \new_[18659]_ ;
  assign \new_[14642]_  = \new_[15162]_  ? \new_[16613]_  : \new_[19479]_ ;
  assign \new_[14643]_  = \new_[15371]_  ? \new_[16613]_  : \new_[19475]_ ;
  assign \new_[14644]_  = \new_[15370]_  ? \new_[16613]_  : \new_[19476]_ ;
  assign \new_[14645]_  = \new_[15375]_  ? \new_[16613]_  : \new_[17899]_ ;
  assign \new_[14646]_  = \new_[15410]_  ? \new_[16613]_  : \new_[19681]_ ;
  assign \new_[14647]_  = \new_[15369]_  ? \new_[16613]_  : \new_[19474]_ ;
  assign \new_[14648]_  = \new_[15367]_  ? \new_[16613]_  : \new_[19471]_ ;
  assign \new_[14649]_  = \new_[15373]_  ? \new_[16613]_  : \new_[17948]_ ;
  assign \new_[14650]_  = \new_[15378]_  ? \new_[16613]_  : \new_[19491]_ ;
  assign \new_[14651]_  = \new_[15372]_  ? \new_[16613]_  : \new_[19520]_ ;
  assign \new_[14652]_  = \new_[15366]_  ? \new_[16613]_  : \new_[18674]_ ;
  assign \new_[14653]_  = \new_[15368]_  ? \new_[16613]_  : \new_[19469]_ ;
  assign \new_[14654]_  = \new_[15365]_  ? \new_[16985]_  : \new_[18405]_ ;
  assign \new_[14655]_  = \new_[15374]_  ? \new_[16985]_  : \new_[19571]_ ;
  assign \new_[14656]_  = \new_[15377]_  ? \new_[16985]_  : \new_[18229]_ ;
  assign \new_[14657]_  = \new_[15376]_  ? \new_[16985]_  : \new_[19146]_ ;
  assign \new_[14658]_  = \new_[15375]_  ? \new_[16985]_  : \new_[18042]_ ;
  assign \new_[14659]_  = \new_[15378]_  ? \new_[16985]_  : \new_[18280]_ ;
  assign \new_[14660]_  = \new_[15372]_  ? \new_[16985]_  : \new_[18145]_ ;
  assign \new_[14661]_  = \new_[15377]_  ? \new_[17067]_  : \new_[19413]_ ;
  assign \new_[14662]_  = \new_[15374]_  ? \new_[16888]_  : \new_[18859]_ ;
  assign \new_[14663]_  = \new_[15365]_  ? \new_[16881]_  : \new_[19505]_ ;
  assign \new_[14664]_  = \new_[15162]_  ? \new_[16888]_  : \new_[18656]_ ;
  assign \new_[14665]_  = \new_[15377]_  ? \new_[16888]_  : \new_[19464]_ ;
  assign \new_[14666]_  = \new_[15370]_  ? \new_[16888]_  : \new_[18842]_ ;
  assign \new_[14667]_  = \new_[15376]_  ? \new_[16888]_  : \new_[19215]_ ;
  assign \new_[14668]_  = \new_[15375]_  ? \new_[16888]_  : \new_[18698]_ ;
  assign \new_[14669]_  = \new_[15410]_  ? \new_[16888]_  : \new_[19220]_ ;
  assign \new_[14670]_  = \new_[15373]_  ? \new_[16888]_  : \new_[19328]_ ;
  assign \new_[14671]_  = \new_[15372]_  ? \new_[16888]_  : \new_[19329]_ ;
  assign \new_[14672]_  = \new_[15366]_  ? \new_[16888]_  : \new_[19330]_ ;
  assign \new_[14673]_  = \new_[15365]_  ? \new_[16864]_  : \new_[18916]_ ;
  assign \new_[14674]_  = \new_[15162]_  ? \new_[16864]_  : \new_[18008]_ ;
  assign \new_[14675]_  = \new_[15377]_  ? \new_[16864]_  : \new_[18009]_ ;
  assign \new_[14676]_  = \new_[15371]_  ? \new_[16864]_  : \new_[19457]_ ;
  assign \new_[14677]_  = \new_[15370]_  ? \new_[16864]_  : \new_[19456]_ ;
  assign \new_[14678]_  = \new_[15375]_  ? \new_[16864]_  : \new_[18013]_ ;
  assign \new_[14679]_  = \new_[15410]_  ? \new_[16864]_  : \new_[19037]_ ;
  assign \new_[14680]_  = \new_[15369]_  ? \new_[16864]_  : \new_[18131]_ ;
  assign \new_[14681]_  = \new_[15367]_  ? \new_[16864]_  : \new_[18965]_ ;
  assign \new_[14682]_  = \new_[15373]_  ? \new_[16864]_  : \new_[19831]_ ;
  assign \new_[14683]_  = \new_[15378]_  ? \new_[16864]_  : \new_[19228]_ ;
  assign \new_[14684]_  = \new_[15366]_  ? \new_[16864]_  : \new_[19229]_ ;
  assign \new_[14685]_  = \new_[15368]_  ? \new_[16864]_  : \new_[18383]_ ;
  assign \new_[14686]_  = \new_[15366]_  ? \new_[17013]_  : \new_[19483]_ ;
  assign \new_[14687]_  = \new_[15368]_  ? \new_[17013]_  : \new_[19482]_ ;
  assign \new_[14688]_  = \new_[15372]_  ? \new_[17013]_  : \new_[18078]_ ;
  assign \new_[14689]_  = \new_[15371]_  ? \new_[17067]_  : \new_[19415]_ ;
  assign \new_[14690]_  = \new_[15370]_  ? \new_[17013]_  : \new_[17808]_ ;
  assign \new_[14691]_  = \new_[15373]_  ? \new_[16615]_  : \new_[19525]_ ;
  assign \new_[14692]_  = \new_[15367]_  ? \new_[16615]_  : \new_[19515]_ ;
  assign \new_[14693]_  = \new_[15378]_  ? \new_[17013]_  : \new_[17975]_ ;
  assign \new_[14694]_  = \new_[15365]_  ? \new_[17013]_  : \new_[19430]_ ;
  assign \new_[14695]_  = \new_[15372]_  ? \new_[16997]_  : \new_[19004]_ ;
  assign \new_[14696]_  = \new_[15374]_  ? \new_[16864]_  : \new_[19458]_ ;
  assign \new_[14697]_  = \new_[15378]_  ? \new_[16997]_  : \new_[18395]_ ;
  assign \new_[14698]_  = \new_[15376]_  ? \new_[16615]_  : \new_[18650]_ ;
  assign \new_[14699]_  = \new_[15367]_  ? \new_[16997]_  : \new_[18998]_ ;
  assign \new_[14700]_  = \new_[15368]_  ? \new_[16888]_  : \new_[18620]_ ;
  assign \new_[14701]_  = \new_[15378]_  ? \new_[16888]_  : \new_[18558]_ ;
  assign \new_[14702]_  = \new_[15410]_  ? \new_[16997]_  : \new_[19225]_ ;
  assign \new_[14703]_  = \new_[15370]_  ? \new_[16615]_  : \new_[18611]_ ;
  assign \new_[14704]_  = \new_[15375]_  ? \new_[16997]_  : \new_[19437]_ ;
  assign \new_[14705]_  = \new_[15367]_  ? \new_[16888]_  : \new_[18831]_ ;
  assign \new_[14706]_  = \new_[15410]_  ? \new_[16615]_  : \new_[17905]_ ;
  assign \new_[14707]_  = \new_[15370]_  ? \new_[16997]_  : \new_[19871]_ ;
  assign \new_[14708]_  = \new_[15368]_  ? \new_[16985]_  : \new_[18686]_ ;
  assign \new_[14709]_  = \new_[15377]_  ? \new_[16997]_  : \new_[17869]_ ;
  assign \new_[14710]_  = \new_[15366]_  ? \new_[16985]_  : \new_[18109]_ ;
  assign \new_[14711]_  = \new_[15374]_  ? \new_[16997]_  : \new_[19398]_ ;
  assign \new_[14712]_  = \new_[15368]_  ? \new_[16881]_  : \new_[18345]_ ;
  assign \new_[14713]_  = \new_[15377]_  ? \new_[16613]_  : \new_[18782]_ ;
  assign \new_[14714]_  = \new_[15366]_  ? \new_[16881]_  : \new_[18902]_ ;
  assign \new_[14715]_  = \new_[15367]_  ? \new_[16985]_  : \new_[18060]_ ;
  assign \new_[14716]_  = \new_[15378]_  ? \new_[16881]_  : \new_[18593]_ ;
  assign \new_[14717]_  = \new_[15373]_  ? \new_[16881]_  : \new_[17941]_ ;
  assign \new_[14718]_  = \new_[15369]_  ? \new_[16888]_  : \new_[18721]_ ;
  assign \new_[14719]_  = \new_[15367]_  ? \new_[16881]_  : \new_[18793]_ ;
  assign \new_[14720]_  = \new_[15369]_  ? \new_[16985]_  : \new_[18044]_ ;
  assign \new_[14721]_  = \new_[15410]_  ? \new_[16985]_  : \new_[18043]_ ;
  assign \new_[14722]_  = \new_[15370]_  ? \new_[16881]_  : \new_[18880]_ ;
  assign \new_[14723]_  = \new_[15410]_  ? \new_[16881]_  : \new_[19502]_ ;
  assign \new_[14724]_  = \new_[15376]_  ? \new_[16613]_  : \new_[19119]_ ;
  assign \new_[14725]_  = \new_[15372]_  ? \new_[16864]_  : \new_[18138]_ ;
  assign \new_[14726]_  = \new_[15162]_  ? \new_[17067]_  : \new_[19585]_ ;
  assign \new_[14727]_  = \new_[15376]_  ? \new_[17067]_  : \new_[18146]_ ;
  assign \new_[14728]_  = \new_[15370]_  ? \new_[16985]_  : \new_[19170]_ ;
  assign \new_[14729]_  = \new_[15374]_  ? \new_[17067]_  : \new_[17874]_ ;
  assign \new_[14730]_  = \new_[15371]_  ? \new_[16615]_  : \new_[18834]_ ;
  assign \new_[14731]_  = \new_[15365]_  ? \new_[17067]_  : \new_[18136]_ ;
  assign \new_[14732]_  = \new_[15375]_  ? \new_[17067]_  : \new_[19231]_ ;
  assign \new_[14733]_  = \new_[15371]_  ? \new_[16881]_  : \new_[19304]_ ;
  assign \new_[14734]_  = \new_[15410]_  ? \new_[17067]_  : \new_[19234]_ ;
  assign \new_[14735]_  = \new_[15374]_  ? \new_[16991]_  : \new_[19521]_ ;
  assign \new_[14736]_  = \new_[15377]_  ? \new_[16615]_  : \new_[18371]_ ;
  assign \new_[14737]_  = \new_[15369]_  ? \new_[16991]_  : \new_[17932]_ ;
  assign \new_[14738]_  = \new_[15162]_  ? \new_[16615]_  : \new_[18763]_ ;
  assign \new_[14739]_  = \new_[15365]_  ? \new_[16888]_  : \new_[18867]_ ;
  assign \new_[14740]_  = \new_[15376]_  ? \new_[16991]_  : \new_[18546]_ ;
  assign \new_[14741]_  = \new_[15162]_  ? \new_[16881]_  : \new_[19504]_ ;
  assign \new_[14742]_  = \new_[15371]_  ? \new_[16985]_  : \new_[19586]_ ;
  assign \new_[14743]_  = \new_[15375]_  ? \new_[16991]_  : \new_[19295]_ ;
  assign \new_[14744]_  = \new_[15371]_  ? \new_[16888]_  : \new_[18114]_ ;
  assign \new_[14745]_  = \new_[15365]_  ? \new_[16615]_  : \new_[18365]_ ;
  assign \new_[14746]_  = \new_[15162]_  ? \new_[16985]_  : \new_[18209]_ ;
  assign \new_[14747]_  = \new_[15373]_  ? \new_[17067]_  : \new_[18246]_ ;
  assign \new_[14748]_  = \new_[15372]_  ? \new_[16998]_  : \new_[19532]_ ;
  assign \new_[14749]_  = ~\new_[14961]_ ;
  assign \new_[14750]_  = (~\new_[4136]_  | ~\new_[15382]_ ) & (~\new_[20158]_  | ~\new_[17690]_ );
  assign \new_[14751]_  = \new_[15364]_  ? \new_[16795]_  : \new_[18167]_ ;
  assign \new_[14752]_  = \new_[15364]_  ? \new_[16794]_  : \new_[19209]_ ;
  assign \new_[14753]_  = \new_[15364]_  ? \new_[16783]_  : \new_[18709]_ ;
  assign \new_[14754]_  = \new_[15364]_  ? \new_[16803]_  : \new_[18803]_ ;
  assign \new_[14755]_  = \new_[17999]_  ? \new_[16987]_  : \new_[15365]_ ;
  assign \new_[14756]_  = \new_[19451]_  ? \new_[16987]_  : \new_[15162]_ ;
  assign \new_[14757]_  = \new_[19067]_  ? \new_[16987]_  : \new_[15371]_ ;
  assign \new_[14758]_  = \new_[18538]_  ? \new_[16987]_  : \new_[15370]_ ;
  assign \new_[14759]_  = \new_[17859]_  ? \new_[16987]_  : \new_[15410]_ ;
  assign \new_[14760]_  = \new_[18439]_  ? \new_[16987]_  : \new_[15369]_ ;
  assign \new_[14761]_  = \new_[18582]_  ? \new_[16987]_  : \new_[15367]_ ;
  assign \new_[14762]_  = \new_[19813]_  ? \new_[16987]_  : \new_[15373]_ ;
  assign \new_[14763]_  = \new_[18379]_  ? \new_[16987]_  : \new_[15378]_ ;
  assign \new_[14764]_  = \new_[19431]_  ? \new_[16987]_  : \new_[15366]_ ;
  assign \new_[14765]_  = \new_[19130]_  ? \new_[16792]_  : \new_[15365]_ ;
  assign \new_[14766]_  = \new_[17987]_  ? \new_[16792]_  : \new_[15162]_ ;
  assign \new_[14767]_  = \new_[19770]_  ? \new_[16792]_  : \new_[15371]_ ;
  assign \new_[14768]_  = \new_[17847]_  ? \new_[16792]_  : \new_[15410]_ ;
  assign \new_[14769]_  = \new_[19613]_  ? \new_[16792]_  : \new_[15369]_ ;
  assign \new_[14770]_  = \new_[18417]_  ? \new_[16792]_  : \new_[15367]_ ;
  assign \new_[14771]_  = \new_[18648]_  ? \new_[16792]_  : \new_[15373]_ ;
  assign \new_[14772]_  = \new_[19609]_  ? \new_[16792]_  : \new_[15378]_ ;
  assign \new_[14773]_  = \new_[18450]_  ? \new_[16792]_  : \new_[15366]_ ;
  assign \new_[14774]_  = \new_[18068]_  ? \new_[16792]_  : \new_[15368]_ ;
  assign \new_[14775]_  = \new_[18875]_  ? \new_[16983]_  : \new_[15374]_ ;
  assign \new_[14776]_  = \new_[19040]_  ? \new_[16983]_  : \new_[15371]_ ;
  assign \new_[14777]_  = \new_[18564]_  ? \new_[16983]_  : \new_[15370]_ ;
  assign \new_[14778]_  = \new_[17828]_  ? \new_[16983]_  : \new_[15376]_ ;
  assign \new_[14779]_  = \new_[18728]_  ? \new_[16983]_  : \new_[15410]_ ;
  assign \new_[14780]_  = ~\new_[14997]_  & ~\new_[17121]_ ;
  assign \new_[14781]_  = \new_[18690]_  ? \new_[16983]_  : \new_[15367]_ ;
  assign \new_[14782]_  = \new_[17970]_  ? \new_[16983]_  : \new_[15373]_ ;
  assign \new_[14783]_  = \new_[19486]_  ? \new_[16983]_  : \new_[15372]_ ;
  assign \new_[14784]_  = \new_[19239]_  ? \new_[16983]_  : \new_[15366]_ ;
  assign \new_[14785]_  = ~\new_[15001]_  & ~\new_[16950]_ ;
  assign \new_[14786]_  = \new_[18943]_  ? \new_[17103]_  : \new_[15365]_ ;
  assign \new_[14787]_  = \new_[18407]_  ? \new_[17103]_  : \new_[15162]_ ;
  assign \new_[14788]_  = \new_[18801]_  ? \new_[17103]_  : \new_[15371]_ ;
  assign \new_[14789]_  = \new_[19632]_  ? \new_[17103]_  : \new_[15370]_ ;
  assign \new_[14790]_  = \new_[18737]_  ? \new_[17103]_  : \new_[15410]_ ;
  assign \new_[14791]_  = \new_[18486]_  ? \new_[17103]_  : \new_[15369]_ ;
  assign \new_[14792]_  = \new_[18805]_  ? \new_[17103]_  : \new_[15367]_ ;
  assign \new_[14793]_  = \new_[19417]_  ? \new_[16987]_  : \new_[15377]_ ;
  assign \new_[14794]_  = \new_[17907]_  ? \new_[17103]_  : \new_[15373]_ ;
  assign \new_[14795]_  = \new_[18170]_  ? \new_[17103]_  : \new_[15378]_ ;
  assign \new_[14796]_  = \new_[18340]_  ? \new_[17103]_  : \new_[15366]_ ;
  assign \new_[14797]_  = \new_[18746]_  ? \new_[17103]_  : \new_[15368]_ ;
  assign \new_[14798]_  = \new_[19128]_  ? \new_[16983]_  : \new_[15369]_ ;
  assign \new_[14799]_  = \new_[18533]_  ? \new_[16977]_  : \new_[15365]_ ;
  assign \new_[14800]_  = \new_[17995]_  ? \new_[16977]_  : \new_[15162]_ ;
  assign \new_[14801]_  = \new_[19262]_  ? \new_[16977]_  : \new_[15370]_ ;
  assign \new_[14802]_  = \new_[18663]_  ? \new_[16977]_  : \new_[15376]_ ;
  assign \new_[14803]_  = \new_[18797]_  ? \new_[16977]_  : \new_[15410]_ ;
  assign \new_[14804]_  = \new_[19745]_  ? \new_[16977]_  : \new_[15369]_ ;
  assign \new_[14805]_  = \new_[19856]_  ? \new_[16977]_  : \new_[15373]_ ;
  assign \new_[14806]_  = \new_[19565]_  ? \new_[16977]_  : \new_[15378]_ ;
  assign \new_[14807]_  = \new_[18697]_  ? \new_[16977]_  : \new_[15366]_ ;
  assign \new_[14808]_  = \new_[18352]_  ? \new_[16977]_  : \new_[15368]_ ;
  assign \new_[14809]_  = \new_[17857]_  ? \new_[16987]_  : \new_[15375]_ ;
  assign \new_[14810]_  = \new_[19351]_  ? \new_[16983]_  : \new_[15378]_ ;
  assign \new_[14811]_  = \new_[18087]_  ? \new_[16983]_  : \new_[15368]_ ;
  assign \new_[14812]_  = \new_[19847]_  ? \new_[16792]_  : \new_[15375]_ ;
  assign \new_[14813]_  = \new_[19001]_  ? \new_[16792]_  : \new_[15374]_ ;
  assign \new_[14814]_  = \new_[18806]_  ? \new_[16784]_  : \new_[15364]_ ;
  assign \new_[14815]_  = \new_[19866]_  ? \new_[16983]_  : \new_[15365]_ ;
  assign \new_[14816]_  = \new_[19316]_  ? \new_[16977]_  : \new_[15367]_ ;
  assign \new_[14817]_  = \new_[18240]_  ? \new_[16977]_  : \new_[15375]_ ;
  assign \new_[14818]_  = \new_[18804]_  ? \new_[16984]_  : \new_[15364]_ ;
  assign \new_[14819]_  = \new_[18454]_  ? \new_[16792]_  : \new_[15376]_ ;
  assign \new_[14820]_  = \new_[18551]_  ? \new_[16977]_  : \new_[15371]_ ;
  assign \new_[14821]_  = \new_[18830]_  ? \new_[16977]_  : \new_[15374]_ ;
  assign \new_[14822]_  = \new_[17986]_  ? \new_[16987]_  : \new_[15376]_ ;
  assign \new_[14823]_  = \new_[17835]_  ? \new_[16977]_  : \new_[15372]_ ;
  assign \new_[14824]_  = \new_[19628]_  ? \new_[16792]_  : \new_[15372]_ ;
  assign \new_[14825]_  = \new_[18950]_  ? \new_[17103]_  : \new_[15377]_ ;
  assign \new_[14826]_  = \new_[19419]_  ? \new_[16987]_  : \new_[15374]_ ;
  assign \new_[14827]_  = \new_[18420]_  ? \new_[16987]_  : \new_[15372]_ ;
  assign \new_[14828]_  = \new_[18451]_  ? \new_[16983]_  : \new_[15377]_ ;
  assign \new_[14829]_  = \new_[17923]_  ? \new_[16983]_  : \new_[15375]_ ;
  assign \new_[14830]_  = \new_[19786]_  ? \new_[17103]_  : \new_[15374]_ ;
  assign \new_[14831]_  = \new_[19638]_  ? \new_[16792]_  : \new_[15377]_ ;
  assign \new_[14832]_  = \new_[18802]_  ? \new_[16789]_  : \new_[15364]_ ;
  assign \new_[14833]_  = \new_[19548]_  ? \new_[17103]_  : \new_[15375]_ ;
  assign \new_[14834]_  = \new_[19150]_  ? \new_[17103]_  : \new_[15376]_ ;
  assign \new_[14835]_  = \new_[19365]_  ? \new_[17103]_  : \new_[15372]_ ;
  assign \new_[14836]_  = \new_[18799]_  ? \new_[16883]_  : \new_[15364]_ ;
  assign \new_[14837]_  = ~\new_[15746]_  & ~\new_[15382]_ ;
  assign \new_[14838]_  = ~\new_[16829]_  | ~\new_[16837]_  | ~\new_[16801]_  | ~\new_[16638]_ ;
  assign \new_[14839]_  = ~\new_[15116]_  & ~\new_[19906]_ ;
  assign \new_[14840]_  = ~\new_[15112]_  & ~\new_[19906]_ ;
  assign n15425 = ~\new_[15880]_  | ~\new_[15002]_ ;
  assign n15435 = ~\new_[15111]_  & ~\new_[15836]_ ;
  assign \new_[14843]_  = \new_[4896]_  ^ \new_[15379]_ ;
  assign \new_[14844]_  = \new_[15737]_  ? \new_[15255]_  : \new_[12301]_ ;
  assign \new_[14845]_  = \wbm_adr_o[10]  ? \new_[15502]_  : \new_[15381]_ ;
  assign \new_[14846]_  = \new_[5012]_  ^ \new_[15362]_ ;
  assign \new_[14847]_  = ~\new_[15127]_  | ~\new_[6552]_ ;
  assign n15475 = ~\new_[15144]_  & ~\new_[15836]_ ;
  assign \new_[14849]_  = ~\new_[15128]_  & ~\new_[16807]_ ;
  assign \new_[14850]_  = ~\new_[15135]_  & ~\new_[17200]_ ;
  assign \new_[14851]_  = ~\new_[15122]_  | (~\new_[15583]_  & ~\new_[6328]_ );
  assign \new_[14852]_  = ~\new_[15125]_  | (~\new_[15582]_  & ~\wbm_adr_o[18] );
  assign \new_[14853]_  = ~\new_[15126]_  | (~\new_[15584]_  & ~\wbm_adr_o[22] );
  assign \new_[14854]_  = ~\new_[15124]_  & (~\new_[4975]_  | ~\new_[19906]_ );
  assign \new_[14855]_  = \wbm_adr_o[21]  ? \new_[15502]_  : \new_[15408]_ ;
  assign \new_[14856]_  = \wbm_adr_o[13]  ? \new_[15502]_  : \new_[15158]_ ;
  assign \new_[14857]_  = \new_[15810]_  | \new_[16992]_ ;
  assign \new_[14858]_  = ~\new_[15154]_  & (~\new_[4977]_  | ~\new_[19906]_ );
  assign \new_[14859]_  = ~\new_[15152]_  | (~\new_[15414]_  & ~\wbm_adr_o[25] );
  assign \new_[14860]_  = ~\new_[15153]_  & (~\new_[4962]_  | ~\new_[19906]_ );
  assign \new_[14861]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[10] ;
  assign \new_[14862]_  = \new_[14996]_  | \new_[15426]_ ;
  assign \new_[14863]_  = ~\new_[14994]_  & ~\new_[19906]_ ;
  assign \new_[14864]_  = ~\new_[14999]_  & (~\new_[4966]_  | ~\new_[19906]_ );
  assign \new_[14865]_  = \new_[15431]_  ^ \new_[15430]_ ;
  assign \new_[14866]_  = ~\\pci_target_unit_del_sync_be_out_reg[0] ;
  assign \new_[14867]_  = \\input_register_pci_cbe_reg_out_reg[0] ;
  assign \new_[14868]_  = \wbm_adr_o[28]  ^ \new_[15443]_ ;
  assign \new_[14869]_  = \new_[6326]_  ^ \new_[15440]_ ;
  assign \new_[14870]_  = \new_[15593]_  ? \new_[19906]_  : \new_[5044]_ ;
  assign \new_[14871]_  = \wbm_adr_o[12]  ? \new_[15502]_  : \new_[15609]_ ;
  assign \new_[14872]_  = ~\new_[14996]_ ;
  assign \new_[14873]_  = ~\new_[15246]_  & ~\new_[19906]_ ;
  assign \new_[14874]_  = ~\new_[20120]_  | ~\new_[19924]_ ;
  assign \new_[14875]_  = \new_[4970]_  ^ \new_[15466]_ ;
  assign \new_[14876]_  = \new_[16663]_  ^ \new_[15446]_ ;
  assign \new_[14877]_  = ~\new_[15239]_  | (~\new_[15621]_  & ~\new_[6316]_ );
  assign \new_[14878]_  = ~\new_[15025]_ ;
  assign \new_[14879]_  = ~\new_[13684]_  | ~\new_[15353]_  | ~\new_[13704]_ ;
  assign \new_[14880]_  = ~\new_[18100]_  | ~\new_[15288]_  | ~\new_[18595]_ ;
  assign \new_[14881]_  = ~\new_[15025]_ ;
  assign \new_[14882]_  = \new_[15630]_  ? \new_[19906]_  : \new_[5090]_ ;
  assign \new_[14883]_  = \new_[17357]_  ? \new_[19906]_  : \new_[5041]_ ;
  assign \new_[14884]_  = \new_[15956]_  ? \new_[19906]_  : \new_[5042]_ ;
  assign \new_[14885]_  = \wbm_adr_o[8]  ? \new_[15502]_  : \new_[15957]_ ;
  assign \new_[14886]_  = \wbm_adr_o[4]  ? \new_[15502]_  : \new_[16472]_ ;
  assign \new_[14887]_  = \wbm_adr_o[11]  ? \new_[15502]_  : \new_[15629]_ ;
  assign \new_[14888]_  = ~\new_[15259]_  & ~\new_[20151]_ ;
  assign \new_[14889]_  = ~\new_[15255]_  | ~\new_[11622]_ ;
  assign \new_[14890]_  = ~\new_[20119]_ ;
  assign \new_[14891]_  = \new_[15461]_  & \new_[15262]_ ;
  assign \new_[14892]_  = ~\new_[15816]_  & ~\new_[15279]_ ;
  assign \new_[14893]_  = ~\new_[17305]_  | ~\new_[20415]_  | ~\new_[16729]_ ;
  assign \new_[14894]_  = \new_[15254]_  | \new_[13601]_ ;
  assign \new_[14895]_  = ~\new_[15007]_ ;
  assign \new_[14896]_  = ~\new_[11691]_  | ~\new_[15255]_ ;
  assign \new_[14897]_  = ~\new_[15255]_  | ~\new_[11882]_ ;
  assign \new_[14898]_  = ~\new_[15255]_  | ~\new_[11880]_ ;
  assign \new_[14899]_  = ~\new_[15255]_  | ~\new_[11331]_ ;
  assign \new_[14900]_  = ~\new_[15255]_  | ~\new_[11330]_ ;
  assign \new_[14901]_  = ~\new_[15861]_  | ~\new_[16103]_  | ~\new_[17100]_ ;
  assign \new_[14902]_  = ~\new_[15016]_ ;
  assign \new_[14903]_  = ~\new_[15264]_  & (~\new_[12072]_  | ~\new_[19956]_ );
  assign \new_[14904]_  = ~\new_[15266]_  & (~\new_[12074]_  | ~\new_[19956]_ );
  assign \new_[14905]_  = ~\new_[15263]_  & (~\new_[12523]_  | ~\new_[19956]_ );
  assign \new_[14906]_  = ~\new_[15018]_ ;
  assign \new_[14907]_  = ~\new_[15265]_  & (~\new_[12536]_  | ~\new_[19956]_ );
  assign \new_[14908]_  = ~\new_[15995]_  | (~\new_[15503]_  & ~\new_[17180]_ );
  assign \new_[14909]_  = ~\new_[15267]_  & (~\new_[12524]_  | ~\new_[19956]_ );
  assign \new_[14910]_  = \new_[19308]_  ? \new_[19908]_  : \new_[20500]_ ;
  assign \new_[14911]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[8] ;
  assign \new_[14912]_  = ~\new_[15256]_  & (~\new_[20092]_  | ~\new_[12027]_ );
  assign \new_[14913]_  = \wbm_adr_o[3]  ? \new_[15502]_  : \new_[17284]_ ;
  assign \new_[14914]_  = \wbm_adr_o[7]  ? \new_[15502]_  : \new_[15988]_ ;
  assign \new_[14915]_  = \wbm_adr_o[2]  ^ \new_[15502]_ ;
  assign \new_[14916]_  = ~\new_[15025]_ ;
  assign \new_[14917]_  = ~\new_[15025]_ ;
  assign \new_[14918]_  = ~\new_[15025]_ ;
  assign \new_[14919]_  = ~\new_[15025]_ ;
  assign \new_[14920]_  = ~\new_[15025]_ ;
  assign \new_[14921]_  = ~\new_[15025]_ ;
  assign \new_[14922]_  = ~\new_[15025]_ ;
  assign \new_[14923]_  = \new_[15307]_  & \new_[16076]_ ;
  assign \new_[14924]_  = ~\new_[15279]_  | ~\new_[20509]_ ;
  assign \new_[14925]_  = ~\new_[15026]_ ;
  assign \new_[14926]_  = ~\new_[13219]_  | ~\new_[15488]_ ;
  assign \new_[14927]_  = ~\new_[15488]_  | ~\new_[13437]_ ;
  assign \new_[14928]_  = ~\new_[15488]_  | ~\new_[13218]_ ;
  assign \new_[14929]_  = ~\new_[17654]_  | ~\new_[15488]_ ;
  assign \new_[14930]_  = ~\new_[13217]_  | ~\new_[15488]_ ;
  assign \new_[14931]_  = ~\new_[15980]_  & ~\new_[15281]_ ;
  assign \new_[14932]_  = ~\new_[15488]_  & ~\new_[15330]_ ;
  assign \new_[14933]_  = ~\new_[16674]_  & ~\new_[20528]_ ;
  assign \new_[14934]_  = n17010 & \new_[20528]_ ;
  assign \new_[14935]_  = ~\new_[17180]_  & ~\new_[20528]_ ;
  assign \new_[14936]_  = ~\new_[15314]_  & ~\new_[17122]_ ;
  assign \new_[14937]_  = ~\new_[15283]_  | ~\new_[15357]_ ;
  assign \new_[14938]_  = ~\new_[15290]_  & (~\new_[20375]_  | ~\new_[17799]_ );
  assign \new_[14939]_  = ~\new_[15319]_  & (~\new_[20375]_  | ~\new_[17611]_ );
  assign \new_[14940]_  = ~\new_[17583]_  | ~\new_[15994]_  | ~\new_[15561]_ ;
  assign \new_[14941]_  = ~\new_[15278]_  & (~\new_[15749]_  | ~\new_[9988]_ );
  assign \new_[14942]_  = ~\new_[16678]_  | ~\new_[19360]_  | ~\new_[15354]_  | ~\new_[16706]_ ;
  assign \new_[14943]_  = (~\new_[20298]_  | ~\new_[12025]_ ) & (~\new_[9987]_  | ~\new_[15746]_ );
  assign \new_[14944]_  = ~\new_[15025]_ ;
  assign \new_[14945]_  = ~\new_[15226]_  & (~\new_[15607]_  | ~\new_[19139]_ );
  assign \new_[14946]_  = \new_[15360]_  | \new_[15942]_ ;
  assign \new_[14947]_  = ~\new_[15359]_  & ~\new_[15902]_ ;
  assign \new_[14948]_  = ~\new_[15359]_  & ~\new_[15898]_ ;
  assign \new_[14949]_  = ~\new_[16620]_  | ~\new_[15572]_  | ~\new_[20081]_ ;
  assign \new_[14950]_  = ~\new_[15572]_  & ~\new_[16706]_ ;
  assign \new_[14951]_  = ~\new_[15359]_  & ~\new_[15905]_ ;
  assign \new_[14952]_  = ~\new_[15359]_  & ~\new_[15900]_ ;
  assign \new_[14953]_  = \new_[15359]_  | \new_[17258]_ ;
  assign n15545 = ~\new_[18082]_  & (~\new_[15576]_  | ~n16775);
  assign \new_[14955]_  = \new_[15205]_  & \new_[15354]_ ;
  assign \new_[14956]_  = ~\new_[17476]_  | ~\new_[15356]_  | ~\new_[17318]_ ;
  assign \new_[14957]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[13] ;
  assign \new_[14958]_  = ~\new_[15234]_  & ~\new_[19906]_ ;
  assign \new_[14959]_  = ~\new_[15235]_  & ~\new_[19906]_ ;
  assign \new_[14960]_  = (~\new_[20092]_  | ~\new_[12405]_ ) & (~\new_[15569]_  | ~\new_[9992]_ );
  assign \new_[14961]_  = \new_[15384]_  | \new_[17310]_ ;
  assign \new_[14962]_  = (~\new_[15749]_  | ~\new_[9996]_ ) & (~\new_[15569]_  | ~\new_[9986]_ );
  assign \new_[14963]_  = (~\new_[10069]_  | ~\new_[15746]_ ) & (~\new_[16077]_  | ~n17350);
  assign \new_[14964]_  = (~\new_[10263]_  | ~\new_[15746]_ ) & (~\new_[16077]_  | ~n17335);
  assign \new_[14965]_  = (~\new_[15569]_  | ~\new_[9991]_ ) & (~\new_[20375]_  | ~\new_[10528]_ );
  assign \new_[14966]_  = (~\new_[16191]_  | ~\new_[9985]_ ) & (~\new_[9993]_  | ~\new_[15746]_ );
  assign \new_[14967]_  = ~\new_[15738]_  | ~\new_[17266]_  | ~\new_[17750]_  | ~wbs_we_i;
  assign n15555 = ~\new_[15868]_  | ~\new_[15225]_ ;
  assign \new_[14969]_  = wishbone_slave_unit_pci_initiator_if_last_transfered_reg;
  assign \new_[14970]_  = \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[0] ;
  assign \new_[14971]_  = ~\new_[15572]_  & (~\new_[16786]_  | ~\new_[16465]_ );
  assign \new_[14972]_  = \new_[15570]_  ? \new_[19906]_  : \new_[5043]_ ;
  assign \new_[14973]_  = ~\new_[17184]_  | ~\new_[15363]_  | ~\new_[17077]_ ;
  assign \new_[14974]_  = \new_[6306]_  ^ \new_[15579]_ ;
  assign \new_[14975]_  = \wbm_adr_o[14]  ^ \new_[15580]_ ;
  assign \new_[14976]_  = \wbm_adr_o[6]  ? \new_[15502]_  : \new_[15790]_ ;
  assign n15550 = ~\new_[15394]_  & ~\new_[15836]_ ;
  assign \new_[14978]_  = ~\new_[15409]_  & ~\new_[19906]_ ;
  assign \new_[14979]_  = ~\new_[17462]_  | ~\new_[17573]_  | ~\new_[15403]_  | ~\new_[16979]_ ;
  assign \new_[14980]_  = \new_[5010]_  ^ \new_[15413]_ ;
  assign \new_[14981]_  = ~\new_[15404]_  | (~\new_[15638]_  & ~\new_[6315]_ );
  assign \new_[14982]_  = ~\new_[15405]_  | (~\new_[15706]_  & ~\wbm_adr_o[17] );
  assign \new_[14983]_  = \wbm_adr_o[9]  ? \new_[15502]_  : \new_[15596]_ ;
  assign \new_[14984]_  = \wbm_adr_o[5]  ? \new_[15502]_  : \new_[15947]_ ;
  assign \new_[14985]_  = \new_[5040]_  ^ \new_[15586]_ ;
  assign \new_[14986]_  = \new_[6309]_  ^ \new_[15425]_ ;
  assign \new_[14987]_  = \new_[5038]_  ^ \new_[15937]_ ;
  assign \new_[14988]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[7] ;
  assign \new_[14989]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[9] ;
  assign \new_[14990]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[4] ;
  assign \new_[14991]_  = \\pci_target_unit_pci_target_if_strd_address_reg[1] ;
  assign \new_[14992]_  = \\pci_target_unit_pci_target_if_strd_address_reg[8] ;
  assign \new_[14993]_  = \\pci_target_unit_pci_target_if_strd_address_reg[6] ;
  assign \new_[14994]_  = \new_[4971]_  ^ \new_[15606]_ ;
  assign \new_[14995]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[6] ;
  assign \new_[14996]_  = \new_[15426]_  & \new_[15740]_ ;
  assign \new_[14997]_  = \new_[15844]_  | \new_[15845]_  | \new_[17422]_  | \new_[17127]_ ;
  assign \new_[14998]_  = ~\new_[15445]_  & ~\new_[19906]_ ;
  assign \new_[14999]_  = ~\new_[15444]_  & ~\new_[19906]_ ;
  assign \new_[15000]_  = ~\new_[15442]_  & ~\new_[17323]_ ;
  assign \new_[15001]_  = ~\new_[16505]_  | ~\new_[16504]_  | ~\new_[15622]_  | ~\new_[15623]_ ;
  assign \new_[15002]_  = ~\new_[15840]_  | ~\new_[16214]_  | ~\new_[16379]_  | ~\new_[15849]_ ;
  assign \new_[15003]_  = (~\new_[15952]_  | ~\new_[15976]_ ) & (~\new_[15617]_  | ~\new_[16863]_ );
  assign \new_[15004]_  = ~\new_[16995]_  | (~\new_[15601]_  & ~\new_[15821]_ );
  assign \new_[15005]_  = ~\new_[15435]_  | (~\new_[15823]_  & ~\new_[6314]_ );
  assign \new_[15006]_  = ~\new_[15439]_  | (~\new_[15824]_  & ~\wbm_adr_o[24] );
  assign \new_[15007]_  = ~\new_[15447]_  & ~\new_[20290]_ ;
  assign \new_[15008]_  = \new_[13801]_  ^ \new_[15680]_ ;
  assign \new_[15009]_  = \new_[18189]_  ^ \new_[15681]_ ;
  assign \new_[15010]_  = ~\new_[19940]_  & ~\new_[15548]_ ;
  assign \new_[15011]_  = ~\new_[5008]_  | ~\new_[19906]_ ;
  assign \new_[15012]_  = ~\new_[16473]_  & ~\new_[19906]_ ;
  assign \new_[15013]_  = ~\new_[15453]_  | ~\wbm_adr_o[27] ;
  assign \new_[15014]_  = ~\new_[15852]_  & ~\new_[19906]_ ;
  assign \new_[15015]_  = pci_target_unit_pci_target_sm_cnf_progress_reg;
  assign \new_[15016]_  = ~\new_[19924]_ ;
  assign \new_[15017]_  = ~\new_[15460]_  | ~\new_[15686]_ ;
  assign \new_[15018]_  = ~\new_[9282]_  | ~\new_[16890]_  | ~\new_[15634]_ ;
  assign \new_[15019]_  = ~\new_[17145]_  & ~\new_[15447]_ ;
  assign \new_[15020]_  = ~\new_[15454]_  & ~\new_[17195]_ ;
  assign \new_[15021]_  = ~\new_[15450]_  | (~\new_[15838]_  & ~\wbm_adr_o[19] );
  assign \new_[15022]_  = (~\new_[16905]_  | ~\new_[16194]_ ) & (~\new_[16079]_  | ~\new_[18968]_ );
  assign n15560 = pci_inta_oe_o ? \new_[17707]_  : \new_[15631]_ ;
  assign \new_[15024]_  = ~wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg;
  assign \new_[15025]_  = ~\new_[15561]_  | ~\new_[15634]_ ;
  assign \new_[15026]_  = \new_[20198]_  & \new_[16988]_ ;
  assign \new_[15027]_  = ~\new_[15518]_  | ~\new_[15510]_ ;
  assign \new_[15028]_  = ~\new_[15539]_  | ~\new_[15540]_ ;
  assign \new_[15029]_  = ~\new_[15848]_  & ~\new_[15501]_ ;
  assign \new_[15030]_  = ~\new_[15503]_  | ~\new_[20211]_ ;
  assign \new_[15031]_  = ~\new_[15526]_  | ~\new_[15690]_ ;
  assign \new_[15032]_  = ~\new_[20091]_  | ~\new_[15412]_ ;
  assign \new_[15033]_  = ~\new_[16345]_  | ~\new_[15862]_  | ~\new_[15720]_  | ~\new_[16038]_ ;
  assign \new_[15034]_  = (~\new_[20298]_  | ~\new_[12417]_ ) & (~\new_[10066]_  | ~\new_[15746]_ );
  assign \new_[15035]_  = (~\new_[20298]_  | ~\new_[12428]_ ) & (~\new_[9994]_  | ~\new_[15746]_ );
  assign \new_[15036]_  = (~\new_[20298]_  | ~\new_[12422]_ ) & (~\new_[10068]_  | ~\new_[15746]_ );
  assign \new_[15037]_  = (~\new_[20298]_  | ~\new_[12022]_ ) & (~\new_[9989]_  | ~\new_[15746]_ );
  assign \new_[15038]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[3] ;
  assign \new_[15039]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[0] ;
  assign \new_[15040]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[1] ;
  assign \new_[15041]_  = wishbone_slave_unit_pci_initiator_if_rdy_out_reg;
  assign \new_[15042]_  = ~\new_[15543]_  | ~\new_[10401]_ ;
  assign \new_[15043]_  = ~\new_[15543]_  | ~\new_[10484]_ ;
  assign \new_[15044]_  = \new_[15994]_  & \new_[15561]_ ;
  assign \new_[15045]_  = ~\new_[15543]_  | ~\new_[10403]_ ;
  assign \new_[15046]_  = ~\new_[15543]_  | ~\new_[10409]_ ;
  assign \new_[15047]_  = ~\new_[15543]_  | ~\new_[10411]_ ;
  assign \new_[15048]_  = ~\new_[15543]_  | ~\new_[10410]_ ;
  assign \new_[15049]_  = ~\new_[15543]_  | ~\new_[10408]_ ;
  assign \new_[15050]_  = ~\new_[15543]_  | ~\new_[10356]_ ;
  assign \new_[15051]_  = \new_[15550]_  | \new_[16677]_ ;
  assign \new_[15052]_  = ~\new_[15564]_  & ~\new_[15900]_ ;
  assign \new_[15053]_  = ~\new_[15564]_  & ~\new_[15902]_ ;
  assign \new_[15054]_  = ~\new_[15564]_  & ~\new_[15905]_ ;
  assign \new_[15055]_  = \new_[15699]_  & \new_[16837]_ ;
  assign \new_[15056]_  = \new_[15564]_  | \new_[17258]_ ;
  assign \new_[15057]_  = ~\new_[15547]_  | ~\new_[17123]_ ;
  assign n15575 = ~\new_[15548]_  | ~\new_[15897]_ ;
  assign \new_[15059]_  = ~\new_[15564]_  & ~\new_[15898]_ ;
  assign \new_[15060]_  = \new_[16147]_  | \new_[15563]_ ;
  assign \new_[15061]_  = ~\new_[15544]_  | ~\new_[16678]_ ;
  assign \new_[15062]_  = (~\new_[15742]_  | ~\new_[9906]_ ) & (~\new_[15876]_  | ~\new_[15892]_ );
  assign \new_[15063]_  = \new_[16424]_  | \new_[15563]_ ;
  assign \new_[15064]_  = \new_[15563]_  | \new_[16146]_ ;
  assign \new_[15065]_  = \new_[15563]_  | \new_[16418]_ ;
  assign \new_[15066]_  = \new_[16152]_  | \new_[15563]_ ;
  assign \new_[15067]_  = \new_[16151]_  | \new_[15563]_ ;
  assign \new_[15068]_  = (~\new_[16191]_  | ~\new_[16573]_ ) & (~\new_[15744]_  | ~\new_[10002]_ );
  assign \new_[15069]_  = ~\new_[15542]_  & (~\new_[10412]_  | ~\new_[16079]_ );
  assign \new_[15070]_  = (~\new_[16575]_  | ~\new_[15735]_ ) & (~\new_[15744]_  | ~\new_[9997]_ );
  assign \new_[15071]_  = (~n17430 | ~\new_[15744]_ ) & (~\new_[15735]_  | ~\new_[16574]_ );
  assign \new_[15072]_  = ~\\pci_target_unit_pci_target_if_norm_address_reg[1] ;
  assign \new_[15073]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[2] ;
  assign \new_[15074]_  = (~\new_[10010]_  | ~\new_[15735]_ ) & (~\new_[15744]_  | ~\new_[9998]_ );
  assign \new_[15075]_  = (~\new_[3738]_  | ~\new_[15744]_ ) & (~\new_[20158]_  | ~\new_[17525]_ );
  assign \new_[15076]_  = (~\new_[20092]_  | ~\new_[12340]_ ) & (~\new_[12266]_  | ~\new_[20450]_ );
  assign \new_[15077]_  = (~\new_[10005]_  | ~\new_[15744]_ ) & (~\new_[20158]_  | ~\new_[17563]_ );
  assign \new_[15078]_  = (~\new_[20092]_  | ~\new_[11960]_ ) & (~\new_[11963]_  | ~\new_[20450]_ );
  assign \new_[15079]_  = (~\new_[10009]_  | ~\new_[15744]_ ) & (~\new_[20158]_  | ~\new_[17491]_ );
  assign \new_[15080]_  = (~\new_[20092]_  | ~\new_[12035]_ ) & (~\new_[12198]_  | ~\new_[20450]_ );
  assign \new_[15081]_  = (~\new_[4267]_  | ~\new_[15744]_ ) & (~\new_[20158]_  | ~\new_[17783]_ );
  assign \new_[15082]_  = (~\new_[20092]_  | ~\new_[12305]_ ) & (~\new_[11957]_  | ~\new_[20450]_ );
  assign \new_[15083]_  = (~\new_[12040]_  | ~\new_[20450]_ ) & (~\new_[15888]_  | ~\new_[10407]_ );
  assign \new_[15084]_  = (~\new_[11981]_  | ~\new_[20056]_ ) & (~\new_[15744]_  | ~\new_[10046]_ );
  assign \new_[15085]_  = (~\new_[10007]_  | ~\new_[15744]_ ) & (~\new_[20158]_  | ~\new_[17739]_ );
  assign \new_[15086]_  = (~\new_[12268]_  | ~\new_[20450]_ ) & (~\new_[15888]_  | ~\new_[10483]_ );
  assign \new_[15087]_  = (~\new_[20092]_  | ~\new_[12367]_ ) & (~\new_[12267]_  | ~\new_[20450]_ );
  assign \new_[15088]_  = (~\new_[20092]_  | ~\new_[12036]_ ) & (~\new_[12042]_  | ~\new_[20450]_ );
  assign \new_[15089]_  = (~\new_[9907]_  | ~\new_[20450]_ ) & (~\new_[15749]_  | ~\new_[9995]_ );
  assign \new_[15090]_  = ~\new_[15320]_ ;
  assign \new_[15091]_  = ~\\pci_target_unit_pci_target_if_norm_address_reg[3] ;
  assign \new_[15092]_  = \\pci_target_unit_pci_target_if_norm_bc_reg[1] ;
  assign \new_[15093]_  = \new_[10534]_  ^ \new_[16194]_ ;
  assign \new_[15094]_  = ~\new_[15330]_ ;
  assign \new_[15095]_  = \\pci_target_unit_wishbone_master_pcir_fifo_control_out_reg[1] ;
  assign \new_[15096]_  = ~\new_[15588]_  & ~n16755;
  assign \new_[15097]_  = \\pci_target_unit_pci_target_if_strd_address_reg[4] ;
  assign \new_[15098]_  = ~\new_[15572]_  | ~\new_[17971]_ ;
  assign n15580 = n15710 | \new_[16194]_ ;
  assign \new_[15100]_  = ~\new_[15578]_  | ~\new_[16078]_ ;
  assign n15565 = ~\new_[15874]_  | ~\new_[15568]_ ;
  assign n15585 = ~\new_[15568]_  | (~\new_[16852]_  & ~\new_[16572]_ );
  assign n15570 = ~\new_[15575]_  | ~\new_[16064]_ ;
  assign \new_[15104]_  = \new_[15783]_  ? \new_[16795]_  : \new_[19274]_ ;
  assign \new_[15105]_  = \\pci_target_unit_pci_target_if_strd_address_reg[7] ;
  assign \new_[15106]_  = \new_[15783]_  ? \new_[16794]_  : \new_[18228]_ ;
  assign \new_[15107]_  = \\pci_target_unit_pci_target_if_strd_address_reg[9] ;
  assign \new_[15108]_  = \new_[15783]_  ? \new_[16803]_  : \new_[18725]_ ;
  assign \new_[15109]_  = \new_[15783]_  ? \new_[16783]_  : \new_[18807]_ ;
  assign \new_[15110]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[5] ;
  assign \new_[15111]_  = \new_[13684]_  ^ \new_[15787]_ ;
  assign \new_[15112]_  = \new_[4967]_  ^ \new_[15786]_ ;
  assign \new_[15113]_  = \new_[18100]_  ^ \new_[15788]_ ;
  assign \new_[15114]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[1] ;
  assign \new_[15115]_  = \new_[18215]_  ? \new_[16784]_  : \new_[15783]_ ;
  assign \new_[15116]_  = \new_[4963]_  ^ \new_[15785]_ ;
  assign \new_[15117]_  = \new_[18188]_  ? \new_[16984]_  : \new_[15783]_ ;
  assign \new_[15118]_  = ~\\pci_target_unit_pci_target_if_norm_address_reg[6] ;
  assign \new_[15119]_  = \new_[19261]_  ? \new_[16789]_  : \new_[15783]_ ;
  assign \new_[15120]_  = \\pci_target_unit_pci_target_if_strd_address_reg[5] ;
  assign \new_[15121]_  = \new_[15579]_  & \new_[17119]_ ;
  assign \new_[15122]_  = ~\new_[15583]_  | ~\new_[6328]_ ;
  assign \new_[15123]_  = \\pci_target_unit_del_sync_comp_cycle_count_reg[0] ;
  assign \new_[15124]_  = ~\new_[15585]_  & ~\new_[19906]_ ;
  assign \new_[15125]_  = ~\new_[15582]_  | ~\wbm_adr_o[18] ;
  assign \new_[15126]_  = ~\new_[15584]_  | ~\wbm_adr_o[22] ;
  assign \new_[15127]_  = ~\new_[17156]_  | ~\new_[17186]_  | ~\new_[15579]_  | ~\new_[17119]_ ;
  assign \new_[15128]_  = ~\new_[17186]_  | ~\new_[15579]_  | ~\new_[16737]_ ;
  assign \new_[15129]_  = \new_[16013]_  | \new_[15810]_ ;
  assign \new_[15130]_  = \new_[16384]_  | \new_[15810]_ ;
  assign \new_[15131]_  = \new_[16100]_  | \new_[15810]_ ;
  assign \new_[15132]_  = \new_[15928]_  | \new_[15810]_ ;
  assign \new_[15133]_  = ~\new_[15582]_  & ~\new_[16756]_ ;
  assign \new_[15134]_  = \new_[16435]_  | \new_[15810]_ ;
  assign \new_[15135]_  = ~\new_[17120]_  | ~\new_[15580]_  | ~\new_[16842]_ ;
  assign \new_[15136]_  = \new_[15941]_  | \new_[15810]_ ;
  assign \new_[15137]_  = \new_[16144]_  | \new_[15810]_ ;
  assign \new_[15138]_  = \new_[16440]_  | \new_[15810]_ ;
  assign \new_[15139]_  = \new_[16210]_  | \new_[15810]_ ;
  assign \new_[15140]_  = \new_[15989]_  | \new_[15810]_ ;
  assign \new_[15141]_  = \new_[15924]_  | \new_[15810]_ ;
  assign \new_[15142]_  = \new_[15927]_  | \new_[15810]_ ;
  assign \new_[15143]_  = \new_[16032]_  | \new_[15810]_ ;
  assign \new_[15144]_  = \new_[13704]_  ^ \new_[15796]_ ;
  assign \new_[15145]_  = \new_[16443]_  | \new_[15810]_ ;
  assign \new_[15146]_  = \new_[18595]_  ^ \new_[15798]_ ;
  assign \new_[15147]_  = \new_[16369]_  | \new_[15810]_ ;
  assign \new_[15148]_  = \new_[16143]_  | \new_[15810]_ ;
  assign \new_[15149]_  = ~\\pci_target_unit_pci_target_if_norm_address_reg[2] ;
  assign \new_[15150]_  = ~\new_[17136]_  | ~\new_[17177]_  | ~\new_[15422]_  | ~\new_[17078]_ ;
  assign \new_[15151]_  = \new_[18711]_  ? \new_[16883]_  : \new_[15783]_ ;
  assign \new_[15152]_  = ~\new_[15414]_  | ~\wbm_adr_o[25] ;
  assign \new_[15153]_  = ~\new_[15946]_  & ~\new_[19906]_ ;
  assign \new_[15154]_  = ~\new_[15415]_  & ~\new_[19906]_ ;
  assign n15590 = ~\new_[15428]_  & ~\new_[15836]_ ;
  assign \new_[15156]_  = ~\new_[15504]_  & ~\new_[16758]_ ;
  assign \new_[15157]_  = \new_[6305]_  ^ \new_[15803]_ ;
  assign \new_[15158]_  = \wbm_adr_o[13]  ^ \new_[15804]_ ;
  assign \new_[15159]_  = \new_[6312]_  ^ \new_[15805]_ ;
  assign \new_[15160]_  = \\pci_target_unit_pci_target_if_norm_address_reg[11] ;
  assign \new_[15161]_  = \\pci_target_unit_del_sync_addr_out_reg[22] ;
  assign \new_[15162]_  = \new_[15985]_  | \new_[16171]_ ;
  assign \new_[15163]_  = \\pci_target_unit_del_sync_addr_out_reg[21] ;
  assign \new_[15164]_  = \\pci_target_unit_del_sync_bc_out_reg[1] ;
  assign \new_[15165]_  = \\pci_target_unit_pci_target_if_norm_address_reg[16] ;
  assign \new_[15166]_  = \\pci_target_unit_pci_target_if_norm_address_reg[22] ;
  assign \new_[15167]_  = \\pci_target_unit_pci_target_if_norm_address_reg[23] ;
  assign \new_[15168]_  = \\pci_target_unit_pci_target_if_norm_address_reg[24] ;
  assign \new_[15169]_  = \\pci_target_unit_pci_target_if_norm_address_reg[25] ;
  assign \new_[15170]_  = \\pci_target_unit_del_sync_addr_out_reg[16] ;
  assign \new_[15171]_  = \\pci_target_unit_pci_target_if_norm_address_reg[17] ;
  assign \new_[15172]_  = \\pci_target_unit_pci_target_if_norm_address_reg[10] ;
  assign \new_[15173]_  = ~\\pci_target_unit_del_sync_be_out_reg[1] ;
  assign \new_[15174]_  = \\pci_target_unit_pci_target_if_norm_address_reg[30] ;
  assign \new_[15175]_  = \\input_register_pci_cbe_reg_out_reg[3] ;
  assign \new_[15176]_  = \\pci_target_unit_pci_target_if_norm_address_reg[14] ;
  assign \new_[15177]_  = \\input_register_pci_cbe_reg_out_reg[2] ;
  assign \new_[15178]_  = \\pci_target_unit_pci_target_if_norm_address_reg[28] ;
  assign \new_[15179]_  = \\pci_target_unit_pci_target_if_norm_address_reg[27] ;
  assign \new_[15180]_  = \\pci_target_unit_pci_target_if_norm_address_reg[13] ;
  assign \new_[15181]_  = \\pci_target_unit_pci_target_if_norm_bc_reg[3] ;
  assign \new_[15182]_  = \\pci_target_unit_pci_target_if_norm_bc_reg[2] ;
  assign \new_[15183]_  = \\pci_target_unit_del_sync_addr_out_reg[2] ;
  assign n16745 = wishbone_slave_unit_pci_initiator_sm_mabort1_reg;
  assign \new_[15185]_  = \\pci_target_unit_del_sync_addr_out_reg[26] ;
  assign \new_[15186]_  = \\pci_target_unit_del_sync_addr_out_reg[25] ;
  assign \new_[15187]_  = \\pci_target_unit_del_sync_addr_out_reg[24] ;
  assign \new_[15188]_  = \\pci_target_unit_del_sync_addr_out_reg[23] ;
  assign \new_[15189]_  = \\pci_target_unit_del_sync_addr_out_reg[28] ;
  assign \new_[15190]_  = \\pci_target_unit_del_sync_addr_out_reg[20] ;
  assign \new_[15191]_  = pci_target_unit_del_sync_burst_out_reg;
  assign \new_[15192]_  = \\pci_target_unit_del_sync_addr_out_reg[4] ;
  assign \new_[15193]_  = ~\\pci_target_unit_pci_target_if_norm_address_reg[5] ;
  assign \new_[15194]_  = \\pci_target_unit_del_sync_addr_out_reg[7] ;
  assign \new_[15195]_  = \\pci_target_unit_pci_target_if_norm_address_reg[21] ;
  assign \new_[15196]_  = \\pci_target_unit_pci_target_if_norm_address_reg[12] ;
  assign \new_[15197]_  = \\pci_target_unit_pci_target_if_norm_address_reg[31] ;
  assign \new_[15198]_  = \\pci_target_unit_pci_target_if_norm_address_reg[26] ;
  assign \new_[15199]_  = input_register_pci_trdy_reg_out_reg;
  assign \new_[15200]_  = \\pci_target_unit_pci_target_if_norm_address_reg[15] ;
  assign \new_[15201]_  = \\pci_target_unit_del_sync_addr_out_reg[27] ;
  assign \new_[15202]_  = ~\new_[16194]_  | ~\new_[17455]_ ;
  assign \new_[15203]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[13] ;
  assign \new_[15204]_  = \\pci_target_unit_del_sync_addr_out_reg[9] ;
  assign \new_[15205]_  = \new_[15743]_  | \new_[16618]_ ;
  assign \new_[15206]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[21] ;
  assign \new_[15207]_  = \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[3] ;
  assign \new_[15208]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[20] ;
  assign \new_[15209]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[27] ;
  assign \new_[15210]_  = \\pci_target_unit_del_sync_addr_out_reg[31] ;
  assign \new_[15211]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[8] ;
  assign \new_[15212]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[4] ;
  assign \new_[15213]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[6] ;
  assign \new_[15214]_  = \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[1] ;
  assign \new_[15215]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[29] ;
  assign \new_[15216]_  = \\input_register_pci_cbe_reg_out_reg[1] ;
  assign \new_[15217]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[30] ;
  assign \new_[15218]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[26] ;
  assign \new_[15219]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[22] ;
  assign \new_[15220]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[18] ;
  assign \new_[15221]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[12] ;
  assign \new_[15222]_  = \\pci_target_unit_pci_target_if_norm_address_reg[29] ;
  assign n15610 = ~\new_[15608]_  & ~\new_[15836]_ ;
  assign \new_[15224]_  = ~\\pci_target_unit_del_sync_be_out_reg[2] ;
  assign \new_[15225]_  = ~\new_[20151]_  | ~\new_[15605]_  | ~\new_[16572]_ ;
  assign \new_[15226]_  = \new_[15607]_  & \new_[9676]_ ;
  assign \new_[15227]_  = ~\new_[15603]_  & (~\new_[16774]_  | ~wbm_rty_i);
  assign \new_[15228]_  = ~\new_[15603]_  & (~\new_[15930]_  | ~wbm_rty_i);
  assign \new_[15229]_  = ~\new_[15603]_  & (~\new_[15851]_  | ~wbm_rty_i);
  assign \new_[15230]_  = \\pci_target_unit_pci_target_if_norm_address_reg[20] ;
  assign \new_[15231]_  = \\pci_target_unit_del_sync_addr_out_reg[1] ;
  assign \new_[15232]_  = \\pci_target_unit_del_sync_addr_out_reg[14] ;
  assign \new_[15233]_  = \\pci_target_unit_del_sync_addr_out_reg[6] ;
  assign \new_[15234]_  = \new_[4969]_  ^ \new_[15822]_ ;
  assign \new_[15235]_  = \new_[4964]_  ^ \new_[15818]_ ;
  assign \new_[15236]_  = \\pci_target_unit_del_sync_addr_out_reg[11] ;
  assign \new_[15237]_  = \wbm_adr_o[16]  ^ \new_[15815]_ ;
  assign \new_[15238]_  = \new_[6308]_  ^ \new_[15817]_ ;
  assign \new_[15239]_  = ~\new_[15621]_  | ~\new_[6316]_ ;
  assign \new_[15240]_  = ~\new_[16645]_  | ~\new_[17188]_  | ~\new_[16999]_  | ~\new_[15834]_ ;
  assign \new_[15241]_  = ~\new_[17104]_  | ~\new_[17170]_  | ~\new_[16515]_  | ~\new_[15830]_ ;
  assign \new_[15242]_  = ~\new_[15614]_  | (~\new_[15970]_  & ~\new_[6310]_ );
  assign \new_[15243]_  = ~\new_[15615]_  | (~\new_[15977]_  & ~\new_[6311]_ );
  assign \new_[15244]_  = ~\new_[15616]_  | (~\new_[15971]_  & ~\new_[6313]_ );
  assign \new_[15245]_  = ~\new_[15620]_  | (~\new_[15978]_  & ~\wbm_adr_o[20] );
  assign \new_[15246]_  = \new_[4968]_  ^ \new_[15850]_ ;
  assign \new_[15247]_  = ~\\pci_target_unit_del_sync_be_out_reg[3] ;
  assign \new_[15248]_  = \wbm_adr_o[23]  ^ \new_[15835]_ ;
  assign \new_[15249]_  = \wbm_adr_o[15]  ^ \new_[15831]_ ;
  assign \new_[15250]_  = \new_[6307]_  ^ \new_[15834]_ ;
  assign \new_[15251]_  = \new_[5039]_  ^ \new_[15830]_ ;
  assign \new_[15252]_  = ~wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg;
  assign \new_[15253]_  = \new_[17207]_  | \new_[15488]_ ;
  assign \new_[15254]_  = ~\new_[9617]_  & ~\new_[15632]_ ;
  assign \new_[15255]_  = ~\new_[16221]_  | ~\new_[15633]_ ;
  assign \new_[15256]_  = ~\new_[16076]_  | ~\new_[15745]_  | ~\new_[15855]_ ;
  assign \new_[15257]_  = ~\new_[19201]_  | ~\new_[16577]_  | ~\new_[15683]_  | ~\new_[20421]_ ;
  assign \new_[15258]_  = ~\new_[15488]_  & (~\new_[17095]_  | ~\new_[17255]_ );
  assign \new_[15259]_  = ~n16095 & (~\new_[15994]_  | ~\new_[16171]_ );
  assign n15600 = \new_[17258]_  ? \new_[17707]_  : \new_[17403]_ ;
  assign \new_[15261]_  = (~\new_[15854]_  | ~\new_[10063]_ ) & (~\new_[12299]_  | ~\new_[19956]_ );
  assign \new_[15262]_  = (~\new_[15854]_  | ~\new_[10365]_ ) & (~\new_[12076]_  | ~\new_[19956]_ );
  assign \new_[15263]_  = ~\new_[15465]_ ;
  assign \new_[15264]_  = ~\new_[15469]_ ;
  assign \new_[15265]_  = ~\new_[15470]_ ;
  assign \new_[15266]_  = ~\new_[15471]_ ;
  assign \new_[15267]_  = ~\new_[15473]_ ;
  assign \new_[15268]_  = \\pci_target_unit_del_sync_addr_out_reg[19] ;
  assign \new_[15269]_  = (~\new_[15854]_  | ~\new_[10064]_ ) & (~\new_[12075]_  | ~\new_[19956]_ );
  assign \new_[15270]_  = \\pci_target_unit_del_sync_addr_out_reg[15] ;
  assign \new_[15271]_  = \new_[15791]_  & \new_[16073]_ ;
  assign \new_[15272]_  = \\pci_target_unit_del_sync_addr_out_reg[30] ;
  assign \new_[15273]_  = ~\new_[15487]_ ;
  assign \new_[15274]_  = ~\new_[15487]_ ;
  assign \new_[15275]_  = ~\new_[15487]_ ;
  assign \new_[15276]_  = ~\new_[15699]_  | ~\new_[17033]_ ;
  assign \new_[15277]_  = \new_[15994]_  | \new_[17793]_ ;
  assign \new_[15278]_  = ~\new_[15684]_  | ~\new_[15856]_ ;
  assign \new_[15279]_  = ~\new_[17272]_  | ~wbs_stb_i | ~\new_[15739]_  | ~\new_[17266]_ ;
  assign n15615 = \new_[15912]_  & \new_[15994]_ ;
  assign \new_[15281]_  = ~\new_[16915]_  | ~\new_[16072]_  | ~\new_[16922]_  | ~\new_[16913]_ ;
  assign \new_[15282]_  = ~\new_[15889]_  & (~\new_[20158]_  | ~\new_[17611]_ );
  assign \new_[15283]_  = (~\new_[15890]_  | ~\new_[9905]_ ) & (~\new_[12059]_  | ~\new_[20056]_ );
  assign \new_[15284]_  = \\pci_target_unit_del_sync_addr_out_reg[8] ;
  assign \new_[15285]_  = \\pci_target_unit_del_sync_addr_out_reg[3] ;
  assign \new_[15286]_  = ~\new_[15603]_  & (~\new_[16483]_  | ~wbm_rty_i);
  assign \new_[15287]_  = \\pci_target_unit_pci_target_if_norm_address_reg[19] ;
  assign \new_[15288]_  = ~\new_[15681]_  & ~\new_[17472]_ ;
  assign \new_[15289]_  = (~\new_[11964]_  | ~\new_[19956]_ ) & (~\new_[20158]_  | ~\new_[17677]_ );
  assign \new_[15290]_  = ~\new_[15505]_ ;
  assign \new_[15291]_  = (~\new_[10858]_  | ~\new_[20506]_ ) & (~\new_[20175]_  | ~\new_[10491]_ );
  assign \new_[15292]_  = (~\new_[15888]_  | ~\new_[10399]_ ) & (~\new_[20494]_  | ~\new_[10520]_ );
  assign \new_[15293]_  = (~\new_[12331]_  | ~\new_[19956]_ ) & (~\new_[20158]_  | ~\new_[17594]_ );
  assign \new_[15294]_  = (~\new_[10864]_  | ~\new_[20506]_ ) & (~\new_[20494]_  | ~\new_[10493]_ );
  assign \new_[15295]_  = (~\new_[12069]_  | ~\new_[19956]_ ) & (~\new_[20158]_  | ~\new_[17541]_ );
  assign \new_[15296]_  = (~\new_[15888]_  | ~\new_[10402]_ ) & (~\new_[20175]_  | ~\new_[10521]_ );
  assign \new_[15297]_  = (~\new_[12070]_  | ~\new_[19956]_ ) & (~\new_[20158]_  | ~\new_[17530]_ );
  assign \new_[15298]_  = (~\new_[15888]_  | ~\new_[10486]_ ) & (~\new_[20494]_  | ~\new_[10523]_ );
  assign \new_[15299]_  = (~\new_[12071]_  | ~\new_[19956]_ ) & (~\new_[20158]_  | ~\new_[17784]_ );
  assign \new_[15300]_  = \\pci_target_unit_del_sync_addr_out_reg[13] ;
  assign \new_[15301]_  = (~\new_[10857]_  | ~\new_[20506]_ ) & (~\new_[20494]_  | ~\new_[10527]_ );
  assign \new_[15302]_  = (~\new_[10866]_  | ~\new_[20506]_ ) & (~\new_[20494]_  | ~\new_[10529]_ );
  assign \new_[15303]_  = \\pci_target_unit_pci_target_if_norm_address_reg[18] ;
  assign \new_[15304]_  = (~\new_[12080]_  | ~\new_[19956]_ ) & (~\new_[20158]_  | ~\new_[17481]_ );
  assign \new_[15305]_  = (~\new_[12067]_  | ~\new_[19956]_ ) & (~\new_[20158]_  | ~\new_[17718]_ );
  assign \new_[15306]_  = (~\new_[15888]_  | ~\new_[10404]_ ) & (~\new_[20494]_  | ~\new_[10519]_ );
  assign \new_[15307]_  = (~\new_[20092]_  | ~\new_[12366]_ ) & (~\new_[20175]_  | ~\new_[10845]_ );
  assign \new_[15308]_  = (~\new_[15888]_  | ~\new_[10481]_ ) & (~\new_[20175]_  | ~\new_[10528]_ );
  assign \new_[15309]_  = \\pci_target_unit_del_sync_addr_out_reg[12] ;
  assign \new_[15310]_  = (~\new_[20158]_  | ~\new_[17504]_ ) & (~\new_[19956]_  | ~\new_[12494]_ );
  assign \new_[15311]_  = (~\new_[11067]_  | ~\new_[20506]_ ) & (~\new_[20494]_  | ~\new_[10848]_ );
  assign \new_[15312]_  = (~\new_[15888]_  | ~\new_[10405]_ ) & (~\new_[20175]_  | ~\new_[10492]_ );
  assign \new_[15313]_  = (~\new_[15888]_  | ~\new_[10485]_ ) & (~\new_[20175]_  | ~\new_[10514]_ );
  assign \new_[15314]_  = (~\new_[16852]_  | ~\new_[9287]_ ) & (~\new_[16446]_  | ~\new_[5047]_ );
  assign \new_[15315]_  = (~\new_[10394]_  | ~\new_[16077]_ ) & (~\new_[20158]_  | ~\new_[10528]_ );
  assign \new_[15316]_  = (~\new_[12420]_  | ~\new_[19957]_ ) & (~\new_[20158]_  | ~\new_[17542]_ );
  assign \new_[15317]_  = (~\new_[20092]_  | ~\new_[12413]_ ) & (~\new_[20175]_  | ~\new_[10515]_ );
  assign \new_[15318]_  = (~\new_[12064]_  | ~\new_[19957]_ ) & (~\new_[20158]_  | ~\new_[17570]_ );
  assign \new_[15319]_  = ~\new_[15535]_ ;
  assign \new_[15320]_  = (~\new_[11954]_  | ~\new_[19957]_ ) & (~\new_[20158]_  | ~\new_[17697]_ );
  assign \new_[15321]_  = (~\new_[10867]_  | ~\new_[20506]_ ) & (~\new_[20175]_  | ~\new_[10530]_ );
  assign \new_[15322]_  = (~\new_[10865]_  | ~\new_[20506]_ ) & (~\new_[20494]_  | ~\new_[10524]_ );
  assign \new_[15323]_  = (~\new_[11036]_  | ~\new_[20506]_ ) & (~\new_[20175]_  | ~\new_[10516]_ );
  assign \new_[15324]_  = (~\new_[12065]_  | ~\new_[19957]_ ) & (~\new_[20158]_  | ~\new_[20378]_ );
  assign \new_[15325]_  = (~\new_[15888]_  | ~\new_[10398]_ ) & (~\new_[20175]_  | ~\new_[10518]_ );
  assign \new_[15326]_  = (~\new_[12066]_  | ~\new_[19957]_ ) & (~\new_[20158]_  | ~\new_[17485]_ );
  assign \new_[15327]_  = (~\new_[15888]_  | ~\new_[10395]_ ) & (~\new_[20494]_  | ~\new_[10522]_ );
  assign n15595 = \new_[17258]_  ? \new_[16362]_  : \new_[18583]_ ;
  assign \new_[15329]_  = \\pci_target_unit_del_sync_addr_out_reg[10] ;
  assign \new_[15330]_  = ~\\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0] ;
  assign \new_[15331]_  = ~pci_target_unit_pci_target_sm_state_backoff_reg_reg;
  assign \new_[15332]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[10] ;
  assign \new_[15333]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[11] ;
  assign \new_[15334]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[16] ;
  assign \new_[15335]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[19] ;
  assign \new_[15336]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[23] ;
  assign \new_[15337]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[28] ;
  assign \new_[15338]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[2] ;
  assign \new_[15339]_  = \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[2] ;
  assign \new_[15340]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[3] ;
  assign \new_[15341]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[5] ;
  assign \new_[15342]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[7] ;
  assign \new_[15343]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[9] ;
  assign \new_[15344]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[31] ;
  assign \new_[15345]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[24] ;
  assign \new_[15346]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[14] ;
  assign \new_[15347]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[15] ;
  assign \new_[15348]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[25] ;
  assign \new_[15349]_  = \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[17] ;
  assign n15605 = ~\new_[15794]_  & ~\new_[15836]_ ;
  assign \new_[15351]_  = \new_[15885]_  & \new_[15741]_ ;
  assign \new_[15352]_  = ~\new_[15889]_  & ~\new_[15746]_ ;
  assign \new_[15353]_  = ~\new_[15680]_  & ~\new_[17649]_ ;
  assign \new_[15354]_  = \new_[20081]_  | \new_[15743]_ ;
  assign \new_[15355]_  = ~\new_[15743]_  & ~\new_[17971]_ ;
  assign \new_[15356]_  = ~\new_[15784]_  & ~\new_[16949]_ ;
  assign \new_[15357]_  = \new_[16069]_  & \new_[15745]_ ;
  assign \new_[15358]_  = ~\new_[10000]_  | ~\new_[16404]_  | ~\new_[19886]_ ;
  assign \new_[15359]_  = ~\new_[20128]_  | ~\new_[20488]_  | ~\new_[15734]_  | ~\new_[16836]_ ;
  assign \new_[15360]_  = (~\new_[16402]_  | ~\new_[17680]_ ) & (~\new_[20161]_  | ~\new_[9879]_ );
  assign \new_[15361]_  = \\pci_target_unit_del_sync_bc_out_reg[3] ;
  assign \new_[15362]_  = ~\new_[15785]_  & ~\new_[16972]_ ;
  assign \new_[15363]_  = ~\new_[16708]_  & ~\new_[15785]_ ;
  assign \new_[15364]_  = \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[2] ;
  assign \new_[15365]_  = \new_[15948]_  | \new_[16171]_ ;
  assign \new_[15366]_  = \new_[15923]_  | \new_[16171]_ ;
  assign \new_[15367]_  = \new_[15925]_  | \new_[16171]_ ;
  assign \new_[15368]_  = \new_[16027]_  | \new_[16171]_ ;
  assign \new_[15369]_  = \new_[16107]_  | \new_[16171]_ ;
  assign \new_[15370]_  = \new_[16354]_  | \new_[16171]_ ;
  assign \new_[15371]_  = \new_[15926]_  | \new_[16171]_ ;
  assign \new_[15372]_  = \new_[16150]_  | \new_[16171]_ ;
  assign \new_[15373]_  = \new_[15986]_  | \new_[16171]_ ;
  assign \new_[15374]_  = \new_[16405]_  | \new_[16171]_ ;
  assign \new_[15375]_  = \new_[16382]_  | \new_[16171]_ ;
  assign \new_[15376]_  = \new_[16134]_  | \new_[16171]_ ;
  assign \new_[15377]_  = \new_[16127]_  | \new_[16171]_ ;
  assign \new_[15378]_  = \new_[16414]_  | \new_[16171]_ ;
  assign \new_[15379]_  = ~\new_[17184]_  | ~\new_[16132]_  | ~\new_[16585]_  | ~\new_[17176]_ ;
  assign \new_[15380]_  = \new_[6304]_  ^ \new_[15909]_ ;
  assign \new_[15381]_  = \wbm_adr_o[10]  ^ \new_[15910]_ ;
  assign \new_[15382]_  = ~\new_[15573]_ ;
  assign \new_[15383]_  = ~\new_[15746]_ ;
  assign \new_[15384]_  = ~\new_[16103]_  & (~\new_[17304]_  | ~\new_[10371]_ );
  assign \new_[15385]_  = ~\\pci_target_unit_pci_target_if_norm_address_reg[9] ;
  assign n15620 = \new_[14208]_  ? \new_[16415]_  : \new_[17258]_ ;
  assign \new_[15387]_  = \\pci_target_unit_del_sync_addr_out_reg[5] ;
  assign \new_[15388]_  = ~\new_[15792]_  & ~\new_[12039]_ ;
  assign \new_[15389]_  = ~\\pci_target_unit_pci_target_if_norm_address_reg[4] ;
  assign \new_[15390]_  = ~\\pci_target_unit_pci_target_if_norm_address_reg[0] ;
  assign \new_[15391]_  = ~\new_[15603]_  & (~\new_[15932]_  | ~wbm_rty_i);
  assign \new_[15392]_  = ~\\pci_target_unit_pci_target_if_norm_address_reg[8] ;
  assign \new_[15393]_  = \\pci_target_unit_pci_target_if_strd_address_reg[0] ;
  assign \new_[15394]_  = \new_[13821]_  ^ \new_[15828]_ ;
  assign \new_[15395]_  = \new_[18509]_  ^ \new_[15825]_ ;
  assign \new_[15396]_  = ~\\pci_target_unit_pci_target_if_norm_address_reg[7] ;
  assign \new_[15397]_  = ~\new_[17033]_  & ~\new_[16836]_ ;
  assign \new_[15398]_  = \\pci_target_unit_del_sync_bc_out_reg[0] ;
  assign \new_[15399]_  = \\pci_target_unit_del_sync_bc_out_reg[2] ;
  assign \new_[15400]_  = \\pci_target_unit_del_sync_addr_out_reg[29] ;
  assign \new_[15401]_  = \\pci_target_unit_del_sync_addr_out_reg[18] ;
  assign \new_[15402]_  = \\pci_target_unit_del_sync_addr_out_reg[0] ;
  assign \new_[15403]_  = ~\new_[15797]_  & ~\new_[16892]_ ;
  assign \new_[15404]_  = ~\new_[15638]_  | ~\new_[6315]_ ;
  assign \new_[15405]_  = ~\new_[15706]_  | ~\wbm_adr_o[17] ;
  assign \new_[15406]_  = \\pci_target_unit_del_sync_addr_out_reg[17] ;
  assign \new_[15407]_  = ~\new_[15603]_  & (~\new_[15811]_  | ~wbm_rty_i);
  assign \new_[15408]_  = \wbm_adr_o[21]  ^ \new_[15808]_ ;
  assign \new_[15409]_  = \new_[5009]_  ^ \new_[15807]_ ;
  assign \new_[15410]_  = \new_[16130]_  | \new_[16171]_ ;
  assign \new_[15411]_  = input_register_pci_frame_reg_out_reg;
  assign \new_[15412]_  = ~\new_[20494]_  | ~\new_[10847]_ ;
  assign \new_[15413]_  = ~\new_[16979]_  | ~\new_[16184]_  | ~\new_[16503]_  | ~\new_[17276]_ ;
  assign \new_[15414]_  = ~\new_[17167]_  | ~\new_[16185]_  | ~\new_[16748]_  | ~\new_[17154]_ ;
  assign \new_[15415]_  = \new_[4977]_  ^ \new_[16476]_ ;
  assign n15655 = ~\new_[16186]_  & ~\new_[15836]_ ;
  assign \new_[15417]_  = input_register_pci_devsel_reg_out_reg;
  assign \new_[15418]_  = ~\new_[15800]_  & (~\new_[16368]_  | ~\new_[17747]_ );
  assign n15680 = ~\new_[15704]_ ;
  assign \new_[15420]_  = (~\new_[16099]_  | ~\new_[9908]_ ) & (~\new_[19886]_  | ~\new_[17737]_ );
  assign pci_irdy_o = pci_io_mux_irdy_iob_dat_out_reg;
  assign \new_[15422]_  = \new_[17199]_  & \new_[15803]_ ;
  assign \new_[15423]_  = (~\new_[16191]_  | ~\new_[12006]_ ) & (~\new_[16077]_  | ~\new_[10358]_ );
  assign \new_[15424]_  = input_register_pci_irdy_reg_out_reg;
  assign \new_[15425]_  = \new_[17078]_  & \new_[15803]_ ;
  assign \new_[15426]_  = \new_[19940]_  | \new_[15897]_ ;
  assign \new_[15427]_  = \new_[9791]_  ^ \new_[15954]_ ;
  assign \new_[15428]_  = \new_[18971]_  ^ \new_[15953]_ ;
  assign \new_[15429]_  = \new_[15960]_  ^ \new_[15965]_ ;
  assign \new_[15430]_  = \new_[15961]_  ^ \new_[15963]_ ;
  assign \new_[15431]_  = \new_[15962]_  ^ \new_[15959]_ ;
  assign \new_[15432]_  = ~\new_[15821]_  & ~\new_[15837]_ ;
  assign \new_[15433]_  = ~\new_[15603]_ ;
  assign \new_[15434]_  = ~\new_[15604]_ ;
  assign \new_[15435]_  = ~\new_[15823]_  | ~\new_[6314]_ ;
  assign n15695 = ~\new_[16693]_  & ~\new_[15836]_ ;
  assign n15630 = ~\new_[15826]_  & ~\new_[15836]_ ;
  assign \new_[15438]_  = ~\new_[17181]_  | ~\new_[15814]_ ;
  assign \new_[15439]_  = ~\new_[15824]_  | ~\wbm_adr_o[24] ;
  assign \new_[15440]_  = ~\new_[15820]_  & ~\new_[16744]_ ;
  assign n15660 = ~\new_[20331]_  | (~\new_[19201]_  & ~\new_[16572]_ );
  assign \new_[15442]_  = ~\new_[15607]_ ;
  assign \new_[15443]_  = ~\new_[15819]_  & ~\new_[16736]_ ;
  assign \new_[15444]_  = \new_[4966]_  ^ \new_[15983]_ ;
  assign \new_[15445]_  = \new_[4965]_  ^ \new_[15951]_ ;
  assign \new_[15446]_  = \new_[15984]_  ^ \new_[16717]_ ;
  assign \new_[15447]_  = ~\new_[15612]_ ;
  assign n15735 = ~\new_[17112]_  & ~\new_[15836]_ ;
  assign n15730 = ~\new_[16455]_  & ~\new_[15836]_ ;
  assign \new_[15450]_  = ~\new_[15838]_  | ~\wbm_adr_o[19] ;
  assign \new_[15451]_  = \new_[15846]_  | \new_[15847]_ ;
  assign n15750 = ~\new_[15836]_  & ~\new_[15123]_ ;
  assign \new_[15453]_  = ~\new_[17168]_  | ~\new_[17161]_  | ~\new_[15831]_  | ~\new_[17162]_ ;
  assign \new_[15454]_  = ~\new_[17161]_  | ~\new_[15831]_  | ~\new_[16844]_ ;
  assign \new_[15455]_  = (~\new_[20298]_  | ~\new_[12436]_ ) & (~\new_[12068]_  | ~\new_[19957]_ );
  assign \new_[15456]_  = (~\new_[20298]_  | ~\new_[12019]_ ) & (~\new_[20049]_  | ~\new_[10486]_ );
  assign \new_[15457]_  = (~\new_[20298]_  | ~\new_[12434]_ ) & (~\new_[20049]_  | ~\new_[10399]_ );
  assign \new_[15458]_  = (~\new_[20298]_  | ~\new_[12433]_ ) & (~\new_[20049]_  | ~\new_[10404]_ );
  assign \new_[15459]_  = (~\new_[20298]_  | ~\new_[12429]_ ) & (~\new_[12509]_  | ~\new_[19957]_ );
  assign \new_[15460]_  = (~\new_[20298]_  | ~\new_[12427]_ ) & (~\new_[16191]_  | ~\new_[12412]_ );
  assign \new_[15461]_  = (~\new_[20298]_  | ~\new_[12023]_ ) & (~\new_[16191]_  | ~\new_[12437]_ );
  assign \new_[15462]_  = (~\new_[20092]_  | ~\new_[12311]_ ) & (~\new_[20298]_  | ~\new_[12024]_ );
  assign \new_[15463]_  = (~\new_[20092]_  | ~\new_[12038]_ ) & (~\new_[20298]_  | ~\new_[12383]_ );
  assign \new_[15464]_  = (~\new_[20298]_  | ~\new_[12431]_ ) & (~\new_[20049]_  | ~\new_[10485]_ );
  assign \new_[15465]_  = (~\new_[20298]_  | ~\new_[12423]_ ) & (~\new_[16191]_  | ~\new_[12008]_ );
  assign \new_[15466]_  = ~\new_[17104]_  | ~\new_[16226]_  | ~\new_[16644]_  | ~\new_[17094]_ ;
  assign \new_[15467]_  = (~\new_[20298]_  | ~\new_[12018]_ ) & (~\new_[20049]_  | ~\new_[10402]_ );
  assign \new_[15468]_  = (~\new_[20298]_  | ~\new_[12026]_ ) & (~\new_[16077]_  | ~\new_[10387]_ );
  assign \new_[15469]_  = (~\new_[20298]_  | ~\new_[12430]_ ) & (~\new_[16191]_  | ~\new_[12410]_ );
  assign \new_[15470]_  = (~\new_[20298]_  | ~\new_[12425]_ ) & (~\new_[16191]_  | ~\new_[12416]_ );
  assign \new_[15471]_  = (~\new_[20298]_  | ~\new_[12021]_ ) & (~\new_[16191]_  | ~\new_[12009]_ );
  assign \new_[15472]_  = (~\new_[20298]_  | ~\new_[12013]_ ) & (~\new_[11329]_  | ~\new_[19957]_ );
  assign \new_[15473]_  = (~\new_[20298]_  | ~\new_[12426]_ ) & (~\new_[16191]_  | ~\new_[12010]_ );
  assign \new_[15474]_  = (~\new_[20298]_  | ~\new_[12014]_ ) & (~\new_[16077]_  | ~\new_[10389]_ );
  assign \new_[15475]_  = (~\new_[20298]_  | ~\new_[12015]_ ) & (~\new_[16077]_  | ~\new_[10390]_ );
  assign \new_[15476]_  = (~\new_[20298]_  | ~\new_[12432]_ ) & (~\new_[16077]_  | ~\new_[10391]_ );
  assign \new_[15477]_  = (~\new_[20298]_  | ~\new_[12435]_ ) & (~\new_[16077]_  | ~\new_[10392]_ );
  assign \new_[15478]_  = (~\new_[20298]_  | ~\new_[12020]_ ) & (~\new_[16191]_  | ~\new_[12415]_ );
  assign \new_[15479]_  = (~\new_[20298]_  | ~\new_[12016]_ ) & (~\new_[16077]_  | ~\new_[10393]_ );
  assign \new_[15480]_  = output_backup_irdy_out_reg;
  assign n15665 = \\wishbone_slave_unit_del_sync_rty_exp_back_prop_sync_sync_data_out_reg[0] ;
  assign \new_[15482]_  = ~\new_[15854]_  | ~\new_[10062]_ ;
  assign \new_[15483]_  = ~\new_[19921]_  & ~\new_[17033]_ ;
  assign \new_[15484]_  = ~\new_[15829]_ ;
  assign \new_[15485]_  = ~\new_[15829]_ ;
  assign \new_[15486]_  = ~\new_[15795]_ ;
  assign \new_[15487]_  = ~\new_[15488]_ ;
  assign \new_[15488]_  = ~\new_[15829]_ ;
  assign \new_[15489]_  = ~\new_[15829]_ ;
  assign n16690 = pci_target_unit_del_sync_req_req_pending_reg;
  assign \new_[15491]_  = ~\new_[15795]_ ;
  assign \new_[15492]_  = ~\new_[15795]_ ;
  assign \new_[15493]_  = ~\new_[15795]_ ;
  assign \new_[15494]_  = ~\new_[15795]_ ;
  assign \new_[15495]_  = ~\new_[15795]_ ;
  assign \new_[15496]_  = ~\new_[15634]_ ;
  assign \new_[15497]_  = ~\new_[15802]_  & ~\new_[17549]_ ;
  assign \new_[15498]_  = ~\new_[19907]_ ;
  assign \new_[15499]_  = ~\new_[16106]_  & (~\new_[16577]_  | ~\new_[16734]_ );
  assign \new_[15500]_  = ~\new_[15637]_ ;
  assign \new_[15501]_  = ~\new_[16640]_  | ~\new_[16381]_  | ~\new_[16732]_  | ~\new_[16760]_ ;
  assign \new_[15502]_  = (~\new_[16374]_  & ~\new_[20218]_ ) | (~\new_[20212]_  & ~\new_[16079]_ );
  assign \new_[15503]_  = ~\new_[16596]_  | ~\new_[16193]_  | ~\new_[15918]_ ;
  assign \new_[15504]_  = ~\new_[17108]_  | ~\new_[15804]_  | ~\new_[17154]_ ;
  assign \new_[15505]_  = (~\new_[20092]_  | ~\new_[12411]_ ) & (~\new_[12048]_  | ~\new_[20056]_ );
  assign \new_[15506]_  = (~\new_[12287]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17594]_ );
  assign \new_[15507]_  = (~\new_[20092]_  | ~\new_[12404]_ ) & (~\new_[10861]_  | ~\new_[20094]_ );
  assign \new_[15508]_  = (~\new_[12049]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17541]_ );
  assign \new_[15509]_  = (~\new_[12053]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17784]_ );
  assign \new_[15510]_  = (~\new_[12050]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[20023]_ );
  assign \new_[15511]_  = (~\new_[20092]_  | ~\new_[12033]_ ) & (~\new_[10863]_  | ~\new_[20506]_ );
  assign \new_[15512]_  = (~\new_[20092]_  | ~\new_[12407]_ ) & (~\new_[11070]_  | ~\new_[20506]_ );
  assign \new_[15513]_  = (~\new_[20092]_  | ~\new_[12031]_ ) & (~\new_[10860]_  | ~\new_[20506]_ );
  assign \new_[15514]_  = (~\new_[12056]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17686]_ );
  assign \new_[15515]_  = (~\new_[12058]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17491]_ );
  assign \new_[15516]_  = (~\new_[12060]_  | ~\new_[20056]_ ) & (~\new_[12508]_  | ~\new_[19957]_ );
  assign \new_[15517]_  = (~\new_[11986]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17783]_ );
  assign \new_[15518]_  = (~\new_[20092]_  | ~\new_[12032]_ ) & (~\new_[11071]_  | ~\new_[20506]_ );
  assign \new_[15519]_  = (~\new_[11987]_  | ~\new_[20056]_ ) & (~\new_[12077]_  | ~\new_[19957]_ );
  assign \new_[15520]_  = (~\new_[12061]_  | ~\new_[20056]_ ) & (~\new_[12495]_  | ~\new_[19957]_ );
  assign \new_[15521]_  = (~\new_[20092]_  | ~\new_[12310]_ ) & (~\new_[12078]_  | ~\new_[19957]_ );
  assign \new_[15522]_  = (~\new_[12063]_  | ~\new_[20056]_ ) & (~\new_[12079]_  | ~\new_[19957]_ );
  assign \new_[15523]_  = (~\new_[11984]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17481]_ );
  assign \new_[15524]_  = (~\new_[20092]_  | ~\new_[12034]_ ) & (~\new_[20049]_  | ~\new_[10407]_ );
  assign \new_[15525]_  = (~\new_[11991]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17563]_ );
  assign \new_[15526]_  = (~\new_[11988]_  | ~\new_[20056]_ ) & (~\new_[10868]_  | ~\new_[20506]_ );
  assign \new_[15527]_  = (~\new_[20375]_  | ~\new_[17504]_ ) & (~\new_[20056]_  | ~\new_[12062]_ );
  assign \new_[15528]_  = (~\new_[12004]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17530]_ );
  assign \new_[15529]_  = (~\new_[12055]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17766]_ );
  assign \new_[15530]_  = (~\new_[11068]_  | ~\new_[20506]_ ) & (~\new_[20049]_  | ~\new_[10483]_ );
  assign \new_[15531]_  = (~\new_[12052]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17542]_ );
  assign \new_[15532]_  = (~\new_[11990]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17739]_ );
  assign \new_[15533]_  = (~\new_[16191]_  | ~\new_[12007]_ ) & (~\new_[16077]_  | ~\new_[10388]_ );
  assign \new_[15534]_  = (~\new_[12043]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17570]_ );
  assign \new_[15535]_  = (~\new_[20092]_  | ~\new_[12323]_ ) & (~\new_[12054]_  | ~\new_[20056]_ );
  assign \new_[15536]_  = (~\new_[20092]_  | ~\new_[12028]_ ) & (~\new_[10972]_  | ~\new_[20094]_ );
  assign \new_[15537]_  = (~\new_[12044]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17697]_ );
  assign \new_[15538]_  = (~\new_[11993]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17525]_ );
  assign \new_[15539]_  = (~\new_[20092]_  | ~\new_[12029]_ ) & (~\new_[11029]_  | ~\new_[20506]_ );
  assign \new_[15540]_  = (~\new_[12259]_  | ~\new_[20056]_ ) & (~\new_[20375]_  | ~\new_[17485]_ );
  assign \new_[15541]_  = ~\new_[16079]_  | ~\new_[10855]_ ;
  assign \new_[15542]_  = ~\new_[17090]_  & ~\new_[16079]_ ;
  assign \new_[15543]_  = \new_[15888]_  | \new_[20049]_ ;
  assign \new_[15544]_  = ~\new_[16446]_  | ~\new_[16618]_ ;
  assign \new_[15545]_  = ~\new_[20494]_  | ~\new_[10525]_ ;
  assign n15685 = \new_[15878]_  | \new_[17323]_ ;
  assign \new_[15547]_  = ~\new_[16577]_  & ~\new_[18325]_ ;
  assign \new_[15548]_  = ~\new_[16603]_  | ~\new_[20205]_  | ~\new_[4627]_ ;
  assign \new_[15549]_  = ~\new_[20494]_  | ~\new_[10517]_ ;
  assign \new_[15550]_  = ~\new_[16426]_  | ~\new_[20128]_  | ~\new_[15903]_  | ~\new_[16608]_ ;
  assign n15690 = ~\new_[16067]_  | (~\new_[15072]_  & ~\new_[16572]_ );
  assign n15705 = ~\new_[16432]_  | (~\new_[17383]_  & ~\new_[19929]_ );
  assign n15755 = ~\new_[16065]_  | (~\new_[15149]_  & ~\new_[16572]_ );
  assign n15700 = ~\new_[16064]_  | (~\new_[15091]_  & ~\new_[16572]_ );
  assign n15740 = ~\new_[16066]_  | (~\new_[15118]_  & ~\new_[16572]_ );
  assign n15645 = ~\new_[15877]_  | ~\new_[16063]_ ;
  assign n15725 = ~\new_[15870]_  | ~\new_[16062]_ ;
  assign n15650 = ~\new_[15872]_  | ~\new_[16066]_ ;
  assign n15745 = ~\new_[15873]_  | ~\new_[15917]_ ;
  assign n15715 = ~\new_[15871]_  | ~\new_[15914]_ ;
  assign \new_[15561]_  = \new_[15886]_  | \new_[20089]_ ;
  assign n15640 = ~\new_[16067]_  | (~\new_[20173]_  & ~\new_[16572]_ );
  assign \new_[15563]_  = ~\new_[15884]_  | ~\new_[15903]_ ;
  assign \new_[15564]_  = ~\new_[16836]_  | ~\new_[15884]_  | ~\new_[17033]_ ;
  assign n15675 = ~\new_[15599]_ ;
  assign \new_[15566]_  = (~\new_[20092]_  | ~\new_[12406]_ ) & (~\new_[10862]_  | ~\new_[20506]_ );
  assign n15635 = ~\new_[15895]_  & ~\new_[15836]_ ;
  assign \new_[15568]_  = ~\new_[17258]_  | ~\new_[16572]_ ;
  assign \new_[15569]_  = \new_[20451]_  & \new_[15892]_ ;
  assign \new_[15570]_  = \new_[5043]_  ^ \new_[16132]_ ;
  assign n15710 = ~\new_[16674]_  & ~\new_[16839]_ ;
  assign \new_[15572]_  = ~\new_[15743]_ ;
  assign \new_[15573]_  = ~\new_[15744]_ ;
  assign \new_[15574]_  = ~\new_[15747]_ ;
  assign \new_[15575]_  = ~\new_[16836]_  | ~\new_[19929]_ ;
  assign \new_[15576]_  = (~\new_[16630]_  | ~\new_[13813]_ ) & (~\new_[4092]_  | ~\new_[18584]_ );
  assign \new_[15577]_  = \new_[15907]_  & \new_[19201]_ ;
  assign \new_[15578]_  = \new_[16115]_  & \new_[16837]_ ;
  assign \new_[15579]_  = \new_[15909]_  & \new_[17109]_ ;
  assign \new_[15580]_  = \new_[15910]_  & \new_[17157]_ ;
  assign n15625 = ~\new_[15911]_  & ~\new_[15836]_ ;
  assign \new_[15582]_  = ~\new_[17155]_  | ~\new_[15910]_  | ~\new_[17157]_ ;
  assign \new_[15583]_  = ~\new_[16737]_  | ~\new_[16181]_  | ~\new_[17116]_  | ~\new_[17109]_ ;
  assign \new_[15584]_  = ~\new_[16842]_  | ~\new_[16182]_  | ~\new_[17165]_  | ~\new_[17157]_ ;
  assign \new_[15585]_  = \new_[4975]_  ^ \new_[16475]_ ;
  assign \new_[15586]_  = ~\new_[16892]_  & ~\new_[15806]_ ;
  assign n15670 = ~\new_[16173]_  & ~\new_[15836]_ ;
  assign \new_[15588]_  = ~\new_[15736]_ ;
  assign n15720 = ~\new_[15883]_  | ~\new_[15915]_ ;
  assign \new_[15590]_  = ~\new_[15795]_ ;
  assign \new_[15591]_  = ~\new_[15795]_ ;
  assign \new_[15592]_  = ~\new_[15829]_ ;
  assign \new_[15593]_  = \new_[5044]_  ^ \new_[16195]_ ;
  assign \new_[15594]_  = input_register_pci_stop_reg_out_reg;
  assign \new_[15595]_  = \new_[6325]_  ^ \new_[16183]_ ;
  assign \new_[15596]_  = \wbm_adr_o[9]  ^ \new_[16185]_ ;
  assign n16270 = ~\new_[15914]_  | (~\new_[15389]_  & ~\new_[16572]_ );
  assign \new_[15598]_  = \new_[18256]_  ^ \new_[16202]_ ;
  assign \new_[15599]_  = (~\new_[18649]_  | ~\new_[16403]_ ) & (~\new_[16878]_  | ~\new_[15928]_ );
  assign n16255 = ~n16380 & ~n16500;
  assign \new_[15601]_  = ~\new_[15976]_  | ~\new_[17038]_ ;
  assign \new_[15602]_  = ~\new_[13689]_  & (~\new_[16890]_  | ~\new_[16157]_ );
  assign \new_[15603]_  = ~\new_[19940]_  & ~\new_[18523]_ ;
  assign \new_[15604]_  = ~\new_[19940]_  & ~\new_[16912]_ ;
  assign \new_[15605]_  = ~\new_[20192]_  & ~\new_[17254]_ ;
  assign \new_[15606]_  = ~\new_[17160]_  | ~\new_[17190]_  | ~\new_[16754]_  | ~\new_[16195]_ ;
  assign \new_[15607]_  = ~\new_[10870]_  & ~\new_[20192]_  & ~\new_[10448]_ ;
  assign \new_[15608]_  = \new_[14957]_  ^ \new_[16203]_ ;
  assign \new_[15609]_  = \wbm_adr_o[12]  ^ \new_[16200]_ ;
  assign \new_[15610]_  = \new_[6317]_  ^ \new_[16197]_ ;
  assign n15950 = \new_[15199]_  ? \new_[17707]_  : \new_[17122]_ ;
  assign \new_[15612]_  = \\configuration_sync_cache_lsize_to_wb_bits_reg[8] ;
  assign \new_[15613]_  = ~\new_[15814]_ ;
  assign \new_[15614]_  = ~\new_[15970]_  | ~\new_[6310]_ ;
  assign \new_[15615]_  = ~\new_[15977]_  | ~\new_[6311]_ ;
  assign \new_[15616]_  = ~\new_[15971]_  | ~\new_[6313]_ ;
  assign \new_[15617]_  = \new_[15976]_  & \new_[5048]_ ;
  assign \new_[15618]_  = ~\new_[15982]_  & ~\new_[15981]_ ;
  assign \new_[15619]_  = ~\new_[19012]_  | ~\new_[18023]_  | ~\new_[16227]_  | ~\new_[16224]_ ;
  assign \new_[15620]_  = ~\new_[15978]_  | ~\wbm_adr_o[20] ;
  assign \new_[15621]_  = ~\new_[17159]_  | ~\new_[17188]_  | ~\new_[16739]_  | ~\new_[16222]_ ;
  assign \new_[15622]_  = ~\new_[15972]_  & ~\new_[15973]_ ;
  assign \new_[15623]_  = ~\new_[15974]_  & ~\new_[15975]_ ;
  assign \new_[15624]_  = ~\new_[16578]_  | ~\new_[17180]_  | ~\new_[15995]_  | ~\new_[16674]_ ;
  assign \new_[15625]_  = (~\new_[16161]_  | ~\new_[10000]_ ) & (~\new_[16215]_  | ~\new_[10001]_ );
  assign \new_[15626]_  = (~\new_[16161]_  | ~\new_[9992]_ ) & (~\new_[16215]_  | ~\new_[9988]_ );
  assign \new_[15627]_  = (~\new_[16161]_  | ~\new_[9991]_ ) & (~\new_[16215]_  | ~\new_[9995]_ );
  assign \new_[15628]_  = \new_[6303]_  ^ \new_[16222]_ ;
  assign \new_[15629]_  = \wbm_adr_o[11]  ^ \new_[16217]_ ;
  assign \new_[15630]_  = \new_[5090]_  ^ \new_[16226]_ ;
  assign \new_[15631]_  = ~configuration_interrupt_out_reg;
  assign \new_[15632]_  = ~\new_[15993]_  | ~pci_gnt_i;
  assign \new_[15633]_  = ~\new_[15743]_  | ~\new_[16678]_ ;
  assign \new_[15634]_  = \new_[15994]_  & \new_[9903]_ ;
  assign n16095 = \new_[15994]_  & \new_[17310]_ ;
  assign n15875 = \new_[16129]_  & \new_[16620]_ ;
  assign \new_[15637]_  = ~\new_[4008]_  & (~n16520 | ~\new_[16142]_ );
  assign \new_[15638]_  = ~\new_[16183]_  | ~\new_[16220]_  | ~\new_[17177]_ ;
  assign n15805 = \new_[15165]_  ? \new_[16362]_  : \new_[15170]_ ;
  assign n16250 = \new_[15181]_  ? \new_[16362]_  : \new_[15361]_ ;
  assign n15910 = \new_[16729]_  ? \new_[16362]_  : \new_[15191]_ ;
  assign n15900 = \new_[15178]_  ? \new_[16362]_  : \new_[15189]_ ;
  assign n16105 = \new_[15200]_  ? \new_[16362]_  : \new_[15270]_ ;
  assign n16315 = \new_[18649]_  ? \new_[16362]_  : \new_[15402]_ ;
  assign n15960 = \new_[15179]_  ? \new_[16362]_  : \new_[15201]_ ;
  assign n15880 = \new_[15198]_  ? \new_[16362]_  : \new_[15185]_ ;
  assign n16075 = \new_[15176]_  ? \new_[16362]_  : \new_[15232]_ ;
  assign n16115 = \new_[19199]_  ? \new_[16362]_  : \new_[15284]_ ;
  assign n15885 = \new_[15169]_  ? \new_[16362]_  : \new_[15186]_ ;
  assign n15890 = \new_[15168]_  ? \new_[16362]_  : \new_[15187]_ ;
  assign n15895 = \new_[15167]_  ? \new_[16362]_  : \new_[15188]_ ;
  assign n15925 = \new_[18088]_  ? \new_[16362]_  : \new_[15194]_ ;
  assign n16300 = \new_[15182]_  ? \new_[16362]_  : \new_[15399]_ ;
  assign n15770 = \new_[15195]_  ? \new_[16362]_  : \new_[15163]_ ;
  assign n16140 = \new_[15196]_  ? \new_[16362]_  : \new_[15309]_ ;
  assign n15765 = \new_[15166]_  ? \new_[16362]_  : \new_[15161]_ ;
  assign n16130 = \new_[15180]_  ? \new_[16362]_  : \new_[15300]_ ;
  assign n15775 = \new_[15092]_  ? \new_[16362]_  : \new_[17746]_ ;
  assign n15995 = \new_[15197]_  ? \new_[16362]_  : \new_[15210]_ ;
  assign n16120 = \new_[18609]_  ? \new_[16362]_  : \new_[15285]_ ;
  assign n15970 = \new_[18888]_  ? \new_[16362]_  : \new_[15204]_ ;
  assign n16070 = \new_[19255]_  ? \new_[16362]_  : \new_[15231]_ ;
  assign n15820 = \new_[16838]_  ? \new_[16362]_  : \new_[18300]_ ;
  assign n16060 = \new_[17318]_  ? \new_[16362]_  : \new_[19074]_ ;
  assign n15905 = \new_[15230]_  ? \new_[16362]_  : \new_[15190]_ ;
  assign n16080 = \new_[18624]_  ? \new_[16362]_  : \new_[15233]_ ;
  assign n16295 = \new_[14208]_  ? \new_[16362]_  : \new_[17794]_ ;
  assign n16090 = \new_[17476]_  ? \new_[16362]_  : \new_[19634]_ ;
  assign n16110 = \new_[15174]_  ? \new_[16362]_  : \new_[15272]_ ;
  assign n15870 = \new_[18428]_  ? \new_[16362]_  : \new_[15183]_ ;
  assign n15915 = \new_[18642]_  ? \new_[16362]_  : \new_[15192]_ ;
  assign n16100 = \new_[15287]_  ? \new_[16362]_  : \new_[15268]_ ;
  assign n16305 = \new_[15222]_  ? \new_[16362]_  : \new_[15400]_ ;
  assign n16320 = \new_[15171]_  ? \new_[16362]_  : \new_[15406]_ ;
  assign n16085 = \new_[15160]_  ? \new_[16362]_  : \new_[15236]_ ;
  assign n16310 = \new_[15303]_  ? \new_[16362]_  : \new_[15401]_ ;
  assign n16265 = \new_[18289]_  ? \new_[16362]_  : \new_[15387]_ ;
  assign n16145 = \new_[15172]_  ? \new_[16362]_  : \new_[15329]_ ;
  assign \new_[15679]_  = \new_[18438]_  ^ \new_[16336]_ ;
  assign \new_[15680]_  = ~\new_[17667]_  | ~\new_[13821]_  | ~\new_[16031]_  | ~\new_[14861]_ ;
  assign \new_[15681]_  = ~\new_[17698]_  | ~\new_[18509]_  | ~\new_[16035]_  | ~\new_[18756]_ ;
  assign \new_[15682]_  = \new_[16729]_  ? \new_[16436]_  : \new_[20319]_ ;
  assign \new_[15683]_  = ~\new_[15802]_ ;
  assign \new_[15684]_  = ~\new_[12051]_  | ~\new_[20056]_ ;
  assign \new_[15685]_  = ~\new_[12073]_  | ~\new_[19957]_ ;
  assign \new_[15686]_  = ~\new_[12532]_  | ~\new_[19957]_ ;
  assign \new_[15687]_  = ~\new_[16077]_  | ~n16995;
  assign \new_[15688]_  = \new_[16577]_  | \new_[15411]_ ;
  assign \new_[15689]_  = ~\new_[10396]_  | ~\new_[16077]_ ;
  assign \new_[15690]_  = ~\new_[20049]_  | ~\new_[10481]_ ;
  assign \new_[15691]_  = ~\new_[16077]_  | ~n17500;
  assign \new_[15692]_  = \new_[16577]_  | \new_[18584]_ ;
  assign \new_[15693]_  = ~\new_[19029]_  | ~\new_[19948]_  | ~\new_[16436]_ ;
  assign \new_[15694]_  = ~\new_[16077]_  | ~n17220;
  assign \new_[15695]_  = ~\new_[10854]_  | ~\new_[20506]_ ;
  assign \new_[15696]_  = \new_[17032]_  & \new_[16073]_ ;
  assign n16260 = ~\new_[16062]_  | (~\new_[15385]_  & ~\new_[16572]_ );
  assign n16280 = ~\new_[16063]_  | (~\new_[15392]_  & ~\new_[16572]_ );
  assign \new_[15699]_  = \new_[16073]_  & \new_[16115]_ ;
  assign n16290 = ~\new_[15915]_  | (~\new_[15396]_  & ~\new_[16572]_ );
  assign n15920 = ~\new_[15917]_  | (~\new_[15193]_  & ~\new_[16572]_ );
  assign n16275 = ~\new_[16068]_  | (~\new_[15390]_  & ~\new_[16572]_ );
  assign n16285 = ~\new_[16068]_  | (~\new_[20352]_  & ~\new_[16572]_ );
  assign \new_[15704]_  = (~\new_[16403]_  | ~\new_[19255]_ ) & (~\new_[16878]_  | ~\new_[16354]_ );
  assign pci_req_o = pci_io_mux_req_iob_dat_out_reg;
  assign \new_[15706]_  = ~\new_[16185]_  | ~\new_[17182]_  | ~\new_[17108]_ ;
  assign n15760 = \new_[16405]_  ? \new_[19929]_  : \new_[15160]_ ;
  assign n16135 = \new_[16369]_  ? \new_[19929]_  : \new_[15303]_ ;
  assign n15855 = \new_[15989]_  ? \new_[19929]_  : \new_[15180]_ ;
  assign n15815 = \new_[15948]_  ? \new_[19929]_  : \new_[15172]_ ;
  assign n15785 = \new_[16382]_  ? \new_[19929]_  : \new_[15166]_ ;
  assign n16125 = \new_[16440]_  ? \new_[19929]_  : \new_[15287]_ ;
  assign n15825 = \new_[15925]_  ? \new_[19929]_  : \new_[15174]_ ;
  assign n15940 = \new_[16144]_  ? \new_[19929]_  : \new_[15197]_ ;
  assign n15845 = \new_[15927]_  ? \new_[19929]_  : \new_[15178]_ ;
  assign n15850 = \new_[16443]_  ? \new_[19929]_  : \new_[15179]_ ;
  assign n15945 = \new_[16143]_  ? \new_[19929]_  : \new_[15198]_ ;
  assign n15800 = \new_[16107]_  ? \new_[19929]_  : \new_[15169]_ ;
  assign n15930 = \new_[16210]_  ? \new_[19929]_  : \new_[15195]_ ;
  assign \new_[15720]_  = \new_[17405]_  ^ \new_[20143]_ ;
  assign n15860 = \new_[15181]_  ? \new_[16572]_  : \new_[17476]_ ;
  assign n15780 = \new_[15926]_  ? \new_[19929]_  : \new_[15165]_ ;
  assign n15935 = \new_[15985]_  ? \new_[19929]_  : \new_[15196]_ ;
  assign n15865 = \new_[15182]_  ? \new_[16572]_  : \new_[17318]_ ;
  assign n15955 = \new_[16127]_  ? \new_[19929]_  : \new_[15200]_ ;
  assign n15835 = \new_[16032]_  ? \new_[19929]_  : \new_[15176]_ ;
  assign n15795 = \new_[15941]_  ? \new_[19929]_  : \new_[15168]_ ;
  assign n16065 = \new_[16134]_  ? \new_[19929]_  : \new_[15230]_ ;
  assign n15810 = \new_[15924]_  ? \new_[19929]_  : \new_[15171]_ ;
  assign n16055 = \new_[16100]_  ? \new_[19929]_  : \new_[15222]_ ;
  assign n15840 = \new_[17318]_  ? n16645 : \new_[17380]_ ;
  assign n15830 = \new_[17476]_  ? \new_[17707]_  : \new_[17405]_ ;
  assign n16025 = \new_[16838]_  ? \new_[17707]_  : \new_[17404]_ ;
  assign \new_[15734]_  = \new_[20125]_  & \new_[17033]_ ;
  assign \new_[15735]_  = \new_[16099]_  & \new_[16617]_ ;
  assign \new_[15736]_  = ~\new_[16658]_  | ~\new_[13813]_  | ~\new_[16153]_ ;
  assign \new_[15737]_  = \new_[12301]_  ^ \new_[16445]_ ;
  assign \new_[15738]_  = \new_[16098]_  & \new_[17473]_ ;
  assign \new_[15739]_  = wbs_cyc_i & \new_[16098]_ ;
  assign \new_[15740]_  = ~\new_[16990]_  | ~\new_[20212]_ ;
  assign \new_[15741]_  = ~\new_[16164]_  & ~\new_[15920]_ ;
  assign \new_[15742]_  = \new_[16402]_  & \new_[20451]_ ;
  assign \new_[15743]_  = ~\new_[16446]_ ;
  assign \new_[15744]_  = ~\new_[16101]_  & ~\new_[19912]_ ;
  assign \new_[15745]_  = \new_[16619]_  | \new_[16101]_ ;
  assign \new_[15746]_  = ~\new_[16619]_  & ~\new_[16104]_ ;
  assign \new_[15747]_  = ~\new_[15889]_ ;
  assign n16150 = ~n16380 & (~\new_[17249]_  | ~\new_[19930]_ );
  assign \new_[15749]_  = \new_[20451]_  & \new_[20161]_ ;
  assign n16050 = \new_[15196]_  ? \new_[16415]_  : \new_[15985]_ ;
  assign n16205 = \new_[18289]_  ? \new_[16415]_  : \new_[16414]_ ;
  assign n15990 = \new_[15179]_  ? \new_[16415]_  : \new_[16443]_ ;
  assign n16210 = \new_[18088]_  ? \new_[16415]_  : \new_[15923]_ ;
  assign n15985 = \new_[15230]_  ? \new_[16415]_  : \new_[16134]_ ;
  assign n16180 = \new_[15167]_  ? \new_[16415]_  : \new_[16130]_ ;
  assign n16170 = \new_[15165]_  ? \new_[16415]_  : \new_[15926]_ ;
  assign n16245 = \new_[15171]_  ? \new_[16415]_  : \new_[15924]_ ;
  assign n15965 = \new_[15180]_  ? \new_[16415]_  : \new_[15989]_ ;
  assign n16035 = \new_[15198]_  ? \new_[16415]_  : \new_[16143]_ ;
  assign n15975 = \new_[15195]_  ? \new_[16415]_  : \new_[16210]_ ;
  assign n16045 = \new_[15303]_  ? \new_[16415]_  : \new_[16369]_ ;
  assign n16175 = \new_[15287]_  ? \new_[16415]_  : \new_[16440]_ ;
  assign n16005 = \new_[18642]_  ? \new_[16415]_  : \new_[16013]_ ;
  assign n16195 = \new_[15182]_  ? \new_[16415]_  : \new_[17318]_ ;
  assign n16240 = \new_[15169]_  ? \new_[16415]_  : \new_[16107]_ ;
  assign n15980 = \new_[15181]_  ? \new_[16415]_  : \new_[17476]_ ;
  assign n16160 = \new_[15172]_  ? \new_[16415]_  : \new_[15948]_ ;
  assign n16185 = \new_[15178]_  ? \new_[16415]_  : \new_[15927]_ ;
  assign n16165 = \new_[15160]_  ? \new_[16415]_  : \new_[16405]_ ;
  assign n16190 = \new_[18428]_  ? \new_[16415]_  : \new_[16384]_ ;
  assign n16040 = \new_[15166]_  ? \new_[16415]_  : \new_[16382]_ ;
  assign n16010 = \new_[18624]_  ? \new_[16415]_  : \new_[16150]_ ;
  assign n16030 = \new_[15174]_  ? \new_[16415]_  : \new_[15925]_ ;
  assign n16000 = \new_[19199]_  ? \new_[16415]_  : \new_[16435]_ ;
  assign n16020 = \new_[15222]_  ? \new_[16415]_  : \new_[16100]_ ;
  assign n16215 = \new_[18888]_  ? \new_[16415]_  : \new_[16027]_ ;
  assign n16225 = \new_[15168]_  ? \new_[16415]_  : \new_[15941]_ ;
  assign n16015 = \new_[15092]_  ? \new_[16415]_  : \new_[16838]_ ;
  assign n16200 = \new_[18609]_  ? \new_[16415]_  : \new_[15986]_ ;
  assign n16235 = \new_[15200]_  ? \new_[16415]_  : \new_[16127]_ ;
  assign n16220 = \new_[15197]_  ? \new_[16415]_  : \new_[16144]_ ;
  assign n16230 = \new_[15176]_  ? \new_[16415]_  : \new_[16032]_ ;
  assign \new_[15783]_  = \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[3] ;
  assign \new_[15784]_  = ~\new_[16108]_  | ~\new_[19928]_ ;
  assign \new_[15785]_  = ~\new_[17134]_  | ~\new_[16132]_ ;
  assign \new_[15786]_  = ~\new_[16165]_  | ~\new_[16219]_  | ~\new_[17184]_ ;
  assign \new_[15787]_  = ~\new_[14957]_  | ~\new_[13704]_  | ~\new_[15922]_  | ~\new_[17741]_ ;
  assign \new_[15788]_  = ~\new_[18256]_  | ~\new_[18595]_  | ~\new_[15943]_  | ~\new_[17259]_ ;
  assign \new_[15789]_  = \new_[6323]_  ^ \new_[16181]_ ;
  assign \new_[15790]_  = \wbm_adr_o[6]  ^ \new_[16182]_ ;
  assign \new_[15791]_  = ~\new_[17385]_  & ~\new_[20128]_ ;
  assign \new_[15792]_  = ~\new_[15908]_ ;
  assign n15790 = \new_[16130]_  ? \new_[19929]_  : \new_[15167]_ ;
  assign \new_[15794]_  = \new_[14911]_  ^ \new_[16329]_ ;
  assign \new_[15795]_  = \new_[15829]_ ;
  assign \new_[15796]_  = ~\new_[13821]_  | ~\new_[17465]_  | ~\new_[15953]_  | ~\new_[14861]_ ;
  assign \new_[15797]_  = ~\new_[15937]_  | ~\new_[17276]_ ;
  assign \new_[15798]_  = ~\new_[18509]_  | ~\new_[17270]_  | ~\new_[15954]_  | ~\new_[18756]_ ;
  assign n16340 = \new_[15424]_  ? \new_[17707]_  : \new_[16889]_ ;
  assign \new_[15800]_  = ~\new_[16368]_  & ~\new_[16820]_ ;
  assign \new_[15801]_  = ~\new_[15934]_ ;
  assign \new_[15802]_  = ~pci_target_unit_pci_target_sm_state_transfere_reg_reg;
  assign \new_[15803]_  = \new_[17166]_  & \new_[16183]_ ;
  assign \new_[15804]_  = \new_[17182]_  & \new_[16185]_ ;
  assign \new_[15805]_  = \new_[16220]_  & \new_[16183]_ ;
  assign \new_[15806]_  = ~\new_[15937]_ ;
  assign \new_[15807]_  = ~\new_[16979]_  | ~\new_[16184]_  | ~\new_[16503]_ ;
  assign \new_[15808]_  = \new_[16223]_  & \new_[16185]_ ;
  assign \new_[15809]_  = \new_[14969]_  ? \new_[16613]_  : \new_[18268]_ ;
  assign \new_[15810]_  = ~\new_[16103]_ ;
  assign \new_[15811]_  = ~\new_[16176]_  | (~\new_[16682]_  & ~\new_[9647]_ );
  assign \new_[15812]_  = ~\new_[19909]_  & (~\new_[16606]_  | ~\new_[16781]_ );
  assign n16355 = \new_[17374]_  & \new_[16361]_ ;
  assign \new_[15814]_  = ~\new_[16474]_  & ~\new_[16201]_ ;
  assign \new_[15815]_  = \new_[16200]_  & \new_[17178]_ ;
  assign \new_[15816]_  = ~\new_[16479]_  & ~\new_[16199]_ ;
  assign \new_[15817]_  = \new_[16197]_  & \new_[17189]_ ;
  assign \new_[15818]_  = ~\new_[16195]_  | ~\new_[17190]_ ;
  assign \new_[15819]_  = ~\new_[17178]_  | ~\new_[16200]_  | ~\new_[17135]_ ;
  assign \new_[15820]_  = ~\new_[17189]_  | ~\new_[16197]_  | ~\new_[17172]_ ;
  assign \new_[15821]_  = (~\new_[17059]_  | ~\new_[16511]_ ) & (~\new_[16863]_  | ~\new_[5096]_ );
  assign \new_[15822]_  = ~\new_[17187]_  | ~\new_[16704]_  | ~\new_[16731]_  | ~\new_[17160]_ ;
  assign \new_[15823]_  = ~\new_[17138]_  | ~\new_[16703]_  | ~\new_[16809]_  | ~\new_[17172]_ ;
  assign \new_[15824]_  = ~\new_[17164]_  | ~\new_[16705]_  | ~\new_[16835]_  | ~\new_[17135]_ ;
  assign \new_[15825]_  = ~\new_[15943]_ ;
  assign \new_[15826]_  = \new_[14989]_  ^ \new_[16508]_ ;
  assign \new_[15827]_  = \new_[18247]_  ^ \new_[16509]_ ;
  assign \new_[15828]_  = ~\new_[15922]_ ;
  assign \new_[15829]_  = \new_[16212]_  & \new_[9800]_ ;
  assign \new_[15830]_  = \new_[17196]_  & \new_[16226]_ ;
  assign \new_[15831]_  = \new_[16217]_  & \new_[17179]_ ;
  assign \new_[15832]_  = ~\new_[16148]_  | (~\new_[17086]_  & ~\new_[17793]_ );
  assign \new_[15833]_  = \new_[16211]_  | \new_[16684]_ ;
  assign \new_[15834]_  = \new_[16222]_  & \new_[17083]_ ;
  assign \new_[15835]_  = ~\new_[16204]_  & ~\new_[16743]_ ;
  assign \new_[15836]_  = ~\new_[16230]_  | ~n16575;
  assign \new_[15837]_  = ~\new_[15976]_ ;
  assign \new_[15838]_  = ~\wbm_adr_o[2]  | ~\new_[16218]_  | ~\new_[17162]_ ;
  assign n16345 = ~\new_[16618]_  | (~\new_[20081]_  & ~\new_[17971]_ );
  assign \new_[15840]_  = ~\new_[16213]_  & (~\new_[17254]_  | ~n16690);
  assign \new_[15841]_  = ~\new_[16353]_  & ~\new_[16355]_ ;
  assign \new_[15842]_  = ~\new_[16148]_  | (~\new_[12448]_  & ~\new_[17793]_ );
  assign \new_[15843]_  = ~\new_[16148]_  | (~\new_[18445]_  & ~\new_[17323]_ );
  assign \new_[15844]_  = ~\new_[16738]_  | ~\new_[16818]_  | ~\new_[16742]_  | ~\new_[16741]_ ;
  assign \new_[15845]_  = ~\new_[16746]_  | ~\new_[16834]_  | ~\new_[16773]_  | ~\new_[16750]_ ;
  assign \new_[15846]_  = ~\new_[16757]_  | ~\new_[16769]_  | ~\new_[16767]_  | ~\new_[16831]_ ;
  assign \new_[15847]_  = ~\new_[16830]_  | ~\new_[16765]_  | ~\new_[16768]_  | ~\new_[16766]_ ;
  assign \new_[15848]_  = ~\new_[16686]_  | ~\new_[16761]_  | ~\new_[16759]_  | ~\new_[16749]_ ;
  assign \new_[15849]_  = \new_[16212]_  & \new_[16216]_ ;
  assign \new_[15850]_  = ~\new_[17104]_  | ~\new_[16647]_  | ~\new_[17089]_  | ~\new_[16644]_ ;
  assign \new_[15851]_  = ~\new_[16192]_  | (~\new_[16770]_  & ~\new_[9619]_ );
  assign \new_[15852]_  = \new_[4976]_  ^ \new_[16576]_ ;
  assign \new_[15853]_  = \new_[16674]_  & \new_[16578]_ ;
  assign \new_[15854]_  = ~\new_[16367]_  & ~\new_[19901]_ ;
  assign \new_[15855]_  = ~\new_[10001]_  | ~\new_[16402]_  | ~\new_[19886]_ ;
  assign \new_[15856]_  = ~\new_[9904]_  | ~\new_[16402]_  | ~\new_[20377]_ ;
  assign \new_[15857]_  = ~\new_[15995]_ ;
  assign n16350 = ~\new_[16954]_  & ~\new_[16142]_ ;
  assign \new_[15859]_  = ~\new_[10528]_  | ~\new_[16179]_  | ~\new_[16411]_  | ~\new_[9997]_ ;
  assign \new_[15860]_  = \new_[14969]_  ? \new_[16615]_  : \new_[19506]_ ;
  assign \new_[15861]_  = ~\new_[13601]_  | ~\new_[13689]_  | ~\new_[16376]_  | ~\new_[15594]_ ;
  assign \new_[15862]_  = \new_[17403]_  ^ \new_[20340]_ ;
  assign \new_[15863]_  = \new_[8390]_  ^ \new_[16600]_ ;
  assign n16330 = \new_[15417]_  ? n16645 : \new_[16620]_ ;
  assign n16325 = n16500 ? n16645 : \new_[20082]_ ;
  assign \new_[15866]_  = ~\new_[12302]_  | ~\new_[19929]_ ;
  assign \new_[15867]_  = ~\new_[17122]_  & ~\new_[16782]_ ;
  assign \new_[15868]_  = ~\new_[13869]_  | ~\new_[19929]_ ;
  assign \new_[15869]_  = ~\new_[9877]_  | ~\new_[19929]_ ;
  assign \new_[15870]_  = ~\new_[17802]_  | ~\new_[19929]_ ;
  assign \new_[15871]_  = ~\new_[20128]_  | ~\new_[19929]_ ;
  assign \new_[15872]_  = ~\new_[20159]_  | ~\new_[19929]_ ;
  assign \new_[15873]_  = ~\new_[20488]_  | ~\new_[19929]_ ;
  assign \new_[15874]_  = ~\new_[14208]_  | ~\new_[19929]_ ;
  assign \new_[15875]_  = ~\new_[12039]_  | ~\new_[19929]_ ;
  assign \new_[15876]_  = \new_[19886]_  & \new_[9880]_ ;
  assign \new_[15877]_  = ~\new_[17636]_  | ~\new_[19929]_ ;
  assign \new_[15878]_  = ~\new_[16398]_  & ~\new_[17062]_ ;
  assign \new_[15879]_  = ~n16690 & ~\new_[19929]_ ;
  assign \new_[15880]_  = ~\new_[19929]_  | ~\new_[13678]_ ;
  assign \new_[15881]_  = ~\new_[9884]_  | ~\new_[19929]_ ;
  assign \new_[15882]_  = ~\new_[9765]_  | ~\new_[19929]_ ;
  assign \new_[15883]_  = ~\new_[17474]_  | ~\new_[19929]_ ;
  assign \new_[15884]_  = \new_[16833]_  & \new_[20125]_ ;
  assign \new_[15885]_  = ~\new_[16158]_  & ~\new_[16409]_ ;
  assign \new_[15886]_  = \new_[16171]_  | \new_[17310]_ ;
  assign \new_[15887]_  = ~\new_[16400]_  & ~\new_[11328]_ ;
  assign \new_[15888]_  = \new_[20377]_  & \new_[16401]_ ;
  assign \new_[15889]_  = \new_[16404]_  & \new_[20178]_ ;
  assign \new_[15890]_  = \new_[16402]_  & \new_[20377]_ ;
  assign \new_[15891]_  = ~\new_[16399]_  | ~n16575;
  assign \new_[15892]_  = ~\new_[16101]_ ;
  assign \new_[15893]_  = ~\new_[16430]_  & ~\new_[20128]_ ;
  assign \new_[15894]_  = ~\new_[16105]_ ;
  assign \new_[15895]_  = \new_[14990]_  ^ \new_[16461]_ ;
  assign \new_[15896]_  = \new_[9808]_  ^ \new_[16460]_ ;
  assign \new_[15897]_  = ~\new_[20205]_  | ~\new_[20212]_ ;
  assign \new_[15898]_  = ~\new_[20340]_  | ~\new_[15923]_ ;
  assign \new_[15899]_  = ~\new_[15931]_ ;
  assign \new_[15900]_  = ~\new_[20340]_  | ~\new_[15986]_ ;
  assign \new_[15901]_  = ~\new_[16122]_ ;
  assign \new_[15902]_  = ~\new_[20340]_  | ~\new_[16414]_ ;
  assign \new_[15903]_  = ~\new_[16837]_  & ~\new_[16836]_ ;
  assign \new_[15904]_  = ~\new_[9884]_  & ~\new_[16852]_ ;
  assign \new_[15905]_  = ~\new_[20340]_  | ~\new_[16013]_ ;
  assign \new_[15906]_  = ~\new_[16436]_  & ~\new_[12039]_ ;
  assign \new_[15907]_  = ~\new_[16852]_  & ~\new_[19029]_ ;
  assign \new_[15908]_  = ~\new_[9884]_  & ~\new_[16436]_ ;
  assign \new_[15909]_  = \new_[17116]_  & \new_[16181]_ ;
  assign \new_[15910]_  = \new_[17165]_  & \new_[16182]_ ;
  assign \new_[15911]_  = \new_[14988]_  ^ \new_[16462]_ ;
  assign \new_[15912]_  = ~\new_[17122]_  & ~\new_[19742]_ ;
  assign \new_[15913]_  = \new_[9798]_  ^ \new_[16463]_ ;
  assign \new_[15914]_  = ~\new_[16572]_  | ~\new_[16013]_ ;
  assign \new_[15915]_  = ~\new_[16572]_  | ~\new_[15923]_ ;
  assign \new_[15916]_  = \new_[19774]_  ? \new_[16785]_  : \new_[17694]_ ;
  assign \new_[15917]_  = ~\new_[16572]_  | ~\new_[16414]_ ;
  assign \new_[15918]_  = ~\new_[16616]_  | ~\new_[10855]_ ;
  assign \new_[15919]_  = pci_target_unit_pci_target_sm_previous_frame_reg;
  assign \new_[15920]_  = \new_[17794]_  ^ \new_[17258]_ ;
  assign \new_[15921]_  = \new_[16589]_  | pci_gnt_i;
  assign \new_[15922]_  = ~\new_[16730]_  & ~\new_[16462]_ ;
  assign \new_[15923]_  = \\input_register_pci_ad_reg_out_reg[7] ;
  assign \new_[15924]_  = \\input_register_pci_ad_reg_out_reg[17] ;
  assign \new_[15925]_  = \\input_register_pci_ad_reg_out_reg[30] ;
  assign \new_[15926]_  = \\input_register_pci_ad_reg_out_reg[16] ;
  assign \new_[15927]_  = \\input_register_pci_ad_reg_out_reg[28] ;
  assign \new_[15928]_  = \\input_register_pci_ad_reg_out_reg[0] ;
  assign \new_[15929]_  = \new_[17561]_  ? \new_[16787]_  : \new_[19865]_ ;
  assign \new_[15930]_  = \new_[9618]_  ^ \new_[16657]_ ;
  assign \new_[15931]_  = \new_[20340]_  & \new_[15928]_ ;
  assign \new_[15932]_  = \new_[9623]_  ^ \new_[16816]_ ;
  assign \new_[15933]_  = ~\new_[16416]_ ;
  assign \new_[15934]_  = ~\new_[20340]_  | ~\new_[16354]_ ;
  assign \new_[15935]_  = ~\new_[16889]_  & ~\new_[20082]_ ;
  assign n16370 = \\configuration_int_pin_sync_sync_data_out_reg[0] ;
  assign \new_[15937]_  = ~\new_[17000]_  & ~\new_[16476]_ ;
  assign \new_[15938]_  = ~n16380 & ~n16775;
  assign \new_[15939]_  = ~\new_[16499]_  | ~\new_[17370]_ ;
  assign \new_[15940]_  = ~\new_[17851]_  | ~\new_[12039]_  | ~\new_[16904]_  | ~\new_[17467]_ ;
  assign \new_[15941]_  = \\input_register_pci_ad_reg_out_reg[24] ;
  assign \new_[15942]_  = ~\new_[19886]_ ;
  assign \new_[15943]_  = ~\new_[16727]_  & ~\new_[16463]_ ;
  assign \new_[15944]_  = \new_[9626]_  ^ \new_[16700]_ ;
  assign \new_[15945]_  = \new_[6322]_  ^ \new_[16699]_ ;
  assign \new_[15946]_  = \new_[4962]_  ^ \new_[16661]_ ;
  assign \new_[15947]_  = \wbm_adr_o[5]  ^ \new_[16701]_ ;
  assign \new_[15948]_  = \\input_register_pci_ad_reg_out_reg[10] ;
  assign \new_[15949]_  = \new_[19023]_  ^ \new_[16846]_ ;
  assign \new_[15950]_  = ~\new_[16477]_  | ~n16910;
  assign \new_[15951]_  = ~\new_[5008]_  | ~\new_[16755]_  | ~\new_[16644]_ ;
  assign \new_[15952]_  = (~\new_[16863]_  & ~\new_[18152]_  & ~\new_[11133]_ ) | (~\new_[17442]_  & ~\new_[16863]_  & ~\new_[18152]_ );
  assign \new_[15953]_  = ~\new_[16642]_  & ~\new_[16897]_ ;
  assign \new_[15954]_  = ~\new_[16641]_  & ~\new_[16898]_ ;
  assign \new_[15955]_  = \new_[11330]_  ^ \new_[16702]_ ;
  assign \new_[15956]_  = \new_[5042]_  ^ \new_[16704]_ ;
  assign \new_[15957]_  = \wbm_adr_o[8]  ^ \new_[16705]_ ;
  assign \new_[15958]_  = \new_[6551]_  ^ \new_[16703]_ ;
  assign \new_[15959]_  = \new_[16720]_  ^ \new_[16721]_ ;
  assign \new_[15960]_  = \new_[16723]_  ^ \new_[16712]_ ;
  assign \new_[15961]_  = \new_[16713]_  ^ \new_[16719]_ ;
  assign \new_[15962]_  = \new_[16716]_  ^ \new_[16718]_ ;
  assign \new_[15963]_  = \new_[16669]_  ^ \new_[16711]_ ;
  assign \new_[15964]_  = \new_[16714]_  ^ \new_[16715]_ ;
  assign \new_[15965]_  = \new_[16722]_  ^ \new_[16680]_ ;
  assign n16365 = \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[6] ;
  assign \new_[15967]_  = \new_[16514]_  | \new_[17169]_ ;
  assign \new_[15968]_  = \new_[16513]_  | \new_[16789]_ ;
  assign n16375 = ~\new_[16196]_ ;
  assign \new_[15970]_  = ~\new_[6554]_  | ~\new_[16752]_  | ~\new_[16646]_ ;
  assign \new_[15971]_  = ~\new_[16726]_  | ~\new_[16646]_  | ~\new_[16645]_ ;
  assign \new_[15972]_  = ~\new_[16928]_  | ~\new_[16937]_  | ~\new_[16927]_  | ~\new_[16946]_ ;
  assign \new_[15973]_  = ~\new_[16943]_  | ~\new_[16929]_  | ~\new_[16945]_  | ~\new_[16947]_ ;
  assign \new_[15974]_  = ~\new_[16942]_  | ~\new_[16934]_  | ~\new_[16926]_  | ~\new_[16941]_ ;
  assign \new_[15975]_  = ~\new_[16930]_  | ~\new_[16931]_  | ~\new_[16939]_  | ~\new_[16938]_ ;
  assign \new_[15976]_  = ~\new_[16545]_  & (~\new_[17293]_  | ~\new_[17453]_ );
  assign \new_[15977]_  = ~\new_[17138]_  | ~\new_[17285]_  | ~\new_[17192]_  | ~\new_[16809]_ ;
  assign \new_[15978]_  = ~\new_[17164]_  | ~\new_[17283]_  | ~\new_[17074]_  | ~\new_[16835]_ ;
  assign \new_[15979]_  = ~\new_[16451]_  & (~n17220 | ~\new_[17793]_ );
  assign \new_[15980]_  = ~\new_[16895]_  | ~\new_[16869]_  | ~\new_[17035]_  | ~\new_[16914]_ ;
  assign \new_[15981]_  = ~\new_[17016]_  | ~\new_[16916]_  | ~\new_[16870]_  | ~\new_[16865]_ ;
  assign \new_[15982]_  = ~\new_[16924]_  | ~\new_[17023]_  | ~\new_[16917]_  | ~\new_[16919]_ ;
  assign \new_[15983]_  = ~\new_[17187]_  | ~\new_[17438]_  | ~\new_[17197]_  | ~\new_[16731]_ ;
  assign \new_[15984]_  = \new_[17015]_  ^ \new_[16811]_ ;
  assign \new_[15985]_  = \\input_register_pci_ad_reg_out_reg[12] ;
  assign \new_[15986]_  = \\input_register_pci_ad_reg_out_reg[3] ;
  assign \new_[15987]_  = \new_[6324]_  ^ \new_[16726]_ ;
  assign \new_[15988]_  = \wbm_adr_o[7]  ^ \new_[16648]_ ;
  assign \new_[15989]_  = \\input_register_pci_ad_reg_out_reg[13] ;
  assign \new_[15990]_  = (~\new_[16810]_  | ~wbm_rty_i) & (~\new_[9621]_  | ~\new_[18523]_ );
  assign \new_[15991]_  = ~parity_checker_master_perr_report_reg;
  assign \new_[15992]_  = ~\new_[15015]_  & ~\new_[16734]_ ;
  assign \new_[15993]_  = ~\new_[16221]_ ;
  assign \new_[15994]_  = \new_[20090]_ ;
  assign \new_[15995]_  = ~\new_[17180]_  | ~\new_[16912]_  | ~\new_[16674]_ ;
  assign \new_[15996]_  = \new_[17712]_  ? \new_[16787]_  : \new_[18774]_ ;
  assign \new_[15997]_  = \new_[17608]_  ? \new_[16787]_  : \new_[18542]_ ;
  assign \new_[15998]_  = \new_[17639]_  ? \new_[16787]_  : \new_[18900]_ ;
  assign \new_[15999]_  = \new_[17694]_  ? \new_[16787]_  : \new_[19595]_ ;
  assign \new_[16000]_  = \new_[17700]_  ? \new_[16787]_  : \new_[19183]_ ;
  assign \new_[16001]_  = \new_[17734]_  ? \new_[16787]_  : \new_[18940]_ ;
  assign \new_[16002]_  = \new_[17758]_  ? \new_[16787]_  : \new_[18194]_ ;
  assign \new_[16003]_  = \new_[17728]_  ? \new_[16787]_  : \new_[18874]_ ;
  assign \new_[16004]_  = \new_[17719]_  ? \new_[16787]_  : \new_[19121]_ ;
  assign \new_[16005]_  = \new_[17641]_  ? \new_[16787]_  : \new_[18069]_ ;
  assign \new_[16006]_  = \new_[17613]_  ? \new_[16787]_  : \new_[18312]_ ;
  assign \new_[16007]_  = \new_[17642]_  ? \new_[16787]_  : \new_[19487]_ ;
  assign \new_[16008]_  = \new_[17760]_  ? \new_[16787]_  : \new_[17839]_ ;
  assign \new_[16009]_  = \new_[17755]_  ? \new_[16787]_  : \new_[18539]_ ;
  assign \new_[16010]_  = \new_[17688]_  ? \new_[16787]_  : \new_[19399]_ ;
  assign \new_[16011]_  = \new_[17723]_  ? \new_[16787]_  : \new_[19678]_ ;
  assign \new_[16012]_  = \new_[17645]_  ? \new_[16787]_  : \new_[18935]_ ;
  assign \new_[16013]_  = \\input_register_pci_ad_reg_out_reg[4] ;
  assign \new_[16014]_  = \new_[17591]_  ? \new_[16787]_  : \new_[18920]_ ;
  assign \new_[16015]_  = \new_[17703]_  ? \new_[16787]_  : \new_[18476]_ ;
  assign \new_[16016]_  = \new_[17702]_  ? \new_[16787]_  : \new_[18547]_ ;
  assign \new_[16017]_  = \new_[17633]_  ? \new_[16787]_  : \new_[18197]_ ;
  assign \new_[16018]_  = \new_[17564]_  ? \new_[16787]_  : \new_[18788]_ ;
  assign \new_[16019]_  = \new_[17560]_  ? \new_[16787]_  : \new_[18617]_ ;
  assign \new_[16020]_  = \new_[17650]_  ? \new_[16787]_  : \new_[18522]_ ;
  assign \new_[16021]_  = \new_[17708]_  ? \new_[16787]_  : \new_[19258]_ ;
  assign \new_[16022]_  = \new_[17612]_  ? \new_[16787]_  : \new_[18941]_ ;
  assign \new_[16023]_  = \new_[17599]_  ? \new_[16787]_  : \new_[17919]_ ;
  assign \new_[16024]_  = \new_[19297]_  ? \new_[16785]_  : \new_[17700]_ ;
  assign \new_[16025]_  = \new_[19780]_  ? \new_[16785]_  : \new_[17692]_ ;
  assign \new_[16026]_  = \new_[19776]_  ? \new_[16785]_  : \new_[17564]_ ;
  assign \new_[16027]_  = \\input_register_pci_ad_reg_out_reg[9] ;
  assign \new_[16028]_  = \new_[18588]_  ? \new_[16785]_  : \new_[17723]_ ;
  assign \new_[16029]_  = \new_[18036]_  ? \new_[16785]_  : \new_[17645]_ ;
  assign \new_[16030]_  = \new_[18629]_  ? \new_[16792]_  : \new_[14969]_ ;
  assign \new_[16031]_  = ~\new_[16329]_ ;
  assign \new_[16032]_  = \\input_register_pci_ad_reg_out_reg[14] ;
  assign \new_[16033]_  = \new_[19772]_  ? \new_[16785]_  : \new_[17758]_ ;
  assign \new_[16034]_  = \new_[19771]_  ? \new_[16785]_  : \new_[17627]_ ;
  assign \new_[16035]_  = ~\new_[16336]_ ;
  assign \new_[16036]_  = \new_[18253]_  ? \new_[16785]_  : \new_[17591]_ ;
  assign \new_[16037]_  = \new_[19438]_  ? \new_[16785]_  : \new_[17728]_ ;
  assign \new_[16038]_  = \new_[17380]_  ^ \new_[17080]_ ;
  assign \new_[16039]_  = \new_[18380]_  ? \new_[16785]_  : \new_[17703]_ ;
  assign \new_[16040]_  = \new_[19685]_  ? \new_[16785]_  : \new_[17760]_ ;
  assign \new_[16041]_  = \new_[18938]_  ? \new_[16785]_  : \new_[17608]_ ;
  assign \new_[16042]_  = \new_[18350]_  ? \new_[16785]_  : \new_[17755]_ ;
  assign \new_[16043]_  = \new_[19779]_  ? \new_[16785]_  : \new_[17561]_ ;
  assign \new_[16044]_  = \new_[19768]_  ? \new_[16785]_  : \new_[17560]_ ;
  assign \new_[16045]_  = \new_[18579]_  ? \new_[16785]_  : \new_[17712]_ ;
  assign \new_[16046]_  = \new_[18619]_  ? \new_[16785]_  : \new_[17639]_ ;
  assign \new_[16047]_  = \new_[19302]_  ? \new_[16785]_  : \new_[17641]_ ;
  assign \new_[16048]_  = \new_[19710]_  ? \new_[16785]_  : \new_[17734]_ ;
  assign \new_[16049]_  = \new_[18263]_  ? \new_[16785]_  : \new_[17612]_ ;
  assign \new_[16050]_  = \new_[19400]_  ? \new_[16785]_  : \new_[17650]_ ;
  assign \new_[16051]_  = \new_[18422]_  ? \new_[16785]_  : \new_[17688]_ ;
  assign \new_[16052]_  = \new_[19008]_  ? \new_[16785]_  : \new_[17753]_ ;
  assign \new_[16053]_  = \new_[19773]_  ? \new_[16785]_  : \new_[17759]_ ;
  assign \new_[16054]_  = \new_[18356]_  ? \new_[16785]_  : \new_[17613]_ ;
  assign \new_[16055]_  = \new_[19732]_  ? \new_[16785]_  : \new_[17719]_ ;
  assign \new_[16056]_  = \new_[18367]_  ? \new_[16785]_  : \new_[17599]_ ;
  assign \new_[16057]_  = \new_[19347]_  ? \new_[16785]_  : \new_[17708]_ ;
  assign \new_[16058]_  = \new_[18370]_  ? \new_[16785]_  : \new_[17633]_ ;
  assign \new_[16059]_  = \new_[19435]_  ? \new_[16785]_  : \new_[17702]_ ;
  assign n16360 = \new_[15594]_  ? n16645 : \new_[16668]_ ;
  assign \new_[16061]_  = ~pci_target_unit_del_sync_comp_done_reg_clr_reg;
  assign \new_[16062]_  = ~\new_[16572]_  | ~\new_[16027]_ ;
  assign \new_[16063]_  = ~\new_[16572]_  | ~\new_[16435]_ ;
  assign \new_[16064]_  = ~\new_[16572]_  | ~\new_[15986]_ ;
  assign \new_[16065]_  = ~\new_[16572]_  | ~\new_[16384]_ ;
  assign \new_[16066]_  = ~\new_[16572]_  | ~\new_[16150]_ ;
  assign \new_[16067]_  = ~\new_[16572]_  | ~\new_[16354]_ ;
  assign \new_[16068]_  = ~\new_[16572]_  | ~\new_[15928]_ ;
  assign \new_[16069]_  = \new_[16607]_  | \new_[19912]_ ;
  assign \new_[16070]_  = ~\new_[17908]_  | ~\new_[16615]_ ;
  assign \new_[16071]_  = ~\new_[20082]_  & ~n16775;
  assign \new_[16072]_  = ~\new_[16621]_  & ~\new_[17317]_ ;
  assign \new_[16073]_  = \new_[16827]_  & \new_[16608]_ ;
  assign \new_[16074]_  = ~\new_[19909]_  & ~\new_[16609]_ ;
  assign \new_[16075]_  = ~\new_[17951]_  | ~\new_[16613]_ ;
  assign \new_[16076]_  = \new_[16607]_  | \new_[16793]_ ;
  assign \new_[16077]_  = ~\new_[16605]_  & ~\new_[16793]_ ;
  assign \new_[16078]_  = \new_[16638]_  & \new_[16608]_ ;
  assign \new_[16079]_  = ~\new_[16194]_ ;
  assign \new_[16080]_  = (~\new_[16826]_  | ~\new_[5042]_ ) & (~\new_[17454]_  | ~\new_[10352]_ );
  assign \new_[16081]_  = (~\new_[17038]_  | ~\new_[4962]_ ) & (~\new_[17454]_  | ~\new_[10350]_ );
  assign \new_[16082]_  = (~\new_[17038]_  | ~\new_[5008]_ ) & (~\new_[17454]_  | ~\new_[10431]_ );
  assign \new_[16083]_  = (~\new_[17038]_  | ~\new_[5043]_ ) & (~\new_[17454]_  | ~\new_[10417]_ );
  assign \new_[16084]_  = (~\new_[17038]_  | ~\new_[5012]_ ) & (~\new_[17454]_  | ~\new_[10422]_ );
  assign \new_[16085]_  = (~\new_[16826]_  | ~\new_[4967]_ ) & (~\new_[17454]_  | ~\new_[10425]_ );
  assign \new_[16086]_  = (~\new_[17038]_  | ~\new_[4964]_ ) & (~\new_[17454]_  | ~\new_[10363]_ );
  assign \new_[16087]_  = (~\new_[17038]_  | ~\new_[4966]_ ) & (~\new_[17454]_  | ~\new_[10424]_ );
  assign \new_[16088]_  = (~\new_[17038]_  | ~\new_[5044]_ ) & (~\new_[17454]_  | ~\new_[10359]_ );
  assign \new_[16089]_  = (~\new_[17038]_  | ~\new_[5041]_ ) & (~\new_[17454]_  | ~\new_[10432]_ );
  assign \new_[16090]_  = (~\new_[17038]_  | ~\new_[5010]_ ) & (~\new_[17454]_  | ~\new_[10427]_ );
  assign \new_[16091]_  = (~\new_[17038]_  | ~\new_[4896]_ ) & (~\new_[17454]_  | ~\new_[10428]_ );
  assign \new_[16092]_  = (~\new_[17038]_  | ~\new_[4970]_ ) & (~\new_[17454]_  | ~\new_[10357]_ );
  assign \new_[16093]_  = (~\new_[17038]_  | ~\new_[5009]_ ) & (~\new_[17454]_  | ~\new_[10361]_ );
  assign \new_[16094]_  = (~\new_[16826]_  | ~\new_[4975]_ ) & (~\new_[17454]_  | ~\new_[10433]_ );
  assign \new_[16095]_  = (~\new_[16826]_  | ~\new_[4972]_ ) & (~\new_[17454]_  | ~\new_[10430]_ );
  assign \new_[16096]_  = (~\new_[17038]_  | ~\new_[5090]_ ) & (~\new_[17454]_  | ~\new_[10418]_ );
  assign \new_[16097]_  = (~\new_[17038]_  | ~\new_[5038]_ ) & (~\new_[17454]_  | ~\new_[10419]_ );
  assign \new_[16098]_  = configuration_wb_init_complete_out_reg;
  assign \new_[16099]_  = ~\new_[20456]_  & ~\new_[20305]_ ;
  assign \new_[16100]_  = \\input_register_pci_ad_reg_out_reg[29] ;
  assign \new_[16101]_  = ~\new_[16401]_ ;
  assign \new_[16102]_  = ~\new_[17558]_  | ~\new_[20515]_  | ~\new_[20513]_  | ~\new_[19922]_ ;
  assign \new_[16103]_  = ~\new_[16171]_ ;
  assign \new_[16104]_  = ~\new_[20161]_ ;
  assign \new_[16105]_  = ~\new_[17583]_  & (~\new_[19308]_  | ~\new_[20153]_ );
  assign \new_[16106]_  = ~\new_[16630]_  & (~\new_[15199]_  | ~\new_[15594]_ );
  assign \new_[16107]_  = \\input_register_pci_ad_reg_out_reg[25] ;
  assign \new_[16108]_  = parity_checker_frame_dec2_reg;
  assign \new_[16109]_  = ~\new_[16156]_ ;
  assign \new_[16110]_  = ~\new_[16155]_ ;
  assign \new_[16111]_  = ~\new_[16417]_ ;
  assign \new_[16112]_  = ~\new_[16418]_ ;
  assign \new_[16113]_  = ~\new_[16152]_ ;
  assign \new_[16114]_  = ~\new_[16151]_ ;
  assign \new_[16115]_  = \new_[17385]_  & \new_[20128]_ ;
  assign \new_[16116]_  = ~\new_[16420]_ ;
  assign \new_[16117]_  = ~\new_[16421]_ ;
  assign \new_[16118]_  = ~\new_[16422]_ ;
  assign \new_[16119]_  = ~\new_[16423]_ ;
  assign \new_[16120]_  = \new_[20340]_  & \new_[16150]_ ;
  assign \new_[16121]_  = ~\new_[16424]_ ;
  assign \new_[16122]_  = ~\new_[20340]_  | ~\new_[16384]_ ;
  assign \new_[16123]_  = ~\new_[16147]_ ;
  assign \new_[16124]_  = ~\new_[16428]_ ;
  assign \new_[16125]_  = ~\new_[16146]_ ;
  assign \new_[16126]_  = ~\new_[16429]_ ;
  assign \new_[16127]_  = \\input_register_pci_ad_reg_out_reg[15] ;
  assign \new_[16128]_  = \new_[17692]_  ? \new_[16787]_  : \new_[18840]_ ;
  assign \new_[16129]_  = \new_[20081]_  & \new_[17546]_ ;
  assign \new_[16130]_  = \\input_register_pci_ad_reg_out_reg[23] ;
  assign \new_[16131]_  = \new_[17753]_  ? \new_[16787]_  : \new_[18353]_ ;
  assign \new_[16132]_  = ~\new_[16918]_  & ~\new_[16475]_ ;
  assign \new_[16133]_  = \new_[17759]_  ? \new_[16787]_  : \new_[18944]_ ;
  assign \new_[16134]_  = \\input_register_pci_ad_reg_out_reg[20] ;
  assign \new_[16135]_  = \new_[19777]_  ? \new_[16785]_  : \new_[17642]_ ;
  assign \new_[16136]_  = \new_[17627]_  ? \new_[16787]_  : \new_[18925]_ ;
  assign \new_[16137]_  = ~\new_[16777]_  | ~\new_[17434]_ ;
  assign n16155 = ~\new_[16577]_ ;
  assign \new_[16139]_  = \new_[17758]_  ? \new_[16989]_  : \new_[19833]_ ;
  assign \new_[16140]_  = \new_[18373]_  ? \new_[16971]_  : \new_[17564]_ ;
  assign \new_[16141]_  = ~\new_[16636]_ ;
  assign \new_[16142]_  = ~wishbone_slave_unit_del_sync_req_rty_exp_clr_reg;
  assign \new_[16143]_  = \\input_register_pci_ad_reg_out_reg[26] ;
  assign \new_[16144]_  = \\input_register_pci_ad_reg_out_reg[31] ;
  assign \new_[16145]_  = ~\new_[16772]_  | ~\new_[17443]_ ;
  assign \new_[16146]_  = ~\new_[20143]_  | ~\new_[15941]_ ;
  assign \new_[16147]_  = ~\new_[20143]_  | ~\new_[15925]_ ;
  assign \new_[16148]_  = ~\new_[16451]_ ;
  assign \new_[16149]_  = \new_[17561]_  ? \new_[16973]_  : \new_[18061]_ ;
  assign \new_[16150]_  = \\input_register_pci_ad_reg_out_reg[6] ;
  assign \new_[16151]_  = ~\new_[20143]_  | ~\new_[15927]_ ;
  assign \new_[16152]_  = ~\new_[20143]_  | ~\new_[16443]_ ;
  assign \new_[16153]_  = ~\new_[16630]_ ;
  assign \new_[16154]_  = \new_[17688]_  ? \new_[16989]_  : \new_[18331]_ ;
  assign \new_[16155]_  = \new_[20143]_  & \new_[16107]_ ;
  assign \new_[16156]_  = \new_[17080]_  & \new_[15924]_ ;
  assign \new_[16157]_  = ~\new_[16620]_ ;
  assign \new_[16158]_  = \new_[15361]_  ^ \new_[17476]_ ;
  assign \new_[16159]_  = ~\new_[16457]_ ;
  assign \new_[16160]_  = ~\new_[16458]_ ;
  assign \new_[16161]_  = \new_[16776]_  & \new_[9880]_ ;
  assign \new_[16162]_  = \new_[17719]_  ? \new_[16973]_  : \new_[19737]_ ;
  assign \new_[16163]_  = \new_[18111]_  ? \new_[16910]_  : \new_[17612]_ ;
  assign \new_[16164]_  = \new_[15399]_  ^ \new_[17318]_ ;
  assign \new_[16165]_  = ~\new_[16475]_ ;
  assign \new_[16166]_  = ~\new_[16845]_  & (~\new_[17061]_  | ~\new_[11622]_ );
  assign \new_[16167]_  = \new_[17712]_  ? \new_[16973]_  : \new_[18076]_ ;
  assign \new_[16168]_  = \new_[19747]_  ? \new_[16971]_  : \new_[17650]_ ;
  assign \new_[16169]_  = \new_[14969]_  ? \new_[16997]_  : \new_[18265]_ ;
  assign \new_[16170]_  = ~\new_[16851]_  & ~\new_[16837]_ ;
  assign \new_[16171]_  = \new_[16665]_  & n16745;
  assign \new_[16172]_  = ~\new_[18523]_  | ~\new_[4627]_  | ~\new_[17576]_ ;
  assign \new_[16173]_  = \new_[15038]_  ^ \new_[16894]_ ;
  assign \new_[16174]_  = \new_[9795]_  ^ \new_[16861]_ ;
  assign \new_[16175]_  = \new_[8622]_  ^ \new_[16860]_ ;
  assign \new_[16176]_  = ~\new_[16682]_  | ~\new_[9647]_ ;
  assign \new_[16177]_  = \new_[19232]_  ? \new_[16910]_  : \new_[17759]_ ;
  assign \new_[16178]_  = \new_[19217]_  ? \new_[16910]_  : \new_[17641]_ ;
  assign \new_[16179]_  = configuration_init_complete_reg;
  assign \new_[16180]_  = \new_[19420]_  ^ \new_[16859]_ ;
  assign \new_[16181]_  = \new_[16699]_  & \new_[6322]_ ;
  assign \new_[16182]_  = \new_[16701]_  & \wbm_adr_o[5] ;
  assign \new_[16183]_  = \new_[16699]_  & \new_[17111]_ ;
  assign \new_[16184]_  = ~\new_[16476]_ ;
  assign \new_[16185]_  = \new_[16701]_  & \new_[16974]_ ;
  assign \new_[16186]_  = \new_[14995]_  ^ \new_[16897]_ ;
  assign \new_[16187]_  = \new_[9807]_  ^ \new_[16898]_ ;
  assign \new_[16188]_  = \new_[17591]_  ? \new_[16973]_  : \new_[18262]_ ;
  assign \new_[16189]_  = ~\new_[16697]_  | ~\new_[16857]_ ;
  assign \new_[16190]_  = \new_[17694]_  ? \new_[16989]_  : \new_[19819]_ ;
  assign \new_[16191]_  = \new_[16671]_  & \new_[19891]_ ;
  assign \new_[16192]_  = ~\new_[16770]_  | ~\new_[9619]_ ;
  assign \new_[16193]_  = ~\new_[16683]_  | (~\new_[16855]_  & ~\new_[17568]_ );
  assign \new_[16194]_  = ~\new_[16839]_  & ~\new_[17180]_ ;
  assign \new_[16195]_  = \new_[17194]_  & \new_[16704]_ ;
  assign \new_[16196]_  = ~\new_[16706]_  & ~\new_[16782]_ ;
  assign \new_[16197]_  = \new_[17132]_  & \new_[16703]_ ;
  assign \new_[16198]_  = \new_[17650]_  ? \new_[16989]_  : \new_[19459]_ ;
  assign \new_[16199]_  = (~\new_[17681]_  & ~\new_[19493]_  & ~\wbs_bte_i[1] ) | (~\new_[17555]_  & ~\wbs_adr_i[5]  & ~\new_[17274]_ );
  assign \new_[16200]_  = \new_[17099]_  & \new_[16705]_ ;
  assign \new_[16201]_  = ~\new_[16706]_  & ~\new_[16673]_ ;
  assign \new_[16202]_  = ~\new_[18756]_  | ~\new_[18247]_  | ~\new_[16691]_  | ~\new_[17259]_ ;
  assign \new_[16203]_  = ~\new_[14861]_  | ~\new_[14989]_  | ~\new_[16692]_  | ~\new_[17741]_ ;
  assign \new_[16204]_  = ~\new_[16844]_  | ~\new_[16648]_ ;
  assign \new_[16205]_  = input_register_pci_idsel_reg_out_reg;
  assign \new_[16206]_  = \new_[17599]_  ? \new_[16989]_  : \new_[19670]_ ;
  assign \new_[16207]_  = ~\new_[17602]_  | ~\new_[17476]_  | ~\new_[16205]_  | ~\new_[17022]_ ;
  assign \new_[16208]_  = \new_[16672]_  & \new_[5297]_ ;
  assign \new_[16209]_  = \new_[19872]_  ? \new_[20151]_  : \new_[16951]_ ;
  assign \new_[16210]_  = \\input_register_pci_ad_reg_out_reg[21] ;
  assign \new_[16211]_  = ~\new_[14614]_  & ~\new_[16734]_ ;
  assign \new_[16212]_  = \new_[16745]_  | \new_[17411]_ ;
  assign \new_[16213]_  = ~\new_[16763]_  & ~\new_[17351]_ ;
  assign \new_[16214]_  = \new_[16753]_  | \new_[17364]_ ;
  assign \new_[16215]_  = \new_[16775]_  & \new_[9879]_ ;
  assign \new_[16216]_  = \new_[16764]_  | \new_[17417]_ ;
  assign \new_[16217]_  = \new_[17097]_  & \new_[16648]_ ;
  assign \new_[16218]_  = ~\new_[17130]_  & ~\new_[16743]_ ;
  assign \new_[16219]_  = ~\new_[16918]_  & ~\new_[16819]_ ;
  assign \new_[16220]_  = \new_[17199]_  & \new_[16728]_ ;
  assign \new_[16221]_  = ~\new_[17273]_  | ~\new_[18590]_  | ~\new_[19542]_  | ~\new_[17721]_ ;
  assign \new_[16222]_  = \new_[17185]_  & \new_[16726]_ ;
  assign \new_[16223]_  = \new_[16748]_  & \new_[17167]_ ;
  assign \new_[16224]_  = ~\new_[16751]_  | ~\new_[16747]_ ;
  assign \new_[16225]_  = ~\new_[16771]_  | ~\new_[17437]_ ;
  assign \new_[16226]_  = \new_[17089]_  & \new_[16647]_ ;
  assign \new_[16227]_  = \new_[17203]_  | \new_[17228]_  | \new_[17057]_  | \new_[17214]_ ;
  assign \new_[16228]_  = \new_[19948]_  & \new_[9672]_ ;
  assign \new_[16229]_  = ~wbs_ack_o | ~\new_[16762]_  | ~\new_[20509]_ ;
  assign \new_[16230]_  = ~n16755 & (~\new_[16967]_  | ~\new_[12302]_ );
  assign \new_[16231]_  = \new_[14969]_  ? \new_[16998]_  : \new_[18689]_ ;
  assign \new_[16232]_  = \new_[14969]_  ? \new_[16864]_  : \new_[18739]_ ;
  assign \new_[16233]_  = \new_[14969]_  ? \new_[16985]_  : \new_[18832]_ ;
  assign \new_[16234]_  = \new_[17728]_  ? \new_[16989]_  : \new_[18302]_ ;
  assign \new_[16235]_  = \new_[17692]_  ? \new_[16973]_  : \new_[18510]_ ;
  assign \new_[16236]_  = \new_[17759]_  ? \new_[16989]_  : \new_[19812]_ ;
  assign \new_[16237]_  = \new_[17642]_  ? \new_[16973]_  : \new_[19826]_ ;
  assign \new_[16238]_  = \new_[17564]_  ? \new_[16973]_  : \new_[18083]_ ;
  assign \new_[16239]_  = \new_[17759]_  ? \new_[16973]_  : \new_[18161]_ ;
  assign \new_[16240]_  = \new_[17612]_  ? \new_[16989]_  : \new_[19124]_ ;
  assign \new_[16241]_  = \new_[17723]_  ? \new_[16989]_  : \new_[19679]_ ;
  assign \new_[16242]_  = \new_[17613]_  ? \new_[16973]_  : \new_[18580]_ ;
  assign \new_[16243]_  = \new_[17639]_  ? \new_[16989]_  : \new_[18203]_ ;
  assign \new_[16244]_  = \new_[17753]_  ? \new_[16989]_  : \new_[19334]_ ;
  assign \new_[16245]_  = \new_[17599]_  ? \new_[16973]_  : \new_[19021]_ ;
  assign \new_[16246]_  = \new_[17708]_  ? \new_[16973]_  : \new_[19820]_ ;
  assign \new_[16247]_  = \new_[17702]_  ? \new_[16973]_  : \new_[17900]_ ;
  assign \new_[16248]_  = \new_[17723]_  ? \new_[16973]_  : \new_[18293]_ ;
  assign \new_[16249]_  = \new_[17760]_  ? \new_[16973]_  : \new_[19114]_ ;
  assign \new_[16250]_  = \new_[17627]_  ? \new_[16989]_  : \new_[19317]_ ;
  assign \new_[16251]_  = \new_[17708]_  ? \new_[16989]_  : \new_[18284]_ ;
  assign \new_[16252]_  = \new_[17591]_  ? \new_[16989]_  : \new_[17924]_ ;
  assign \new_[16253]_  = \new_[17702]_  ? \new_[16989]_  : \new_[17853]_ ;
  assign \new_[16254]_  = \new_[17760]_  ? \new_[16989]_  : \new_[19108]_ ;
  assign \new_[16255]_  = \new_[17564]_  ? \new_[16989]_  : \new_[19739]_ ;
  assign \new_[16256]_  = \new_[17758]_  ? \new_[16973]_  : \new_[19309]_ ;
  assign \new_[16257]_  = \new_[17734]_  ? \new_[16973]_  : \new_[19000]_ ;
  assign \new_[16258]_  = \new_[17627]_  ? \new_[16973]_  : \new_[18096]_ ;
  assign \new_[16259]_  = \new_[17719]_  ? \new_[16989]_  : \new_[19726]_ ;
  assign \new_[16260]_  = \new_[17712]_  ? \new_[16989]_  : \new_[17909]_ ;
  assign \new_[16261]_  = \new_[17703]_  ? \new_[16989]_  : \new_[19818]_ ;
  assign \new_[16262]_  = \new_[17613]_  ? \new_[16989]_  : \new_[19815]_ ;
  assign \new_[16263]_  = \new_[17641]_  ? \new_[16989]_  : \new_[19026]_ ;
  assign \new_[16264]_  = \new_[17560]_  ? \new_[16989]_  : \new_[19821]_ ;
  assign \new_[16265]_  = \new_[17633]_  ? \new_[16989]_  : \new_[17955]_ ;
  assign \new_[16266]_  = \new_[17755]_  ? \new_[16973]_  : \new_[18160]_ ;
  assign \new_[16267]_  = \new_[17700]_  ? \new_[16989]_  : \new_[19741]_ ;
  assign \new_[16268]_  = \new_[17753]_  ? \new_[16973]_  : \new_[18168]_ ;
  assign \new_[16269]_  = \new_[17560]_  ? \new_[16973]_  : \new_[19017]_ ;
  assign \new_[16270]_  = \new_[17692]_  ? \new_[16989]_  : \new_[17912]_ ;
  assign \new_[16271]_  = \new_[17734]_  ? \new_[16989]_  : \new_[19463]_ ;
  assign \new_[16272]_  = \new_[17633]_  ? \new_[16973]_  : \new_[18924]_ ;
  assign \new_[16273]_  = \new_[17608]_  ? \new_[16973]_  : \new_[18175]_ ;
  assign \new_[16274]_  = \new_[17645]_  ? \new_[16973]_  : \new_[18169]_ ;
  assign \new_[16275]_  = \new_[17650]_  ? \new_[16973]_  : \new_[18179]_ ;
  assign \new_[16276]_  = \new_[17645]_  ? \new_[16989]_  : \new_[19816]_ ;
  assign \new_[16277]_  = \new_[17612]_  ? \new_[16973]_  : \new_[18107]_ ;
  assign \new_[16278]_  = \new_[17641]_  ? \new_[16973]_  : \new_[18932]_ ;
  assign \new_[16279]_  = \new_[17728]_  ? \new_[16973]_  : \new_[17892]_ ;
  assign \new_[16280]_  = \new_[17561]_  ? \new_[16989]_  : \new_[19043]_ ;
  assign \new_[16281]_  = \new_[17642]_  ? \new_[16989]_  : \new_[19342]_ ;
  assign \new_[16282]_  = \new_[17639]_  ? \new_[16973]_  : \new_[18597]_ ;
  assign \new_[16283]_  = \new_[17703]_  ? \new_[16973]_  : \new_[18174]_ ;
  assign \new_[16284]_  = \new_[17694]_  ? \new_[16973]_  : \new_[18835]_ ;
  assign \new_[16285]_  = \new_[17755]_  ? \new_[16989]_  : \new_[19807]_ ;
  assign \new_[16286]_  = \new_[17688]_  ? \new_[16973]_  : \new_[18178]_ ;
  assign \new_[16287]_  = \new_[19801]_  ? \new_[16971]_  : \new_[17591]_ ;
  assign \new_[16288]_  = \new_[19643]_  ? \new_[16971]_  : \new_[17612]_ ;
  assign \new_[16289]_  = \new_[19169]_  ? \new_[16971]_  : \new_[17642]_ ;
  assign \new_[16290]_  = \new_[18067]_  ? \new_[16971]_  : \new_[17688]_ ;
  assign \new_[16291]_  = \new_[19799]_  ? \new_[16971]_  : \new_[17703]_ ;
  assign \new_[16292]_  = \new_[18055]_  ? \new_[16971]_  : \new_[17608]_ ;
  assign \new_[16293]_  = \new_[19672]_  ? \new_[16971]_  : \new_[17753]_ ;
  assign \new_[16294]_  = \new_[19653]_  ? \new_[16971]_  : \new_[17760]_ ;
  assign \new_[16295]_  = \new_[19182]_  ? \new_[16971]_  : \new_[17613]_ ;
  assign \new_[16296]_  = \new_[19186]_  ? \new_[16971]_  : \new_[17719]_ ;
  assign \new_[16297]_  = \new_[19202]_  ? \new_[16971]_  : \new_[17627]_ ;
  assign \new_[16298]_  = \new_[19617]_  ? \new_[16971]_  : \new_[17599]_ ;
  assign \new_[16299]_  = \new_[18871]_  ? \new_[16910]_  : \new_[17723]_ ;
  assign \new_[16300]_  = \new_[19210]_  ? \new_[16910]_  : \new_[17692]_ ;
  assign \new_[16301]_  = \new_[18868]_  ? \new_[16910]_  : \new_[17560]_ ;
  assign \new_[16302]_  = \new_[19752]_  ? \new_[16910]_  : \new_[17712]_ ;
  assign \new_[16303]_  = \new_[18110]_  ? \new_[16910]_  : \new_[17591]_ ;
  assign \new_[16304]_  = \new_[19211]_  ? \new_[16910]_  : \new_[17639]_ ;
  assign \new_[16305]_  = \new_[18113]_  ? \new_[16910]_  : \new_[17734]_ ;
  assign \new_[16306]_  = \new_[19212]_  ? \new_[16910]_  : \new_[17642]_ ;
  assign \new_[16307]_  = \new_[19863]_  ? \new_[16910]_  : \new_[17700]_ ;
  assign \new_[16308]_  = \new_[19598]_  ? \new_[16910]_  : \new_[17688]_ ;
  assign \new_[16309]_  = \new_[18126]_  ? \new_[16910]_  : \new_[17608]_ ;
  assign \new_[16310]_  = \new_[18120]_  ? \new_[16910]_  : \new_[17645]_ ;
  assign \new_[16311]_  = \new_[19584]_  ? \new_[16910]_  : \new_[17753]_ ;
  assign \new_[16312]_  = \new_[18306]_  ? \new_[16910]_  : \new_[17760]_ ;
  assign \new_[16313]_  = \new_[19577]_  ? \new_[16910]_  : \new_[17719]_ ;
  assign \new_[16314]_  = \new_[19716]_  ? \new_[16910]_  : \new_[17627]_ ;
  assign \new_[16315]_  = \new_[19792]_  ? \new_[16910]_  : \new_[17599]_ ;
  assign \new_[16316]_  = \new_[18212]_  ? \new_[16910]_  : \new_[17708]_ ;
  assign \new_[16317]_  = \new_[19246]_  ? \new_[16910]_  : \new_[17633]_ ;
  assign \new_[16318]_  = \new_[18419]_  ? \new_[16971]_  : \new_[17561]_ ;
  assign \new_[16319]_  = \new_[19016]_  ? \new_[16910]_  : \new_[17564]_ ;
  assign \new_[16320]_  = \new_[19575]_  ? \new_[16987]_  : \new_[14969]_ ;
  assign \new_[16321]_  = \new_[19756]_  ? \new_[16910]_  : \new_[17758]_ ;
  assign \new_[16322]_  = \new_[19791]_  ? \new_[16910]_  : \new_[17702]_ ;
  assign \new_[16323]_  = \new_[19709]_  ? \new_[16971]_  : \new_[17723]_ ;
  assign \new_[16324]_  = \new_[18147]_  ? \new_[16971]_  : \new_[17702]_ ;
  assign \new_[16325]_  = \new_[19363]_  ? \new_[16971]_  : \new_[17633]_ ;
  assign \new_[16326]_  = \new_[18092]_  ? \new_[16971]_  : \new_[17708]_ ;
  assign \new_[16327]_  = \new_[17889]_  ? \new_[16971]_  : \new_[17758]_ ;
  assign \new_[16328]_  = \new_[19623]_  ? \new_[16971]_  : \new_[17728]_ ;
  assign \new_[16329]_  = ~\new_[17762]_  | ~\new_[14988]_  | ~\new_[16681]_  | ~\new_[14990]_ ;
  assign \new_[16330]_  = \new_[18159]_  ? \new_[16910]_  : \new_[17755]_ ;
  assign \new_[16331]_  = \new_[14969]_  ? \new_[16991]_  : \new_[19553]_ ;
  assign \new_[16332]_  = \new_[14969]_  ? \new_[16881]_  : \new_[18918]_ ;
  assign \new_[16333]_  = \new_[18166]_  ? \new_[16910]_  : \new_[17728]_ ;
  assign \new_[16334]_  = \new_[19168]_  ? \new_[16971]_  : \new_[17639]_ ;
  assign \new_[16335]_  = \new_[19784]_  ? \new_[16910]_  : \new_[17650]_ ;
  assign \new_[16336]_  = ~\new_[17678]_  | ~\new_[9798]_  | ~\new_[16649]_  | ~\new_[9808]_ ;
  assign \new_[16337]_  = \new_[18062]_  ? \new_[16971]_  : \new_[17759]_ ;
  assign \new_[16338]_  = \new_[19748]_  ? \new_[16971]_  : \new_[17755]_ ;
  assign \new_[16339]_  = \new_[19174]_  ? \new_[16971]_  : \new_[17645]_ ;
  assign \new_[16340]_  = \new_[17985]_  ? \new_[16971]_  : \new_[17734]_ ;
  assign \new_[16341]_  = \new_[18616]_  ? \new_[16983]_  : \new_[14969]_ ;
  assign \new_[16342]_  = \new_[18038]_  ? \new_[16971]_  : \new_[17641]_ ;
  assign \new_[16343]_  = \new_[14969]_  ? \new_[16888]_  : \new_[18414]_ ;
  assign \new_[16344]_  = \new_[14969]_  ? \new_[17013]_  : \new_[18970]_ ;
  assign \new_[16345]_  = \new_[17404]_  ^ \new_[17383]_ ;
  assign \new_[16346]_  = \new_[19795]_  ? \new_[16910]_  : \new_[17561]_ ;
  assign \new_[16347]_  = \new_[17978]_  ? \new_[16971]_  : \new_[17700]_ ;
  assign \new_[16348]_  = \new_[19802]_  ? \new_[16971]_  : \new_[17694]_ ;
  assign \new_[16349]_  = \new_[19686]_  ? \new_[16971]_  : \new_[17692]_ ;
  assign \new_[16350]_  = \new_[19354]_  ? \new_[16971]_  : \new_[17560]_ ;
  assign \new_[16351]_  = \new_[17896]_  ? \new_[16971]_  : \new_[17712]_ ;
  assign \new_[16352]_  = \new_[8391]_  ^ \new_[17011]_ ;
  assign \new_[16353]_  = \new_[16962]_  ^ \new_[18681]_ ;
  assign \new_[16354]_  = \\input_register_pci_ad_reg_out_reg[1] ;
  assign \new_[16355]_  = \new_[16961]_  ^ \new_[19171]_ ;
  assign \new_[16356]_  = \new_[8603]_  ^ \new_[16963]_ ;
  assign \new_[16357]_  = \new_[8392]_  ^ \new_[16958]_ ;
  assign \new_[16358]_  = \new_[16956]_  ^ \new_[9803]_ ;
  assign \new_[16359]_  = \new_[17018]_  ^ \new_[9624]_ ;
  assign \new_[16360]_  = ~\new_[20532]_  | ~\new_[9676]_  | ~\new_[17019]_ ;
  assign \new_[16361]_  = \new_[16798]_  | n16690;
  assign \new_[16362]_  = ~\new_[19343]_  | ~\new_[16798]_  | ~\new_[17254]_ ;
  assign \new_[16363]_  = ~\new_[9672]_  | ~\new_[19929]_ ;
  assign \new_[16364]_  = ~\new_[19763]_  | ~\new_[16796]_ ;
  assign \new_[16365]_  = ~\new_[18409]_  | ~\new_[16790]_ ;
  assign \new_[16366]_  = ~\new_[17943]_  | ~\new_[16805]_ ;
  assign \new_[16367]_  = \new_[20305]_  | \new_[19910]_ ;
  assign \new_[16368]_  = ~\new_[18023]_  | ~\new_[16843]_  | ~\new_[18251]_ ;
  assign \new_[16369]_  = \\input_register_pci_ad_reg_out_reg[18] ;
  assign \new_[16370]_  = ~\new_[16795]_  | ~\new_[18561]_ ;
  assign \new_[16371]_  = ~\new_[18382]_  | ~\new_[16679]_ ;
  assign \new_[16372]_  = \new_[16801]_  & \new_[16827]_ ;
  assign \new_[16373]_  = ~\new_[19590]_  | ~\new_[16797]_ ;
  assign \new_[16374]_  = ~\new_[16839]_  | ~\new_[20211]_ ;
  assign \new_[16375]_  = ~\new_[19285]_  | ~\new_[16662]_ ;
  assign \new_[16376]_  = ~\new_[16589]_ ;
  assign \new_[16377]_  = ~\new_[19284]_  | ~\new_[16783]_ ;
  assign \new_[16378]_  = ~\new_[19436]_  | ~\new_[16803]_ ;
  assign \new_[16379]_  = ~\new_[19929]_  & ~n16890;
  assign \new_[16380]_  = ~\new_[18475]_  | ~\new_[16804]_ ;
  assign \new_[16381]_  = ~\new_[16659]_  & ~\new_[17039]_ ;
  assign \new_[16382]_  = \\input_register_pci_ad_reg_out_reg[22] ;
  assign \new_[16383]_  = \new_[16670]_  | \new_[17747]_ ;
  assign \new_[16384]_  = \\input_register_pci_ad_reg_out_reg[2] ;
  assign \new_[16385]_  = ~\new_[18249]_  | ~\new_[16794]_ ;
  assign \new_[16386]_  = (~\new_[17038]_  | ~\new_[5039]_ ) & (~\new_[17454]_  | ~\new_[10420]_ );
  assign \new_[16387]_  = (~\new_[17038]_  | ~\new_[4971]_ ) & (~\new_[17454]_  | ~\new_[10429]_ );
  assign \new_[16388]_  = (~\new_[17038]_  | ~\new_[4965]_ ) & (~\new_[17454]_  | ~\new_[10423]_ );
  assign \new_[16389]_  = (~\new_[17038]_  | ~\new_[5011]_ ) & (~\new_[17454]_  | ~\new_[10435]_ );
  assign \new_[16390]_  = (~\new_[17038]_  | ~\new_[18791]_ ) & (~\new_[17454]_  | ~\new_[10355]_ );
  assign \new_[16391]_  = (~\new_[17038]_  | ~\new_[4976]_ ) & (~\new_[17454]_  | ~\new_[10351]_ );
  assign \new_[16392]_  = (~\new_[17038]_  | ~\new_[5040]_ ) & (~\new_[17454]_  | ~\new_[10421]_ );
  assign \new_[16393]_  = (~\new_[17038]_  | ~\new_[4974]_ ) & (~\new_[17454]_  | ~\new_[10354]_ );
  assign \new_[16394]_  = (~\new_[17038]_  | ~\new_[4977]_ ) & (~\new_[17454]_  | ~\new_[10434]_ );
  assign \new_[16395]_  = (~\new_[17038]_  | ~\new_[4969]_ ) & (~\new_[17454]_  | ~\new_[10426]_ );
  assign \new_[16396]_  = (~\new_[17038]_  | ~\new_[4968]_ ) & (~\new_[17454]_  | ~\new_[10353]_ );
  assign \new_[16397]_  = (~\new_[17038]_  | ~\new_[4963]_ ) & (~\new_[17454]_  | ~\new_[10362]_ );
  assign \new_[16398]_  = ~\new_[16599]_ ;
  assign \new_[16399]_  = ~pci_target_unit_pci_target_sm_read_completed_reg_reg;
  assign \new_[16400]_  = ~\new_[16602]_ ;
  assign \new_[16401]_  = ~\new_[16605]_ ;
  assign \new_[16402]_  = ~\new_[19967]_ ;
  assign \new_[16403]_  = ~\new_[16878]_  & ~\new_[17305]_ ;
  assign \new_[16404]_  = ~\new_[16607]_ ;
  assign \new_[16405]_  = \\input_register_pci_ad_reg_out_reg[11] ;
  assign \new_[16406]_  = ~\new_[16612]_ ;
  assign \new_[16407]_  = \new_[19682]_  ? \new_[16910]_  : \new_[17694]_ ;
  assign \new_[16408]_  = ~\new_[16821]_  & (~\new_[10004]_  | ~\new_[19859]_ );
  assign \new_[16409]_  = \new_[17746]_  ^ \new_[16838]_ ;
  assign \new_[16410]_  = ~\new_[16666]_  & (~\new_[13598]_  | ~\new_[18338]_ );
  assign \new_[16411]_  = ~\new_[17258]_  | ~\new_[17476]_  | ~\new_[17383]_  | ~\new_[17318]_ ;
  assign \new_[16412]_  = \new_[12012]_  ^ \new_[16909]_ ;
  assign \new_[16413]_  = \new_[17608]_  ? \new_[16989]_  : \new_[18323]_ ;
  assign \new_[16414]_  = \\input_register_pci_ad_reg_out_reg[5] ;
  assign \new_[16415]_  = ~n16380;
  assign \new_[16416]_  = \new_[20143]_  & \new_[16143]_ ;
  assign \new_[16417]_  = \new_[17080]_  & \new_[16382]_ ;
  assign \new_[16418]_  = ~\new_[20143]_  | ~\new_[16144]_ ;
  assign \new_[16419]_  = ~\new_[16631]_ ;
  assign \new_[16420]_  = \new_[17080]_  & \new_[16134]_ ;
  assign \new_[16421]_  = \new_[17080]_  & \new_[16130]_ ;
  assign \new_[16422]_  = \new_[17080]_  & \new_[16369]_ ;
  assign \new_[16423]_  = \new_[17080]_  & \new_[15926]_ ;
  assign \new_[16424]_  = ~\new_[20143]_  | ~\new_[16100]_ ;
  assign \new_[16425]_  = ~\new_[16633]_ ;
  assign \new_[16426]_  = \new_[20487]_  & \new_[20159]_ ;
  assign \new_[16427]_  = ~\new_[16634]_ ;
  assign \new_[16428]_  = \new_[17080]_  & \new_[16210]_ ;
  assign \new_[16429]_  = \new_[17080]_  & \new_[16440]_ ;
  assign \new_[16430]_  = \new_[20487]_  | \new_[20159]_ ;
  assign \new_[16431]_  = ~\new_[16635]_ ;
  assign \new_[16432]_  = ~\new_[20183]_ ;
  assign \new_[16433]_  = ~\new_[16901]_ ;
  assign \new_[16434]_  = ~\new_[16901]_ ;
  assign \new_[16435]_  = \\input_register_pci_ad_reg_out_reg[8] ;
  assign \new_[16436]_  = ~\new_[16852]_ ;
  assign \new_[16437]_  = \new_[17700]_  ? \new_[16973]_  : \new_[19407]_ ;
  assign \new_[16438]_  = ~\new_[19410]_  | ~\new_[20509]_  | ~\new_[18458]_  | ~\new_[19194]_ ;
  assign n16385 = ~\new_[16734]_ ;
  assign \new_[16440]_  = \\input_register_pci_ad_reg_out_reg[19] ;
  assign \new_[16441]_  = \new_[19218]_  ? \new_[16910]_  : \new_[17703]_ ;
  assign \new_[16442]_  = \new_[18787]_  ? \new_[16977]_  : \new_[14969]_ ;
  assign \new_[16443]_  = \\input_register_pci_ad_reg_out_reg[27] ;
  assign \new_[16444]_  = \new_[19838]_  ? \new_[16910]_  : \new_[17613]_ ;
  assign \new_[16445]_  = \new_[17273]_  & \new_[16845]_ ;
  assign \new_[16446]_  = ~\new_[16799]_  & ~\new_[20512]_ ;
  assign \new_[16447]_  = \new_[19562]_  ? \new_[17169]_  : \new_[17561]_ ;
  assign \new_[16448]_  = \new_[18086]_  ? \new_[17169]_  : \new_[17692]_ ;
  assign \new_[16449]_  = \new_[19765]_  ? \new_[17169]_  : \new_[17708]_ ;
  assign n16460 = parity_checker_frame_and_irdy_en_prev_prev_reg;
  assign \new_[16451]_  = ~\new_[17323]_  & (~\new_[17463]_  | ~\new_[17140]_ );
  assign n16495 = \new_[16107]_  ? \new_[17707]_  : \pci_ad_i[25] ;
  assign n17480 = wishbone_slave_unit_del_sync_comp_done_reg_main_reg;
  assign \new_[16454]_  = \new_[19538]_  ? \new_[17169]_  : \new_[17760]_ ;
  assign \new_[16455]_  = \new_[15110]_  ^ \new_[17141]_ ;
  assign \new_[16456]_  = \new_[17633]_  ? \new_[17150]_  : \new_[19650]_ ;
  assign \new_[16457]_  = \new_[17383]_  & \new_[16405]_ ;
  assign \new_[16458]_  = \new_[17383]_  & \new_[15985]_ ;
  assign \new_[16459]_  = \new_[16923]_  & \new_[10448]_ ;
  assign \new_[16460]_  = ~\new_[16649]_ ;
  assign \new_[16461]_  = ~\new_[16681]_ ;
  assign \new_[16462]_  = ~\new_[17486]_  | ~\new_[17762]_  | ~\new_[17128]_ ;
  assign \new_[16463]_  = ~\new_[17488]_  | ~\new_[17678]_  | ~\new_[17129]_ ;
  assign \new_[16464]_  = \new_[11880]_  ^ \new_[17058]_ ;
  assign \new_[16465]_  = ~\new_[20512]_  & (~\new_[17592]_  | ~\new_[17558]_ );
  assign n16455 = \new_[15989]_  ? n16645 : \pci_ad_i[13] ;
  assign n16465 = \new_[16013]_  ? n16645 : \pci_ad_i[4] ;
  assign n16510 = \new_[16130]_  ? \new_[17707]_  : \pci_ad_i[23] ;
  assign \new_[16469]_  = \new_[6553]_  ^ \new_[17285]_ ;
  assign \new_[16470]_  = \new_[9625]_  ^ \new_[17281]_ ;
  assign n16490 = \new_[16100]_  ? n16645 : \pci_ad_i[29] ;
  assign \new_[16472]_  = \wbm_adr_o[4]  ^ \new_[17283]_ ;
  assign \new_[16473]_  = \new_[4974]_  ^ \new_[17484]_ ;
  assign \new_[16474]_  = ~\new_[16678]_ ;
  assign \new_[16475]_  = ~\new_[16906]_  | ~\new_[4962]_ ;
  assign \new_[16476]_  = ~\new_[17671]_  | ~\new_[16906]_  | ~\new_[17489]_ ;
  assign \new_[16477]_  = ~pci_target_unit_del_sync_comp_rty_exp_clr_reg;
  assign \new_[16478]_  = \new_[17702]_  ? \new_[17150]_  : \new_[18024]_ ;
  assign \new_[16479]_  = ~\wbs_bte_i[0]  & (~\new_[17274]_  | ~\wbs_bte_i[1] );
  assign \new_[16480]_  = \new_[17688]_  ? \new_[17150]_  : \new_[19725]_ ;
  assign \new_[16481]_  = \new_[17599]_  ? \new_[17150]_  : \new_[19803]_ ;
  assign \new_[16482]_  = \new_[17627]_  ? \new_[17150]_  : \new_[19164]_ ;
  assign \new_[16483]_  = \new_[9644]_  ^ \new_[17102]_ ;
  assign \new_[16484]_  = ~\new_[16859]_  & (~\new_[10859]_  | ~\new_[17359]_ );
  assign \new_[16485]_  = ~\new_[16907]_  & (~\new_[17795]_  | ~\new_[11331]_ );
  assign \new_[16486]_  = \new_[19673]_  ? \new_[17169]_  : \new_[17694]_ ;
  assign \new_[16487]_  = \new_[9796]_  ^ \new_[17139]_ ;
  assign \new_[16488]_  = \new_[19235]_  ? \new_[17169]_  : \new_[17723]_ ;
  assign n16420 = \new_[15928]_  ? n16645 : \pci_ad_i[0] ;
  assign \new_[16490]_  = \new_[17933]_  ? \new_[17169]_  : \new_[17650]_ ;
  assign n16400 = \new_[15924]_  ? n16645 : \pci_ad_i[17] ;
  assign \new_[16492]_  = \new_[17612]_  ? \new_[17150]_  : \new_[18162]_ ;
  assign n16450 = \new_[15986]_  ? \new_[17707]_  : \pci_ad_i[3] ;
  assign \new_[16494]_  = \new_[19764]_  ? \new_[17169]_  : \new_[17599]_ ;
  assign n16445 = \new_[15985]_  ? \new_[17707]_  : \pci_ad_i[12] ;
  assign \new_[16496]_  = \new_[17700]_  ? \new_[17150]_  : \new_[19148]_ ;
  assign \new_[16497]_  = ~\new_[19933]_  & ~\new_[5297]_ ;
  assign \new_[16498]_  = \new_[17561]_  ? \new_[17150]_  : \new_[19291]_ ;
  assign \new_[16499]_  = \new_[17256]_  ? \new_[11345]_  : \new_[11344]_ ;
  assign \new_[16500]_  = ~\new_[20336]_  | ~\new_[16881]_ ;
  assign n16470 = \new_[16027]_  ? \new_[17707]_  : \pci_ad_i[9] ;
  assign n16405 = \new_[15925]_  ? n16645 : \pci_ad_i[30] ;
  assign \new_[16503]_  = ~\new_[16892]_  & ~\new_[17000]_ ;
  assign \new_[16504]_  = ~\new_[16936]_  & ~\new_[16933]_ ;
  assign \new_[16505]_  = ~\new_[16932]_  & ~\new_[16925]_ ;
  assign \new_[16506]_  = ~\new_[16923]_  & ~\new_[16868]_ ;
  assign n16505 = \new_[16127]_  ? \new_[17707]_  : \pci_ad_i[15] ;
  assign \new_[16508]_  = ~\new_[16692]_ ;
  assign \new_[16509]_  = ~\new_[16691]_ ;
  assign \new_[16510]_  = ~\new_[16948]_  & (~\new_[8385]_  | ~\new_[8387]_ );
  assign \new_[16511]_  = ~\new_[16863]_  & (~\new_[4459]_  | ~\new_[4460]_ );
  assign n16440 = ~\new_[17483]_  & (~\new_[17261]_  | ~\new_[17140]_ );
  assign \new_[16513]_  = ~\new_[16848]_  | (~\new_[17654]_  & ~\new_[18338]_ );
  assign \new_[16514]_  = ~\new_[17020]_  | (~\new_[17656]_  & ~\new_[19859]_ );
  assign \new_[16515]_  = ~\new_[16676]_ ;
  assign \new_[16516]_  = ~\new_[13869]_  | ~\new_[12039]_  | ~\new_[16903]_  | ~\new_[17467]_ ;
  assign \new_[16517]_  = ~\new_[13869]_  | ~\new_[16852]_  | ~\new_[16903]_  | ~\new_[17365]_ ;
  assign n16395 = \new_[15923]_  ? n16645 : \pci_ad_i[7] ;
  assign \new_[16519]_  = \new_[17608]_  ? \new_[17150]_  : \new_[19806]_ ;
  assign \new_[16520]_  = \new_[17760]_  ? \new_[17150]_  : \new_[19151]_ ;
  assign \new_[16521]_  = \new_[17692]_  ? \new_[17150]_  : \new_[19292]_ ;
  assign \new_[16522]_  = \new_[17694]_  ? \new_[17150]_  : \new_[17998]_ ;
  assign \new_[16523]_  = \new_[8394]_  ^ \new_[17175]_ ;
  assign \new_[16524]_  = \new_[17753]_  ? \new_[17150]_  : \new_[18157]_ ;
  assign \new_[16525]_  = \new_[17560]_  ? \new_[17150]_  : \new_[18562]_ ;
  assign \new_[16526]_  = \new_[17723]_  ? \new_[17150]_  : \new_[19743]_ ;
  assign \new_[16527]_  = \new_[17564]_  ? \new_[17150]_  : \new_[17964]_ ;
  assign \new_[16528]_  = \new_[17759]_  ? \new_[17150]_  : \new_[18989]_ ;
  assign \new_[16529]_  = \new_[17650]_  ? \new_[17150]_  : \new_[17997]_ ;
  assign \new_[16530]_  = \new_[17708]_  ? \new_[17150]_  : \new_[19162]_ ;
  assign \new_[16531]_  = \new_[17642]_  ? \new_[17150]_  : \new_[17994]_ ;
  assign \new_[16532]_  = \new_[17645]_  ? \new_[17150]_  : \new_[19512]_ ;
  assign \new_[16533]_  = \new_[17728]_  ? \new_[17150]_  : \new_[19158]_ ;
  assign \new_[16534]_  = \new_[17719]_  ? \new_[17150]_  : \new_[19669]_ ;
  assign \new_[16535]_  = \new_[17734]_  ? \new_[17150]_  : \new_[19808]_ ;
  assign \new_[16536]_  = \new_[17758]_  ? \new_[17150]_  : \new_[19160]_ ;
  assign \new_[16537]_  = \new_[17641]_  ? \new_[17150]_  : \new_[19266]_ ;
  assign \new_[16538]_  = \new_[17703]_  ? \new_[17150]_  : \new_[19560]_ ;
  assign \new_[16539]_  = \new_[17639]_  ? \new_[17150]_  : \new_[19138]_ ;
  assign \new_[16540]_  = \new_[17591]_  ? \new_[17150]_  : \new_[19811]_ ;
  assign \new_[16541]_  = \new_[17755]_  ? \new_[17150]_  : \new_[19582]_ ;
  assign \new_[16542]_  = \new_[17712]_  ? \new_[17150]_  : \new_[19810]_ ;
  assign \new_[16543]_  = \new_[11343]_  ^ \new_[17173]_ ;
  assign \new_[16544]_  = \new_[17613]_  ? \new_[17150]_  : \new_[19724]_ ;
  assign \new_[16545]_  = (~\new_[17580]_  & ~\new_[5047]_  & ~\new_[10371]_ ) | (~\new_[17241]_  & ~\new_[19136]_  & ~\new_[5046]_ );
  assign \new_[16546]_  = \new_[19208]_  ? \new_[17169]_  : \new_[17564]_ ;
  assign \new_[16547]_  = \new_[19015]_  ? \new_[17169]_  : \new_[17560]_ ;
  assign \new_[16548]_  = \new_[19785]_  ? \new_[17169]_  : \new_[17591]_ ;
  assign \new_[16549]_  = \new_[18200]_  ? \new_[17169]_  : \new_[17734]_ ;
  assign \new_[16550]_  = \new_[18201]_  ? \new_[17169]_  : \new_[17642]_ ;
  assign \new_[16551]_  = \new_[18223]_  ? \new_[17169]_  : \new_[17613]_ ;
  assign \new_[16552]_  = \new_[18222]_  ? \new_[17169]_  : \new_[17719]_ ;
  assign \new_[16553]_  = \new_[18258]_  ? \new_[17169]_  : \new_[17728]_ ;
  assign \new_[16554]_  = \new_[19782]_  ? \new_[17169]_  : \new_[17627]_ ;
  assign \new_[16555]_  = \new_[19082]_  ? \new_[17169]_  : \new_[17712]_ ;
  assign \new_[16556]_  = \new_[19256]_  ? \new_[17169]_  : \new_[17641]_ ;
  assign \new_[16557]_  = \new_[14969]_  ? \new_[17067]_  : \new_[18754]_ ;
  assign \new_[16558]_  = \new_[19190]_  ? \new_[17103]_  : \new_[14969]_ ;
  assign \new_[16559]_  = \new_[19137]_  ? \new_[17169]_  : \new_[17639]_ ;
  assign \new_[16560]_  = \new_[18202]_  ? \new_[17169]_  : \new_[17700]_ ;
  assign \new_[16561]_  = \new_[19864]_  ? \new_[17169]_  : \new_[17702]_ ;
  assign \new_[16562]_  = \new_[19013]_  ? \new_[17169]_  : \new_[17755]_ ;
  assign \new_[16563]_  = \new_[17838]_  ? \new_[17169]_  : \new_[17633]_ ;
  assign \new_[16564]_  = \new_[19790]_  ? \new_[17169]_  : \new_[17612]_ ;
  assign \new_[16565]_  = \new_[19117]_  ? \new_[17169]_  : \new_[17753]_ ;
  assign \new_[16566]_  = \new_[19759]_  ? \new_[17169]_  : \new_[17645]_ ;
  assign \new_[16567]_  = \new_[19271]_  ? \new_[17169]_  : \new_[17759]_ ;
  assign \new_[16568]_  = \new_[19789]_  ? \new_[17169]_  : \new_[17608]_ ;
  assign \new_[16569]_  = \new_[19783]_  ? \new_[17169]_  : \new_[17758]_ ;
  assign \new_[16570]_  = \new_[19120]_  ? \new_[17169]_  : \new_[17703]_ ;
  assign \new_[16571]_  = \new_[18213]_  ? \new_[17169]_  : \new_[17688]_ ;
  assign \new_[16572]_  = ~\new_[19929]_ ;
  assign \new_[16573]_  = configuration_pci_err_cs_bit8_reg;
  assign \new_[16574]_  = \\configuration_isr_bit2_0_reg[2] ;
  assign \new_[16575]_  = \\configuration_isr_bit2_0_reg[0] ;
  assign \new_[16576]_  = ~\new_[16647]_ ;
  assign \new_[16577]_  = ~\new_[16886]_  | ~\new_[3944]_ ;
  assign \new_[16578]_  = \new_[16912]_  | \new_[4627]_ ;
  assign \new_[16579]_  = ~\new_[19484]_  | ~\new_[17013]_ ;
  assign \new_[16580]_  = ~\new_[16955]_  & ~\new_[9801]_ ;
  assign \new_[16581]_  = \new_[16992]_  | \new_[17793]_ ;
  assign \new_[16582]_  = ~\new_[19173]_  | ~\new_[16985]_ ;
  assign \new_[16583]_  = ~\new_[19403]_  | ~\new_[16864]_ ;
  assign \new_[16584]_  = ~\new_[20082]_  | ~\new_[16886]_ ;
  assign \new_[16585]_  = ~\new_[16819]_ ;
  assign \new_[16586]_  = ~\new_[19671]_  | ~\new_[16997]_ ;
  assign \new_[16587]_  = ~\new_[18144]_  | ~\new_[16888]_ ;
  assign n16425 = ~\new_[16970]_  | ~\new_[17565]_ ;
  assign \new_[16589]_  = ~\new_[20515]_  | ~\new_[20512]_  | ~\new_[20043]_ ;
  assign \new_[16590]_  = ~\new_[18492]_  | ~\new_[17001]_ ;
  assign \new_[16591]_  = \new_[16858]_  | \new_[17233]_ ;
  assign \new_[16592]_  = ~\new_[18427]_  | ~\new_[16896]_ ;
  assign \new_[16593]_  = ~n17360 & ~\new_[16964]_ ;
  assign \new_[16594]_  = ~\new_[16966]_  | ~\new_[19909]_ ;
  assign \new_[16595]_  = ~\new_[17934]_  | ~\new_[16991]_ ;
  assign \new_[16596]_  = ~\new_[17292]_  | ~\new_[15191]_  | ~\new_[20292]_  | ~\new_[10855]_ ;
  assign \new_[16597]_  = n16685 ? n16930 : \new_[13688]_ ;
  assign \new_[16598]_  = n16675 ? n16750 : \new_[4008]_ ;
  assign \new_[16599]_  = wishbone_slave_unit_pci_initiator_if_write_req_int_reg;
  assign \new_[16600]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[0] ;
  assign n16480 = ~\new_[16843]_ ;
  assign \new_[16602]_  = ~\new_[19885]_ ;
  assign \new_[16603]_  = ~\new_[16839]_ ;
  assign \new_[16604]_  = ~\new_[16877]_  & ~\new_[19416]_ ;
  assign \new_[16605]_  = ~\new_[19903]_  | ~\new_[19911]_ ;
  assign \new_[16606]_  = ~\new_[16788]_ ;
  assign \new_[16607]_  = ~\new_[20071]_  | ~\new_[19911]_ ;
  assign \new_[16608]_  = \new_[16885]_  & \new_[17474]_ ;
  assign \new_[16609]_  = ~\new_[16687]_ ;
  assign \new_[16610]_  = ~\new_[16673]_ ;
  assign \new_[16611]_  = ~\new_[17305]_  | ~\new_[20319]_ ;
  assign \new_[16612]_  = ~\new_[17249]_  & ~\new_[17030]_ ;
  assign \new_[16613]_  = ~\new_[17063]_  | ~\new_[17300]_ ;
  assign \new_[16614]_  = \new_[17368]_  | \new_[17063]_ ;
  assign \new_[16615]_  = ~\new_[17063]_  | ~\new_[17433]_ ;
  assign \new_[16616]_  = ~\new_[16683]_ ;
  assign \new_[16617]_  = ~\new_[16851]_  & ~\new_[17251]_ ;
  assign \new_[16618]_  = ~\new_[16871]_  & (~n16745 | ~\new_[9617]_ );
  assign \new_[16619]_  = ~\new_[19393]_  | ~\new_[17024]_  | ~\new_[20488]_ ;
  assign \new_[16620]_  = ~\new_[17030]_  | (~\new_[9287]_  & ~\new_[19312]_ );
  assign \new_[16621]_  = \new_[15272]_  ^ \new_[15925]_ ;
  assign n16430 = \new_[15941]_  ? \new_[17707]_  : \pci_ad_i[24] ;
  assign n16475 = \new_[16032]_  ? \new_[17707]_  : \pci_ad_i[14] ;
  assign n16415 = \new_[15927]_  ? \new_[17707]_  : \pci_ad_i[28] ;
  assign n16410 = \new_[15926]_  ? \new_[17707]_  : \pci_ad_i[16] ;
  assign n16435 = \new_[15948]_  ? \new_[17707]_  : \pci_ad_i[10] ;
  assign n16380 = ~\new_[16878]_ ;
  assign n16485 = \\configuration_i_wb_init_complete_sync_sync_data_out_reg[0] ;
  assign n16515 = \new_[16134]_  ? \new_[17707]_  : \pci_ad_i[20] ;
  assign \new_[16630]_  = ~\new_[19781]_  | ~n16500;
  assign \new_[16631]_  = \new_[17383]_  & \new_[15989]_ ;
  assign \new_[16632]_  = ~\new_[16677]_ ;
  assign \new_[16633]_  = \new_[17383]_  & \new_[15948]_ ;
  assign \new_[16634]_  = \new_[17383]_  & \new_[16127]_ ;
  assign \new_[16635]_  = \new_[17383]_  & \new_[16027]_ ;
  assign \new_[16636]_  = \new_[17383]_  & \new_[16032]_ ;
  assign \new_[16637]_  = ~\new_[18967]_  | ~\new_[17003]_ ;
  assign \new_[16638]_  = ~\new_[20487]_  & ~\new_[20068]_ ;
  assign \new_[16639]_  = ~\new_[19277]_  | ~\new_[16998]_ ;
  assign \new_[16640]_  = ~\new_[17006]_  & ~\new_[17222]_ ;
  assign \new_[16641]_  = ~\new_[16969]_  | ~\new_[9807]_ ;
  assign \new_[16642]_  = ~\new_[16968]_  | ~\new_[14995]_ ;
  assign n16600 = \new_[16443]_  ? \new_[17707]_  : \pci_ad_i[27] ;
  assign \new_[16644]_  = \new_[17196]_  & \new_[17170]_ ;
  assign \new_[16645]_  = \new_[17091]_  & \new_[17159]_ ;
  assign \new_[16646]_  = \new_[17083]_  & \new_[17185]_ ;
  assign \new_[16647]_  = \new_[17082]_  & \new_[5008]_ ;
  assign \new_[16648]_  = ~\new_[17130]_  & ~\new_[19345]_ ;
  assign \new_[16649]_  = \new_[17129]_  & \new_[9795]_ ;
  assign \new_[16650]_  = ~\new_[9623]_  | ~\new_[18523]_ ;
  assign n16565 = \new_[16382]_  ? n16645 : \pci_ad_i[22] ;
  assign n17340 = configuration_sync_isr_2_sync_del_bit_reg;
  assign pci_req_oe_o = pci_io_mux_req_iob_en_out_reg;
  assign \new_[16654]_  = (~\new_[17452]_  | ~\new_[13134]_ ) & (~\new_[17817]_  | ~\new_[17546]_ );
  assign \new_[16655]_  = ~\new_[16901]_ ;
  assign n16530 = \new_[16144]_  ? \new_[16179]_  : \pci_ad_i[31] ;
  assign \new_[16657]_  = ~\new_[17152]_  & ~\new_[17800]_ ;
  assign \new_[16658]_  = ~\new_[16901]_ ;
  assign \new_[16659]_  = \new_[19282]_  ^ \new_[18545]_ ;
  assign \new_[16660]_  = \new_[8394]_  ^ \new_[8548]_ ;
  assign \new_[16661]_  = ~\new_[16906]_ ;
  assign \new_[16662]_  = ~\new_[17777]_  | ~\new_[17268]_ ;
  assign \new_[16663]_  = \new_[17429]_  ^ \new_[17423]_ ;
  assign \new_[16664]_  = ~\new_[16868]_ ;
  assign \new_[16665]_  = ~\new_[16871]_ ;
  assign \new_[16666]_  = ~\new_[16848]_ ;
  assign n16545 = \new_[16205]_  ? \new_[17707]_  : pci_idsel_i;
  assign \new_[16668]_  = ~\new_[17012]_ ;
  assign \new_[16669]_  = \new_[17425]_  ^ \new_[17427]_ ;
  assign \new_[16670]_  = ~\new_[16882]_ ;
  assign \new_[16671]_  = ~\new_[20305]_  & ~\new_[20303]_ ;
  assign \new_[16672]_  = ~\new_[19933]_ ;
  assign \new_[16673]_  = ~\new_[19159]_  | ~\new_[15424]_  | ~n16500;
  assign \new_[16674]_  = ~\new_[16990]_ ;
  assign n16525 = \new_[16143]_  ? \new_[17707]_  : \pci_ad_i[26] ;
  assign \new_[16676]_  = ~\new_[4972]_  | ~\new_[5011]_  | ~\new_[17094]_  | ~\new_[17573]_ ;
  assign \new_[16677]_  = ~\new_[17383]_  | ~\new_[16435]_ ;
  assign \new_[16678]_  = ~\new_[19923]_  | ~\new_[20529]_  | ~\new_[17592]_ ;
  assign \new_[16679]_  = ~\new_[17367]_  | ~\new_[17777]_ ;
  assign \new_[16680]_  = \new_[17346]_  ^ \new_[17413]_ ;
  assign \new_[16681]_  = \new_[17128]_  & \new_[15038]_ ;
  assign \new_[16682]_  = ~\new_[9619]_  | ~\new_[9618]_  | ~\new_[17102]_  | ~\new_[17495]_ ;
  assign \new_[16683]_  = ~\new_[15399]_  | ~\new_[17253]_  | ~\new_[17746]_ ;
  assign \new_[16684]_  = ~\new_[17181]_  & ~\new_[14614]_ ;
  assign \new_[16685]_  = ~\new_[17231]_  & ~\new_[17137]_ ;
  assign \new_[16686]_  = ~\new_[17126]_  & ~\new_[17220]_ ;
  assign \new_[16687]_  = \new_[17264]_  & \new_[4009]_ ;
  assign n16550 = \new_[16210]_  ? \new_[16179]_  : \pci_ad_i[21] ;
  assign n16580 = \new_[16405]_  ? \new_[16179]_  : \pci_ad_i[11] ;
  assign n16560 = \new_[16369]_  ? \new_[16179]_  : \pci_ad_i[18] ;
  assign \new_[16691]_  = ~\new_[17139]_  & ~\new_[17193]_ ;
  assign \new_[16692]_  = ~\new_[17141]_  & ~\new_[17198]_ ;
  assign \new_[16693]_  = \new_[15073]_  ^ \new_[17291]_ ;
  assign \new_[16694]_  = \new_[9275]_  ^ \new_[17449]_ ;
  assign \new_[16695]_  = \new_[9810]_  ^ \new_[17440]_ ;
  assign \new_[16696]_  = \new_[8389]_  ^ \new_[17470]_ ;
  assign \new_[16697]_  = \new_[17664]_  ? \new_[8548]_  : \new_[17640]_ ;
  assign n16935 = pci_target_unit_del_sync_req_rty_exp_reg_reg;
  assign \new_[16699]_  = \new_[17285]_  & \new_[6553]_ ;
  assign \new_[16700]_  = \new_[17281]_  & \new_[9625]_ ;
  assign \new_[16701]_  = \new_[17283]_  & \wbm_adr_o[4] ;
  assign \new_[16702]_  = ~\new_[17445]_  | ~\new_[17384]_  | ~\new_[17721]_ ;
  assign \new_[16703]_  = \new_[17192]_  & \new_[17285]_ ;
  assign \new_[16704]_  = \new_[17197]_  & \new_[17438]_ ;
  assign \new_[16705]_  = \new_[17074]_  & \new_[17283]_ ;
  assign \new_[16706]_  = ~\new_[17558]_  | ~\new_[20529]_  | ~\new_[19922]_ ;
  assign n16585 = \new_[16414]_  ? \new_[17707]_  : \pci_ad_i[5] ;
  assign \new_[16708]_  = ~\new_[4971]_  | ~\new_[4972]_  | ~\new_[17176]_  | ~\new_[17461]_ ;
  assign \new_[16709]_  = \new_[17404]_  ^ \new_[17403]_ ;
  assign \new_[16710]_  = \new_[17405]_  ^ \new_[17380]_ ;
  assign \new_[16711]_  = \new_[17418]_  ^ \new_[17426]_ ;
  assign \new_[16712]_  = \new_[17345]_  ^ \new_[17415]_ ;
  assign \new_[16713]_  = \new_[17347]_  ^ \new_[17421]_ ;
  assign \new_[16714]_  = \new_[17416]_  ^ \new_[17356]_ ;
  assign \new_[16715]_  = \new_[17339]_  ^ \new_[17355]_ ;
  assign \new_[16716]_  = \new_[17410]_  ^ \new_[17353]_ ;
  assign \new_[16717]_  = \new_[17420]_  ^ \new_[17362]_ ;
  assign \new_[16718]_  = \new_[17352]_  ^ \new_[17408]_ ;
  assign \new_[16719]_  = \new_[17349]_  ^ \new_[17366]_ ;
  assign \new_[16720]_  = \new_[17369]_  ^ \new_[17430]_ ;
  assign \new_[16721]_  = \new_[17407]_  ^ \new_[17428]_ ;
  assign \new_[16722]_  = \new_[17419]_  ^ \new_[17340]_ ;
  assign \new_[16723]_  = \new_[17343]_  ^ \new_[17406]_ ;
  assign \new_[16724]_  = ~configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg;
  assign \new_[16725]_  = ~configuration_sync_isr_2_delayed_bckp_bit_reg;
  assign \new_[16726]_  = \new_[17201]_  & \new_[6554]_ ;
  assign \new_[16727]_  = \new_[17153]_  | \new_[9791]_ ;
  assign \new_[16728]_  = \new_[17078]_  & \new_[17166]_ ;
  assign \new_[16729]_  = ~\new_[17382]_  & ~\new_[17044]_ ;
  assign \new_[16730]_  = \new_[17142]_  | \new_[18971]_ ;
  assign \new_[16731]_  = \new_[17194]_  & \new_[17190]_ ;
  assign \new_[16732]_  = ~\new_[17206]_  & ~\new_[17056]_ ;
  assign n16540 = \new_[17144]_  | n16645;
  assign \new_[16734]_  = \new_[17098]_  | \new_[3944]_ ;
  assign \new_[16735]_  = ~\new_[17163]_  | ~\new_[17257]_ ;
  assign \new_[16736]_  = ~\new_[17699]_  | ~\new_[17164]_  | ~\new_[17451]_ ;
  assign \new_[16737]_  = \new_[17119]_  & \new_[17156]_ ;
  assign \new_[16738]_  = ~\new_[17050]_  & ~\new_[17239]_ ;
  assign \new_[16739]_  = \new_[17083]_  & \new_[17091]_ ;
  assign \new_[16740]_  = ~\new_[19690]_  | ~\new_[17067]_ ;
  assign \new_[16741]_  = ~\new_[17225]_  & ~\new_[17051]_ ;
  assign \new_[16742]_  = ~\new_[17227]_  & ~\new_[17219]_ ;
  assign \new_[16743]_  = ~\new_[17097]_  | ~\new_[17179]_ ;
  assign \new_[16744]_  = ~\new_[17533]_  | ~\new_[17138]_  | ~\new_[17471]_ ;
  assign \new_[16745]_  = \new_[17224]_  | \new_[17223]_ ;
  assign \new_[16746]_  = ~\new_[17216]_  & ~\new_[17202]_ ;
  assign \new_[16747]_  = ~\new_[17226]_  & ~\new_[17217]_ ;
  assign \new_[16748]_  = \new_[17182]_  & \new_[17108]_ ;
  assign \new_[16749]_  = ~\new_[17060]_  & ~\new_[17208]_ ;
  assign \new_[16750]_  = ~\new_[17041]_  & ~\new_[17213]_ ;
  assign \new_[16751]_  = ~\new_[17042]_  & ~\new_[17205]_ ;
  assign \new_[16752]_  = \new_[17201]_  & \new_[17091]_ ;
  assign \new_[16753]_  = \new_[17118]_  | \new_[17070]_ ;
  assign \new_[16754]_  = \new_[17110]_  & \new_[17187]_ ;
  assign \new_[16755]_  = \new_[17082]_  & \new_[17089]_ ;
  assign \new_[16756]_  = ~\new_[17171]_  | ~\new_[17120]_ ;
  assign \new_[16757]_  = ~\new_[17229]_  & ~\new_[17235]_ ;
  assign \new_[16758]_  = ~\new_[17789]_  | ~\new_[17167]_  | ~\new_[17469]_ ;
  assign \new_[16759]_  = ~\new_[17280]_  & ~\new_[17204]_ ;
  assign \new_[16760]_  = ~\new_[17209]_  & ~\new_[17114]_ ;
  assign \new_[16761]_  = ~\new_[17073]_  & ~\new_[17117]_ ;
  assign \new_[16762]_  = \new_[20536]_  & \new_[17750]_ ;
  assign \new_[16763]_  = \new_[17124]_  | \new_[17424]_ ;
  assign \new_[16764]_  = \new_[17232]_  | \new_[17230]_ ;
  assign \new_[16765]_  = ~\new_[17210]_  & ~\new_[17277]_ ;
  assign \new_[16766]_  = ~\new_[17234]_  & ~\new_[17278]_ ;
  assign \new_[16767]_  = ~\new_[17237]_  & ~\new_[17275]_ ;
  assign \new_[16768]_  = ~\new_[17236]_  & ~\new_[17066]_ ;
  assign \new_[16769]_  = ~\new_[17068]_  & ~\new_[17240]_ ;
  assign \new_[16770]_  = ~\new_[9618]_  | ~\new_[17174]_  | ~\new_[9623]_ ;
  assign \new_[16771]_  = (~\new_[17306]_  | ~\new_[18798]_ ) & (~\new_[9799]_  | ~\new_[19224]_ );
  assign \new_[16772]_  = (~\new_[17439]_  | ~\new_[17812]_ ) & (~\new_[9268]_  | ~\new_[19273]_ );
  assign \new_[16773]_  = ~\new_[17053]_  & ~\new_[17055]_ ;
  assign \new_[16774]_  = ~\new_[17133]_  | (~\new_[17800]_  & ~\new_[9622]_ );
  assign \new_[16775]_  = \new_[17680]_  ^ \new_[17456]_ ;
  assign \new_[16776]_  = \new_[17737]_  ^ \new_[17448]_ ;
  assign \new_[16777]_  = (~\new_[18901]_  | ~\new_[13771]_ ) & (~\new_[13219]_  | ~\new_[17303]_ );
  assign \new_[16778]_  = ~wishbone_slave_unit_del_sync_req_comp_pending_sample_reg;
  assign \new_[16779]_  = ~\\configuration_sync_cache_lsize_to_wb_bits_reg[3] ;
  assign \new_[16780]_  = ~pci_target_unit_del_sync_req_comp_pending_sample_reg;
  assign \new_[16781]_  = ~\new_[16966]_ ;
  assign \new_[16782]_  = \new_[20146]_ ;
  assign \new_[16783]_  = ~\new_[17262]_  | ~\new_[13720]_ ;
  assign \new_[16784]_  = \new_[17271]_  & \new_[18338]_ ;
  assign \new_[16785]_  = \new_[17260]_  & \new_[19859]_ ;
  assign \new_[16786]_  = ~\new_[20043]_  & ~\new_[20514]_ ;
  assign \new_[16787]_  = ~\new_[17260]_  | ~\new_[10074]_ ;
  assign \new_[16788]_  = ~\new_[17269]_  & ~\new_[3995]_ ;
  assign \new_[16789]_  = \new_[17262]_  & \new_[18338]_ ;
  assign \new_[16790]_  = ~\new_[17299]_  | ~\new_[17268]_ ;
  assign \new_[16791]_  = ~\new_[20398]_ ;
  assign \new_[16792]_  = \new_[17063]_  & \new_[17557]_ ;
  assign \new_[16793]_  = \new_[20177]_  | \new_[17450]_ ;
  assign \new_[16794]_  = \new_[18338]_  | \new_[17095]_ ;
  assign \new_[16795]_  = \new_[18338]_  | \new_[17255]_ ;
  assign \new_[16796]_  = ~\new_[17341]_  | ~\new_[17268]_ ;
  assign \new_[16797]_  = ~\new_[17268]_  | ~\new_[17603]_ ;
  assign \new_[16798]_  = \new_[17267]_  & \new_[9910]_ ;
  assign \new_[16799]_  = ~\new_[20043]_  | ~\new_[20514]_ ;
  assign \new_[16800]_  = ~\new_[16978]_ ;
  assign \new_[16801]_  = ~\new_[17474]_  & ~\new_[17054]_ ;
  assign \new_[16802]_  = ~n16770 & ~\new_[17308]_ ;
  assign \new_[16803]_  = ~\new_[17271]_  | ~\new_[13720]_ ;
  assign \new_[16804]_  = ~\new_[17367]_  | ~\new_[17341]_ ;
  assign \new_[16805]_  = ~\new_[17367]_  | ~\new_[17299]_ ;
  assign \new_[16806]_  = \new_[17436]_  | \new_[17367]_ ;
  assign \new_[16807]_  = ~\new_[6326]_  | ~\new_[17533]_  | ~\new_[18545]_ ;
  assign \new_[16808]_  = ~\new_[17434]_  | ~\new_[17252]_ ;
  assign \new_[16809]_  = \new_[17132]_  & \new_[17189]_ ;
  assign \new_[16810]_  = ~\new_[17049]_  | (~\new_[17878]_  & ~\new_[9621]_ );
  assign \new_[16811]_  = ~\new_[20174]_  & (~\new_[15216]_  | ~\new_[20340]_ );
  assign n16570 = \new_[16384]_  ? \new_[17707]_  : \pci_ad_i[2] ;
  assign n16535 = \new_[16150]_  ? \new_[16179]_  : \pci_ad_i[6] ;
  assign n16590 = \new_[16435]_  ? \new_[16179]_  : \pci_ad_i[8] ;
  assign n16595 = \new_[16440]_  ? \new_[16179]_  : \pci_ad_i[19] ;
  assign \new_[16816]_  = \new_[17102]_  & \new_[9644]_ ;
  assign n16555 = \new_[16354]_  ? \new_[16179]_  : \pci_ad_i[1] ;
  assign \new_[16818]_  = ~\new_[17238]_  & ~\new_[17048]_ ;
  assign \new_[16819]_  = ~\new_[17134]_  | ~\new_[17077]_ ;
  assign \new_[16820]_  = ~\\pci_target_unit_del_sync_req_sync_sync_data_out_reg[0] ;
  assign \new_[16821]_  = ~\new_[17020]_ ;
  assign \new_[16822]_  = ~\new_[9622]_  | ~\new_[18523]_ ;
  assign \new_[16823]_  = ~\new_[9647]_  | ~\new_[18523]_ ;
  assign \new_[16824]_  = ~\new_[9619]_  | ~\new_[18523]_ ;
  assign \new_[16825]_  = ~\new_[9644]_  | ~\new_[18523]_ ;
  assign \new_[16826]_  = ~\new_[17027]_ ;
  assign \new_[16827]_  = ~\new_[20489]_  & ~\new_[20159]_ ;
  assign \new_[16828]_  = ~\new_[20159]_  & ~\new_[17474]_ ;
  assign \new_[16829]_  = ~\new_[17748]_  & ~\new_[20128]_ ;
  assign \new_[16830]_  = ~\new_[17125]_  & ~\new_[17037]_ ;
  assign \new_[16831]_  = ~\new_[17065]_  & ~\new_[17211]_ ;
  assign \new_[16832]_  = ~\new_[14614]_  & ~n16500;
  assign \new_[16833]_  = ~\new_[20128]_  & ~\new_[20488]_ ;
  assign \new_[16834]_  = ~\new_[17215]_  & ~\new_[17218]_ ;
  assign \new_[16835]_  = \new_[17099]_  & \new_[17178]_ ;
  assign \new_[16836]_  = ~\new_[17385]_ ;
  assign \new_[16837]_  = ~\new_[17033]_ ;
  assign \new_[16838]_  = ~\new_[17383]_ ;
  assign \new_[16839]_  = ~\new_[17084]_  | ~\new_[17544]_ ;
  assign \new_[16840]_  = ~\new_[17040]_  & ~\new_[17212]_ ;
  assign \new_[16841]_  = ~\new_[19750]_  | ~\new_[17131]_ ;
  assign \new_[16842]_  = \new_[17155]_  & \new_[17171]_ ;
  assign \new_[16843]_  = ~pci_target_unit_del_sync_comp_done_reg_main_reg;
  assign \new_[16844]_  = \new_[17162]_  & \new_[17168]_ ;
  assign \new_[16845]_  = ~\new_[17061]_  & ~\new_[11622]_ ;
  assign \new_[16846]_  = \new_[17880]_  & \new_[20229]_ ;
  assign \new_[16847]_  = \new_[17880]_  ^ \new_[20229]_ ;
  assign \new_[16848]_  = \new_[13598]_  | \new_[18338]_ ;
  assign \new_[16849]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2] ;
  assign \new_[16850]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[0] ;
  assign \new_[16851]_  = ~\new_[20072]_ ;
  assign \new_[16852]_  = ~\new_[14614]_ ;
  assign \new_[16853]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0] ;
  assign pci_irdy_oe_o = pci_io_mux_irdy_iob_en_out_reg;
  assign \new_[16855]_  = ~\new_[17253]_ ;
  assign n16615 = \\pci_target_unit_del_sync_rty_exp_back_prop_sync_sync_data_out_reg[0] ;
  assign \new_[16857]_  = ~\new_[17367]_ ;
  assign \new_[16858]_  = \new_[17515]_  ^ \new_[18789]_ ;
  assign \new_[16859]_  = ~\new_[10859]_  & ~\new_[17359]_ ;
  assign \new_[16860]_  = \new_[17470]_  | \new_[8389]_ ;
  assign \new_[16861]_  = ~\new_[17129]_ ;
  assign n16640 = \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[0] ;
  assign \new_[16863]_  = ~\new_[17638]_  | ~\new_[17293]_ ;
  assign \new_[16864]_  = ~\new_[17457]_  | ~\new_[17557]_ ;
  assign \new_[16865]_  = ~\new_[17379]_  & ~\new_[17397]_ ;
  assign \new_[16866]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1] ;
  assign \new_[16867]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1] ;
  assign \new_[16868]_  = \\wishbone_slave_unit_del_sync_req_sync_sync_data_out_reg[0] ;
  assign \new_[16869]_  = ~\new_[17394]_  & ~\new_[17375]_ ;
  assign \new_[16870]_  = ~\new_[17396]_  & ~\new_[17399]_ ;
  assign \new_[16871]_  = wishbone_slave_unit_pci_initiator_sm_mabort2_reg;
  assign n16610 = \\wishbone_slave_unit_del_sync_done_sync_sync_data_out_reg[0] ;
  assign \new_[16873]_  = ~pci_target_unit_del_sync_comp_flush_out_reg;
  assign \new_[16874]_  = ~\new_[17579]_  & (~\new_[13612]_  | ~\new_[13221]_ );
  assign \new_[16875]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[2] ;
  assign \new_[16876]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0] ;
  assign \new_[16877]_  = wishbone_slave_unit_del_sync_comp_flush_out_reg;
  assign \new_[16878]_  = ~pci_target_unit_pci_target_sm_bckp_trdy_reg_reg;
  assign \new_[16879]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2] ;
  assign \new_[16880]_  = ~\new_[17454]_  | ~\new_[4460]_ ;
  assign \new_[16881]_  = ~\new_[17368]_  | ~\new_[17446]_ ;
  assign \new_[16882]_  = ~\new_[17460]_  & ~\new_[18615]_ ;
  assign \new_[16883]_  = \new_[17296]_  & \new_[18338]_ ;
  assign \new_[16884]_  = \new_[11345]_  ^ \new_[11343]_ ;
  assign \new_[16885]_  = ~\new_[17054]_ ;
  assign \new_[16886]_  = ~\new_[17098]_ ;
  assign \new_[16887]_  = \new_[10876]_  ^ \new_[11344]_ ;
  assign \new_[16888]_  = ~\new_[17433]_  | ~\new_[17457]_ ;
  assign \new_[16889]_  = ~\new_[17113]_ ;
  assign \new_[16890]_  = ~\new_[17122]_ ;
  assign \new_[16891]_  = ~\new_[13150]_  & (~\new_[17756]_  | ~n17495);
  assign \new_[16892]_  = ~\new_[17548]_  | ~\new_[5038]_  | ~\new_[4963]_ ;
  assign \new_[16893]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3] ;
  assign \new_[16894]_  = ~\new_[17128]_ ;
  assign \new_[16895]_  = ~\new_[17314]_  & ~\new_[17372]_ ;
  assign \new_[16896]_  = ~\new_[17436]_  | ~\new_[17777]_ ;
  assign \new_[16897]_  = ~\new_[15073]_  | ~\new_[15110]_  | ~\new_[17588]_  | ~\new_[17486]_ ;
  assign \new_[16898]_  = ~\new_[9810]_  | ~\new_[9796]_  | ~\new_[17492]_  | ~\new_[17488]_ ;
  assign \new_[16899]_  = ~\new_[17576]_  | ~n17010 | ~\new_[17722]_ ;
  assign \new_[16900]_  = \new_[17587]_  & \new_[17341]_ ;
  assign \new_[16901]_  = ~\new_[17549]_ ;
  assign n17495 = configuration_sync_pci_err_cs_8_sync_del_bit_reg;
  assign \new_[16903]_  = ~\new_[17441]_  & ~\new_[15199]_ ;
  assign \new_[16904]_  = ~\new_[17181]_ ;
  assign \new_[16905]_  = \new_[18968]_  ^ \new_[17523]_ ;
  assign \new_[16906]_  = \new_[17438]_  & \new_[4974]_ ;
  assign \new_[16907]_  = ~\new_[17061]_ ;
  assign \new_[16908]_  = ~\new_[17344]_  | ~\new_[9623]_ ;
  assign \new_[16909]_  = \new_[17384]_  & \new_[17721]_ ;
  assign \new_[16910]_  = \new_[17324]_  & \new_[19859]_ ;
  assign \new_[16911]_  = \new_[17587]_  & \new_[17299]_ ;
  assign \new_[16912]_  = ~\new_[20205]_ ;
  assign \new_[16913]_  = ~\new_[17387]_  & ~\new_[17378]_ ;
  assign \new_[16914]_  = ~\new_[17393]_  & ~\new_[17391]_ ;
  assign \new_[16915]_  = ~\new_[17288]_  & ~\new_[17381]_ ;
  assign \new_[16916]_  = ~\new_[17309]_  & ~\new_[17371]_ ;
  assign \new_[16917]_  = ~\new_[17389]_  & ~\new_[17398]_ ;
  assign \new_[16918]_  = ~\new_[4977]_  | ~\new_[4975]_  | ~\new_[17671]_ ;
  assign \new_[16919]_  = ~\new_[17301]_  & ~\new_[17361]_ ;
  assign \new_[16920]_  = ~\new_[17302]_  & ~\new_[17400]_ ;
  assign \new_[16921]_  = ~\new_[17402]_  & ~\new_[17307]_ ;
  assign \new_[16922]_  = ~\new_[17386]_  & ~\new_[17390]_ ;
  assign \new_[16923]_  = \new_[17447]_  | n17480;
  assign \new_[16924]_  = ~\new_[17298]_  & ~\new_[17392]_ ;
  assign \new_[16925]_  = \new_[17769]_  ^ \new_[17783]_ ;
  assign \new_[16926]_  = \new_[17542]_  ^ \new_[17798]_ ;
  assign \new_[16927]_  = \new_[17677]_  ^ \new_[17672]_ ;
  assign \new_[16928]_  = \new_[17485]_  ^ \new_[17547]_ ;
  assign \new_[16929]_  = \new_[17799]_  ^ \new_[17691]_ ;
  assign \new_[16930]_  = \new_[17504]_  ^ \new_[17682]_ ;
  assign \new_[16931]_  = \new_[17481]_  ^ \new_[17569]_ ;
  assign \new_[16932]_  = \new_[17690]_  ^ \new_[17575]_ ;
  assign \new_[16933]_  = \new_[17739]_  ^ \new_[17673]_ ;
  assign \new_[16934]_  = \new_[17530]_  ^ \new_[17514]_ ;
  assign \new_[16935]_  = \new_[17766]_  ^ \new_[17663]_ ;
  assign \new_[16936]_  = \new_[17491]_  ^ \new_[17716]_ ;
  assign \new_[16937]_  = \new_[20378]_  ^ \new_[17683]_ ;
  assign \new_[16938]_  = \new_[17570]_  ^ \new_[17478]_ ;
  assign \new_[16939]_  = \new_[17697]_  ^ \new_[17772]_ ;
  assign \new_[16940]_  = \new_[17563]_  ^ \new_[17554]_ ;
  assign \new_[16941]_  = \new_[17784]_  ^ \new_[17480]_ ;
  assign \new_[16942]_  = \new_[17611]_  ^ \new_[17590]_ ;
  assign \new_[16943]_  = \new_[17594]_  ^ \new_[17705]_ ;
  assign \new_[16944]_  = \new_[17686]_  ^ \new_[17630]_ ;
  assign \new_[16945]_  = \new_[20023]_  ^ \new_[17584]_ ;
  assign \new_[16946]_  = \new_[17718]_  ^ \new_[17518]_ ;
  assign \new_[16947]_  = \new_[17541]_  ^ \new_[17676]_ ;
  assign \new_[16948]_  = \new_[17805]_  ? \new_[8387]_  : \new_[8386]_ ;
  assign \new_[16949]_  = ~\new_[20174]_ ;
  assign \new_[16950]_  = \new_[17525]_  ^ \new_[17781]_ ;
  assign \new_[16951]_  = \new_[19498]_  ? \new_[11961]_  : \new_[17764]_ ;
  assign n16605 = parity_checker_frame_and_irdy_en_prev_reg;
  assign n16630 = \\configuration_isr_bit0_sync_sync_data_out_reg[0] ;
  assign \new_[16954]_  = ~n16520;
  assign \new_[16955]_  = ~\\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[2] ;
  assign \new_[16956]_  = \\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[1] ;
  assign n16620 = \\configuration_pci_err_cs_bits_sync_sync_data_out_reg[0] ;
  assign \new_[16958]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[3] ;
  assign \new_[16959]_  = ~\new_[17147]_ ;
  assign \new_[16960]_  = ~\new_[17148]_ ;
  assign \new_[16961]_  = \\pci_target_unit_fifos_wb_clk_inGreyCount_reg[0] ;
  assign \new_[16962]_  = \\pci_target_unit_fifos_wb_clk_inGreyCount_reg[1] ;
  assign \new_[16963]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[2] ;
  assign \new_[16964]_  = ~\\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[1] ;
  assign \new_[16965]_  = ~\new_[17183]_ ;
  assign \new_[16966]_  = ~\new_[17567]_  & ~\new_[18502]_ ;
  assign \new_[16967]_  = ~\new_[16901]_  & ~n16775;
  assign \new_[16968]_  = ~\new_[17142]_ ;
  assign \new_[16969]_  = ~\new_[17153]_ ;
  assign \new_[16970]_  = ~n16845 & ~\new_[10010]_ ;
  assign \new_[16971]_  = \new_[17313]_  & \new_[19859]_ ;
  assign \new_[16972]_  = ~\new_[17077]_ ;
  assign \new_[16973]_  = ~\new_[17313]_  | ~\new_[10074]_ ;
  assign \new_[16974]_  = ~\new_[17444]_  & ~\new_[17780]_ ;
  assign \new_[16975]_  = \new_[17436]_  & \new_[17603]_ ;
  assign \new_[16976]_  = \new_[17367]_  & \new_[17603]_ ;
  assign \new_[16977]_  = \new_[17771]_  & \new_[17300]_ ;
  assign \new_[16978]_  = ~\new_[17468]_  | ~\new_[8385]_ ;
  assign \new_[16979]_  = \new_[17459]_  & \new_[17662]_ ;
  assign \new_[16980]_  = ~\new_[17454]_  | ~\new_[4458]_ ;
  assign \new_[16981]_  = ~\new_[17664]_  | (~\new_[8224]_  & ~\new_[17640]_ );
  assign \new_[16982]_  = ~\new_[17454]_  | ~\new_[4459]_ ;
  assign \new_[16983]_  = \new_[17771]_  & \new_[17433]_ ;
  assign \new_[16984]_  = \new_[17435]_  & \new_[18338]_ ;
  assign \new_[16985]_  = ~\new_[17446]_  | ~\new_[17771]_ ;
  assign \new_[16986]_  = ~\new_[17454]_  | ~\new_[11133]_ ;
  assign \new_[16987]_  = \new_[17368]_  & \new_[17557]_ ;
  assign \new_[16988]_  = ~\new_[17334]_  & ~\new_[17544]_ ;
  assign \new_[16989]_  = ~\new_[17324]_  | ~\new_[10074]_ ;
  assign \new_[16990]_  = ~\new_[17311]_  & ~wbm_ack_i;
  assign \new_[16991]_  = ~\new_[17300]_  | ~\new_[17457]_ ;
  assign \new_[16992]_  = \new_[14969]_  | \new_[17310]_ ;
  assign \new_[16993]_  = \new_[17750]_  & \new_[20508]_ ;
  assign \new_[16994]_  = ~\new_[17305]_  | ~\new_[18729]_ ;
  assign \new_[16995]_  = ~\new_[17454]_  | ~\new_[10360]_ ;
  assign \new_[16996]_  = ~\new_[17384]_  & (~\new_[11691]_  | ~\new_[11882]_ );
  assign \new_[16997]_  = ~\new_[17368]_  | ~\new_[17300]_ ;
  assign \new_[16998]_  = ~\new_[17368]_  | ~\new_[17433]_ ;
  assign \new_[16999]_  = ~\new_[17464]_  & ~\new_[17574]_ ;
  assign \new_[17000]_  = ~\new_[4977]_  | ~\new_[17466]_  | ~\new_[5044]_ ;
  assign \new_[17001]_  = ~\new_[17436]_  | ~\new_[17299]_ ;
  assign \new_[17002]_  = \new_[17313]_  | \new_[17324]_ ;
  assign \new_[17003]_  = ~\new_[17436]_  | ~\new_[17341]_ ;
  assign \new_[17004]_  = (~\new_[9677]_  | ~\new_[9799]_ ) & (~\new_[18798]_  | ~\new_[18199]_ );
  assign \new_[17005]_  = ~\new_[17437]_  | (~\new_[9677]_  & ~\new_[19224]_ );
  assign \new_[17006]_  = \new_[17854]_  ^ \new_[17959]_ ;
  assign \new_[17007]_  = ~\new_[17441]_  | (~\new_[19583]_  & ~\new_[15199]_ );
  assign \new_[17008]_  = \new_[17589]_  ^ \new_[17866]_ ;
  assign \new_[17009]_  = (~\new_[8688]_  | ~\new_[9268]_ ) & (~\new_[17812]_  | ~\new_[18890]_ );
  assign n16625 = \\configuration_isr_bit2_sync_sync_data_out_reg[0] ;
  assign \new_[17011]_  = ~\\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[1] ;
  assign \new_[17012]_  = (~pci_stop_i | ~\new_[17509]_ ) & (~\new_[18325]_  | ~\new_[9287]_ );
  assign \new_[17013]_  = \new_[17370]_  | \new_[17715]_ ;
  assign \new_[17014]_  = \new_[8599]_  ^ \new_[8201]_ ;
  assign \new_[17015]_  = \new_[20101]_  ^ \new_[20143]_ ;
  assign \new_[17016]_  = ~\new_[17395]_  & ~\new_[17377]_ ;
  assign \new_[17017]_  = \new_[9488]_  ^ \new_[18056]_ ;
  assign \new_[17018]_  = \\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[0] ;
  assign \new_[17019]_  = ~\new_[17308]_ ;
  assign \new_[17020]_  = \new_[10004]_  | \new_[19859]_ ;
  assign \new_[17021]_  = ~\new_[9618]_  | ~\new_[18523]_ ;
  assign \new_[17022]_  = ~\new_[20156]_ ;
  assign \new_[17023]_  = ~\new_[17388]_  & ~\new_[17401]_ ;
  assign \new_[17024]_  = ~\new_[20177]_ ;
  assign \new_[17025]_  = ~\new_[15015]_  & ~\new_[16852]_ ;
  assign \new_[17026]_  = ~\new_[18729]_  & ~\new_[12039]_ ;
  assign \new_[17027]_  = ~\new_[17038]_ ;
  assign \new_[17028]_  = \new_[13678]_  & \new_[19781]_ ;
  assign \new_[17029]_  = ~wbm_ack_i & ~wbm_err_i;
  assign \new_[17030]_  = ~\new_[18584]_  | ~\new_[9287]_ ;
  assign \new_[17031]_  = ~\new_[17383]_  | ~\new_[20143]_ ;
  assign \new_[17032]_  = ~\new_[17385]_  & ~\new_[20131]_ ;
  assign \new_[17033]_  = ~\new_[20127]_ ;
  assign \new_[17034]_  = ~\new_[17443]_  | (~\new_[8688]_  & ~\new_[19273]_ );
  assign \new_[17035]_  = ~\new_[17294]_  & ~\new_[17290]_ ;
  assign \new_[17036]_  = \new_[17409]_  | \new_[17412]_ ;
  assign \new_[17037]_  = \new_[18047]_  ^ \new_[6325]_ ;
  assign \new_[17038]_  = ~\new_[18392]_  & ~\new_[17646]_ ;
  assign \new_[17039]_  = \new_[19610]_  ^ \new_[6319]_ ;
  assign \new_[17040]_  = ~\new_[17731]_  & (~\new_[17052]_  | ~\new_[9637]_ );
  assign \new_[17041]_  = ~\new_[17751]_  & (~\new_[10485]_  | ~\new_[16210]_ );
  assign \new_[17042]_  = ~\new_[17526]_  & (~\new_[16893]_  | ~n17250);
  assign \new_[17043]_  = \\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[0] ;
  assign \new_[17044]_  = ~\new_[20319]_ ;
  assign \new_[17045]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0] ;
  assign \new_[17046]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[0] ;
  assign \new_[17047]_  = output_backup_irdy_en_out_reg;
  assign \new_[17048]_  = ~\new_[17535]_  & (~\new_[10399]_  | ~\new_[15924]_ );
  assign \new_[17049]_  = ~\new_[17344]_ ;
  assign \new_[17050]_  = ~\new_[17593]_  & (~\new_[10401]_  | ~\new_[15926]_ );
  assign \new_[17051]_  = ~\new_[17787]_  & (~\new_[10398]_  | ~\new_[15989]_ );
  assign \new_[17052]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[3] ;
  assign \new_[17053]_  = ~\new_[17506]_  & (~\new_[10403]_  | ~\new_[16130]_ );
  assign \new_[17054]_  = \new_[19393]_  | \new_[17802]_ ;
  assign \new_[17055]_  = ~\new_[17786]_  & (~\new_[10486]_  | ~\new_[16382]_ );
  assign \new_[17056]_  = \new_[19366]_  ^ \new_[6552]_ ;
  assign \new_[17057]_  = ~\new_[17528]_  & (~\new_[8395]_  | ~\new_[16853]_ );
  assign \new_[17058]_  = \new_[11331]_  | \new_[12012]_  | \new_[17795]_  | \new_[11622]_ ;
  assign \new_[17059]_  = \new_[4458]_  & \new_[11133]_ ;
  assign \new_[17060]_  = \new_[18987]_  ^ \new_[6310]_ ;
  assign \new_[17061]_  = \new_[17795]_  | \new_[11331]_ ;
  assign \new_[17062]_  = ~n16635;
  assign \new_[17063]_  = ~\new_[17370]_ ;
  assign \new_[17064]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1] ;
  assign \new_[17065]_  = \new_[13679]_  ^ \new_[18020]_ ;
  assign \new_[17066]_  = \new_[19564]_  ^ \new_[6306]_ ;
  assign \new_[17067]_  = \new_[17715]_  | \new_[17740]_ ;
  assign \new_[17068]_  = \new_[18748]_  ^ \new_[6323]_ ;
  assign n16675 = \\wishbone_slave_unit_del_sync_comp_sync_sync_data_out_reg[0] ;
  assign \new_[17070]_  = ~\new_[17792]_  & (~\new_[13437]_  | ~\new_[16867]_ );
  assign n16685 = \\pci_target_unit_del_sync_comp_sync_sync_data_out_reg[0] ;
  assign \new_[17072]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[1] ;
  assign \new_[17073]_  = \new_[19572]_  ^ \new_[6328]_ ;
  assign \new_[17074]_  = ~\new_[17531]_  & ~\new_[17729]_ ;
  assign \new_[17075]_  = \new_[19869]_  ^ \new_[18046]_ ;
  assign \new_[17076]_  = \\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[1] ;
  assign \new_[17077]_  = ~\new_[17516]_  & ~\new_[17767]_ ;
  assign \new_[17078]_  = ~\new_[17803]_  & ~\new_[17730]_ ;
  assign n16660 = \\pci_target_unit_del_sync_rty_exp_sync_sync_data_out_reg[0] ;
  assign \new_[17080]_  = ~\new_[17318]_ ;
  assign \new_[17081]_  = \\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2] ;
  assign \new_[17082]_  = \new_[17571]_  & \new_[17489]_ ;
  assign \new_[17083]_  = ~\new_[17532]_  & ~\new_[17537]_ ;
  assign \new_[17084]_  = ~\new_[17334]_ ;
  assign n16650 = \\configuration_sync_isr_2_delete_sync_sync_data_out_reg[0] ;
  assign \new_[17086]_  = ~\new_[17628]_  & (~\new_[12448]_  | ~\new_[12011]_ );
  assign \new_[17087]_  = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[2] ;
  assign n16695 = \\pci_target_unit_del_sync_done_sync_sync_data_out_reg[0] ;
  assign \new_[17089]_  = \new_[17521]_  & \new_[17671]_ ;
  assign \new_[17090]_  = ~\new_[17523]_  & (~\new_[10412]_  | ~\new_[10534]_ );
  assign \new_[17091]_  = ~\new_[17572]_  & ~\new_[17607]_ ;
  assign \new_[17092]_  = \new_[9794]_  ^ \new_[19126]_ ;
  assign \new_[17093]_  = \new_[19392]_  ^ \new_[18084]_ ;
  assign \new_[17094]_  = ~\new_[17768]_  & ~\new_[17679]_ ;
  assign \new_[17095]_  = ~\new_[17435]_ ;
  assign \new_[17096]_  = \new_[14614]_  & \new_[13678]_ ;
  assign \new_[17097]_  = ~\new_[17512]_  & ~\new_[17780]_ ;
  assign \new_[17098]_  = ~\new_[17805]_  | ~\new_[8387]_ ;
  assign \new_[17099]_  = ~\new_[17674]_  & ~\new_[17742]_ ;
  assign \new_[17100]_  = ~\new_[13689]_  | ~\new_[18962]_  | ~\new_[19011]_ ;
  assign \new_[17101]_  = \new_[10410]_  ^ \new_[18437]_ ;
  assign \new_[17102]_  = ~\new_[17800]_  & ~\new_[18786]_ ;
  assign \new_[17103]_  = \new_[17771]_  & \new_[17557]_ ;
  assign \new_[17104]_  = ~\new_[17727]_  & ~\new_[17713]_ ;
  assign \new_[17105]_  = \new_[18680]_  ^ \new_[18027]_ ;
  assign \new_[17106]_  = \new_[20230]_  ^ \new_[19272]_ ;
  assign \new_[17107]_  = \new_[19163]_  ^ \new_[20189]_ ;
  assign \new_[17108]_  = ~\new_[17556]_  & ~\new_[17801]_ ;
  assign \new_[17109]_  = ~\new_[17601]_  & ~\new_[17706]_ ;
  assign \new_[17110]_  = ~\new_[17666]_  & ~\new_[17709]_ ;
  assign \new_[17111]_  = ~\new_[17562]_  & ~\new_[17717]_ ;
  assign \new_[17112]_  = \new_[15114]_  ^ \new_[18122]_ ;
  assign \new_[17113]_  = (~pci_irdy_i | ~\new_[19583]_ ) & (~\new_[17047]_  | ~\new_[15480]_ );
  assign \new_[17114]_  = \new_[19409]_  ^ \new_[6315]_ ;
  assign \new_[17115]_  = ~pci_target_unit_del_sync_req_rty_exp_clr_reg;
  assign \new_[17116]_  = ~\new_[17493]_  & ~\new_[17524]_ ;
  assign \new_[17117]_  = \new_[18568]_  ^ \new_[6311]_ ;
  assign \new_[17118]_  = ~\new_[17775]_  & (~\new_[13216]_  | ~\new_[16876]_ );
  assign \new_[17119]_  = ~\new_[17730]_  & ~\new_[17607]_ ;
  assign \new_[17120]_  = ~\new_[17494]_  & ~\new_[17763]_ ;
  assign \new_[17121]_  = ~\new_[17545]_  & (~\new_[10481]_  | ~\new_[16144]_ );
  assign \new_[17122]_  = pci_trdy_i ? \new_[9287]_  : n16775;
  assign \new_[17123]_  = ~\new_[20082]_ ;
  assign \new_[17124]_  = ~\new_[17487]_  & (~\new_[13761]_  | ~\new_[16867]_ );
  assign \new_[17125]_  = \new_[17821]_  ^ \new_[6303]_ ;
  assign \new_[17126]_  = \new_[19576]_  ^ \new_[6313]_ ;
  assign \new_[17127]_  = ~\new_[17782]_  & (~\new_[10409]_  | ~\new_[15927]_ );
  assign \new_[17128]_  = \new_[17588]_  & \new_[15073]_ ;
  assign \new_[17129]_  = \new_[17492]_  & \new_[9810]_ ;
  assign \new_[17130]_  = ~\wbm_adr_o[4]  | ~\new_[17490]_  | ~\wbm_adr_o[3] ;
  assign \new_[17131]_  = ~\new_[17777]_  | ~\new_[17587]_ ;
  assign \new_[17132]_  = ~\new_[17493]_  & ~\new_[17601]_ ;
  assign \new_[17133]_  = ~\new_[17800]_  | ~\new_[9622]_ ;
  assign \new_[17134]_  = ~\new_[17635]_  & ~\new_[17779]_ ;
  assign \new_[17135]_  = ~\new_[17778]_  & ~\new_[17494]_ ;
  assign \new_[17136]_  = ~\new_[17704]_  & ~\new_[17574]_ ;
  assign \new_[17137]_  = ~\new_[17655]_  & (~\new_[17046]_  | ~\new_[9635]_ );
  assign \new_[17138]_  = ~\new_[17582]_  & ~\new_[17607]_ ;
  assign \new_[17139]_  = ~\new_[9810]_  | ~\new_[9790]_  | ~\new_[17488]_  | ~\new_[9794]_ ;
  assign \new_[17140]_  = \new_[17744]_  & \new_[17505]_ ;
  assign \new_[17141]_  = ~\new_[15073]_  | ~\new_[15123]_  | ~\new_[17486]_  | ~\new_[15114]_ ;
  assign \new_[17142]_  = ~\new_[17667]_  | ~\new_[14988]_ ;
  assign \new_[17143]_  = \\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[2] ;
  assign \new_[17144]_  = configuration_rst_inactive_reg;
  assign \new_[17145]_  = ~\\configuration_sync_cache_lsize_to_wb_bits_reg[2] ;
  assign \new_[17146]_  = ~\\configuration_sync_cache_lsize_to_wb_bits_reg[4] ;
  assign \new_[17147]_  = \\configuration_sync_cache_lsize_to_wb_bits_reg[7] ;
  assign \new_[17148]_  = \\configuration_sync_cache_lsize_to_wb_bits_reg[5] ;
  assign \new_[17149]_  = configuration_sync_command_bit_reg;
  assign \new_[17150]_  = \new_[17622]_  | \new_[19859]_ ;
  assign \new_[17151]_  = ~\new_[17520]_  & ~\new_[11326]_ ;
  assign \new_[17152]_  = ~\new_[17495]_  | ~\new_[9622]_ ;
  assign \new_[17153]_  = ~\new_[17698]_  | ~\new_[9798]_ ;
  assign \new_[17154]_  = ~\new_[17791]_  & ~\new_[17597]_ ;
  assign \new_[17155]_  = ~\new_[17585]_  & ~\new_[17714]_ ;
  assign \new_[17156]_  = ~\new_[17582]_  & ~\new_[17732]_ ;
  assign \new_[17157]_  = ~\new_[17742]_  & ~\new_[17733]_ ;
  assign \new_[17158]_  = ~\new_[17648]_  | ~n17340;
  assign \new_[17159]_  = ~\new_[17785]_  & ~\new_[17661]_ ;
  assign \new_[17160]_  = ~\new_[17550]_  & ~\new_[17620]_ ;
  assign \new_[17161]_  = ~\new_[17597]_  & ~\new_[17675]_ ;
  assign \new_[17162]_  = ~\new_[17801]_  & ~\new_[17684]_ ;
  assign \new_[17163]_  = ~\new_[17805]_  & ~\new_[8387]_ ;
  assign \new_[17164]_  = ~\new_[17714]_  & ~\new_[17551]_ ;
  assign \new_[17165]_  = ~\new_[17674]_  & ~\new_[17729]_ ;
  assign \new_[17166]_  = ~\new_[17539]_  & ~\new_[17537]_ ;
  assign \new_[17167]_  = ~\new_[17684]_  & ~\new_[17522]_ ;
  assign \new_[17168]_  = ~\new_[17522]_  & ~\new_[17791]_ ;
  assign \new_[17169]_  = ~\new_[17622]_  & ~\new_[10074]_ ;
  assign \new_[17170]_  = \new_[17548]_  & \new_[17662]_ ;
  assign \new_[17171]_  = ~\new_[17551]_  & ~\new_[17778]_ ;
  assign \new_[17172]_  = ~\new_[17732]_  & ~\new_[17659]_ ;
  assign \new_[17173]_  = \new_[17771]_  & \new_[11344]_ ;
  assign \new_[17174]_  = ~\new_[17800]_  & ~\new_[17540]_ ;
  assign \new_[17175]_  = \new_[17587]_  & \new_[8226]_ ;
  assign \new_[17176]_  = ~\new_[17550]_  & ~\new_[17666]_ ;
  assign \new_[17177]_  = ~\new_[17661]_  & ~\new_[17773]_ ;
  assign \new_[17178]_  = ~\new_[17733]_  & ~\new_[17585]_ ;
  assign \new_[17179]_  = ~\new_[17507]_  & ~\new_[17556]_ ;
  assign \new_[17180]_  = ~\new_[17722]_  | ~wbm_ack_i;
  assign \new_[17181]_  = ~\new_[19058]_  | ~\new_[19088]_  | ~\new_[8386]_ ;
  assign \new_[17182]_  = ~\new_[17512]_  & ~\new_[17507]_ ;
  assign \new_[17183]_  = \\configuration_sync_cache_lsize_to_wb_bits_reg[6] ;
  assign \new_[17184]_  = ~\new_[17788]_  & ~\new_[17620]_ ;
  assign \new_[17185]_  = ~\new_[17539]_  & ~\new_[17717]_ ;
  assign \new_[17186]_  = ~\new_[17659]_  & ~\new_[17670]_ ;
  assign \new_[17187]_  = ~\new_[17767]_  & ~\new_[17788]_ ;
  assign \new_[17188]_  = ~\new_[17773]_  & ~\new_[17704]_ ;
  assign \new_[17189]_  = ~\new_[17706]_  & ~\new_[17730]_ ;
  assign \new_[17190]_  = ~\new_[17516]_  & ~\new_[17779]_ ;
  assign \new_[17191]_  = \new_[17587]_  & \new_[17603]_ ;
  assign \new_[17192]_  = ~\new_[17508]_  & ~\new_[17524]_ ;
  assign \new_[17193]_  = ~\new_[18438]_  | ~\new_[17678]_  | ~\new_[9798]_ ;
  assign \new_[17194]_  = ~\new_[17770]_  & ~\new_[17635]_ ;
  assign \new_[17195]_  = ~\wbm_adr_o[30]  | ~\new_[17789]_  | ~\wbm_adr_o[29] ;
  assign \new_[17196]_  = ~\new_[17665]_  & ~\new_[17779]_ ;
  assign \new_[17197]_  = \new_[17637]_  & \new_[17489]_ ;
  assign \new_[17198]_  = ~\new_[14911]_  | ~\new_[17762]_  | ~\new_[14988]_ ;
  assign \new_[17199]_  = ~\new_[17669]_  & ~\new_[17785]_ ;
  assign \new_[17200]_  = ~\wbm_adr_o[29]  | ~\new_[17699]_  | ~\wbm_adr_o[28] ;
  assign \new_[17201]_  = ~\new_[17598]_  & ~\new_[17562]_ ;
  assign \new_[17202]_  = ~\new_[17776]_  & (~\new_[10483]_  | ~\new_[16143]_ );
  assign \new_[17203]_  = ~\new_[17605]_  & (~\new_[8397]_  | ~\new_[16849]_ );
  assign \new_[17204]_  = \new_[17891]_  ^ \new_[6308]_ ;
  assign \new_[17205]_  = ~\new_[17604]_  & (~\new_[16849]_  | ~n17285);
  assign \new_[17206]_  = \new_[19349]_  ^ \new_[6316]_ ;
  assign \new_[17207]_  = \new_[18901]_  ^ \new_[13217]_ ;
  assign \new_[17208]_  = \new_[18779]_  ^ \new_[6309]_ ;
  assign \new_[17209]_  = \new_[18150]_  ^ \new_[6314]_ ;
  assign \new_[17210]_  = \new_[17876]_  ^ \new_[6304]_ ;
  assign \new_[17211]_  = \new_[13686]_  ^ \new_[18917]_ ;
  assign \new_[17212]_  = ~\new_[17566]_  & (~\new_[17087]_  | ~\new_[9636]_ );
  assign \new_[17213]_  = ~\new_[17479]_  & (~\new_[10402]_  | ~\new_[16134]_ );
  assign \new_[17214]_  = ~\new_[17631]_  & (~\new_[8398]_  | ~\new_[16893]_ );
  assign \new_[17215]_  = ~\new_[17668]_  & (~\new_[10484]_  | ~\new_[15941]_ );
  assign \new_[17216]_  = ~\new_[17738]_  & (~\new_[10407]_  | ~\new_[16107]_ );
  assign \new_[17217]_  = ~\new_[17581]_  & (~\new_[16853]_  | ~n17435);
  assign \new_[17218]_  = ~\new_[17543]_  & (~\new_[10408]_  | ~\new_[16443]_ );
  assign \new_[17219]_  = ~\new_[17735]_  & (~\new_[10356]_  | ~\new_[15985]_ );
  assign \new_[17220]_  = \new_[17863]_  ^ \new_[6312]_ ;
  assign \new_[17221]_  = \new_[12548]_  ^ \new_[17868]_ ;
  assign \new_[17222]_  = \new_[18357]_  ^ \new_[6326]_ ;
  assign \new_[17223]_  = ~\new_[17527]_  & (~\new_[13774]_  | ~\new_[16867]_ );
  assign \new_[17224]_  = ~\new_[17774]_  & (~\new_[13799]_  | ~\new_[16876]_ );
  assign \new_[17225]_  = ~\new_[17685]_  & (~\new_[10405]_  | ~\new_[16127]_ );
  assign \new_[17226]_  = ~\new_[17606]_  & (~\new_[16866]_  | ~n17450);
  assign \new_[17227]_  = ~\new_[17517]_  & (~\new_[10395]_  | ~\new_[16032]_ );
  assign \new_[17228]_  = ~\new_[17765]_  & (~\new_[8396]_  | ~\new_[16866]_ );
  assign \new_[17229]_  = \new_[17844]_  ^ \new_[6322]_ ;
  assign \new_[17230]_  = ~\new_[17553]_  & (~\new_[16867]_  | ~n17355);
  assign \new_[17231]_  = ~\new_[17652]_  & (~\new_[17072]_  | ~\new_[9639]_ );
  assign \new_[17232]_  = ~\new_[17513]_  & (~\new_[16876]_  | ~n17395);
  assign \new_[17233]_  = \new_[17045]_  ^ \new_[19070]_ ;
  assign \new_[17234]_  = \new_[17816]_  ^ \new_[6307]_ ;
  assign \new_[17235]_  = \new_[19614]_  ^ \new_[6553]_ ;
  assign \new_[17236]_  = \new_[19563]_  ^ \new_[6305]_ ;
  assign \new_[17237]_  = \new_[19296]_  ^ \new_[6554]_ ;
  assign \new_[17238]_  = ~\new_[17736]_  & (~\new_[10404]_  | ~\new_[16369]_ );
  assign \new_[17239]_  = ~\new_[17482]_  & (~\new_[10406]_  | ~\new_[16440]_ );
  assign \new_[17240]_  = \new_[19604]_  ^ \new_[6324]_ ;
  assign \new_[17241]_  = ~\new_[17293]_ ;
  assign n16670 = configuration_sync_isr_2_sync_bckp_bit_reg;
  assign \new_[17243]_  = \new_[17826]_  ^ \new_[19272]_ ;
  assign \new_[17244]_  = \new_[18085]_  ^ \new_[18084]_ ;
  assign n16520 = wishbone_slave_unit_del_sync_req_rty_exp_reg_reg;
  assign n16665 = configuration_sync_pci_err_cs_8_sync_bckp_bit_reg;
  assign \new_[17247]_  = ~\new_[17319]_ ;
  assign n16680 = \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[1] ;
  assign \new_[17249]_  = ~\new_[4092]_  | ~n16775;
  assign \new_[17250]_  = ~\new_[20521]_  | ~\new_[17544]_ ;
  assign \new_[17251]_  = ~\new_[20127]_  | ~\new_[20159]_ ;
  assign \new_[17252]_  = ~\new_[17303]_ ;
  assign \new_[17253]_  = ~\new_[17794]_  & ~\new_[19140]_ ;
  assign \new_[17254]_  = ~n16575;
  assign \new_[17255]_  = ~\new_[17296]_ ;
  assign \new_[17256]_  = ~\new_[10876]_  | ~\new_[11344]_ ;
  assign \new_[17257]_  = ~\new_[8385]_  | ~\new_[8386]_ ;
  assign \new_[17258]_  = ~\new_[20340]_ ;
  assign \new_[17259]_  = ~\new_[9792]_  & ~\new_[9764]_ ;
  assign \new_[17260]_  = ~\new_[10008]_  & ~\new_[10004]_ ;
  assign \new_[17261]_  = ~n17220 & ~n16995;
  assign \new_[17262]_  = \new_[13490]_  & \new_[13598]_ ;
  assign \new_[17263]_  = ~\new_[17460]_ ;
  assign \new_[17264]_  = ~\new_[3995]_  & ~\new_[10853]_ ;
  assign \new_[17265]_  = ~\new_[17636]_  & ~\new_[17802]_ ;
  assign \new_[17266]_  = ~wbs_err_o & ~wbs_rty_o;
  assign \new_[17267]_  = ~n16690 & ~\new_[15424]_ ;
  assign \new_[17268]_  = ~\new_[8548]_  & ~\new_[8224]_ ;
  assign \new_[17269]_  = ~\new_[10853]_  | ~\new_[4009]_ ;
  assign \new_[17270]_  = ~\new_[17472]_ ;
  assign \new_[17271]_  = ~\new_[17654]_  & ~\new_[13598]_ ;
  assign \new_[17272]_  = ~\new_[20479]_  & ~wbs_ack_o;
  assign \new_[17273]_  = ~\new_[17632]_  & ~\new_[11330]_ ;
  assign \new_[17274]_  = \new_[17681]_  | \wbs_adr_i[4] ;
  assign \new_[17275]_  = \new_[18116]_  ^ \new_[6321]_ ;
  assign \new_[17276]_  = ~\new_[17768]_  & ~\new_[17713]_ ;
  assign \new_[17277]_  = \new_[17841]_  ^ \new_[6551]_ ;
  assign \new_[17278]_  = \new_[17810]_  ^ \new_[6317]_ ;
  assign \new_[17279]_  = ~\new_[18928]_ ;
  assign \new_[17280]_  = \new_[19578]_  ^ \new_[6329]_ ;
  assign \new_[17281]_  = \new_[9565]_  & \new_[9627]_ ;
  assign \new_[17282]_  = \new_[9565]_  ^ \new_[9627]_ ;
  assign \new_[17283]_  = \wbm_adr_o[2]  & \wbm_adr_o[3] ;
  assign \new_[17284]_  = \wbm_adr_o[2]  ^ \wbm_adr_o[3] ;
  assign \new_[17285]_  = \new_[6321]_  & \new_[6554]_ ;
  assign \new_[17286]_  = \new_[6321]_  ^ \new_[6554]_ ;
  assign n16720 = ~\new_[19762]_  & ~\new_[17115]_ ;
  assign \new_[17288]_  = \new_[15210]_  ^ \new_[16144]_ ;
  assign n16815 = ~\new_[13150]_  & ~n17085;
  assign \new_[17290]_  = \new_[15406]_  ^ \new_[15924]_ ;
  assign \new_[17291]_  = ~\new_[17588]_ ;
  assign \new_[17292]_  = ~\new_[17568]_ ;
  assign \new_[17293]_  = \new_[10371]_  ? \new_[5047]_  : \new_[10371]_ ;
  assign \new_[17294]_  = \new_[15268]_  ^ \new_[16440]_ ;
  assign n16795 = ~\new_[19583]_  & ~n16715;
  assign \new_[17296]_  = \new_[18810]_  & \new_[13598]_ ;
  assign n16575 = \new_[13688]_  & \new_[19343]_ ;
  assign \new_[17298]_  = \new_[15231]_  ^ \new_[16354]_ ;
  assign \new_[17299]_  = ~\new_[19857]_  & ~\new_[8394]_ ;
  assign \new_[17300]_  = \new_[11344]_  & \new_[18910]_ ;
  assign \new_[17301]_  = \new_[15309]_  ^ \new_[15985]_ ;
  assign \new_[17302]_  = \new_[9675]_  ^ \new_[13763]_ ;
  assign \new_[17303]_  = ~\new_[18098]_  & ~\new_[13771]_ ;
  assign \new_[17304]_  = \new_[19136]_  & \new_[5046]_ ;
  assign \new_[17305]_  = ~\new_[20184]_ ;
  assign \new_[17306]_  = ~\new_[9799]_  & ~\new_[19224]_ ;
  assign \new_[17307]_  = \new_[9673]_  ^ \new_[13794]_ ;
  assign \new_[17308]_  = ~\new_[4008]_  | ~\new_[19012]_ ;
  assign \new_[17309]_  = \new_[15387]_  ^ \new_[16414]_ ;
  assign \new_[17310]_  = ~\new_[15594]_  & ~\new_[19011]_ ;
  assign \new_[17311]_  = ~\new_[18523]_  | ~wbm_err_i;
  assign \new_[17312]_  = ~\new_[12005]_  | ~\new_[9903]_ ;
  assign \new_[17313]_  = ~\new_[19567]_  & ~\new_[10004]_ ;
  assign \new_[17314]_  = \new_[15163]_  ^ \new_[16210]_ ;
  assign n16735 = \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg[1] ;
  assign n16805 = \\wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[2] ;
  assign \new_[17317]_  = \new_[15400]_  ^ \new_[16100]_ ;
  assign \new_[17318]_  = ~\new_[20101]_ ;
  assign \new_[17319]_  = ~pci_target_unit_wishbone_master_burst_chopped_delayed_reg;
  assign n16810 = \\wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[1] ;
  assign n16760 = \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[2] ;
  assign n16730 = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[1] ;
  assign \new_[17323]_  = ~\new_[17793]_ ;
  assign \new_[17324]_  = \new_[19567]_  & \new_[10004]_ ;
  assign n16780 = \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg[2] ;
  assign n16840 = \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[1] ;
  assign n16820 = \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[3] ;
  assign n16785 = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[3] ;
  assign n16850 = \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[1] ;
  assign n16830 = \\pci_target_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[1] ;
  assign n16765 = \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg[0] ;
  assign n16705 = \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[0] ;
  assign n16825 = \\pci_target_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[0] ;
  assign \new_[17334]_  = ~\new_[18615]_  | ~\new_[20520]_ ;
  assign n16845 = ~\new_[11325]_  & ~n16920;
  assign n16700 = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[2] ;
  assign n16835 = \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[2] ;
  assign n16790 = \\configuration_sync_pci_err_cs_8_delete_sync_sync_data_out_reg[0] ;
  assign \new_[17339]_  = \new_[16027]_  ^ \new_[16435]_ ;
  assign \new_[17340]_  = \new_[16440]_  ^ \new_[16369]_ ;
  assign \new_[17341]_  = \new_[19857]_  & \new_[8394]_ ;
  assign \new_[17342]_  = \new_[4178]_  ^ \new_[9902]_ ;
  assign \new_[17343]_  = \new_[16107]_  ^ \new_[15941]_ ;
  assign \new_[17344]_  = \new_[17878]_  & \new_[9621]_ ;
  assign \new_[17345]_  = \new_[16130]_  ^ \new_[16382]_ ;
  assign \new_[17346]_  = \new_[15989]_  ^ \new_[15985]_ ;
  assign \new_[17347]_  = \new_[4228]_  ^ \new_[4226]_ ;
  assign \new_[17348]_  = ~\new_[17819]_  & ~\new_[15399]_ ;
  assign \new_[17349]_  = \new_[4180]_  ^ \new_[4211]_ ;
  assign \new_[17350]_  = \new_[9641]_  ^ \new_[9628]_ ;
  assign \new_[17351]_  = \new_[13687]_  ^ \new_[16879]_ ;
  assign \new_[17352]_  = \new_[4185]_  ^ \new_[4184]_ ;
  assign \new_[17353]_  = \new_[4456]_  ^ \new_[4182]_ ;
  assign \new_[17354]_  = ~\new_[19194]_  & ~\new_[19410]_ ;
  assign \new_[17355]_  = \new_[16405]_  ^ \new_[15948]_ ;
  assign \new_[17356]_  = \new_[16414]_  ^ \new_[16013]_ ;
  assign \new_[17357]_  = \new_[5008]_  ^ \new_[5041]_ ;
  assign \new_[17358]_  = ~\new_[18825]_  & ~\new_[15399]_ ;
  assign \new_[17359]_  = ~\new_[17628]_ ;
  assign \new_[17360]_  = \new_[17043]_  ^ \new_[10012]_ ;
  assign \new_[17361]_  = \new_[15300]_  ^ \new_[15989]_ ;
  assign \new_[17362]_  = \new_[16100]_  ^ \new_[15927]_ ;
  assign \new_[17363]_  = \new_[9628]_  ^ \new_[9678]_ ;
  assign \new_[17364]_  = \new_[13685]_  ^ \new_[16879]_ ;
  assign \new_[17365]_  = \new_[19201]_  & \new_[12039]_ ;
  assign \new_[17366]_  = \new_[4210]_  ^ \new_[4229]_ ;
  assign \new_[17367]_  = ~\new_[17873]_  & ~\new_[8224]_ ;
  assign \new_[17368]_  = ~\new_[11345]_  & ~\new_[18123]_ ;
  assign \new_[17369]_  = \new_[4213]_  ^ \new_[4212]_ ;
  assign \new_[17370]_  = ~\new_[11345]_  | ~\new_[18123]_ ;
  assign \new_[17371]_  = \new_[15192]_  ^ \new_[16013]_ ;
  assign \new_[17372]_  = \new_[15188]_  ^ \new_[16130]_ ;
  assign wb_rst_o = ~\new_[18317]_  | ~pci_rst_i;
  assign \new_[17374]_  = ~\new_[13688]_  & (~n16935 | ~\new_[17115]_ );
  assign \new_[17375]_  = \new_[15190]_  ^ \new_[16134]_ ;
  assign n16710 = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[0] ;
  assign \new_[17377]_  = \new_[15233]_  ^ \new_[16150]_ ;
  assign \new_[17378]_  = \new_[15187]_  ^ \new_[15941]_ ;
  assign \new_[17379]_  = \new_[15329]_  ^ \new_[15948]_ ;
  assign \new_[17380]_  = \pci_cbe_i[2]  ? \new_[11095]_  : \new_[4178]_ ;
  assign \new_[17381]_  = \new_[15189]_  ^ \new_[15927]_ ;
  assign \new_[17382]_  = ~\new_[15181]_  & (~\new_[9765]_  | ~\new_[15182]_ );
  assign \new_[17383]_  = ~\new_[15216]_ ;
  assign \new_[17384]_  = ~\new_[17795]_ ;
  assign \new_[17385]_  = ~\new_[17748]_ ;
  assign \new_[17386]_  = \new_[15201]_  ^ \new_[16443]_ ;
  assign \new_[17387]_  = \new_[15186]_  ^ \new_[16107]_ ;
  assign \new_[17388]_  = \new_[15183]_  ^ \new_[16384]_ ;
  assign \new_[17389]_  = \new_[15232]_  ^ \new_[16032]_ ;
  assign \new_[17390]_  = \new_[15185]_  ^ \new_[16143]_ ;
  assign \new_[17391]_  = \new_[15170]_  ^ \new_[15926]_ ;
  assign \new_[17392]_  = \new_[15402]_  ^ \new_[15928]_ ;
  assign \new_[17393]_  = \new_[15401]_  ^ \new_[16369]_ ;
  assign \new_[17394]_  = \new_[15161]_  ^ \new_[16382]_ ;
  assign \new_[17395]_  = \new_[15194]_  ^ \new_[15923]_ ;
  assign \new_[17396]_  = \new_[15236]_  ^ \new_[16405]_ ;
  assign \new_[17397]_  = \new_[15204]_  ^ \new_[16027]_ ;
  assign \new_[17398]_  = \new_[15270]_  ^ \new_[16127]_ ;
  assign \new_[17399]_  = \new_[15284]_  ^ \new_[16435]_ ;
  assign \new_[17400]_  = \new_[9679]_  ^ \new_[13809]_ ;
  assign \new_[17401]_  = \new_[15285]_  ^ \new_[15986]_ ;
  assign \new_[17402]_  = \new_[9674]_  ^ \new_[13802]_ ;
  assign \new_[17403]_  = \pci_cbe_i[0]  ? \new_[11095]_  : \new_[4174]_ ;
  assign \new_[17404]_  = \pci_cbe_i[1]  ? \new_[11095]_  : \new_[9902]_ ;
  assign \new_[17405]_  = \pci_cbe_i[3]  ? \new_[11095]_  : \new_[4175]_ ;
  assign \new_[17406]_  = \new_[16443]_  ^ \new_[16143]_ ;
  assign \new_[17407]_  = \new_[4181]_  ^ \new_[4217]_ ;
  assign \new_[17408]_  = \new_[4130]_  ^ \new_[4261]_ ;
  assign \new_[17409]_  = \new_[17076]_  ^ \new_[10006]_ ;
  assign \new_[17410]_  = \new_[4183]_  ^ \new_[4268]_ ;
  assign \new_[17411]_  = \new_[13672]_  ^ \new_[16879]_ ;
  assign \new_[17412]_  = \new_[17143]_  ^ \new_[10077]_ ;
  assign \new_[17413]_  = \new_[16127]_  ^ \new_[16032]_ ;
  assign \new_[17414]_  = \new_[9616]_  ^ \new_[9678]_ ;
  assign \new_[17415]_  = \new_[16210]_  ^ \new_[16134]_ ;
  assign \new_[17416]_  = \new_[15923]_  ^ \new_[16150]_ ;
  assign \new_[17417]_  = \new_[16879]_  ^ n17165;
  assign \new_[17418]_  = \new_[4189]_  ^ \new_[4188]_ ;
  assign \new_[17419]_  = \new_[15924]_  ^ \new_[15926]_ ;
  assign \new_[17420]_  = \new_[15925]_  ^ \new_[16144]_ ;
  assign \new_[17421]_  = \new_[4218]_  ^ \new_[4192]_ ;
  assign \new_[17422]_  = \new_[10411]_  ^ \new_[16100]_ ;
  assign \new_[17423]_  = \new_[16354]_  ^ \new_[15928]_ ;
  assign \new_[17424]_  = \new_[13218]_  ^ \new_[16876]_ ;
  assign \new_[17425]_  = \new_[4187]_  ^ \new_[4186]_ ;
  assign \new_[17426]_  = \new_[4191]_  ^ \new_[4190]_ ;
  assign \new_[17427]_  = \new_[4260]_  ^ \new_[4345]_ ;
  assign \new_[17428]_  = \new_[4265]_  ^ \new_[4216]_ ;
  assign \new_[17429]_  = \new_[15986]_  ^ \new_[16384]_ ;
  assign \new_[17430]_  = \new_[4215]_  ^ \new_[4214]_ ;
  assign \new_[17431]_  = \new_[8203]_  ^ \new_[8202]_ ;
  assign n16855 = \\wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[0] ;
  assign \new_[17433]_  = ~\new_[11344]_  & ~\new_[18910]_ ;
  assign \new_[17434]_  = ~\new_[18098]_  | ~\new_[13771]_ ;
  assign \new_[17435]_  = ~\new_[18810]_  & ~\new_[13598]_ ;
  assign \new_[17436]_  = \new_[17873]_  & \new_[8224]_ ;
  assign \new_[17437]_  = ~\new_[9677]_  | ~\new_[19224]_ ;
  assign \new_[17438]_  = ~\new_[17484]_ ;
  assign \new_[17439]_  = ~\new_[9268]_  & ~\new_[19273]_ ;
  assign \new_[17440]_  = ~\new_[17492]_ ;
  assign \new_[17441]_  = ~\new_[19781]_  | ~\new_[9287]_ ;
  assign \new_[17442]_  = ~\new_[4459]_  | ~\new_[19077]_ ;
  assign \new_[17443]_  = ~\new_[8688]_  | ~\new_[19273]_ ;
  assign \new_[17444]_  = ~\new_[17490]_ ;
  assign \new_[17445]_  = ~\new_[17632]_ ;
  assign \new_[17446]_  = ~\new_[17715]_ ;
  assign \new_[17447]_  = n16890 | n17365;
  assign \new_[17448]_  = ~\new_[17959]_  | ~\new_[9880]_ ;
  assign \new_[17449]_  = ~\new_[18056]_  | ~\new_[9488]_ ;
  assign \new_[17450]_  = ~\new_[20490]_  | ~\new_[19393]_ ;
  assign \new_[17451]_  = ~\new_[17763]_ ;
  assign \new_[17452]_  = ~\new_[17579]_ ;
  assign \new_[17453]_  = ~\new_[17580]_ ;
  assign \new_[17454]_  = \new_[18392]_  & \new_[18928]_ ;
  assign \new_[17455]_  = ~\new_[10534]_  & ~\new_[18968]_ ;
  assign \new_[17456]_  = ~\new_[9879]_  | ~\new_[17959]_ ;
  assign \new_[17457]_  = ~\new_[17740]_ ;
  assign n16800 = ~\new_[17565]_ ;
  assign \new_[17459]_  = ~\new_[17727]_ ;
  assign \new_[17460]_  = ~\new_[20521]_  | ~\new_[19192]_ ;
  assign \new_[17461]_  = ~\new_[17709]_ ;
  assign \new_[17462]_  = ~\new_[17679]_ ;
  assign \new_[17463]_  = \new_[18190]_  | \new_[18515]_ ;
  assign \new_[17464]_  = ~\new_[6319]_  | ~\new_[18545]_ ;
  assign \new_[17465]_  = ~\new_[17649]_ ;
  assign \new_[17466]_  = ~\new_[17635]_ ;
  assign \new_[17467]_  = \new_[19201]_  & \new_[16852]_ ;
  assign \new_[17468]_  = ~\new_[8386]_  & ~\new_[8387]_ ;
  assign \new_[17469]_  = ~\new_[17675]_ ;
  assign \new_[17470]_  = ~\new_[19683]_  | ~\new_[20188]_ ;
  assign \new_[17471]_  = ~\new_[17670]_ ;
  assign \new_[17472]_  = ~\new_[18189]_  | ~\new_[18256]_ ;
  assign \new_[17473]_  = ~wbs_ack_o;
  assign \new_[17474]_  = ~\new_[20300]_ ;
  assign \new_[17475]_  = ~wbs_err_o;
  assign \new_[17476]_  = ~\new_[20143]_ ;
  assign n17100 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[18] ;
  assign \new_[17478]_  = ~\new_[10515]_  | ~\new_[15948]_ ;
  assign \new_[17479]_  = ~\new_[10402]_  & ~\new_[16134]_ ;
  assign \new_[17480]_  = ~\new_[10523]_  | ~\new_[16382]_ ;
  assign \new_[17481]_  = \new_[10773]_  & \new_[10846]_ ;
  assign \new_[17482]_  = ~\new_[10406]_  & ~\new_[16440]_ ;
  assign \new_[17483]_  = \new_[10394]_  | \new_[10396]_ ;
  assign \new_[17484]_  = ~\new_[5041]_  | ~\new_[5008]_ ;
  assign \new_[17485]_  = \new_[10510]_  & \new_[10518]_ ;
  assign \new_[17486]_  = \new_[15038]_  & \new_[14990]_ ;
  assign \new_[17487]_  = ~\new_[13761]_  & ~\new_[16867]_ ;
  assign \new_[17488]_  = \new_[9795]_  & \new_[9808]_ ;
  assign \new_[17489]_  = \new_[4962]_  & \new_[4975]_ ;
  assign \new_[17490]_  = \wbm_adr_o[5]  & \wbm_adr_o[6] ;
  assign \new_[17491]_  = \new_[10506]_  & \new_[10527]_ ;
  assign \new_[17492]_  = \new_[9794]_  & \new_[9790]_ ;
  assign \new_[17493]_  = ~\new_[6551]_  | ~\new_[6325]_ ;
  assign \new_[17494]_  = ~\wbm_adr_o[22]  | ~\wbm_adr_o[23] ;
  assign \new_[17495]_  = \new_[9644]_  & \new_[9623]_ ;
  assign n17105 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[31] ;
  assign n17110 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[3] ;
  assign n17115 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[4] ;
  assign n17120 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[25] ;
  assign n17125 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[6] ;
  assign n17130 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[16] ;
  assign n17135 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[11] ;
  assign n17140 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[2] ;
  assign \new_[17504]_  = \new_[10774]_  & \new_[10847]_ ;
  assign \new_[17505]_  = ~n17500 & ~n17350;
  assign \new_[17506]_  = ~\new_[10403]_  & ~\new_[16130]_ ;
  assign \new_[17507]_  = ~\wbm_adr_o[11]  | ~\wbm_adr_o[12] ;
  assign \new_[17508]_  = ~\new_[6553]_  | ~\new_[6322]_ ;
  assign \new_[17509]_  = ~\new_[9287]_ ;
  assign \new_[17510]_  = ~\new_[19904]_ ;
  assign n17145 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[1] ;
  assign \new_[17512]_  = ~\wbm_adr_o[9]  | ~\wbm_adr_o[10] ;
  assign \new_[17513]_  = ~\new_[16876]_  & ~n17395;
  assign \new_[17514]_  = ~\new_[10521]_  | ~\new_[16134]_ ;
  assign \new_[17515]_  = ~\new_[20225]_ ;
  assign \new_[17516]_  = ~\new_[4963]_  | ~\new_[5039]_ ;
  assign \new_[17517]_  = ~\new_[10395]_  & ~\new_[16032]_ ;
  assign \new_[17518]_  = ~\new_[10522]_  | ~\new_[16032]_ ;
  assign \new_[17519]_  = \new_[10046]_  & \new_[16179]_ ;
  assign \new_[17520]_  = \new_[10759]_  | \new_[10824]_ ;
  assign \new_[17521]_  = \new_[4977]_  & \new_[5043]_ ;
  assign \new_[17522]_  = ~\wbm_adr_o[19]  | ~\wbm_adr_o[20] ;
  assign \new_[17523]_  = ~\new_[10412]_  & ~\new_[10534]_ ;
  assign \new_[17524]_  = ~\new_[6323]_  | ~\new_[6324]_ ;
  assign \new_[17525]_  = \new_[10816]_  & \new_[10493]_ ;
  assign \new_[17526]_  = ~\new_[16893]_  & ~n17250;
  assign \new_[17527]_  = ~\new_[13774]_  & ~\new_[16867]_ ;
  assign \new_[17528]_  = ~\new_[8395]_  & ~\new_[16853]_ ;
  assign \new_[17529]_  = ~\new_[20224]_ ;
  assign \new_[17530]_  = \new_[10500]_  & \new_[10521]_ ;
  assign \new_[17531]_  = ~\wbm_adr_o[4]  | ~\wbm_adr_o[5] ;
  assign \new_[17532]_  = ~\new_[6305]_  | ~\new_[6306]_ ;
  assign \new_[17533]_  = \new_[6316]_  & \new_[6552]_ ;
  assign n17150 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[15] ;
  assign \new_[17535]_  = ~\new_[10399]_  & ~\new_[15924]_ ;
  assign \new_[17536]_  = ~\new_[9282]_  & ~\new_[9679]_ ;
  assign \new_[17537]_  = ~\new_[6317]_  | ~\new_[6303]_ ;
  assign n17155 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[14] ;
  assign \new_[17539]_  = ~\new_[6304]_  | ~\new_[6325]_ ;
  assign \new_[17540]_  = ~\new_[9622]_  | ~\new_[9644]_ ;
  assign \new_[17541]_  = \new_[10498]_  & \new_[10519]_ ;
  assign \new_[17542]_  = \new_[10501]_  & \new_[10514]_ ;
  assign \new_[17543]_  = ~\new_[10408]_  & ~\new_[16443]_ ;
  assign \new_[17544]_  = ~\new_[19192]_ ;
  assign \new_[17545]_  = ~\new_[10481]_  & ~\new_[16144]_ ;
  assign \new_[17546]_  = ~\new_[13221]_  & ~\new_[13134]_ ;
  assign \new_[17547]_  = ~\new_[10518]_  | ~\new_[15989]_ ;
  assign \new_[17548]_  = \new_[5039]_  & \new_[4964]_ ;
  assign \new_[17549]_  = ~\new_[15015]_  & ~\new_[9884]_ ;
  assign \new_[17550]_  = ~\new_[4968]_  | ~\new_[4967]_ ;
  assign \new_[17551]_  = ~\wbm_adr_o[18]  | ~\wbm_adr_o[19] ;
  assign n16860 = \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg[0] ;
  assign \new_[17553]_  = ~\new_[16867]_  & ~n17355;
  assign \new_[17554]_  = ~\new_[10848]_  | ~\new_[16443]_ ;
  assign \new_[17555]_  = ~\wbs_bte_i[0]  | ~\wbs_bte_i[1] ;
  assign \new_[17556]_  = ~\wbm_adr_o[13]  | ~\wbm_adr_o[14] ;
  assign \new_[17557]_  = \new_[11344]_  & \new_[11343]_ ;
  assign \new_[17558]_  = ~\new_[19923]_ ;
  assign n16915 = \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[2] ;
  assign \new_[17560]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[13] ;
  assign \new_[17561]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[11] ;
  assign \new_[17562]_  = ~\new_[6322]_  | ~\new_[6323]_ ;
  assign \new_[17563]_  = \new_[10505]_  & \new_[10848]_ ;
  assign \new_[17564]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[10] ;
  assign \new_[17565]_  = ~wb_int_i | ~\new_[10062]_ ;
  assign \new_[17566]_  = ~\new_[17087]_  & ~\new_[9636]_ ;
  assign \new_[17567]_  = ~\new_[3995]_  | ~\new_[10853]_ ;
  assign \new_[17568]_  = ~\new_[15399]_  | ~\new_[15361]_ ;
  assign \new_[17569]_  = ~\new_[10846]_  | ~\new_[16435]_ ;
  assign \new_[17570]_  = \new_[10508]_  & \new_[10515]_ ;
  assign \new_[17571]_  = \new_[5041]_  & \new_[4974]_ ;
  assign \new_[17572]_  = ~\new_[6329]_  | ~\new_[6307]_ ;
  assign \new_[17573]_  = \new_[4970]_  & \new_[4971]_ ;
  assign \new_[17574]_  = ~\new_[6326]_  | ~\new_[6316]_ ;
  assign \new_[17575]_  = \new_[10528]_  & \new_[16144]_ ;
  assign \new_[17576]_  = ~wbm_ack_i;
  assign \new_[17577]_  = ~\new_[11282]_  & ~\new_[11327]_ ;
  assign \new_[17578]_  = ~\new_[9907]_  | ~\new_[10063]_ ;
  assign \new_[17579]_  = ~\new_[13612]_  & ~\new_[13221]_ ;
  assign \new_[17580]_  = ~\new_[5045]_  | ~\new_[5046]_ ;
  assign \new_[17581]_  = ~\new_[16853]_  & ~n17435;
  assign \new_[17582]_  = ~\new_[6329]_  | ~\new_[6310]_ ;
  assign \new_[17583]_  = ~\new_[20105]_ ;
  assign \new_[17584]_  = ~\new_[10526]_  | ~\new_[16440]_ ;
  assign \new_[17585]_  = ~\wbm_adr_o[14]  | ~\wbm_adr_o[15] ;
  assign n16940 = \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg[2] ;
  assign \new_[17587]_  = \new_[8548]_  & \new_[8224]_ ;
  assign \new_[17588]_  = \new_[15114]_  & \new_[15123]_ ;
  assign \new_[17589]_  = ~\new_[20405]_ ;
  assign \new_[17590]_  = ~\new_[16130]_  | ~\new_[10524]_ ;
  assign \new_[17591]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[15] ;
  assign \new_[17592]_  = ~\new_[19922]_ ;
  assign \new_[17593]_  = ~\new_[10401]_  & ~\new_[15926]_ ;
  assign \new_[17594]_  = \new_[10822]_  & \new_[10520]_ ;
  assign n17195 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[8] ;
  assign n17200 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[0] ;
  assign \new_[17597]_  = ~\wbm_adr_o[23]  | ~\wbm_adr_o[24] ;
  assign \new_[17598]_  = ~\new_[6553]_  | ~\new_[6321]_ ;
  assign \new_[17599]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[6] ;
  assign n17210 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[21] ;
  assign \new_[17601]_  = ~\new_[6304]_  | ~\new_[6303]_ ;
  assign \new_[17602]_  = ~\new_[15928]_  & ~\new_[16354]_ ;
  assign \new_[17603]_  = \new_[8226]_  & \new_[8394]_ ;
  assign \new_[17604]_  = ~\new_[16849]_  & ~n17285;
  assign \new_[17605]_  = ~\new_[8397]_  & ~\new_[16849]_ ;
  assign \new_[17606]_  = ~\new_[16866]_  & ~n17450;
  assign \new_[17607]_  = ~\new_[6309]_  | ~\new_[6308]_ ;
  assign \new_[17608]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[25] ;
  assign n16950 = \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[0] ;
  assign n16980 = \\configuration_sync_isr_2_clear_delete_sync_sync_data_out_reg[0] ;
  assign \new_[17611]_  = \new_[10502]_  & \new_[10524]_ ;
  assign \new_[17612]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[19] ;
  assign \new_[17613]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[30] ;
  assign n17240 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[27] ;
  assign n17245 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[29] ;
  assign n16880 = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[3] ;
  assign n17255 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[19] ;
  assign n17260 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[23] ;
  assign n17265 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[22] ;
  assign \new_[17620]_  = ~\new_[4966]_  | ~\new_[5009]_ ;
  assign n17270 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[28] ;
  assign \new_[17622]_  = ~\new_[10008]_  | ~\new_[10004]_ ;
  assign n17275 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[24] ;
  assign n16975 = \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[4] ;
  assign n16925 = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[2] ;
  assign n17290 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[5] ;
  assign \new_[17627]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[4] ;
  assign \new_[17628]_  = ~\new_[12448]_  & ~\new_[12011]_ ;
  assign n17300 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[13] ;
  assign \new_[17630]_  = ~\new_[10845]_  | ~\new_[16143]_ ;
  assign \new_[17631]_  = ~\new_[8398]_  & ~\new_[16893]_ ;
  assign \new_[17632]_  = \new_[12012]_  | \new_[11880]_ ;
  assign \new_[17633]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[8] ;
  assign n16875 = ~n16715;
  assign \new_[17635]_  = ~\new_[5043]_  | ~\new_[5090]_ ;
  assign \new_[17636]_  = ~\new_[19393]_ ;
  assign \new_[17637]_  = \new_[4974]_  & \new_[4976]_ ;
  assign \new_[17638]_  = ~\new_[5045]_  & ~\new_[5046]_ ;
  assign \new_[17639]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[16] ;
  assign \new_[17640]_  = ~\new_[19857]_ ;
  assign \new_[17641]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[17] ;
  assign \new_[17642]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[1] ;
  assign n16945 = configuration_rst_inactive_sync_reg;
  assign wbs_ack_o = ~\new_[19204]_ ;
  assign \new_[17645]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[26] ;
  assign \new_[17646]_  = ~\new_[18928]_ ;
  assign n16960 = \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[5] ;
  assign \new_[17648]_  = ~configuration_sync_isr_2_delayed_del_bit_reg;
  assign \new_[17649]_  = ~\new_[13801]_  | ~\new_[14957]_ ;
  assign \new_[17650]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[22] ;
  assign n16955 = \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[2] ;
  assign \new_[17652]_  = ~\new_[17072]_  & ~\new_[9639]_ ;
  assign \new_[17653]_  = ~\new_[10370]_  | ~\new_[10372]_ ;
  assign \new_[17654]_  = ~\new_[18810]_ ;
  assign \new_[17655]_  = ~\new_[17046]_  & ~\new_[9635]_ ;
  assign \new_[17656]_  = ~\new_[19567]_ ;
  assign n16885 = \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[1] ;
  assign n16905 = \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg[1] ;
  assign \new_[17659]_  = ~\new_[6328]_  | ~\new_[6313]_ ;
  assign n16985 = \\wishbone_slave_unit_del_sync_rty_exp_sync_sync_data_out_reg[0] ;
  assign \new_[17661]_  = ~\new_[6328]_  | ~\new_[6312]_ ;
  assign \new_[17662]_  = \new_[5040]_  & \new_[5012]_ ;
  assign \new_[17663]_  = ~\new_[10525]_  | ~\new_[16107]_ ;
  assign \new_[17664]_  = ~\new_[8224]_  | ~\new_[8226]_ ;
  assign \new_[17665]_  = ~\new_[4963]_  | ~\new_[5090]_ ;
  assign \new_[17666]_  = ~\new_[4969]_  | ~\new_[5010]_ ;
  assign \new_[17667]_  = \new_[14911]_  & \new_[14989]_ ;
  assign \new_[17668]_  = ~\new_[10484]_  & ~\new_[15941]_ ;
  assign \new_[17669]_  = ~\new_[6309]_  | ~\new_[6329]_ ;
  assign \new_[17670]_  = ~\new_[6315]_  | ~\new_[6314]_ ;
  assign \new_[17671]_  = \new_[4976]_  & \new_[5042]_ ;
  assign \new_[17672]_  = ~\new_[10492]_  | ~\new_[16127]_ ;
  assign \new_[17673]_  = \new_[10530]_  & \new_[15927]_ ;
  assign \new_[17674]_  = ~\wbm_adr_o[8]  | ~\wbm_adr_o[9] ;
  assign \new_[17675]_  = ~\wbm_adr_o[25]  | ~\wbm_adr_o[26] ;
  assign \new_[17676]_  = ~\new_[10519]_  | ~\new_[16369]_ ;
  assign \new_[17677]_  = \new_[10495]_  & \new_[10492]_ ;
  assign \new_[17678]_  = \new_[9796]_  & \new_[9807]_ ;
  assign \new_[17679]_  = ~\new_[5010]_  | ~\new_[4896]_ ;
  assign \new_[17680]_  = \new_[10042]_  & \new_[9879]_ ;
  assign \new_[17681]_  = \wbs_adr_i[2]  | \wbs_adr_i[3] ;
  assign \new_[17682]_  = ~\new_[10847]_  | ~\new_[16027]_ ;
  assign \new_[17683]_  = ~\new_[10516]_  | ~\new_[15985]_ ;
  assign \new_[17684]_  = ~\wbm_adr_o[17]  | ~\wbm_adr_o[18] ;
  assign \new_[17685]_  = ~\new_[10405]_  & ~\new_[16127]_ ;
  assign \new_[17686]_  = \new_[10504]_  & \new_[10845]_ ;
  assign \new_[17687]_  = ~\new_[9282]_  & ~\new_[9673]_ ;
  assign \new_[17688]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[23] ;
  assign n17375 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[20] ;
  assign \new_[17690]_  = \new_[10744]_  & \new_[10528]_ ;
  assign \new_[17691]_  = ~\new_[10491]_  | ~\new_[15926]_ ;
  assign \new_[17692]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[12] ;
  assign n17385 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[12] ;
  assign \new_[17694]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[21] ;
  assign n16865 = \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[0] ;
  assign n17400 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[7] ;
  assign \new_[17697]_  = \new_[10494]_  & \new_[10517]_ ;
  assign \new_[17698]_  = ~\new_[9828]_  & ~\new_[9797]_ ;
  assign \new_[17699]_  = \wbm_adr_o[26]  & \wbm_adr_o[27] ;
  assign \new_[17700]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[20] ;
  assign n17410 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[26] ;
  assign \new_[17702]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[9] ;
  assign \new_[17703]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[24] ;
  assign \new_[17704]_  = ~\new_[6315]_  | ~\new_[6552]_ ;
  assign \new_[17705]_  = ~\new_[10520]_  | ~\new_[15924]_ ;
  assign \new_[17706]_  = ~\new_[6317]_  | ~\new_[6305]_ ;
  assign \new_[17707]_  = ~n16655;
  assign \new_[17708]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[7] ;
  assign \new_[17709]_  = ~\new_[4896]_  | ~\new_[4970]_ ;
  assign n16970 = \\configuration_command_bit_sync_sync_data_out_reg[0] ;
  assign n16870 = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[0] ;
  assign \new_[17712]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[14] ;
  assign \new_[17713]_  = ~\new_[5009]_  | ~\new_[4967]_ ;
  assign \new_[17714]_  = ~\wbm_adr_o[16]  | ~\wbm_adr_o[17] ;
  assign \new_[17715]_  = \new_[11344]_  | \new_[11343]_ ;
  assign \new_[17716]_  = \new_[10527]_  & \new_[16100]_ ;
  assign \new_[17717]_  = ~\new_[6551]_  | ~\new_[6324]_ ;
  assign \new_[17718]_  = \new_[10511]_  & \new_[10522]_ ;
  assign \new_[17719]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[31] ;
  assign n16900 = \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[1] ;
  assign \new_[17721]_  = ~\new_[11622]_  & ~\new_[11331]_ ;
  assign \new_[17722]_  = ~wbm_rty_i & ~wbm_err_i;
  assign \new_[17723]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[0] ;
  assign n17460 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[10] ;
  assign n16990 = \\configuration_sync_pci_err_cs_8_clear_delete_sync_sync_data_out_reg[0] ;
  assign \new_[17726]_  = ~\wbs_cti_i[0]  & ~\wbs_cti_i[2] ;
  assign \new_[17727]_  = ~\new_[4965]_  | ~\new_[4966]_ ;
  assign \new_[17728]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[3] ;
  assign \new_[17729]_  = ~\wbm_adr_o[6]  | ~\wbm_adr_o[7] ;
  assign \new_[17730]_  = ~\new_[6307]_  | ~\new_[6306]_ ;
  assign \new_[17731]_  = ~\new_[17052]_  & ~\new_[9637]_ ;
  assign \new_[17732]_  = ~\new_[6311]_  | ~\new_[6312]_ ;
  assign \new_[17733]_  = ~\wbm_adr_o[12]  | ~\wbm_adr_o[13] ;
  assign \new_[17734]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[18] ;
  assign \new_[17735]_  = ~\new_[10356]_  & ~\new_[15985]_ ;
  assign \new_[17736]_  = ~\new_[10404]_  & ~\new_[16369]_ ;
  assign \new_[17737]_  = \new_[10043]_  & \new_[9880]_ ;
  assign \new_[17738]_  = ~\new_[10407]_  & ~\new_[16107]_ ;
  assign \new_[17739]_  = \new_[10794]_  & \new_[10530]_ ;
  assign \new_[17740]_  = \new_[11345]_  | \new_[10876]_ ;
  assign \new_[17741]_  = \new_[13821]_  & \new_[13801]_ ;
  assign \new_[17742]_  = ~\wbm_adr_o[10]  | ~\wbm_adr_o[11] ;
  assign \new_[17743]_  = ~wishbone_slave_unit_del_sync_comp_done_reg_clr_reg;
  assign \new_[17744]_  = ~n17335 & ~n17280;
  assign wbs_err_o = ~\new_[19900]_ ;
  assign \new_[17746]_  = ~\new_[20296]_ ;
  assign \new_[17747]_  = ~\new_[18066]_ ;
  assign \new_[17748]_  = ~\new_[20301]_ ;
  assign \new_[17749]_  = ~\new_[20284]_ ;
  assign \new_[17750]_  = wbs_cyc_i & wbs_stb_i;
  assign \new_[17751]_  = ~\new_[10485]_  & ~\new_[16210]_ ;
  assign \new_[17752]_  = ~\new_[19905]_ ;
  assign \new_[17753]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[27] ;
  assign n16645 = ~n16655;
  assign \new_[17755]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[28] ;
  assign \new_[17756]_  = ~configuration_sync_pci_err_cs_8_delayed_del_bit_reg;
  assign n16965 = \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[3] ;
  assign \new_[17758]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[5] ;
  assign \new_[17759]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[29] ;
  assign \new_[17760]_  = \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[2] ;
  assign \new_[17761]_  = ~\new_[9282]_  & ~\new_[9675]_ ;
  assign \new_[17762]_  = \new_[15110]_  & \new_[14995]_ ;
  assign \new_[17763]_  = ~\wbm_adr_o[24]  | ~\wbm_adr_o[25] ;
  assign \new_[17764]_  = ~\new_[9282]_  & ~\new_[9674]_ ;
  assign \new_[17765]_  = ~\new_[8396]_  & ~\new_[16866]_ ;
  assign \new_[17766]_  = \new_[10503]_  & \new_[10525]_ ;
  assign \new_[17767]_  = ~\new_[4964]_  | ~\new_[5040]_ ;
  assign \new_[17768]_  = ~\new_[4968]_  | ~\new_[4969]_ ;
  assign \new_[17769]_  = \new_[10529]_  & \new_[15925]_ ;
  assign \new_[17770]_  = ~\new_[5042]_  | ~\new_[4977]_ ;
  assign \new_[17771]_  = \new_[11345]_  & \new_[10876]_ ;
  assign \new_[17772]_  = ~\new_[10517]_  | ~\new_[16405]_ ;
  assign \new_[17773]_  = ~\new_[6314]_  | ~\new_[6313]_ ;
  assign \new_[17774]_  = ~\new_[13799]_  & ~\new_[16876]_ ;
  assign \new_[17775]_  = ~\new_[13216]_  & ~\new_[16876]_ ;
  assign \new_[17776]_  = ~\new_[10483]_  & ~\new_[16143]_ ;
  assign \new_[17777]_  = ~\new_[8226]_  & ~\new_[8394]_ ;
  assign \new_[17778]_  = ~\wbm_adr_o[20]  | ~\wbm_adr_o[21] ;
  assign \new_[17779]_  = ~\new_[5044]_  | ~\new_[5038]_ ;
  assign \new_[17780]_  = ~\wbm_adr_o[7]  | ~\wbm_adr_o[8] ;
  assign \new_[17781]_  = \new_[10493]_  & \new_[15941]_ ;
  assign \new_[17782]_  = ~\new_[10409]_  & ~\new_[15927]_ ;
  assign \new_[17783]_  = \new_[10507]_  & \new_[10529]_ ;
  assign \new_[17784]_  = \new_[10775]_  & \new_[10523]_ ;
  assign \new_[17785]_  = ~\new_[6311]_  | ~\new_[6310]_ ;
  assign \new_[17786]_  = ~\new_[10486]_  & ~\new_[16382]_ ;
  assign \new_[17787]_  = ~\new_[10398]_  & ~\new_[15989]_ ;
  assign \new_[17788]_  = ~\new_[4965]_  | ~\new_[5012]_ ;
  assign \new_[17789]_  = \wbm_adr_o[27]  & \wbm_adr_o[28] ;
  assign n17520 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[17] ;
  assign \new_[17791]_  = ~\wbm_adr_o[21]  | ~\wbm_adr_o[22] ;
  assign \new_[17792]_  = ~\new_[13437]_  & ~\new_[16867]_ ;
  assign \new_[17793]_  = ~\new_[9903]_ ;
  assign \new_[17794]_  = ~\new_[20297]_ ;
  assign \new_[17795]_  = \new_[11691]_  | \new_[11882]_ ;
  assign n17525 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[9] ;
  assign \new_[17797]_  = \new_[9672]_  & \new_[12039]_ ;
  assign \new_[17798]_  = ~\new_[10514]_  | ~\new_[16210]_ ;
  assign \new_[17799]_  = \new_[10512]_  & \new_[10491]_ ;
  assign \new_[17800]_  = ~\new_[9562]_  | ~\new_[9621]_ ;
  assign \new_[17801]_  = ~\wbm_adr_o[15]  | ~\wbm_adr_o[16] ;
  assign \new_[17802]_  = ~\new_[18903]_ ;
  assign \new_[17803]_  = ~\new_[6308]_  | ~\new_[6305]_ ;
  assign n17530 = \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[30] ;
  assign \new_[17805]_  = ~\new_[8385]_  & ~\new_[8386]_ ;
  assign \new_[17806]_  = ~\new_[6701]_ ;
  assign \new_[17807]_  = ~\new_[6916]_ ;
  assign \new_[17808]_  = ~\new_[11456]_ ;
  assign \new_[17809]_  = ~\new_[11545]_ ;
  assign \new_[17810]_  = ~\new_[8689]_ ;
  assign \new_[17811]_  = ~\new_[12140]_ ;
  assign \new_[17812]_  = ~\new_[8688]_ ;
  assign \new_[17813]_  = ~\new_[6966]_ ;
  assign \new_[17814]_  = ~\new_[9771]_ ;
  assign \new_[17815]_  = ~\new_[7245]_ ;
  assign \new_[17816]_  = ~\new_[8208]_ ;
  assign \new_[17817]_  = ~\new_[13612]_ ;
  assign \new_[17818]_  = ~\new_[11336]_ ;
  assign \new_[17819]_  = ~\new_[15402]_ ;
  assign \new_[17820]_  = ~\new_[12272]_ ;
  assign \new_[17821]_  = ~\new_[8206]_ ;
  assign \new_[17822]_  = ~\new_[11091]_ ;
  assign \new_[17823]_  = ~\new_[6629]_ ;
  assign \new_[17824]_  = ~\new_[9779]_ ;
  assign \new_[17825]_  = ~\new_[5472]_ ;
  assign \new_[17826]_  = ~\new_[5110]_ ;
  assign \new_[17827]_  = ~\new_[11606]_ ;
  assign \new_[17828]_  = ~\new_[11548]_ ;
  assign \new_[17829]_  = ~\new_[12134]_ ;
  assign n17015 = ~\new_[9192]_ ;
  assign \new_[17831]_  = ~\new_[5413]_ ;
  assign \new_[17832]_  = ~\new_[7432]_ ;
  assign \new_[17833]_  = ~\new_[7499]_ ;
  assign \new_[17834]_  = ~\new_[6899]_ ;
  assign \new_[17835]_  = ~\new_[11572]_ ;
  assign \new_[17836]_  = ~\new_[11276]_ ;
  assign \new_[17837]_  = ~\new_[11465]_ ;
  assign \new_[17838]_  = ~\new_[10219]_ ;
  assign \new_[17839]_  = ~\new_[10335]_ ;
  assign \new_[17840]_  = ~\new_[5024]_ ;
  assign \new_[17841]_  = ~\new_[8222]_ ;
  assign \new_[17842]_  = ~\new_[11732]_ ;
  assign \new_[17843]_  = ~\new_[9671]_ ;
  assign \new_[17844]_  = ~\new_[8692]_ ;
  assign \new_[17845]_  = ~\new_[11463]_ ;
  assign \new_[17846]_  = ~\new_[11703]_ ;
  assign \new_[17847]_  = ~\new_[11539]_ ;
  assign \new_[17848]_  = ~\new_[6906]_ ;
  assign \new_[17849]_  = ~\new_[11666]_ ;
  assign \new_[17850]_  = ~\new_[6636]_ ;
  assign \new_[17851]_  = ~\new_[9672]_ ;
  assign \new_[17852]_  = ~\new_[7447]_ ;
  assign \new_[17853]_  = ~\new_[10274]_ ;
  assign \new_[17854]_  = ~\new_[8220]_ ;
  assign \new_[17855]_  = ~\new_[5476]_ ;
  assign \new_[17856]_  = ~\new_[11072]_ ;
  assign \new_[17857]_  = ~\new_[11576]_ ;
  assign \new_[17858]_  = ~\new_[9769]_ ;
  assign \new_[17859]_  = ~\new_[11484]_ ;
  assign \new_[17860]_  = ~\new_[9780]_ ;
  assign \new_[17861]_  = ~\new_[12236]_ ;
  assign \new_[17862]_  = ~\new_[12528]_ ;
  assign \new_[17863]_  = ~\new_[8274]_ ;
  assign \new_[17864]_  = ~\new_[6975]_ ;
  assign \new_[17865]_  = ~\new_[12379]_ ;
  assign \new_[17866]_  = ~\new_[5063]_ ;
  assign \new_[17867]_  = ~\new_[5023]_ ;
  assign \new_[17868]_  = ~\new_[12081]_ ;
  assign \new_[17869]_  = ~\new_[11434]_ ;
  assign \new_[17870]_  = ~\new_[11464]_ ;
  assign \new_[17871]_  = ~\new_[12529]_ ;
  assign \new_[17872]_  = ~\new_[12277]_ ;
  assign \new_[17873]_  = ~\new_[8548]_ ;
  assign \new_[17874]_  = ~\new_[11754]_ ;
  assign \new_[17875]_  = ~\new_[12478]_ ;
  assign \new_[17876]_  = ~\new_[8205]_ ;
  assign \new_[17877]_  = ~\new_[7229]_ ;
  assign \new_[17878]_  = ~\new_[9562]_ ;
  assign \new_[17879]_  = ~\new_[6951]_ ;
  assign \new_[17880]_  = ~\new_[5051]_ ;
  assign \new_[17881]_  = ~\new_[11698]_ ;
  assign \new_[17882]_  = ~\new_[5478]_ ;
  assign \new_[17883]_  = ~\new_[11660]_ ;
  assign \new_[17884]_  = ~\new_[9822]_ ;
  assign \new_[17885]_  = ~\new_[11265]_ ;
  assign \new_[17886]_  = ~\new_[6659]_ ;
  assign \new_[17887]_  = ~\new_[11116]_ ;
  assign \new_[17888]_  = ~\new_[6962]_ ;
  assign \new_[17889]_  = ~\new_[10259]_ ;
  assign \new_[17890]_  = ~\new_[11301]_ ;
  assign \new_[17891]_  = ~\new_[8209]_ ;
  assign \new_[17892]_  = ~\new_[10113]_ ;
  assign \new_[17893]_  = ~\new_[7459]_ ;
  assign \new_[17894]_  = ~\new_[9770]_ ;
  assign \new_[17895]_  = ~\new_[6947]_ ;
  assign \new_[17896]_  = ~\new_[10162]_ ;
  assign \new_[17897]_  = ~\new_[6726]_ ;
  assign \new_[17898]_  = ~\new_[11309]_ ;
  assign \new_[17899]_  = ~\new_[11478]_ ;
  assign \new_[17900]_  = ~\new_[10118]_ ;
  assign \new_[17901]_  = ~\new_[6872]_ ;
  assign \new_[17902]_  = ~\new_[11477]_ ;
  assign \new_[17903]_  = ~\new_[7704]_ ;
  assign \new_[17904]_  = ~\new_[6837]_ ;
  assign \new_[17905]_  = ~\new_[11306]_ ;
  assign \new_[17906]_  = ~\new_[11305]_ ;
  assign \new_[17907]_  = ~\new_[11853]_ ;
  assign \new_[17908]_  = ~\new_[10879]_ ;
  assign \new_[17909]_  = ~\new_[10122]_ ;
  assign \new_[17910]_  = ~\new_[6695]_ ;
  assign \new_[17911]_  = ~\new_[6967]_ ;
  assign \new_[17912]_  = ~\new_[10121]_ ;
  assign \new_[17913]_  = ~\new_[6780]_ ;
  assign \new_[17914]_  = ~\new_[6164]_ ;
  assign \new_[17915]_  = ~\new_[6777]_ ;
  assign \new_[17916]_  = ~\new_[6776]_ ;
  assign \new_[17917]_  = ~\new_[11399]_ ;
  assign \new_[17918]_  = ~\new_[7474]_ ;
  assign \new_[17919]_  = ~\new_[10095]_ ;
  assign \new_[17920]_  = ~\new_[11079]_ ;
  assign \new_[17921]_  = ~\new_[10938]_ ;
  assign \new_[17922]_  = ~\new_[6774]_ ;
  assign \new_[17923]_  = ~\new_[11549]_ ;
  assign \new_[17924]_  = ~\new_[10291]_ ;
  assign \new_[17925]_  = ~\new_[6592]_ ;
  assign \new_[17926]_  = ~\new_[6769]_ ;
  assign \new_[17927]_  = ~\new_[6767]_ ;
  assign \new_[17928]_  = ~\new_[7961]_ ;
  assign \new_[17929]_  = ~\new_[6766]_ ;
  assign \new_[17930]_  = ~\new_[6968]_ ;
  assign \new_[17931]_  = ~\new_[11480]_ ;
  assign \new_[17932]_  = ~\new_[11410]_ ;
  assign \new_[17933]_  = ~\new_[10054]_ ;
  assign \new_[17934]_  = ~\new_[10882]_ ;
  assign \new_[17935]_  = ~\new_[12154]_ ;
  assign \new_[17936]_  = ~\new_[12281]_ ;
  assign \new_[17937]_  = ~\new_[11559]_ ;
  assign \new_[17938]_  = ~\new_[11733]_ ;
  assign \new_[17939]_  = ~\new_[6792]_ ;
  assign \new_[17940]_  = ~\new_[11725]_ ;
  assign \new_[17941]_  = ~\new_[11721]_ ;
  assign \new_[17942]_  = ~\new_[6943]_ ;
  assign \new_[17943]_  = ~\new_[9230]_ ;
  assign \new_[17944]_  = ~\new_[7926]_ ;
  assign \new_[17945]_  = ~\new_[6717]_ ;
  assign \new_[17946]_  = ~\new_[10448]_ ;
  assign \new_[17947]_  = ~\new_[9283]_ ;
  assign \new_[17948]_  = ~\new_[11751]_ ;
  assign \new_[17949]_  = ~\new_[6791]_ ;
  assign \new_[17950]_  = ~\new_[12344]_ ;
  assign \new_[17951]_  = ~\new_[10934]_ ;
  assign \new_[17952]_  = ~\new_[6608]_ ;
  assign \new_[17953]_  = ~\new_[12245]_ ;
  assign \new_[17954]_  = ~\new_[12142]_ ;
  assign \new_[17955]_  = ~\new_[10139]_ ;
  assign \new_[17956]_  = ~\new_[6960]_ ;
  assign \new_[17957]_  = ~\new_[10853]_ ;
  assign \new_[17958]_  = ~\new_[9983]_ ;
  assign \new_[17959]_  = ~\new_[6320]_ ;
  assign \new_[17960]_  = ~\new_[11441]_ ;
  assign \new_[17961]_  = ~\new_[11770]_ ;
  assign \new_[17962]_  = ~\new_[6694]_ ;
  assign \new_[17963]_  = ~\new_[11765]_ ;
  assign \new_[17964]_  = ~\new_[10141]_ ;
  assign \new_[17965]_  = ~\new_[11750]_ ;
  assign \new_[17966]_  = ~\new_[11452]_ ;
  assign \new_[17967]_  = ~\new_[7450]_ ;
  assign \new_[17968]_  = ~\new_[11458]_ ;
  assign \new_[17969]_  = ~\new_[6589]_ ;
  assign \new_[17970]_  = ~\new_[11552]_ ;
  assign \new_[17971]_  = ~\new_[9617]_ ;
  assign \new_[17972]_  = ~\new_[12319]_ ;
  assign \new_[17973]_  = ~\new_[6853]_ ;
  assign \new_[17974]_  = ~\new_[11603]_ ;
  assign \new_[17975]_  = ~\new_[11611]_ ;
  assign \new_[17976]_  = ~\new_[6721]_ ;
  assign \new_[17977]_  = ~\new_[6722]_ ;
  assign \new_[17978]_  = ~\new_[10265]_ ;
  assign \new_[17979]_  = ~\new_[12274]_ ;
  assign \new_[17980]_  = ~\new_[6697]_ ;
  assign \new_[17981]_  = ~\new_[7486]_ ;
  assign \new_[17982]_  = ~\new_[6912]_ ;
  assign \new_[17983]_  = ~\new_[6819]_ ;
  assign \new_[17984]_  = ~\new_[9620]_ ;
  assign \new_[17985]_  = ~\new_[10165]_ ;
  assign \new_[17986]_  = ~\new_[11530]_ ;
  assign \new_[17987]_  = ~\new_[11881]_ ;
  assign \new_[17988]_  = ~\new_[11535]_ ;
  assign \new_[17989]_  = ~\new_[9640]_ ;
  assign \new_[17990]_  = ~\new_[6892]_ ;
  assign \new_[17991]_  = ~\new_[11134]_ ;
  assign \new_[17992]_  = ~\new_[6790]_ ;
  assign \new_[17993]_  = ~\new_[12271]_ ;
  assign \new_[17994]_  = ~\new_[10047]_ ;
  assign \new_[17995]_  = ~\new_[11816]_ ;
  assign \new_[17996]_  = ~\new_[11690]_ ;
  assign \new_[17997]_  = ~\new_[10149]_ ;
  assign \new_[17998]_  = ~\new_[10256]_ ;
  assign \new_[17999]_  = ~\new_[11592]_ ;
  assign \new_[18000]_  = ~\new_[11779]_ ;
  assign \new_[18001]_  = ~\new_[11105]_ ;
  assign \new_[18002]_  = ~\new_[5056]_ ;
  assign \new_[18003]_  = ~\new_[11581]_ ;
  assign \new_[18004]_  = ~\new_[6556]_ ;
  assign \new_[18005]_  = ~\new_[12242]_ ;
  assign \new_[18006]_  = ~\new_[11967]_ ;
  assign \new_[18007]_  = ~\new_[7476]_ ;
  assign \new_[18008]_  = ~\new_[11879]_ ;
  assign \new_[18009]_  = ~\new_[11665]_ ;
  assign \new_[18010]_  = ~\new_[11689]_ ;
  assign \new_[18011]_  = ~\new_[11634]_ ;
  assign \new_[18012]_  = ~\new_[11644]_ ;
  assign \new_[18013]_  = ~\new_[11649]_ ;
  assign \new_[18014]_  = ~\new_[6908]_ ;
  assign \new_[18015]_  = ~\new_[11566]_ ;
  assign \new_[18016]_  = ~\new_[11339]_ ;
  assign \new_[18017]_  = ~\new_[11337]_ ;
  assign \new_[18018]_  = ~\new_[6643]_ ;
  assign \new_[18019]_  = ~\new_[6789]_ ;
  assign \new_[18020]_  = ~\new_[8204]_ ;
  assign \new_[18021]_  = ~\new_[10157]_ ;
  assign \new_[18022]_  = ~\new_[7456]_ ;
  assign \new_[18023]_  = ~n16895;
  assign \new_[18024]_  = ~\new_[10161]_ ;
  assign \new_[18025]_  = ~\new_[11692]_ ;
  assign \new_[18026]_  = ~\new_[11704]_ ;
  assign \new_[18027]_  = ~\new_[8203]_ ;
  assign \new_[18028]_  = ~\new_[11686]_ ;
  assign \new_[18029]_  = ~\new_[6705]_ ;
  assign \new_[18030]_  = ~\new_[6724]_ ;
  assign \new_[18031]_  = ~\new_[9629]_ ;
  assign \new_[18032]_  = ~\new_[12094]_ ;
  assign \new_[18033]_  = ~\new_[11128]_ ;
  assign \new_[18034]_  = ~\new_[6890]_ ;
  assign \new_[18035]_  = ~\new_[9821]_ ;
  assign \new_[18036]_  = ~\new_[10231]_ ;
  assign \new_[18037]_  = ~\new_[5486]_ ;
  assign \new_[18038]_  = ~\new_[10266]_ ;
  assign \new_[18039]_  = ~\new_[11467]_ ;
  assign \new_[18040]_  = ~\new_[7288]_ ;
  assign \new_[18041]_  = ~\new_[9766]_ ;
  assign \new_[18042]_  = ~\new_[11609]_ ;
  assign \new_[18043]_  = ~\new_[11296]_ ;
  assign \new_[18044]_  = ~\new_[11295]_ ;
  assign \new_[18045]_  = ~\new_[11446]_ ;
  assign \new_[18046]_  = ~\new_[4979]_ ;
  assign \new_[18047]_  = ~\new_[8223]_ ;
  assign \new_[18048]_  = ~\new_[11491]_ ;
  assign \new_[18049]_  = ~\new_[11114]_ ;
  assign \new_[18050]_  = ~\new_[11789]_ ;
  assign \new_[18051]_  = ~\new_[12109]_ ;
  assign \new_[18052]_  = ~\new_[6759]_ ;
  assign \new_[18053]_  = ~\new_[12110]_ ;
  assign \new_[18054]_  = ~\new_[7455]_ ;
  assign \new_[18055]_  = ~\new_[10170]_ ;
  assign \new_[18056]_  = ~\new_[8681]_ ;
  assign \new_[18057]_  = ~\new_[7819]_ ;
  assign \new_[18058]_  = ~\new_[7453]_ ;
  assign \new_[18059]_  = ~\new_[11784]_ ;
  assign \new_[18060]_  = ~\new_[11492]_ ;
  assign \new_[18061]_  = ~\new_[10098]_ ;
  assign \new_[18062]_  = ~\new_[10172]_ ;
  assign \new_[18063]_  = ~\new_[9768]_ ;
  assign \new_[18064]_  = ~\new_[6848]_ ;
  assign n16775 = ~\new_[4084]_ ;
  assign \new_[18066]_  = ~\new_[10374]_ ;
  assign \new_[18067]_  = ~\new_[10169]_ ;
  assign \new_[18068]_  = ~\new_[11268]_ ;
  assign \new_[18069]_  = ~\new_[10343]_ ;
  assign \new_[18070]_  = ~\new_[6866]_ ;
  assign \new_[18071]_  = ~\new_[6742]_ ;
  assign \new_[18072]_  = ~\new_[7738]_ ;
  assign \new_[18073]_  = ~\new_[11117]_ ;
  assign \new_[18074]_  = ~\new_[12336]_ ;
  assign \new_[18075]_  = ~\new_[9824]_ ;
  assign \new_[18076]_  = ~\new_[10317]_ ;
  assign \new_[18077]_  = ~\new_[6846]_ ;
  assign \new_[18078]_  = ~\new_[11466]_ ;
  assign \new_[18079]_  = ~\new_[10175]_ ;
  assign \new_[18080]_  = ~\new_[5500]_ ;
  assign \new_[18081]_  = ~\new_[7783]_ ;
  assign \new_[18082]_  = ~\new_[12302]_ ;
  assign \new_[18083]_  = ~\new_[10318]_ ;
  assign \new_[18084]_  = ~\new_[9276]_ ;
  assign \new_[18085]_  = ~\new_[9277]_ ;
  assign \new_[18086]_  = ~\new_[10201]_ ;
  assign \new_[18087]_  = ~\new_[11289]_ ;
  assign \new_[18088]_  = ~\new_[15396]_ ;
  assign \new_[18089]_  = ~\new_[7438]_ ;
  assign \new_[18090]_  = ~\new_[7642]_ ;
  assign \new_[18091]_  = ~\new_[11543]_ ;
  assign \new_[18092]_  = ~\new_[10178]_ ;
  assign \new_[18093]_  = ~\new_[6930]_ ;
  assign \new_[18094]_  = ~\new_[12356]_ ;
  assign \new_[18095]_  = ~\new_[11826]_ ;
  assign \new_[18096]_  = ~\new_[10114]_ ;
  assign \new_[18097]_  = ~\new_[11582]_ ;
  assign \new_[18098]_  = ~\new_[13217]_ ;
  assign \new_[18099]_  = ~\new_[9775]_ ;
  assign \new_[18100]_  = ~\new_[9811]_ ;
  assign \new_[18101]_  = ~\new_[7012]_ ;
  assign \new_[18102]_  = ~\new_[9774]_ ;
  assign \new_[18103]_  = ~\new_[6905]_ ;
  assign \new_[18104]_  = ~\new_[12351]_ ;
  assign \new_[18105]_  = ~\new_[5499]_ ;
  assign \new_[18106]_  = ~\new_[6830]_ ;
  assign \new_[18107]_  = ~\new_[10104]_ ;
  assign \new_[18108]_  = ~\new_[7248]_ ;
  assign \new_[18109]_  = ~\new_[11761]_ ;
  assign \new_[18110]_  = ~\new_[10184]_ ;
  assign \new_[18111]_  = ~\new_[10187]_ ;
  assign \new_[18112]_  = ~\new_[6887]_ ;
  assign \new_[18113]_  = ~\new_[10186]_ ;
  assign \new_[18114]_  = ~\new_[11497]_ ;
  assign \new_[18115]_  = ~\new_[7480]_ ;
  assign \new_[18116]_  = ~\new_[8261]_ ;
  assign \new_[18117]_  = ~\new_[7015]_ ;
  assign \new_[18118]_  = ~\new_[11712]_ ;
  assign n16770 = ~\new_[9812]_ ;
  assign \new_[18120]_  = ~\new_[10191]_ ;
  assign \new_[18121]_  = ~\new_[6834]_ ;
  assign \new_[18122]_  = ~\new_[15123]_ ;
  assign \new_[18123]_  = ~\new_[10876]_ ;
  assign \new_[18124]_  = ~\new_[7944]_ ;
  assign \new_[18125]_  = ~\new_[11523]_ ;
  assign \new_[18126]_  = ~\new_[10245]_ ;
  assign \new_[18127]_  = ~\new_[11560]_ ;
  assign \new_[18128]_  = ~\new_[11664]_ ;
  assign \new_[18129]_  = ~\new_[11648]_ ;
  assign \new_[18130]_  = ~\new_[11508]_ ;
  assign \new_[18131]_  = ~\new_[11647]_ ;
  assign \new_[18132]_  = ~\new_[11509]_ ;
  assign n17040 = ~\new_[11346]_ ;
  assign n17080 = ~\new_[11756]_ ;
  assign \new_[18135]_  = ~\new_[6620]_ ;
  assign \new_[18136]_  = ~\new_[11348]_ ;
  assign \new_[18137]_  = ~\new_[11641]_ ;
  assign \new_[18138]_  = ~\new_[11515]_ ;
  assign \new_[18139]_  = ~\new_[11747]_ ;
  assign \new_[18140]_  = ~\new_[6661]_ ;
  assign \new_[18141]_  = ~\new_[11353]_ ;
  assign \new_[18142]_  = ~\new_[11638]_ ;
  assign \new_[18143]_  = ~\new_[11354]_ ;
  assign \new_[18144]_  = ~\new_[10887]_ ;
  assign \new_[18145]_  = ~\new_[11730]_ ;
  assign \new_[18146]_  = ~\new_[11727]_ ;
  assign \new_[18147]_  = ~\new_[10252]_ ;
  assign \new_[18148]_  = ~\new_[6693]_ ;
  assign \new_[18149]_  = ~\new_[11090]_ ;
  assign \new_[18150]_  = ~\new_[8215]_ ;
  assign \new_[18151]_  = ~\new_[7250]_ ;
  assign \new_[18152]_  = ~\new_[4458]_ ;
  assign \new_[18153]_  = ~\new_[7496]_ ;
  assign \new_[18154]_  = ~\new_[11602]_ ;
  assign \new_[18155]_  = ~\new_[12197]_ ;
  assign \new_[18156]_  = ~\new_[9825]_ ;
  assign \new_[18157]_  = ~\new_[10271]_ ;
  assign \new_[18158]_  = ~\new_[8160]_ ;
  assign \new_[18159]_  = ~\new_[10192]_ ;
  assign \new_[18160]_  = ~\new_[10110]_ ;
  assign \new_[18161]_  = ~\new_[10292]_ ;
  assign \new_[18162]_  = ~\new_[10147]_ ;
  assign \new_[18163]_  = ~\new_[12084]_ ;
  assign \new_[18164]_  = ~\new_[6957]_ ;
  assign \new_[18165]_  = ~\new_[11357]_ ;
  assign \new_[18166]_  = ~\new_[10196]_ ;
  assign \new_[18167]_  = ~\new_[12537]_ ;
  assign \new_[18168]_  = ~\new_[10307]_ ;
  assign \new_[18169]_  = ~\new_[10109]_ ;
  assign \new_[18170]_  = ~\new_[11851]_ ;
  assign \new_[18171]_  = ~\new_[7478]_ ;
  assign \new_[18172]_  = ~\new_[12300]_ ;
  assign \new_[18173]_  = ~\new_[11131]_ ;
  assign \new_[18174]_  = ~\new_[10108]_ ;
  assign \new_[18175]_  = ~\new_[10304]_ ;
  assign \new_[18176]_  = ~\new_[11106]_ ;
  assign \new_[18177]_  = ~\new_[12294]_ ;
  assign \new_[18178]_  = ~\new_[10310]_ ;
  assign \new_[18179]_  = ~\new_[10107]_ ;
  assign \new_[18180]_  = ~\new_[11359]_ ;
  assign \new_[18181]_  = ~\new_[6785]_ ;
  assign \new_[18182]_  = ~\new_[11833]_ ;
  assign \new_[18183]_  = ~\new_[11653]_ ;
  assign \new_[18184]_  = ~\new_[7460]_ ;
  assign \new_[18185]_  = ~\new_[8622]_ ;
  assign \new_[18186]_  = ~\new_[6886]_ ;
  assign \new_[18187]_  = ~\new_[11077]_ ;
  assign \new_[18188]_  = ~\new_[13616]_ ;
  assign \new_[18189]_  = ~\new_[9764]_ ;
  assign \new_[18190]_  = ~\new_[9804]_ ;
  assign \new_[18191]_  = ~\new_[6637]_ ;
  assign \new_[18192]_  = ~\new_[6738]_ ;
  assign \new_[18193]_  = ~\new_[12172]_ ;
  assign \new_[18194]_  = ~\new_[10094]_ ;
  assign \new_[18195]_  = ~\new_[6704]_ ;
  assign \new_[18196]_  = ~\new_[11529]_ ;
  assign \new_[18197]_  = ~\new_[10096]_ ;
  assign \new_[18198]_  = ~\new_[6913]_ ;
  assign \new_[18199]_  = ~\new_[9799]_ ;
  assign \new_[18200]_  = ~\new_[10206]_ ;
  assign \new_[18201]_  = ~\new_[10207]_ ;
  assign \new_[18202]_  = ~\new_[10057]_ ;
  assign \new_[18203]_  = ~\new_[10123]_ ;
  assign \new_[18204]_  = ~\new_[7658]_ ;
  assign \new_[18205]_  = ~\new_[8078]_ ;
  assign \new_[18206]_  = ~\new_[11772]_ ;
  assign \new_[18207]_  = ~\new_[11567]_ ;
  assign \new_[18208]_  = ~\new_[11533]_ ;
  assign \new_[18209]_  = ~\new_[11487]_ ;
  assign \new_[18210]_  = ~\new_[12315]_ ;
  assign \new_[18211]_  = ~\new_[11738]_ ;
  assign \new_[18212]_  = ~\new_[10198]_ ;
  assign \new_[18213]_  = ~\new_[10209]_ ;
  assign \new_[18214]_  = ~\new_[6744]_ ;
  assign \new_[18215]_  = ~\new_[13621]_ ;
  assign \new_[18216]_  = ~\new_[6740]_ ;
  assign \new_[18217]_  = ~\new_[11769]_ ;
  assign \new_[18218]_  = ~\new_[6884]_ ;
  assign \new_[18219]_  = ~\new_[6933]_ ;
  assign \new_[18220]_  = ~\new_[6583]_ ;
  assign \new_[18221]_  = ~\new_[11355]_ ;
  assign \new_[18222]_  = ~\new_[10052]_ ;
  assign \new_[18223]_  = ~\new_[10214]_ ;
  assign \new_[18224]_  = ~\new_[5014]_ ;
  assign \new_[18225]_  = ~\new_[6942]_ ;
  assign \new_[18226]_  = ~\new_[11358]_ ;
  assign \new_[18227]_  = ~\new_[9776]_ ;
  assign \new_[18228]_  = ~\new_[13622]_ ;
  assign \new_[18229]_  = ~\new_[11711]_ ;
  assign \new_[18230]_  = ~\new_[6689]_ ;
  assign \new_[18231]_  = ~\new_[6815]_ ;
  assign \new_[18232]_  = ~\new_[11962]_ ;
  assign \new_[18233]_  = ~\new_[12147]_ ;
  assign \new_[18234]_  = ~\new_[7707]_ ;
  assign \new_[18235]_  = ~\new_[12088]_ ;
  assign \new_[18236]_  = ~\new_[11362]_ ;
  assign \new_[18237]_  = ~\new_[12087]_ ;
  assign \new_[18238]_  = ~\new_[6732]_ ;
  assign \new_[18239]_  = ~\new_[5485]_ ;
  assign \new_[18240]_  = ~\new_[11821]_ ;
  assign \new_[18241]_  = ~\new_[11294]_ ;
  assign \new_[18242]_  = ~\new_[6844]_ ;
  assign \new_[18243]_  = ~\new_[11831]_ ;
  assign \new_[18244]_  = ~\new_[11402]_ ;
  assign \new_[18245]_  = ~\new_[7788]_ ;
  assign \new_[18246]_  = ~\new_[11651]_ ;
  assign \new_[18247]_  = ~\new_[9797]_ ;
  assign \new_[18248]_  = ~\new_[11364]_ ;
  assign \new_[18249]_  = ~\new_[11519]_ ;
  assign \new_[18250]_  = ~\new_[11616]_ ;
  assign \new_[18251]_  = ~n16910;
  assign \new_[18252]_  = ~\new_[12205]_ ;
  assign \new_[18253]_  = ~\new_[10224]_ ;
  assign n17065 = ~\new_[10075]_ ;
  assign \new_[18255]_  = ~\new_[12481]_ ;
  assign \new_[18256]_  = ~\new_[9809]_ ;
  assign \new_[18257]_  = ~\new_[6822]_ ;
  assign \new_[18258]_  = ~\new_[10049]_ ;
  assign \new_[18259]_  = ~\new_[11366]_ ;
  assign \new_[18260]_  = ~\new_[9815]_ ;
  assign \new_[18261]_  = ~\new_[5016]_ ;
  assign \new_[18262]_  = ~\new_[10101]_ ;
  assign \new_[18263]_  = ~\new_[10226]_ ;
  assign \new_[18264]_  = ~\new_[7262]_ ;
  assign \new_[18265]_  = ~\new_[11520]_ ;
  assign \new_[18266]_  = ~\new_[11297]_ ;
  assign \new_[18267]_  = ~\new_[11283]_ ;
  assign \new_[18268]_  = ~\new_[11521]_ ;
  assign \new_[18269]_  = ~\new_[12380]_ ;
  assign \new_[18270]_  = ~\new_[12328]_ ;
  assign \new_[18271]_  = ~\new_[12000]_ ;
  assign \new_[18272]_  = ~\new_[7679]_ ;
  assign \new_[18273]_  = ~\new_[12096]_ ;
  assign \new_[18274]_  = ~\new_[12098]_ ;
  assign \new_[18275]_  = ~\new_[12099]_ ;
  assign \new_[18276]_  = ~\new_[11351]_ ;
  assign \new_[18277]_  = ~\new_[9787]_ ;
  assign \new_[18278]_  = ~\new_[12365]_ ;
  assign \new_[18279]_  = ~\new_[11892]_ ;
  assign \new_[18280]_  = ~\new_[11783]_ ;
  assign \new_[18281]_  = ~\new_[11777]_ ;
  assign \new_[18282]_  = ~\new_[11475]_ ;
  assign \new_[18283]_  = ~\new_[12248]_ ;
  assign \new_[18284]_  = ~\new_[10138]_ ;
  assign \new_[18285]_  = ~\new_[6833]_ ;
  assign \new_[18286]_  = ~\new_[7503]_ ;
  assign \new_[18287]_  = ~\new_[6650]_ ;
  assign \new_[18288]_  = ~\new_[9784]_ ;
  assign \new_[18289]_  = ~\new_[15193]_ ;
  assign \new_[18290]_  = ~\new_[9818]_ ;
  assign \new_[18291]_  = ~\new_[11323]_ ;
  assign \new_[18292]_  = ~\new_[6607]_ ;
  assign \new_[18293]_  = ~\new_[10097]_ ;
  assign \new_[18294]_  = ~\new_[11656]_ ;
  assign \new_[18295]_  = ~\new_[8159]_ ;
  assign \new_[18296]_  = ~\new_[7806]_ ;
  assign \new_[18297]_  = ~\new_[7641]_ ;
  assign n16890 = ~\new_[10011]_ ;
  assign \new_[18299]_  = ~\new_[6651]_ ;
  assign \new_[18300]_  = ~\new_[15173]_ ;
  assign \new_[18301]_  = ~\new_[7434]_ ;
  assign \new_[18302]_  = ~\new_[10135]_ ;
  assign \new_[18303]_  = ~\new_[7764]_ ;
  assign \new_[18304]_  = ~\new_[11481]_ ;
  assign \new_[18305]_  = ~\new_[11372]_ ;
  assign \new_[18306]_  = ~\new_[10194]_ ;
  assign \new_[18307]_  = ~\new_[12001]_ ;
  assign \new_[18308]_  = ~\new_[5103]_ ;
  assign \new_[18309]_  = ~\new_[12163]_ ;
  assign \new_[18310]_  = ~\new_[11081]_ ;
  assign \new_[18311]_  = ~\new_[6737]_ ;
  assign \new_[18312]_  = ~\new_[10091]_ ;
  assign \new_[18313]_  = ~\new_[12175]_ ;
  assign \new_[18314]_  = ~\new_[6926]_ ;
  assign \new_[18315]_  = ~\new_[6642]_ ;
  assign \new_[18316]_  = ~\new_[12176]_ ;
  assign \new_[18317]_  = ~\new_[10365]_ ;
  assign \new_[18318]_  = ~\new_[11811]_ ;
  assign \new_[18319]_  = ~\new_[11604]_ ;
  assign \new_[18320]_  = ~\new_[11318]_ ;
  assign \new_[18321]_  = ~\new_[5017]_ ;
  assign \new_[18322]_  = ~\new_[7746]_ ;
  assign \new_[18323]_  = ~\new_[10129]_ ;
  assign \new_[18324]_  = ~\new_[6617]_ ;
  assign \new_[18325]_  = ~\new_[4092]_ ;
  assign \new_[18326]_  = ~\new_[6857]_ ;
  assign \new_[18327]_  = ~\new_[11373]_ ;
  assign n17020 = ~\new_[10076]_ ;
  assign \new_[18329]_  = ~\new_[6840]_ ;
  assign \new_[18330]_  = ~\new_[11377]_ ;
  assign \new_[18331]_  = ~\new_[10128]_ ;
  assign \new_[18332]_  = ~\new_[7293]_ ;
  assign \new_[18333]_  = ~\new_[11846]_ ;
  assign \new_[18334]_  = ~\new_[12159]_ ;
  assign \new_[18335]_  = ~\new_[7442]_ ;
  assign \new_[18336]_  = ~\new_[11435]_ ;
  assign \new_[18337]_  = ~\new_[5026]_ ;
  assign \new_[18338]_  = ~\new_[13720]_ ;
  assign \new_[18339]_  = ~\new_[6591]_ ;
  assign \new_[18340]_  = ~\new_[11844]_ ;
  assign \new_[18341]_  = ~\new_[6688]_ ;
  assign \new_[18342]_  = ~\new_[6618]_ ;
  assign \new_[18343]_  = ~\new_[7461]_ ;
  assign \new_[18344]_  = ~\new_[12136]_ ;
  assign \new_[18345]_  = ~\new_[11432]_ ;
  assign \new_[18346]_  = ~\new_[11110]_ ;
  assign \new_[18347]_  = ~\new_[9281]_ ;
  assign \new_[18348]_  = ~\new_[12335]_ ;
  assign \new_[18349]_  = ~\new_[11450]_ ;
  assign \new_[18350]_  = ~\new_[10233]_ ;
  assign \new_[18351]_  = ~\new_[6622]_ ;
  assign \new_[18352]_  = ~\new_[11693]_ ;
  assign \new_[18353]_  = ~\new_[10089]_ ;
  assign \new_[18354]_  = ~\new_[6719]_ ;
  assign \new_[18355]_  = ~\new_[11479]_ ;
  assign \new_[18356]_  = ~\new_[10298]_ ;
  assign \new_[18357]_  = ~\new_[8218]_ ;
  assign \new_[18358]_  = ~\new_[11379]_ ;
  assign \new_[18359]_  = ~\new_[6700]_ ;
  assign \new_[18360]_  = ~\new_[12258]_ ;
  assign \new_[18361]_  = ~\new_[11314]_ ;
  assign \new_[18362]_  = ~\new_[4978]_ ;
  assign \new_[18363]_  = ~\new_[11383]_ ;
  assign \new_[18364]_  = ~\new_[12105]_ ;
  assign \new_[18365]_  = ~\new_[11311]_ ;
  assign \new_[18366]_  = ~\new_[6602]_ ;
  assign \new_[18367]_  = ~\new_[10294]_ ;
  assign \new_[18368]_  = ~\new_[11312]_ ;
  assign \new_[18369]_  = ~\new_[11384]_ ;
  assign \new_[18370]_  = ~\new_[10273]_ ;
  assign \new_[18371]_  = ~\new_[11387]_ ;
  assign \new_[18372]_  = ~\new_[12244]_ ;
  assign \new_[18373]_  = ~\new_[10241]_ ;
  assign \new_[18374]_  = ~\new_[11842]_ ;
  assign \new_[18375]_  = ~\new_[12250]_ ;
  assign \new_[18376]_  = ~\new_[12246]_ ;
  assign \new_[18377]_  = ~\new_[12108]_ ;
  assign \new_[18378]_  = ~\new_[12102]_ ;
  assign \new_[18379]_  = ~\new_[11534]_ ;
  assign \new_[18380]_  = ~\new_[10230]_ ;
  assign \new_[18381]_  = ~\new_[6879]_ ;
  assign \new_[18382]_  = ~\new_[9231]_ ;
  assign \new_[18383]_  = ~\new_[11517]_ ;
  assign \new_[18384]_  = ~\new_[6923]_ ;
  assign \new_[18385]_  = ~\new_[6686]_ ;
  assign \new_[18386]_  = ~\new_[5483]_ ;
  assign \new_[18387]_  = ~\new_[12341]_ ;
  assign \new_[18388]_  = ~\new_[6762]_ ;
  assign \new_[18389]_  = ~\new_[11126]_ ;
  assign \new_[18390]_  = ~\new_[7441]_ ;
  assign \new_[18391]_  = ~\new_[11717]_ ;
  assign \new_[18392]_  = ~\new_[10386]_ ;
  assign \new_[18393]_  = ~\new_[12346]_ ;
  assign \new_[18394]_  = ~\new_[6646]_ ;
  assign \new_[18395]_  = ~\new_[11445]_ ;
  assign \new_[18396]_  = ~\new_[11130]_ ;
  assign \new_[18397]_  = ~\new_[11300]_ ;
  assign \new_[18398]_  = ~\new_[12212]_ ;
  assign \new_[18399]_  = ~\new_[6765]_ ;
  assign \new_[18400]_  = ~\new_[12126]_ ;
  assign \new_[18401]_  = ~\new_[6764]_ ;
  assign \new_[18402]_  = ~\new_[8144]_ ;
  assign \new_[18403]_  = ~\new_[11617]_ ;
  assign \new_[18404]_  = ~\new_[7440]_ ;
  assign \new_[18405]_  = ~\new_[11486]_ ;
  assign \new_[18406]_  = ~\new_[9782]_ ;
  assign \new_[18407]_  = ~\new_[11285]_ ;
  assign \new_[18408]_  = ~\new_[12168]_ ;
  assign \new_[18409]_  = ~\new_[9194]_ ;
  assign \new_[18410]_  = ~\new_[12320]_ ;
  assign \new_[18411]_  = ~\new_[12297]_ ;
  assign \new_[18412]_  = ~\new_[7251]_ ;
  assign \new_[18413]_  = ~\new_[12381]_ ;
  assign \new_[18414]_  = ~\new_[11694]_ ;
  assign \new_[18415]_  = ~\new_[12157]_ ;
  assign \new_[18416]_  = ~\new_[6980]_ ;
  assign \new_[18417]_  = ~\new_[11808]_ ;
  assign \new_[18418]_  = ~\new_[12186]_ ;
  assign \new_[18419]_  = ~\new_[10287]_ ;
  assign \new_[18420]_  = ~\new_[11271]_ ;
  assign \new_[18421]_  = ~\new_[7471]_ ;
  assign \new_[18422]_  = ~\new_[10303]_ ;
  assign \new_[18423]_  = ~\new_[12260]_ ;
  assign \new_[18424]_  = ~\new_[11716]_ ;
  assign \new_[18425]_  = ~\new_[5030]_ ;
  assign \new_[18426]_  = ~\new_[11292]_ ;
  assign \new_[18427]_  = ~\new_[9195]_ ;
  assign \new_[18428]_  = ~\new_[15149]_ ;
  assign \new_[18429]_  = ~\new_[11096]_ ;
  assign \new_[18430]_  = ~\new_[12170]_ ;
  assign \new_[18431]_  = ~\new_[12117]_ ;
  assign \new_[18432]_  = ~\new_[12116]_ ;
  assign \new_[18433]_  = ~\new_[11997]_ ;
  assign \new_[18434]_  = ~\new_[7665]_ ;
  assign \new_[18435]_  = ~\new_[5031]_ ;
  assign \new_[18436]_  = ~\new_[6931]_ ;
  assign \new_[18437]_  = ~\new_[15925]_ ;
  assign \new_[18438]_  = ~\new_[9828]_ ;
  assign \new_[18439]_  = ~\new_[11280]_ ;
  assign \new_[18440]_  = ~\new_[7954]_ ;
  assign \new_[18441]_  = ~\new_[9781]_ ;
  assign \new_[18442]_  = ~\new_[12152]_ ;
  assign \new_[18443]_  = ~\new_[6959]_ ;
  assign \new_[18444]_  = ~\new_[6827]_ ;
  assign \new_[18445]_  = ~n16995;
  assign \new_[18446]_  = ~\new_[11392]_ ;
  assign \new_[18447]_  = ~\new_[11910]_ ;
  assign \new_[18448]_  = ~\new_[10881]_ ;
  assign \new_[18449]_  = ~\new_[11400]_ ;
  assign \new_[18450]_  = ~\new_[11267]_ ;
  assign \new_[18451]_  = ~\new_[11601]_ ;
  assign \new_[18452]_  = ~\new_[12003]_ ;
  assign \new_[18453]_  = ~\new_[6775]_ ;
  assign \new_[18454]_  = ~\new_[11896]_ ;
  assign \new_[18455]_  = ~\new_[6770]_ ;
  assign \new_[18456]_  = ~\new_[11510]_ ;
  assign \new_[18457]_  = ~\new_[7953]_ ;
  assign \new_[18458]_  = ~\new_[10497]_ ;
  assign \new_[18459]_  = ~\new_[7443]_ ;
  assign \new_[18460]_  = ~\new_[7966]_ ;
  assign \new_[18461]_  = ~\new_[12241]_ ;
  assign \new_[18462]_  = ~\new_[5174]_ ;
  assign \new_[18463]_  = ~\new_[11823]_ ;
  assign \new_[18464]_  = ~\new_[11992]_ ;
  assign \new_[18465]_  = ~\new_[12121]_ ;
  assign \new_[18466]_  = ~\new_[11980]_ ;
  assign \new_[18467]_  = ~\new_[11405]_ ;
  assign \new_[18468]_  = ~\new_[11764]_ ;
  assign \new_[18469]_  = ~\new_[6808]_ ;
  assign \new_[18470]_  = ~\new_[11810]_ ;
  assign n17030 = ~\new_[5060]_ ;
  assign \new_[18472]_  = ~\new_[6797]_ ;
  assign \new_[18473]_  = ~\new_[11409]_ ;
  assign \new_[18474]_  = ~\new_[11436]_ ;
  assign \new_[18475]_  = ~\new_[9201]_ ;
  assign \new_[18476]_  = ~\new_[10340]_ ;
  assign \new_[18477]_  = ~\new_[12119]_ ;
  assign \new_[18478]_  = ~\new_[11411]_ ;
  assign \new_[18479]_  = ~\new_[11406]_ ;
  assign \new_[18480]_  = ~\new_[5484]_ ;
  assign \new_[18481]_  = ~\new_[5034]_ ;
  assign \new_[18482]_  = ~\new_[12527]_ ;
  assign \new_[18483]_  = ~\new_[6656]_ ;
  assign \new_[18484]_  = ~\new_[6843]_ ;
  assign \new_[18485]_  = ~\new_[12424]_ ;
  assign \new_[18486]_  = ~\new_[11557]_ ;
  assign \new_[18487]_  = ~\new_[7669]_ ;
  assign \new_[18488]_  = ~\wbm_cti_o[1] ;
  assign \new_[18489]_  = ~\new_[11370]_ ;
  assign \new_[18490]_  = ~\new_[12333]_ ;
  assign \new_[18491]_  = ~\new_[5013]_ ;
  assign \new_[18492]_  = ~\new_[9196]_ ;
  assign \new_[18493]_  = ~\new_[12129]_ ;
  assign \new_[18494]_  = ~\new_[12131]_ ;
  assign \new_[18495]_  = ~\new_[11418]_ ;
  assign \new_[18496]_  = ~\new_[12130]_ ;
  assign \new_[18497]_  = ~\new_[12486]_ ;
  assign \new_[18498]_  = ~\new_[12388]_ ;
  assign \new_[18499]_  = ~\new_[6585]_ ;
  assign \new_[18500]_  = ~\new_[12185]_ ;
  assign \new_[18501]_  = ~\new_[6653]_ ;
  assign \new_[18502]_  = ~\new_[4009]_ ;
  assign \new_[18503]_  = ~\new_[7869]_ ;
  assign \new_[18504]_  = ~\new_[6826]_ ;
  assign \new_[18505]_  = ~\new_[12326]_ ;
  assign \new_[18506]_  = ~\new_[7470]_ ;
  assign \new_[18507]_  = ~\new_[7510]_ ;
  assign \new_[18508]_  = ~\new_[11994]_ ;
  assign \new_[18509]_  = ~\new_[9792]_ ;
  assign \new_[18510]_  = ~\new_[10099]_ ;
  assign \new_[18511]_  = ~\new_[7751]_ ;
  assign \new_[18512]_  = ~\new_[5057]_ ;
  assign \new_[18513]_  = ~\new_[6786]_ ;
  assign \new_[18514]_  = ~\new_[10092]_ ;
  assign \new_[18515]_  = ~\new_[9680]_ ;
  assign \new_[18516]_  = ~\new_[6958]_ ;
  assign \new_[18517]_  = ~\new_[5036]_ ;
  assign \new_[18518]_  = ~\new_[9229]_ ;
  assign \new_[18519]_  = ~\new_[11454]_ ;
  assign \new_[18520]_  = ~\new_[9786]_ ;
  assign \new_[18521]_  = ~\new_[5482]_ ;
  assign \new_[18522]_  = ~\new_[10339]_ ;
  assign \new_[18523]_  = ~wbm_rty_i;
  assign \new_[18524]_  = ~\new_[11959]_ ;
  assign \new_[18525]_  = ~\new_[11790]_ ;
  assign \new_[18526]_  = ~\new_[6654]_ ;
  assign \new_[18527]_  = ~\new_[12135]_ ;
  assign \new_[18528]_  = ~\new_[6630]_ ;
  assign \new_[18529]_  = ~\new_[6612]_ ;
  assign \new_[18530]_  = ~\new_[6882]_ ;
  assign \new_[18531]_  = ~\new_[11719]_ ;
  assign \new_[18532]_  = ~\new_[6708]_ ;
  assign \new_[18533]_  = ~\new_[11565]_ ;
  assign \new_[18534]_  = ~\new_[5105]_ ;
  assign \new_[18535]_  = ~\new_[11855]_ ;
  assign \new_[18536]_  = ~\new_[6929]_ ;
  assign \new_[18537]_  = ~\new_[6603]_ ;
  assign \new_[18538]_  = ~\new_[11579]_ ;
  assign \new_[18539]_  = ~\new_[10331]_ ;
  assign \new_[18540]_  = ~\new_[7281]_ ;
  assign \new_[18541]_  = ~\new_[7473]_ ;
  assign \new_[18542]_  = ~\new_[10088]_ ;
  assign \new_[18543]_  = ~\new_[12120]_ ;
  assign \new_[18544]_  = ~\new_[6885]_ ;
  assign \new_[18545]_  = ~\new_[6318]_ ;
  assign \new_[18546]_  = ~\new_[11407]_ ;
  assign \new_[18547]_  = ~\new_[10319]_ ;
  assign \new_[18548]_  = ~\new_[7406]_ ;
  assign \new_[18549]_  = ~\new_[12330]_ ;
  assign \new_[18550]_  = ~\new_[11419]_ ;
  assign \new_[18551]_  = ~\new_[11836]_ ;
  assign \new_[18552]_  = ~\new_[12522]_ ;
  assign \new_[18553]_  = ~\new_[7275]_ ;
  assign \new_[18554]_  = ~\new_[7866]_ ;
  assign \new_[18555]_  = ~\new_[11108]_ ;
  assign \new_[18556]_  = ~\new_[11792]_ ;
  assign \new_[18557]_  = ~\new_[6626]_ ;
  assign \new_[18558]_  = ~\new_[11610]_ ;
  assign \new_[18559]_  = ~\new_[6954]_ ;
  assign \new_[18560]_  = ~\new_[11084]_ ;
  assign \new_[18561]_  = ~\new_[11524]_ ;
  assign \new_[18562]_  = ~\new_[10143]_ ;
  assign \new_[18563]_  = ~\new_[6813]_ ;
  assign \new_[18564]_  = ~\new_[11580]_ ;
  assign \new_[18565]_  = ~\new_[5032]_ ;
  assign \new_[18566]_  = ~\new_[11422]_ ;
  assign \new_[18567]_  = ~\new_[6877]_ ;
  assign \new_[18568]_  = ~\new_[8213]_ ;
  assign \new_[18569]_  = ~\new_[6725]_ ;
  assign \new_[18570]_  = ~\new_[12173]_ ;
  assign \new_[18571]_  = ~\new_[6805]_ ;
  assign \new_[18572]_  = ~\new_[12256]_ ;
  assign \new_[18573]_  = ~\new_[6599]_ ;
  assign \new_[18574]_  = ~\new_[11092]_ ;
  assign \new_[18575]_  = ~\new_[11999]_ ;
  assign \new_[18576]_  = ~\new_[11817]_ ;
  assign \new_[18577]_  = ~\new_[12202]_ ;
  assign \new_[18578]_  = ~\new_[6836]_ ;
  assign \new_[18579]_  = ~\new_[10313]_ ;
  assign \new_[18580]_  = ~\new_[10300]_ ;
  assign \new_[18581]_  = ~\new_[6918]_ ;
  assign \new_[18582]_  = ~\new_[11279]_ ;
  assign \new_[18583]_  = ~\new_[14866]_ ;
  assign \new_[18584]_  = ~\new_[4094]_ ;
  assign \new_[18585]_  = ~\new_[6924]_ ;
  assign \new_[18586]_  = ~\new_[11093]_ ;
  assign \new_[18587]_  = ~\new_[11507]_ ;
  assign \new_[18588]_  = ~\new_[10221]_ ;
  assign \new_[18589]_  = ~\new_[9783]_ ;
  assign \new_[18590]_  = ~\new_[12301]_ ;
  assign \new_[18591]_  = ~\new_[11431]_ ;
  assign \new_[18592]_  = ~\new_[12337]_ ;
  assign \new_[18593]_  = ~\new_[11701]_ ;
  assign \new_[18594]_  = ~\new_[9817]_ ;
  assign \new_[18595]_  = ~\new_[9793]_ ;
  assign \new_[18596]_  = ~\new_[9785]_ ;
  assign \new_[18597]_  = ~\new_[10102]_ ;
  assign \new_[18598]_  = ~\new_[5415]_ ;
  assign \new_[18599]_  = ~\new_[12278]_ ;
  assign \new_[18600]_  = ~\new_[5503]_ ;
  assign \new_[18601]_  = ~\new_[6874]_ ;
  assign \new_[18602]_  = ~\new_[11748]_ ;
  assign \new_[18603]_  = ~\new_[5501]_ ;
  assign \new_[18604]_  = ~\new_[6782]_ ;
  assign \new_[18605]_  = ~\new_[11781]_ ;
  assign \new_[18606]_  = ~\new_[11097]_ ;
  assign \new_[18607]_  = ~\new_[5471]_ ;
  assign \new_[18608]_  = ~\new_[7463]_ ;
  assign \new_[18609]_  = ~\new_[15091]_ ;
  assign \new_[18610]_  = ~\new_[12357]_ ;
  assign \new_[18611]_  = ~\new_[11303]_ ;
  assign \new_[18612]_  = ~\new_[11978]_ ;
  assign \new_[18613]_  = ~\new_[11394]_ ;
  assign \new_[18614]_  = ~\new_[6707]_ ;
  assign \new_[18615]_  = ~\new_[10375]_ ;
  assign \new_[18616]_  = ~\new_[11578]_ ;
  assign \new_[18617]_  = ~\new_[10341]_ ;
  assign \new_[18618]_  = ~\new_[8142]_ ;
  assign \new_[18619]_  = ~\new_[10308]_ ;
  assign \new_[18620]_  = ~\new_[11605]_ ;
  assign \new_[18621]_  = ~\new_[6855]_ ;
  assign \new_[18622]_  = ~\new_[12100]_ ;
  assign \new_[18623]_  = ~\new_[12252]_ ;
  assign \new_[18624]_  = ~\new_[15118]_ ;
  assign \new_[18625]_  = ~\new_[12097]_ ;
  assign \new_[18626]_  = ~\new_[12123]_ ;
  assign \new_[18627]_  = ~\new_[6616]_ ;
  assign \new_[18628]_  = ~\new_[9778]_ ;
  assign \new_[18629]_  = ~\new_[11791]_ ;
  assign \new_[18630]_  = ~\new_[6878]_ ;
  assign \new_[18631]_  = ~\new_[6639]_ ;
  assign \new_[18632]_  = ~\new_[11453]_ ;
  assign \new_[18633]_  = ~\new_[6601]_ ;
  assign \new_[18634]_  = ~\new_[12270]_ ;
  assign \new_[18635]_  = ~\new_[12234]_ ;
  assign \new_[18636]_  = ~\new_[6839]_ ;
  assign \new_[18637]_  = ~\new_[6714]_ ;
  assign \new_[18638]_  = ~\new_[12282]_ ;
  assign \new_[18639]_  = ~\new_[7458]_ ;
  assign \new_[18640]_  = ~\new_[7241]_ ;
  assign \new_[18641]_  = ~\new_[6645]_ ;
  assign \new_[18642]_  = ~\new_[15389]_ ;
  assign \new_[18643]_  = ~\new_[11746]_ ;
  assign \new_[18644]_  = ~\new_[11538]_ ;
  assign \new_[18645]_  = ~\new_[11820]_ ;
  assign \new_[18646]_  = ~\new_[11415]_ ;
  assign \new_[18647]_  = ~\new_[11983]_ ;
  assign \new_[18648]_  = ~\new_[11799]_ ;
  assign \new_[18649]_  = ~\new_[15390]_ ;
  assign \new_[18650]_  = ~\new_[11391]_ ;
  assign \new_[18651]_  = ~\new_[12307]_ ;
  assign \new_[18652]_  = ~\new_[12199]_ ;
  assign \new_[18653]_  = ~\new_[11839]_ ;
  assign \new_[18654]_  = ~\new_[6597]_ ;
  assign \new_[18655]_  = ~\new_[6823]_ ;
  assign \new_[18656]_  = ~\new_[11495]_ ;
  assign \new_[18657]_  = ~\new_[7258]_ ;
  assign \new_[18658]_  = ~\new_[11550]_ ;
  assign \new_[18659]_  = ~\new_[11469]_ ;
  assign \new_[18660]_  = ~\new_[12249]_ ;
  assign \new_[18661]_  = ~\new_[11100]_ ;
  assign \new_[18662]_  = ~\new_[12146]_ ;
  assign \new_[18663]_  = ~\new_[11812]_ ;
  assign \new_[18664]_  = ~\new_[5033]_ ;
  assign \new_[18665]_  = ~\new_[7771]_ ;
  assign \new_[18666]_  = ~\new_[7483]_ ;
  assign \new_[18667]_  = ~\new_[6709]_ ;
  assign \new_[18668]_  = ~\new_[6606]_ ;
  assign \new_[18669]_  = ~\new_[12348]_ ;
  assign \new_[18670]_  = ~\new_[6735]_ ;
  assign n17035 = ~\new_[10050]_ ;
  assign \new_[18672]_  = ~\new_[11768]_ ;
  assign \new_[18673]_  = ~\new_[5414]_ ;
  assign \new_[18674]_  = ~\new_[11729]_ ;
  assign \new_[18675]_  = ~\new_[6691]_ ;
  assign \new_[18676]_  = ~\new_[7631]_ ;
  assign \new_[18677]_  = ~\new_[5064]_ ;
  assign \new_[18678]_  = ~\new_[9773]_ ;
  assign \new_[18679]_  = ~\new_[11388]_ ;
  assign \new_[18680]_  = ~\new_[8687]_ ;
  assign \new_[18681]_  = ~\new_[5050]_ ;
  assign \new_[18682]_  = ~\new_[6680]_ ;
  assign \new_[18683]_  = ~\new_[11829]_ ;
  assign \new_[18684]_  = ~\new_[7451]_ ;
  assign \new_[18685]_  = ~\new_[7448]_ ;
  assign \new_[18686]_  = ~\new_[11774]_ ;
  assign \new_[18687]_  = ~\new_[6873]_ ;
  assign \new_[18688]_  = ~\new_[11574]_ ;
  assign \new_[18689]_  = ~\new_[11938]_ ;
  assign \new_[18690]_  = ~\new_[11575]_ ;
  assign \new_[18691]_  = ~\new_[6715]_ ;
  assign \new_[18692]_  = ~\new_[6746]_ ;
  assign \new_[18693]_  = ~\new_[7437]_ ;
  assign \new_[18694]_  = ~\new_[6755]_ ;
  assign \new_[18695]_  = ~\new_[6672]_ ;
  assign \new_[18696]_  = ~\new_[7446]_ ;
  assign \new_[18697]_  = ~\new_[11700]_ ;
  assign \new_[18698]_  = ~\new_[11316]_ ;
  assign \new_[18699]_  = ~\new_[12104]_ ;
  assign \new_[18700]_  = ~\new_[11363]_ ;
  assign \new_[18701]_  = ~\new_[6587]_ ;
  assign \new_[18702]_  = ~\new_[12095]_ ;
  assign \new_[18703]_  = ~\new_[11074]_ ;
  assign \new_[18704]_  = ~\new_[11385]_ ;
  assign \new_[18705]_  = ~\new_[7230]_ ;
  assign \new_[18706]_  = ~\new_[12526]_ ;
  assign \new_[18707]_  = ~\new_[6624]_ ;
  assign \new_[18708]_  = ~\new_[12124]_ ;
  assign \new_[18709]_  = ~\new_[12421]_ ;
  assign \new_[18710]_  = ~\new_[12092]_ ;
  assign \new_[18711]_  = ~\new_[13618]_ ;
  assign \new_[18712]_  = ~\new_[12141]_ ;
  assign \new_[18713]_  = ~\new_[12257]_ ;
  assign \new_[18714]_  = ~\new_[11715]_ ;
  assign \new_[18715]_  = ~\new_[10376]_ ;
  assign \new_[18716]_  = ~\new_[11381]_ ;
  assign \new_[18717]_  = ~\new_[12151]_ ;
  assign \new_[18718]_  = ~\new_[6758]_ ;
  assign \new_[18719]_  = ~\new_[11367]_ ;
  assign \new_[18720]_  = ~\new_[6600]_ ;
  assign \new_[18721]_  = ~\new_[11503]_ ;
  assign \new_[18722]_  = ~\new_[6898]_ ;
  assign \new_[18723]_  = ~\new_[6949]_ ;
  assign \new_[18724]_  = ~\new_[8046]_ ;
  assign \new_[18725]_  = ~\new_[13633]_ ;
  assign n16715 = ~\new_[11332]_ ;
  assign \new_[18727]_  = ~\new_[11269]_ ;
  assign \new_[18728]_  = ~\new_[11593]_ ;
  assign \new_[18729]_  = ~\new_[9884]_ ;
  assign \new_[18730]_  = ~\new_[6666]_ ;
  assign \new_[18731]_  = ~\new_[12363]_ ;
  assign \new_[18732]_  = ~\new_[10378]_ ;
  assign \new_[18733]_  = ~\new_[9789]_ ;
  assign \new_[18734]_  = ~\new_[11805]_ ;
  assign \new_[18735]_  = ~\new_[11998]_ ;
  assign \new_[18736]_  = ~\new_[7234]_ ;
  assign \new_[18737]_  = ~\new_[11899]_ ;
  assign \new_[18738]_  = ~\new_[7494]_ ;
  assign \new_[18739]_  = ~\new_[11522]_ ;
  assign \new_[18740]_  = ~\new_[11720]_ ;
  assign \new_[18741]_  = ~\new_[7468]_ ;
  assign \new_[18742]_  = ~\new_[11299]_ ;
  assign \new_[18743]_  = ~\new_[11695]_ ;
  assign \new_[18744]_  = ~\new_[11471]_ ;
  assign \new_[18745]_  = ~\new_[12255]_ ;
  assign \new_[18746]_  = ~\new_[11837]_ ;
  assign \new_[18747]_  = ~\new_[6584]_ ;
  assign \new_[18748]_  = ~\new_[8902]_ ;
  assign \new_[18749]_  = ~\new_[7236]_ ;
  assign \new_[18750]_  = ~\new_[11763]_ ;
  assign \new_[18751]_  = ~\new_[11270]_ ;
  assign \new_[18752]_  = ~\new_[6614]_ ;
  assign \new_[18753]_  = ~\new_[6904]_ ;
  assign \new_[18754]_  = ~\new_[11526]_ ;
  assign \new_[18755]_  = ~\new_[11386]_ ;
  assign \new_[18756]_  = ~\new_[9791]_ ;
  assign \new_[18757]_  = ~\new_[12374]_ ;
  assign \new_[18758]_  = ~\new_[7705]_ ;
  assign \new_[18759]_  = ~\new_[7431]_ ;
  assign \new_[18760]_  = ~\new_[12361]_ ;
  assign \new_[18761]_  = ~\new_[12325]_ ;
  assign \new_[18762]_  = ~\new_[7491]_ ;
  assign \new_[18763]_  = ~\new_[11310]_ ;
  assign \new_[18764]_  = ~\new_[12194]_ ;
  assign \new_[18765]_  = ~\new_[11499]_ ;
  assign \new_[18766]_  = ~\new_[11490]_ ;
  assign \new_[18767]_  = ~\new_[11281]_ ;
  assign \new_[18768]_  = ~\new_[11426]_ ;
  assign \new_[18769]_  = ~\new_[7505]_ ;
  assign \new_[18770]_  = ~\new_[11111]_ ;
  assign \new_[18771]_  = ~\new_[6664]_ ;
  assign \new_[18772]_  = ~\new_[11827]_ ;
  assign \new_[18773]_  = ~\new_[12106]_ ;
  assign \new_[18774]_  = ~\new_[10081]_ ;
  assign \new_[18775]_  = ~\new_[7967]_ ;
  assign \new_[18776]_  = ~\new_[6690]_ ;
  assign \new_[18777]_  = ~\new_[6611]_ ;
  assign \new_[18778]_  = ~\new_[12402]_ ;
  assign \new_[18779]_  = ~\new_[8210]_ ;
  assign \new_[18780]_  = ~\new_[11722]_ ;
  assign \new_[18781]_  = ~\new_[6799]_ ;
  assign \new_[18782]_  = ~\new_[11472]_ ;
  assign \new_[18783]_  = ~\new_[6795]_ ;
  assign \new_[18784]_  = ~\new_[12103]_ ;
  assign \new_[18785]_  = ~\new_[12518]_ ;
  assign \new_[18786]_  = ~\new_[9622]_ ;
  assign \new_[18787]_  = ~\new_[11571]_ ;
  assign \new_[18788]_  = ~\new_[10079]_ ;
  assign \new_[18789]_  = ~\new_[5062]_ ;
  assign \new_[18790]_  = ~\new_[6806]_ ;
  assign \new_[18791]_  = ~\new_[4973]_ ;
  assign \new_[18792]_  = ~\new_[11380]_ ;
  assign \new_[18793]_  = ~\new_[11428]_ ;
  assign \new_[18794]_  = ~\new_[6683]_ ;
  assign \new_[18795]_  = ~\new_[11501]_ ;
  assign \new_[18796]_  = ~\new_[6796]_ ;
  assign \new_[18797]_  = ~\new_[11569]_ ;
  assign \new_[18798]_  = ~\new_[9677]_ ;
  assign \new_[18799]_  = ~\new_[12373]_ ;
  assign \new_[18800]_  = ~\new_[12535]_ ;
  assign \new_[18801]_  = ~\new_[11275]_ ;
  assign \new_[18802]_  = ~\new_[12385]_ ;
  assign \new_[18803]_  = ~\new_[12178]_ ;
  assign \new_[18804]_  = ~\new_[12180]_ ;
  assign \new_[18805]_  = ~\new_[11561]_ ;
  assign \new_[18806]_  = ~\new_[12179]_ ;
  assign \new_[18807]_  = ~\new_[13617]_ ;
  assign n17085 = ~\new_[10073]_ ;
  assign \new_[18809]_  = ~\new_[12369]_ ;
  assign \new_[18810]_  = ~\new_[13490]_ ;
  assign \new_[18811]_  = ~\new_[6676]_ ;
  assign \new_[18812]_  = ~\new_[11696]_ ;
  assign \new_[18813]_  = ~\new_[11546]_ ;
  assign \new_[18814]_  = ~\new_[9788]_ ;
  assign \new_[18815]_  = ~\new_[10880]_ ;
  assign \new_[18816]_  = ~\new_[12184]_ ;
  assign \new_[18817]_  = ~\new_[11726]_ ;
  assign \new_[18818]_  = ~\new_[6824]_ ;
  assign \new_[18819]_  = ~\new_[11982]_ ;
  assign \new_[18820]_  = ~\new_[6613]_ ;
  assign \new_[18821]_  = ~\new_[12324]_ ;
  assign n16920 = ~\new_[10072]_ ;
  assign n16750 = ~\new_[3994]_ ;
  assign \new_[18824]_  = ~\new_[11583]_ ;
  assign \new_[18825]_  = ~\new_[15231]_ ;
  assign \new_[18826]_  = ~\new_[6632]_ ;
  assign \new_[18827]_  = ~\new_[12298]_ ;
  assign \new_[18828]_  = ~\new_[7488]_ ;
  assign \new_[18829]_  = ~\new_[11597]_ ;
  assign \new_[18830]_  = ~\new_[11838]_ ;
  assign \new_[18831]_  = ~\new_[11699]_ ;
  assign \new_[18832]_  = ~\new_[11947]_ ;
  assign \new_[18833]_  = ~\new_[12352]_ ;
  assign \new_[18834]_  = ~\new_[11308]_ ;
  assign \new_[18835]_  = ~\new_[10316]_ ;
  assign \new_[18836]_  = ~\new_[11504]_ ;
  assign \new_[18837]_  = ~\new_[12107]_ ;
  assign \new_[18838]_  = ~\new_[10379]_ ;
  assign \new_[18839]_  = ~\new_[9823]_ ;
  assign \new_[18840]_  = ~\new_[10080]_ ;
  assign \new_[18841]_  = ~\new_[12368]_ ;
  assign \new_[18842]_  = ~\new_[11500]_ ;
  assign \new_[18843]_  = ~\new_[9816]_ ;
  assign \new_[18844]_  = ~\new_[6941]_ ;
  assign \new_[18845]_  = ~\new_[6648]_ ;
  assign \new_[18846]_  = ~\new_[6625]_ ;
  assign \new_[18847]_  = ~\new_[8149]_ ;
  assign \new_[18848]_  = ~\new_[5481]_ ;
  assign \new_[18849]_  = ~\new_[12492]_ ;
  assign \new_[18850]_  = ~\new_[11948]_ ;
  assign \new_[18851]_  = ~\new_[7445]_ ;
  assign \new_[18852]_  = ~\new_[11083]_ ;
  assign \new_[18853]_  = ~\new_[12253]_ ;
  assign \new_[18854]_  = ~\new_[12419]_ ;
  assign \new_[18855]_  = ~\new_[11496]_ ;
  assign \new_[18856]_  = ~\new_[6665]_ ;
  assign \new_[18857]_  = ~\new_[6677]_ ;
  assign \new_[18858]_  = ~\new_[12342]_ ;
  assign \new_[18859]_  = ~\new_[11773]_ ;
  assign \new_[18860]_  = ~n16930;
  assign n17050 = ~\new_[11782]_ ;
  assign \new_[18862]_  = ~\new_[11753]_ ;
  assign \new_[18863]_  = ~\new_[6862]_ ;
  assign \new_[18864]_  = ~\new_[11608]_ ;
  assign \new_[18865]_  = ~\new_[11657]_ ;
  assign \new_[18866]_  = ~\new_[12525]_ ;
  assign \new_[18867]_  = ~\new_[11494]_ ;
  assign \new_[18868]_  = ~\new_[10182]_ ;
  assign \new_[18869]_  = ~\new_[6948]_ ;
  assign \new_[18870]_  = ~\new_[12128]_ ;
  assign \new_[18871]_  = ~\new_[10180]_ ;
  assign \new_[18872]_  = ~\new_[11767]_ ;
  assign \new_[18873]_  = ~\new_[7508]_ ;
  assign \new_[18874]_  = ~\new_[10336]_ ;
  assign \new_[18875]_  = ~\new_[11594]_ ;
  assign \new_[18876]_  = ~\new_[6596]_ ;
  assign \new_[18877]_  = ~\new_[7464]_ ;
  assign \new_[18878]_  = ~\new_[6852]_ ;
  assign \new_[18879]_  = ~\new_[7242]_ ;
  assign \new_[18880]_  = ~\new_[11425]_ ;
  assign \new_[18881]_  = ~\new_[6865]_ ;
  assign \new_[18882]_  = ~\new_[11757]_ ;
  assign \new_[18883]_  = ~\new_[11815]_ ;
  assign \new_[18884]_  = ~\new_[5477]_ ;
  assign \new_[18885]_  = ~\new_[15097]_ ;
  assign \new_[18886]_  = ~\new_[9199]_ ;
  assign \new_[18887]_  = ~\new_[11304]_ ;
  assign \new_[18888]_  = ~\new_[15385]_ ;
  assign \new_[18889]_  = ~\new_[6673]_ ;
  assign \new_[18890]_  = ~\new_[9268]_ ;
  assign \new_[18891]_  = ~\new_[7235]_ ;
  assign \new_[18892]_  = ~\new_[11537]_ ;
  assign \new_[18893]_  = ~\new_[7822]_ ;
  assign \new_[18894]_  = ~\new_[12166]_ ;
  assign \new_[18895]_  = ~\new_[11506]_ ;
  assign \new_[18896]_  = ~\new_[12101]_ ;
  assign \new_[18897]_  = ~\new_[11089]_ ;
  assign \new_[18898]_  = ~\new_[6864]_ ;
  assign \new_[18899]_  = ~\new_[6647]_ ;
  assign \new_[18900]_  = ~\new_[10082]_ ;
  assign \new_[18901]_  = ~\new_[13219]_ ;
  assign \new_[18902]_  = ~\new_[11708]_ ;
  assign \new_[18903]_  = ~\new_[15107]_ ;
  assign \new_[18904]_  = ~\new_[10444]_ ;
  assign \new_[18905]_  = ~\new_[6847]_ ;
  assign \new_[18906]_  = ~\new_[6750]_ ;
  assign \new_[18907]_  = ~\new_[8017]_ ;
  assign \new_[18908]_  = ~\new_[10301]_ ;
  assign \new_[18909]_  = ~\new_[3883]_ ;
  assign \new_[18910]_  = ~\new_[11343]_ ;
  assign \new_[18911]_  = ~\new_[11775]_ ;
  assign \new_[18912]_  = ~\new_[11976]_ ;
  assign \new_[18913]_  = ~\new_[12408]_ ;
  assign \new_[18914]_  = ~\new_[11430]_ ;
  assign n17060 = ~\new_[5058]_ ;
  assign \new_[18916]_  = ~\new_[11731]_ ;
  assign \new_[18917]_  = ~\new_[8212]_ ;
  assign \new_[18918]_  = ~\new_[11840]_ ;
  assign \new_[18919]_  = ~\new_[11845]_ ;
  assign \new_[18920]_  = ~\new_[10344]_ ;
  assign \new_[18921]_  = ~\new_[7465]_ ;
  assign \new_[18922]_  = ~\new_[12329]_ ;
  assign \new_[18923]_  = ~\new_[7861]_ ;
  assign \new_[18924]_  = ~\new_[10117]_ ;
  assign \new_[18925]_  = ~\new_[10093]_ ;
  assign \new_[18926]_  = ~\new_[5099]_ ;
  assign \new_[18927]_  = ~\new_[11511]_ ;
  assign \new_[18928]_  = ~\new_[10364]_ ;
  assign \new_[18929]_  = ~\new_[6915]_ ;
  assign \new_[18930]_  = ~\new_[6598]_ ;
  assign \new_[18931]_  = ~\new_[6841]_ ;
  assign \new_[18932]_  = ~\new_[10103]_ ;
  assign \new_[18933]_  = ~\new_[11847]_ ;
  assign \new_[18934]_  = ~\new_[5106]_ ;
  assign \new_[18935]_  = ~\new_[10338]_ ;
  assign \new_[18936]_  = ~\new_[5491]_ ;
  assign \new_[18937]_  = ~\new_[11474]_ ;
  assign \new_[18938]_  = ~\new_[10302]_ ;
  assign \new_[18939]_  = ~\new_[7439]_ ;
  assign \new_[18940]_  = ~\new_[10083]_ ;
  assign \new_[18941]_  = ~\new_[10342]_ ;
  assign \new_[18942]_  = ~\new_[11319]_ ;
  assign \new_[18943]_  = ~\new_[11286]_ ;
  assign \new_[18944]_  = ~\new_[10090]_ ;
  assign \new_[18945]_  = ~\new_[6631]_ ;
  assign \new_[18946]_  = ~\new_[5025]_ ;
  assign \new_[18947]_  = ~\new_[6838]_ ;
  assign \new_[18948]_  = ~\new_[5490]_ ;
  assign \new_[18949]_  = ~\new_[12261]_ ;
  assign \new_[18950]_  = ~\new_[11272]_ ;
  assign \new_[18951]_  = ~\new_[5019]_ ;
  assign \new_[18952]_  = ~\new_[6784]_ ;
  assign \new_[18953]_  = ~\new_[11325]_ ;
  assign \new_[18954]_  = ~\new_[7257]_ ;
  assign \new_[18955]_  = ~\new_[11532]_ ;
  assign \new_[18956]_  = ~\new_[6590]_ ;
  assign \new_[18957]_  = ~\new_[12150]_ ;
  assign \new_[18958]_  = ~\new_[11787]_ ;
  assign \new_[18959]_  = ~\new_[6804]_ ;
  assign \new_[18960]_  = ~\new_[6698]_ ;
  assign \new_[18961]_  = ~\new_[6919]_ ;
  assign \new_[18962]_  = ~\new_[15594]_ ;
  assign \new_[18963]_  = ~\new_[6728]_ ;
  assign \new_[18964]_  = ~\new_[6940]_ ;
  assign \new_[18965]_  = ~\new_[11640]_ ;
  assign \new_[18966]_  = ~\new_[7501]_ ;
  assign \new_[18967]_  = ~\new_[9193]_ ;
  assign \new_[18968]_  = ~\new_[10413]_ ;
  assign \new_[18969]_  = ~\new_[6736]_ ;
  assign \new_[18970]_  = ~\new_[11564]_ ;
  assign \new_[18971]_  = ~\new_[14861]_ ;
  assign \new_[18972]_  = ~\new_[6668]_ ;
  assign \new_[18973]_  = ~\new_[6609]_ ;
  assign \new_[18974]_  = ~\new_[12137]_ ;
  assign \new_[18975]_  = ~\new_[6876]_ ;
  assign \new_[18976]_  = ~\new_[7415]_ ;
  assign \new_[18977]_  = ~\new_[7492]_ ;
  assign \new_[18978]_  = ~\new_[7964]_ ;
  assign \new_[18979]_  = ~\new_[6867]_ ;
  assign \new_[18980]_  = ~\new_[12167]_ ;
  assign \new_[18981]_  = ~\new_[6849]_ ;
  assign \new_[18982]_  = ~\new_[7249]_ ;
  assign \new_[18983]_  = ~\new_[6875]_ ;
  assign \new_[18984]_  = ~\new_[12322]_ ;
  assign \new_[18985]_  = ~\new_[11806]_ ;
  assign \new_[18986]_  = ~\new_[6710]_ ;
  assign \new_[18987]_  = ~\new_[8211]_ ;
  assign \new_[18988]_  = ~\new_[7259]_ ;
  assign \new_[18989]_  = ~\new_[10154]_ ;
  assign \new_[18990]_  = ~\new_[11570]_ ;
  assign \new_[18991]_  = ~\new_[11541]_ ;
  assign \new_[18992]_  = ~\new_[5487]_ ;
  assign \new_[18993]_  = ~\new_[6939]_ ;
  assign \new_[18994]_  = ~\new_[7921]_ ;
  assign \new_[18995]_  = ~\new_[11403]_ ;
  assign \new_[18996]_  = ~\new_[12161]_ ;
  assign \new_[18997]_  = ~\new_[6831]_ ;
  assign \new_[18998]_  = ~\new_[11442]_ ;
  assign \new_[18999]_  = ~pci_frame_o;
  assign \new_[19000]_  = ~\new_[10309]_ ;
  assign \new_[19001]_  = ~\new_[11859]_ ;
  assign \new_[19002]_  = ~\new_[7247]_ ;
  assign \new_[19003]_  = ~\new_[12475]_ ;
  assign \new_[19004]_  = ~\new_[11759]_ ;
  assign \new_[19005]_  = ~\new_[12195]_ ;
  assign \new_[19006]_  = ~\new_[6807]_ ;
  assign \new_[19007]_  = ~\new_[6692]_ ;
  assign \new_[19008]_  = ~\new_[10232]_ ;
  assign \new_[19009]_  = ~\new_[5497]_ ;
  assign \new_[19010]_  = ~\new_[6909]_ ;
  assign \new_[19011]_  = ~\new_[15417]_ ;
  assign \new_[19012]_  = ~n16740;
  assign \new_[19013]_  = ~\new_[10212]_ ;
  assign \new_[19014]_  = ~\new_[6743]_ ;
  assign \new_[19015]_  = ~\new_[10202]_ ;
  assign \new_[19016]_  = ~\new_[10253]_ ;
  assign \new_[19017]_  = ~\new_[10100]_ ;
  assign \new_[19018]_  = ~\new_[7741]_ ;
  assign \new_[19019]_  = ~\new_[6671]_ ;
  assign \new_[19020]_  = ~\new_[12127]_ ;
  assign \new_[19021]_  = ~\new_[10295]_ ;
  assign \new_[19022]_  = ~\new_[6811]_ ;
  assign \new_[19023]_  = ~\new_[5052]_ ;
  assign \new_[19024]_  = ~\new_[11786]_ ;
  assign \new_[19025]_  = ~\new_[7420]_ ;
  assign \new_[19026]_  = ~\new_[10289]_ ;
  assign \new_[19027]_  = ~\new_[7484]_ ;
  assign \new_[19028]_  = ~\new_[10447]_ ;
  assign \new_[19029]_  = ~\new_[9877]_ ;
  assign \new_[19030]_  = ~\new_[11347]_ ;
  assign \new_[19031]_  = ~\new_[12138]_ ;
  assign \new_[19032]_  = ~\new_[7253]_ ;
  assign \new_[19033]_  = ~\new_[6935]_ ;
  assign \new_[19034]_  = ~\new_[12372]_ ;
  assign \new_[19035]_  = ~\new_[6868]_ ;
  assign \new_[19036]_  = ~\new_[6950]_ ;
  assign \new_[19037]_  = ~\new_[11646]_ ;
  assign \new_[19038]_  = ~\new_[9772]_ ;
  assign \new_[19039]_  = ~\new_[12384]_ ;
  assign \new_[19040]_  = ~\new_[11595]_ ;
  assign n17025 = ~\new_[9633]_ ;
  assign \new_[19042]_  = ~\new_[5489]_ ;
  assign \new_[19043]_  = ~\new_[10120]_ ;
  assign \new_[19044]_  = ~\new_[5474]_ ;
  assign \new_[19045]_  = ~\new_[11752]_ ;
  assign \new_[19046]_  = ~\new_[12382]_ ;
  assign \new_[19047]_  = ~\new_[6987]_ ;
  assign \new_[19048]_  = ~\new_[9591]_ ;
  assign \new_[19049]_  = ~\new_[11995]_ ;
  assign \new_[19050]_  = ~\new_[11804]_ ;
  assign n17075 = ~\new_[9634]_ ;
  assign \new_[19052]_  = ~\new_[7252]_ ;
  assign \new_[19053]_  = ~\new_[6679]_ ;
  assign \new_[19054]_  = ~\new_[10215]_ ;
  assign \new_[19055]_  = ~\new_[6644]_ ;
  assign \new_[19056]_  = ~\new_[7482]_ ;
  assign \new_[19057]_  = ~\new_[6856]_ ;
  assign \new_[19058]_  = ~\new_[8387]_ ;
  assign \new_[19059]_  = ~\new_[6818]_ ;
  assign \new_[19060]_  = ~\new_[12321]_ ;
  assign \new_[19061]_  = ~\new_[6675]_ ;
  assign \new_[19062]_  = ~\new_[10377]_ ;
  assign \new_[19063]_  = ~\new_[7263]_ ;
  assign \new_[19064]_  = ~\new_[11333]_ ;
  assign \new_[19065]_  = ~\new_[6896]_ ;
  assign \new_[19066]_  = ~\new_[6685]_ ;
  assign \new_[19067]_  = ~\new_[11573]_ ;
  assign \new_[19068]_  = ~\new_[11551]_ ;
  assign \new_[19069]_  = ~\new_[9802]_ ;
  assign \new_[19070]_  = ~\new_[5061]_ ;
  assign \new_[19071]_  = ~\new_[10446]_ ;
  assign \new_[19072]_  = ~\new_[11861]_ ;
  assign \new_[19073]_  = ~\new_[6859]_ ;
  assign \new_[19074]_  = ~\new_[15224]_ ;
  assign \new_[19075]_  = ~\new_[5502]_ ;
  assign \new_[19076]_  = ~\new_[12377]_ ;
  assign \new_[19077]_  = ~\new_[4460]_ ;
  assign \new_[19078]_  = ~\new_[12316]_ ;
  assign \new_[19079]_  = ~\new_[6821]_ ;
  assign \new_[19080]_  = ~\new_[7404]_ ;
  assign \new_[19081]_  = ~\new_[12190]_ ;
  assign \new_[19082]_  = ~\new_[10203]_ ;
  assign \new_[19083]_  = ~\new_[5101]_ ;
  assign \new_[19084]_  = ~\new_[11455]_ ;
  assign \new_[19085]_  = ~\new_[6869]_ ;
  assign \new_[19086]_  = ~\new_[6900]_ ;
  assign \new_[19087]_  = ~\new_[6851]_ ;
  assign \new_[19088]_  = ~\new_[8385]_ ;
  assign \new_[19089]_  = ~\new_[6610]_ ;
  assign \new_[19090]_  = ~\new_[12165]_ ;
  assign \new_[19091]_  = ~\new_[7730]_ ;
  assign \new_[19092]_  = ~\new_[6953]_ ;
  assign \new_[19093]_  = ~\new_[11706]_ ;
  assign \new_[19094]_  = ~\new_[7472]_ ;
  assign \new_[19095]_  = ~\new_[11338]_ ;
  assign \new_[19096]_  = ~\new_[11340]_ ;
  assign \new_[19097]_  = ~\new_[6910]_ ;
  assign \new_[19098]_  = ~\new_[12314]_ ;
  assign \new_[19099]_  = ~\new_[11460]_ ;
  assign \new_[19100]_  = ~\new_[12171]_ ;
  assign \new_[19101]_  = ~\new_[6881]_ ;
  assign \new_[19102]_  = ~\new_[12169]_ ;
  assign \new_[19103]_  = ~\new_[6820]_ ;
  assign \new_[19104]_  = ~\new_[11934]_ ;
  assign \new_[19105]_  = ~\new_[12303]_ ;
  assign \new_[19106]_  = ~\new_[6781]_ ;
  assign \new_[19107]_  = ~\new_[6604]_ ;
  assign \new_[19108]_  = ~\new_[10280]_ ;
  assign \new_[19109]_  = ~\new_[6727]_ ;
  assign \new_[19110]_  = ~\new_[6928]_ ;
  assign \new_[19111]_  = ~\new_[5022]_ ;
  assign \new_[19112]_  = ~\new_[12149]_ ;
  assign \new_[19113]_  = ~\new_[6605]_ ;
  assign \new_[19114]_  = ~\new_[10111]_ ;
  assign \new_[19115]_  = ~\new_[12534]_ ;
  assign \new_[19116]_  = ~\new_[3885]_ ;
  assign \new_[19117]_  = ~\new_[10211]_ ;
  assign \new_[19118]_  = ~\new_[6615]_ ;
  assign \new_[19119]_  = ~\new_[11476]_ ;
  assign \new_[19120]_  = ~\new_[10055]_ ;
  assign \new_[19121]_  = ~\new_[10337]_ ;
  assign \new_[19122]_  = ~\new_[11856]_ ;
  assign \new_[19123]_  = ~\new_[9826]_ ;
  assign \new_[19124]_  = ~\new_[10125]_ ;
  assign \new_[19125]_  = ~\new_[7444]_ ;
  assign \new_[19126]_  = ~\new_[9790]_ ;
  assign \new_[19127]_  = ~\new_[11589]_ ;
  assign \new_[19128]_  = ~\new_[11588]_ ;
  assign \new_[19129]_  = ~\new_[11793]_ ;
  assign \new_[19130]_  = ~\new_[11536]_ ;
  assign \new_[19131]_  = ~\new_[11483]_ ;
  assign \new_[19132]_  = ~\new_[8158]_ ;
  assign \new_[19133]_  = ~\new_[11828]_ ;
  assign \new_[19134]_  = ~\new_[12114]_ ;
  assign \new_[19135]_  = ~\new_[11742]_ ;
  assign \new_[19136]_  = ~\new_[5045]_ ;
  assign \new_[19137]_  = ~\new_[10204]_ ;
  assign \new_[19138]_  = ~\new_[10277]_ ;
  assign \new_[19139]_  = ~\new_[9676]_ ;
  assign \new_[19140]_  = ~\new_[15191]_ ;
  assign n17090 = ~\new_[9632]_ ;
  assign \new_[19142]_  = ~\new_[11429]_ ;
  assign \new_[19143]_  = ~\new_[9827]_ ;
  assign \new_[19144]_  = ~\new_[6640]_ ;
  assign \new_[19145]_  = ~\new_[9280]_ ;
  assign \new_[19146]_  = ~\new_[11607]_ ;
  assign \new_[19147]_  = ~\new_[11277]_ ;
  assign \new_[19148]_  = ~\new_[10148]_ ;
  assign \new_[19149]_  = ~\new_[6749]_ ;
  assign \new_[19150]_  = ~\new_[11795]_ ;
  assign \new_[19151]_  = ~\new_[10155]_ ;
  assign \new_[19152]_  = ~\new_[6963]_ ;
  assign \new_[19153]_  = ~\new_[11334]_ ;
  assign \new_[19154]_  = ~\new_[8401]_ ;
  assign \new_[19155]_  = ~\new_[11414]_ ;
  assign \new_[19156]_  = ~\new_[6660]_ ;
  assign \new_[19157]_  = ~\new_[6635]_ ;
  assign \new_[19158]_  = ~\new_[10158]_ ;
  assign \new_[19159]_  = ~pci_gnt_i;
  assign \new_[19160]_  = ~\new_[10159]_ ;
  assign \new_[19161]_  = ~\new_[11291]_ ;
  assign \new_[19162]_  = ~\new_[10160]_ ;
  assign \new_[19163]_  = ~\new_[8200]_ ;
  assign \new_[19164]_  = ~\new_[10267]_ ;
  assign \new_[19165]_  = ~\new_[6674]_ ;
  assign \new_[19166]_  = ~\new_[9631]_ ;
  assign \new_[19167]_  = ~\new_[9630]_ ;
  assign \new_[19168]_  = ~\new_[10164]_ ;
  assign \new_[19169]_  = ~\new_[10166]_ ;
  assign \new_[19170]_  = ~\new_[11488]_ ;
  assign \new_[19171]_  = ~\new_[4980]_ ;
  assign \new_[19172]_  = ~\new_[6588]_ ;
  assign \new_[19173]_  = ~\new_[10936]_ ;
  assign \new_[19174]_  = ~\new_[10255]_ ;
  assign \new_[19175]_  = ~\new_[9985]_ ;
  assign \new_[19176]_  = ~\new_[6883]_ ;
  assign \new_[19177]_  = ~\new_[11709]_ ;
  assign \new_[19178]_  = ~\new_[5021]_ ;
  assign \new_[19179]_  = ~\new_[6678]_ ;
  assign \new_[19180]_  = ~\new_[7260]_ ;
  assign \new_[19181]_  = ~\new_[7747]_ ;
  assign \new_[19182]_  = ~\new_[10174]_ ;
  assign \new_[19183]_  = ~\new_[10085]_ ;
  assign \new_[19184]_  = ~\new_[11542]_ ;
  assign \new_[19185]_  = ~\new_[12334]_ ;
  assign \new_[19186]_  = ~\new_[10260]_ ;
  assign \new_[19187]_  = ~\new_[10445]_ ;
  assign \new_[19188]_  = ~\new_[6652]_ ;
  assign \new_[19189]_  = ~\new_[7777]_ ;
  assign \new_[19190]_  = ~\new_[11562]_ ;
  assign \new_[19191]_  = ~\new_[7965]_ ;
  assign \new_[19192]_  = ~\new_[5888]_ ;
  assign \new_[19193]_  = ~\new_[11136]_ ;
  assign \new_[19194]_  = ~\new_[10368]_ ;
  assign \new_[19195]_  = ~\new_[12160]_ ;
  assign \new_[19196]_  = ~\new_[11659]_ ;
  assign \new_[19197]_  = ~\new_[9767]_ ;
  assign \new_[19198]_  = ~\new_[6772]_ ;
  assign \new_[19199]_  = ~\new_[15392]_ ;
  assign \new_[19200]_  = ~\new_[6687]_ ;
  assign \new_[19201]_  = ~\new_[15015]_ ;
  assign \new_[19202]_  = ~\new_[10176]_ ;
  assign \new_[19203]_  = ~\new_[6703]_ ;
  assign \new_[19204]_  = ~\new_[7433]_ ;
  assign \new_[19205]_  = ~\new_[6927]_ ;
  assign \new_[19206]_  = ~\new_[6829]_ ;
  assign \new_[19207]_  = ~\new_[11558]_ ;
  assign \new_[19208]_  = ~\new_[10200]_ ;
  assign \new_[19209]_  = ~\new_[12177]_ ;
  assign \new_[19210]_  = ~\new_[10254]_ ;
  assign \new_[19211]_  = ~\new_[10251]_ ;
  assign \new_[19212]_  = ~\new_[10250]_ ;
  assign \new_[19213]_  = ~\new_[11736]_ ;
  assign \new_[19214]_  = ~\new_[6903]_ ;
  assign \new_[19215]_  = ~\new_[11745]_ ;
  assign n16755 = ~\new_[11324]_ ;
  assign \new_[19217]_  = ~\new_[10185]_ ;
  assign \new_[19218]_  = ~\new_[10190]_ ;
  assign \new_[19219]_  = ~\new_[3884]_ ;
  assign \new_[19220]_  = ~\new_[11502]_ ;
  assign \new_[19221]_  = ~\new_[11505]_ ;
  assign n17070 = ~\new_[12082]_ ;
  assign \new_[19223]_  = ~\new_[6800]_ ;
  assign \new_[19224]_  = ~\new_[9805]_ ;
  assign \new_[19225]_  = ~\new_[11438]_ ;
  assign \new_[19226]_  = ~\new_[5035]_ ;
  assign \new_[19227]_  = ~\new_[7264]_ ;
  assign \new_[19228]_  = ~\new_[11514]_ ;
  assign \new_[19229]_  = ~\new_[11516]_ ;
  assign \new_[19230]_  = ~\new_[6702]_ ;
  assign \new_[19231]_  = ~\new_[11714]_ ;
  assign \new_[19232]_  = ~\new_[10193]_ ;
  assign \new_[19233]_  = ~\new_[10244]_ ;
  assign \new_[19234]_  = ~\new_[11356]_ ;
  assign \new_[19235]_  = ~\new_[10059]_ ;
  assign \new_[19236]_  = ~\new_[6731]_ ;
  assign \new_[19237]_  = ~\new_[12355]_ ;
  assign \new_[19238]_  = ~\new_[6920]_ ;
  assign \new_[19239]_  = ~\new_[11278]_ ;
  assign \new_[19240]_  = ~\new_[12164]_ ;
  assign \new_[19241]_  = ~\new_[7237]_ ;
  assign \new_[19242]_  = ~\new_[7498]_ ;
  assign \new_[19243]_  = ~\new_[6863]_ ;
  assign \new_[19244]_  = ~\new_[12144]_ ;
  assign \new_[19245]_  = ~\new_[8081]_ ;
  assign \new_[19246]_  = ~\new_[10060]_ ;
  assign \new_[19247]_  = ~\new_[6748]_ ;
  assign \new_[19248]_  = ~\new_[11707]_ ;
  assign \new_[19249]_  = ~\new_[6783]_ ;
  assign \new_[19250]_  = ~\new_[9777]_ ;
  assign \new_[19251]_  = ~\new_[6619]_ ;
  assign \new_[19252]_  = ~\new_[6932]_ ;
  assign \new_[19253]_  = ~\new_[6787]_ ;
  assign \new_[19254]_  = ~\new_[7254]_ ;
  assign \new_[19255]_  = ~\new_[15072]_ ;
  assign \new_[19256]_  = ~\new_[10205]_ ;
  assign \new_[19257]_  = ~\new_[7734]_ ;
  assign \new_[19258]_  = ~\new_[10327]_ ;
  assign \new_[19259]_  = ~\new_[11360]_ ;
  assign \new_[19260]_  = ~\new_[6641]_ ;
  assign \new_[19261]_  = ~\new_[13615]_ ;
  assign \new_[19262]_  = ~\new_[11568]_ ;
  assign \new_[19263]_  = ~\new_[6638]_ ;
  assign n16725 = ~\new_[11094]_ ;
  assign \new_[19265]_  = ~\new_[6649]_ ;
  assign \new_[19266]_  = ~\new_[10145]_ ;
  assign \new_[19267]_  = ~\new_[6861]_ ;
  assign \new_[19268]_  = ~\new_[6794]_ ;
  assign \new_[19269]_  = ~\new_[11554]_ ;
  assign \new_[19270]_  = ~\new_[7477]_ ;
  assign \new_[19271]_  = ~\new_[10213]_ ;
  assign \new_[19272]_  = ~\new_[5109]_ ;
  assign \new_[19273]_  = ~\new_[9191]_ ;
  assign \new_[19274]_  = ~\new_[13628]_ ;
  assign \new_[19275]_  = ~\new_[11322]_ ;
  assign \new_[19276]_  = ~\new_[6733]_ ;
  assign \new_[19277]_  = ~\new_[10877]_ ;
  assign \new_[19278]_  = ~\new_[12247]_ ;
  assign \new_[19279]_  = ~\new_[6663]_ ;
  assign \new_[19280]_  = ~\new_[12251]_ ;
  assign \new_[19281]_  = ~\new_[12243]_ ;
  assign \new_[19282]_  = ~\new_[8262]_ ;
  assign \new_[19283]_  = ~\new_[11302]_ ;
  assign \new_[19284]_  = ~\new_[11518]_ ;
  assign \new_[19285]_  = ~\new_[8694]_ ;
  assign \new_[19286]_  = ~\new_[12090]_ ;
  assign \new_[19287]_  = ~\new_[11365]_ ;
  assign \new_[19288]_  = ~\new_[7935]_ ;
  assign \new_[19289]_  = ~\new_[7844]_ ;
  assign \new_[19290]_  = ~\new_[12091]_ ;
  assign \new_[19291]_  = ~\new_[10142]_ ;
  assign \new_[19292]_  = ~\new_[10278]_ ;
  assign \new_[19293]_  = ~\new_[12308]_ ;
  assign \new_[19294]_  = ~\new_[12371]_ ;
  assign \new_[19295]_  = ~\new_[11408]_ ;
  assign \new_[19296]_  = ~\new_[8691]_ ;
  assign \new_[19297]_  = ~\new_[10228]_ ;
  assign \new_[19298]_  = ~\new_[12498]_ ;
  assign \new_[19299]_  = ~\new_[12093]_ ;
  assign \new_[19300]_  = ~\new_[6870]_ ;
  assign \new_[19301]_  = ~\new_[12254]_ ;
  assign \new_[19302]_  = ~\new_[10225]_ ;
  assign \new_[19303]_  = ~\new_[11423]_ ;
  assign \new_[19304]_  = ~\new_[11424]_ ;
  assign \new_[19305]_  = ~\new_[7009]_ ;
  assign \new_[19306]_  = ~\new_[11132]_ ;
  assign \new_[19307]_  = ~\new_[11688]_ ;
  assign \new_[19308]_  = ~\new_[5781]_ ;
  assign \new_[19309]_  = ~\new_[10115]_ ;
  assign \new_[19310]_  = ~\new_[11755]_ ;
  assign \new_[19311]_  = ~\new_[11444]_ ;
  assign \new_[19312]_  = ~pci_devsel_i;
  assign \new_[19313]_  = ~\new_[7895]_ ;
  assign \new_[19314]_  = ~\new_[11710]_ ;
  assign \new_[19315]_  = ~\new_[11320]_ ;
  assign \new_[19316]_  = ~\new_[11762]_ ;
  assign \new_[19317]_  = ~\new_[10136]_ ;
  assign \new_[19318]_  = ~\new_[5020]_ ;
  assign \new_[19319]_  = ~\new_[11468]_ ;
  assign \new_[19320]_  = ~\new_[6669]_ ;
  assign \new_[19321]_  = ~\new_[5473]_ ;
  assign \new_[19322]_  = ~\new_[11078]_ ;
  assign \new_[19323]_  = ~\new_[11771]_ ;
  assign \new_[19324]_  = ~\new_[11685]_ ;
  assign \new_[19325]_  = ~\new_[11723]_ ;
  assign \new_[19326]_  = ~\new_[11739]_ ;
  assign \new_[19327]_  = ~\new_[11317]_ ;
  assign \new_[19328]_  = ~\new_[11663]_ ;
  assign \new_[19329]_  = ~\new_[11624]_ ;
  assign \new_[19330]_  = ~\new_[11630]_ ;
  assign \new_[19331]_  = ~\new_[7449]_ ;
  assign \new_[19332]_  = ~\new_[6720]_ ;
  assign \new_[19333]_  = ~\new_[11085]_ ;
  assign \new_[19334]_  = ~\new_[10131]_ ;
  assign \new_[19335]_  = ~\new_[6961]_ ;
  assign \new_[19336]_  = ~\new_[8151]_ ;
  assign \new_[19337]_  = ~\new_[7803]_ ;
  assign \new_[19338]_  = ~\new_[6788]_ ;
  assign \new_[19339]_  = ~\new_[11794]_ ;
  assign \new_[19340]_  = ~\new_[11416]_ ;
  assign \new_[19341]_  = ~\new_[5027]_ ;
  assign \new_[19342]_  = ~\new_[10126]_ ;
  assign \new_[19343]_  = ~n16690;
  assign \new_[19344]_  = ~\new_[6756]_ ;
  assign \new_[19345]_  = ~\wbm_adr_o[2] ;
  assign \new_[19346]_  = ~\new_[10878]_ ;
  assign \new_[19347]_  = ~\new_[10239]_ ;
  assign \new_[19348]_  = ~\new_[11389]_ ;
  assign \new_[19349]_  = ~\new_[8217]_ ;
  assign \new_[19350]_  = ~\new_[11393]_ ;
  assign \new_[19351]_  = ~\new_[11553]_ ;
  assign \new_[19352]_  = ~\new_[6835]_ ;
  assign \new_[19353]_  = ~\new_[6734]_ ;
  assign \new_[19354]_  = ~\new_[10290]_ ;
  assign \new_[19355]_  = ~\new_[12201]_ ;
  assign \new_[19356]_  = ~\new_[12083]_ ;
  assign \new_[19357]_  = ~\new_[12112]_ ;
  assign \new_[19358]_  = ~\new_[6763]_ ;
  assign \new_[19359]_  = ~\new_[12235]_ ;
  assign \new_[19360]_  = ~n16745;
  assign \new_[19361]_  = ~\new_[6699]_ ;
  assign \new_[19362]_  = ~\new_[5029]_ ;
  assign \new_[19363]_  = ~\new_[10179]_ ;
  assign \new_[19364]_  = ~\new_[6667]_ ;
  assign \new_[19365]_  = ~\new_[11843]_ ;
  assign \new_[19366]_  = ~\new_[8216]_ ;
  assign \new_[19367]_  = ~\new_[11555]_ ;
  assign \new_[19368]_  = ~\new_[6760]_ ;
  assign \new_[19369]_  = ~\new_[6593]_ ;
  assign \new_[19370]_  = ~\new_[6817]_ ;
  assign \new_[19371]_  = ~\new_[7674]_ ;
  assign \new_[19372]_  = ~\new_[6621]_ ;
  assign \new_[19373]_  = ~\new_[6771]_ ;
  assign \new_[19374]_  = ~\new_[11825]_ ;
  assign \new_[19375]_  = ~\new_[11743]_ ;
  assign \new_[19376]_  = ~\new_[11818]_ ;
  assign \new_[19377]_  = ~\new_[11985]_ ;
  assign \new_[19378]_  = ~\new_[8079]_ ;
  assign \new_[19379]_  = ~\new_[12118]_ ;
  assign \new_[19380]_  = ~\new_[7409]_ ;
  assign \new_[19381]_  = ~\new_[5028]_ ;
  assign \new_[19382]_  = ~\new_[11404]_ ;
  assign \new_[19383]_  = ~\new_[6778]_ ;
  assign \new_[19384]_  = ~\new_[12378]_ ;
  assign \new_[19385]_  = ~\new_[11979]_ ;
  assign \new_[19386]_  = ~\new_[6907]_ ;
  assign \new_[19387]_  = ~\new_[12125]_ ;
  assign \new_[19388]_  = ~\new_[6557]_ ;
  assign \new_[19389]_  = ~\new_[11087]_ ;
  assign \new_[19390]_  = ~\new_[7475]_ ;
  assign \new_[19391]_  = ~\new_[6816]_ ;
  assign \new_[19392]_  = ~\new_[9289]_ ;
  assign \new_[19393]_  = ~\new_[14992]_ ;
  assign \new_[19394]_  = ~\new_[6752]_ ;
  assign \new_[19395]_  = ~\new_[6757]_ ;
  assign \new_[19396]_  = ~\new_[6779]_ ;
  assign \new_[19397]_  = ~\new_[12115]_ ;
  assign \new_[19398]_  = ~\new_[11654]_ ;
  assign \new_[19399]_  = ~\new_[10087]_ ;
  assign \new_[19400]_  = ~\new_[10229]_ ;
  assign \new_[19401]_  = ~\new_[12490]_ ;
  assign \new_[19402]_  = ~\new_[12122]_ ;
  assign \new_[19403]_  = ~\new_[10888]_ ;
  assign \new_[19404]_  = ~\new_[7497]_ ;
  assign \new_[19405]_  = ~\new_[6741]_ ;
  assign \new_[19406]_  = ~\new_[6798]_ ;
  assign \new_[19407]_  = ~\new_[10106]_ ;
  assign \new_[19408]_  = ~\new_[6773]_ ;
  assign \new_[19409]_  = ~\new_[8698]_ ;
  assign \new_[19410]_  = ~\new_[10369]_ ;
  assign \new_[19411]_  = ~\new_[12327]_ ;
  assign \new_[19412]_  = ~\new_[11350]_ ;
  assign \new_[19413]_  = ~\new_[11658]_ ;
  assign \new_[19414]_  = ~\new_[6768]_ ;
  assign \new_[19415]_  = ~\new_[11352]_ ;
  assign \new_[19416]_  = ~\new_[4137]_ ;
  assign \new_[19417]_  = ~\new_[11528]_ ;
  assign \new_[19418]_  = ~\new_[7457]_ ;
  assign \new_[19419]_  = ~\new_[11590]_ ;
  assign \new_[19420]_  = ~\new_[10496]_ ;
  assign \new_[19421]_  = ~\new_[6845]_ ;
  assign \new_[19422]_  = ~\new_[11397]_ ;
  assign \new_[19423]_  = ~\new_[11637]_ ;
  assign \new_[19424]_  = ~\new_[11531]_ ;
  assign \new_[19425]_  = ~\new_[7016]_ ;
  assign \new_[19426]_  = ~\new_[12350]_ ;
  assign \new_[19427]_  = ~\new_[11687]_ ;
  assign \new_[19428]_  = ~\new_[6761]_ ;
  assign \new_[19429]_  = ~\new_[11862]_ ;
  assign \new_[19430]_  = ~\new_[11449]_ ;
  assign \new_[19431]_  = ~\new_[11274]_ ;
  assign \new_[19432]_  = ~\new_[11390]_ ;
  assign \new_[19433]_  = ~\new_[12132]_ ;
  assign \new_[19434]_  = ~\new_[10296]_ ;
  assign \new_[19435]_  = ~\new_[10240]_ ;
  assign \new_[19436]_  = ~\new_[11525]_ ;
  assign \new_[19437]_  = ~\new_[11437]_ ;
  assign \new_[19438]_  = ~\new_[10236]_ ;
  assign \new_[19439]_  = ~\new_[11315]_ ;
  assign \new_[19440]_  = ~\new_[7454]_ ;
  assign \new_[19441]_  = ~\new_[6888]_ ;
  assign \new_[19442]_  = ~\new_[11956]_ ;
  assign \new_[19443]_  = ~\new_[6889]_ ;
  assign \new_[19444]_  = ~\new_[6662]_ ;
  assign \new_[19445]_  = ~\new_[12318]_ ;
  assign \new_[19446]_  = ~\new_[6946]_ ;
  assign \new_[19447]_  = ~\new_[12174]_ ;
  assign \new_[19448]_  = ~\new_[12086]_ ;
  assign \new_[19449]_  = ~\new_[7261]_ ;
  assign \new_[19450]_  = ~\new_[6891]_ ;
  assign \new_[19451]_  = ~\new_[11586]_ ;
  assign \new_[19452]_  = ~\new_[12515]_ ;
  assign \new_[19453]_  = ~\new_[11433]_ ;
  assign \new_[19454]_  = ~\new_[7479]_ ;
  assign \new_[19455]_  = ~\new_[11498]_ ;
  assign \new_[19456]_  = ~\new_[11645]_ ;
  assign \new_[19457]_  = ~\new_[11652]_ ;
  assign \new_[19458]_  = ~\new_[11878]_ ;
  assign \new_[19459]_  = ~\new_[10283]_ ;
  assign \new_[19460]_  = ~\new_[6871]_ ;
  assign \new_[19461]_  = ~\new_[11705]_ ;
  assign \new_[19462]_  = ~\new_[10886]_ ;
  assign \new_[19463]_  = ~\new_[10124]_ ;
  assign \new_[19464]_  = ~\new_[11766]_ ;
  assign \new_[19465]_  = ~\new_[12343]_ ;
  assign \new_[19466]_  = ~\new_[9907]_ ;
  assign \new_[19467]_  = ~\new_[11780]_ ;
  assign \new_[19468]_  = ~\new_[11891]_ ;
  assign \new_[19469]_  = ~\new_[11485]_ ;
  assign \new_[19470]_  = ~\new_[11101]_ ;
  assign \new_[19471]_  = ~\new_[11758]_ ;
  assign \new_[19472]_  = ~\new_[11734]_ ;
  assign \new_[19473]_  = ~\new_[11482]_ ;
  assign \new_[19474]_  = ~\new_[11776]_ ;
  assign \new_[19475]_  = ~\new_[11785]_ ;
  assign \new_[19476]_  = ~\new_[11760]_ ;
  assign \new_[19477]_  = ~\new_[8080]_ ;
  assign \new_[19478]_  = ~\new_[11473]_ ;
  assign \new_[19479]_  = ~\new_[11801]_ ;
  assign \new_[19480]_  = ~\new_[11470]_ ;
  assign \new_[19481]_  = ~\new_[11459]_ ;
  assign \new_[19482]_  = ~\new_[11741]_ ;
  assign \new_[19483]_  = ~\new_[11293]_ ;
  assign \new_[19484]_  = ~\new_[10885]_ ;
  assign \new_[19485]_  = ~\new_[11462]_ ;
  assign \new_[19486]_  = ~\new_[11263]_ ;
  assign \new_[19487]_  = ~\new_[10084]_ ;
  assign \new_[19488]_  = ~\new_[11457]_ ;
  assign \new_[19489]_  = ~\new_[11451]_ ;
  assign \new_[19490]_  = ~\new_[6893]_ ;
  assign \new_[19491]_  = ~\new_[11749]_ ;
  assign \new_[19492]_  = ~\new_[12345]_ ;
  assign \new_[19493]_  = ~\wbs_bte_i[0] ;
  assign \new_[19494]_  = ~\new_[7962]_ ;
  assign \new_[19495]_  = ~\new_[6828]_ ;
  assign \new_[19496]_  = ~\new_[12133]_ ;
  assign \new_[19497]_  = ~\new_[5037]_ ;
  assign \new_[19498]_  = ~\new_[5780]_ ;
  assign \new_[19499]_  = ~\new_[11655]_ ;
  assign \new_[19500]_  = ~\new_[11427]_ ;
  assign \new_[19501]_  = ~\new_[11113]_ ;
  assign \new_[19502]_  = ~\new_[11684]_ ;
  assign \new_[19503]_  = ~\new_[11417]_ ;
  assign \new_[19504]_  = ~\new_[11421]_ ;
  assign \new_[19505]_  = ~\new_[11420]_ ;
  assign \new_[19506]_  = ~\new_[11894]_ ;
  assign \new_[19507]_  = ~\new_[11413]_ ;
  assign \new_[19508]_  = ~\new_[12483]_ ;
  assign \new_[19509]_  = ~\new_[11369]_ ;
  assign \new_[19510]_  = ~\new_[11800]_ ;
  assign \new_[19511]_  = ~\new_[11412]_ ;
  assign \new_[19512]_  = ~\new_[10152]_ ;
  assign \new_[19513]_  = ~\new_[11819]_ ;
  assign \new_[19514]_  = ~\new_[6793]_ ;
  assign \new_[19515]_  = ~\new_[11807]_ ;
  assign \new_[19516]_  = ~\new_[11822]_ ;
  assign \new_[19517]_  = ~\new_[5015]_ ;
  assign \new_[19518]_  = ~\new_[6895]_ ;
  assign \new_[19519]_  = ~\new_[7462]_ ;
  assign \new_[19520]_  = ~\new_[11744]_ ;
  assign \new_[19521]_  = ~\new_[11401]_ ;
  assign \new_[19522]_  = ~\new_[11809]_ ;
  assign \new_[19523]_  = ~\new_[11832]_ ;
  assign \new_[19524]_  = ~\new_[11398]_ ;
  assign \new_[19525]_  = ~\new_[11396]_ ;
  assign \new_[19526]_  = ~\new_[11728]_ ;
  assign \new_[19527]_  = ~\new_[11395]_ ;
  assign \new_[19528]_  = ~\new_[12503]_ ;
  assign \new_[19529]_  = ~\new_[8121]_ ;
  assign \new_[19530]_  = ~\new_[5018]_ ;
  assign \new_[19531]_  = ~\new_[12312]_ ;
  assign \new_[19532]_  = ~\new_[11298]_ ;
  assign \new_[19533]_  = ~\new_[11378]_ ;
  assign \new_[19534]_  = ~\new_[11313]_ ;
  assign \new_[19535]_  = ~\new_[11375]_ ;
  assign \new_[19536]_  = ~\new_[11374]_ ;
  assign \new_[19537]_  = ~\new_[6952]_ ;
  assign \new_[19538]_  = ~\new_[10053]_ ;
  assign \new_[19539]_  = ~\new_[11371]_ ;
  assign \new_[19540]_  = ~\new_[11368]_ ;
  assign \new_[19541]_  = ~\new_[11361]_ ;
  assign \new_[19542]_  = ~\new_[11882]_ ;
  assign \new_[19543]_  = ~\new_[6897]_ ;
  assign \new_[19544]_  = ~\new_[11080]_ ;
  assign \new_[19545]_  = ~\new_[6802]_ ;
  assign \new_[19546]_  = ~\new_[7910]_ ;
  assign \new_[19547]_  = ~\new_[6729]_ ;
  assign \new_[19548]_  = ~\new_[11886]_ ;
  assign \new_[19549]_  = ~\new_[6696]_ ;
  assign \new_[19550]_  = ~\new_[12085]_ ;
  assign \new_[19551]_  = ~\new_[12162]_ ;
  assign n17095 = ~\new_[9141]_ ;
  assign \new_[19553]_  = ~\new_[11563]_ ;
  assign \new_[19554]_  = ~\new_[12139]_ ;
  assign \new_[19555]_  = ~\new_[9282]_ ;
  assign \new_[19556]_  = ~\new_[12196]_ ;
  assign \new_[19557]_  = ~\new_[12148]_ ;
  assign \new_[19558]_  = ~\new_[7507]_ ;
  assign \new_[19559]_  = ~\new_[12493]_ ;
  assign \new_[19560]_  = ~\new_[10150]_ ;
  assign \new_[19561]_  = ~\new_[6634]_ ;
  assign \new_[19562]_  = ~\new_[10058]_ ;
  assign \new_[19563]_  = ~\new_[8207]_ ;
  assign \new_[19564]_  = ~\new_[9138]_ ;
  assign \new_[19565]_  = ~\new_[11683]_ ;
  assign \new_[19566]_  = ~\new_[6850]_ ;
  assign \new_[19567]_  = ~\new_[10008]_ ;
  assign \new_[19568]_  = ~\new_[11989]_ ;
  assign \new_[19569]_  = ~\new_[7900]_ ;
  assign \new_[19570]_  = ~\new_[12153]_ ;
  assign \new_[19571]_  = ~\new_[11697]_ ;
  assign \new_[19572]_  = ~\new_[8690]_ ;
  assign \new_[19573]_  = ~\new_[3886]_ ;
  assign \new_[19574]_  = ~\new_[11860]_ ;
  assign \new_[19575]_  = ~\new_[11287]_ ;
  assign \new_[19576]_  = ~\new_[8214]_ ;
  assign \new_[19577]_  = ~\new_[10195]_ ;
  assign \new_[19578]_  = ~\new_[8271]_ ;
  assign \new_[19579]_  = ~\new_[11798]_ ;
  assign \new_[19580]_  = ~\new_[8055]_ ;
  assign \new_[19581]_  = ~\new_[6832]_ ;
  assign \new_[19582]_  = ~\new_[10153]_ ;
  assign \new_[19583]_  = ~\new_[17047]_ ;
  assign \new_[19584]_  = ~\new_[10246]_ ;
  assign \new_[19585]_  = ~\new_[11349]_ ;
  assign \new_[19586]_  = ~\new_[11718]_ ;
  assign \new_[19587]_  = ~\new_[11512]_ ;
  assign \new_[19588]_  = ~\new_[11633]_ ;
  assign \new_[19589]_  = ~\new_[11290]_ ;
  assign \new_[19590]_  = ~\new_[8400]_ ;
  assign \new_[19591]_  = ~\new_[7648]_ ;
  assign \new_[19592]_  = ~\new_[6739]_ ;
  assign \new_[19593]_  = ~\new_[5496]_ ;
  assign \new_[19594]_  = ~\new_[7256]_ ;
  assign \new_[19595]_  = ~\new_[10086]_ ;
  assign \new_[19596]_  = ~\new_[11307]_ ;
  assign \new_[19597]_  = ~\new_[12273]_ ;
  assign \new_[19598]_  = ~\new_[10247]_ ;
  assign \new_[19599]_  = ~\new_[11702]_ ;
  assign \new_[19600]_  = ~\new_[6914]_ ;
  assign \new_[19601]_  = ~\new_[12317]_ ;
  assign \new_[19602]_  = ~\new_[6684]_ ;
  assign \new_[19603]_  = ~\new_[12111]_ ;
  assign \new_[19604]_  = ~\new_[8221]_ ;
  assign \new_[19605]_  = ~\new_[12192]_ ;
  assign \new_[19606]_  = ~\new_[12332]_ ;
  assign \new_[19607]_  = ~\new_[6842]_ ;
  assign \new_[19608]_  = ~\new_[5100]_ ;
  assign \new_[19609]_  = ~\new_[11661]_ ;
  assign \new_[19610]_  = ~\new_[8219]_ ;
  assign \new_[19611]_  = ~\new_[6682]_ ;
  assign \new_[19612]_  = ~\new_[6814]_ ;
  assign \new_[19613]_  = ~\new_[11797]_ ;
  assign \new_[19614]_  = ~\new_[8693]_ ;
  assign \new_[19615]_  = ~\new_[7255]_ ;
  assign \new_[19616]_  = ~\new_[11082]_ ;
  assign \new_[19617]_  = ~\new_[10177]_ ;
  assign \new_[19618]_  = ~\new_[12113]_ ;
  assign \new_[19619]_  = ~\new_[11584]_ ;
  assign \new_[19620]_  = ~\new_[11668]_ ;
  assign \new_[19621]_  = ~\new_[11854]_ ;
  assign \new_[19622]_  = ~\new_[12143]_ ;
  assign \new_[19623]_  = ~\new_[10258]_ ;
  assign \new_[19624]_  = ~\new_[6747]_ ;
  assign \new_[19625]_  = ~\new_[6633]_ ;
  assign \new_[19626]_  = ~\new_[6586]_ ;
  assign n17005 = ~\new_[9232]_ ;
  assign \new_[19628]_  = ~\new_[11544]_ ;
  assign \new_[19629]_  = ~\new_[11439]_ ;
  assign \new_[19630]_  = ~\new_[7802]_ ;
  assign \new_[19631]_  = ~\new_[11461]_ ;
  assign \new_[19632]_  = ~\new_[11556]_ ;
  assign \new_[19633]_  = ~\new_[11599]_ ;
  assign \new_[19634]_  = ~\new_[15247]_ ;
  assign \new_[19635]_  = ~\new_[6880]_ ;
  assign \new_[19636]_  = ~\new_[5104]_ ;
  assign \new_[19637]_  = ~\new_[11440]_ ;
  assign \new_[19638]_  = ~\new_[11949]_ ;
  assign \new_[19639]_  = ~\new_[5479]_ ;
  assign \new_[19640]_  = ~\new_[9198]_ ;
  assign \new_[19641]_  = ~\new_[12156]_ ;
  assign \new_[19642]_  = ~\new_[12145]_ ;
  assign \new_[19643]_  = ~\new_[10264]_ ;
  assign \new_[19644]_  = ~\new_[11489]_ ;
  assign \new_[19645]_  = ~\new_[6730]_ ;
  assign \new_[19646]_  = ~\new_[12353]_ ;
  assign \new_[19647]_  = ~\new_[9275]_ ;
  assign \new_[19648]_  = ~\new_[6658]_ ;
  assign \new_[19649]_  = ~\new_[7509]_ ;
  assign \new_[19650]_  = ~\new_[10268]_ ;
  assign \new_[19651]_  = ~\new_[11547]_ ;
  assign \new_[19652]_  = ~\new_[6922]_ ;
  assign \new_[19653]_  = ~\new_[10173]_ ;
  assign \new_[19654]_  = ~\new_[11788]_ ;
  assign \new_[19655]_  = ~\new_[7467]_ ;
  assign \new_[19656]_  = ~\new_[7469]_ ;
  assign \new_[19657]_  = ~\new_[6657]_ ;
  assign \new_[19658]_  = ~\new_[6803]_ ;
  assign \new_[19659]_  = ~\new_[6825]_ ;
  assign \new_[19660]_  = ~\new_[12182]_ ;
  assign \new_[19661]_  = ~\new_[12269]_ ;
  assign \new_[19662]_  = ~\new_[7504]_ ;
  assign \new_[19663]_  = ~\new_[10859]_ ;
  assign \new_[19664]_  = ~\new_[6594]_ ;
  assign \new_[19665]_  = ~\new_[6801]_ ;
  assign \new_[19666]_  = ~\new_[11443]_ ;
  assign \new_[19667]_  = ~\new_[12354]_ ;
  assign \new_[19668]_  = ~\new_[6754]_ ;
  assign \new_[19669]_  = ~\new_[10156]_ ;
  assign \new_[19670]_  = ~\new_[10137]_ ;
  assign \new_[19671]_  = ~\new_[10884]_ ;
  assign \new_[19672]_  = ~\new_[10171]_ ;
  assign \new_[19673]_  = ~\new_[10208]_ ;
  assign \new_[19674]_  = ~\new_[11112]_ ;
  assign \new_[19675]_  = ~\new_[11587]_ ;
  assign \new_[19676]_  = ~\new_[11598]_ ;
  assign \new_[19677]_  = ~\new_[6925]_ ;
  assign \new_[19678]_  = ~\new_[10078]_ ;
  assign \new_[19679]_  = ~\new_[10284]_ ;
  assign \new_[19680]_  = ~\new_[6860]_ ;
  assign \new_[19681]_  = ~\new_[11778]_ ;
  assign \new_[19682]_  = ~\new_[10249]_ ;
  assign \new_[19683]_  = ~\new_[8201]_ ;
  assign \new_[19684]_  = ~\new_[9487]_ ;
  assign \new_[19685]_  = ~\new_[10234]_ ;
  assign \new_[19686]_  = ~\new_[10242]_ ;
  assign \new_[19687]_  = ~\new_[7246]_ ;
  assign \new_[19688]_  = ~\new_[12155]_ ;
  assign \new_[19689]_  = ~\new_[6911]_ ;
  assign \new_[19690]_  = ~\new_[10933]_ ;
  assign \new_[19691]_  = ~\new_[12181]_ ;
  assign \new_[19692]_  = ~\new_[8696]_ ;
  assign \new_[19693]_  = ~\new_[6858]_ ;
  assign \new_[19694]_  = ~\new_[11650]_ ;
  assign \new_[19695]_  = ~\new_[11740]_ ;
  assign \new_[19696]_  = ~\new_[7968]_ ;
  assign \new_[19697]_  = ~\new_[6945]_ ;
  assign \new_[19698]_  = ~\new_[11796]_ ;
  assign \new_[19699]_  = ~\new_[6558]_ ;
  assign \new_[19700]_  = ~\new_[6999]_ ;
  assign \new_[19701]_  = ~\new_[11600]_ ;
  assign \new_[19702]_  = ~\new_[11493]_ ;
  assign \new_[19703]_  = ~\new_[11376]_ ;
  assign \new_[19704]_  = ~\new_[10134]_ ;
  assign \new_[19705]_  = ~\new_[11901]_ ;
  assign \new_[19706]_  = ~\new_[11996]_ ;
  assign \new_[19707]_  = ~\new_[6965]_ ;
  assign \new_[19708]_  = ~\new_[11527]_ ;
  assign \new_[19709]_  = ~\new_[10285]_ ;
  assign \new_[19710]_  = ~\new_[10306]_ ;
  assign \new_[19711]_  = ~\new_[11086]_ ;
  assign \new_[19712]_  = ~\new_[7481]_ ;
  assign \new_[19713]_  = ~\new_[11830]_ ;
  assign \new_[19714]_  = ~\new_[6711]_ ;
  assign \new_[19715]_  = ~\new_[12339]_ ;
  assign \new_[19716]_  = ~\new_[10065]_ ;
  assign \new_[19717]_  = ~\new_[12223]_ ;
  assign \new_[19718]_  = ~\new_[6753]_ ;
  assign \new_[19719]_  = ~\new_[7424]_ ;
  assign \new_[19720]_  = ~\new_[11109]_ ;
  assign \new_[19721]_  = ~\new_[5488]_ ;
  assign \new_[19722]_  = ~\new_[6810]_ ;
  assign \new_[19723]_  = ~\new_[12473]_ ;
  assign \new_[19724]_  = ~\new_[10270]_ ;
  assign \new_[19725]_  = ~\new_[10272]_ ;
  assign \new_[19726]_  = ~\new_[10281]_ ;
  assign \new_[19727]_  = ~\new_[6812]_ ;
  assign n17055 = ~\new_[12549]_ ;
  assign \new_[19729]_  = ~\new_[11737]_ ;
  assign \new_[19730]_  = ~\new_[12183]_ ;
  assign \new_[19731]_  = ~\new_[11098]_ ;
  assign \new_[19732]_  = ~\new_[10235]_ ;
  assign \new_[19733]_  = ~\new_[8155]_ ;
  assign \new_[19734]_  = ~\new_[12376]_ ;
  assign \new_[19735]_  = ~\new_[5475]_ ;
  assign \new_[19736]_  = ~\new_[12291]_ ;
  assign \new_[19737]_  = ~\new_[10112]_ ;
  assign \new_[19738]_  = ~\new_[11088]_ ;
  assign \new_[19739]_  = ~\new_[10119]_ ;
  assign \new_[19740]_  = ~\new_[12349]_ ;
  assign \new_[19741]_  = ~\new_[10286]_ ;
  assign \new_[19742]_  = ~\new_[10823]_ ;
  assign \new_[19743]_  = ~\new_[10140]_ ;
  assign \new_[19744]_  = ~\new_[12375]_ ;
  assign \new_[19745]_  = ~\new_[11814]_ ;
  assign \new_[19746]_  = ~\new_[11577]_ ;
  assign \new_[19747]_  = ~\new_[10168]_ ;
  assign \new_[19748]_  = ~\new_[10261]_ ;
  assign \new_[19749]_  = ~\new_[6894]_ ;
  assign \new_[19750]_  = ~\new_[9197]_ ;
  assign \new_[19751]_  = ~\new_[11099]_ ;
  assign \new_[19752]_  = ~\new_[10183]_ ;
  assign \new_[19753]_  = ~\new_[6745]_ ;
  assign \new_[19754]_  = ~\new_[6670]_ ;
  assign \new_[19755]_  = ~\new_[7960]_ ;
  assign \new_[19756]_  = ~\new_[10197]_ ;
  assign \new_[19757]_  = ~\new_[6902]_ ;
  assign n16655 = ~\new_[16179]_ ;
  assign \new_[19759]_  = ~\new_[10051]_ ;
  assign \new_[19760]_  = ~\new_[7500]_ ;
  assign \new_[19761]_  = ~\new_[12347]_ ;
  assign \new_[19762]_  = ~n16935;
  assign \new_[19763]_  = ~\new_[8695]_ ;
  assign \new_[19764]_  = ~\new_[10218]_ ;
  assign \new_[19765]_  = ~\new_[10325]_ ;
  assign \new_[19766]_  = ~\new_[11835]_ ;
  assign \new_[19767]_  = ~\new_[6706]_ ;
  assign \new_[19768]_  = ~\new_[10223]_ ;
  assign \new_[19769]_  = ~\new_[12360]_ ;
  assign \new_[19770]_  = ~\new_[11953]_ ;
  assign \new_[19771]_  = ~\new_[10237]_ ;
  assign \new_[19772]_  = ~\new_[10238]_ ;
  assign \new_[19773]_  = ~\new_[10299]_ ;
  assign \new_[19774]_  = ~\new_[10297]_ ;
  assign \new_[19775]_  = ~\new_[7435]_ ;
  assign \new_[19776]_  = ~\new_[10305]_ ;
  assign \new_[19777]_  = ~\new_[10227]_ ;
  assign \new_[19778]_  = ~\new_[11858]_ ;
  assign \new_[19779]_  = ~\new_[10222]_ ;
  assign \new_[19780]_  = ~\new_[10311]_ ;
  assign \new_[19781]_  = ~\new_[15424]_ ;
  assign \new_[19782]_  = ~\new_[10216]_ ;
  assign \new_[19783]_  = ~\new_[10217]_ ;
  assign \new_[19784]_  = ~\new_[10189]_ ;
  assign \new_[19785]_  = ~\new_[10061]_ ;
  assign \new_[19786]_  = ~\new_[11288]_ ;
  assign \new_[19787]_  = ~\new_[6955]_ ;
  assign \new_[19788]_  = ~\new_[6809]_ ;
  assign \new_[19789]_  = ~\new_[10210]_ ;
  assign \new_[19790]_  = ~\new_[10056]_ ;
  assign \new_[19791]_  = ~\new_[10199]_ ;
  assign \new_[19792]_  = ~\new_[10048]_ ;
  assign \new_[19793]_  = ~\new_[7969]_ ;
  assign \new_[19794]_  = ~\new_[6716]_ ;
  assign \new_[19795]_  = ~\new_[10181]_ ;
  assign \new_[19796]_  = ~\new_[6627]_ ;
  assign \new_[19797]_  = ~\new_[6628]_ ;
  assign \new_[19798]_  = ~\new_[6934]_ ;
  assign \new_[19799]_  = ~\new_[10262]_ ;
  assign \new_[19800]_  = ~\new_[6712]_ ;
  assign \new_[19801]_  = ~\new_[10163]_ ;
  assign \new_[19802]_  = ~\new_[10167]_ ;
  assign \new_[19803]_  = ~\new_[10269]_ ;
  assign \new_[19804]_  = ~\new_[11977]_ ;
  assign \new_[19805]_  = ~\new_[11670]_ ;
  assign \new_[19806]_  = ~\new_[10151]_ ;
  assign \new_[19807]_  = ~\new_[10275]_ ;
  assign \new_[19808]_  = ~\new_[10146]_ ;
  assign \new_[19809]_  = ~\new_[7436]_ ;
  assign \new_[19810]_  = ~\new_[10276]_ ;
  assign \new_[19811]_  = ~\new_[10144]_ ;
  assign \new_[19812]_  = ~\new_[10132]_ ;
  assign \new_[19813]_  = ~\new_[11284]_ ;
  assign \new_[19814]_  = ~\new_[12158]_ ;
  assign \new_[19815]_  = ~\new_[10133]_ ;
  assign \new_[19816]_  = ~\new_[10130]_ ;
  assign \new_[19817]_  = ~\new_[7466]_ ;
  assign \new_[19818]_  = ~\new_[10282]_ ;
  assign \new_[19819]_  = ~\new_[10127]_ ;
  assign \new_[19820]_  = ~\new_[10116]_ ;
  assign \new_[19821]_  = ~\new_[10288]_ ;
  assign \new_[19822]_  = ~\new_[7265]_ ;
  assign \new_[19823]_  = ~\new_[7688]_ ;
  assign \new_[19824]_  = ~\new_[6751]_ ;
  assign \new_[19825]_  = ~\new_[6595]_ ;
  assign \new_[19826]_  = ~\new_[10105]_ ;
  assign \new_[19827]_  = ~\new_[11834]_ ;
  assign \new_[19828]_  = ~\new_[7452]_ ;
  assign n17000 = ~\new_[5059]_ ;
  assign n17045 = ~\new_[9638]_ ;
  assign \new_[19831]_  = ~\new_[11513]_ ;
  assign \new_[19832]_  = ~\new_[6723]_ ;
  assign \new_[19833]_  = ~\new_[10279]_ ;
  assign \new_[19834]_  = ~\new_[6713]_ ;
  assign \new_[19835]_  = ~\new_[11107]_ ;
  assign \new_[19836]_  = ~\new_[11591]_ ;
  assign \new_[19837]_  = ~\new_[11264]_ ;
  assign \new_[19838]_  = ~\new_[10243]_ ;
  assign \new_[19839]_  = ~\new_[12517]_ ;
  assign \new_[19840]_  = ~\new_[7238]_ ;
  assign \new_[19841]_  = ~\new_[12362]_ ;
  assign \new_[19842]_  = ~\new_[7489]_ ;
  assign \new_[19843]_  = ~\new_[12313]_ ;
  assign \new_[19844]_  = ~\new_[5480]_ ;
  assign \new_[19845]_  = ~\new_[5102]_ ;
  assign \new_[19846]_  = ~\new_[7963]_ ;
  assign \new_[19847]_  = ~\new_[11857]_ ;
  assign \new_[19848]_  = ~\new_[11448]_ ;
  assign \new_[19849]_  = ~\new_[5498]_ ;
  assign \new_[19850]_  = ~\new_[11447]_ ;
  assign \new_[19851]_  = ~\new_[11540]_ ;
  assign \new_[19852]_  = ~\new_[7244]_ ;
  assign \new_[19853]_  = ~\new_[6718]_ ;
  assign \new_[19854]_  = ~\new_[6623]_ ;
  assign \new_[19855]_  = ~\new_[6655]_ ;
  assign \new_[19856]_  = ~\new_[11266]_ ;
  assign \new_[19857]_  = ~\new_[8226]_ ;
  assign \new_[19858]_  = ~\new_[6956]_ ;
  assign \new_[19859]_  = ~\new_[10074]_ ;
  assign \new_[19860]_  = ~\new_[11824]_ ;
  assign \new_[19861]_  = ~\new_[12089]_ ;
  assign \new_[19862]_  = ~\new_[11724]_ ;
  assign \new_[19863]_  = ~\new_[10188]_ ;
  assign \new_[19864]_  = ~\new_[10220]_ ;
  assign \new_[19865]_  = ~\new_[10349]_ ;
  assign \new_[19866]_  = ~\new_[11585]_ ;
  assign \new_[19867]_  = ~\new_[6921]_ ;
  assign \new_[19868]_  = ~\new_[11321]_ ;
  assign \new_[19869]_  = ~\new_[5049]_ ;
  assign \new_[19870]_  = ~\new_[7243]_ ;
  assign \new_[19871]_  = ~\new_[11735]_ ;
  assign \new_[19872]_  = ~\new_[10381]_ ;
  assign \new_[19873]_  = ~\new_[19874]_ ;
  assign \new_[19874]_  = \new_[20285]_ ;
  assign \new_[19875]_  = \new_[20478]_ ;
  assign \new_[19876]_  = \new_[19881]_ ;
  assign \new_[19877]_  = ~\new_[19880]_ ;
  assign \new_[19878]_  = \new_[19880]_ ;
  assign \new_[19879]_  = ~\new_[19877]_ ;
  assign \new_[19880]_  = ~\new_[19881]_ ;
  assign \new_[19881]_  = ~\new_[8557]_ ;
  assign \new_[19882]_  = \new_[14874]_ ;
  assign \new_[19883]_  = ~\new_[20425]_  | ~\new_[20407]_ ;
  assign \new_[19884]_  = \new_[15041]_  & \new_[19908]_ ;
  assign \new_[19885]_  = \new_[18458]_  | \new_[19909]_ ;
  assign \new_[19886]_  = ~\new_[20454]_  & ~\new_[19901]_ ;
  assign \new_[19887]_  = ~\new_[20318]_  | ~\new_[20347]_ ;
  assign \new_[19888]_  = ~\new_[19889]_  | ~\new_[5295]_  | ~\new_[20543]_ ;
  assign \new_[19889]_  = ~\new_[20542]_ ;
  assign \new_[19890]_  = ~\new_[19883]_  | ~\new_[17947]_ ;
  assign \new_[19891]_  = ~\new_[20302]_  & ~\new_[17251]_ ;
  assign \new_[19892]_  = ~\new_[20177]_  & ~\new_[20305]_ ;
  assign \new_[19893]_  = ~\new_[20201]_  | ~\new_[19939]_ ;
  assign n780 = ~\new_[19899]_  | (~\new_[19895]_  & ~\new_[20313]_ );
  assign \new_[19895]_  = ~\new_[3948]_  & (~\new_[5299]_  | ~\wbm_dat_o[10] );
  assign \new_[19896]_  = ~\new_[19897]_ ;
  assign \new_[19897]_  = ~\new_[11175]_  | ~\new_[11137]_ ;
  assign n9175 = ~\new_[13629]_  | ~\new_[13845]_  | ~\new_[13705]_ ;
  assign \new_[19899]_  = ~\new_[5631]_  | ~\wbm_dat_o[10] ;
  assign \new_[19900]_  = ~\new_[9269]_ ;
  assign \new_[19901]_  = \new_[20301]_  | \new_[20300]_ ;
  assign \new_[19902]_  = ~\new_[19937]_ ;
  assign \new_[19903]_  = ~\new_[20127]_  & ~\new_[20159]_ ;
  assign \new_[19904]_  = ~\new_[6327]_ ;
  assign \new_[19905]_  = ~\new_[9878]_ ;
  assign \new_[19906]_  = ~\new_[19907]_  | ~\new_[11075]_ ;
  assign \new_[19907]_  = \new_[20090]_  & \new_[20089]_ ;
  assign \new_[19908]_  = ~\new_[19907]_ ;
  assign \new_[19909]_  = ~\new_[20509]_  | ~\new_[20479]_ ;
  assign \new_[19910]_  = ~\new_[19911]_  | ~\new_[20155]_ ;
  assign \new_[19911]_  = ~\new_[20302]_ ;
  assign \new_[19912]_  = ~\new_[20162]_ ;
  assign \new_[19913]_  = ~\new_[14893]_  | ~\new_[16832]_ ;
  assign \new_[19914]_  = ~\new_[20031]_  | ~\new_[19913]_ ;
  assign n16500 = ~\new_[19930]_ ;
  assign \new_[19916]_  = ~\new_[19917]_  | ~\new_[11890]_ ;
  assign \new_[19917]_  = ~\new_[19918]_  & ~\new_[20536]_ ;
  assign \new_[19918]_  = ~wbs_stb_i;
  assign \new_[19919]_  = ~\new_[19900]_  | ~\new_[20523]_  | ~\new_[19204]_ ;
  assign \new_[19920]_  = ~\new_[19921]_  & ~\new_[20127]_  & ~\new_[20130]_ ;
  assign \new_[19921]_  = ~\new_[16372]_  | ~\new_[17032]_ ;
  assign \new_[19922]_  = ~\new_[10382]_ ;
  assign \new_[19923]_  = ~\new_[10383]_ ;
  assign \new_[19924]_  = ~\new_[19949]_  | ~\new_[20511]_ ;
  assign \new_[19925]_  = \new_[20095]_  & \new_[19926]_ ;
  assign \new_[19926]_  = ~\new_[19959]_ ;
  assign \new_[19927]_  = ~\new_[19928]_  | ~\new_[15919]_ ;
  assign \new_[19928]_  = ~\new_[11332]_  & ~\new_[15411]_ ;
  assign \new_[19929]_  = \new_[19927]_ ;
  assign \new_[19930]_  = ~\new_[15411]_ ;
  assign \new_[19931]_  = ~\new_[20466]_  | ~\new_[19932]_ ;
  assign \new_[19932]_  = ~\new_[19933]_  & ~\new_[19934]_ ;
  assign \new_[19933]_  = ~\new_[3995]_  | ~\new_[4009]_  | ~\new_[17957]_ ;
  assign \new_[19934]_  = \new_[19909]_ ;
  assign \new_[19935]_  = ~\new_[19936]_  | ~\new_[14250]_  | ~\new_[20466]_ ;
  assign \new_[19936]_  = ~\new_[19934]_ ;
  assign \new_[19937]_  = ~n17010 | ~\new_[20201]_  | ~\new_[19939]_ ;
  assign \new_[19938]_  = \new_[9647]_  & \new_[9618]_ ;
  assign \new_[19939]_  = ~\new_[16990]_  | ~\new_[20550]_ ;
  assign \new_[19940]_  = ~\new_[20206]_  | ~\new_[20204]_ ;
  assign \new_[19941]_  = ~\new_[20415]_ ;
  assign \new_[19942]_  = ~\new_[19945]_  & (~\new_[19887]_  | ~\new_[19943]_ );
  assign \new_[19943]_  = ~\new_[19944]_  & ~\new_[17181]_ ;
  assign \new_[19944]_  = ~\new_[12039]_  | ~\new_[13869]_  | ~\new_[16852]_  | ~\new_[19201]_ ;
  assign \new_[19945]_  = ~\new_[16516]_  | ~\new_[15891]_ ;
  assign \new_[19946]_  = \new_[16852]_  & \new_[12039]_ ;
  assign \new_[19947]_  = \new_[13869]_  & \new_[19887]_ ;
  assign \new_[19948]_  = ~\new_[15015]_  & ~\new_[17181]_ ;
  assign \new_[19949]_  = ~\new_[19950]_  | ~\new_[19952]_ ;
  assign \new_[19950]_  = ~\new_[19951]_  | ~\new_[20510]_ ;
  assign \new_[19951]_  = ~\new_[19916]_  | ~\new_[19919]_ ;
  assign \new_[19952]_  = ~\new_[6327]_  | ~\new_[20479]_  | ~\new_[20534]_ ;
  assign \new_[19953]_  = ~\new_[19954]_  | ~\new_[20510]_ ;
  assign \new_[19954]_  = ~\new_[19916]_  | ~\new_[19919]_ ;
  assign \new_[19955]_  = ~\new_[19958]_  & ~\new_[19965]_ ;
  assign \new_[19956]_  = \new_[19886]_  & \new_[16617]_ ;
  assign \new_[19957]_  = \new_[19886]_  & \new_[16617]_ ;
  assign \new_[19958]_  = ~\new_[19885]_  | ~\new_[14874]_  | ~\new_[20172]_ ;
  assign \new_[19959]_  = \new_[17045]_  & \new_[20284]_ ;
  assign \new_[19960]_  = \new_[20197]_  & \new_[20473]_ ;
  assign \new_[19961]_  = ~\new_[20285]_  | ~\new_[19902]_ ;
  assign \new_[19962]_  = ~\new_[19963]_  & ~\new_[19964]_ ;
  assign \new_[19963]_  = ~\new_[20212]_ ;
  assign \new_[19964]_  = ~\new_[19893]_  & (~\new_[20198]_  | ~\new_[20211]_ );
  assign \new_[19965]_  = ~\new_[20118]_  | ~\new_[20111]_ ;
  assign \new_[19966]_  = ~\new_[20159]_  & ~\new_[20127]_ ;
  assign \new_[19967]_  = ~\new_[20069]_ ;
  assign \new_[19968]_  = ~\new_[19969]_  & ~\new_[19972]_ ;
  assign \new_[19969]_  = ~\new_[19971]_  & (~\new_[9488]_  | ~\new_[19970]_ );
  assign \new_[19970]_  = ~\new_[19942]_  & ~\new_[19941]_ ;
  assign \new_[19971]_  = ~\new_[19970]_  & ~\new_[9276]_ ;
  assign \new_[19972]_  = ~\new_[9919]_  | ~\new_[9915]_ ;
  assign \new_[19973]_  = ~\new_[19969]_ ;
  assign \new_[19974]_  = ~\new_[19975]_ ;
  assign \new_[19975]_  = ~\new_[19941]_  & ~\new_[19942]_ ;
  assign n2845 = ~\new_[19977]_  | ~\new_[19978]_ ;
  assign \new_[19977]_  = ~\new_[6985]_  & ~\new_[8327]_ ;
  assign \new_[19978]_  = ~\new_[19979]_ ;
  assign \new_[19979]_  = ~\new_[19985]_  | ~\new_[19982]_  | ~\new_[19980]_  | ~\new_[19981]_ ;
  assign \new_[19980]_  = (~\new_[18532]_  | ~\new_[9299]_ ) & (~\new_[9290]_  | ~\new_[19107]_ );
  assign \new_[19981]_  = (~\new_[18385]_  | ~\new_[20001]_ ) & (~\new_[19999]_  | ~\new_[19677]_ );
  assign \new_[19982]_  = ~\new_[20551]_  | ~\new_[19984]_ ;
  assign \new_[19983]_  = \new_[20193]_  & \new_[20470]_ ;
  assign \new_[19984]_  = ~\new_[6901]_ ;
  assign \new_[19985]_  = ~\new_[19986]_  | ~\new_[19988]_ ;
  assign \new_[19986]_  = \new_[19987]_ ;
  assign \new_[19987]_  = \new_[20470]_  & \new_[9691]_ ;
  assign \new_[19988]_  = ~\new_[6854]_ ;
  assign \new_[19989]_  = ~\new_[19990]_  & (~\new_[11031]_  | ~\new_[20506]_ );
  assign \new_[19990]_  = ~\new_[19991]_  | ~\new_[19992]_ ;
  assign \new_[19991]_  = (~\new_[17677]_  | ~\new_[20375]_ ) & (~\new_[20092]_  | ~\new_[12030]_ );
  assign \new_[19992]_  = ~\new_[19993]_  & (~\new_[20056]_  | ~\new_[12047]_ );
  assign \new_[19993]_  = \new_[20049]_  & \new_[10405]_ ;
  assign n2815 = \new_[7403]_  | \new_[20005]_ ;
  assign \new_[19995]_  = (~\new_[19996]_  & ~\new_[6681]_ ) | (~\new_[20468]_  & ~\new_[7239]_ );
  assign \new_[19996]_  = ~\new_[19997]_ ;
  assign \new_[19997]_  = \new_[19998]_ ;
  assign \new_[19998]_  = \new_[20471]_  & \new_[9683]_ ;
  assign \new_[19999]_  = ~\new_[20469]_ ;
  assign \new_[20000]_  = ~\new_[7239]_ ;
  assign \new_[20001]_  = ~\new_[19996]_ ;
  assign \new_[20002]_  = ~\new_[6681]_ ;
  assign \new_[20003]_  = ~\new_[20190]_  | ~\new_[20392]_ ;
  assign \new_[20004]_  = ~\new_[20466]_  | ~\new_[20441]_ ;
  assign \new_[20005]_  = ~\new_[20014]_  | ~\new_[20006]_  | ~\new_[20009]_ ;
  assign \new_[20006]_  = ~\new_[20007]_  & ~\new_[19995]_ ;
  assign \new_[20007]_  = ~\new_[20008]_  | ~\new_[9156]_ ;
  assign \new_[20008]_  = ~\new_[9299]_  | ~\new_[19203]_ ;
  assign \new_[20009]_  = ~\new_[20010]_  & (~\new_[9290]_  | ~\new_[18573]_ );
  assign \new_[20010]_  = ~\new_[9157]_  | (~\new_[20011]_  & ~\new_[6964]_ );
  assign \new_[20011]_  = ~\new_[20012]_ ;
  assign \new_[20012]_  = \new_[20013]_ ;
  assign \new_[20013]_  = \new_[9690]_  & \new_[9683]_ ;
  assign \new_[20014]_  = ~\new_[20015]_  & (~\new_[20518]_  | ~\new_[18117]_ );
  assign \new_[20015]_  = ~\new_[8610]_  | ~\new_[8310]_ ;
  assign \new_[20016]_  = ~\new_[6964]_ ;
  assign \new_[20017]_  = ~\new_[15027]_  & ~\new_[20018]_ ;
  assign \new_[20018]_  = ~\new_[20025]_  | ~\new_[20019]_  | ~\new_[20024]_ ;
  assign \new_[20019]_  = ~\new_[20020]_  & (~\new_[20049]_  | ~\new_[10406]_ );
  assign \new_[20020]_  = ~\new_[20021]_  | ~\new_[20022]_ ;
  assign \new_[20021]_  = (~\new_[11958]_  | ~\new_[19957]_ ) & (~\new_[12017]_  | ~\new_[20298]_ );
  assign \new_[20022]_  = ~\new_[20158]_  | ~\new_[20023]_ ;
  assign \new_[20023]_  = \new_[10526]_  & \new_[10499]_ ;
  assign \new_[20024]_  = ~\new_[15888]_  | ~\new_[10406]_ ;
  assign \new_[20025]_  = ~\new_[20494]_  | ~\new_[10526]_ ;
  assign \new_[20026]_  = \new_[20027]_  & \new_[20029]_ ;
  assign \new_[20027]_  = ~\new_[20028]_  | (~\new_[9643]_  & ~\new_[16611]_ );
  assign \new_[20028]_  = \new_[14614]_  & \new_[19930]_ ;
  assign \new_[20029]_  = \new_[19913]_  & \new_[20030]_ ;
  assign \new_[20030]_  = \new_[17549]_  | \new_[17098]_ ;
  assign \new_[20031]_  = ~\new_[20028]_  | (~\new_[9643]_  & ~\new_[16611]_ );
  assign \new_[20032]_  = ~\new_[20033]_  & (~\new_[20506]_  | ~\new_[11046]_ );
  assign \new_[20033]_  = ~\new_[20034]_  | ~\new_[20035]_ ;
  assign \new_[20034]_  = ~\new_[20092]_  | ~\new_[12304]_ ;
  assign \new_[20035]_  = ~\new_[20036]_  & (~\new_[20494]_  | ~\new_[10846]_ );
  assign \new_[20036]_  = ~\new_[20037]_ ;
  assign \new_[20037]_  = ~\new_[20450]_  | ~\new_[10003]_ ;
  assign \new_[20038]_  = ~\new_[19931]_ ;
  assign \new_[20039]_  = ~\new_[20466]_ ;
  assign \new_[20040]_  = ~\new_[20516]_  | ~\new_[20513]_ ;
  assign \new_[20041]_  = ~\new_[10383]_  & ~\new_[10382]_ ;
  assign \new_[20042]_  = ~\new_[10384]_  | ~\new_[10385]_ ;
  assign \new_[20043]_  = \new_[20041]_ ;
  assign \new_[20044]_  = ~\new_[20524]_  & ~\new_[20119]_ ;
  assign \new_[20045]_  = ~\new_[20046]_  & (~\new_[10869]_  | ~\new_[20506]_ );
  assign \new_[20046]_  = ~\new_[20051]_  | ~\new_[20047]_  | ~\new_[20050]_ ;
  assign \new_[20047]_  = ~\new_[20048]_  & (~\new_[20056]_  | ~\new_[12046]_ );
  assign \new_[20048]_  = \new_[20049]_  & \new_[10395]_ ;
  assign \new_[20049]_  = \new_[20069]_  & \new_[20162]_ ;
  assign \new_[20050]_  = ~\new_[20375]_  | ~\new_[17718]_ ;
  assign \new_[20051]_  = ~\new_[20092]_  | ~\new_[12409]_ ;
  assign \new_[20052]_  = ~\new_[20053]_ ;
  assign \new_[20053]_  = ~\new_[20055]_  | ~\new_[20374]_  | ~\new_[20054]_ ;
  assign \new_[20054]_  = ~\new_[20092]_  | ~\new_[12414]_ ;
  assign \new_[20055]_  = ~\new_[20056]_  | ~\new_[12045]_ ;
  assign \new_[20056]_  = \new_[20057]_ ;
  assign \new_[20057]_  = \new_[20058]_  & \new_[20059]_ ;
  assign \new_[20058]_  = ~\new_[20066]_  & ~\new_[20304]_ ;
  assign \new_[20059]_  = ~\new_[20454]_  & ~\new_[19901]_ ;
  assign \new_[20060]_  = ~\new_[20061]_  | ~\new_[20062]_ ;
  assign \new_[20061]_  = ~\new_[16580]_  & (~\new_[16955]_  | ~\new_[9801]_ );
  assign \new_[20062]_  = ~\new_[16358]_  & ~\new_[16359]_ ;
  assign \new_[20063]_  = ~\new_[20103]_  & ~\new_[20064]_ ;
  assign \new_[20064]_  = \new_[9903]_  | \new_[10870]_ ;
  assign \new_[20065]_  = ~\new_[10870]_ ;
  assign \new_[20066]_  = ~\new_[15097]_  | ~\new_[18903]_ ;
  assign \new_[20067]_  = ~\new_[20068]_  | ~\new_[20127]_ ;
  assign \new_[20068]_  = ~\new_[20159]_ ;
  assign \new_[20069]_  = ~\new_[20066]_  & ~\new_[20070]_ ;
  assign \new_[20070]_  = ~\new_[20068]_  | ~\new_[20127]_ ;
  assign \new_[20071]_  = ~\new_[20070]_ ;
  assign \new_[20072]_  = ~\new_[20066]_ ;
  assign \new_[20073]_  = \new_[20074]_ ;
  assign \new_[20074]_  = ~\new_[20075]_  | ~\new_[20079]_ ;
  assign \new_[20075]_  = ~\new_[20078]_  | ~\new_[20076]_  | ~\new_[20077]_ ;
  assign \new_[20076]_  = ~\new_[9615]_ ;
  assign \new_[20077]_  = \new_[13858]_  & \new_[15921]_ ;
  assign \new_[20078]_  = ~\new_[15833]_ ;
  assign \new_[20079]_  = ~\new_[20080]_  | ~\new_[20082]_ ;
  assign \new_[20080]_  = ~\new_[20081]_ ;
  assign \new_[20081]_  = ~\new_[17012]_  & ~\new_[16890]_ ;
  assign \new_[20082]_  = pci_frame_i ? \new_[11332]_  : \new_[9617]_ ;
  assign \new_[20083]_  = ~\new_[20084]_  & ~\new_[15833]_ ;
  assign \new_[20084]_  = ~\new_[20076]_ ;
  assign \new_[20085]_  = ~\new_[15019]_  & ~\new_[20434]_ ;
  assign \new_[20086]_  = ~\new_[15417]_  & ~\new_[10380]_ ;
  assign \new_[20087]_  = ~\new_[15199]_ ;
  assign \new_[20088]_  = \new_[15041]_  | \new_[10380]_ ;
  assign \new_[20089]_  = ~\new_[15199]_  & ~\new_[15417]_ ;
  assign \new_[20090]_  = ~\new_[20154]_  & ~\new_[20529]_ ;
  assign \new_[20091]_  = (~\new_[12306]_  | ~\new_[20092]_ ) & (~\new_[20094]_  | ~\new_[11047]_ );
  assign \new_[20092]_  = \new_[20093]_ ;
  assign \new_[20093]_  = \new_[19892]_  & \new_[19891]_ ;
  assign \new_[20094]_  = ~\new_[20160]_  & ~\new_[20177]_  & ~\new_[20454]_  & ~\new_[20159]_ ;
  assign \new_[20095]_  = ~\new_[20283]_ ;
  assign \new_[20096]_  = ~\new_[20226]_  | ~\new_[20383]_ ;
  assign \new_[20097]_  = ~\new_[20282]_  & ~\new_[20380]_ ;
  assign \new_[20098]_  = \new_[16356]_  & \new_[16357]_ ;
  assign \new_[20099]_  = \new_[15863]_  & \new_[16352]_ ;
  assign \new_[20100]_  = \new_[20465]_ ;
  assign \new_[20101]_  = ~\new_[15177]_ ;
  assign n16635 = \new_[20103]_ ;
  assign \new_[20103]_  = \new_[20104]_ ;
  assign \new_[20104]_  = ~\new_[20152]_  | ~\new_[20105]_ ;
  assign \new_[20105]_  = ~\new_[13158]_ ;
  assign \new_[20106]_  = \new_[20404]_  & \new_[20096]_ ;
  assign \new_[20107]_  = ~\new_[4040]_  & ~\new_[20108]_ ;
  assign \new_[20108]_  = ~\new_[4041]_ ;
  assign \new_[20109]_  = ~\new_[20115]_  | ~\new_[20110]_  | ~\new_[20114]_ ;
  assign \new_[20110]_  = \new_[20111]_  & \new_[20113]_ ;
  assign \new_[20111]_  = ~\new_[20166]_  | ~\new_[20112]_ ;
  assign \new_[20112]_  = ~\new_[10366]_ ;
  assign \new_[20113]_  = ~\new_[17653]_  | ~\new_[15016]_ ;
  assign \new_[20114]_  = \new_[14874]_  & \new_[19885]_ ;
  assign \new_[20115]_  = ~\new_[20164]_ ;
  assign \new_[20116]_  = ~\new_[20117]_ ;
  assign \new_[20117]_  = ~\new_[20172]_  | ~\new_[20165]_  | ~\new_[20171]_ ;
  assign \new_[20118]_  = ~\new_[17653]_  | ~\new_[15016]_ ;
  assign \new_[20119]_  = \new_[20166]_ ;
  assign \new_[20120]_  = ~\new_[20168]_  | ~\new_[20169]_ ;
  assign \new_[20121]_  = \new_[20122]_  & \new_[20129]_ ;
  assign \new_[20122]_  = ~\new_[20123]_  | ~\new_[20124]_ ;
  assign \new_[20123]_  = ~\new_[16829]_  | ~\new_[16372]_  | ~\new_[17033]_ ;
  assign \new_[20124]_  = ~\new_[20128]_  | ~\new_[20127]_  | ~\new_[20125]_  | ~\new_[20126]_ ;
  assign \new_[20125]_  = \new_[16828]_  & \new_[17265]_ ;
  assign \new_[20126]_  = ~\new_[20488]_  & ~\new_[17748]_ ;
  assign \new_[20127]_  = ~\new_[13222]_ ;
  assign \new_[20128]_  = \new_[15097]_ ;
  assign \new_[20129]_  = ~\new_[20130]_ ;
  assign \new_[20130]_  = ~\new_[14614]_  | ~\new_[15497]_  | ~\new_[20421]_ ;
  assign \new_[20131]_  = ~\new_[20128]_ ;
  assign n2515 = ~\new_[20139]_  | ~\new_[20133]_  | ~\new_[20137]_ ;
  assign \new_[20133]_  = ~\new_[20134]_  & ~\new_[20135]_ ;
  assign \new_[20134]_  = ~\new_[7317]_  | ~\new_[6366]_ ;
  assign \new_[20135]_  = ~\new_[7119]_  | ~\new_[6048]_  | ~\new_[20136]_  | ~\new_[6458]_ ;
  assign \new_[20136]_  = ~\new_[7386]_  | ~\new_[19534]_ ;
  assign \new_[20137]_  = ~\new_[6046]_  & ~\new_[20138]_ ;
  assign \new_[20138]_  = ~\new_[5824]_ ;
  assign \new_[20139]_  = ~\new_[6290]_  & ~\new_[6045]_ ;
  assign \new_[20140]_  = ~\new_[15175]_  | ~\new_[15216]_ ;
  assign \new_[20141]_  = ~\new_[20142]_ ;
  assign \new_[20142]_  = \new_[14867]_  & \new_[15177]_ ;
  assign \new_[20143]_  = ~\new_[15175]_ ;
  assign \new_[20144]_  = ~\new_[20335]_  | ~\new_[20458]_ ;
  assign \new_[20145]_  = \new_[20146]_  & \new_[10870]_ ;
  assign \new_[20146]_  = ~\new_[9903]_  & ~\new_[20104]_ ;
  assign \new_[20147]_  = ~\new_[20151]_  & (~\new_[20148]_  | ~\new_[20149]_ );
  assign \new_[20148]_  = \new_[20088]_  & \new_[16599]_ ;
  assign \new_[20149]_  = ~\new_[20087]_  | ~\new_[20040]_  | ~\new_[20150]_  | ~\new_[20086]_ ;
  assign \new_[20150]_  = \new_[20041]_  & \new_[20042]_ ;
  assign \new_[20151]_  = \new_[20152]_ ;
  assign \new_[20152]_  = ~\new_[11075]_ ;
  assign \new_[20153]_  = ~\new_[20151]_ ;
  assign \new_[20154]_  = ~\new_[20150]_ ;
  assign \new_[20155]_  = ~\new_[20304]_ ;
  assign \new_[20156]_  = ~\new_[20157]_  | ~\new_[15216]_ ;
  assign \new_[20157]_  = ~\new_[15177]_ ;
  assign \new_[20158]_  = ~\new_[20160]_  & ~\new_[17450]_  & ~\new_[20159]_  & ~\new_[20303]_ ;
  assign \new_[20159]_  = \new_[14993]_ ;
  assign \new_[20160]_  = \new_[20127]_  | \new_[20066]_ ;
  assign \new_[20161]_  = ~\new_[20159]_  & ~\new_[20160]_ ;
  assign \new_[20162]_  = ~\new_[20303]_  & ~\new_[17450]_ ;
  assign \new_[20163]_  = ~\new_[14993]_ ;
  assign \new_[20164]_  = ~\new_[20165]_  | ~\new_[20170]_ ;
  assign \new_[20165]_  = ~\new_[20166]_ ;
  assign \new_[20166]_  = ~\new_[20167]_ ;
  assign \new_[20167]_  = ~\new_[20168]_  | ~\new_[20169]_ ;
  assign \new_[20168]_  = ~\new_[19953]_  | ~\new_[19952]_ ;
  assign \new_[20169]_  = \new_[20479]_  & \new_[20534]_ ;
  assign \new_[20170]_  = \new_[20171]_  & \new_[20172]_ ;
  assign \new_[20171]_  = ~\new_[11328]_  & ~\new_[20403]_ ;
  assign \new_[20172]_  = ~\new_[17151]_  | ~\new_[17577]_ ;
  assign \new_[20173]_  = ~\new_[14991]_ ;
  assign \new_[20174]_  = ~\new_[20338]_ ;
  assign \new_[20175]_  = ~\new_[20176]_  & ~\new_[20067]_  & ~\new_[20066]_ ;
  assign \new_[20176]_  = \new_[20454]_  | \new_[20177]_ ;
  assign \new_[20177]_  = ~\new_[17748]_  | ~\new_[20300]_ ;
  assign \new_[20178]_  = ~\new_[20176]_ ;
  assign \new_[20179]_  = ~\new_[14991]_  | ~\new_[15216]_  | ~\new_[20142]_  | ~\new_[15393]_ ;
  assign \new_[20180]_  = ~\new_[15182]_  & ~\new_[20181]_ ;
  assign \new_[20181]_  = ~\new_[20182]_  | ~\new_[15092]_ ;
  assign \new_[20182]_  = ~\new_[15181]_ ;
  assign \new_[20183]_  = \new_[19927]_  & \new_[15092]_ ;
  assign \new_[20184]_  = ~\new_[15182]_  & ~\new_[15181]_ ;
  assign \new_[20185]_  = ~\new_[20186]_  | ~\new_[20410]_ ;
  assign \new_[20186]_  = ~\new_[20187]_  | ~\new_[20192]_ ;
  assign \new_[20187]_  = ~\new_[20411]_ ;
  assign \new_[20188]_  = ~\new_[8599]_ ;
  assign \new_[20189]_  = ~\new_[8202]_ ;
  assign \new_[20190]_  = ~\new_[20191]_ ;
  assign \new_[20191]_  = \new_[20188]_  ? \new_[20440]_  : \new_[20189]_ ;
  assign \new_[20192]_  = \new_[20412]_ ;
  assign \new_[20193]_  = ~\new_[20474]_  & ~\new_[20472]_ ;
  assign \new_[20194]_  = \new_[20478]_  | \new_[9626]_ ;
  assign \new_[20195]_  = ~\new_[20196]_  | ~\new_[20478]_ ;
  assign \new_[20196]_  = ~\new_[9641]_ ;
  assign \new_[20197]_  = ~\new_[20472]_ ;
  assign \new_[20198]_  = \new_[20207]_  & \new_[20550]_ ;
  assign \new_[20199]_  = \new_[20546]_ ;
  assign \new_[20200]_  = ~\new_[20109]_  | ~\new_[20444]_ ;
  assign \new_[20201]_  = ~\new_[20550]_  | ~\new_[20202]_  | ~\new_[20206]_ ;
  assign \new_[20202]_  = ~\new_[4042]_  & ~\new_[20203]_ ;
  assign \new_[20203]_  = ~\new_[20204]_  | ~\new_[20205]_ ;
  assign \new_[20204]_  = \new_[19938]_  & \new_[9619]_ ;
  assign \new_[20205]_  = ~\new_[18523]_  & ~wbm_ack_i & ~wbm_err_i;
  assign \new_[20206]_  = ~\new_[17540]_  & ~\new_[16908]_ ;
  assign \new_[20207]_  = ~\new_[4042]_ ;
  assign n3000 = ~\new_[20217]_  | ~\new_[20214]_  | ~\new_[20209]_  | ~\new_[20213]_ ;
  assign \new_[20209]_  = ~\new_[20212]_  | ~\new_[20210]_  | ~\new_[20211]_ ;
  assign \new_[20210]_  = ~\new_[14934]_  | ~\new_[19874]_ ;
  assign \new_[20211]_  = ~\new_[17180]_ ;
  assign \new_[20212]_  = ~\new_[10375]_  & ~\new_[17250]_ ;
  assign \new_[20213]_  = ~\new_[20212]_  | (~\new_[14933]_  & ~\new_[15857]_ );
  assign \new_[20214]_  = ~\new_[20215]_  & (~\new_[15624]_  | ~\new_[16603]_ );
  assign \new_[20215]_  = ~\new_[20216]_ ;
  assign \new_[20216]_  = ~\new_[20407]_  | ~\new_[20497]_ ;
  assign \new_[20217]_  = ~\new_[17752]_  | ~\new_[20499]_  | ~\new_[20407]_ ;
  assign \new_[20218]_  = ~\new_[20212]_ ;
  assign n1160 = ~\new_[20220]_  | ~\new_[20222]_ ;
  assign \new_[20220]_  = ~\new_[4332]_  & ~\new_[20221]_ ;
  assign \new_[20221]_  = ~\new_[4829]_  | ~\new_[4666]_ ;
  assign \new_[20222]_  = ~\new_[20223]_  & ~\new_[4249]_ ;
  assign \new_[20223]_  = ~\new_[4743]_  | ~\new_[4744]_ ;
  assign \new_[20224]_  = ~\new_[5054]_ ;
  assign \new_[20225]_  = ~\new_[17064]_ ;
  assign \new_[20226]_  = ~\new_[20224]_  | ~\new_[20225]_ ;
  assign \new_[20227]_  = ~\new_[20156]_  & ~\new_[20339]_ ;
  assign \new_[20228]_  = ~\new_[20231]_  | ~\new_[20541]_  | ~\new_[20539]_ ;
  assign \new_[20229]_  = ~\new_[4981]_ ;
  assign \new_[20230]_  = ~\new_[5107]_ ;
  assign \new_[20231]_  = ~\new_[20544]_ ;
  assign n1155 = ~\new_[20233]_  | ~\new_[20236]_ ;
  assign \new_[20233]_  = ~\new_[20234]_  & ~\new_[20235]_ ;
  assign \new_[20234]_  = ~\new_[4848]_  | ~\new_[4735]_ ;
  assign \new_[20235]_  = ~\new_[4513]_  | ~\new_[4514]_ ;
  assign \new_[20236]_  = ~\new_[20237]_  & ~\new_[20238]_ ;
  assign \new_[20237]_  = ~\new_[4737]_  | ~\new_[4736]_ ;
  assign \new_[20238]_  = ~\new_[4827]_  | ~\new_[4664]_ ;
  assign n1210 = ~\new_[20240]_  | ~\new_[20242]_ ;
  assign \new_[20240]_  = ~\new_[20241]_ ;
  assign \new_[20241]_  = ~\new_[4702]_  | ~\new_[4640]_  | ~\new_[4701]_  | ~\new_[4480]_ ;
  assign \new_[20242]_  = ~\new_[20243]_ ;
  assign \new_[20243]_  = ~\new_[4641]_  | ~\new_[4808]_  | ~\new_[4549]_  | ~\new_[4548]_ ;
  assign n1240 = ~\new_[20249]_  | ~\new_[20245]_  | ~\new_[20248]_ ;
  assign \new_[20245]_  = ~\new_[20246]_  & ~\new_[20247]_ ;
  assign \new_[20246]_  = ~\new_[4559]_  | ~\new_[4558]_ ;
  assign \new_[20247]_  = ~\new_[4490]_  | ~\new_[4489]_ ;
  assign \new_[20248]_  = \new_[4814]_  & \new_[4649]_ ;
  assign \new_[20249]_  = ~\new_[20250]_ ;
  assign \new_[20250]_  = ~\new_[4712]_  | ~\new_[4713]_ ;
  assign n1315 = ~\new_[20258]_  | ~\new_[20252]_  | ~\new_[20255]_ ;
  assign \new_[20252]_  = ~\new_[20253]_  & ~\new_[20254]_ ;
  assign \new_[20253]_  = ~\new_[4589]_  | ~\new_[4588]_ ;
  assign \new_[20254]_  = ~\new_[4524]_  | ~\new_[4523]_ ;
  assign \new_[20255]_  = ~\new_[20256]_  & ~\new_[20257]_ ;
  assign \new_[20256]_  = ~\new_[4832]_ ;
  assign \new_[20257]_  = ~\new_[4669]_ ;
  assign \new_[20258]_  = ~\new_[20259]_ ;
  assign \new_[20259]_  = ~\new_[4749]_  | ~\new_[4750]_ ;
  assign n1350 = ~\new_[20265]_  | ~\new_[20261]_  | ~\new_[20262]_ ;
  assign \new_[20261]_  = \new_[4473]_  & \new_[4472]_ ;
  assign \new_[20262]_  = ~\new_[20263]_  & ~\new_[20264]_ ;
  assign \new_[20263]_  = ~\new_[4691]_  | ~\new_[4692]_ ;
  assign \new_[20264]_  = ~\new_[4636]_  | ~\new_[4804]_ ;
  assign \new_[20265]_  = ~\new_[20266]_ ;
  assign \new_[20266]_  = ~\new_[4689]_  | ~\new_[4690]_ ;
  assign n1355 = ~\new_[20272]_  | ~\new_[20268]_  | ~\new_[20269]_ ;
  assign \new_[20268]_  = \new_[4479]_  & \new_[4478]_ ;
  assign \new_[20269]_  = ~\new_[20270]_  & ~\new_[20271]_ ;
  assign \new_[20270]_  = ~\new_[4699]_  | ~\new_[4700]_ ;
  assign \new_[20271]_  = ~\new_[4639]_  | ~\new_[4807]_ ;
  assign \new_[20272]_  = ~\new_[20273]_ ;
  assign \new_[20273]_  = ~\new_[4697]_  | ~\new_[4698]_ ;
  assign n1360 = ~\new_[20279]_  | ~\new_[20275]_  | ~\new_[20276]_ ;
  assign \new_[20275]_  = \new_[4529]_  & \new_[4528]_ ;
  assign \new_[20276]_  = ~\new_[20277]_  & ~\new_[20278]_ ;
  assign \new_[20277]_  = ~\new_[4755]_  | ~\new_[4756]_ ;
  assign \new_[20278]_  = ~\new_[4673]_  | ~\new_[4835]_ ;
  assign \new_[20279]_  = ~\new_[20280]_ ;
  assign \new_[20280]_  = ~\new_[4753]_  | ~\new_[4754]_ ;
  assign \new_[20281]_  = ~\new_[20282]_  & ~\new_[20283]_ ;
  assign \new_[20282]_  = ~\new_[10374]_  | ~\new_[19905]_ ;
  assign \new_[20283]_  = ~\new_[17045]_  & ~\new_[20284]_ ;
  assign \new_[20284]_  = ~\new_[5053]_ ;
  assign \new_[20285]_  = ~\new_[20286]_  | ~\new_[20427]_ ;
  assign \new_[20286]_  = ~\new_[20406]_  | ~\new_[20287]_ ;
  assign \new_[20287]_  = \new_[20550]_  & \new_[20107]_ ;
  assign \new_[20288]_  = ~\new_[8389]_ ;
  assign \new_[20289]_  = ~\new_[20200]_  | ~\new_[20466]_ ;
  assign \new_[20290]_  = ~\new_[20291]_  | ~\new_[20294]_ ;
  assign \new_[20291]_  = ~\new_[20292]_  & ~\new_[20293]_ ;
  assign \new_[20292]_  = ~\new_[15164]_  & ~\new_[15398]_ ;
  assign \new_[20293]_  = ~\new_[16779]_ ;
  assign \new_[20294]_  = ~\new_[20295]_ ;
  assign \new_[20295]_  = ~\new_[16960]_  | ~\new_[16959]_  | ~\new_[17146]_  | ~\new_[16965]_ ;
  assign \new_[20296]_  = ~\new_[15164]_ ;
  assign \new_[20297]_  = ~\new_[15398]_ ;
  assign \new_[20298]_  = ~\new_[20302]_  & ~\new_[20299]_  & ~\new_[20127]_  & ~\new_[20163]_ ;
  assign \new_[20299]_  = ~\new_[14992]_  | ~\new_[20491]_  | ~\new_[20300]_  | ~\new_[20301]_ ;
  assign \new_[20300]_  = ~\new_[15105]_ ;
  assign \new_[20301]_  = ~\new_[14209]_ ;
  assign \new_[20302]_  = ~\new_[18885]_  | ~\new_[18903]_ ;
  assign \new_[20303]_  = ~\new_[20300]_  | ~\new_[20301]_ ;
  assign \new_[20304]_  = \new_[20127]_  | \new_[20163]_ ;
  assign \new_[20305]_  = ~\new_[20489]_  | ~\new_[14992]_ ;
  assign n830 = ~\new_[20307]_  | ~\new_[20308]_ ;
  assign \new_[20307]_  = ~\new_[5632]_  | ~\wbm_dat_o[22] ;
  assign \new_[20308]_  = ~\new_[20309]_  | ~\new_[20314]_ ;
  assign \new_[20309]_  = ~\new_[20310]_  | (~\new_[5416]_  & ~\new_[4022]_ );
  assign \new_[20310]_  = ~\new_[5299]_  | ~\wbm_dat_o[22] ;
  assign \new_[20311]_  = ~\new_[20312]_  | ~\new_[17947]_ ;
  assign \new_[20312]_  = \new_[9982]_  | \new_[5886]_ ;
  assign \new_[20313]_  = ~\new_[20314]_ ;
  assign \new_[20314]_  = ~\new_[20315]_ ;
  assign \new_[20315]_  = ~\new_[19896]_  | ~n3000;
  assign \new_[20316]_  = ~\new_[20314]_ ;
  assign \new_[20317]_  = ~\new_[20311]_ ;
  assign \new_[20318]_  = ~\new_[20321]_  & (~\new_[20319]_  | ~\new_[20320]_ );
  assign \new_[20319]_  = \new_[20352]_  & \new_[20173]_ ;
  assign \new_[20320]_  = ~\new_[20341]_  | (~\new_[20140]_  & ~\new_[20141]_ );
  assign \new_[20321]_  = ~\new_[19927]_  | ~\new_[20179]_  | ~\new_[20180]_ ;
  assign \new_[20322]_  = \new_[20323]_  & \new_[20390]_ ;
  assign \new_[20323]_  = \new_[20463]_  & \new_[20461]_ ;
  assign \new_[20324]_  = ~\new_[20467]_  | ~\new_[20466]_ ;
  assign \new_[20325]_  = ~\new_[20331]_  | (~\new_[20326]_  & ~\new_[20330]_ );
  assign \new_[20326]_  = \new_[20327]_  & \new_[20328]_ ;
  assign \new_[20327]_  = ~\new_[9998]_  | ~\new_[16179]_  | ~\new_[12370]_  | ~\new_[16411]_ ;
  assign \new_[20328]_  = \new_[13795]_  | \new_[15859]_  | \new_[20329]_  | \new_[17476]_ ;
  assign \new_[20329]_  = \new_[20156]_ ;
  assign \new_[20330]_  = ~\new_[16207]_  | ~\new_[16572]_ ;
  assign \new_[20331]_  = \new_[19929]_  | \new_[16207]_ ;
  assign \new_[20332]_  = ~\new_[20327]_ ;
  assign \new_[20333]_  = ~\new_[8092]_  | ~\new_[20336]_ ;
  assign \new_[20334]_  = ~\new_[20344]_  | ~\new_[20335]_ ;
  assign \new_[20335]_  = \new_[20462]_  & \new_[20346]_ ;
  assign \new_[20336]_  = ~\new_[10883]_ ;
  assign \new_[20337]_  = \new_[20338]_  & \new_[15393]_ ;
  assign \new_[20338]_  = \new_[15216]_  | \new_[20339]_ ;
  assign \new_[20339]_  = ~\new_[14867]_ ;
  assign \new_[20340]_  = ~\new_[20341]_ ;
  assign \new_[20341]_  = ~\new_[20339]_ ;
  assign \new_[20342]_  = ~\new_[20408]_  | ~\new_[15191]_ ;
  assign \new_[20343]_  = ~\new_[20344]_  | ~\new_[20345]_ ;
  assign \new_[20344]_  = ~\new_[20392]_  & ~\new_[20190]_ ;
  assign \new_[20345]_  = \new_[20463]_  & \new_[20346]_ ;
  assign \new_[20346]_  = \new_[8201]_  ? \new_[20324]_  : \new_[8200]_ ;
  assign \new_[20347]_  = ~\new_[20354]_  | ~\new_[20348]_  | ~\new_[20353]_ ;
  assign \new_[20348]_  = ~\new_[20352]_  | ~\new_[20349]_  | ~\new_[20351]_ ;
  assign \new_[20349]_  = ~\new_[20142]_  | ~\new_[20350]_ ;
  assign \new_[20350]_  = ~\new_[20140]_ ;
  assign \new_[20351]_  = ~\new_[20227]_ ;
  assign \new_[20352]_  = ~\new_[15393]_ ;
  assign \new_[20353]_  = ~\new_[20337]_  | ~\new_[20349]_ ;
  assign \new_[20354]_  = \new_[14991]_  ? \new_[15393]_  : \new_[20173]_ ;
  assign \new_[20355]_  = ~\new_[20356]_  & ~\new_[20360]_ ;
  assign \new_[20356]_  = ~\new_[7227]_  | ~\new_[20357]_  | ~\new_[20358]_ ;
  assign \new_[20357]_  = ~\new_[6157]_ ;
  assign \new_[20358]_  = ~\new_[20359]_  & ~\new_[6160]_ ;
  assign \new_[20359]_  = ~\new_[7226]_ ;
  assign \new_[20360]_  = ~\new_[20361]_ ;
  assign \new_[20361]_  = ~\new_[6159]_  & ~\new_[6158]_ ;
  assign \new_[20362]_  = ~\new_[20363]_  & ~\new_[20365]_ ;
  assign \new_[20363]_  = ~\new_[20364]_  | ~\new_[6281]_ ;
  assign \new_[20364]_  = ~\new_[6011]_ ;
  assign \new_[20365]_  = ~\new_[7308]_  | ~\new_[20366]_  | ~\new_[20367]_ ;
  assign \new_[20366]_  = ~\new_[6013]_ ;
  assign \new_[20367]_  = ~\new_[6010]_  & ~\new_[6012]_ ;
  assign \new_[20368]_  = ~\new_[20369]_  & ~\new_[20370]_ ;
  assign \new_[20369]_  = ~\new_[6286]_  | ~\new_[6379]_ ;
  assign \new_[20370]_  = ~\new_[20373]_  | ~\new_[20371]_  | ~\new_[20372]_ ;
  assign \new_[20371]_  = ~\new_[6074]_  & ~\new_[6249]_ ;
  assign \new_[20372]_  = ~\new_[6073]_ ;
  assign \new_[20373]_  = ~\new_[6072]_ ;
  assign \new_[20374]_  = ~\new_[20375]_  | ~\new_[20378]_ ;
  assign \new_[20375]_  = ~\new_[20376]_ ;
  assign \new_[20376]_  = ~\new_[19966]_  | ~\new_[20072]_  | ~\new_[20377]_ ;
  assign \new_[20377]_  = ~\new_[20454]_  & ~\new_[20303]_ ;
  assign \new_[20378]_  = \new_[10509]_  & \new_[10516]_ ;
  assign \new_[20379]_  = ~\new_[20380]_  & ~\new_[20381]_ ;
  assign \new_[20380]_  = \new_[17045]_  & \new_[20284]_ ;
  assign \new_[20381]_  = ~\new_[20382]_  & (~\new_[20225]_  | ~\new_[20224]_ );
  assign \new_[20382]_  = ~\new_[20383]_ ;
  assign \new_[20383]_  = ~\new_[5054]_  | ~\new_[17064]_ ;
  assign \new_[20384]_  = \new_[20385]_ ;
  assign \new_[20385]_  = ~\new_[20386]_  | ~\new_[20389]_ ;
  assign \new_[20386]_  = \new_[20387]_  | \new_[20388]_ ;
  assign \new_[20387]_  = ~\new_[13648]_  | ~\new_[13818]_ ;
  assign \new_[20388]_  = ~\new_[13716]_  | ~\new_[16687]_ ;
  assign \new_[20389]_  = ~\new_[20525]_  | ~\new_[13716]_  | ~\new_[19955]_ ;
  assign \new_[20390]_  = ~\new_[20391]_  & ~\new_[20392]_ ;
  assign \new_[20391]_  = \new_[20188]_  ? \new_[20440]_  : \new_[20189]_ ;
  assign \new_[20392]_  = ~\new_[20393]_  | ~\new_[20464]_ ;
  assign \new_[20393]_  = ~\new_[20004]_  | ~\new_[18680]_ ;
  assign \new_[20394]_  = \new_[20395]_  | \new_[20400]_ ;
  assign \new_[20395]_  = ~\new_[20398]_  | ~\new_[20396]_  | ~\new_[20397]_ ;
  assign \new_[20396]_  = ~\new_[11328]_  & ~\new_[16602]_ ;
  assign \new_[20397]_  = \new_[14874]_  & \new_[20172]_ ;
  assign \new_[20398]_  = \new_[20399]_ ;
  assign \new_[20399]_  = ~\new_[4009]_  & ~\new_[17567]_ ;
  assign \new_[20400]_  = ~\new_[20401]_  & ~\new_[20402]_ ;
  assign \new_[20401]_  = \new_[13716]_  & \new_[13208]_ ;
  assign \new_[20402]_  = ~\new_[5297]_  & ~\new_[12542]_ ;
  assign \new_[20403]_  = ~\new_[20399]_ ;
  assign \new_[20404]_  = \new_[20405]_  ? \new_[5055]_  : \new_[17081]_ ;
  assign \new_[20405]_  = ~\new_[17081]_ ;
  assign \new_[20406]_  = ~\new_[20435]_  | ~\new_[20407]_ ;
  assign \new_[20407]_  = \new_[20408]_ ;
  assign \new_[20408]_  = \new_[17263]_  & \new_[18615]_ ;
  assign \new_[20409]_  = ~\new_[20410]_  | ~\new_[20411]_ ;
  assign \new_[20410]_  = ~\new_[20145]_  & ~\new_[20147]_ ;
  assign \new_[20411]_  = ~\new_[20063]_  | ~\new_[20060]_ ;
  assign \new_[20412]_  = ~\new_[16685]_  | ~\new_[16840]_ ;
  assign \new_[20413]_  = \new_[20414]_ ;
  assign \new_[20414]_  = ~\new_[20415]_  | ~\new_[20421]_ ;
  assign \new_[20415]_  = ~\new_[20419]_  | ~\new_[20416]_  | ~\new_[20417]_ ;
  assign \new_[20416]_  = ~\new_[16593]_  & (~\new_[16875]_  | ~n17185);
  assign \new_[20417]_  = ~\new_[20418]_  & (~\new_[16850]_  | ~n17160);
  assign \new_[20418]_  = ~n17185 & ~\new_[16875]_ ;
  assign \new_[20419]_  = ~\new_[20420]_  & (~\new_[16964]_  | ~n17360);
  assign \new_[20420]_  = ~n17160 & ~\new_[16850]_ ;
  assign \new_[20421]_  = \new_[16878]_  & \new_[19781]_ ;
  assign \new_[20422]_  = ~\new_[20404]_  | ~\new_[20379]_  | ~\new_[20281]_ ;
  assign \new_[20423]_  = \new_[17319]_  & \new_[20439]_ ;
  assign \new_[20424]_  = \new_[9878]_ ;
  assign \new_[20425]_  = ~\new_[20426]_ ;
  assign \new_[20426]_  = ~\new_[20424]_  | ~\new_[20422]_  | ~\new_[20439]_ ;
  assign \new_[20427]_  = ~\new_[7266]_  & (~\new_[20433]_  | ~\new_[20428]_ );
  assign \new_[20428]_  = \new_[20429]_  & \new_[20430]_ ;
  assign \new_[20429]_  = ~\new_[20342]_  & ~\new_[20438]_ ;
  assign \new_[20430]_  = ~\new_[20431]_  | ~\new_[20432]_ ;
  assign \new_[20431]_  = ~\new_[15019]_  & ~\new_[15007]_ ;
  assign \new_[20432]_  = ~\new_[20290]_  | ~\new_[15612]_ ;
  assign \new_[20433]_  = ~\new_[20436]_  | ~\new_[20437]_ ;
  assign \new_[20434]_  = ~\new_[20432]_ ;
  assign \new_[20435]_  = ~\new_[20437]_  | ~\new_[20436]_ ;
  assign \new_[20436]_  = ~\new_[4042]_  | ~\new_[20424]_  | ~\new_[20422]_  | ~\new_[20423]_ ;
  assign \new_[20437]_  = ~\new_[20496]_  | ~\new_[20439]_ ;
  assign \new_[20438]_  = ~\new_[20096]_  | ~\new_[20404]_  | ~\new_[20097]_  | ~\new_[20095]_ ;
  assign \new_[20439]_  = ~\new_[14278]_ ;
  assign \new_[20440]_  = ~\new_[20441]_  | ~\new_[20466]_ ;
  assign \new_[20441]_  = ~\new_[20442]_  | ~\new_[20443]_ ;
  assign \new_[20442]_  = ~\new_[14250]_  | ~\new_[20038]_ ;
  assign \new_[20443]_  = ~\new_[20111]_  | ~\new_[20118]_  | ~\new_[20114]_  | ~\new_[20116]_ ;
  assign \new_[20444]_  = ~\new_[14250]_  | ~\new_[20038]_ ;
  assign \new_[20445]_  = ~\new_[20446]_  & ~\new_[20447]_ ;
  assign \new_[20446]_  = \new_[9625]_  ? \new_[20478]_  : \new_[9628]_ ;
  assign \new_[20447]_  = \new_[9565]_  ? \new_[20478]_  : \new_[9616]_ ;
  assign \new_[20448]_  = ~\new_[20447]_ ;
  assign \new_[20449]_  = ~\new_[20446]_ ;
  assign \new_[20450]_  = \new_[20451]_  & \new_[20455]_ ;
  assign \new_[20451]_  = ~\new_[20452]_ ;
  assign \new_[20452]_  = ~\new_[20453]_  | ~\new_[17385]_  | ~\new_[17474]_ ;
  assign \new_[20453]_  = ~\new_[20454]_ ;
  assign \new_[20454]_  = ~\new_[14992]_  | ~\new_[20492]_ ;
  assign \new_[20455]_  = ~\new_[20066]_  & ~\new_[20304]_ ;
  assign \new_[20456]_  = ~\new_[17385]_  | ~\new_[17474]_ ;
  assign \new_[20457]_  = ~\new_[20458]_  | ~\new_[20459]_ ;
  assign \new_[20458]_  = \new_[20392]_  & \new_[20391]_ ;
  assign \new_[20459]_  = ~\new_[20460]_ ;
  assign \new_[20460]_  = ~\new_[20461]_  | ~\new_[20462]_ ;
  assign \new_[20461]_  = \new_[19683]_  ? \new_[20324]_  : \new_[19163]_ ;
  assign \new_[20462]_  = \new_[8389]_  ? \new_[20289]_  : \new_[8203]_ ;
  assign \new_[20463]_  = \new_[20288]_  ? \new_[20289]_  : \new_[18027]_ ;
  assign \new_[20464]_  = ~\new_[20465]_  | ~\new_[18185]_ ;
  assign \new_[20465]_  = ~\new_[20039]_  & (~\new_[20444]_  | ~\new_[20109]_ );
  assign \new_[20466]_  = ~\new_[20098]_  | ~\new_[20099]_ ;
  assign \new_[20467]_  = ~\new_[20444]_  | ~\new_[20109]_ ;
  assign \new_[20468]_  = \new_[20469]_ ;
  assign \new_[20469]_  = ~\new_[20470]_  | ~\new_[20471]_ ;
  assign \new_[20470]_  = ~\new_[20449]_  & ~\new_[20448]_ ;
  assign \new_[20471]_  = \new_[20472]_  & \new_[20473]_ ;
  assign \new_[20472]_  = ~\new_[20194]_  | ~\new_[20195]_ ;
  assign \new_[20473]_  = ~\new_[20474]_ ;
  assign \new_[20474]_  = \new_[20475]_  ? \new_[20477]_  : \new_[20476]_ ;
  assign \new_[20475]_  = ~\new_[9627]_ ;
  assign \new_[20476]_  = ~\new_[9678]_ ;
  assign \new_[20477]_  = ~\new_[20412]_  | ~\new_[20409]_ ;
  assign \new_[20478]_  = ~\new_[20409]_  | ~\new_[20412]_ ;
  assign \new_[20479]_  = \new_[6163]_ ;
  assign \new_[20480]_  = ~\new_[20483]_ ;
  assign \new_[20481]_  = ~\new_[20483]_ ;
  assign \new_[20482]_  = ~\new_[20483]_ ;
  assign \new_[20483]_  = ~\new_[20484]_ ;
  assign \new_[20484]_  = ~\new_[9200]_ ;
  assign \new_[20485]_  = ~\new_[20486]_ ;
  assign \new_[20486]_  = ~\new_[16794]_ ;
  assign \new_[20487]_  = ~\new_[20488]_ ;
  assign \new_[20488]_  = \new_[20489]_ ;
  assign \new_[20489]_  = ~\new_[20490]_ ;
  assign \new_[20490]_  = \new_[20492]_ ;
  assign \new_[20491]_  = ~\new_[20492]_ ;
  assign \new_[20492]_  = ~\new_[15120]_ ;
  assign \new_[20493]_  = ~\new_[9491]_ ;
  assign \new_[20494]_  = ~\new_[20495]_ ;
  assign \new_[20495]_  = ~\new_[20175]_ ;
  assign \new_[20496]_  = ~\new_[20438]_ ;
  assign \new_[20497]_  = ~\new_[20499]_ ;
  assign \new_[20498]_  = ~\new_[20497]_ ;
  assign \new_[20499]_  = \new_[20438]_ ;
  assign \new_[20500]_  = \new_[10380]_ ;
  assign \new_[20501]_  = ~\new_[20502]_ ;
  assign \new_[20502]_  = ~\new_[20504]_ ;
  assign \new_[20503]_  = \new_[20504]_ ;
  assign \new_[20504]_  = ~\new_[9273]_ ;
  assign \new_[20505]_  = \new_[19887]_ ;
  assign \new_[20506]_  = ~\new_[20507]_ ;
  assign \new_[20507]_  = ~\new_[20094]_ ;
  assign \new_[20508]_  = ~\new_[20509]_ ;
  assign \new_[20509]_  = \new_[11890]_ ;
  assign \new_[20510]_  = \new_[20535]_  & \new_[6163]_ ;
  assign \new_[20511]_  = \new_[20533]_  & \new_[6163]_ ;
  assign \new_[20512]_  = ~\new_[20513]_ ;
  assign \new_[20513]_  = ~\new_[10385]_ ;
  assign \new_[20514]_  = ~\new_[20515]_ ;
  assign \new_[20515]_  = \new_[20516]_ ;
  assign \new_[20516]_  = ~\new_[10384]_ ;
  assign \new_[20517]_  = ~\new_[20549]_ ;
  assign \new_[20518]_  = ~\new_[20519]_ ;
  assign \new_[20519]_  = \new_[9569]_ ;
  assign \new_[20520]_  = ~\new_[20521]_ ;
  assign \new_[20521]_  = ~\new_[10513]_ ;
  assign wbs_rty_o = ~\new_[20523]_ ;
  assign \new_[20523]_  = ~\new_[9806]_ ;
  assign \new_[20524]_  = ~\new_[20525]_ ;
  assign \new_[20525]_  = \new_[20171]_ ;
  assign \new_[20526]_  = ~\new_[20527]_ ;
  assign \new_[20527]_  = ~\new_[13841]_ ;
  assign \new_[20528]_  = \new_[20198]_ ;
  assign \new_[20529]_  = ~\new_[20530]_ ;
  assign \new_[20530]_  = \new_[20040]_ ;
  assign \new_[20531]_  = ~\new_[20532]_ ;
  assign \new_[20532]_  = \new_[20533]_ ;
  assign \new_[20533]_  = ~\new_[20534]_ ;
  assign \new_[20534]_  = ~\new_[20535]_ ;
  assign \new_[20535]_  = ~\new_[13810]_ ;
  assign \new_[20536]_  = ~\new_[20555]_  & ~\new_[20537]_ ;
  assign \new_[20537]_  = ~\wbs_cti_i[0]  | ~\wbs_cti_i[2] ;
  assign \new_[20538]_  = ~\new_[20543]_  | ~\new_[5295]_  | ~\new_[20541]_ ;
  assign \new_[20539]_  = ~\new_[20540]_ ;
  assign \new_[20540]_  = \new_[17880]_  ? \new_[20545]_  : \new_[19272]_ ;
  assign \new_[20541]_  = \new_[20542]_ ;
  assign \new_[20542]_  = \new_[20229]_  ? \new_[20545]_  : \new_[20230]_ ;
  assign \new_[20543]_  = \new_[20544]_ ;
  assign \new_[20544]_  = \new_[19023]_  ? \new_[20545]_  : \new_[17826]_ ;
  assign \new_[20545]_  = ~\new_[20546]_  | ~\new_[20549]_ ;
  assign \new_[20546]_  = ~\new_[20547]_  | ~\new_[20548]_ ;
  assign \new_[20547]_  = ~\new_[19961]_  | ~\new_[19962]_ ;
  assign \new_[20548]_  = ~\new_[19890]_  & ~\new_[15026]_ ;
  assign \new_[20549]_  = \new_[20550]_ ;
  assign \new_[20550]_  = ~\new_[20106]_  | ~\new_[19925]_ ;
  assign \new_[20551]_  = \new_[19983]_ ;
  assign \new_[20552]_  = ~\new_[20553]_ ;
  assign \new_[20553]_  = ~\new_[19983]_ ;
  assign \new_[20554]_  = ~\new_[20555]_ ;
  assign \new_[20555]_  = ~\wbs_cti_i[1] ;
  assign n1340 = n1345;
  assign n1365 = n1370;
  assign n1375 = n1380;
  assign n1835 = n1855;
  assign n1845 = n1860;
  assign n2435 = n2440;
  assign n3335 = n5435;
  assign n3340 = n3450;
  assign n3345 = n3360;
  assign n3350 = n3375;
  assign n3355 = n5405;
  assign n3365 = n3425;
  assign n3370 = n3410;
  assign n3380 = n3425;
  assign n3385 = n3425;
  assign n3390 = n3450;
  assign n3395 = n5430;
  assign n3400 = n3435;
  assign n3405 = n5390;
  assign n3415 = n3450;
  assign n3420 = n5395;
  assign n3430 = n5430;
  assign n3440 = n5435;
  assign n3445 = n5410;
  assign n5380 = n5430;
  assign n5415 = n5435;
  assign n6865 = n6875;
  assign n6870 = n6875;
  assign n7470 = n7475;
  assign n10645 = n12765;
  assign n10650 = n12765;
  assign n12760 = n12765;
  assign n16335 = n16345;
  assign n16390 = n16500;
  assign n17170 = \wbm_dat_i[13] ;
  assign n17175 = \wbm_dat_i[11] ;
  assign n17180 = \wbm_dat_i[10] ;
  assign n17190 = \wbm_dat_i[15] ;
  assign n17205 = \wbm_dat_i[6] ;
  assign n17215 = \wbm_dat_i[25] ;
  assign n17225 = n17340;
  assign n17230 = \wbm_dat_i[19] ;
  assign n17235 = \wbm_dat_i[30] ;
  assign n17295 = \wbm_dat_i[4] ;
  assign n17305 = \wbm_dat_i[8] ;
  assign n17310 = \wbm_dat_i[16] ;
  assign n17315 = \wbm_dat_i[17] ;
  assign n17320 = \wbm_dat_i[1] ;
  assign n17330 = \wbm_dat_i[26] ;
  assign n17345 = \wbm_dat_i[22] ;
  assign n17370 = \wbm_dat_i[23] ;
  assign n17380 = \wbm_dat_i[12] ;
  assign n17390 = \wbm_dat_i[21] ;
  assign n17405 = \wbm_dat_i[20] ;
  assign n17415 = \wbm_dat_i[9] ;
  assign n17420 = \wbm_dat_i[24] ;
  assign n17425 = \wbm_dat_i[7] ;
  assign n17440 = \wbm_dat_i[14] ;
  assign n17445 = \wbm_dat_i[31] ;
  assign n17455 = \wbm_dat_i[0] ;
  assign n17465 = n17495;
  assign n17470 = \wbm_dat_i[3] ;
  assign n17475 = \wbm_dat_i[18] ;
  assign n17485 = \wbm_dat_i[27] ;
  assign n17490 = \wbm_dat_i[28] ;
  assign n17505 = \wbm_dat_i[5] ;
  assign n17510 = \wbm_dat_i[29] ;
  assign n17515 = \wbm_dat_i[2] ;
  assign n17325 = 1'b1;
  always @ (posedge clock) begin
    \\pci_target_unit_wishbone_master_wb_cti_o_reg[0]  <= n740;
    \\pci_target_unit_wishbone_master_wb_cti_o_reg[2]  <= n745;
    configuration_status_bit8_reg <= n750;
    \\pci_target_unit_wishbone_master_wb_sel_o_reg[0]  <= n755;
    \\pci_target_unit_wishbone_master_wb_sel_o_reg[1]  <= n760;
    \\pci_target_unit_wishbone_master_wb_sel_o_reg[2]  <= n765;
    \\pci_target_unit_wishbone_master_wb_sel_o_reg[3]  <= n770;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[0]  <= n775;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[10]  <= n780;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[11]  <= n785;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[12]  <= n790;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[13]  <= n795;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[16]  <= n800;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[17]  <= n805;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[19]  <= n810;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[1]  <= n815;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[20]  <= n820;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[21]  <= n825;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[22]  <= n830;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[23]  <= n835;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[24]  <= n840;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[25]  <= n845;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[26]  <= n850;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[27]  <= n855;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[28]  <= n860;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[29]  <= n865;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[2]  <= n870;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[31]  <= n875;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[3]  <= n880;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[4]  <= n885;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[5]  <= n890;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[6]  <= n895;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[8]  <= n900;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[9]  <= n905;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[30]  <= n910;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[14]  <= n915;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[18]  <= n920;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[7]  <= n925;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[15]  <= n930;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[19]  <= n935;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[22]  <= n940;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[24]  <= n945;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[20]  <= n950;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[27]  <= n955;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[21]  <= n960;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[30]  <= n965;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[25]  <= n970;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[28]  <= n975;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[31]  <= n980;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[29]  <= n985;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[17]  <= n990;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[10]  <= n995;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[11]  <= n1000;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[12]  <= n1005;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[16]  <= n1010;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[14]  <= n1015;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[13]  <= n1020;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[23]  <= n1025;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[26]  <= n1030;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[3]  <= n1035;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[4]  <= n1040;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[5]  <= n1045;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[6]  <= n1050;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[8]  <= n1055;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[9]  <= n1060;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[2]  <= n1065;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[18]  <= n1070;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[15]  <= n1075;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[7]  <= n1080;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[0]  <= n1085;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[1]  <= n1090;
    parity_checker_perr_sampled_reg <= n1095;
    \\pci_target_unit_wishbone_master_bc_register_reg[0]  <= n1100;
    \\pci_target_unit_wishbone_master_bc_register_reg[1]  <= n1105;
    \\pci_target_unit_wishbone_master_bc_register_reg[2]  <= n1110;
    \\pci_target_unit_wishbone_master_bc_register_reg[3]  <= n1115;
    pci_target_unit_wishbone_master_burst_chopped_reg <= n1120;
    pci_target_unit_pci_target_sm_backoff_reg <= n1125;
    wishbone_slave_unit_del_sync_req_done_reg_reg <= n1130;
    \\wishbone_slave_unit_wishbone_slave_c_state_reg[0]  <= n1135;
    \\pci_target_unit_wishbone_master_wb_cti_o_reg[1]  <= n1140;
    wishbone_slave_unit_del_sync_req_comp_pending_reg <= n1145;
    \\wishbone_slave_unit_wishbone_slave_c_state_reg[2]  <= n1150;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[36]  <= n1155;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[38]  <= n1160;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[39]  <= n1165;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[10]  <= n1170;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[11]  <= n1175;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[12]  <= n1180;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[0]  <= n1185;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[13]  <= n1190;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[16]  <= n1195;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[14]  <= n1200;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[17]  <= n1205;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[19]  <= n1210;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[1]  <= n1215;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[20]  <= n1220;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[21]  <= n1225;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[22]  <= n1230;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[23]  <= n1235;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[24]  <= n1240;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[25]  <= n1245;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[26]  <= n1250;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[27]  <= n1255;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[28]  <= n1260;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[29]  <= n1265;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[2]  <= n1270;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[30]  <= n1275;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[31]  <= n1280;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[32]  <= n1285;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[33]  <= n1290;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[34]  <= n1295;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[35]  <= n1300;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[37]  <= n1305;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[3]  <= n1310;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[4]  <= n1315;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[5]  <= n1320;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[6]  <= n1325;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[8]  <= n1330;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[9]  <= n1335;
    output_backup_trdy_out_reg <= n1340;
    pci_io_mux_trdy_iob_dat_out_reg <= n1345;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[15]  <= n1350;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[18]  <= n1355;
    \\pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg[7]  <= n1360;
    pci_io_mux_stop_iob_dat_out_reg <= n1365;
    output_backup_stop_out_reg <= n1370;
    pci_io_mux_devsel_iob_dat_out_reg <= n1375;
    output_backup_devsel_out_reg <= n1380;
    output_backup_perr_en_out_reg <= n1385;
    \\output_backup_ad_out_reg[31]  <= n1390;
    pci_io_mux_ad_iob31_dat_out_reg <= n1395;
    pci_io_mux_perr_iob_en_out_reg <= n1400;
    \\configuration_status_bit15_11_reg[15]  <= n1405;
    wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg <= n1410;
    \\output_backup_cbe_out_reg[0]  <= n1415;
    \\output_backup_cbe_out_reg[3]  <= n1420;
    pci_io_mux_cbe_iob0_dat_out_reg <= n1425;
    pci_io_mux_cbe_iob2_dat_out_reg <= n1430;
    \\output_backup_cbe_out_reg[2]  <= n1435;
    pci_io_mux_cbe_iob3_dat_out_reg <= n1440;
    \\output_backup_ad_out_reg[15]  <= n1445;
    \\output_backup_ad_out_reg[23]  <= n1450;
    \\output_backup_ad_out_reg[24]  <= n1455;
    \\output_backup_ad_out_reg[27]  <= n1460;
    \\output_backup_ad_out_reg[28]  <= n1465;
    \\output_backup_ad_out_reg[29]  <= n1470;
    \\output_backup_ad_out_reg[2]  <= n1475;
    \\output_backup_ad_out_reg[3]  <= n1480;
    \\output_backup_ad_out_reg[4]  <= n1485;
    \\output_backup_ad_out_reg[5]  <= n1490;
    \\output_backup_ad_out_reg[6]  <= n1495;
    \\output_backup_ad_out_reg[7]  <= n1500;
    \\output_backup_ad_out_reg[8]  <= n1505;
    pci_io_mux_ad_iob11_dat_out_reg <= n1510;
    pci_io_mux_ad_iob12_dat_out_reg <= n1515;
    pci_io_mux_ad_iob13_dat_out_reg <= n1520;
    pci_io_mux_ad_iob14_dat_out_reg <= n1525;
    pci_io_mux_ad_iob15_dat_out_reg <= n1530;
    pci_io_mux_ad_iob24_dat_out_reg <= n1535;
    pci_io_mux_ad_iob27_dat_out_reg <= n1540;
    pci_io_mux_ad_iob29_dat_out_reg <= n1545;
    pci_io_mux_ad_iob28_dat_out_reg <= n1550;
    pci_io_mux_ad_iob2_dat_out_reg <= n1555;
    pci_io_mux_ad_iob4_dat_out_reg <= n1560;
    pci_io_mux_ad_iob5_dat_out_reg <= n1565;
    pci_io_mux_ad_iob6_dat_out_reg <= n1570;
    pci_io_mux_ad_iob7_dat_out_reg <= n1575;
    pci_io_mux_ad_iob23_dat_out_reg <= n1580;
    pci_io_mux_ad_iob8_dat_out_reg <= n1585;
    pci_io_mux_ad_iob3_dat_out_reg <= n1590;
    \\output_backup_ad_out_reg[13]  <= n1595;
    \\output_backup_ad_out_reg[14]  <= n1600;
    \\output_backup_ad_out_reg[16]  <= n1605;
    \\output_backup_ad_out_reg[17]  <= n1610;
    \\output_backup_ad_out_reg[18]  <= n1615;
    \\output_backup_ad_out_reg[19]  <= n1620;
    \\output_backup_ad_out_reg[20]  <= n1625;
    \\output_backup_ad_out_reg[22]  <= n1630;
    \\output_backup_ad_out_reg[9]  <= n1635;
    pci_io_mux_ad_iob10_dat_out_reg <= n1640;
    pci_io_mux_ad_iob16_dat_out_reg <= n1645;
    pci_io_mux_ad_iob17_dat_out_reg <= n1650;
    pci_io_mux_ad_iob18_dat_out_reg <= n1655;
    pci_io_mux_ad_iob19_dat_out_reg <= n1660;
    pci_io_mux_ad_iob22_dat_out_reg <= n1665;
    pci_io_mux_ad_iob20_dat_out_reg <= n1670;
    \\output_backup_ad_out_reg[10]  <= n1675;
    pci_io_mux_ad_iob9_dat_out_reg <= n1680;
    \\output_backup_ad_out_reg[11]  <= n1685;
    \\output_backup_ad_out_reg[12]  <= n1690;
    \\output_backup_ad_out_reg[1]  <= n1695;
    \\output_backup_ad_out_reg[30]  <= n1700;
    pci_io_mux_ad_iob1_dat_out_reg <= n1705;
    pci_io_mux_ad_iob30_dat_out_reg <= n1710;
    \\output_backup_ad_out_reg[21]  <= n1715;
    pci_io_mux_ad_iob21_dat_out_reg <= n1720;
    \\configuration_status_bit15_11_reg[14]  <= n1725;
    \\output_backup_ad_out_reg[26]  <= n1730;
    pci_io_mux_ad_iob26_dat_out_reg <= n1735;
    pci_io_mux_ad_iob0_dat_out_reg <= n1740;
    \\output_backup_ad_out_reg[0]  <= n1745;
    parity_checker_perr_en_crit_gen_perr_en_reg_out_reg <= n1750;
    \\output_backup_ad_out_reg[25]  <= n1755;
    pci_io_mux_ad_iob25_dat_out_reg <= n1760;
    \\wishbone_slave_unit_pci_initiator_if_be_out_reg[0]  <= n1765;
    \\wishbone_slave_unit_pci_initiator_if_be_out_reg[2]  <= n1770;
    \\wishbone_slave_unit_pci_initiator_if_be_out_reg[3]  <= n1775;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[10]  <= n1780;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[11]  <= n1785;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[16]  <= n1790;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[18]  <= n1795;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[19]  <= n1800;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[1]  <= n1805;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[21]  <= n1810;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[22]  <= n1815;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[30]  <= n1820;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[5]  <= n1825;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[6]  <= n1830;
    pci_io_mux_perr_iob_dat_out_reg <= n1835;
    pci_io_mux_serr_iob_en_out_reg <= n1840;
    pci_io_mux_serr_iob_dat_out_reg <= n1845;
    pci_target_unit_wishbone_master_first_wb_data_access_reg <= n1850;
    output_backup_perr_out_reg <= n1855;
    output_backup_serr_out_reg <= n1860;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[15]  <= n1865;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[24]  <= n1870;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[25]  <= n1875;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[27]  <= n1880;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[2]  <= n1885;
    output_backup_serr_en_out_reg <= n1890;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[0]  <= n1895;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[12]  <= n1900;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[13]  <= n1905;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[14]  <= n1910;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[17]  <= n1915;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[20]  <= n1920;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[23]  <= n1925;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[26]  <= n1930;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[28]  <= n1935;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[29]  <= n1940;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[31]  <= n1945;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[3]  <= n1950;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[4]  <= n1955;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[7]  <= n1960;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[8]  <= n1965;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[9]  <= n1970;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]  <= n1975;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]  <= n1980;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]  <= n1985;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]  <= n1990;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]  <= n1995;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]  <= n2000;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]  <= n2005;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]  <= n2010;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]  <= n2015;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]  <= n2020;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]  <= n2025;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]  <= n2030;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29]  <= n2035;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2]  <= n2040;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4]  <= n2045;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]  <= n2050;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]  <= n2055;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[26]  <= n2060;
    \\pci_target_unit_fifos_pciw_outTransactionCount_reg[1]  <= n2065;
    \\pci_target_unit_fifos_outGreyCount_reg[0]  <= n2070;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]  <= n2075;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0]  <= n2080;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]  <= n2085;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]  <= n2090;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]  <= n2095;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]  <= n2100;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[0]  <= n2105;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[2]  <= n2110;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[0]  <= n2115;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[10]  <= n2120;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[11]  <= n2125;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[12]  <= n2130;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[13]  <= n2135;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[14]  <= n2140;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[15]  <= n2145;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[17]  <= n2150;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[18]  <= n2155;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[19]  <= n2160;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[20]  <= n2165;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[22]  <= n2170;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[24]  <= n2175;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[27]  <= n2180;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[28]  <= n2185;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[29]  <= n2190;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[2]  <= n2195;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[31]  <= n2200;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[3]  <= n2205;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[4]  <= n2210;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[6]  <= n2215;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[7]  <= n2220;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[8]  <= n2225;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]  <= n2230;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]  <= n2235;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]  <= n2240;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]  <= n2245;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]  <= n2250;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]  <= n2255;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]  <= n2260;
    \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]  <= n2265;
    \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]  <= n2270;
    \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]  <= n2275;
    \\wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[0]  <= n2280;
    \\pci_target_unit_fifos_pciw_outTransactionCount_reg[0]  <= n2285;
    \\pci_target_unit_fifos_outGreyCount_reg[1]  <= n2290;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1]  <= n2295;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2]  <= n2300;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[0]  <= n2305;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[1]  <= n2310;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[2]  <= n2315;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg[0]  <= n2320;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg[2]  <= n2325;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg[0]  <= n2330;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg[1]  <= n2335;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg[2]  <= n2340;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[0]  <= n2345;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[1]  <= n2350;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[2]  <= n2355;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg[1]  <= n2360;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9]  <= n2365;
    \\wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[1]  <= n2370;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[5]  <= n2375;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[9]  <= n2380;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[1]  <= n2385;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[23]  <= n2390;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[16]  <= n2395;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[3]  <= n2400;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[21]  <= n2405;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[25]  <= n2410;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0]  <= n2415;
    pci_target_unit_wishbone_master_wb_we_o_reg <= n2420;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]  <= n2425;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2]  <= n2430;
    pci_target_unit_wishbone_master_wb_cyc_o_reg <= n2435;
    pci_target_unit_wishbone_master_wb_stb_o_reg <= n2440;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[10]  <= n2445;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[11]  <= n2450;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[16]  <= n2455;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[18]  <= n2460;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[19]  <= n2465;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[1]  <= n2470;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[21]  <= n2475;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[22]  <= n2480;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[30]  <= n2485;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[5]  <= n2490;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[6]  <= n2495;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[30]  <= n2500;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[15]  <= n2505;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[24]  <= n2510;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[25]  <= n2515;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[27]  <= n2520;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[2]  <= n2525;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[36]  <= n2530;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[37]  <= n2535;
    \\pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_reg[1]  <= n2540;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[0]  <= n2545;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[12]  <= n2550;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[13]  <= n2555;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[14]  <= n2560;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[17]  <= n2565;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[20]  <= n2570;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[23]  <= n2575;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[26]  <= n2580;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[28]  <= n2585;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[29]  <= n2590;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[31]  <= n2595;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[3]  <= n2600;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[4]  <= n2605;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[7]  <= n2610;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[8]  <= n2615;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg[9]  <= n2620;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[15]  <= n2625;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[25]  <= n2630;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[7]  <= n2635;
    parity_checker_check_perr_reg <= n2640;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[0]  <= n2645;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[10]  <= n2650;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[11]  <= n2655;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[13]  <= n2660;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[14]  <= n2665;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[17]  <= n2670;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[18]  <= n2675;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[19]  <= n2680;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[21]  <= n2685;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[22]  <= n2690;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[20]  <= n2695;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[24]  <= n2700;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[26]  <= n2705;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[28]  <= n2710;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[29]  <= n2715;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[2]  <= n2720;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[31]  <= n2725;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[3]  <= n2730;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[4]  <= n2735;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[6]  <= n2740;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[8]  <= n2745;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[9]  <= n2750;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[5]  <= n2755;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[30]  <= n2760;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[27]  <= n2765;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[23]  <= n2770;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[12]  <= n2775;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[1]  <= n2780;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[16]  <= n2785;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[26]  <= n2790;
    output_backup_par_en_out_reg <= n2795;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[15]  <= n2800;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[16]  <= n2805;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[17]  <= n2810;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[18]  <= n2815;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[19]  <= n2820;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[1]  <= n2825;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[20]  <= n2830;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[22]  <= n2835;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[23]  <= n2840;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[24]  <= n2845;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[27]  <= n2850;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[28]  <= n2855;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[29]  <= n2860;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[2]  <= n2865;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[31]  <= n2870;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[3]  <= n2875;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[4]  <= n2880;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[5]  <= n2885;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[6]  <= n2890;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[7]  <= n2895;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[8]  <= n2900;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[9]  <= n2905;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[32]  <= n2910;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[34]  <= n2915;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[35]  <= n2920;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[0]  <= n2925;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[10]  <= n2930;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[11]  <= n2935;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[12]  <= n2940;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[13]  <= n2945;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[14]  <= n2950;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[33]  <= n2955;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[36]  <= n2960;
    pci_io_mux_par_iob_en_out_reg <= n2965;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[21]  <= n2970;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[25]  <= n2975;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg[30]  <= n2980;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[25]  <= n2985;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[15]  <= n2990;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[7]  <= n2995;
    \\pci_target_unit_wishbone_master_c_state_reg[0]  <= n3000;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[17]  <= n3005;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[18]  <= n3010;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[16]  <= n3015;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[19]  <= n3020;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[1]  <= n3025;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[20]  <= n3030;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[21]  <= n3035;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[23]  <= n3040;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[24]  <= n3045;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[22]  <= n3050;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[26]  <= n3055;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[27]  <= n3060;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[28]  <= n3065;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[29]  <= n3070;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[2]  <= n3075;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[30]  <= n3080;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[31]  <= n3085;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[3]  <= n3090;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[4]  <= n3095;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[5]  <= n3100;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[6]  <= n3105;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[8]  <= n3110;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[9]  <= n3115;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[37]  <= n3120;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[0]  <= n3125;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[10]  <= n3130;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[11]  <= n3135;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[12]  <= n3140;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[13]  <= n3145;
    \\pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg[14]  <= n3150;
    i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg <= n3155;
    pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg <= n3160;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]  <= n3165;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]  <= n3170;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]  <= n3175;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]  <= n3180;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]  <= n3185;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]  <= n3190;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]  <= n3195;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]  <= n3200;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]  <= n3205;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]  <= n3210;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]  <= n3215;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]  <= n3220;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]  <= n3225;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]  <= n3230;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]  <= n3235;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]  <= n3240;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]  <= n3245;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]  <= n3250;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]  <= n3255;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]  <= n3260;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]  <= n3265;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]  <= n3270;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]  <= n3275;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]  <= n3280;
    i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg <= n3285;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]  <= n3290;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]  <= n3295;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]  <= n3300;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]  <= n3305;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]  <= n3310;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]  <= n3315;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][11]  <= n3320;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][19]  <= n3325;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][19]  <= n3330;
    pci_io_mux_ad_iob23_en_out_reg <= n3335;
    pci_io_mux_ad_iob22_en_out_reg <= n3340;
    pci_io_mux_ad_iob21_en_out_reg <= n3345;
    pci_io_mux_ad_iob19_en_out_reg <= n3350;
    pci_io_mux_ad_iob17_en_out_reg <= n3355;
    pci_io_mux_ad_iob18_en_out_reg <= n3360;
    pci_io_mux_ad_iob15_en_out_reg <= n3365;
    pci_io_mux_ad_iob14_en_out_reg <= n3370;
    pci_io_mux_ad_iob13_en_out_reg <= n3375;
    pci_io_mux_ad_iob11_en_out_reg <= n3380;
    pci_io_mux_ad_iob25_en_out_reg <= n3385;
    pci_io_mux_ad_iob8_en_out_reg <= n3390;
    pci_io_mux_ad_iob7_en_out_reg <= n3395;
    pci_io_mux_ad_iob9_en_out_reg <= n3400;
    pci_io_mux_ad_iob5_en_out_reg <= n3405;
    pci_io_mux_ad_iob3_en_out_reg <= n3410;
    pci_io_mux_ad_iob4_en_out_reg <= n3415;
    pci_io_mux_ad_iob1_en_out_reg <= n3420;
    pci_io_mux_ad_iob2_en_out_reg <= n3425;
    pci_io_mux_ad_iob26_en_out_reg <= n3430;
    pci_io_mux_ad_iob31_en_out_reg <= n3435;
    pci_io_mux_ad_iob29_en_out_reg <= n3440;
    pci_io_mux_ad_iob28_en_out_reg <= n3445;
    pci_io_mux_ad_iob27_en_out_reg <= n3450;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][35]  <= n3455;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][35]  <= n3460;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][35]  <= n3465;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][35]  <= n3470;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][35]  <= n3475;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][35]  <= n3480;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][35]  <= n3485;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][35]  <= n3490;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][35]  <= n3495;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][0]  <= n3500;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][10]  <= n3505;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][11]  <= n3510;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][13]  <= n3515;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][15]  <= n3520;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][16]  <= n3525;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][17]  <= n3530;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][18]  <= n3535;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][19]  <= n3540;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][20]  <= n3545;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][21]  <= n3550;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][23]  <= n3555;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][24]  <= n3560;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][26]  <= n3565;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][28]  <= n3570;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][29]  <= n3575;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][30]  <= n3580;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][31]  <= n3585;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][3]  <= n3590;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][7]  <= n3595;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][8]  <= n3600;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][9]  <= n3605;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][10]  <= n3610;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][11]  <= n3615;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][13]  <= n3620;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][15]  <= n3625;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][16]  <= n3630;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][18]  <= n3635;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][19]  <= n3640;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][20]  <= n3645;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][23]  <= n3650;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][24]  <= n3655;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][26]  <= n3660;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][27]  <= n3665;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][1]  <= n3670;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][30]  <= n3675;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][31]  <= n3680;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][3]  <= n3685;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][7]  <= n3690;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][8]  <= n3695;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][9]  <= n3700;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][0]  <= n3705;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][11]  <= n3710;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][13]  <= n3715;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][15]  <= n3720;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][16]  <= n3725;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][17]  <= n3730;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][18]  <= n3735;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][19]  <= n3740;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][1]  <= n3745;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][20]  <= n3750;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][23]  <= n3755;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][24]  <= n3760;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][26]  <= n3765;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][27]  <= n3770;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][28]  <= n3775;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][30]  <= n3780;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][31]  <= n3785;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][3]  <= n3790;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][7]  <= n3795;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][8]  <= n3800;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][9]  <= n3805;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][0]  <= n3810;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][10]  <= n3815;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][13]  <= n3820;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][15]  <= n3825;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][16]  <= n3830;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][17]  <= n3835;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][18]  <= n3840;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][1]  <= n3845;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][20]  <= n3850;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][21]  <= n3855;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][23]  <= n3860;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][24]  <= n3865;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][26]  <= n3870;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][27]  <= n3875;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][28]  <= n3880;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][29]  <= n3885;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][30]  <= n3890;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][31]  <= n3895;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][3]  <= n3900;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][7]  <= n3905;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][8]  <= n3910;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][0]  <= n3915;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][10]  <= n3920;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][11]  <= n3925;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][13]  <= n3930;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][15]  <= n3935;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][17]  <= n3940;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][18]  <= n3945;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][19]  <= n3950;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][20]  <= n3955;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][21]  <= n3960;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][23]  <= n3965;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][24]  <= n3970;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][26]  <= n3975;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][27]  <= n3980;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][28]  <= n3985;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][29]  <= n3990;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][30]  <= n3995;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][31]  <= n4000;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][3]  <= n4005;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][7]  <= n4010;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][8]  <= n4015;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][9]  <= n4020;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][10]  <= n4025;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][11]  <= n4030;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][13]  <= n4035;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][15]  <= n4040;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][16]  <= n4045;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][17]  <= n4050;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][18]  <= n4055;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][19]  <= n4060;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][1]  <= n4065;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][21]  <= n4070;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][23]  <= n4075;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][24]  <= n4080;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][26]  <= n4085;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][27]  <= n4090;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][29]  <= n4095;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][30]  <= n4100;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][31]  <= n4105;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][3]  <= n4110;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][7]  <= n4115;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][8]  <= n4120;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][9]  <= n4125;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][0]  <= n4130;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][11]  <= n4135;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][13]  <= n4140;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][15]  <= n4145;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][16]  <= n4150;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][17]  <= n4155;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][19]  <= n4160;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][1]  <= n4165;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][20]  <= n4170;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][21]  <= n4175;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][23]  <= n4180;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][24]  <= n4185;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][26]  <= n4190;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][27]  <= n4195;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][28]  <= n4200;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][30]  <= n4205;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][31]  <= n4210;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][7]  <= n4215;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][8]  <= n4220;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][9]  <= n4225;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][0]  <= n4230;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][11]  <= n4235;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][13]  <= n4240;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][15]  <= n4245;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][16]  <= n4250;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][17]  <= n4255;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][19]  <= n4260;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][1]  <= n4265;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][20]  <= n4270;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][21]  <= n4275;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][23]  <= n4280;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][24]  <= n4285;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][26]  <= n4290;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][27]  <= n4295;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][28]  <= n4300;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][30]  <= n4305;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][31]  <= n4310;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][7]  <= n4315;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][8]  <= n4320;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][9]  <= n4325;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][0]  <= n4330;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][11]  <= n4335;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][13]  <= n4340;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][15]  <= n4345;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][16]  <= n4350;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][18]  <= n4355;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][1]  <= n4360;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][20]  <= n4365;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][21]  <= n4370;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][23]  <= n4375;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][24]  <= n4380;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][26]  <= n4385;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][27]  <= n4390;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][28]  <= n4395;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][29]  <= n4400;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][30]  <= n4405;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][31]  <= n4410;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][3]  <= n4415;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][7]  <= n4420;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][8]  <= n4425;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][17]  <= n4430;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][9]  <= n4435;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][0]  <= n4440;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][11]  <= n4445;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][13]  <= n4450;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][15]  <= n4455;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][16]  <= n4460;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][17]  <= n4465;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][19]  <= n4470;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][1]  <= n4475;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][20]  <= n4480;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][23]  <= n4485;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][24]  <= n4490;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][26]  <= n4495;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][27]  <= n4500;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][28]  <= n4505;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][30]  <= n4510;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][31]  <= n4515;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][7]  <= n4520;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][8]  <= n4525;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][9]  <= n4530;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][0]  <= n4535;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][11]  <= n4540;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][13]  <= n4545;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][15]  <= n4550;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][16]  <= n4555;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][17]  <= n4560;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][19]  <= n4565;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][1]  <= n4570;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][20]  <= n4575;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][21]  <= n4580;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][23]  <= n4585;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][24]  <= n4590;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][26]  <= n4595;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][27]  <= n4600;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][28]  <= n4605;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][30]  <= n4610;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][31]  <= n4615;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][7]  <= n4620;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][8]  <= n4625;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][9]  <= n4630;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][0]  <= n4635;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][10]  <= n4640;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][11]  <= n4645;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][13]  <= n4650;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][15]  <= n4655;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][16]  <= n4660;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][17]  <= n4665;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][18]  <= n4670;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][1]  <= n4675;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][20]  <= n4680;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][21]  <= n4685;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][23]  <= n4690;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][24]  <= n4695;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][26]  <= n4700;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][27]  <= n4705;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][28]  <= n4710;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][29]  <= n4715;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][30]  <= n4720;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][31]  <= n4725;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][35]  <= n4730;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][3]  <= n4735;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][7]  <= n4740;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][9]  <= n4745;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][8]  <= n4750;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][0]  <= n4755;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][10]  <= n4760;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][13]  <= n4765;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][15]  <= n4770;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][16]  <= n4775;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][17]  <= n4780;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][18]  <= n4785;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][1]  <= n4790;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][20]  <= n4795;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][21]  <= n4800;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][23]  <= n4805;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][24]  <= n4810;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][26]  <= n4815;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][27]  <= n4820;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][28]  <= n4825;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][29]  <= n4830;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][30]  <= n4835;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][31]  <= n4840;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][35]  <= n4845;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][3]  <= n4850;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][7]  <= n4855;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][8]  <= n4860;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][9]  <= n4865;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][0]  <= n4870;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][10]  <= n4875;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][11]  <= n4880;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][13]  <= n4885;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][15]  <= n4890;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][16]  <= n4895;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][17]  <= n4900;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][18]  <= n4905;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][1]  <= n4910;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][20]  <= n4915;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][21]  <= n4920;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][23]  <= n4925;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][24]  <= n4930;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][26]  <= n4935;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][27]  <= n4940;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][28]  <= n4945;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][29]  <= n4950;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][30]  <= n4955;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][31]  <= n4960;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][35]  <= n4965;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][3]  <= n4970;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][7]  <= n4975;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][8]  <= n4980;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][9]  <= n4985;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][0]  <= n4990;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][10]  <= n4995;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][13]  <= n5000;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][15]  <= n5005;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][16]  <= n5010;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][17]  <= n5015;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][18]  <= n5020;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][1]  <= n5025;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][20]  <= n5030;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][21]  <= n5035;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][23]  <= n5040;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][24]  <= n5045;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][26]  <= n5050;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][27]  <= n5055;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][28]  <= n5060;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][29]  <= n5065;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][30]  <= n5070;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][31]  <= n5075;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][35]  <= n5080;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][3]  <= n5085;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][7]  <= n5090;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][8]  <= n5095;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][9]  <= n5100;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][0]  <= n5105;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][10]  <= n5110;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][11]  <= n5115;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][13]  <= n5120;
    output_backup_mas_ad_en_out_reg <= n5125;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][15]  <= n5130;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][16]  <= n5135;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][17]  <= n5140;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][19]  <= n5145;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][1]  <= n5150;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][20]  <= n5155;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][23]  <= n5160;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][24]  <= n5165;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][26]  <= n5170;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][27]  <= n5175;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][28]  <= n5180;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][30]  <= n5185;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][31]  <= n5190;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][35]  <= n5195;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][3]  <= n5200;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][7]  <= n5205;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][8]  <= n5210;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][9]  <= n5215;
    output_backup_tar_ad_en_out_reg <= n5220;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][10]  <= n5225;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][19]  <= n5230;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][11]  <= n5235;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][29]  <= n5240;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][21]  <= n5245;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][19]  <= n5250;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][11]  <= n5255;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][28]  <= n5260;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][29]  <= n5265;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][21]  <= n5270;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][17]  <= n5275;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][19]  <= n5280;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][0]  <= n5285;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][29]  <= n5290;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][3]  <= n5295;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][28]  <= n5300;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][27]  <= n5305;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][10]  <= n5310;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][18]  <= n5315;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][1]  <= n5320;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][3]  <= n5325;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][21]  <= n5330;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][29]  <= n5335;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][35]  <= n5340;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][18]  <= n5345;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][10]  <= n5350;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][35]  <= n5355;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][10]  <= n5360;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][19]  <= n5365;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][29]  <= n5370;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][3]  <= n5375;
    pci_io_mux_ad_iob30_en_out_reg <= n5380;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][29]  <= n5385;
    pci_io_mux_ad_iob0_en_out_reg <= n5390;
    pci_io_mux_ad_iob6_en_out_reg <= n5395;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][18]  <= n5400;
    pci_io_mux_ad_iob12_en_out_reg <= n5405;
    pci_io_mux_ad_iob10_en_out_reg <= n5410;
    pci_io_mux_ad_iob16_en_out_reg <= n5415;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][10]  <= n5420;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][3]  <= n5425;
    pci_io_mux_ad_iob20_en_out_reg <= n5430;
    pci_io_mux_ad_iob24_en_out_reg <= n5435;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][18]  <= n5440;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][10]  <= n5445;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][20]  <= n5450;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][0]  <= n5455;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][1]  <= n5460;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][16]  <= n5465;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][9]  <= n5470;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][29]  <= n5475;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][21]  <= n5480;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][18]  <= n5485;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][33]  <= n5490;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][32]  <= n5495;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][33]  <= n5500;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][33]  <= n5505;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][32]  <= n5510;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][32]  <= n5515;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][33]  <= n5520;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][32]  <= n5525;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][32]  <= n5530;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][33]  <= n5535;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][33]  <= n5540;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][32]  <= n5545;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][32]  <= n5550;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][32]  <= n5555;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][32]  <= n5560;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][32]  <= n5565;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][32]  <= n5570;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][32]  <= n5575;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][33]  <= n5580;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][32]  <= n5585;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][33]  <= n5590;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][32]  <= n5595;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][33]  <= n5600;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][32]  <= n5605;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][32]  <= n5610;
    pci_target_unit_wishbone_master_first_data_is_burst_reg_reg <= n5615;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][33]  <= n5620;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][33]  <= n5625;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][33]  <= n5630;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][33]  <= n5635;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][33]  <= n5640;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][33]  <= n5645;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][33]  <= n5650;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][34]  <= n5655;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][5]  <= n5660;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][4]  <= n5665;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][2]  <= n5670;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][25]  <= n5675;
    i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg <= n5680;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][14]  <= n5685;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][22]  <= n5690;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][25]  <= n5695;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][4]  <= n5700;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][5]  <= n5705;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][14]  <= n5710;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][22]  <= n5715;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][2]  <= n5720;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][5]  <= n5725;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][4]  <= n5730;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][12]  <= n5735;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][22]  <= n5740;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][2]  <= n5745;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][34]  <= n5750;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][5]  <= n5755;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][12]  <= n5760;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][34]  <= n5765;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][4]  <= n5770;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][6]  <= n5775;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][12]  <= n5780;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][14]  <= n5785;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][4]  <= n5790;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][5]  <= n5795;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][22]  <= n5800;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][25]  <= n5805;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][4]  <= n5810;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][5]  <= n5815;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][12]  <= n5820;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][14]  <= n5825;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][22]  <= n5830;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][2]  <= n5835;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][4]  <= n5840;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][6]  <= n5845;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][5]  <= n5850;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][12]  <= n5855;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][22]  <= n5860;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][2]  <= n5865;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][4]  <= n5870;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][5]  <= n5875;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][12]  <= n5880;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][5]  <= n5885;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][12]  <= n5890;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][22]  <= n5895;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][2]  <= n5900;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][4]  <= n5905;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][5]  <= n5910;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][12]  <= n5915;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][22]  <= n5920;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][2]  <= n5925;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][4]  <= n5930;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][5]  <= n5935;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][12]  <= n5940;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][5]  <= n5945;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][12]  <= n5950;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][34]  <= n5955;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][6]  <= n5960;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][12]  <= n5965;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][5]  <= n5970;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][6]  <= n5975;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][12]  <= n5980;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][22]  <= n5985;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][34]  <= n5990;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][6]  <= n5995;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][34]  <= n6000;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][12]  <= n6005;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][22]  <= n6010;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][34]  <= n6015;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][4]  <= n6020;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][5]  <= n6025;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][34]  <= n6030;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][34]  <= n6035;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][4]  <= n6040;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][14]  <= n6045;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][6]  <= n6050;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][2]  <= n6055;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][25]  <= n6060;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][4]  <= n6065;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][22]  <= n6070;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][4]  <= n6075;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][14]  <= n6080;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][25]  <= n6085;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][5]  <= n6090;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][22]  <= n6095;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][2]  <= n6100;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][14]  <= n6105;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][25]  <= n6110;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][25]  <= n6115;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][6]  <= n6120;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][6]  <= n6125;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][2]  <= n6130;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][14]  <= n6135;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][34]  <= n6140;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][25]  <= n6145;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][34]  <= n6150;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][4]  <= n6155;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][25]  <= n6160;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][2]  <= n6165;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][34]  <= n6170;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][22]  <= n6175;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][12]  <= n6180;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][14]  <= n6185;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][6]  <= n6190;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][6]  <= n6195;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][34]  <= n6200;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][14]  <= n6205;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][6]  <= n6210;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][14]  <= n6215;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][12]  <= n6220;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][25]  <= n6225;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][14]  <= n6230;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][4]  <= n6235;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][6]  <= n6240;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][2]  <= n6245;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][25]  <= n6250;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][22]  <= n6255;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][14]  <= n6260;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][6]  <= n6265;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][25]  <= n6270;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][14]  <= n6275;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][25]  <= n6280;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][6]  <= n6285;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][34]  <= n6290;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][2]  <= n6295;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][22]  <= n6300;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][25]  <= n6305;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][14]  <= n6310;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][12]  <= n6315;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][34]  <= n6320;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][6]  <= n6325;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][2]  <= n6330;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][22]  <= n6335;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][2]  <= n6340;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][6]  <= n6345;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][5]  <= n6350;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][34]  <= n6355;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][25]  <= n6360;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][14]  <= n6365;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][25]  <= n6370;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][2]  <= n6375;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0]  <= n6380;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]  <= n6385;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]  <= n6390;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]  <= n6395;
    \\wishbone_slave_unit_del_sync_addr_out_reg[0]  <= n6400;
    \\wishbone_slave_unit_del_sync_addr_out_reg[10]  <= n6405;
    \\wishbone_slave_unit_del_sync_addr_out_reg[11]  <= n6410;
    \\wishbone_slave_unit_del_sync_addr_out_reg[13]  <= n6415;
    \\wishbone_slave_unit_del_sync_addr_out_reg[15]  <= n6420;
    \\wishbone_slave_unit_del_sync_addr_out_reg[16]  <= n6425;
    \\wishbone_slave_unit_del_sync_addr_out_reg[17]  <= n6430;
    \\wishbone_slave_unit_del_sync_addr_out_reg[19]  <= n6435;
    \\wishbone_slave_unit_del_sync_addr_out_reg[1]  <= n6440;
    \\wishbone_slave_unit_del_sync_addr_out_reg[20]  <= n6445;
    \\wishbone_slave_unit_del_sync_addr_out_reg[23]  <= n6450;
    \\wishbone_slave_unit_del_sync_addr_out_reg[24]  <= n6455;
    \\wishbone_slave_unit_del_sync_addr_out_reg[26]  <= n6460;
    \\wishbone_slave_unit_del_sync_addr_out_reg[27]  <= n6465;
    \\wishbone_slave_unit_del_sync_addr_out_reg[28]  <= n6470;
    \\wishbone_slave_unit_del_sync_addr_out_reg[30]  <= n6475;
    \\wishbone_slave_unit_del_sync_addr_out_reg[31]  <= n6480;
    \\wishbone_slave_unit_del_sync_addr_out_reg[7]  <= n6485;
    \\wishbone_slave_unit_del_sync_addr_out_reg[8]  <= n6490;
    \\wishbone_slave_unit_del_sync_addr_out_reg[9]  <= n6495;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]  <= n6500;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[0]  <= n6505;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]  <= n6510;
    \\wishbone_slave_unit_del_sync_addr_out_reg[3]  <= n6515;
    \\wishbone_slave_unit_del_sync_addr_out_reg[29]  <= n6520;
    \\wishbone_slave_unit_del_sync_addr_out_reg[18]  <= n6525;
    \\wishbone_slave_unit_del_sync_addr_out_reg[21]  <= n6530;
    \\pci_target_unit_pci_target_sm_c_state_reg[0]  <= n6535;
    \\pci_target_unit_pci_target_sm_c_state_reg[1]  <= n6540;
    \\pci_target_unit_pci_target_sm_c_state_reg[2]  <= n6545;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]  <= n6550;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0]  <= n6555;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1]  <= n6560;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3]  <= n6565;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[1]  <= n6570;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]  <= n6575;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[0]  <= n6580;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[1]  <= n6585;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[2]  <= n6590;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[3]  <= n6595;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[2]  <= n6600;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[9][36]  <= n6605;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[7][36]  <= n6610;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[3]  <= n6615;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]  <= n6620;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]  <= n6625;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2]  <= n6630;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3]  <= n6635;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[0]  <= n6640;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]  <= n6645;
    \\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[1]  <= n6650;
    \\wishbone_slave_unit_del_sync_addr_out_reg[12]  <= n6655;
    \\wishbone_slave_unit_del_sync_addr_out_reg[22]  <= n6660;
    \\wishbone_slave_unit_del_sync_addr_out_reg[2]  <= n6665;
    \\wishbone_slave_unit_del_sync_addr_out_reg[5]  <= n6670;
    \\wishbone_slave_unit_del_sync_addr_out_reg[4]  <= n6675;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[0][36]  <= n6680;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[8][36]  <= n6685;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[11][36]  <= n6690;
    \\wishbone_slave_unit_del_sync_addr_out_reg[25]  <= n6695;
    \\wishbone_slave_unit_del_sync_addr_out_reg[6]  <= n6700;
    \\wishbone_slave_unit_del_sync_addr_out_reg[14]  <= n6705;
    \\wishbone_slave_unit_fifos_inGreyCount_reg[0]  <= n6710;
    \\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2]  <= n6715;
    \\wishbone_slave_unit_fifos_inGreyCount_reg[1]  <= n6720;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[10][36]  <= n6725;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[1][36]  <= n6730;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[2][36]  <= n6735;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[3][36]  <= n6740;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[6][36]  <= n6745;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[13][36]  <= n6750;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[14][36]  <= n6755;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[12][36]  <= n6760;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[15][36]  <= n6765;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[5][36]  <= n6770;
    \\wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg[4][36]  <= n6775;
    \\wishbone_slave_unit_fifos_inGreyCount_reg[2]  <= n6780;
    \\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0]  <= n6785;
    i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg <= n6790;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2]  <= n6795;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]  <= n6800;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]  <= n6805;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0]  <= n6810;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1]  <= n6815;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[0]  <= n6820;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[1]  <= n6825;
    wishbone_slave_unit_del_sync_burst_out_reg <= n6830;
    pci_target_unit_wishbone_master_addr_into_cnt_reg_reg <= n6835;
    output_backup_trdy_en_out_reg <= n6840;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0]  <= n6845;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2]  <= n6850;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[2]  <= n6855;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1]  <= n6860;
    pci_io_mux_trdy_iob_en_out_reg <= n6865;
    pci_io_mux_stop_iob_en_out_reg <= n6870;
    pci_io_mux_devsel_iob_en_out_reg <= n6875;
    \\pci_target_unit_wishbone_master_rty_counter_reg[0]  <= n6880;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]  <= n6885;
    \\wishbone_slave_unit_del_sync_bc_out_reg[3]  <= n6890;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0]  <= n6895;
    output_backup_frame_out_reg <= n6900;
    \\pci_target_unit_wishbone_master_rty_counter_reg[5]  <= n6905;
    \\pci_target_unit_wishbone_master_rty_counter_reg[6]  <= n6910;
    \\wishbone_slave_unit_del_sync_bc_out_reg[2]  <= n6915;
    \\pci_target_unit_wishbone_master_rty_counter_reg[1]  <= n6920;
    \\pci_target_unit_wishbone_master_rty_counter_reg[2]  <= n6925;
    \\pci_target_unit_wishbone_master_rty_counter_reg[4]  <= n6930;
    \\wishbone_slave_unit_fifos_outGreyCount_reg[0]  <= n6935;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2]  <= n6940;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3]  <= n6945;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]  <= n6950;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]  <= n6955;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[0]  <= n6960;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[1]  <= n6965;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[2]  <= n6970;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[0]  <= n6975;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[1]  <= n6980;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[2]  <= n6985;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[0]  <= n6990;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[2]  <= n6995;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[3]  <= n7000;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[3]  <= n7005;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[1]  <= n7010;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[3]  <= n7015;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3]  <= n7020;
    \\pci_target_unit_wishbone_master_rty_counter_reg[3]  <= n7025;
    \\pci_target_unit_wishbone_master_rty_counter_reg[7]  <= n7030;
    pci_io_mux_frame_iob_dat_out_reg <= n7035;
    pci_target_unit_pci_target_sm_rd_request_reg <= n7040;
    pci_target_unit_pci_target_sm_rd_progress_reg <= n7045;
    \\wishbone_slave_unit_del_sync_be_out_reg[0]  <= n7050;
    \\wishbone_slave_unit_del_sync_be_out_reg[1]  <= n7055;
    \\wishbone_slave_unit_del_sync_be_out_reg[2]  <= n7060;
    wishbone_slave_unit_del_sync_we_out_reg <= n7065;
    \\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[1]  <= n7070;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]  <= n7075;
    \\wishbone_slave_unit_del_sync_be_out_reg[3]  <= n7080;
    \\wishbone_slave_unit_del_sync_bc_out_reg[1]  <= n7085;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[12]  <= n7090;
    pci_target_unit_pci_target_if_norm_prf_en_reg <= n7095;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[0]  <= n7100;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[10]  <= n7105;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[11]  <= n7110;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[13]  <= n7115;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[14]  <= n7120;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[15]  <= n7125;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[17]  <= n7130;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[18]  <= n7135;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[1]  <= n7140;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[21]  <= n7145;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[23]  <= n7150;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[25]  <= n7155;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[26]  <= n7160;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[27]  <= n7165;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[29]  <= n7170;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[2]  <= n7175;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[30]  <= n7180;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[32]  <= n7185;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[33]  <= n7190;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[34]  <= n7195;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[3]  <= n7200;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[5]  <= n7205;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[8]  <= n7210;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[7]  <= n7215;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]  <= n7220;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[10]  <= n7225;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[11]  <= n7230;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[14]  <= n7235;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[1]  <= n7240;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[3]  <= n7245;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[5]  <= n7250;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[9]  <= n7255;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[7]  <= n7260;
    \\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0]  <= n7265;
    pci_target_unit_pci_target_if_pciw_fifo_wenable_out_reg <= n7270;
    \\wishbone_slave_unit_fifos_outGreyCount_reg[2]  <= n7275;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[6]  <= n7280;
    \\wishbone_slave_unit_fifos_outGreyCount_reg[1]  <= n7285;
    \\wishbone_slave_unit_del_sync_bc_out_reg[0]  <= n7290;
    \\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2]  <= n7295;
    i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg <= n7300;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[6]  <= n7305;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[4]  <= n7310;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[13]  <= n7315;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[2]  <= n7320;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[15]  <= n7325;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[16]  <= n7330;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[9]  <= n7335;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[4]  <= n7340;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[35]  <= n7345;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[31]  <= n7350;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[22]  <= n7355;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[28]  <= n7360;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[24]  <= n7365;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[16]  <= n7370;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[20]  <= n7375;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[12]  <= n7380;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[19]  <= n7385;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[8]  <= n7390;
    pci_target_unit_pci_target_sm_wr_progress_reg <= n7395;
    pci_target_unit_wishbone_master_w_attempt_reg <= n7400;
    \\configuration_wb_am2_reg[31]  <= n7405;
    \\configuration_wb_am1_reg[31]  <= n7410;
    pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg <= n7415;
    \\output_backup_cbe_out_reg[1]  <= n7420;
    wishbone_slave_unit_pci_initiator_if_del_read_req_reg <= n7425;
    \\configuration_pci_img_ctrl1_bit2_1_reg[1]  <= n7430;
    \\configuration_pci_img_ctrl1_bit2_1_reg[2]  <= n7435;
    \\configuration_wb_ta1_reg[31]  <= n7440;
    configuration_wb_err_cs_bit0_reg <= n7445;
    \\configuration_wb_ta2_reg[31]  <= n7450;
    pci_io_mux_cbe_iob1_dat_out_reg <= n7455;
    pci_target_unit_pci_target_sm_master_will_request_read_reg <= n7460;
    wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg <= n7465;
    output_backup_par_out_reg <= n7470;
    pci_io_mux_par_iob_dat_out_reg <= n7475;
    configuration_pci_err_cs_bit0_reg <= n7480;
    \\configuration_wb_img_ctrl1_bit2_0_reg[2]  <= n7485;
    \\configuration_interrupt_line_reg[6]  <= n7490;
    \\configuration_wb_img_ctrl2_bit2_0_reg[1]  <= n7495;
    \\configuration_interrupt_line_reg[2]  <= n7500;
    wishbone_slave_unit_del_sync_req_req_pending_reg <= n7505;
    \\configuration_wb_img_ctrl1_bit2_0_reg[0]  <= n7510;
    \\configuration_wb_img_ctrl1_bit2_0_reg[1]  <= n7515;
    \\configuration_interrupt_line_reg[0]  <= n7520;
    \\configuration_interrupt_line_reg[1]  <= n7525;
    \\configuration_wb_img_ctrl2_bit2_0_reg[0]  <= n7530;
    \\configuration_wb_img_ctrl2_bit2_0_reg[2]  <= n7535;
    \\configuration_command_bit2_0_reg[0]  <= n7540;
    \\configuration_command_bit2_0_reg[1]  <= n7545;
    \\configuration_command_bit2_0_reg[2]  <= n7550;
    configuration_wb_ba1_bit0_reg <= n7555;
    configuration_wb_ba2_bit0_reg <= n7560;
    configuration_command_bit8_reg <= n7565;
    configuration_wb_err_cs_bit8_reg <= n7570;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]  <= n7575;
    \\configuration_status_bit15_11_reg[11]  <= n7580;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]  <= n7585;
    \\configuration_status_bit15_11_reg[12]  <= n7590;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]  <= n7595;
    \\configuration_status_bit15_11_reg[13]  <= n7600;
    \\configuration_isr_bit2_0_reg[1]  <= n7605;
    wishbone_slave_unit_del_sync_comp_comp_pending_reg <= n7610;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[0]  <= n7615;
    pci_target_unit_wishbone_master_reset_rty_cnt_reg <= n7620;
    \\configuration_wb_ba2_bit31_12_reg[31]  <= n7625;
    \\configuration_wb_ba1_bit31_12_reg[31]  <= n7630;
    configuration_command_bit6_reg <= n7635;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][1]  <= n7640;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][6]  <= n7645;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][3]  <= n7650;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[1]  <= n7655;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][26]  <= n7660;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][31]  <= n7665;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][2]  <= n7670;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][22]  <= n7675;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][24]  <= n7680;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][19]  <= n7685;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][20]  <= n7690;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][11]  <= n7695;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][0]  <= n7700;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][8]  <= n7705;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][15]  <= n7710;
    \\configuration_icr_bit2_0_reg[0]  <= n7715;
    \\configuration_icr_bit2_0_reg[1]  <= n7720;
    \\configuration_icr_bit2_0_reg[2]  <= n7725;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][4]  <= n7730;
    \\configuration_interrupt_line_reg[3]  <= n7735;
    \\configuration_cache_line_size_reg_reg[3]  <= n7740;
    \\configuration_interrupt_line_reg[5]  <= n7745;
    \\configuration_interrupt_line_reg[4]  <= n7750;
    \\configuration_cache_line_size_reg_reg[5]  <= n7755;
    \\configuration_cache_line_size_reg_reg[4]  <= n7760;
    configuration_sync_isr_2_del_bit_reg <= n7765;
    configuration_sync_pci_err_cs_8_del_bit_reg <= n7770;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]  <= n7775;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[0]  <= n7780;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[2]  <= n7785;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2]  <= n7790;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][0]  <= n7795;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][10]  <= n7800;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][12]  <= n7805;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][14]  <= n7810;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][16]  <= n7815;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][18]  <= n7820;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][1]  <= n7825;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][20]  <= n7830;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][21]  <= n7835;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][23]  <= n7840;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][25]  <= n7845;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][27]  <= n7850;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][29]  <= n7855;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][30]  <= n7860;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][37]  <= n7865;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][4]  <= n7870;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][5]  <= n7875;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][6]  <= n7880;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][8]  <= n7885;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][0]  <= n7890;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][11]  <= n7895;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][12]  <= n7900;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][13]  <= n7905;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][15]  <= n7910;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][16]  <= n7915;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][17]  <= n7920;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][19]  <= n7925;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][1]  <= n7930;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][20]  <= n7935;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][22]  <= n7940;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][24]  <= n7945;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][26]  <= n7950;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][28]  <= n7955;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][2]  <= n7960;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][31]  <= n7965;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][3]  <= n7970;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][4]  <= n7975;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][5]  <= n7980;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][7]  <= n7985;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][8]  <= n7990;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][9]  <= n7995;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][10]  <= n8000;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][11]  <= n8005;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][12]  <= n8010;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][14]  <= n8015;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][16]  <= n8020;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][18]  <= n8025;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][19]  <= n8030;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][1]  <= n8035;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][21]  <= n8040;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][23]  <= n8045;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][25]  <= n8050;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][26]  <= n8055;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][27]  <= n8060;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][29]  <= n8065;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][30]  <= n8070;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][37]  <= n8075;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][3]  <= n8080;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][4]  <= n8085;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][6]  <= n8090;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][7]  <= n8095;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][8]  <= n8100;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][0]  <= n8105;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][10]  <= n8110;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][11]  <= n8115;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][13]  <= n8120;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][15]  <= n8125;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][17]  <= n8130;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][18]  <= n8135;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][19]  <= n8140;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][20]  <= n8145;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][22]  <= n8150;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][24]  <= n8155;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][25]  <= n8160;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][26]  <= n8165;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][28]  <= n8170;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][29]  <= n8175;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][2]  <= n8180;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][31]  <= n8185;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][37]  <= n8190;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][3]  <= n8195;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][5]  <= n8200;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][7]  <= n8205;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][9]  <= n8210;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][14]  <= n8215;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][15]  <= n8220;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][16]  <= n8225;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][18]  <= n8230;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][1]  <= n8235;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][21]  <= n8240;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][22]  <= n8245;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][23]  <= n8250;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][25]  <= n8255;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][27]  <= n8260;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][29]  <= n8265;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][2]  <= n8270;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][30]  <= n8275;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][37]  <= n8280;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][4]  <= n8285;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][6]  <= n8290;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][7]  <= n8295;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][8]  <= n8300;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][0]  <= n8305;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][11]  <= n8310;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][13]  <= n8315;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][14]  <= n8320;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][15]  <= n8325;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][17]  <= n8330;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][18]  <= n8335;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][19]  <= n8340;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][20]  <= n8345;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][22]  <= n8350;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][24]  <= n8355;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][26]  <= n8360;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][28]  <= n8365;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][29]  <= n8370;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][2]  <= n8375;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][31]  <= n8380;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][3]  <= n8385;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][5]  <= n8390;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][7]  <= n8395;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][9]  <= n8400;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][10]  <= n8405;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][12]  <= n8410;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][13]  <= n8415;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][14]  <= n8420;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][16]  <= n8425;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][17]  <= n8430;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][18]  <= n8435;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][1]  <= n8440;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][21]  <= n8445;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][23]  <= n8450;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][25]  <= n8455;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][27]  <= n8460;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][28]  <= n8465;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][29]  <= n8470;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][30]  <= n8475;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][37]  <= n8480;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][4]  <= n8485;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][5]  <= n8490;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][6]  <= n8495;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][8]  <= n8500;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][9]  <= n8505;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][0]  <= n8510;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][11]  <= n8515;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][13]  <= n8520;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][15]  <= n8525;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][17]  <= n8530;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][19]  <= n8535;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][1]  <= n8540;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][20]  <= n8545;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][22]  <= n8550;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][24]  <= n8555;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][26]  <= n8560;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][27]  <= n8565;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][28]  <= n8570;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][2]  <= n8575;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][31]  <= n8580;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][3]  <= n8585;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][4]  <= n8590;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][5]  <= n8595;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][7]  <= n8600;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][9]  <= n8605;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][10]  <= n8610;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][12]  <= n8615;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][30]  <= n8620;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][37]  <= n8625;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][25]  <= n8630;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][27]  <= n8635;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][23]  <= n8640;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][21]  <= n8645;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][1]  <= n8650;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][16]  <= n8655;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][9]  <= n8660;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][10]  <= n8665;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[2][12]  <= n8670;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][26]  <= n8675;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][21]  <= n8680;
    \\configuration_cache_line_size_reg_reg[7]  <= n8685;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][3]  <= n8690;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][5]  <= n8695;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][31]  <= n8700;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][28]  <= n8705;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][24]  <= n8710;
    \\configuration_interrupt_line_reg[7]  <= n8715;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][19]  <= n8720;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][20]  <= n8725;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][17]  <= n8730;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][4]  <= n8735;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][8]  <= n8740;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][6]  <= n8745;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][30]  <= n8750;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][27]  <= n8755;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][23]  <= n8760;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][8]  <= n8765;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][9]  <= n8770;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][28]  <= n8775;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][14]  <= n8780;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][16]  <= n8785;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[7][12]  <= n8790;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][5]  <= n8795;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][2]  <= n8800;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][31]  <= n8805;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][24]  <= n8810;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][22]  <= n8815;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][0]  <= n8820;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][0]  <= n8825;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][20]  <= n8830;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][11]  <= n8835;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][13]  <= n8840;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][17]  <= n8845;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[1][13]  <= n8850;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[6][15]  <= n8855;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][29]  <= n8860;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][6]  <= n8865;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][6]  <= n8870;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][37]  <= n8875;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][21]  <= n8880;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][30]  <= n8885;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][29]  <= n8890;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][30]  <= n8895;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][37]  <= n8900;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][25]  <= n8905;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][23]  <= n8910;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][25]  <= n8915;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][10]  <= n8920;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][18]  <= n8925;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][27]  <= n8930;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][16]  <= n8935;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][18]  <= n8940;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][23]  <= n8945;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][12]  <= n8950;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[0][14]  <= n8955;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][21]  <= n8960;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][14]  <= n8965;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[5][10]  <= n8970;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][9]  <= n8975;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[3][7]  <= n8980;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][7]  <= n8985;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][28]  <= n8990;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][2]  <= n8995;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][3]  <= n9000;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][31]  <= n9005;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][26]  <= n9010;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][22]  <= n9015;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][24]  <= n9020;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][13]  <= n9025;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][19]  <= n9030;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][17]  <= n9035;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][15]  <= n9040;
    \\pci_target_unit_fifos_pcir_fifo_storage_mem_reg[4][11]  <= n9045;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[5]  <= n9050;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[7]  <= n9055;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[8]  <= n9060;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[23]  <= n9065;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[4]  <= n9070;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[31]  <= n9075;
    \\configuration_pci_ba0_bit31_8_reg[12]  <= n9080;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[27]  <= n9085;
    \\configuration_latency_timer_reg[1]  <= n9090;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[12]  <= n9095;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[1]  <= n9100;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[21]  <= n9105;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[14]  <= n9110;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[16]  <= n9115;
    \\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]  <= n9120;
    configuration_icr_bit31_reg <= n9125;
    wishbone_slave_unit_wishbone_slave_img_wallow_reg <= n9130;
    wishbone_slave_unit_wishbone_slave_do_del_request_reg <= n9135;
    wishbone_slave_unit_wishbone_slave_mrl_en_reg <= n9140;
    wishbone_slave_unit_wishbone_slave_pref_en_reg <= n9145;
    wishbone_slave_unit_wishbone_slave_del_addr_hit_reg <= n9150;
    \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]  <= n9155;
    wishbone_slave_unit_wishbone_slave_del_completion_allow_reg <= n9160;
    pci_target_unit_del_sync_comp_comp_pending_reg <= n9165;
    pci_target_unit_del_sync_comp_req_pending_reg <= n9170;
    \\pci_target_unit_wishbone_master_c_state_reg[2]  <= n9175;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][37]  <= n9180;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][37]  <= n9185;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][37]  <= n9190;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][37]  <= n9195;
    wishbone_slave_unit_pci_initiator_if_intermediate_last_reg <= n9200;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[1]  <= n9205;
    \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]  <= n9210;
    \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]  <= n9215;
    \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]  <= n9220;
    \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]  <= n9225;
    \\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]  <= n9230;
    \\configuration_latency_timer_reg[0]  <= n9235;
    \\configuration_latency_timer_reg[2]  <= n9240;
    \\configuration_latency_timer_reg[3]  <= n9245;
    \\configuration_latency_timer_reg[4]  <= n9250;
    \\configuration_latency_timer_reg[5]  <= n9255;
    \\configuration_latency_timer_reg[6]  <= n9260;
    \\configuration_latency_timer_reg[7]  <= n9265;
    \\configuration_cache_line_size_reg_reg[0]  <= n9270;
    \\configuration_pci_ba0_bit31_8_reg[14]  <= n9275;
    \\configuration_cache_line_size_reg_reg[1]  <= n9280;
    \\configuration_cache_line_size_reg_reg[2]  <= n9285;
    \\configuration_pci_ba0_bit31_8_reg[13]  <= n9290;
    \\configuration_pci_ba0_bit31_8_reg[17]  <= n9295;
    \\configuration_cache_line_size_reg_reg[6]  <= n9300;
    \\configuration_pci_ba0_bit31_8_reg[16]  <= n9305;
    \\configuration_pci_ba0_bit31_8_reg[20]  <= n9310;
    \\configuration_pci_ba0_bit31_8_reg[23]  <= n9315;
    \\configuration_pci_ba0_bit31_8_reg[18]  <= n9320;
    \\configuration_pci_ba0_bit31_8_reg[15]  <= n9325;
    \\configuration_pci_ba0_bit31_8_reg[19]  <= n9330;
    \\configuration_pci_ba0_bit31_8_reg[25]  <= n9335;
    \\configuration_pci_ba0_bit31_8_reg[27]  <= n9340;
    \\configuration_pci_ba0_bit31_8_reg[28]  <= n9345;
    \\configuration_pci_ba0_bit31_8_reg[30]  <= n9350;
    \\configuration_pci_ba0_bit31_8_reg[29]  <= n9355;
    \\pci_target_unit_wishbone_master_read_count_reg[1]  <= n9360;
    \\pci_target_unit_wishbone_master_read_count_reg[2]  <= n9365;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[0]  <= n9370;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[10]  <= n9375;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[11]  <= n9380;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[13]  <= n9385;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[15]  <= n9390;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[17]  <= n9395;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[18]  <= n9400;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[19]  <= n9405;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[20]  <= n9410;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[22]  <= n9415;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[24]  <= n9420;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[25]  <= n9425;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[26]  <= n9430;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[28]  <= n9435;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[29]  <= n9440;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[2]  <= n9445;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[3]  <= n9450;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[6]  <= n9455;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[9]  <= n9460;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[30]  <= n9465;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][37]  <= n9470;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][37]  <= n9475;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][37]  <= n9480;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][37]  <= n9485;
    wishbone_slave_unit_del_sync_comp_req_pending_reg <= n9490;
    \\configuration_pci_ba0_bit31_8_reg[31]  <= n9495;
    \\configuration_pci_ba0_bit31_8_reg[26]  <= n9500;
    \\configuration_pci_ba0_bit31_8_reg[24]  <= n9505;
    \\configuration_pci_ba0_bit31_8_reg[21]  <= n9510;
    \\configuration_pci_ba0_bit31_8_reg[22]  <= n9515;
    \\configuration_pci_am1_reg[16]  <= n9520;
    \\configuration_pci_am1_reg[15]  <= n9525;
    \\configuration_pci_am1_reg[24]  <= n9530;
    \\configuration_pci_ba1_bit31_8_reg[11]  <= n9535;
    \\configuration_pci_ba1_bit31_8_reg[15]  <= n9540;
    \\wishbone_slave_unit_pci_initiator_if_read_count_reg[3]  <= n9545;
    wishbone_slave_unit_wishbone_slave_map_reg <= n9550;
    \\configuration_pci_ba1_bit31_8_reg[18]  <= n9555;
    \\configuration_pci_ba1_bit31_8_reg[19]  <= n9560;
    \\configuration_pci_ba1_bit31_8_reg[20]  <= n9565;
    \\configuration_pci_ba1_bit31_8_reg[21]  <= n9570;
    \\configuration_pci_ba1_bit31_8_reg[23]  <= n9575;
    \\configuration_pci_ba1_bit31_8_reg[25]  <= n9580;
    \\configuration_pci_ba1_bit31_8_reg[26]  <= n9585;
    \\configuration_pci_ba1_bit31_8_reg[27]  <= n9590;
    \\configuration_pci_ba1_bit31_8_reg[29]  <= n9595;
    \\configuration_pci_ba1_bit31_8_reg[30]  <= n9600;
    \\configuration_pci_ba1_bit31_8_reg[10]  <= n9605;
    \\configuration_pci_ba1_bit31_8_reg[12]  <= n9610;
    \\configuration_pci_ba1_bit31_8_reg[13]  <= n9615;
    \\configuration_pci_ba1_bit31_8_reg[14]  <= n9620;
    \\configuration_pci_ba1_bit31_8_reg[16]  <= n9625;
    \\pci_target_unit_wishbone_master_c_state_reg[1]  <= n9630;
    \\configuration_pci_am1_reg[21]  <= n9635;
    \\configuration_pci_am1_reg[10]  <= n9640;
    \\configuration_pci_am1_reg[12]  <= n9645;
    \\configuration_pci_am1_reg[11]  <= n9650;
    \\configuration_pci_am1_reg[13]  <= n9655;
    \\configuration_pci_am1_reg[18]  <= n9660;
    \\configuration_pci_am1_reg[17]  <= n9665;
    \\configuration_pci_am1_reg[20]  <= n9670;
    \\configuration_pci_am1_reg[14]  <= n9675;
    \\configuration_pci_am1_reg[22]  <= n9680;
    \\configuration_pci_am1_reg[23]  <= n9685;
    \\configuration_pci_am1_reg[25]  <= n9690;
    \\configuration_pci_am1_reg[19]  <= n9695;
    \\configuration_pci_am1_reg[29]  <= n9700;
    \\configuration_pci_am1_reg[31]  <= n9705;
    \\configuration_pci_am1_reg[30]  <= n9710;
    \\configuration_pci_am1_reg[28]  <= n9715;
    \\pci_target_unit_wishbone_master_read_count_reg[0]  <= n9720;
    \\configuration_pci_ba1_bit31_8_reg[31]  <= n9725;
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[1]  <= n9730;
    \\configuration_pci_ba1_bit31_8_reg[8]  <= n9735;
    \\configuration_pci_ba1_bit31_8_reg[9]  <= n9740;
    \\configuration_pci_ba1_bit31_8_reg[22]  <= n9745;
    \\configuration_pci_ba1_bit31_8_reg[28]  <= n9750;
    \\configuration_pci_ba1_bit31_8_reg[24]  <= n9755;
    \\configuration_pci_ba1_bit31_8_reg[17]  <= n9760;
    wishbone_slave_unit_pci_initiator_if_current_last_reg <= n9765;
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[0]  <= n9770;
    \\configuration_pci_am1_reg[26]  <= n9775;
    \\configuration_pci_am1_reg[8]  <= n9780;
    \\configuration_pci_am1_reg[9]  <= n9785;
    \\configuration_pci_am1_reg[27]  <= n9790;
    \\wishbone_slave_unit_wishbone_slave_c_state_reg[1]  <= n9795;
    \\configuration_pci_ta1_reg[10]  <= n9800;
    pci_target_unit_wishbone_master_read_bound_reg <= n9805;
    \\configuration_pci_ta1_reg[29]  <= n9810;
    \\configuration_pci_ta1_reg[16]  <= n9815;
    \\wishbone_slave_unit_pci_initiator_if_read_count_reg[2]  <= n9820;
    \\configuration_pci_ta1_reg[17]  <= n9825;
    \\configuration_pci_ta1_reg[18]  <= n9830;
    \\configuration_pci_ta1_reg[20]  <= n9835;
    \\configuration_pci_ta1_reg[21]  <= n9840;
    \\configuration_pci_ta1_reg[24]  <= n9845;
    \\configuration_pci_ta1_reg[23]  <= n9850;
    \\configuration_pci_ta1_reg[30]  <= n9855;
    \\configuration_pci_ta1_reg[28]  <= n9860;
    \\configuration_pci_ta1_reg[31]  <= n9865;
    \\configuration_pci_ta1_reg[14]  <= n9870;
    wishbone_slave_unit_pci_initiator_if_err_recovery_reg <= n9875;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]  <= n9880;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][37]  <= n9885;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][37]  <= n9890;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][37]  <= n9895;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][37]  <= n9900;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][37]  <= n9905;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][37]  <= n9910;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][37]  <= n9915;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][37]  <= n9920;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][37]  <= n9925;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][37]  <= n9930;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][37]  <= n9935;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][37]  <= n9940;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][37]  <= n9945;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][37]  <= n9950;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][37]  <= n9955;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][37]  <= n9960;
    \\configuration_pci_ta1_reg[11]  <= n9965;
    \\configuration_pci_ta1_reg[13]  <= n9970;
    \\configuration_pci_ta1_reg[15]  <= n9975;
    \\configuration_pci_ta1_reg[12]  <= n9980;
    \\configuration_pci_ta1_reg[8]  <= n9985;
    \\configuration_pci_ta1_reg[9]  <= n9990;
    \\configuration_pci_ta1_reg[27]  <= n9995;
    \\configuration_pci_ta1_reg[26]  <= n10000;
    \\configuration_pci_ta1_reg[25]  <= n10005;
    \\configuration_pci_ta1_reg[22]  <= n10010;
    \\configuration_pci_ta1_reg[19]  <= n10015;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][32]  <= n10020;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][32]  <= n10025;
    wishbone_slave_unit_pci_initiator_if_posted_write_req_reg <= n10030;
    pci_io_mux_frame_iob_en_out_reg <= n10035;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[27]  <= n10040;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[17]  <= n10045;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[19]  <= n10050;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[20]  <= n10055;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[22]  <= n10060;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[23]  <= n10065;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[24]  <= n10070;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[28]  <= n10075;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[29]  <= n10080;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[2]  <= n10085;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[31]  <= n10090;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[3]  <= n10095;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[4]  <= n10100;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[6]  <= n10105;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[8]  <= n10110;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[16]  <= n10115;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[14]  <= n10120;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[0]  <= n10125;
    output_backup_cbe_en_out_reg <= n10130;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][32]  <= n10135;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][32]  <= n10140;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][32]  <= n10145;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][32]  <= n10150;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][36]  <= n10155;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][32]  <= n10160;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[13]  <= n10165;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[15]  <= n10170;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[9]  <= n10175;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[5]  <= n10180;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[7]  <= n10185;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][36]  <= n10190;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[26]  <= n10195;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[30]  <= n10200;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[18]  <= n10205;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[21]  <= n10210;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[1]  <= n10215;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[12]  <= n10220;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[25]  <= n10225;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[11]  <= n10230;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[0]  <= n10235;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[10]  <= n10240;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][36]  <= n10245;
    \\wishbone_slave_unit_pci_initiator_if_be_out_reg[1]  <= n10250;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][32]  <= n10255;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][36]  <= n10260;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][6]  <= n10265;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][4]  <= n10270;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][13]  <= n10275;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][3]  <= n10280;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][7]  <= n10285;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][9]  <= n10290;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][0]  <= n10295;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][19]  <= n10300;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][6]  <= n10305;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][15]  <= n10310;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][7]  <= n10315;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][16]  <= n10320;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][8]  <= n10325;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][17]  <= n10330;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][7]  <= n10335;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][30]  <= n10340;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][25]  <= n10345;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][0]  <= n10350;
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[4]  <= n10355;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][12]  <= n10360;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][3]  <= n10365;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][12]  <= n10370;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][10]  <= n10375;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][36]  <= n10380;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][11]  <= n10385;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][9]  <= n10390;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][2]  <= n10395;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][29]  <= n10400;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][8]  <= n10405;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][7]  <= n10410;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][8]  <= n10415;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][25]  <= n10420;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][23]  <= n10425;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][14]  <= n10430;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][6]  <= n10435;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][16]  <= n10440;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][27]  <= n10445;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][13]  <= n10450;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][28]  <= n10455;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][1]  <= n10460;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][25]  <= n10465;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][26]  <= n10470;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][23]  <= n10475;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][16]  <= n10480;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][16]  <= n10485;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][8]  <= n10490;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][12]  <= n10495;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][10]  <= n10500;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][9]  <= n10505;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][25]  <= n10510;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][31]  <= n10515;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][4]  <= n10520;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][22]  <= n10525;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][18]  <= n10530;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][27]  <= n10535;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][29]  <= n10540;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][21]  <= n10545;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][27]  <= n10550;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][23]  <= n10555;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][1]  <= n10560;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[16]  <= n10565;
    configuration_set_isr_bit2_reg <= n10570;
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[2]  <= n10575;
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[3]  <= n10580;
    wishbone_slave_unit_wishbone_slave_wb_conf_hit_reg <= n10585;
    \\configuration_wb_err_addr_reg[0]  <= n10590;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6]  <= n10595;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2]  <= n10600;
    output_backup_frame_en_out_reg <= n10605;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][0]  <= n10610;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][0]  <= n10615;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][0]  <= n10620;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][0]  <= n10625;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][1]  <= n10630;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][0]  <= n10635;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][0]  <= n10640;
    pci_io_mux_cbe_iob3_en_out_reg <= n10645;
    pci_io_mux_cbe_iob2_en_out_reg <= n10650;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]  <= n10655;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]  <= n10660;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]  <= n10665;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[3]  <= n10670;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][0]  <= n10675;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][10]  <= n10680;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][12]  <= n10685;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][14]  <= n10690;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][10]  <= n10695;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][16]  <= n10700;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][18]  <= n10705;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][1]  <= n10710;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][21]  <= n10715;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][23]  <= n10720;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][24]  <= n10725;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][25]  <= n10730;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][27]  <= n10735;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][28]  <= n10740;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][29]  <= n10745;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][30]  <= n10750;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][4]  <= n10755;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][6]  <= n10760;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][8]  <= n10765;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][0]  <= n10770;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][11]  <= n10775;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][13]  <= n10780;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][15]  <= n10785;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][17]  <= n10790;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][19]  <= n10795;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][20]  <= n10800;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][22]  <= n10805;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][24]  <= n10810;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][26]  <= n10815;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][28]  <= n10820;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][30]  <= n10825;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][2]  <= n10830;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][3]  <= n10835;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][5]  <= n10840;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][7]  <= n10845;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][0]  <= n10850;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][11]  <= n10855;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][13]  <= n10860;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][14]  <= n10865;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][15]  <= n10870;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][17]  <= n10875;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][18]  <= n10880;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][19]  <= n10885;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][20]  <= n10890;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][21]  <= n10895;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][22]  <= n10900;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][24]  <= n10905;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][2]  <= n10910;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][3]  <= n10915;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][5]  <= n10920;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][7]  <= n10925;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][9]  <= n10930;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][0]  <= n10935;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][11]  <= n10940;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][13]  <= n10945;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][15]  <= n10950;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][17]  <= n10955;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][18]  <= n10960;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][19]  <= n10965;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][20]  <= n10970;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][22]  <= n10975;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][24]  <= n10980;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][25]  <= n10985;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][26]  <= n10990;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][28]  <= n10995;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][2]  <= n11000;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][31]  <= n11005;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][3]  <= n11010;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][5]  <= n11015;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][6]  <= n11020;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][7]  <= n11025;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][9]  <= n11030;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][10]  <= n11035;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][12]  <= n11040;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][13]  <= n11045;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][14]  <= n11050;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][16]  <= n11055;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][1]  <= n11060;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][27]  <= n11065;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][31]  <= n11070;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][30]  <= n11075;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][4]  <= n11080;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][6]  <= n11085;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][8]  <= n11090;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][9]  <= n11095;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][0]  <= n11100;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][15]  <= n11105;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][19]  <= n11110;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][20]  <= n11115;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][22]  <= n11120;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][23]  <= n11125;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][24]  <= n11130;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][26]  <= n11135;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][28]  <= n11140;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][30]  <= n11145;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][2]  <= n11150;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][3]  <= n11155;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][5]  <= n11160;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][24]  <= n11165;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][7]  <= n11170;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][9]  <= n11175;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][10]  <= n11180;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][12]  <= n11185;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][14]  <= n11190;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][15]  <= n11195;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][16]  <= n11200;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][18]  <= n11205;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][19]  <= n11210;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][1]  <= n11215;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][21]  <= n11220;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][22]  <= n11225;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][23]  <= n11230;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][25]  <= n11235;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][27]  <= n11240;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][29]  <= n11245;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][2]  <= n11250;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][30]  <= n11255;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][4]  <= n11260;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][6]  <= n11265;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][8]  <= n11270;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][0]  <= n11275;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][11]  <= n11280;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][13]  <= n11285;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][14]  <= n11290;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][15]  <= n11295;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][17]  <= n11300;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][18]  <= n11305;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][19]  <= n11310;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][20]  <= n11315;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][21]  <= n11320;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][22]  <= n11325;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][24]  <= n11330;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][26]  <= n11335;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][28]  <= n11340;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][29]  <= n11345;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][2]  <= n11350;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][23]  <= n11355;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][9]  <= n11360;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][10]  <= n11365;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][12]  <= n11370;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][1]  <= n11375;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][21]  <= n11380;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][17]  <= n11385;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][27]  <= n11390;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][30]  <= n11395;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][4]  <= n11400;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][10]  <= n11405;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][12]  <= n11410;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][14]  <= n11415;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][16]  <= n11420;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][18]  <= n11425;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][19]  <= n11430;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][1]  <= n11435;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][21]  <= n11440;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][23]  <= n11445;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][25]  <= n11450;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][29]  <= n11455;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][4]  <= n11460;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][0]  <= n11465;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][13]  <= n11470;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][24]  <= n11475;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][26]  <= n11480;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][28]  <= n11485;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][29]  <= n11490;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][2]  <= n11495;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][3]  <= n11500;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][5]  <= n11505;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][6]  <= n11510;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][7]  <= n11515;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][9]  <= n11520;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][36]  <= n11525;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][36]  <= n11530;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][36]  <= n11535;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][36]  <= n11540;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][36]  <= n11545;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][14]  <= n11550;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][36]  <= n11555;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][36]  <= n11560;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][36]  <= n11565;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][13]  <= n11570;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][15]  <= n11575;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][19]  <= n11580;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][20]  <= n11585;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][24]  <= n11590;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][28]  <= n11595;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][31]  <= n11600;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][5]  <= n11605;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][9]  <= n11610;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][10]  <= n11615;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][14]  <= n11620;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][1]  <= n11625;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][23]  <= n11630;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][4]  <= n11635;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][27]  <= n11640;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][29]  <= n11645;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][4]  <= n11650;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][6]  <= n11655;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][8]  <= n11660;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][0]  <= n11665;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][19]  <= n11670;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][20]  <= n11675;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][22]  <= n11680;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][2]  <= n11685;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][31]  <= n11690;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][3]  <= n11695;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][5]  <= n11700;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][14]  <= n11705;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][18]  <= n11710;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][1]  <= n11715;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][25]  <= n11720;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][27]  <= n11725;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][29]  <= n11730;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][29]  <= n11735;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][30]  <= n11740;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][36]  <= n11745;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][36]  <= n11750;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][36]  <= n11755;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][10]  <= n11760;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][14]  <= n11765;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][18]  <= n11770;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][1]  <= n11775;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][23]  <= n11780;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][29]  <= n11785;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][36]  <= n11790;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][6]  <= n11795;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][16]  <= n11800;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][18]  <= n11805;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][30]  <= n11810;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][22]  <= n11815;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][21]  <= n11820;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][36]  <= n11825;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][1]  <= n11830;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][1]  <= n11835;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][26]  <= n11840;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][14]  <= n11845;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][27]  <= n11850;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][28]  <= n11855;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][10]  <= n11860;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][12]  <= n11865;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][24]  <= n11870;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][25]  <= n11875;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][0]  <= n11880;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][11]  <= n11885;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][21]  <= n11890;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][10]  <= n11895;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][23]  <= n11900;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][11]  <= n11905;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][16]  <= n11910;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][17]  <= n11915;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][18]  <= n11920;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][14]  <= n11925;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][12]  <= n11930;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][15]  <= n11935;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[14][13]  <= n11940;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][3]  <= n11945;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][8]  <= n11950;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][9]  <= n11955;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][14]  <= n11960;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][20]  <= n11965;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][9]  <= n11970;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][22]  <= n11975;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][5]  <= n11980;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][5]  <= n11985;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][5]  <= n11990;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][7]  <= n11995;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]  <= n12000;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][6]  <= n12005;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][7]  <= n12010;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][27]  <= n12015;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][19]  <= n12020;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][8]  <= n12025;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][4]  <= n12030;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][30]  <= n12035;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][31]  <= n12040;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][20]  <= n12045;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][1]  <= n12050;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][23]  <= n12055;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][25]  <= n12060;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][21]  <= n12065;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][22]  <= n12070;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][31]  <= n12075;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][3]  <= n12080;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][16]  <= n12085;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][10]  <= n12090;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][11]  <= n12095;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][12]  <= n12100;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][17]  <= n12105;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][24]  <= n12110;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][15]  <= n12115;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][31]  <= n12120;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][2]  <= n12125;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][5]  <= n12130;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][3]  <= n12135;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][18]  <= n12140;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][15]  <= n12145;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][17]  <= n12150;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][4]  <= n12155;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][1]  <= n12160;
    configuration_wb_err_cs_bit9_reg <= n12165;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][5]  <= n12170;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][23]  <= n12175;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][0]  <= n12180;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][0]  <= n12185;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][17]  <= n12190;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][26]  <= n12195;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][0]  <= n12200;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][1]  <= n12205;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[0]  <= n12210;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][1]  <= n12215;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][9]  <= n12220;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][36]  <= n12225;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][26]  <= n12230;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][25]  <= n12235;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][11]  <= n12240;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][17]  <= n12245;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][30]  <= n12250;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][7]  <= n12255;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][5]  <= n12260;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][24]  <= n12265;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][28]  <= n12270;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][18]  <= n12275;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][31]  <= n12280;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][26]  <= n12285;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][26]  <= n12290;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][7]  <= n12295;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][19]  <= n12300;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][20]  <= n12305;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][15]  <= n12310;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][2]  <= n12315;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][22]  <= n12320;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][28]  <= n12325;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][8]  <= n12330;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][19]  <= n12335;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][16]  <= n12340;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][24]  <= n12345;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][27]  <= n12350;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][3]  <= n12355;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][29]  <= n12360;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][13]  <= n12365;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][14]  <= n12370;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][2]  <= n12375;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][28]  <= n12380;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][20]  <= n12385;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][29]  <= n12390;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][7]  <= n12395;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][6]  <= n12400;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][10]  <= n12405;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][11]  <= n12410;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][20]  <= n12415;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][31]  <= n12420;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][1]  <= n12425;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][17]  <= n12430;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][27]  <= n12435;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][26]  <= n12440;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][26]  <= n12445;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][0]  <= n12450;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][9]  <= n12455;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][28]  <= n12460;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][18]  <= n12465;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][6]  <= n12470;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][20]  <= n12475;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][21]  <= n12480;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][13]  <= n12485;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][22]  <= n12490;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][5]  <= n12495;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][13]  <= n12500;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][3]  <= n12505;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[4][11]  <= n12510;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][17]  <= n12515;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[0][11]  <= n12520;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][4]  <= n12525;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[2]  <= n12530;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][18]  <= n12535;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][30]  <= n12540;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][6]  <= n12545;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][1]  <= n12550;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][7]  <= n12555;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][30]  <= n12560;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][13]  <= n12565;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][19]  <= n12570;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][8]  <= n12575;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][15]  <= n12580;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][4]  <= n12585;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][8]  <= n12590;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][17]  <= n12595;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][29]  <= n12600;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][27]  <= n12605;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][31]  <= n12610;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][11]  <= n12615;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][9]  <= n12620;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][31]  <= n12625;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][25]  <= n12630;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][15]  <= n12635;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][23]  <= n12640;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[8][0]  <= n12645;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][2]  <= n12650;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][31]  <= n12655;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[1]  <= n12660;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][5]  <= n12665;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][3]  <= n12670;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][16]  <= n12675;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][8]  <= n12680;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][10]  <= n12685;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][25]  <= n12690;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][29]  <= n12695;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][0]  <= n12700;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][36]  <= n12705;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][27]  <= n12710;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][31]  <= n12715;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][4]  <= n12720;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][20]  <= n12725;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][28]  <= n12730;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][25]  <= n12735;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[3][21]  <= n12740;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][3]  <= n12745;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][27]  <= n12750;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[5][12]  <= n12755;
    pci_io_mux_cbe_iob1_en_out_reg <= n12760;
    pci_io_mux_cbe_iob0_en_out_reg <= n12765;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][2]  <= n12770;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][29]  <= n12775;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][30]  <= n12780;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][30]  <= n12785;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][30]  <= n12790;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][31]  <= n12795;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][21]  <= n12800;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][2]  <= n12805;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][20]  <= n12810;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][25]  <= n12815;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][23]  <= n12820;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][12]  <= n12825;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][24]  <= n12830;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][12]  <= n12835;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][1]  <= n12840;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][21]  <= n12845;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][22]  <= n12850;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][14]  <= n12855;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][16]  <= n12860;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[11][26]  <= n12865;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[1][10]  <= n12870;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][13]  <= n12875;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][19]  <= n12880;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][8]  <= n12885;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][17]  <= n12890;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][4]  <= n12895;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][1]  <= n12900;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][6]  <= n12905;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][1]  <= n12910;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][15]  <= n12915;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][1]  <= n12920;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][16]  <= n12925;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][9]  <= n12930;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][11]  <= n12935;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[7][0]  <= n12940;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[2][36]  <= n12945;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][31]  <= n12950;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][6]  <= n12955;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][7]  <= n12960;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][28]  <= n12965;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][26]  <= n12970;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][8]  <= n12975;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][5]  <= n12980;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][3]  <= n12985;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][2]  <= n12990;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][4]  <= n12995;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][28]  <= n13000;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][22]  <= n13005;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][26]  <= n13010;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][11]  <= n13015;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][24]  <= n13020;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][21]  <= n13025;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][21]  <= n13030;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][11]  <= n13035;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[9][12]  <= n13040;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]  <= n13045;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][12]  <= n13050;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]  <= n13055;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][22]  <= n13060;
    i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg <= n13065;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][18]  <= n13070;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][1]  <= n13075;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[12][36]  <= n13080;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][20]  <= n13085;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][23]  <= n13090;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][13]  <= n13095;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][19]  <= n13100;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[15][24]  <= n13105;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[10][36]  <= n13110;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[6][36]  <= n13115;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][17]  <= n13120;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][15]  <= n13125;
    \\wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg[13][16]  <= n13130;
    \\configuration_wb_err_addr_reg[11]  <= n13135;
    \\configuration_wb_err_data_reg[0]  <= n13140;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][20]  <= n13145;
    \\configuration_wb_err_cs_bit31_24_reg[30]  <= n13150;
    \\configuration_wb_err_addr_reg[19]  <= n13155;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][25]  <= n13160;
    \\configuration_pci_err_data_reg[28]  <= n13165;
    wishbone_slave_unit_pci_initiator_if_data_source_reg <= n13170;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][9]  <= n13175;
    \\configuration_wb_err_cs_bit31_24_reg[28]  <= n13180;
    \\configuration_wb_err_addr_reg[15]  <= n13185;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][16]  <= n13190;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][4]  <= n13195;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][14]  <= n13200;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][22]  <= n13205;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][4]  <= n13210;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][30]  <= n13215;
    \\configuration_wb_err_data_reg[6]  <= n13220;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][21]  <= n13225;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][24]  <= n13230;
    \\configuration_wb_err_data_reg[8]  <= n13235;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][27]  <= n13240;
    \\configuration_wb_err_data_reg[30]  <= n13245;
    \\configuration_wb_err_data_reg[4]  <= n13250;
    \\configuration_wb_err_data_reg[31]  <= n13255;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][15]  <= n13260;
    \\configuration_wb_err_data_reg[28]  <= n13265;
    \\configuration_wb_err_data_reg[27]  <= n13270;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][29]  <= n13275;
    \\configuration_wb_err_data_reg[24]  <= n13280;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][23]  <= n13285;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][22]  <= n13290;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][18]  <= n13295;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][21]  <= n13300;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][21]  <= n13305;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][16]  <= n13310;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][12]  <= n13315;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][35]  <= n13320;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][26]  <= n13325;
    \\configuration_wb_err_data_reg[20]  <= n13330;
    wishbone_slave_unit_pci_initiator_if_read_bound_reg <= n13335;
    configuration_pci_err_cs_bit9_reg <= n13340;
    configuration_pci_err_cs_bit10_reg <= n13345;
    \\configuration_pci_err_cs_bit31_24_reg[30]  <= n13350;
    \\configuration_pci_err_cs_bit31_24_reg[28]  <= n13355;
    \\configuration_pci_err_cs_bit31_24_reg[29]  <= n13360;
    \\wishbone_slave_unit_pci_initiator_if_read_count_reg[1]  <= n13365;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4]  <= n13370;
    \\configuration_pci_err_addr_reg[0]  <= n13375;
    \\configuration_pci_err_addr_reg[11]  <= n13380;
    \\configuration_pci_err_addr_reg[12]  <= n13385;
    \\configuration_pci_err_addr_reg[15]  <= n13390;
    \\configuration_pci_err_addr_reg[19]  <= n13395;
    \\configuration_pci_err_addr_reg[20]  <= n13400;
    \\configuration_pci_err_addr_reg[22]  <= n13405;
    \\configuration_pci_err_addr_reg[26]  <= n13410;
    \\configuration_pci_err_addr_reg[28]  <= n13415;
    \\configuration_pci_err_addr_reg[2]  <= n13420;
    \\configuration_pci_err_addr_reg[31]  <= n13425;
    \\configuration_pci_err_addr_reg[4]  <= n13430;
    \\configuration_pci_err_addr_reg[6]  <= n13435;
    \\configuration_pci_err_addr_reg[8]  <= n13440;
    \\configuration_pci_err_data_reg[0]  <= n13445;
    \\configuration_pci_err_data_reg[11]  <= n13450;
    \\configuration_pci_err_data_reg[13]  <= n13455;
    \\configuration_pci_err_data_reg[15]  <= n13460;
    \\configuration_pci_err_data_reg[17]  <= n13465;
    \\configuration_pci_err_data_reg[19]  <= n13470;
    \\configuration_pci_err_data_reg[21]  <= n13475;
    \\configuration_pci_err_data_reg[25]  <= n13480;
    \\configuration_pci_err_data_reg[29]  <= n13485;
    \\configuration_pci_err_data_reg[31]  <= n13490;
    \\configuration_pci_err_data_reg[3]  <= n13495;
    \\configuration_pci_err_data_reg[7]  <= n13500;
    pci_target_unit_pci_target_sm_same_read_reg_reg <= n13505;
    \\configuration_wb_err_cs_bit31_24_reg[25]  <= n13510;
    \\configuration_wb_err_cs_bit31_24_reg[31]  <= n13515;
    \\configuration_wb_err_data_reg[10]  <= n13520;
    \\configuration_wb_err_data_reg[11]  <= n13525;
    \\configuration_wb_err_data_reg[12]  <= n13530;
    \\configuration_wb_err_data_reg[14]  <= n13535;
    \\configuration_wb_err_data_reg[15]  <= n13540;
    \\configuration_wb_err_data_reg[16]  <= n13545;
    \\configuration_wb_err_data_reg[18]  <= n13550;
    \\configuration_wb_err_data_reg[19]  <= n13555;
    \\configuration_wb_err_data_reg[1]  <= n13560;
    \\configuration_wb_err_data_reg[21]  <= n13565;
    \\configuration_wb_err_data_reg[22]  <= n13570;
    \\configuration_wb_err_data_reg[23]  <= n13575;
    \\configuration_wb_err_data_reg[25]  <= n13580;
    \\configuration_wb_err_data_reg[26]  <= n13585;
    \\configuration_wb_err_data_reg[29]  <= n13590;
    \\configuration_wb_err_data_reg[2]  <= n13595;
    \\configuration_wb_err_data_reg[3]  <= n13600;
    \\configuration_wb_err_data_reg[5]  <= n13605;
    \\configuration_wb_err_data_reg[9]  <= n13610;
    \\configuration_wb_err_data_reg[7]  <= n13615;
    \\configuration_wb_err_addr_reg[10]  <= n13620;
    \\configuration_wb_err_addr_reg[12]  <= n13625;
    \\configuration_wb_err_addr_reg[13]  <= n13630;
    \\configuration_wb_err_addr_reg[14]  <= n13635;
    \\configuration_wb_err_addr_reg[16]  <= n13640;
    \\configuration_wb_err_addr_reg[18]  <= n13645;
    \\configuration_wb_err_addr_reg[20]  <= n13650;
    \\configuration_wb_err_addr_reg[22]  <= n13655;
    \\configuration_wb_err_addr_reg[24]  <= n13660;
    \\configuration_wb_err_addr_reg[26]  <= n13665;
    \\configuration_wb_err_addr_reg[28]  <= n13670;
    \\configuration_wb_err_addr_reg[2]  <= n13675;
    \\configuration_wb_err_addr_reg[31]  <= n13680;
    \\configuration_wb_err_addr_reg[4]  <= n13685;
    \\configuration_wb_err_addr_reg[6]  <= n13690;
    \\configuration_wb_err_addr_reg[7]  <= n13695;
    \\configuration_wb_err_addr_reg[8]  <= n13700;
    \\pci_target_unit_fifos_pciw_inTransactionCount_reg[1]  <= n13705;
    \\pci_target_unit_fifos_inGreyCount_reg[0]  <= n13710;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][17]  <= n13715;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][12]  <= n13720;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][11]  <= n13725;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][20]  <= n13730;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][7]  <= n13735;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][24]  <= n13740;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][3]  <= n13745;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][34]  <= n13750;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][33]  <= n13755;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][15]  <= n13760;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][29]  <= n13765;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][11]  <= n13770;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][13]  <= n13775;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][15]  <= n13780;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][17]  <= n13785;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][20]  <= n13790;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][23]  <= n13795;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][25]  <= n13800;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][28]  <= n13805;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][18]  <= n13810;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][30]  <= n13815;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][34]  <= n13820;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][35]  <= n13825;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][5]  <= n13830;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][7]  <= n13835;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][10]  <= n13840;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][12]  <= n13845;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][17]  <= n13850;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][22]  <= n13855;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][24]  <= n13860;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][31]  <= n13865;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][8]  <= n13870;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][16]  <= n13875;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][19]  <= n13880;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][22]  <= n13885;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][26]  <= n13890;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][2]  <= n13895;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][34]  <= n13900;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][33]  <= n13905;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][5]  <= n13910;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][7]  <= n13915;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][9]  <= n13920;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][14]  <= n13925;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][10]  <= n13930;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][17]  <= n13935;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][20]  <= n13940;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][22]  <= n13945;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][24]  <= n13950;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][23]  <= n13955;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][21]  <= n13960;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][25]  <= n13965;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][12]  <= n13970;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][34]  <= n13975;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][5]  <= n13980;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][7]  <= n13985;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][16]  <= n13990;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][23]  <= n13995;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][21]  <= n14000;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][14]  <= n14005;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][11]  <= n14010;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][13]  <= n14015;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][15]  <= n14020;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][17]  <= n14025;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][19]  <= n14030;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][27]  <= n14035;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][2]  <= n14040;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][3]  <= n14045;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][4]  <= n14050;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][6]  <= n14055;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][7]  <= n14060;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][16]  <= n14065;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][20]  <= n14070;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][22]  <= n14075;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][27]  <= n14080;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][29]  <= n14085;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][33]  <= n14090;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][6]  <= n14095;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][8]  <= n14100;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][10]  <= n14105;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][14]  <= n14110;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][9]  <= n14115;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][19]  <= n14120;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][23]  <= n14125;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][28]  <= n14130;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][8]  <= n14135;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][11]  <= n14140;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][21]  <= n14145;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][24]  <= n14150;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][27]  <= n14155;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][2]  <= n14160;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][18]  <= n14165;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][29]  <= n14170;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][35]  <= n14175;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][26]  <= n14180;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][38]  <= n14185;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][38]  <= n14190;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][38]  <= n14195;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][38]  <= n14200;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][13]  <= n14205;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][18]  <= n14210;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][13]  <= n14215;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][25]  <= n14220;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][19]  <= n14225;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][15]  <= n14230;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][20]  <= n14235;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][28]  <= n14240;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][12]  <= n14245;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][14]  <= n14250;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][9]  <= n14255;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][18]  <= n14260;
    \\configuration_wb_err_cs_bit31_24_reg[29]  <= n14265;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][33]  <= n14270;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][27]  <= n14275;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][6]  <= n14280;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][35]  <= n14285;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][5]  <= n14290;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][6]  <= n14295;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][6]  <= n14300;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][3]  <= n14305;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][8]  <= n14310;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][23]  <= n14315;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][22]  <= n14320;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][4]  <= n14325;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][9]  <= n14330;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][6]  <= n14335;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][15]  <= n14340;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][30]  <= n14345;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][8]  <= n14350;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][11]  <= n14355;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][13]  <= n14360;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][9]  <= n14365;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][14]  <= n14370;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][19]  <= n14375;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][4]  <= n14380;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][3]  <= n14385;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][33]  <= n14390;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][2]  <= n14395;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][31]  <= n14400;
    \\configuration_wb_err_data_reg[13]  <= n14405;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][27]  <= n14410;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][29]  <= n14415;
    \\configuration_wb_err_cs_bit31_24_reg[24]  <= n14420;
    \\configuration_wb_err_cs_bit31_24_reg[27]  <= n14425;
    \\configuration_wb_err_cs_bit31_24_reg[26]  <= n14430;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][12]  <= n14435;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][3]  <= n14440;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][10]  <= n14445;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][7]  <= n14450;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][4]  <= n14455;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][29]  <= n14460;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][11]  <= n14465;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][28]  <= n14470;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][5]  <= n14475;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][16]  <= n14480;
    \\configuration_wb_err_data_reg[17]  <= n14485;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][4]  <= n14490;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][31]  <= n14495;
    \\configuration_pci_err_data_reg[2]  <= n14500;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][35]  <= n14505;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][31]  <= n14510;
    \\configuration_wb_err_addr_reg[1]  <= n14515;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][22]  <= n14520;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[7]  <= n14525;
    pci_target_unit_pci_target_if_same_read_reg_reg <= n14530;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][34]  <= n14535;
    \\configuration_pci_err_data_reg[8]  <= n14540;
    \\configuration_pci_err_data_reg[30]  <= n14545;
    \\configuration_pci_err_data_reg[9]  <= n14550;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][13]  <= n14555;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][20]  <= n14560;
    \\configuration_pci_err_data_reg[5]  <= n14565;
    \\configuration_pci_err_data_reg[6]  <= n14570;
    \\configuration_pci_err_data_reg[4]  <= n14575;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][6]  <= n14580;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][2]  <= n14585;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][30]  <= n14590;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][23]  <= n14595;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][4]  <= n14600;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][26]  <= n14605;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][7]  <= n14610;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][24]  <= n14615;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][26]  <= n14620;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][31]  <= n14625;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][29]  <= n14630;
    \\configuration_pci_err_data_reg[23]  <= n14635;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][26]  <= n14640;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][25]  <= n14645;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][23]  <= n14650;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][5]  <= n14655;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][10]  <= n14660;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][31]  <= n14665;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][2]  <= n14670;
    \\configuration_wb_err_addr_reg[17]  <= n14675;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][25]  <= n14680;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][9]  <= n14685;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][6]  <= n14690;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][24]  <= n14695;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][8]  <= n14700;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][17]  <= n14705;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][31]  <= n14710;
    \\configuration_pci_err_data_reg[24]  <= n14715;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][33]  <= n14720;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][9]  <= n14725;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][18]  <= n14730;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][21]  <= n14735;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][19]  <= n14740;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][33]  <= n14745;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][10]  <= n14750;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][15]  <= n14755;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][3]  <= n14760;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][15]  <= n14765;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][14]  <= n14770;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][34]  <= n14775;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][11]  <= n14780;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][12]  <= n14785;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][34]  <= n14790;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][13]  <= n14795;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][8]  <= n14800;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][19]  <= n14805;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][25]  <= n14810;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][17]  <= n14815;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][30]  <= n14820;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][5]  <= n14825;
    \\configuration_pci_err_data_reg[26]  <= n14830;
    \\configuration_pci_err_data_reg[27]  <= n14835;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][34]  <= n14840;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][35]  <= n14845;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][28]  <= n14850;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][35]  <= n14855;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][38]  <= n14860;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][28]  <= n14865;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][16]  <= n14870;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][26]  <= n14875;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][27]  <= n14880;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][10]  <= n14885;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][7]  <= n14890;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][8]  <= n14895;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][18]  <= n14900;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][18]  <= n14905;
    \\configuration_pci_err_addr_reg[7]  <= n14910;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][20]  <= n14915;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][38]  <= n14920;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][14]  <= n14925;
    \\configuration_pci_err_addr_reg[9]  <= n14930;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][12]  <= n14935;
    \\configuration_pci_err_data_reg[18]  <= n14940;
    \\configuration_pci_err_data_reg[1]  <= n14945;
    \\configuration_pci_err_data_reg[20]  <= n14950;
    \\configuration_pci_err_data_reg[22]  <= n14955;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][10]  <= n14960;
    \\configuration_pci_err_data_reg[14]  <= n14965;
    \\configuration_pci_err_cs_bit31_24_reg[24]  <= n14970;
    \\configuration_pci_err_data_reg[16]  <= n14975;
    \\configuration_pci_err_cs_bit31_24_reg[25]  <= n14980;
    \\configuration_pci_err_data_reg[10]  <= n14985;
    \\configuration_pci_err_data_reg[12]  <= n14990;
    \\configuration_pci_err_cs_bit31_24_reg[26]  <= n14995;
    \\configuration_pci_err_cs_bit31_24_reg[27]  <= n15000;
    \\configuration_pci_err_addr_reg[3]  <= n15005;
    \\configuration_pci_err_addr_reg[10]  <= n15010;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][5]  <= n15015;
    \\configuration_wb_err_addr_reg[21]  <= n15020;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][38]  <= n15025;
    \\configuration_pci_err_addr_reg[5]  <= n15030;
    \\configuration_pci_err_addr_reg[30]  <= n15035;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][11]  <= n15040;
    \\configuration_pci_err_addr_reg[27]  <= n15045;
    \\configuration_pci_err_addr_reg[29]  <= n15050;
    \\configuration_pci_err_addr_reg[25]  <= n15055;
    \\configuration_pci_err_addr_reg[1]  <= n15060;
    \\configuration_pci_err_addr_reg[23]  <= n15065;
    \\configuration_pci_err_addr_reg[24]  <= n15070;
    \\configuration_pci_err_addr_reg[21]  <= n15075;
    \\configuration_pci_err_addr_reg[13]  <= n15080;
    \\configuration_pci_err_addr_reg[18]  <= n15085;
    \\configuration_pci_err_addr_reg[17]  <= n15090;
    \\configuration_pci_err_addr_reg[14]  <= n15095;
    \\configuration_pci_err_addr_reg[16]  <= n15100;
    \\configuration_pci_err_cs_bit31_24_reg[31]  <= n15105;
    \\wishbone_slave_unit_pci_initiator_if_read_count_reg[0]  <= n15110;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][3]  <= n15115;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][25]  <= n15120;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][33]  <= n15125;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][31]  <= n15130;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][2]  <= n15135;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][24]  <= n15140;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][13]  <= n15145;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][21]  <= n15150;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][26]  <= n15155;
    \\configuration_wb_err_addr_reg[9]  <= n15160;
    \\configuration_wb_err_addr_reg[5]  <= n15165;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][30]  <= n15170;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][30]  <= n15175;
    \\configuration_wb_err_addr_reg[3]  <= n15180;
    \\configuration_wb_err_addr_reg[23]  <= n15185;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][27]  <= n15190;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][30]  <= n15195;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][28]  <= n15200;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][29]  <= n15205;
    \\configuration_wb_err_addr_reg[30]  <= n15210;
    \\configuration_wb_err_addr_reg[29]  <= n15215;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][19]  <= n15220;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][35]  <= n15225;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][16]  <= n15230;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][28]  <= n15235;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][17]  <= n15240;
    \\configuration_wb_err_addr_reg[25]  <= n15245;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][2]  <= n15250;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][3]  <= n15255;
    \\configuration_wb_err_addr_reg[27]  <= n15260;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][38]  <= n15265;
    \\pci_target_unit_fifos_pciw_inTransactionCount_reg[0]  <= n15270;
    \\pci_target_unit_fifos_inGreyCount_reg[1]  <= n15275;
    pci_target_unit_del_sync_comp_rty_exp_reg_reg <= n15280;
    \\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2]  <= n15285;
    configuration_set_pci_err_cs_bit8_reg <= n15290;
    wishbone_slave_unit_pci_initiator_if_del_write_req_reg <= n15295;
    pci_target_unit_wishbone_master_wb_read_done_out_reg <= n15300;
    pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg <= n15305;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[0]  <= n15310;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]  <= n15315;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[0]  <= n15320;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]  <= n15325;
    pci_target_unit_del_sync_req_done_reg_reg <= n15330;
    \\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1]  <= n15335;
    \\pci_target_unit_pci_target_if_strd_address_reg[2]  <= n15340;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1]  <= n15345;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]  <= n15350;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]  <= n15355;
    wishbone_slave_unit_pci_initiator_sm_timeout_reg <= n15360;
    \\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0]  <= n15365;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[3][39]  <= n15370;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[1][39]  <= n15375;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[7][39]  <= n15380;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[2][39]  <= n15385;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[0][39]  <= n15390;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[5][39]  <= n15395;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[6][39]  <= n15400;
    \\pci_target_unit_fifos_pciw_fifo_storage_mem_reg[4][39]  <= n15405;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[2]  <= n15410;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[0]  <= n15415;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[2]  <= n15420;
    pci_target_unit_pci_target_sm_wr_to_fifo_reg <= n15425;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0]  <= n15430;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[15]  <= n15435;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[2]  <= n15440;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1]  <= n15445;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[2]  <= n15450;
    pci_target_unit_del_sync_req_comp_pending_reg <= n15455;
    wishbone_slave_unit_pci_initiator_sm_transfer_reg <= n15460;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[1]  <= n15465;
    \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[1]  <= n15470;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[14]  <= n15475;
    wishbone_slave_unit_del_sync_comp_rty_exp_reg_reg <= n15480;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]  <= n15485;
    parity_checker_check_for_serr_on_second_reg <= n15490;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[1]  <= n15495;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[2]  <= n15500;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2]  <= n15505;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[1]  <= n15510;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[0]  <= n15515;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[0]  <= n15520;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[12]  <= n15525;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[1]  <= n15530;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[3]  <= n15535;
    i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg <= n15540;
    pci_target_unit_pci_target_if_target_rd_reg <= n15545;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[11]  <= n15550;
    pci_target_unit_pci_target_sm_rd_from_fifo_reg <= n15555;
    pci_resets_and_interrupts_inta_en_out_reg <= n15560;
    \\pci_target_unit_pci_target_if_norm_bc_reg[0]  <= n15565;
    \\pci_target_unit_pci_target_if_strd_address_reg[3]  <= n15570;
    pci_target_unit_wishbone_master_retried_reg <= n15575;
    pci_target_unit_wishbone_master_pcir_fifo_wenable_out_reg <= n15580;
    pci_target_unit_pci_target_sm_rw_cbe0_reg <= n15585;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[10]  <= n15590;
    \\pci_target_unit_del_sync_be_out_reg[0]  <= n15595;
    \\input_register_pci_cbe_reg_out_reg[0]  <= n15600;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[8]  <= n15605;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[13]  <= n15610;
    wishbone_slave_unit_pci_initiator_if_last_transfered_reg <= n15615;
    \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[0]  <= n15620;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[7]  <= n15625;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[9]  <= n15630;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[4]  <= n15635;
    \\pci_target_unit_pci_target_if_strd_address_reg[1]  <= n15640;
    \\pci_target_unit_pci_target_if_strd_address_reg[8]  <= n15645;
    \\pci_target_unit_pci_target_if_strd_address_reg[6]  <= n15650;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[6]  <= n15655;
    pci_target_unit_pci_target_sm_cnf_progress_reg <= n15660;
    wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg <= n15665;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[3]  <= n15670;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[0]  <= n15675;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[1]  <= n15680;
    wishbone_slave_unit_pci_initiator_if_rdy_out_reg <= n15685;
    \\pci_target_unit_pci_target_if_norm_address_reg[1]  <= n15690;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[2]  <= n15695;
    \\pci_target_unit_pci_target_if_norm_address_reg[3]  <= n15700;
    \\pci_target_unit_pci_target_if_norm_bc_reg[1]  <= n15705;
    \\pci_target_unit_wishbone_master_pcir_fifo_control_out_reg[1]  <= n15710;
    \\pci_target_unit_pci_target_if_strd_address_reg[4]  <= n15715;
    \\pci_target_unit_pci_target_if_strd_address_reg[7]  <= n15720;
    \\pci_target_unit_pci_target_if_strd_address_reg[9]  <= n15725;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[5]  <= n15730;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[1]  <= n15735;
    \\pci_target_unit_pci_target_if_norm_address_reg[6]  <= n15740;
    \\pci_target_unit_pci_target_if_strd_address_reg[5]  <= n15745;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[0]  <= n15750;
    \\pci_target_unit_pci_target_if_norm_address_reg[2]  <= n15755;
    \\pci_target_unit_pci_target_if_norm_address_reg[11]  <= n15760;
    \\pci_target_unit_del_sync_addr_out_reg[22]  <= n15765;
    \\pci_target_unit_del_sync_addr_out_reg[21]  <= n15770;
    \\pci_target_unit_del_sync_bc_out_reg[1]  <= n15775;
    \\pci_target_unit_pci_target_if_norm_address_reg[16]  <= n15780;
    \\pci_target_unit_pci_target_if_norm_address_reg[22]  <= n15785;
    \\pci_target_unit_pci_target_if_norm_address_reg[23]  <= n15790;
    \\pci_target_unit_pci_target_if_norm_address_reg[24]  <= n15795;
    \\pci_target_unit_pci_target_if_norm_address_reg[25]  <= n15800;
    \\pci_target_unit_del_sync_addr_out_reg[16]  <= n15805;
    \\pci_target_unit_pci_target_if_norm_address_reg[17]  <= n15810;
    \\pci_target_unit_pci_target_if_norm_address_reg[10]  <= n15815;
    \\pci_target_unit_del_sync_be_out_reg[1]  <= n15820;
    \\pci_target_unit_pci_target_if_norm_address_reg[30]  <= n15825;
    \\input_register_pci_cbe_reg_out_reg[3]  <= n15830;
    \\pci_target_unit_pci_target_if_norm_address_reg[14]  <= n15835;
    \\input_register_pci_cbe_reg_out_reg[2]  <= n15840;
    \\pci_target_unit_pci_target_if_norm_address_reg[28]  <= n15845;
    \\pci_target_unit_pci_target_if_norm_address_reg[27]  <= n15850;
    \\pci_target_unit_pci_target_if_norm_address_reg[13]  <= n15855;
    \\pci_target_unit_pci_target_if_norm_bc_reg[3]  <= n15860;
    \\pci_target_unit_pci_target_if_norm_bc_reg[2]  <= n15865;
    \\pci_target_unit_del_sync_addr_out_reg[2]  <= n15870;
    wishbone_slave_unit_pci_initiator_sm_mabort1_reg <= n15875;
    \\pci_target_unit_del_sync_addr_out_reg[26]  <= n15880;
    \\pci_target_unit_del_sync_addr_out_reg[25]  <= n15885;
    \\pci_target_unit_del_sync_addr_out_reg[24]  <= n15890;
    \\pci_target_unit_del_sync_addr_out_reg[23]  <= n15895;
    \\pci_target_unit_del_sync_addr_out_reg[28]  <= n15900;
    \\pci_target_unit_del_sync_addr_out_reg[20]  <= n15905;
    pci_target_unit_del_sync_burst_out_reg <= n15910;
    \\pci_target_unit_del_sync_addr_out_reg[4]  <= n15915;
    \\pci_target_unit_pci_target_if_norm_address_reg[5]  <= n15920;
    \\pci_target_unit_del_sync_addr_out_reg[7]  <= n15925;
    \\pci_target_unit_pci_target_if_norm_address_reg[21]  <= n15930;
    \\pci_target_unit_pci_target_if_norm_address_reg[12]  <= n15935;
    \\pci_target_unit_pci_target_if_norm_address_reg[31]  <= n15940;
    \\pci_target_unit_pci_target_if_norm_address_reg[26]  <= n15945;
    input_register_pci_trdy_reg_out_reg <= n15950;
    \\pci_target_unit_pci_target_if_norm_address_reg[15]  <= n15955;
    \\pci_target_unit_del_sync_addr_out_reg[27]  <= n15960;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[13]  <= n15965;
    \\pci_target_unit_del_sync_addr_out_reg[9]  <= n15970;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[21]  <= n15975;
    \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[3]  <= n15980;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[20]  <= n15985;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[27]  <= n15990;
    \\pci_target_unit_del_sync_addr_out_reg[31]  <= n15995;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[8]  <= n16000;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[4]  <= n16005;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[6]  <= n16010;
    \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[1]  <= n16015;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[29]  <= n16020;
    \\input_register_pci_cbe_reg_out_reg[1]  <= n16025;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[30]  <= n16030;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[26]  <= n16035;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[22]  <= n16040;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[18]  <= n16045;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[12]  <= n16050;
    \\pci_target_unit_pci_target_if_norm_address_reg[29]  <= n16055;
    \\pci_target_unit_del_sync_be_out_reg[2]  <= n16060;
    \\pci_target_unit_pci_target_if_norm_address_reg[20]  <= n16065;
    \\pci_target_unit_del_sync_addr_out_reg[1]  <= n16070;
    \\pci_target_unit_del_sync_addr_out_reg[14]  <= n16075;
    \\pci_target_unit_del_sync_addr_out_reg[6]  <= n16080;
    \\pci_target_unit_del_sync_addr_out_reg[11]  <= n16085;
    \\pci_target_unit_del_sync_be_out_reg[3]  <= n16090;
    wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg <= n16095;
    \\pci_target_unit_del_sync_addr_out_reg[19]  <= n16100;
    \\pci_target_unit_del_sync_addr_out_reg[15]  <= n16105;
    \\pci_target_unit_del_sync_addr_out_reg[30]  <= n16110;
    \\pci_target_unit_del_sync_addr_out_reg[8]  <= n16115;
    \\pci_target_unit_del_sync_addr_out_reg[3]  <= n16120;
    \\pci_target_unit_pci_target_if_norm_address_reg[19]  <= n16125;
    \\pci_target_unit_del_sync_addr_out_reg[13]  <= n16130;
    \\pci_target_unit_pci_target_if_norm_address_reg[18]  <= n16135;
    \\pci_target_unit_del_sync_addr_out_reg[12]  <= n16140;
    \\pci_target_unit_del_sync_addr_out_reg[10]  <= n16145;
    \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]  <= n16150;
    pci_target_unit_pci_target_sm_state_backoff_reg_reg <= n16155;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[10]  <= n16160;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[11]  <= n16165;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[16]  <= n16170;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[19]  <= n16175;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[23]  <= n16180;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[28]  <= n16185;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[2]  <= n16190;
    \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[2]  <= n16195;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[3]  <= n16200;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[5]  <= n16205;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[7]  <= n16210;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[9]  <= n16215;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[31]  <= n16220;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[24]  <= n16225;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[14]  <= n16230;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[15]  <= n16235;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[25]  <= n16240;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[17]  <= n16245;
    \\pci_target_unit_del_sync_bc_out_reg[3]  <= n16250;
    \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[2]  <= n16255;
    \\pci_target_unit_pci_target_if_norm_address_reg[9]  <= n16260;
    \\pci_target_unit_del_sync_addr_out_reg[5]  <= n16265;
    \\pci_target_unit_pci_target_if_norm_address_reg[4]  <= n16270;
    \\pci_target_unit_pci_target_if_norm_address_reg[0]  <= n16275;
    \\pci_target_unit_pci_target_if_norm_address_reg[8]  <= n16280;
    \\pci_target_unit_pci_target_if_strd_address_reg[0]  <= n16285;
    \\pci_target_unit_pci_target_if_norm_address_reg[7]  <= n16290;
    \\pci_target_unit_del_sync_bc_out_reg[0]  <= n16295;
    \\pci_target_unit_del_sync_bc_out_reg[2]  <= n16300;
    \\pci_target_unit_del_sync_addr_out_reg[29]  <= n16305;
    \\pci_target_unit_del_sync_addr_out_reg[18]  <= n16310;
    \\pci_target_unit_del_sync_addr_out_reg[0]  <= n16315;
    \\pci_target_unit_del_sync_addr_out_reg[17]  <= n16320;
    input_register_pci_frame_reg_out_reg <= n16325;
    input_register_pci_devsel_reg_out_reg <= n16330;
    pci_io_mux_irdy_iob_dat_out_reg <= n16335;
    input_register_pci_irdy_reg_out_reg <= n16340;
    output_backup_irdy_out_reg <= n16345;
    \\wishbone_slave_unit_del_sync_rty_exp_back_prop_sync_sync_data_out_reg[0]  <= n16350;
    pci_target_unit_del_sync_req_req_pending_reg <= n16355;
    input_register_pci_stop_reg_out_reg <= n16360;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[8]  <= n16365;
    configuration_interrupt_out_reg <= n16370;
    pci_io_mux_req_iob_dat_out_reg <= n16375;
    \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[3]  <= n16380;
    pci_target_unit_pci_target_sm_state_transfere_reg_reg <= n16385;
    pci_target_unit_pci_target_sm_previous_frame_reg <= n16390;
    \\input_register_pci_ad_reg_out_reg[7]  <= n16395;
    \\input_register_pci_ad_reg_out_reg[17]  <= n16400;
    \\input_register_pci_ad_reg_out_reg[30]  <= n16405;
    \\input_register_pci_ad_reg_out_reg[16]  <= n16410;
    \\input_register_pci_ad_reg_out_reg[28]  <= n16415;
    \\input_register_pci_ad_reg_out_reg[0]  <= n16420;
    \\configuration_int_pin_sync_sync_data_out_reg[0]  <= n16425;
    \\input_register_pci_ad_reg_out_reg[24]  <= n16430;
    \\input_register_pci_ad_reg_out_reg[10]  <= n16435;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[6]  <= n16440;
    \\input_register_pci_ad_reg_out_reg[12]  <= n16445;
    \\input_register_pci_ad_reg_out_reg[3]  <= n16450;
    \\input_register_pci_ad_reg_out_reg[13]  <= n16455;
    parity_checker_master_perr_report_reg <= n16460;
    \\input_register_pci_ad_reg_out_reg[4]  <= n16465;
    \\input_register_pci_ad_reg_out_reg[9]  <= n16470;
    \\input_register_pci_ad_reg_out_reg[14]  <= n16475;
    pci_target_unit_del_sync_comp_done_reg_clr_reg <= n16480;
    configuration_wb_init_complete_out_reg <= n16485;
    \\input_register_pci_ad_reg_out_reg[29]  <= n16490;
    \\input_register_pci_ad_reg_out_reg[25]  <= n16495;
    parity_checker_frame_dec2_reg <= n16500;
    \\input_register_pci_ad_reg_out_reg[15]  <= n16505;
    \\input_register_pci_ad_reg_out_reg[23]  <= n16510;
    \\input_register_pci_ad_reg_out_reg[20]  <= n16515;
    wishbone_slave_unit_del_sync_req_rty_exp_clr_reg <= n16520;
    \\input_register_pci_ad_reg_out_reg[26]  <= n16525;
    \\input_register_pci_ad_reg_out_reg[31]  <= n16530;
    \\input_register_pci_ad_reg_out_reg[6]  <= n16535;
    configuration_init_complete_reg <= n16540;
    input_register_pci_idsel_reg_out_reg <= n16545;
    \\input_register_pci_ad_reg_out_reg[21]  <= n16550;
    \\input_register_pci_ad_reg_out_reg[1]  <= n16555;
    \\input_register_pci_ad_reg_out_reg[18]  <= n16560;
    \\input_register_pci_ad_reg_out_reg[22]  <= n16565;
    \\input_register_pci_ad_reg_out_reg[2]  <= n16570;
    pci_target_unit_pci_target_sm_read_completed_reg_reg <= n16575;
    \\input_register_pci_ad_reg_out_reg[11]  <= n16580;
    \\input_register_pci_ad_reg_out_reg[5]  <= n16585;
    \\input_register_pci_ad_reg_out_reg[8]  <= n16590;
    \\input_register_pci_ad_reg_out_reg[19]  <= n16595;
    \\input_register_pci_ad_reg_out_reg[27]  <= n16600;
    parity_checker_frame_and_irdy_en_prev_prev_reg <= n16605;
    wishbone_slave_unit_del_sync_comp_done_reg_main_reg <= n16610;
    pci_target_unit_del_sync_comp_rty_exp_clr_reg <= n16615;
    configuration_pci_err_cs_bit8_reg <= n16620;
    \\configuration_isr_bit2_0_reg[2]  <= n16625;
    \\configuration_isr_bit2_0_reg[0]  <= n16630;
    wishbone_slave_unit_pci_initiator_if_write_req_int_reg <= n16635;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[0]  <= n16640;
    \\configuration_i_wb_init_complete_sync_sync_data_out_reg[0]  <= n16645;
    configuration_sync_isr_2_sync_del_bit_reg <= n16650;
    pci_io_mux_req_iob_en_out_reg <= n16655;
    pci_target_unit_del_sync_req_rty_exp_reg_reg <= n16660;
    configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg <= n16665;
    configuration_sync_isr_2_delayed_bckp_bit_reg <= n16670;
    wishbone_slave_unit_del_sync_req_comp_pending_sample_reg <= n16675;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[3]  <= n16680;
    pci_target_unit_del_sync_req_comp_pending_sample_reg <= n16685;
    \\pci_target_unit_del_sync_req_sync_sync_data_out_reg[0]  <= n16690;
    pci_target_unit_del_sync_comp_done_reg_main_reg <= n16695;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2]  <= n16700;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[0]  <= n16705;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0]  <= n16710;
    pci_io_mux_irdy_iob_en_out_reg <= n16715;
    \\pci_target_unit_del_sync_rty_exp_back_prop_sync_sync_data_out_reg[0]  <= n16720;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[0]  <= n16725;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1]  <= n16730;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]  <= n16735;
    \\wishbone_slave_unit_del_sync_req_sync_sync_data_out_reg[0]  <= n16740;
    wishbone_slave_unit_pci_initiator_sm_mabort2_reg <= n16745;
    \\wishbone_slave_unit_del_sync_done_sync_sync_data_out_reg[0]  <= n16750;
    pci_target_unit_del_sync_comp_flush_out_reg <= n16755;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[2]  <= n16760;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]  <= n16765;
    wishbone_slave_unit_del_sync_comp_flush_out_reg <= n16770;
    pci_target_unit_pci_target_sm_bckp_trdy_reg_reg <= n16775;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]  <= n16780;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3]  <= n16785;
    configuration_sync_pci_err_cs_8_sync_del_bit_reg <= n16790;
    parity_checker_frame_and_irdy_en_prev_reg <= n16795;
    \\configuration_isr_bit0_sync_sync_data_out_reg[0]  <= n16800;
    \\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[2]  <= n16805;
    \\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[1]  <= n16810;
    \\configuration_pci_err_cs_bits_sync_sync_data_out_reg[0]  <= n16815;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[3]  <= n16820;
    \\pci_target_unit_fifos_wb_clk_inGreyCount_reg[0]  <= n16825;
    \\pci_target_unit_fifos_wb_clk_inGreyCount_reg[1]  <= n16830;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[2]  <= n16835;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[1]  <= n16840;
    \\configuration_isr_bit2_sync_sync_data_out_reg[0]  <= n16845;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[1]  <= n16850;
    \\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[0]  <= n16855;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[0]  <= n16860;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]  <= n16865;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[0]  <= n16870;
    output_backup_irdy_en_out_reg <= n16875;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[3]  <= n16880;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1]  <= n16885;
    \\wishbone_slave_unit_del_sync_comp_sync_sync_data_out_reg[0]  <= n16890;
    \\pci_target_unit_del_sync_comp_sync_sync_data_out_reg[0]  <= n16895;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[1]  <= n16900;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[1]  <= n16905;
    \\pci_target_unit_del_sync_rty_exp_sync_sync_data_out_reg[0]  <= n16910;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]  <= n16915;
    \\configuration_sync_isr_2_delete_sync_sync_data_out_reg[0]  <= n16920;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[2]  <= n16925;
    \\pci_target_unit_del_sync_done_sync_sync_data_out_reg[0]  <= n16930;
    pci_target_unit_del_sync_req_rty_exp_clr_reg <= n16935;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[2]  <= n16940;
    configuration_rst_inactive_reg <= n16945;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[2]  <= n16950;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[4]  <= n16955;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[7]  <= n16960;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[5]  <= n16965;
    configuration_sync_command_bit_reg <= n16970;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[6]  <= n16975;
    configuration_sync_isr_2_sync_bckp_bit_reg <= n16980;
    wishbone_slave_unit_del_sync_req_rty_exp_reg_reg <= n16985;
    configuration_sync_pci_err_cs_8_sync_bckp_bit_reg <= n16990;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[1]  <= n16995;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg[1]  <= n17000;
    \\wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[2]  <= n17005;
    pci_target_unit_wishbone_master_burst_chopped_delayed_reg <= n17010;
    \\wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[1]  <= n17015;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[2]  <= n17020;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[1]  <= n17025;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg[2]  <= n17030;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[1]  <= n17035;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[3]  <= n17040;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[3]  <= n17045;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[1]  <= n17050;
    \\pci_target_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[1]  <= n17055;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg[0]  <= n17060;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[0]  <= n17065;
    \\pci_target_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[0]  <= n17070;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[2]  <= n17075;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[2]  <= n17080;
    \\configuration_sync_pci_err_cs_8_delete_sync_sync_data_out_reg[0]  <= n17085;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[0]  <= n17090;
    \\wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[0]  <= n17095;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[18]  <= n17100;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[31]  <= n17105;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[3]  <= n17110;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[4]  <= n17115;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[25]  <= n17120;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[6]  <= n17125;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[16]  <= n17130;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[11]  <= n17135;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[2]  <= n17140;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[1]  <= n17145;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[15]  <= n17150;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[14]  <= n17155;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg[0]  <= n17160;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[2]  <= n17165;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[13]  <= n17170;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[11]  <= n17175;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[10]  <= n17180;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg[2]  <= n17185;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[15]  <= n17190;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[8]  <= n17195;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[0]  <= n17200;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[6]  <= n17205;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[21]  <= n17210;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[25]  <= n17215;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[0]  <= n17220;
    \\configuration_sync_isr_2_clear_delete_sync_sync_data_out_reg[0]  <= n17225;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[19]  <= n17230;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[30]  <= n17235;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[27]  <= n17240;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[29]  <= n17245;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[3]  <= n17250;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[19]  <= n17255;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[23]  <= n17260;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[22]  <= n17265;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[28]  <= n17270;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[24]  <= n17275;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[4]  <= n17280;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[2]  <= n17285;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[5]  <= n17290;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[4]  <= n17295;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[13]  <= n17300;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[8]  <= n17305;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[16]  <= n17310;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[17]  <= n17315;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[1]  <= n17320;
    configuration_rst_inactive_sync_reg <= n17325;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[26]  <= n17330;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[5]  <= n17335;
    configuration_sync_isr_2_delayed_del_bit_reg <= n17340;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[22]  <= n17345;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[2]  <= n17350;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[1]  <= n17355;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg[1]  <= n17360;
    \\wishbone_slave_unit_del_sync_rty_exp_sync_sync_data_out_reg[0]  <= n17365;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[23]  <= n17370;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[20]  <= n17375;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[12]  <= n17380;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[12]  <= n17385;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[21]  <= n17390;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[0]  <= n17395;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[7]  <= n17400;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[20]  <= n17405;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[26]  <= n17410;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[9]  <= n17415;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[24]  <= n17420;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[7]  <= n17425;
    \\configuration_command_bit_sync_sync_data_out_reg[0]  <= n17430;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[0]  <= n17435;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[14]  <= n17440;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[31]  <= n17445;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[1]  <= n17450;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[0]  <= n17455;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[10]  <= n17460;
    \\configuration_sync_pci_err_cs_8_clear_delete_sync_sync_data_out_reg[0]  <= n17465;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[3]  <= n17470;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[18]  <= n17475;
    wishbone_slave_unit_del_sync_comp_done_reg_clr_reg <= n17480;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[27]  <= n17485;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[28]  <= n17490;
    configuration_sync_pci_err_cs_8_delayed_del_bit_reg <= n17495;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[3]  <= n17500;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[5]  <= n17505;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[29]  <= n17510;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[2]  <= n17515;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[17]  <= n17520;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[9]  <= n17525;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[30]  <= n17530;
  end
  initial begin
    \\pci_target_unit_wishbone_master_wb_cti_o_reg[0]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_cti_o_reg[2]  <= 1'b0;
    configuration_status_bit8_reg <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_sel_o_reg[0]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_sel_o_reg[1]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_sel_o_reg[2]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_sel_o_reg[3]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[0]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[10]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[11]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[12]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[13]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[16]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[17]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[19]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[1]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[20]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[21]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[22]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[23]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[24]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[25]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[26]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[27]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[28]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[29]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[2]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[31]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[3]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[4]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[5]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[6]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[8]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[9]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[30]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[14]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[18]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[7]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_dat_o_reg[15]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[19]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[22]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[24]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[20]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[27]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[21]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[30]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[25]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[28]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[31]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[29]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[17]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[10]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[11]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[12]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[16]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[14]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[13]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[23]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[26]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[3]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[4]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[5]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[6]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[8]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[9]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[2]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[18]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[15]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[7]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[0]  <= 1'b0;
    \\pci_target_unit_wishbone_master_addr_cnt_out_reg[1]  <= 1'b0;
    parity_checker_perr_sampled_reg <= 1'b0;
    \\pci_target_unit_wishbone_master_bc_register_reg[0]  <= 1'b0;
    \\pci_target_unit_wishbone_master_bc_register_reg[1]  <= 1'b0;
    \\pci_target_unit_wishbone_master_bc_register_reg[2]  <= 1'b0;
    \\pci_target_unit_wishbone_master_bc_register_reg[3]  <= 1'b0;
    pci_target_unit_wishbone_master_burst_chopped_reg <= 1'b0;
    pci_target_unit_pci_target_sm_backoff_reg <= 1'b0;
    wishbone_slave_unit_del_sync_req_done_reg_reg <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_c_state_reg[0]  <= 1'b0;
    \\pci_target_unit_wishbone_master_wb_cti_o_reg[1]  <= 1'b1;
    wishbone_slave_unit_del_sync_req_comp_pending_reg <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_c_state_reg[2]  <= 1'b0;
    output_backup_trdy_out_reg <= 1'b1;
    pci_io_mux_trdy_iob_dat_out_reg <= 1'b0;
    pci_io_mux_stop_iob_dat_out_reg <= 1'b0;
    output_backup_stop_out_reg <= 1'b1;
    pci_io_mux_devsel_iob_dat_out_reg <= 1'b0;
    output_backup_devsel_out_reg <= 1'b1;
    output_backup_perr_en_out_reg <= 1'b0;
    \\output_backup_ad_out_reg[31]  <= 1'b0;
    pci_io_mux_ad_iob31_dat_out_reg <= 1'b0;
    pci_io_mux_perr_iob_en_out_reg <= 1'b1;
    \\configuration_status_bit15_11_reg[15]  <= 1'b0;
    wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg <= 1'b0;
    \\output_backup_cbe_out_reg[0]  <= 1'b1;
    \\output_backup_cbe_out_reg[3]  <= 1'b1;
    pci_io_mux_cbe_iob0_dat_out_reg <= 1'b0;
    pci_io_mux_cbe_iob2_dat_out_reg <= 1'b0;
    \\output_backup_cbe_out_reg[2]  <= 1'b1;
    pci_io_mux_cbe_iob3_dat_out_reg <= 1'b0;
    \\output_backup_ad_out_reg[15]  <= 1'b0;
    \\output_backup_ad_out_reg[23]  <= 1'b0;
    \\output_backup_ad_out_reg[24]  <= 1'b0;
    \\output_backup_ad_out_reg[27]  <= 1'b0;
    \\output_backup_ad_out_reg[28]  <= 1'b0;
    \\output_backup_ad_out_reg[29]  <= 1'b0;
    \\output_backup_ad_out_reg[2]  <= 1'b0;
    \\output_backup_ad_out_reg[3]  <= 1'b0;
    \\output_backup_ad_out_reg[4]  <= 1'b0;
    \\output_backup_ad_out_reg[5]  <= 1'b0;
    \\output_backup_ad_out_reg[6]  <= 1'b0;
    \\output_backup_ad_out_reg[7]  <= 1'b0;
    \\output_backup_ad_out_reg[8]  <= 1'b0;
    pci_io_mux_ad_iob11_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob12_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob13_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob14_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob15_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob24_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob27_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob29_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob28_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob2_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob4_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob5_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob6_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob7_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob23_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob8_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob3_dat_out_reg <= 1'b0;
    \\output_backup_ad_out_reg[13]  <= 1'b0;
    \\output_backup_ad_out_reg[14]  <= 1'b0;
    \\output_backup_ad_out_reg[16]  <= 1'b0;
    \\output_backup_ad_out_reg[17]  <= 1'b0;
    \\output_backup_ad_out_reg[18]  <= 1'b0;
    \\output_backup_ad_out_reg[19]  <= 1'b0;
    \\output_backup_ad_out_reg[20]  <= 1'b0;
    \\output_backup_ad_out_reg[22]  <= 1'b0;
    \\output_backup_ad_out_reg[9]  <= 1'b0;
    pci_io_mux_ad_iob10_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob16_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob17_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob18_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob19_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob22_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob20_dat_out_reg <= 1'b0;
    \\output_backup_ad_out_reg[10]  <= 1'b0;
    pci_io_mux_ad_iob9_dat_out_reg <= 1'b0;
    \\output_backup_ad_out_reg[11]  <= 1'b0;
    \\output_backup_ad_out_reg[12]  <= 1'b0;
    \\output_backup_ad_out_reg[1]  <= 1'b0;
    \\output_backup_ad_out_reg[30]  <= 1'b0;
    pci_io_mux_ad_iob1_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob30_dat_out_reg <= 1'b0;
    \\output_backup_ad_out_reg[21]  <= 1'b0;
    pci_io_mux_ad_iob21_dat_out_reg <= 1'b0;
    \\configuration_status_bit15_11_reg[14]  <= 1'b0;
    \\output_backup_ad_out_reg[26]  <= 1'b0;
    pci_io_mux_ad_iob26_dat_out_reg <= 1'b0;
    pci_io_mux_ad_iob0_dat_out_reg <= 1'b0;
    \\output_backup_ad_out_reg[0]  <= 1'b0;
    parity_checker_perr_en_crit_gen_perr_en_reg_out_reg <= 1'b0;
    \\output_backup_ad_out_reg[25]  <= 1'b0;
    pci_io_mux_ad_iob25_dat_out_reg <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_be_out_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_pci_initiator_if_be_out_reg[2]  <= 1'b1;
    \\wishbone_slave_unit_pci_initiator_if_be_out_reg[3]  <= 1'b1;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[10]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[11]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[16]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[18]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[19]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[1]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[21]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[22]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[30]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[5]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[6]  <= 1'b0;
    pci_io_mux_perr_iob_dat_out_reg <= 1'b0;
    pci_io_mux_serr_iob_en_out_reg <= 1'b1;
    pci_io_mux_serr_iob_dat_out_reg <= 1'b0;
    pci_target_unit_wishbone_master_first_wb_data_access_reg <= 1'b1;
    output_backup_perr_out_reg <= 1'b1;
    output_backup_serr_out_reg <= 1'b1;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[15]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[24]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[25]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[27]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[2]  <= 1'b0;
    output_backup_serr_en_out_reg <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[0]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[12]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[13]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[14]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[17]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[20]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[23]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[26]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[28]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[29]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[31]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[3]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[4]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[7]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[8]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg[9]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[24]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[12]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[14]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[17]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[18]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[20]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[21]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[22]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[25]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[26]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[27]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[29]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[4]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[5]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[7]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[26]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_outTransactionCount_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_outGreyCount_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[19]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[23]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[28]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[16]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[10]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[11]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[12]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[13]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[14]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[15]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[17]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[18]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[19]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[20]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[22]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[24]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[27]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[28]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[29]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[31]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[4]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[6]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[7]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[8]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[11]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[13]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[15]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[6]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[8]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[10]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[2]  <= 1'b1;
    \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_outTransactionCount_reg[0]  <= 1'b1;
    \\pci_target_unit_fifos_outGreyCount_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg[2]  <= 1'b1;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[0]  <= 1'b1;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[1]  <= 1'b1;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg[0]  <= 1'b1;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[1]  <= 1'b1;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_dword_address_reg[9]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_current_byte_address_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[5]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[9]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[23]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[16]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[21]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[25]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[0]  <= 1'b0;
    pci_target_unit_wishbone_master_wb_we_o_reg <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg[2]  <= 1'b1;
    pci_target_unit_wishbone_master_wb_cyc_o_reg <= 1'b0;
    pci_target_unit_wishbone_master_wb_stb_o_reg <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_data_reg[30]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_reg[1]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[15]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[25]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[7]  <= 1'b0;
    parity_checker_check_perr_reg <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[0]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[10]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[11]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[13]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[14]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[17]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[18]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[19]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[21]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[22]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[20]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[24]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[26]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[28]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[29]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[2]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[31]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[3]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[4]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[6]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[8]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[9]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[5]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[30]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[27]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[23]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[12]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[1]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg[16]  <= 1'b0;
    output_backup_par_en_out_reg <= 1'b0;
    pci_io_mux_par_iob_en_out_reg <= 1'b1;
    \\pci_target_unit_wishbone_master_c_state_reg[0]  <= 1'b0;
    i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg <= 1'b0;
    pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[11]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[10]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[13]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[14]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[15]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[16]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[17]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[19]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[20]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[21]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[23]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[24]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[25]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[27]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[12]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[29]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[30]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[31]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[3]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[5]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[6]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[7]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[9]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[28]  <= 1'b0;
    i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[22]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[18]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[8]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[26]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[4]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[2]  <= 1'b0;
    pci_io_mux_ad_iob23_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob22_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob21_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob19_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob17_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob18_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob15_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob14_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob13_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob11_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob25_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob8_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob7_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob9_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob5_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob3_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob4_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob1_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob2_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob26_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob31_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob29_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob28_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob27_en_out_reg <= 1'b1;
    output_backup_mas_ad_en_out_reg <= 1'b0;
    output_backup_tar_ad_en_out_reg <= 1'b0;
    pci_io_mux_ad_iob30_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob0_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob6_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob12_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob10_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob16_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob20_en_out_reg <= 1'b1;
    pci_io_mux_ad_iob24_en_out_reg <= 1'b1;
    pci_target_unit_wishbone_master_first_data_is_burst_reg_reg <= 1'b0;
    i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[10]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[11]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[13]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[15]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[16]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[17]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[19]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[20]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[23]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[24]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[26]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[27]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[28]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[30]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[31]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[7]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[8]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[9]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[1]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_del_sync_addr_out_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[29]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[18]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[21]  <= 1'b0;
    \\pci_target_unit_pci_target_sm_c_state_reg[0]  <= 1'b1;
    \\pci_target_unit_pci_target_sm_c_state_reg[1]  <= 1'b0;
    \\pci_target_unit_pci_target_sm_c_state_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[1]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[1]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg[3]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[12]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[22]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[5]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[4]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[25]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[6]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_addr_out_reg[14]  <= 1'b0;
    \\wishbone_slave_unit_fifos_inGreyCount_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_inGreyCount_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_fifos_inGreyCount_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_inTransactionCount_reg[0]  <= 1'b1;
    i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[1]  <= 1'b1;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[0]  <= 1'b1;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[1]  <= 1'b0;
    wishbone_slave_unit_del_sync_burst_out_reg <= 1'b0;
    pci_target_unit_wishbone_master_addr_into_cnt_reg_reg <= 1'b0;
    output_backup_trdy_en_out_reg <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg[1]  <= 1'b1;
    pci_io_mux_trdy_iob_en_out_reg <= 1'b1;
    pci_io_mux_stop_iob_en_out_reg <= 1'b1;
    pci_io_mux_devsel_iob_en_out_reg <= 1'b1;
    \\pci_target_unit_wishbone_master_rty_counter_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_bc_out_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[0]  <= 1'b1;
    output_backup_frame_out_reg <= 1'b1;
    \\pci_target_unit_wishbone_master_rty_counter_reg[5]  <= 1'b0;
    \\pci_target_unit_wishbone_master_rty_counter_reg[6]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_bc_out_reg[2]  <= 1'b1;
    \\pci_target_unit_wishbone_master_rty_counter_reg[1]  <= 1'b0;
    \\pci_target_unit_wishbone_master_rty_counter_reg[2]  <= 1'b0;
    \\pci_target_unit_wishbone_master_rty_counter_reg[4]  <= 1'b0;
    \\wishbone_slave_unit_fifos_outGreyCount_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[2]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg[1]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[3]  <= 1'b0;
    \\pci_target_unit_wishbone_master_rty_counter_reg[3]  <= 1'b0;
    \\pci_target_unit_wishbone_master_rty_counter_reg[7]  <= 1'b0;
    pci_io_mux_frame_iob_dat_out_reg <= 1'b0;
    pci_target_unit_pci_target_sm_rd_request_reg <= 1'b0;
    pci_target_unit_pci_target_sm_rd_progress_reg <= 1'b0;
    \\wishbone_slave_unit_del_sync_be_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_be_out_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_be_out_reg[2]  <= 1'b0;
    wishbone_slave_unit_del_sync_we_out_reg <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg[1]  <= 1'b1;
    \\wishbone_slave_unit_del_sync_be_out_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_bc_out_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[12]  <= 1'b0;
    pci_target_unit_pci_target_if_norm_prf_en_reg <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[10]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[11]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[13]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[14]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[15]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[17]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[18]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[21]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[23]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[25]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[26]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[27]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[29]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[30]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[32]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[33]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[34]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[5]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[8]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[7]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[10]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[11]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[14]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[5]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[9]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[7]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[0]  <= 1'b1;
    pci_target_unit_pci_target_if_pciw_fifo_wenable_out_reg <= 1'b0;
    \\wishbone_slave_unit_fifos_outGreyCount_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[6]  <= 1'b0;
    \\wishbone_slave_unit_fifos_outGreyCount_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_bc_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_outTransactionCount_reg[2]  <= 1'b0;
    i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[6]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[4]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[13]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[15]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[16]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[9]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[4]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[35]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[31]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[22]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[28]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[24]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[16]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[20]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[12]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_d_incoming_reg[19]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_comp_cycle_count_reg[8]  <= 1'b0;
    pci_target_unit_pci_target_sm_wr_progress_reg <= 1'b0;
    pci_target_unit_wishbone_master_w_attempt_reg <= 1'b0;
    \\configuration_wb_am2_reg[31]  <= 1'b1;
    \\configuration_wb_am1_reg[31]  <= 1'b1;
    pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg <= 1'b0;
    \\output_backup_cbe_out_reg[1]  <= 1'b1;
    wishbone_slave_unit_pci_initiator_if_del_read_req_reg <= 1'b0;
    \\configuration_pci_img_ctrl1_bit2_1_reg[1]  <= 1'b0;
    \\configuration_pci_img_ctrl1_bit2_1_reg[2]  <= 1'b0;
    \\configuration_wb_ta1_reg[31]  <= 1'b0;
    configuration_wb_err_cs_bit0_reg <= 1'b0;
    \\configuration_wb_ta2_reg[31]  <= 1'b0;
    pci_io_mux_cbe_iob1_dat_out_reg <= 1'b0;
    pci_target_unit_pci_target_sm_master_will_request_read_reg <= 1'b0;
    wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg <= 1'b1;
    output_backup_par_out_reg <= 1'b0;
    pci_io_mux_par_iob_dat_out_reg <= 1'b0;
    configuration_pci_err_cs_bit0_reg <= 1'b0;
    \\configuration_wb_img_ctrl1_bit2_0_reg[2]  <= 1'b0;
    \\configuration_interrupt_line_reg[6]  <= 1'b0;
    \\configuration_wb_img_ctrl2_bit2_0_reg[1]  <= 1'b0;
    \\configuration_interrupt_line_reg[2]  <= 1'b0;
    wishbone_slave_unit_del_sync_req_req_pending_reg <= 1'b0;
    \\configuration_wb_img_ctrl1_bit2_0_reg[0]  <= 1'b0;
    \\configuration_wb_img_ctrl1_bit2_0_reg[1]  <= 1'b0;
    \\configuration_interrupt_line_reg[0]  <= 1'b0;
    \\configuration_interrupt_line_reg[1]  <= 1'b0;
    \\configuration_wb_img_ctrl2_bit2_0_reg[0]  <= 1'b0;
    \\configuration_wb_img_ctrl2_bit2_0_reg[2]  <= 1'b0;
    \\configuration_command_bit2_0_reg[0]  <= 1'b0;
    \\configuration_command_bit2_0_reg[1]  <= 1'b0;
    \\configuration_command_bit2_0_reg[2]  <= 1'b0;
    configuration_wb_ba1_bit0_reg <= 1'b0;
    configuration_wb_ba2_bit0_reg <= 1'b0;
    configuration_command_bit8_reg <= 1'b0;
    configuration_wb_err_cs_bit8_reg <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[1]  <= 1'b1;
    \\configuration_status_bit15_11_reg[11]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[1]  <= 1'b0;
    \\configuration_status_bit15_11_reg[12]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[0]  <= 1'b0;
    \\configuration_status_bit15_11_reg[13]  <= 1'b0;
    \\configuration_isr_bit2_0_reg[1]  <= 1'b0;
    wishbone_slave_unit_del_sync_comp_comp_pending_reg <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[0]  <= 1'b1;
    pci_target_unit_wishbone_master_reset_rty_cnt_reg <= 1'b1;
    \\configuration_wb_ba2_bit31_12_reg[31]  <= 1'b1;
    \\configuration_wb_ba1_bit31_12_reg[31]  <= 1'b0;
    configuration_command_bit6_reg <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[1]  <= 1'b0;
    \\configuration_icr_bit2_0_reg[0]  <= 1'b0;
    \\configuration_icr_bit2_0_reg[1]  <= 1'b0;
    \\configuration_icr_bit2_0_reg[2]  <= 1'b0;
    \\configuration_interrupt_line_reg[3]  <= 1'b0;
    \\configuration_cache_line_size_reg_reg[3]  <= 1'b0;
    \\configuration_interrupt_line_reg[5]  <= 1'b0;
    \\configuration_interrupt_line_reg[4]  <= 1'b0;
    \\configuration_cache_line_size_reg_reg[5]  <= 1'b0;
    \\configuration_cache_line_size_reg_reg[4]  <= 1'b0;
    configuration_sync_isr_2_del_bit_reg <= 1'b0;
    configuration_sync_pci_err_cs_8_del_bit_reg <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg[2]  <= 1'b0;
    \\configuration_cache_line_size_reg_reg[7]  <= 1'b0;
    \\configuration_interrupt_line_reg[7]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[5]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[7]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[8]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[23]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[4]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[31]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[12]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[27]  <= 1'b0;
    \\configuration_latency_timer_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[12]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[21]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[14]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[16]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[1]  <= 1'b0;
    configuration_icr_bit31_reg <= 1'b0;
    wishbone_slave_unit_wishbone_slave_img_wallow_reg <= 1'b0;
    wishbone_slave_unit_wishbone_slave_do_del_request_reg <= 1'b0;
    wishbone_slave_unit_wishbone_slave_mrl_en_reg <= 1'b0;
    wishbone_slave_unit_wishbone_slave_pref_en_reg <= 1'b0;
    wishbone_slave_unit_wishbone_slave_del_addr_hit_reg <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_bc_out_reg[1]  <= 1'b0;
    wishbone_slave_unit_wishbone_slave_del_completion_allow_reg <= 1'b0;
    pci_target_unit_del_sync_comp_comp_pending_reg <= 1'b0;
    pci_target_unit_del_sync_comp_req_pending_reg <= 1'b0;
    \\pci_target_unit_wishbone_master_c_state_reg[2]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_if_intermediate_last_reg <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_intermediate_be_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_cur_state_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg[0]  <= 1'b1;
    \\configuration_latency_timer_reg[0]  <= 1'b0;
    \\configuration_latency_timer_reg[2]  <= 1'b0;
    \\configuration_latency_timer_reg[3]  <= 1'b0;
    \\configuration_latency_timer_reg[4]  <= 1'b0;
    \\configuration_latency_timer_reg[5]  <= 1'b0;
    \\configuration_latency_timer_reg[6]  <= 1'b0;
    \\configuration_latency_timer_reg[7]  <= 1'b0;
    \\configuration_cache_line_size_reg_reg[0]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[14]  <= 1'b0;
    \\configuration_cache_line_size_reg_reg[1]  <= 1'b0;
    \\configuration_cache_line_size_reg_reg[2]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[13]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[17]  <= 1'b0;
    \\configuration_cache_line_size_reg_reg[6]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[16]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[20]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[23]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[18]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[15]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[19]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[25]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[27]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[28]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[30]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[29]  <= 1'b0;
    \\pci_target_unit_wishbone_master_read_count_reg[1]  <= 1'b0;
    \\pci_target_unit_wishbone_master_read_count_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[10]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[11]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[13]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[15]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[17]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[18]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[19]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[20]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[22]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[24]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[25]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[26]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[28]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[29]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[6]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[9]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_data_out_reg[30]  <= 1'b0;
    wishbone_slave_unit_del_sync_comp_req_pending_reg <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[31]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[26]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[24]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[21]  <= 1'b0;
    \\configuration_pci_ba0_bit31_8_reg[22]  <= 1'b0;
    \\configuration_pci_am1_reg[16]  <= 1'b1;
    \\configuration_pci_am1_reg[15]  <= 1'b1;
    \\configuration_pci_am1_reg[24]  <= 1'b1;
    \\configuration_pci_ba1_bit31_8_reg[11]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[15]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_read_count_reg[3]  <= 1'b0;
    wishbone_slave_unit_wishbone_slave_map_reg <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[18]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[19]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[20]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[21]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[23]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[25]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[26]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[27]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[29]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[30]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[10]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[12]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[13]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[14]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[16]  <= 1'b0;
    \\pci_target_unit_wishbone_master_c_state_reg[1]  <= 1'b0;
    \\configuration_pci_am1_reg[21]  <= 1'b1;
    \\configuration_pci_am1_reg[10]  <= 1'b1;
    \\configuration_pci_am1_reg[12]  <= 1'b1;
    \\configuration_pci_am1_reg[11]  <= 1'b1;
    \\configuration_pci_am1_reg[13]  <= 1'b1;
    \\configuration_pci_am1_reg[18]  <= 1'b1;
    \\configuration_pci_am1_reg[17]  <= 1'b1;
    \\configuration_pci_am1_reg[20]  <= 1'b1;
    \\configuration_pci_am1_reg[14]  <= 1'b1;
    \\configuration_pci_am1_reg[22]  <= 1'b1;
    \\configuration_pci_am1_reg[23]  <= 1'b1;
    \\configuration_pci_am1_reg[25]  <= 1'b1;
    \\configuration_pci_am1_reg[19]  <= 1'b1;
    \\configuration_pci_am1_reg[29]  <= 1'b1;
    \\configuration_pci_am1_reg[31]  <= 1'b1;
    \\configuration_pci_am1_reg[30]  <= 1'b1;
    \\configuration_pci_am1_reg[28]  <= 1'b1;
    \\pci_target_unit_wishbone_master_read_count_reg[0]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[31]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[1]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[8]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[9]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[22]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[28]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[24]  <= 1'b0;
    \\configuration_pci_ba1_bit31_8_reg[17]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_if_current_last_reg <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[0]  <= 1'b0;
    \\configuration_pci_am1_reg[26]  <= 1'b1;
    \\configuration_pci_am1_reg[8]  <= 1'b1;
    \\configuration_pci_am1_reg[9]  <= 1'b1;
    \\configuration_pci_am1_reg[27]  <= 1'b1;
    \\wishbone_slave_unit_wishbone_slave_c_state_reg[1]  <= 1'b0;
    \\configuration_pci_ta1_reg[10]  <= 1'b0;
    pci_target_unit_wishbone_master_read_bound_reg <= 1'b0;
    \\configuration_pci_ta1_reg[29]  <= 1'b0;
    \\configuration_pci_ta1_reg[16]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_read_count_reg[2]  <= 1'b0;
    \\configuration_pci_ta1_reg[17]  <= 1'b0;
    \\configuration_pci_ta1_reg[18]  <= 1'b0;
    \\configuration_pci_ta1_reg[20]  <= 1'b0;
    \\configuration_pci_ta1_reg[21]  <= 1'b0;
    \\configuration_pci_ta1_reg[24]  <= 1'b0;
    \\configuration_pci_ta1_reg[23]  <= 1'b0;
    \\configuration_pci_ta1_reg[30]  <= 1'b0;
    \\configuration_pci_ta1_reg[28]  <= 1'b0;
    \\configuration_pci_ta1_reg[31]  <= 1'b0;
    \\configuration_pci_ta1_reg[14]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_if_err_recovery_reg <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[1]  <= 1'b0;
    \\configuration_pci_ta1_reg[11]  <= 1'b0;
    \\configuration_pci_ta1_reg[13]  <= 1'b0;
    \\configuration_pci_ta1_reg[15]  <= 1'b0;
    \\configuration_pci_ta1_reg[12]  <= 1'b0;
    \\configuration_pci_ta1_reg[8]  <= 1'b0;
    \\configuration_pci_ta1_reg[9]  <= 1'b0;
    \\configuration_pci_ta1_reg[27]  <= 1'b0;
    \\configuration_pci_ta1_reg[26]  <= 1'b0;
    \\configuration_pci_ta1_reg[25]  <= 1'b0;
    \\configuration_pci_ta1_reg[22]  <= 1'b0;
    \\configuration_pci_ta1_reg[19]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_if_posted_write_req_reg <= 1'b0;
    pci_io_mux_frame_iob_en_out_reg <= 1'b1;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[27]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[17]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[19]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[20]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[22]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[23]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[24]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[28]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[29]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[2]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[31]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[3]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[4]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[6]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[8]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[16]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[14]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[0]  <= 1'b0;
    output_backup_cbe_en_out_reg <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[13]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[15]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[9]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[5]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[7]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[26]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[30]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[18]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[21]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[1]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[12]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[25]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[11]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[0]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg[10]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_be_out_reg[1]  <= 1'b1;
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[4]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[16]  <= 1'b0;
    configuration_set_isr_bit2_reg <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_wishbone_slave_img_hit_reg[3]  <= 1'b0;
    wishbone_slave_unit_wishbone_slave_wb_conf_hit_reg <= 1'b0;
    \\configuration_wb_err_addr_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[6]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[2]  <= 1'b0;
    output_backup_frame_en_out_reg <= 1'b0;
    pci_io_mux_cbe_iob3_en_out_reg <= 1'b1;
    pci_io_mux_cbe_iob2_en_out_reg <= 1'b1;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[3]  <= 1'b0;
    configuration_wb_err_cs_bit9_reg <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg[1]  <= 1'b0;
    pci_io_mux_cbe_iob1_en_out_reg <= 1'b1;
    pci_io_mux_cbe_iob0_en_out_reg <= 1'b1;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[5]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[1]  <= 1'b0;
    i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg <= 1'b0;
    \\configuration_wb_err_addr_reg[11]  <= 1'b0;
    \\configuration_wb_err_data_reg[0]  <= 1'b0;
    \\configuration_wb_err_cs_bit31_24_reg[30]  <= 1'b0;
    \\configuration_wb_err_addr_reg[19]  <= 1'b0;
    \\configuration_pci_err_data_reg[28]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_if_data_source_reg <= 1'b0;
    \\configuration_wb_err_cs_bit31_24_reg[28]  <= 1'b0;
    \\configuration_wb_err_addr_reg[15]  <= 1'b0;
    \\configuration_wb_err_data_reg[6]  <= 1'b0;
    \\configuration_wb_err_data_reg[8]  <= 1'b0;
    \\configuration_wb_err_data_reg[30]  <= 1'b0;
    \\configuration_wb_err_data_reg[4]  <= 1'b0;
    \\configuration_wb_err_data_reg[31]  <= 1'b0;
    \\configuration_wb_err_data_reg[28]  <= 1'b0;
    \\configuration_wb_err_data_reg[27]  <= 1'b0;
    \\configuration_wb_err_data_reg[24]  <= 1'b0;
    \\configuration_wb_err_data_reg[20]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_if_read_bound_reg <= 1'b0;
    configuration_pci_err_cs_bit9_reg <= 1'b0;
    configuration_pci_err_cs_bit10_reg <= 1'b0;
    \\configuration_pci_err_cs_bit31_24_reg[30]  <= 1'b0;
    \\configuration_pci_err_cs_bit31_24_reg[28]  <= 1'b0;
    \\configuration_pci_err_cs_bit31_24_reg[29]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_read_count_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[4]  <= 1'b0;
    \\configuration_pci_err_addr_reg[0]  <= 1'b0;
    \\configuration_pci_err_addr_reg[11]  <= 1'b0;
    \\configuration_pci_err_addr_reg[12]  <= 1'b0;
    \\configuration_pci_err_addr_reg[15]  <= 1'b0;
    \\configuration_pci_err_addr_reg[19]  <= 1'b0;
    \\configuration_pci_err_addr_reg[20]  <= 1'b0;
    \\configuration_pci_err_addr_reg[22]  <= 1'b0;
    \\configuration_pci_err_addr_reg[26]  <= 1'b0;
    \\configuration_pci_err_addr_reg[28]  <= 1'b0;
    \\configuration_pci_err_addr_reg[2]  <= 1'b0;
    \\configuration_pci_err_addr_reg[31]  <= 1'b0;
    \\configuration_pci_err_addr_reg[4]  <= 1'b0;
    \\configuration_pci_err_addr_reg[6]  <= 1'b0;
    \\configuration_pci_err_addr_reg[8]  <= 1'b0;
    \\configuration_pci_err_data_reg[0]  <= 1'b0;
    \\configuration_pci_err_data_reg[11]  <= 1'b0;
    \\configuration_pci_err_data_reg[13]  <= 1'b0;
    \\configuration_pci_err_data_reg[15]  <= 1'b0;
    \\configuration_pci_err_data_reg[17]  <= 1'b0;
    \\configuration_pci_err_data_reg[19]  <= 1'b0;
    \\configuration_pci_err_data_reg[21]  <= 1'b0;
    \\configuration_pci_err_data_reg[25]  <= 1'b0;
    \\configuration_pci_err_data_reg[29]  <= 1'b0;
    \\configuration_pci_err_data_reg[31]  <= 1'b0;
    \\configuration_pci_err_data_reg[3]  <= 1'b0;
    \\configuration_pci_err_data_reg[7]  <= 1'b0;
    pci_target_unit_pci_target_sm_same_read_reg_reg <= 1'b0;
    \\configuration_wb_err_cs_bit31_24_reg[25]  <= 1'b0;
    \\configuration_wb_err_cs_bit31_24_reg[31]  <= 1'b0;
    \\configuration_wb_err_data_reg[10]  <= 1'b0;
    \\configuration_wb_err_data_reg[11]  <= 1'b0;
    \\configuration_wb_err_data_reg[12]  <= 1'b0;
    \\configuration_wb_err_data_reg[14]  <= 1'b0;
    \\configuration_wb_err_data_reg[15]  <= 1'b0;
    \\configuration_wb_err_data_reg[16]  <= 1'b0;
    \\configuration_wb_err_data_reg[18]  <= 1'b0;
    \\configuration_wb_err_data_reg[19]  <= 1'b0;
    \\configuration_wb_err_data_reg[1]  <= 1'b0;
    \\configuration_wb_err_data_reg[21]  <= 1'b0;
    \\configuration_wb_err_data_reg[22]  <= 1'b0;
    \\configuration_wb_err_data_reg[23]  <= 1'b0;
    \\configuration_wb_err_data_reg[25]  <= 1'b0;
    \\configuration_wb_err_data_reg[26]  <= 1'b0;
    \\configuration_wb_err_data_reg[29]  <= 1'b0;
    \\configuration_wb_err_data_reg[2]  <= 1'b0;
    \\configuration_wb_err_data_reg[3]  <= 1'b0;
    \\configuration_wb_err_data_reg[5]  <= 1'b0;
    \\configuration_wb_err_data_reg[9]  <= 1'b0;
    \\configuration_wb_err_data_reg[7]  <= 1'b0;
    \\configuration_wb_err_addr_reg[10]  <= 1'b0;
    \\configuration_wb_err_addr_reg[12]  <= 1'b0;
    \\configuration_wb_err_addr_reg[13]  <= 1'b0;
    \\configuration_wb_err_addr_reg[14]  <= 1'b0;
    \\configuration_wb_err_addr_reg[16]  <= 1'b0;
    \\configuration_wb_err_addr_reg[18]  <= 1'b0;
    \\configuration_wb_err_addr_reg[20]  <= 1'b0;
    \\configuration_wb_err_addr_reg[22]  <= 1'b0;
    \\configuration_wb_err_addr_reg[24]  <= 1'b0;
    \\configuration_wb_err_addr_reg[26]  <= 1'b0;
    \\configuration_wb_err_addr_reg[28]  <= 1'b0;
    \\configuration_wb_err_addr_reg[2]  <= 1'b0;
    \\configuration_wb_err_addr_reg[31]  <= 1'b0;
    \\configuration_wb_err_addr_reg[4]  <= 1'b0;
    \\configuration_wb_err_addr_reg[6]  <= 1'b0;
    \\configuration_wb_err_addr_reg[7]  <= 1'b0;
    \\configuration_wb_err_addr_reg[8]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_inTransactionCount_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_inGreyCount_reg[0]  <= 1'b0;
    \\configuration_wb_err_cs_bit31_24_reg[29]  <= 1'b0;
    \\configuration_wb_err_data_reg[13]  <= 1'b0;
    \\configuration_wb_err_cs_bit31_24_reg[24]  <= 1'b0;
    \\configuration_wb_err_cs_bit31_24_reg[27]  <= 1'b0;
    \\configuration_wb_err_cs_bit31_24_reg[26]  <= 1'b0;
    \\configuration_wb_err_data_reg[17]  <= 1'b0;
    \\configuration_pci_err_data_reg[2]  <= 1'b0;
    \\configuration_wb_err_addr_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_latency_timer_reg[7]  <= 1'b0;
    pci_target_unit_pci_target_if_same_read_reg_reg <= 1'b0;
    \\configuration_pci_err_data_reg[8]  <= 1'b0;
    \\configuration_pci_err_data_reg[30]  <= 1'b0;
    \\configuration_pci_err_data_reg[9]  <= 1'b0;
    \\configuration_pci_err_data_reg[5]  <= 1'b0;
    \\configuration_pci_err_data_reg[6]  <= 1'b0;
    \\configuration_pci_err_data_reg[4]  <= 1'b0;
    \\configuration_pci_err_data_reg[23]  <= 1'b0;
    \\configuration_wb_err_addr_reg[17]  <= 1'b0;
    \\configuration_pci_err_data_reg[24]  <= 1'b0;
    \\configuration_pci_err_data_reg[26]  <= 1'b0;
    \\configuration_pci_err_data_reg[27]  <= 1'b0;
    \\configuration_pci_err_addr_reg[7]  <= 1'b0;
    \\configuration_pci_err_addr_reg[9]  <= 1'b0;
    \\configuration_pci_err_data_reg[18]  <= 1'b0;
    \\configuration_pci_err_data_reg[1]  <= 1'b0;
    \\configuration_pci_err_data_reg[20]  <= 1'b0;
    \\configuration_pci_err_data_reg[22]  <= 1'b0;
    \\configuration_pci_err_data_reg[14]  <= 1'b0;
    \\configuration_pci_err_cs_bit31_24_reg[24]  <= 1'b0;
    \\configuration_pci_err_data_reg[16]  <= 1'b0;
    \\configuration_pci_err_cs_bit31_24_reg[25]  <= 1'b0;
    \\configuration_pci_err_data_reg[10]  <= 1'b0;
    \\configuration_pci_err_data_reg[12]  <= 1'b0;
    \\configuration_pci_err_cs_bit31_24_reg[26]  <= 1'b0;
    \\configuration_pci_err_cs_bit31_24_reg[27]  <= 1'b0;
    \\configuration_pci_err_addr_reg[3]  <= 1'b0;
    \\configuration_pci_err_addr_reg[10]  <= 1'b0;
    \\configuration_wb_err_addr_reg[21]  <= 1'b0;
    \\configuration_pci_err_addr_reg[5]  <= 1'b0;
    \\configuration_pci_err_addr_reg[30]  <= 1'b0;
    \\configuration_pci_err_addr_reg[27]  <= 1'b0;
    \\configuration_pci_err_addr_reg[29]  <= 1'b0;
    \\configuration_pci_err_addr_reg[25]  <= 1'b0;
    \\configuration_pci_err_addr_reg[1]  <= 1'b0;
    \\configuration_pci_err_addr_reg[23]  <= 1'b0;
    \\configuration_pci_err_addr_reg[24]  <= 1'b0;
    \\configuration_pci_err_addr_reg[21]  <= 1'b0;
    \\configuration_pci_err_addr_reg[13]  <= 1'b0;
    \\configuration_pci_err_addr_reg[18]  <= 1'b0;
    \\configuration_pci_err_addr_reg[17]  <= 1'b0;
    \\configuration_pci_err_addr_reg[14]  <= 1'b0;
    \\configuration_pci_err_addr_reg[16]  <= 1'b0;
    \\configuration_pci_err_cs_bit31_24_reg[31]  <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_if_read_count_reg[0]  <= 1'b0;
    \\configuration_wb_err_addr_reg[9]  <= 1'b0;
    \\configuration_wb_err_addr_reg[5]  <= 1'b0;
    \\configuration_wb_err_addr_reg[3]  <= 1'b0;
    \\configuration_wb_err_addr_reg[23]  <= 1'b0;
    \\configuration_wb_err_addr_reg[30]  <= 1'b0;
    \\configuration_wb_err_addr_reg[29]  <= 1'b0;
    \\configuration_wb_err_addr_reg[25]  <= 1'b0;
    \\configuration_wb_err_addr_reg[27]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_inTransactionCount_reg[0]  <= 1'b1;
    \\pci_target_unit_fifos_inGreyCount_reg[1]  <= 1'b0;
    pci_target_unit_del_sync_comp_rty_exp_reg_reg <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[2]  <= 1'b1;
    configuration_set_pci_err_cs_bit8_reg <= 1'b0;
    wishbone_slave_unit_pci_initiator_if_del_write_req_reg <= 1'b0;
    pci_target_unit_wishbone_master_wb_read_done_out_reg <= 1'b0;
    pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[0]  <= 1'b1;
    pci_target_unit_del_sync_req_done_reg_reg <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[1]  <= 1'b0;
    \\pci_target_unit_pci_target_if_strd_address_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[1]  <= 1'b1;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[1]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_sm_timeout_reg <= 1'b0;
    \\wishbone_slave_unit_pci_initiator_sm_decode_count_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[0]  <= 1'b1;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[2]  <= 1'b0;
    pci_target_unit_pci_target_sm_wr_to_fifo_reg <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[0]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[15]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg[2]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[2]  <= 1'b1;
    pci_target_unit_del_sync_req_comp_pending_reg <= 1'b0;
    wishbone_slave_unit_pci_initiator_sm_transfer_reg <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg[1]  <= 1'b1;
    \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[1]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[14]  <= 1'b0;
    wishbone_slave_unit_del_sync_comp_rty_exp_reg_reg <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg[2]  <= 1'b1;
    parity_checker_check_for_serr_on_second_reg <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg[1]  <= 1'b1;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg[2]  <= 1'b1;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[1]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg[0]  <= 1'b1;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[12]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[1]  <= 1'b0;
    \\i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg[3]  <= 1'b0;
    i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg <= 1'b0;
    pci_target_unit_pci_target_if_target_rd_reg <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[11]  <= 1'b0;
    pci_target_unit_pci_target_sm_rd_from_fifo_reg <= 1'b0;
    pci_resets_and_interrupts_inta_en_out_reg <= 1'b1;
    \\pci_target_unit_pci_target_if_norm_bc_reg[0]  <= 1'b0;
    \\pci_target_unit_pci_target_if_strd_address_reg[3]  <= 1'b0;
    pci_target_unit_wishbone_master_retried_reg <= 1'b0;
    pci_target_unit_wishbone_master_pcir_fifo_wenable_out_reg <= 1'b0;
    pci_target_unit_pci_target_sm_rw_cbe0_reg <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[10]  <= 1'b0;
    \\pci_target_unit_del_sync_be_out_reg[0]  <= 1'b0;
    \\input_register_pci_cbe_reg_out_reg[0]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[8]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[13]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_if_last_transfered_reg <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[0]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[7]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[9]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[4]  <= 1'b0;
    \\pci_target_unit_pci_target_if_strd_address_reg[1]  <= 1'b0;
    \\pci_target_unit_pci_target_if_strd_address_reg[8]  <= 1'b0;
    \\pci_target_unit_pci_target_if_strd_address_reg[6]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[6]  <= 1'b0;
    pci_target_unit_pci_target_sm_cnf_progress_reg <= 1'b0;
    wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[3]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[0]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[1]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_if_rdy_out_reg <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[1]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[2]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[3]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_bc_reg[1]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_control_out_reg[1]  <= 1'b0;
    \\pci_target_unit_pci_target_if_strd_address_reg[4]  <= 1'b0;
    \\pci_target_unit_pci_target_if_strd_address_reg[7]  <= 1'b0;
    \\pci_target_unit_pci_target_if_strd_address_reg[9]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[5]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[1]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[6]  <= 1'b0;
    \\pci_target_unit_pci_target_if_strd_address_reg[5]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_cycle_count_reg[0]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[2]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[11]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[22]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[21]  <= 1'b0;
    \\pci_target_unit_del_sync_bc_out_reg[1]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[16]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[22]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[23]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[24]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[25]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[16]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[17]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[10]  <= 1'b0;
    \\pci_target_unit_del_sync_be_out_reg[1]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[30]  <= 1'b0;
    \\input_register_pci_cbe_reg_out_reg[3]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[14]  <= 1'b0;
    \\input_register_pci_cbe_reg_out_reg[2]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[28]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[27]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[13]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_bc_reg[3]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_bc_reg[2]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[2]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_sm_mabort1_reg <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[26]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[25]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[24]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[23]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[28]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[20]  <= 1'b0;
    pci_target_unit_del_sync_burst_out_reg <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[4]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[5]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[7]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[21]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[12]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[31]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[26]  <= 1'b0;
    input_register_pci_trdy_reg_out_reg <= 1'b1;
    \\pci_target_unit_pci_target_if_norm_address_reg[15]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[27]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[13]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[9]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[21]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[3]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[20]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[27]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[31]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[8]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[4]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[6]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[1]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[29]  <= 1'b0;
    \\input_register_pci_cbe_reg_out_reg[1]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[30]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[26]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[22]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[18]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[12]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[29]  <= 1'b0;
    \\pci_target_unit_del_sync_be_out_reg[2]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[20]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[1]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[14]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[6]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[11]  <= 1'b0;
    \\pci_target_unit_del_sync_be_out_reg[3]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[19]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[15]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[30]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[8]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[3]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[19]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[13]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[18]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[12]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[10]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[0]  <= 1'b0;
    pci_target_unit_pci_target_sm_state_backoff_reg_reg <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[10]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[11]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[16]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[19]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[23]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[28]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[2]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg[2]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[3]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[5]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[7]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[9]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[31]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[24]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[14]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[15]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[25]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg[17]  <= 1'b0;
    \\pci_target_unit_del_sync_bc_out_reg[3]  <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[2]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[9]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[5]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[4]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[0]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[8]  <= 1'b0;
    \\pci_target_unit_pci_target_if_strd_address_reg[0]  <= 1'b0;
    \\pci_target_unit_pci_target_if_norm_address_reg[7]  <= 1'b0;
    \\pci_target_unit_del_sync_bc_out_reg[0]  <= 1'b0;
    \\pci_target_unit_del_sync_bc_out_reg[2]  <= 1'b1;
    \\pci_target_unit_del_sync_addr_out_reg[29]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[18]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[0]  <= 1'b0;
    \\pci_target_unit_del_sync_addr_out_reg[17]  <= 1'b0;
    input_register_pci_frame_reg_out_reg <= 1'b0;
    input_register_pci_devsel_reg_out_reg <= 1'b1;
    pci_io_mux_irdy_iob_dat_out_reg <= 1'b0;
    input_register_pci_irdy_reg_out_reg <= 1'b1;
    output_backup_irdy_out_reg <= 1'b1;
    \\wishbone_slave_unit_del_sync_rty_exp_back_prop_sync_sync_data_out_reg[0]  <= 1'b0;
    pci_target_unit_del_sync_req_req_pending_reg <= 1'b0;
    input_register_pci_stop_reg_out_reg <= 1'b1;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[8]  <= 1'b0;
    configuration_interrupt_out_reg <= 1'b0;
    pci_io_mux_req_iob_dat_out_reg <= 1'b0;
    \\pci_target_unit_pci_target_if_pciw_fifo_control_out_reg[3]  <= 1'b0;
    pci_target_unit_pci_target_sm_state_transfere_reg_reg <= 1'b0;
    pci_target_unit_pci_target_sm_previous_frame_reg <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[7]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[17]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[30]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[16]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[28]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[0]  <= 1'b0;
    \\configuration_int_pin_sync_sync_data_out_reg[0]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[24]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[10]  <= 1'b0;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[6]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[12]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[3]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[13]  <= 1'b0;
    parity_checker_master_perr_report_reg <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[4]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[9]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[14]  <= 1'b0;
    pci_target_unit_del_sync_comp_done_reg_clr_reg <= 1'b0;
    configuration_wb_init_complete_out_reg <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[29]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[25]  <= 1'b0;
    parity_checker_frame_dec2_reg <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[15]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[23]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[20]  <= 1'b0;
    wishbone_slave_unit_del_sync_req_rty_exp_clr_reg <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[26]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[31]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[6]  <= 1'b0;
    configuration_init_complete_reg <= 1'b0;
    input_register_pci_idsel_reg_out_reg <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[21]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[1]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[18]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[22]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[2]  <= 1'b0;
    pci_target_unit_pci_target_sm_read_completed_reg_reg <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[11]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[5]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[8]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[19]  <= 1'b0;
    \\input_register_pci_ad_reg_out_reg[27]  <= 1'b0;
    parity_checker_frame_and_irdy_en_prev_prev_reg <= 1'b0;
    wishbone_slave_unit_del_sync_comp_done_reg_main_reg <= 1'b0;
    pci_target_unit_del_sync_comp_rty_exp_clr_reg <= 1'b0;
    configuration_pci_err_cs_bit8_reg <= 1'b0;
    \\configuration_isr_bit2_0_reg[2]  <= 1'b0;
    \\configuration_isr_bit2_0_reg[0]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_if_write_req_int_reg <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[0]  <= 1'b0;
    \\configuration_i_wb_init_complete_sync_sync_data_out_reg[0]  <= 1'b0;
    configuration_sync_isr_2_sync_del_bit_reg <= 1'b0;
    pci_io_mux_req_iob_en_out_reg <= 1'b1;
    pci_target_unit_del_sync_req_rty_exp_reg_reg <= 1'b0;
    configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg <= 1'b0;
    configuration_sync_isr_2_delayed_bckp_bit_reg <= 1'b0;
    wishbone_slave_unit_del_sync_req_comp_pending_sample_reg <= 1'b0;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[3]  <= 1'b0;
    pci_target_unit_del_sync_req_comp_pending_sample_reg <= 1'b0;
    \\pci_target_unit_del_sync_req_sync_sync_data_out_reg[0]  <= 1'b0;
    pci_target_unit_del_sync_comp_done_reg_main_reg <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[0]  <= 1'b0;
    pci_io_mux_irdy_iob_en_out_reg <= 1'b1;
    \\pci_target_unit_del_sync_rty_exp_back_prop_sync_sync_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_req_sync_sync_data_out_reg[0]  <= 1'b0;
    wishbone_slave_unit_pci_initiator_sm_mabort2_reg <= 1'b0;
    \\wishbone_slave_unit_del_sync_done_sync_sync_data_out_reg[0]  <= 1'b0;
    pci_target_unit_del_sync_comp_flush_out_reg <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[0]  <= 1'b0;
    wishbone_slave_unit_del_sync_comp_flush_out_reg <= 1'b0;
    pci_target_unit_pci_target_sm_bckp_trdy_reg_reg <= 1'b1;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg[3]  <= 1'b0;
    configuration_sync_pci_err_cs_8_sync_del_bit_reg <= 1'b0;
    parity_checker_frame_and_irdy_en_prev_reg <= 1'b0;
    \\configuration_isr_bit0_sync_sync_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[1]  <= 1'b0;
    \\configuration_pci_err_cs_bits_sync_sync_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[3]  <= 1'b0;
    \\pci_target_unit_fifos_wb_clk_inGreyCount_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_wb_clk_inGreyCount_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg[1]  <= 1'b0;
    \\configuration_isr_bit2_sync_sync_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[0]  <= 1'b1;
    output_backup_irdy_en_out_reg <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[3]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[1]  <= 1'b1;
    \\wishbone_slave_unit_del_sync_comp_sync_sync_data_out_reg[0]  <= 1'b0;
    \\pci_target_unit_del_sync_comp_sync_sync_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[1]  <= 1'b1;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[1]  <= 1'b0;
    \\pci_target_unit_del_sync_rty_exp_sync_sync_data_out_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg[2]  <= 1'b0;
    \\configuration_sync_isr_2_delete_sync_sync_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg[2]  <= 1'b0;
    \\pci_target_unit_del_sync_done_sync_sync_data_out_reg[0]  <= 1'b0;
    pci_target_unit_del_sync_req_rty_exp_clr_reg <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg[2]  <= 1'b0;
    configuration_rst_inactive_reg <= 1'b0;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[2]  <= 1'b0;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[4]  <= 1'b0;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[7]  <= 1'b0;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[5]  <= 1'b0;
    configuration_sync_command_bit_reg <= 1'b0;
    \\configuration_sync_cache_lsize_to_wb_bits_reg[6]  <= 1'b0;
    configuration_sync_isr_2_sync_bckp_bit_reg <= 1'b0;
    wishbone_slave_unit_del_sync_req_rty_exp_reg_reg <= 1'b0;
    configuration_sync_pci_err_cs_8_sync_bckp_bit_reg <= 1'b0;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[2]  <= 1'b0;
    pci_target_unit_wishbone_master_burst_chopped_delayed_reg <= 1'b0;
    \\wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[1]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[2]  <= 1'b0;
    \\configuration_sync_pci_err_cs_8_delete_sync_sync_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[18]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[31]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[4]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[25]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[6]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[16]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[11]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[15]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[14]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg[0]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[2]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[13]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[11]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[10]  <= 1'b0;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg[2]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[15]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[8]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[0]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[6]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[21]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[25]  <= 1'b0;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[0]  <= 1'b0;
    \\configuration_sync_isr_2_clear_delete_sync_sync_data_out_reg[0]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[19]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[30]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[27]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[29]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[3]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[19]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[23]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[22]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[28]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[24]  <= 1'b0;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[4]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[5]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[4]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[13]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[8]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[16]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[17]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[1]  <= 1'b0;
    configuration_rst_inactive_sync_reg <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[26]  <= 1'b0;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[5]  <= 1'b0;
    configuration_sync_isr_2_delayed_del_bit_reg <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[22]  <= 1'b0;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[2]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[1]  <= 1'b1;
    \\pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg[1]  <= 1'b0;
    \\wishbone_slave_unit_del_sync_rty_exp_sync_sync_data_out_reg[0]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[23]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[20]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[12]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[12]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[21]  <= 1'b0;
    \\pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg[0]  <= 1'b1;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[7]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[20]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[26]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[9]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[24]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[7]  <= 1'b0;
    \\configuration_command_bit_sync_sync_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[0]  <= 1'b1;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[14]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[31]  <= 1'b0;
    \\wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg[1]  <= 1'b1;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[0]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[10]  <= 1'b0;
    \\configuration_sync_pci_err_cs_8_clear_delete_sync_sync_data_out_reg[0]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[3]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[18]  <= 1'b0;
    wishbone_slave_unit_del_sync_comp_done_reg_clr_reg <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[27]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[28]  <= 1'b0;
    configuration_sync_pci_err_cs_8_delayed_del_bit_reg <= 1'b0;
    \\configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg[3]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[5]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[29]  <= 1'b0;
    \\pci_target_unit_wishbone_master_pcir_fifo_data_out_reg[2]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[17]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[9]  <= 1'b0;
    \\wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg[30]  <= 1'b0;
  end
endmodule


