// Benchmark "testing" written by ABC on Thu Oct  8 22:16:44 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A109  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A109;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ ,
    \new_[441]_ , \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ ,
    \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[450]_ ,
    \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ , \new_[455]_ ,
    \new_[456]_ , \new_[457]_ , \new_[458]_ , \new_[459]_ , \new_[460]_ ,
    \new_[461]_ , \new_[462]_ , \new_[463]_ , \new_[464]_ , \new_[465]_ ,
    \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[469]_ , \new_[470]_ ,
    \new_[471]_ , \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[477]_ , \new_[478]_ , \new_[479]_ , \new_[480]_ ,
    \new_[481]_ , \new_[482]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ ,
    \new_[486]_ , \new_[487]_ , \new_[488]_ , \new_[489]_ , \new_[490]_ ,
    \new_[491]_ , \new_[492]_ , \new_[493]_ , \new_[494]_ , \new_[495]_ ,
    \new_[496]_ , \new_[497]_ , \new_[498]_ , \new_[499]_ , \new_[500]_ ,
    \new_[501]_ , \new_[502]_ , \new_[503]_ , \new_[504]_ , \new_[505]_ ,
    \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ , \new_[510]_ ,
    \new_[511]_ , \new_[512]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ ,
    \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ ,
    \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ ,
    \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ ,
    \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ ,
    \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ ,
    \new_[686]_ , \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ ,
    \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ ,
    \new_[696]_ , \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ ,
    \new_[701]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ ,
    \new_[706]_ , \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ ,
    \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ ,
    \new_[716]_ , \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[726]_ , \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ ,
    \new_[731]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ ,
    \new_[741]_ , \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[746]_ , \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ ,
    \new_[751]_ , \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ ,
    \new_[756]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ ,
    \new_[766]_ , \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ ,
    \new_[771]_ , \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ ,
    \new_[776]_ , \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ ,
    \new_[781]_ , \new_[782]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ ,
    \new_[786]_ , \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ ,
    \new_[791]_ , \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ ,
    \new_[796]_ , \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ ,
    \new_[801]_ , \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ ,
    \new_[806]_ , \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ ,
    \new_[811]_ , \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ ,
    \new_[816]_ , \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[824]_ , \new_[825]_ ,
    \new_[826]_ , \new_[827]_ , \new_[828]_ , \new_[829]_ , \new_[830]_ ,
    \new_[831]_ , \new_[832]_ , \new_[833]_ , \new_[834]_ , \new_[835]_ ,
    \new_[836]_ , \new_[837]_ , \new_[838]_ , \new_[839]_ , \new_[840]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[845]_ ,
    \new_[846]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ , \new_[850]_ ,
    \new_[851]_ , \new_[852]_ , \new_[853]_ , \new_[854]_ , \new_[855]_ ,
    \new_[856]_ , \new_[857]_ , \new_[858]_ , \new_[859]_ , \new_[860]_ ,
    \new_[861]_ , \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ ,
    \new_[866]_ , \new_[867]_ , \new_[868]_ , \new_[869]_ , \new_[870]_ ,
    \new_[871]_ , \new_[872]_ , \new_[873]_ , \new_[874]_ , \new_[875]_ ,
    \new_[876]_ , \new_[877]_ , \new_[878]_ , \new_[879]_ , \new_[880]_ ,
    \new_[881]_ , \new_[882]_ , \new_[883]_ , \new_[884]_ , \new_[885]_ ,
    \new_[886]_ , \new_[887]_ , \new_[888]_ , \new_[889]_ , \new_[890]_ ,
    \new_[891]_ , \new_[892]_ , \new_[893]_ , \new_[894]_ , \new_[895]_ ,
    \new_[896]_ , \new_[897]_ , \new_[898]_ , \new_[899]_ , \new_[900]_ ,
    \new_[901]_ , \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ ,
    \new_[906]_ , \new_[907]_ , \new_[908]_ , \new_[909]_ , \new_[910]_ ,
    \new_[911]_ , \new_[912]_ , \new_[913]_ , \new_[914]_ , \new_[915]_ ,
    \new_[916]_ , \new_[917]_ , \new_[918]_ , \new_[919]_ , \new_[920]_ ,
    \new_[921]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[925]_ ,
    \new_[926]_ , \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ ,
    \new_[931]_ , \new_[932]_ , \new_[933]_ , \new_[934]_ , \new_[935]_ ,
    \new_[936]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ , \new_[940]_ ,
    \new_[941]_ , \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ ,
    \new_[946]_ , \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ ,
    \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ ,
    \new_[956]_ , \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ ,
    \new_[961]_ , \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ ,
    \new_[966]_ , \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ ,
    \new_[971]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ ,
    \new_[976]_ , \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ ,
    \new_[986]_ , \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ ,
    \new_[996]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1002]_ , \new_[1003]_ , \new_[1004]_ ,
    \new_[1005]_ , \new_[1006]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1009]_ , \new_[1010]_ , \new_[1011]_ , \new_[1012]_ ,
    \new_[1013]_ , \new_[1014]_ , \new_[1015]_ , \new_[1016]_ ,
    \new_[1017]_ , \new_[1018]_ , \new_[1019]_ , \new_[1020]_ ,
    \new_[1021]_ , \new_[1022]_ , \new_[1023]_ , \new_[1024]_ ,
    \new_[1025]_ , \new_[1026]_ , \new_[1027]_ , \new_[1028]_ ,
    \new_[1029]_ , \new_[1030]_ , \new_[1031]_ , \new_[1032]_ ,
    \new_[1033]_ , \new_[1034]_ , \new_[1035]_ , \new_[1036]_ ,
    \new_[1037]_ , \new_[1038]_ , \new_[1039]_ , \new_[1040]_ ,
    \new_[1041]_ , \new_[1042]_ , \new_[1043]_ , \new_[1044]_ ,
    \new_[1045]_ , \new_[1046]_ , \new_[1047]_ , \new_[1048]_ ,
    \new_[1049]_ , \new_[1050]_ , \new_[1051]_ , \new_[1052]_ ,
    \new_[1053]_ , \new_[1054]_ , \new_[1055]_ , \new_[1056]_ ,
    \new_[1057]_ , \new_[1058]_ , \new_[1059]_ , \new_[1060]_ ,
    \new_[1061]_ , \new_[1062]_ , \new_[1063]_ , \new_[1064]_ ,
    \new_[1065]_ , \new_[1066]_ , \new_[1067]_ , \new_[1068]_ ,
    \new_[1069]_ , \new_[1070]_ , \new_[1071]_ , \new_[1072]_ ,
    \new_[1073]_ , \new_[1074]_ , \new_[1075]_ , \new_[1076]_ ,
    \new_[1077]_ , \new_[1078]_ , \new_[1079]_ , \new_[1080]_ ,
    \new_[1081]_ , \new_[1082]_ , \new_[1083]_ , \new_[1084]_ ,
    \new_[1085]_ , \new_[1086]_ , \new_[1087]_ , \new_[1088]_ ,
    \new_[1089]_ , \new_[1090]_ , \new_[1091]_ , \new_[1092]_ ,
    \new_[1093]_ , \new_[1094]_ , \new_[1095]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1098]_ , \new_[1099]_ , \new_[1100]_ ,
    \new_[1101]_ , \new_[1102]_ , \new_[1103]_ , \new_[1104]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1107]_ , \new_[1108]_ ,
    \new_[1109]_ , \new_[1110]_ , \new_[1111]_ , \new_[1112]_ ,
    \new_[1113]_ , \new_[1114]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1118]_ , \new_[1119]_ , \new_[1120]_ ,
    \new_[1121]_ , \new_[1122]_ , \new_[1123]_ , \new_[1124]_ ,
    \new_[1125]_ , \new_[1126]_ , \new_[1127]_ , \new_[1128]_ ,
    \new_[1129]_ , \new_[1130]_ , \new_[1131]_ , \new_[1132]_ ,
    \new_[1133]_ , \new_[1134]_ , \new_[1135]_ , \new_[1136]_ ,
    \new_[1137]_ , \new_[1138]_ , \new_[1139]_ , \new_[1140]_ ,
    \new_[1141]_ , \new_[1142]_ , \new_[1143]_ , \new_[1144]_ ,
    \new_[1145]_ , \new_[1146]_ , \new_[1147]_ , \new_[1148]_ ,
    \new_[1149]_ , \new_[1150]_ , \new_[1151]_ , \new_[1152]_ ,
    \new_[1153]_ , \new_[1154]_ , \new_[1155]_ , \new_[1156]_ ,
    \new_[1157]_ , \new_[1158]_ , \new_[1159]_ , \new_[1160]_ ,
    \new_[1161]_ , \new_[1162]_ , \new_[1163]_ , \new_[1164]_ ,
    \new_[1165]_ , \new_[1166]_ , \new_[1167]_ , \new_[1168]_ ,
    \new_[1169]_ , \new_[1170]_ , \new_[1171]_ , \new_[1172]_ ,
    \new_[1173]_ , \new_[1174]_ , \new_[1175]_ , \new_[1176]_ ,
    \new_[1177]_ , \new_[1178]_ , \new_[1179]_ , \new_[1180]_ ,
    \new_[1181]_ , \new_[1182]_ , \new_[1183]_ , \new_[1184]_ ,
    \new_[1185]_ , \new_[1186]_ , \new_[1187]_ , \new_[1188]_ ,
    \new_[1189]_ , \new_[1190]_ , \new_[1191]_ , \new_[1192]_ ,
    \new_[1193]_ , \new_[1194]_ , \new_[1195]_ , \new_[1196]_ ,
    \new_[1197]_ , \new_[1198]_ , \new_[1199]_ , \new_[1200]_ ,
    \new_[1201]_ , \new_[1202]_ , \new_[1203]_ , \new_[1204]_ ,
    \new_[1205]_ , \new_[1206]_ , \new_[1207]_ , \new_[1208]_ ,
    \new_[1209]_ , \new_[1210]_ , \new_[1211]_ , \new_[1212]_ ,
    \new_[1213]_ , \new_[1214]_ , \new_[1215]_ , \new_[1216]_ ,
    \new_[1217]_ , \new_[1218]_ , \new_[1219]_ , \new_[1220]_ ,
    \new_[1221]_ , \new_[1222]_ , \new_[1223]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1226]_ , \new_[1227]_ , \new_[1228]_ ,
    \new_[1229]_ , \new_[1230]_ , \new_[1231]_ , \new_[1232]_ ,
    \new_[1233]_ , \new_[1234]_ , \new_[1235]_ , \new_[1236]_ ,
    \new_[1237]_ , \new_[1238]_ , \new_[1239]_ , \new_[1240]_ ,
    \new_[1241]_ , \new_[1242]_ , \new_[1243]_ , \new_[1244]_ ,
    \new_[1245]_ , \new_[1246]_ , \new_[1247]_ , \new_[1248]_ ,
    \new_[1249]_ , \new_[1250]_ , \new_[1251]_ , \new_[1252]_ ,
    \new_[1253]_ , \new_[1254]_ , \new_[1255]_ , \new_[1256]_ ,
    \new_[1257]_ , \new_[1258]_ , \new_[1259]_ , \new_[1260]_ ,
    \new_[1261]_ , \new_[1262]_ , \new_[1263]_ , \new_[1264]_ ,
    \new_[1265]_ , \new_[1266]_ , \new_[1267]_ , \new_[1268]_ ,
    \new_[1269]_ , \new_[1270]_ , \new_[1271]_ , \new_[1272]_ ,
    \new_[1273]_ , \new_[1274]_ , \new_[1275]_ , \new_[1276]_ ,
    \new_[1277]_ , \new_[1278]_ , \new_[1279]_ , \new_[1280]_ ,
    \new_[1281]_ , \new_[1282]_ , \new_[1283]_ , \new_[1284]_ ,
    \new_[1285]_ , \new_[1286]_ , \new_[1287]_ , \new_[1288]_ ,
    \new_[1289]_ , \new_[1290]_ , \new_[1291]_ , \new_[1292]_ ,
    \new_[1293]_ , \new_[1294]_ , \new_[1295]_ , \new_[1296]_ ,
    \new_[1297]_ , \new_[1298]_ , \new_[1299]_ , \new_[1300]_ ,
    \new_[1301]_ , \new_[1302]_ , \new_[1303]_ , \new_[1304]_ ,
    \new_[1305]_ , \new_[1306]_ , \new_[1307]_ , \new_[1308]_ ,
    \new_[1309]_ , \new_[1310]_ , \new_[1311]_ , \new_[1312]_ ,
    \new_[1313]_ , \new_[1314]_ , \new_[1315]_ , \new_[1316]_ ,
    \new_[1317]_ , \new_[1318]_ , \new_[1319]_ , \new_[1320]_ ,
    \new_[1321]_ , \new_[1322]_ , \new_[1323]_ , \new_[1324]_ ,
    \new_[1325]_ , \new_[1326]_ , \new_[1327]_ , \new_[1328]_ ,
    \new_[1329]_ , \new_[1330]_ , \new_[1331]_ , \new_[1332]_ ,
    \new_[1333]_ , \new_[1334]_ , \new_[1335]_ , \new_[1336]_ ,
    \new_[1337]_ , \new_[1338]_ , \new_[1339]_ , \new_[1340]_ ,
    \new_[1341]_ , \new_[1342]_ , \new_[1343]_ , \new_[1344]_ ,
    \new_[1345]_ , \new_[1346]_ , \new_[1347]_ , \new_[1348]_ ,
    \new_[1349]_ , \new_[1350]_ , \new_[1351]_ , \new_[1352]_ ,
    \new_[1353]_ , \new_[1354]_ , \new_[1355]_ , \new_[1356]_ ,
    \new_[1357]_ , \new_[1358]_ , \new_[1359]_ , \new_[1360]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1363]_ , \new_[1364]_ ,
    \new_[1365]_ , \new_[1366]_ , \new_[1367]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1370]_ , \new_[1371]_ , \new_[1372]_ ,
    \new_[1373]_ , \new_[1374]_ , \new_[1375]_ , \new_[1376]_ ,
    \new_[1377]_ , \new_[1378]_ , \new_[1379]_ , \new_[1380]_ ,
    \new_[1381]_ , \new_[1382]_ , \new_[1383]_ , \new_[1384]_ ,
    \new_[1385]_ , \new_[1386]_ , \new_[1387]_ , \new_[1388]_ ,
    \new_[1389]_ , \new_[1390]_ , \new_[1391]_ , \new_[1392]_ ,
    \new_[1393]_ , \new_[1394]_ , \new_[1395]_ , \new_[1396]_ ,
    \new_[1397]_ , \new_[1398]_ , \new_[1399]_ , \new_[1400]_ ,
    \new_[1401]_ , \new_[1402]_ , \new_[1403]_ , \new_[1404]_ ,
    \new_[1405]_ , \new_[1406]_ , \new_[1407]_ , \new_[1408]_ ,
    \new_[1409]_ , \new_[1410]_ , \new_[1411]_ , \new_[1412]_ ,
    \new_[1413]_ , \new_[1414]_ , \new_[1415]_ , \new_[1416]_ ,
    \new_[1417]_ , \new_[1418]_ , \new_[1419]_ , \new_[1420]_ ,
    \new_[1421]_ , \new_[1422]_ , \new_[1423]_ , \new_[1424]_ ,
    \new_[1425]_ , \new_[1426]_ , \new_[1427]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1430]_ , \new_[1431]_ , \new_[1432]_ ,
    \new_[1433]_ , \new_[1434]_ , \new_[1435]_ , \new_[1436]_ ,
    \new_[1437]_ , \new_[1438]_ , \new_[1439]_ , \new_[1440]_ ,
    \new_[1441]_ , \new_[1442]_ , \new_[1443]_ , \new_[1444]_ ,
    \new_[1445]_ , \new_[1446]_ , \new_[1447]_ , \new_[1448]_ ,
    \new_[1449]_ , \new_[1450]_ , \new_[1451]_ , \new_[1452]_ ,
    \new_[1453]_ , \new_[1454]_ , \new_[1455]_ , \new_[1456]_ ,
    \new_[1457]_ , \new_[1458]_ , \new_[1459]_ , \new_[1460]_ ,
    \new_[1461]_ , \new_[1462]_ , \new_[1463]_ , \new_[1464]_ ,
    \new_[1465]_ , \new_[1466]_ , \new_[1467]_ , \new_[1468]_ ,
    \new_[1469]_ , \new_[1470]_ , \new_[1471]_ , \new_[1472]_ ,
    \new_[1473]_ , \new_[1474]_ , \new_[1475]_ , \new_[1476]_ ,
    \new_[1477]_ , \new_[1478]_ , \new_[1479]_ , \new_[1480]_ ,
    \new_[1481]_ , \new_[1482]_ , \new_[1483]_ , \new_[1484]_ ,
    \new_[1485]_ , \new_[1486]_ , \new_[1487]_ , \new_[1488]_ ,
    \new_[1489]_ , \new_[1490]_ , \new_[1491]_ , \new_[1492]_ ,
    \new_[1493]_ , \new_[1494]_ , \new_[1495]_ , \new_[1496]_ ,
    \new_[1497]_ , \new_[1498]_ , \new_[1499]_ , \new_[1500]_ ,
    \new_[1501]_ , \new_[1502]_ , \new_[1503]_ , \new_[1504]_ ,
    \new_[1505]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1514]_ , \new_[1515]_ , \new_[1516]_ ,
    \new_[1517]_ , \new_[1518]_ , \new_[1519]_ , \new_[1520]_ ,
    \new_[1521]_ , \new_[1522]_ , \new_[1523]_ , \new_[1524]_ ,
    \new_[1525]_ , \new_[1526]_ , \new_[1527]_ , \new_[1528]_ ,
    \new_[1529]_ , \new_[1530]_ , \new_[1531]_ , \new_[1532]_ ,
    \new_[1533]_ , \new_[1534]_ , \new_[1535]_ , \new_[1536]_ ,
    \new_[1537]_ , \new_[1538]_ , \new_[1539]_ , \new_[1540]_ ,
    \new_[1541]_ , \new_[1542]_ , \new_[1543]_ , \new_[1544]_ ,
    \new_[1545]_ , \new_[1546]_ , \new_[1547]_ , \new_[1548]_ ,
    \new_[1549]_ , \new_[1550]_ , \new_[1551]_ , \new_[1552]_ ,
    \new_[1553]_ , \new_[1554]_ , \new_[1555]_ , \new_[1556]_ ,
    \new_[1557]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1563]_ , \new_[1564]_ ,
    \new_[1565]_ , \new_[1566]_ , \new_[1567]_ , \new_[1568]_ ,
    \new_[1569]_ , \new_[1570]_ , \new_[1571]_ , \new_[1572]_ ,
    \new_[1573]_ , \new_[1574]_ , \new_[1575]_ , \new_[1576]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1579]_ , \new_[1580]_ ,
    \new_[1581]_ , \new_[1582]_ , \new_[1583]_ , \new_[1584]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1587]_ , \new_[1588]_ ,
    \new_[1589]_ , \new_[1590]_ , \new_[1591]_ , \new_[1592]_ ,
    \new_[1593]_ , \new_[1594]_ , \new_[1595]_ , \new_[1596]_ ,
    \new_[1597]_ , \new_[1598]_ , \new_[1599]_ , \new_[1600]_ ,
    \new_[1601]_ , \new_[1602]_ , \new_[1603]_ , \new_[1604]_ ,
    \new_[1605]_ , \new_[1606]_ , \new_[1607]_ , \new_[1608]_ ,
    \new_[1609]_ , \new_[1610]_ , \new_[1611]_ , \new_[1612]_ ,
    \new_[1613]_ , \new_[1614]_ , \new_[1615]_ , \new_[1616]_ ,
    \new_[1617]_ , \new_[1618]_ , \new_[1619]_ , \new_[1620]_ ,
    \new_[1621]_ , \new_[1622]_ , \new_[1623]_ , \new_[1624]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1627]_ , \new_[1628]_ ,
    \new_[1629]_ , \new_[1630]_ , \new_[1631]_ , \new_[1632]_ ,
    \new_[1633]_ , \new_[1634]_ , \new_[1635]_ , \new_[1636]_ ,
    \new_[1637]_ , \new_[1638]_ , \new_[1639]_ , \new_[1640]_ ,
    \new_[1641]_ , \new_[1642]_ , \new_[1643]_ , \new_[1644]_ ,
    \new_[1645]_ , \new_[1646]_ , \new_[1647]_ , \new_[1648]_ ,
    \new_[1649]_ , \new_[1650]_ , \new_[1651]_ , \new_[1652]_ ,
    \new_[1653]_ , \new_[1654]_ , \new_[1655]_ , \new_[1656]_ ,
    \new_[1657]_ , \new_[1658]_ , \new_[1659]_ , \new_[1660]_ ,
    \new_[1661]_ , \new_[1662]_ , \new_[1663]_ , \new_[1664]_ ,
    \new_[1665]_ , \new_[1666]_ , \new_[1667]_ , \new_[1668]_ ,
    \new_[1669]_ , \new_[1670]_ , \new_[1671]_ , \new_[1672]_ ,
    \new_[1673]_ , \new_[1674]_ , \new_[1675]_ , \new_[1676]_ ,
    \new_[1677]_ , \new_[1678]_ , \new_[1679]_ , \new_[1680]_ ,
    \new_[1681]_ , \new_[1682]_ , \new_[1683]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1686]_ , \new_[1687]_ , \new_[1688]_ ,
    \new_[1689]_ , \new_[1690]_ , \new_[1691]_ , \new_[1692]_ ,
    \new_[1693]_ , \new_[1694]_ , \new_[1695]_ , \new_[1696]_ ,
    \new_[1697]_ , \new_[1698]_ , \new_[1699]_ , \new_[1700]_ ,
    \new_[1701]_ , \new_[1702]_ , \new_[1703]_ , \new_[1704]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1707]_ , \new_[1708]_ ,
    \new_[1709]_ , \new_[1710]_ , \new_[1711]_ , \new_[1712]_ ,
    \new_[1713]_ , \new_[1714]_ , \new_[1715]_ , \new_[1716]_ ,
    \new_[1717]_ , \new_[1718]_ , \new_[1719]_ , \new_[1720]_ ,
    \new_[1721]_ , \new_[1722]_ , \new_[1723]_ , \new_[1724]_ ,
    \new_[1725]_ , \new_[1726]_ , \new_[1727]_ , \new_[1728]_ ,
    \new_[1729]_ , \new_[1730]_ , \new_[1731]_ , \new_[1732]_ ,
    \new_[1733]_ , \new_[1734]_ , \new_[1735]_ , \new_[1736]_ ,
    \new_[1737]_ , \new_[1738]_ , \new_[1739]_ , \new_[1740]_ ,
    \new_[1741]_ , \new_[1742]_ , \new_[1743]_ , \new_[1744]_ ,
    \new_[1745]_ , \new_[1746]_ , \new_[1747]_ , \new_[1748]_ ,
    \new_[1749]_ , \new_[1750]_ , \new_[1751]_ , \new_[1752]_ ,
    \new_[1753]_ , \new_[1754]_ , \new_[1755]_ , \new_[1756]_ ,
    \new_[1757]_ , \new_[1758]_ , \new_[1759]_ , \new_[1760]_ ,
    \new_[1761]_ , \new_[1762]_ , \new_[1763]_ , \new_[1764]_ ,
    \new_[1765]_ , \new_[1766]_ , \new_[1767]_ , \new_[1768]_ ,
    \new_[1769]_ , \new_[1770]_ , \new_[1771]_ , \new_[1772]_ ,
    \new_[1773]_ , \new_[1774]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1780]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1783]_ , \new_[1784]_ ,
    \new_[1785]_ , \new_[1786]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1792]_ ,
    \new_[1793]_ , \new_[1794]_ , \new_[1795]_ , \new_[1796]_ ,
    \new_[1797]_ , \new_[1798]_ , \new_[1799]_ , \new_[1800]_ ,
    \new_[1801]_ , \new_[1802]_ , \new_[1803]_ , \new_[1804]_ ,
    \new_[1805]_ , \new_[1806]_ , \new_[1807]_ , \new_[1808]_ ,
    \new_[1809]_ , \new_[1810]_ , \new_[1811]_ , \new_[1812]_ ,
    \new_[1813]_ , \new_[1814]_ , \new_[1815]_ , \new_[1816]_ ,
    \new_[1817]_ , \new_[1818]_ , \new_[1819]_ , \new_[1820]_ ,
    \new_[1821]_ , \new_[1822]_ , \new_[1823]_ , \new_[1824]_ ,
    \new_[1825]_ , \new_[1826]_ , \new_[1827]_ , \new_[1828]_ ,
    \new_[1829]_ , \new_[1830]_ , \new_[1831]_ , \new_[1832]_ ,
    \new_[1833]_ , \new_[1834]_ , \new_[1835]_ , \new_[1836]_ ,
    \new_[1837]_ , \new_[1838]_ , \new_[1839]_ , \new_[1840]_ ,
    \new_[1841]_ , \new_[1842]_ , \new_[1843]_ , \new_[1844]_ ,
    \new_[1845]_ , \new_[1846]_ , \new_[1847]_ , \new_[1848]_ ,
    \new_[1849]_ , \new_[1850]_ , \new_[1851]_ , \new_[1852]_ ,
    \new_[1853]_ , \new_[1854]_ , \new_[1855]_ , \new_[1856]_ ,
    \new_[1857]_ , \new_[1858]_ , \new_[1859]_ , \new_[1860]_ ,
    \new_[1861]_ , \new_[1862]_ , \new_[1863]_ , \new_[1864]_ ,
    \new_[1865]_ , \new_[1866]_ , \new_[1867]_ , \new_[1868]_ ,
    \new_[1869]_ , \new_[1870]_ , \new_[1871]_ , \new_[1872]_ ,
    \new_[1873]_ , \new_[1874]_ , \new_[1875]_ , \new_[1876]_ ,
    \new_[1877]_ , \new_[1878]_ , \new_[1879]_ , \new_[1880]_ ,
    \new_[1881]_ , \new_[1882]_ , \new_[1883]_ , \new_[1884]_ ,
    \new_[1885]_ , \new_[1886]_ , \new_[1887]_ , \new_[1888]_ ,
    \new_[1889]_ , \new_[1890]_ , \new_[1891]_ , \new_[1892]_ ,
    \new_[1893]_ , \new_[1894]_ , \new_[1895]_ , \new_[1896]_ ,
    \new_[1897]_ , \new_[1898]_ , \new_[1899]_ , \new_[1900]_ ,
    \new_[1901]_ , \new_[1902]_ , \new_[1903]_ , \new_[1904]_ ,
    \new_[1905]_ , \new_[1906]_ , \new_[1907]_ , \new_[1908]_ ,
    \new_[1909]_ , \new_[1910]_ , \new_[1911]_ , \new_[1912]_ ,
    \new_[1913]_ , \new_[1914]_ , \new_[1915]_ , \new_[1916]_ ,
    \new_[1917]_ , \new_[1918]_ , \new_[1919]_ , \new_[1920]_ ,
    \new_[1921]_ , \new_[1922]_ , \new_[1923]_ , \new_[1924]_ ,
    \new_[1925]_ , \new_[1926]_ , \new_[1927]_ , \new_[1928]_ ,
    \new_[1929]_ , \new_[1930]_ , \new_[1931]_ , \new_[1932]_ ,
    \new_[1933]_ , \new_[1934]_ , \new_[1935]_ , \new_[1936]_ ,
    \new_[1937]_ , \new_[1938]_ , \new_[1939]_ , \new_[1940]_ ,
    \new_[1941]_ , \new_[1942]_ , \new_[1943]_ , \new_[1944]_ ,
    \new_[1945]_ , \new_[1946]_ , \new_[1947]_ , \new_[1948]_ ,
    \new_[1949]_ , \new_[1950]_ , \new_[1951]_ , \new_[1952]_ ,
    \new_[1953]_ , \new_[1954]_ , \new_[1955]_ , \new_[1956]_ ,
    \new_[1957]_ , \new_[1958]_ , \new_[1959]_ , \new_[1960]_ ,
    \new_[1961]_ , \new_[1962]_ , \new_[1963]_ , \new_[1964]_ ,
    \new_[1965]_ , \new_[1966]_ , \new_[1967]_ , \new_[1968]_ ,
    \new_[1969]_ , \new_[1970]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1978]_ , \new_[1979]_ , \new_[1980]_ ,
    \new_[1981]_ , \new_[1982]_ , \new_[1983]_ , \new_[1984]_ ,
    \new_[1985]_ , \new_[1986]_ , \new_[1987]_ , \new_[1988]_ ,
    \new_[1989]_ , \new_[1990]_ , \new_[1991]_ , \new_[1992]_ ,
    \new_[1993]_ , \new_[1994]_ , \new_[1995]_ , \new_[1996]_ ,
    \new_[1997]_ , \new_[1998]_ , \new_[1999]_ , \new_[2000]_ ,
    \new_[2001]_ , \new_[2002]_ , \new_[2003]_ , \new_[2004]_ ,
    \new_[2005]_ , \new_[2006]_ , \new_[2007]_ , \new_[2008]_ ,
    \new_[2009]_ , \new_[2010]_ , \new_[2011]_ , \new_[2012]_ ,
    \new_[2013]_ , \new_[2014]_ , \new_[2015]_ , \new_[2016]_ ,
    \new_[2017]_ , \new_[2018]_ , \new_[2019]_ , \new_[2020]_ ,
    \new_[2021]_ , \new_[2022]_ , \new_[2023]_ , \new_[2024]_ ,
    \new_[2025]_ , \new_[2026]_ , \new_[2027]_ , \new_[2028]_ ,
    \new_[2029]_ , \new_[2030]_ , \new_[2031]_ , \new_[2032]_ ,
    \new_[2033]_ , \new_[2034]_ , \new_[2035]_ , \new_[2036]_ ,
    \new_[2037]_ , \new_[2038]_ , \new_[2039]_ , \new_[2040]_ ,
    \new_[2041]_ , \new_[2042]_ , \new_[2043]_ , \new_[2044]_ ,
    \new_[2045]_ , \new_[2046]_ , \new_[2047]_ , \new_[2048]_ ,
    \new_[2049]_ , \new_[2050]_ , \new_[2051]_ , \new_[2052]_ ,
    \new_[2053]_ , \new_[2054]_ , \new_[2055]_ , \new_[2056]_ ,
    \new_[2057]_ , \new_[2058]_ , \new_[2059]_ , \new_[2060]_ ,
    \new_[2061]_ , \new_[2062]_ , \new_[2063]_ , \new_[2064]_ ,
    \new_[2065]_ , \new_[2066]_ , \new_[2067]_ , \new_[2068]_ ,
    \new_[2069]_ , \new_[2070]_ , \new_[2071]_ , \new_[2072]_ ,
    \new_[2073]_ , \new_[2074]_ , \new_[2075]_ , \new_[2076]_ ,
    \new_[2077]_ , \new_[2078]_ , \new_[2079]_ , \new_[2080]_ ,
    \new_[2081]_ , \new_[2082]_ , \new_[2083]_ , \new_[2084]_ ,
    \new_[2085]_ , \new_[2086]_ , \new_[2087]_ , \new_[2088]_ ,
    \new_[2089]_ , \new_[2090]_ , \new_[2091]_ , \new_[2092]_ ,
    \new_[2093]_ , \new_[2094]_ , \new_[2095]_ , \new_[2096]_ ,
    \new_[2097]_ , \new_[2098]_ , \new_[2099]_ , \new_[2100]_ ,
    \new_[2101]_ , \new_[2102]_ , \new_[2103]_ , \new_[2104]_ ,
    \new_[2105]_ , \new_[2106]_ , \new_[2107]_ , \new_[2108]_ ,
    \new_[2109]_ , \new_[2110]_ , \new_[2111]_ , \new_[2112]_ ,
    \new_[2113]_ , \new_[2114]_ , \new_[2115]_ , \new_[2116]_ ,
    \new_[2117]_ , \new_[2118]_ , \new_[2119]_ , \new_[2120]_ ,
    \new_[2121]_ , \new_[2122]_ , \new_[2123]_ , \new_[2124]_ ,
    \new_[2125]_ , \new_[2126]_ , \new_[2127]_ , \new_[2128]_ ,
    \new_[2129]_ , \new_[2130]_ , \new_[2131]_ , \new_[2132]_ ,
    \new_[2133]_ , \new_[2134]_ , \new_[2135]_ , \new_[2136]_ ,
    \new_[2137]_ , \new_[2138]_ , \new_[2139]_ , \new_[2140]_ ,
    \new_[2141]_ , \new_[2142]_ , \new_[2143]_ , \new_[2144]_ ,
    \new_[2145]_ , \new_[2146]_ , \new_[2147]_ , \new_[2148]_ ,
    \new_[2149]_ , \new_[2150]_ , \new_[2151]_ , \new_[2152]_ ,
    \new_[2153]_ , \new_[2154]_ , \new_[2155]_ , \new_[2156]_ ,
    \new_[2157]_ , \new_[2158]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2162]_ , \new_[2163]_ , \new_[2164]_ ,
    \new_[2165]_ , \new_[2166]_ , \new_[2167]_ , \new_[2168]_ ,
    \new_[2169]_ , \new_[2170]_ , \new_[2171]_ , \new_[2172]_ ,
    \new_[2173]_ , \new_[2174]_ , \new_[2175]_ , \new_[2176]_ ,
    \new_[2177]_ , \new_[2178]_ , \new_[2179]_ , \new_[2180]_ ,
    \new_[2181]_ , \new_[2182]_ , \new_[2183]_ , \new_[2184]_ ,
    \new_[2185]_ , \new_[2186]_ , \new_[2187]_ , \new_[2188]_ ,
    \new_[2189]_ , \new_[2190]_ , \new_[2191]_ , \new_[2192]_ ,
    \new_[2193]_ , \new_[2194]_ , \new_[2195]_ , \new_[2196]_ ,
    \new_[2197]_ , \new_[2198]_ , \new_[2199]_ , \new_[2200]_ ,
    \new_[2201]_ , \new_[2202]_ , \new_[2203]_ , \new_[2204]_ ,
    \new_[2205]_ , \new_[2206]_ , \new_[2207]_ , \new_[2208]_ ,
    \new_[2209]_ , \new_[2210]_ , \new_[2211]_ , \new_[2212]_ ,
    \new_[2213]_ , \new_[2214]_ , \new_[2215]_ , \new_[2216]_ ,
    \new_[2217]_ , \new_[2218]_ , \new_[2219]_ , \new_[2220]_ ,
    \new_[2221]_ , \new_[2222]_ , \new_[2223]_ , \new_[2224]_ ,
    \new_[2225]_ , \new_[2226]_ , \new_[2227]_ , \new_[2228]_ ,
    \new_[2229]_ , \new_[2230]_ , \new_[2231]_ , \new_[2232]_ ,
    \new_[2233]_ , \new_[2234]_ , \new_[2235]_ , \new_[2236]_ ,
    \new_[2237]_ , \new_[2238]_ , \new_[2239]_ , \new_[2240]_ ,
    \new_[2241]_ , \new_[2242]_ , \new_[2243]_ , \new_[2244]_ ,
    \new_[2245]_ , \new_[2246]_ , \new_[2247]_ , \new_[2248]_ ,
    \new_[2249]_ , \new_[2250]_ , \new_[2251]_ , \new_[2252]_ ,
    \new_[2253]_ , \new_[2254]_ , \new_[2255]_ , \new_[2256]_ ,
    \new_[2257]_ , \new_[2258]_ , \new_[2259]_ , \new_[2260]_ ,
    \new_[2261]_ , \new_[2262]_ , \new_[2263]_ , \new_[2264]_ ,
    \new_[2265]_ , \new_[2266]_ , \new_[2267]_ , \new_[2268]_ ,
    \new_[2269]_ , \new_[2270]_ , \new_[2271]_ , \new_[2272]_ ,
    \new_[2273]_ , \new_[2274]_ , \new_[2275]_ , \new_[2276]_ ,
    \new_[2277]_ , \new_[2278]_ , \new_[2279]_ , \new_[2280]_ ,
    \new_[2281]_ , \new_[2282]_ , \new_[2283]_ , \new_[2284]_ ,
    \new_[2285]_ , \new_[2286]_ , \new_[2287]_ , \new_[2288]_ ,
    \new_[2289]_ , \new_[2290]_ , \new_[2291]_ , \new_[2292]_ ,
    \new_[2293]_ , \new_[2294]_ , \new_[2295]_ , \new_[2296]_ ,
    \new_[2297]_ , \new_[2298]_ , \new_[2299]_ , \new_[2300]_ ,
    \new_[2301]_ , \new_[2302]_ , \new_[2303]_ , \new_[2304]_ ,
    \new_[2305]_ , \new_[2306]_ , \new_[2307]_ , \new_[2308]_ ,
    \new_[2309]_ , \new_[2310]_ , \new_[2311]_ , \new_[2312]_ ,
    \new_[2313]_ , \new_[2314]_ , \new_[2315]_ , \new_[2316]_ ,
    \new_[2317]_ , \new_[2318]_ , \new_[2319]_ , \new_[2320]_ ,
    \new_[2321]_ , \new_[2322]_ , \new_[2323]_ , \new_[2324]_ ,
    \new_[2325]_ , \new_[2326]_ , \new_[2327]_ , \new_[2328]_ ,
    \new_[2329]_ , \new_[2330]_ , \new_[2331]_ , \new_[2332]_ ,
    \new_[2333]_ , \new_[2334]_ , \new_[2335]_ , \new_[2336]_ ,
    \new_[2337]_ , \new_[2338]_ , \new_[2339]_ , \new_[2340]_ ,
    \new_[2341]_ , \new_[2342]_ , \new_[2343]_ , \new_[2344]_ ,
    \new_[2345]_ , \new_[2346]_ , \new_[2347]_ , \new_[2348]_ ,
    \new_[2349]_ , \new_[2350]_ , \new_[2351]_ , \new_[2352]_ ,
    \new_[2353]_ , \new_[2354]_ , \new_[2355]_ , \new_[2356]_ ,
    \new_[2357]_ , \new_[2358]_ , \new_[2359]_ , \new_[2360]_ ,
    \new_[2361]_ , \new_[2362]_ , \new_[2363]_ , \new_[2364]_ ,
    \new_[2365]_ , \new_[2366]_ , \new_[2367]_ , \new_[2368]_ ,
    \new_[2369]_ , \new_[2370]_ , \new_[2371]_ , \new_[2372]_ ,
    \new_[2373]_ , \new_[2374]_ , \new_[2375]_ , \new_[2376]_ ,
    \new_[2377]_ , \new_[2378]_ , \new_[2379]_ , \new_[2380]_ ,
    \new_[2381]_ , \new_[2382]_ , \new_[2383]_ , \new_[2384]_ ,
    \new_[2385]_ , \new_[2386]_ , \new_[2387]_ , \new_[2388]_ ,
    \new_[2389]_ , \new_[2390]_ , \new_[2391]_ , \new_[2392]_ ,
    \new_[2393]_ , \new_[2394]_ , \new_[2395]_ , \new_[2396]_ ,
    \new_[2397]_ , \new_[2398]_ , \new_[2399]_ , \new_[2400]_ ,
    \new_[2401]_ , \new_[2402]_ , \new_[2403]_ , \new_[2404]_ ,
    \new_[2405]_ , \new_[2406]_ , \new_[2407]_ , \new_[2408]_ ,
    \new_[2409]_ , \new_[2410]_ , \new_[2411]_ , \new_[2412]_ ,
    \new_[2413]_ , \new_[2414]_ , \new_[2415]_ , \new_[2416]_ ,
    \new_[2417]_ , \new_[2418]_ , \new_[2419]_ , \new_[2420]_ ,
    \new_[2421]_ , \new_[2422]_ , \new_[2423]_ , \new_[2424]_ ,
    \new_[2425]_ , \new_[2426]_ , \new_[2427]_ , \new_[2428]_ ,
    \new_[2429]_ , \new_[2430]_ , \new_[2431]_ , \new_[2432]_ ,
    \new_[2433]_ , \new_[2434]_ , \new_[2435]_ , \new_[2436]_ ,
    \new_[2437]_ , \new_[2438]_ , \new_[2439]_ , \new_[2440]_ ,
    \new_[2441]_ , \new_[2442]_ , \new_[2443]_ , \new_[2444]_ ,
    \new_[2445]_ , \new_[2446]_ , \new_[2447]_ , \new_[2448]_ ,
    \new_[2449]_ , \new_[2450]_ , \new_[2451]_ , \new_[2452]_ ,
    \new_[2453]_ , \new_[2454]_ , \new_[2455]_ , \new_[2456]_ ,
    \new_[2457]_ , \new_[2458]_ , \new_[2459]_ , \new_[2460]_ ,
    \new_[2461]_ , \new_[2462]_ , \new_[2463]_ , \new_[2464]_ ,
    \new_[2465]_ , \new_[2466]_ , \new_[2467]_ , \new_[2468]_ ,
    \new_[2469]_ , \new_[2470]_ , \new_[2471]_ , \new_[2472]_ ,
    \new_[2473]_ , \new_[2474]_ , \new_[2475]_ , \new_[2476]_ ,
    \new_[2477]_ , \new_[2478]_ , \new_[2479]_ , \new_[2480]_ ,
    \new_[2481]_ , \new_[2482]_ , \new_[2483]_ , \new_[2484]_ ,
    \new_[2485]_ , \new_[2486]_ , \new_[2487]_ , \new_[2488]_ ,
    \new_[2489]_ , \new_[2490]_ , \new_[2491]_ , \new_[2492]_ ,
    \new_[2493]_ , \new_[2494]_ , \new_[2495]_ , \new_[2496]_ ,
    \new_[2497]_ , \new_[2498]_ , \new_[2499]_ , \new_[2500]_ ,
    \new_[2501]_ , \new_[2502]_ , \new_[2503]_ , \new_[2504]_ ,
    \new_[2505]_ , \new_[2506]_ , \new_[2507]_ , \new_[2508]_ ,
    \new_[2509]_ , \new_[2510]_ , \new_[2511]_ , \new_[2512]_ ,
    \new_[2513]_ , \new_[2514]_ , \new_[2515]_ , \new_[2516]_ ,
    \new_[2517]_ , \new_[2518]_ , \new_[2519]_ , \new_[2520]_ ,
    \new_[2521]_ , \new_[2522]_ , \new_[2523]_ , \new_[2524]_ ,
    \new_[2525]_ , \new_[2526]_ , \new_[2527]_ , \new_[2528]_ ,
    \new_[2529]_ , \new_[2530]_ , \new_[2531]_ , \new_[2532]_ ,
    \new_[2533]_ , \new_[2534]_ , \new_[2535]_ , \new_[2536]_ ,
    \new_[2537]_ , \new_[2538]_ , \new_[2539]_ , \new_[2540]_ ,
    \new_[2541]_ , \new_[2542]_ , \new_[2543]_ , \new_[2544]_ ,
    \new_[2545]_ , \new_[2546]_ , \new_[2547]_ , \new_[2548]_ ,
    \new_[2549]_ , \new_[2550]_ , \new_[2551]_ , \new_[2552]_ ,
    \new_[2553]_ , \new_[2554]_ , \new_[2555]_ , \new_[2556]_ ,
    \new_[2557]_ , \new_[2558]_ , \new_[2559]_ , \new_[2560]_ ,
    \new_[2561]_ , \new_[2562]_ , \new_[2563]_ , \new_[2564]_ ,
    \new_[2565]_ , \new_[2566]_ , \new_[2567]_ , \new_[2568]_ ,
    \new_[2569]_ , \new_[2570]_ , \new_[2571]_ , \new_[2572]_ ,
    \new_[2573]_ , \new_[2574]_ , \new_[2575]_ , \new_[2576]_ ,
    \new_[2577]_ , \new_[2578]_ , \new_[2579]_ , \new_[2580]_ ,
    \new_[2581]_ , \new_[2582]_ , \new_[2583]_ , \new_[2584]_ ,
    \new_[2585]_ , \new_[2586]_ , \new_[2587]_ , \new_[2588]_ ,
    \new_[2589]_ , \new_[2590]_ , \new_[2591]_ , \new_[2592]_ ,
    \new_[2593]_ , \new_[2594]_ , \new_[2595]_ , \new_[2596]_ ,
    \new_[2597]_ , \new_[2598]_ , \new_[2599]_ , \new_[2600]_ ,
    \new_[2601]_ , \new_[2602]_ , \new_[2603]_ , \new_[2604]_ ,
    \new_[2605]_ , \new_[2606]_ , \new_[2607]_ , \new_[2608]_ ,
    \new_[2609]_ , \new_[2610]_ , \new_[2611]_ , \new_[2612]_ ,
    \new_[2613]_ , \new_[2614]_ , \new_[2615]_ , \new_[2616]_ ,
    \new_[2617]_ , \new_[2618]_ , \new_[2619]_ , \new_[2620]_ ,
    \new_[2621]_ , \new_[2622]_ , \new_[2623]_ , \new_[2624]_ ,
    \new_[2625]_ , \new_[2626]_ , \new_[2627]_ , \new_[2628]_ ,
    \new_[2629]_ , \new_[2630]_ , \new_[2631]_ , \new_[2632]_ ,
    \new_[2633]_ , \new_[2634]_ , \new_[2635]_ , \new_[2636]_ ,
    \new_[2637]_ , \new_[2638]_ , \new_[2639]_ , \new_[2640]_ ,
    \new_[2641]_ , \new_[2642]_ , \new_[2643]_ , \new_[2644]_ ,
    \new_[2645]_ , \new_[2646]_ , \new_[2647]_ , \new_[2648]_ ,
    \new_[2649]_ , \new_[2650]_ , \new_[2651]_ , \new_[2652]_ ,
    \new_[2653]_ , \new_[2654]_ , \new_[2655]_ , \new_[2656]_ ,
    \new_[2657]_ , \new_[2658]_ , \new_[2659]_ , \new_[2660]_ ,
    \new_[2661]_ , \new_[2662]_ , \new_[2663]_ , \new_[2664]_ ,
    \new_[2665]_ , \new_[2666]_ , \new_[2667]_ , \new_[2668]_ ,
    \new_[2669]_ , \new_[2670]_ , \new_[2671]_ , \new_[2672]_ ,
    \new_[2673]_ , \new_[2674]_ , \new_[2675]_ , \new_[2676]_ ,
    \new_[2677]_ , \new_[2678]_ , \new_[2679]_ , \new_[2680]_ ,
    \new_[2681]_ , \new_[2682]_ , \new_[2683]_ , \new_[2684]_ ,
    \new_[2685]_ , \new_[2686]_ , \new_[2687]_ , \new_[2688]_ ,
    \new_[2689]_ , \new_[2690]_ , \new_[2691]_ , \new_[2692]_ ,
    \new_[2693]_ , \new_[2694]_ , \new_[2695]_ , \new_[2696]_ ,
    \new_[2697]_ , \new_[2698]_ , \new_[2699]_ , \new_[2700]_ ,
    \new_[2701]_ , \new_[2702]_ , \new_[2703]_ , \new_[2704]_ ,
    \new_[2705]_ , \new_[2706]_ , \new_[2707]_ , \new_[2708]_ ,
    \new_[2709]_ , \new_[2710]_ , \new_[2711]_ , \new_[2712]_ ,
    \new_[2713]_ , \new_[2714]_ , \new_[2715]_ , \new_[2716]_ ,
    \new_[2717]_ , \new_[2718]_ , \new_[2719]_ , \new_[2720]_ ,
    \new_[2721]_ , \new_[2722]_ , \new_[2723]_ , \new_[2724]_ ,
    \new_[2725]_ , \new_[2726]_ , \new_[2727]_ , \new_[2728]_ ,
    \new_[2729]_ , \new_[2730]_ , \new_[2731]_ , \new_[2732]_ ,
    \new_[2733]_ , \new_[2734]_ , \new_[2735]_ , \new_[2736]_ ,
    \new_[2737]_ , \new_[2738]_ , \new_[2739]_ , \new_[2740]_ ,
    \new_[2741]_ , \new_[2742]_ , \new_[2743]_ , \new_[2744]_ ,
    \new_[2745]_ , \new_[2746]_ , \new_[2747]_ , \new_[2748]_ ,
    \new_[2749]_ , \new_[2750]_ , \new_[2751]_ , \new_[2752]_ ,
    \new_[2753]_ , \new_[2754]_ , \new_[2755]_ , \new_[2756]_ ,
    \new_[2757]_ , \new_[2758]_ , \new_[2759]_ , \new_[2760]_ ,
    \new_[2761]_ , \new_[2762]_ , \new_[2763]_ , \new_[2764]_ ,
    \new_[2765]_ , \new_[2766]_ , \new_[2767]_ , \new_[2768]_ ,
    \new_[2769]_ , \new_[2770]_ , \new_[2771]_ , \new_[2772]_ ,
    \new_[2773]_ , \new_[2774]_ , \new_[2775]_ , \new_[2776]_ ,
    \new_[2777]_ , \new_[2778]_ , \new_[2779]_ , \new_[2780]_ ,
    \new_[2781]_ , \new_[2782]_ , \new_[2783]_ , \new_[2784]_ ,
    \new_[2785]_ , \new_[2786]_ , \new_[2787]_ , \new_[2788]_ ,
    \new_[2789]_ , \new_[2790]_ , \new_[2791]_ , \new_[2792]_ ,
    \new_[2793]_ , \new_[2794]_ , \new_[2795]_ , \new_[2796]_ ,
    \new_[2797]_ , \new_[2798]_ , \new_[2799]_ , \new_[2800]_ ,
    \new_[2801]_ , \new_[2802]_ , \new_[2803]_ , \new_[2804]_ ,
    \new_[2805]_ , \new_[2806]_ , \new_[2807]_ , \new_[2808]_ ,
    \new_[2809]_ , \new_[2810]_ , \new_[2811]_ , \new_[2812]_ ,
    \new_[2813]_ , \new_[2814]_ , \new_[2815]_ , \new_[2816]_ ,
    \new_[2817]_ , \new_[2818]_ , \new_[2819]_ , \new_[2820]_ ,
    \new_[2821]_ , \new_[2822]_ , \new_[2823]_ , \new_[2824]_ ,
    \new_[2825]_ , \new_[2826]_ , \new_[2827]_ , \new_[2828]_ ,
    \new_[2829]_ , \new_[2830]_ , \new_[2831]_ , \new_[2832]_ ,
    \new_[2833]_ , \new_[2834]_ , \new_[2835]_ , \new_[2836]_ ,
    \new_[2837]_ , \new_[2838]_ , \new_[2839]_ , \new_[2840]_ ,
    \new_[2841]_ , \new_[2842]_ , \new_[2843]_ , \new_[2844]_ ,
    \new_[2845]_ , \new_[2846]_ , \new_[2847]_ , \new_[2848]_ ,
    \new_[2849]_ , \new_[2850]_ , \new_[2851]_ , \new_[2852]_ ,
    \new_[2853]_ , \new_[2854]_ , \new_[2855]_ , \new_[2856]_ ,
    \new_[2857]_ , \new_[2858]_ , \new_[2859]_ , \new_[2860]_ ,
    \new_[2861]_ , \new_[2862]_ , \new_[2863]_ , \new_[2864]_ ,
    \new_[2865]_ , \new_[2866]_ , \new_[2867]_ , \new_[2868]_ ,
    \new_[2869]_ , \new_[2870]_ , \new_[2871]_ , \new_[2872]_ ,
    \new_[2873]_ , \new_[2874]_ , \new_[2875]_ , \new_[2876]_ ,
    \new_[2877]_ , \new_[2878]_ , \new_[2879]_ , \new_[2880]_ ,
    \new_[2881]_ , \new_[2882]_ , \new_[2883]_ , \new_[2884]_ ,
    \new_[2885]_ , \new_[2886]_ , \new_[2887]_ , \new_[2888]_ ,
    \new_[2889]_ , \new_[2890]_ , \new_[2891]_ , \new_[2892]_ ,
    \new_[2893]_ , \new_[2894]_ , \new_[2895]_ , \new_[2896]_ ,
    \new_[2897]_ , \new_[2898]_ , \new_[2899]_ , \new_[2900]_ ,
    \new_[2901]_ , \new_[2902]_ , \new_[2903]_ , \new_[2904]_ ,
    \new_[2905]_ , \new_[2906]_ , \new_[2907]_ , \new_[2908]_ ,
    \new_[2909]_ , \new_[2910]_ , \new_[2911]_ , \new_[2912]_ ,
    \new_[2913]_ , \new_[2914]_ , \new_[2915]_ , \new_[2916]_ ,
    \new_[2917]_ , \new_[2918]_ , \new_[2919]_ , \new_[2920]_ ,
    \new_[2921]_ , \new_[2922]_ , \new_[2923]_ , \new_[2924]_ ,
    \new_[2925]_ , \new_[2926]_ , \new_[2927]_ , \new_[2928]_ ,
    \new_[2929]_ , \new_[2930]_ , \new_[2931]_ , \new_[2932]_ ,
    \new_[2933]_ , \new_[2934]_ , \new_[2935]_ , \new_[2936]_ ,
    \new_[2937]_ , \new_[2938]_ , \new_[2939]_ , \new_[2940]_ ,
    \new_[2941]_ , \new_[2942]_ , \new_[2943]_ , \new_[2944]_ ,
    \new_[2945]_ , \new_[2946]_ , \new_[2947]_ , \new_[2948]_ ,
    \new_[2949]_ , \new_[2950]_ , \new_[2951]_ , \new_[2952]_ ,
    \new_[2953]_ , \new_[2954]_ , \new_[2955]_ , \new_[2956]_ ,
    \new_[2957]_ , \new_[2958]_ , \new_[2959]_ , \new_[2960]_ ,
    \new_[2961]_ , \new_[2962]_ , \new_[2963]_ , \new_[2964]_ ,
    \new_[2965]_ , \new_[2966]_ , \new_[2967]_ , \new_[2968]_ ,
    \new_[2969]_ , \new_[2970]_ , \new_[2971]_ , \new_[2972]_ ,
    \new_[2973]_ , \new_[2974]_ , \new_[2975]_ , \new_[2976]_ ,
    \new_[2977]_ , \new_[2978]_ , \new_[2979]_ , \new_[2980]_ ,
    \new_[2981]_ , \new_[2982]_ , \new_[2983]_ , \new_[2984]_ ,
    \new_[2985]_ , \new_[2986]_ , \new_[2987]_ , \new_[2988]_ ,
    \new_[2989]_ , \new_[2990]_ , \new_[2991]_ , \new_[2992]_ ,
    \new_[2993]_ , \new_[2994]_ , \new_[2995]_ , \new_[2996]_ ,
    \new_[2997]_ , \new_[2998]_ , \new_[2999]_ , \new_[3000]_ ,
    \new_[3001]_ , \new_[3002]_ , \new_[3003]_ , \new_[3004]_ ,
    \new_[3005]_ , \new_[3006]_ , \new_[3007]_ , \new_[3008]_ ,
    \new_[3009]_ , \new_[3010]_ , \new_[3011]_ , \new_[3012]_ ,
    \new_[3013]_ , \new_[3014]_ , \new_[3015]_ , \new_[3016]_ ,
    \new_[3017]_ , \new_[3018]_ , \new_[3019]_ , \new_[3020]_ ,
    \new_[3021]_ , \new_[3022]_ , \new_[3023]_ , \new_[3024]_ ,
    \new_[3025]_ , \new_[3026]_ , \new_[3027]_ , \new_[3028]_ ,
    \new_[3029]_ , \new_[3030]_ , \new_[3031]_ , \new_[3032]_ ,
    \new_[3033]_ , \new_[3034]_ , \new_[3035]_ , \new_[3036]_ ,
    \new_[3037]_ , \new_[3038]_ , \new_[3039]_ , \new_[3040]_ ,
    \new_[3041]_ , \new_[3042]_ , \new_[3043]_ , \new_[3044]_ ,
    \new_[3045]_ , \new_[3046]_ , \new_[3047]_ , \new_[3048]_ ,
    \new_[3049]_ , \new_[3050]_ , \new_[3051]_ , \new_[3052]_ ,
    \new_[3053]_ , \new_[3054]_ , \new_[3055]_ , \new_[3056]_ ,
    \new_[3057]_ , \new_[3058]_ , \new_[3059]_ , \new_[3060]_ ,
    \new_[3061]_ , \new_[3062]_ , \new_[3063]_ , \new_[3064]_ ,
    \new_[3065]_ , \new_[3066]_ , \new_[3067]_ , \new_[3068]_ ,
    \new_[3069]_ , \new_[3070]_ , \new_[3071]_ , \new_[3072]_ ,
    \new_[3073]_ , \new_[3074]_ , \new_[3075]_ , \new_[3076]_ ,
    \new_[3077]_ , \new_[3078]_ , \new_[3079]_ , \new_[3080]_ ,
    \new_[3081]_ , \new_[3082]_ , \new_[3083]_ , \new_[3084]_ ,
    \new_[3085]_ , \new_[3086]_ , \new_[3087]_ , \new_[3088]_ ,
    \new_[3089]_ , \new_[3090]_ , \new_[3091]_ , \new_[3092]_ ,
    \new_[3093]_ , \new_[3094]_ , \new_[3095]_ , \new_[3096]_ ,
    \new_[3097]_ , \new_[3098]_ , \new_[3099]_ , \new_[3100]_ ,
    \new_[3101]_ , \new_[3102]_ , \new_[3103]_ , \new_[3104]_ ,
    \new_[3105]_ , \new_[3106]_ , \new_[3107]_ , \new_[3108]_ ,
    \new_[3109]_ , \new_[3110]_ , \new_[3111]_ , \new_[3112]_ ,
    \new_[3113]_ , \new_[3114]_ , \new_[3115]_ , \new_[3116]_ ,
    \new_[3117]_ , \new_[3118]_ , \new_[3119]_ , \new_[3120]_ ,
    \new_[3121]_ , \new_[3122]_ , \new_[3123]_ , \new_[3124]_ ,
    \new_[3125]_ , \new_[3126]_ , \new_[3127]_ , \new_[3128]_ ,
    \new_[3129]_ , \new_[3130]_ , \new_[3131]_ , \new_[3132]_ ,
    \new_[3133]_ , \new_[3134]_ , \new_[3135]_ , \new_[3136]_ ,
    \new_[3137]_ , \new_[3138]_ , \new_[3139]_ , \new_[3140]_ ,
    \new_[3141]_ , \new_[3142]_ , \new_[3143]_ , \new_[3144]_ ,
    \new_[3145]_ , \new_[3146]_ , \new_[3147]_ , \new_[3148]_ ,
    \new_[3149]_ , \new_[3150]_ , \new_[3151]_ , \new_[3152]_ ,
    \new_[3153]_ , \new_[3154]_ , \new_[3155]_ , \new_[3156]_ ,
    \new_[3157]_ , \new_[3158]_ , \new_[3159]_ , \new_[3160]_ ,
    \new_[3161]_ , \new_[3162]_ , \new_[3163]_ , \new_[3164]_ ,
    \new_[3165]_ , \new_[3166]_ , \new_[3167]_ , \new_[3168]_ ,
    \new_[3169]_ , \new_[3170]_ , \new_[3171]_ , \new_[3172]_ ,
    \new_[3173]_ , \new_[3174]_ , \new_[3175]_ , \new_[3176]_ ,
    \new_[3177]_ , \new_[3178]_ , \new_[3179]_ , \new_[3180]_ ,
    \new_[3181]_ , \new_[3182]_ , \new_[3183]_ , \new_[3184]_ ,
    \new_[3185]_ , \new_[3186]_ , \new_[3187]_ , \new_[3188]_ ,
    \new_[3189]_ , \new_[3190]_ , \new_[3191]_ , \new_[3192]_ ,
    \new_[3193]_ , \new_[3194]_ , \new_[3195]_ , \new_[3196]_ ,
    \new_[3197]_ , \new_[3198]_ , \new_[3199]_ , \new_[3200]_ ,
    \new_[3201]_ , \new_[3202]_ , \new_[3203]_ , \new_[3204]_ ,
    \new_[3205]_ , \new_[3206]_ , \new_[3207]_ , \new_[3208]_ ,
    \new_[3209]_ , \new_[3210]_ , \new_[3211]_ , \new_[3212]_ ,
    \new_[3213]_ , \new_[3214]_ , \new_[3215]_ , \new_[3216]_ ,
    \new_[3217]_ , \new_[3218]_ , \new_[3219]_ , \new_[3220]_ ,
    \new_[3221]_ , \new_[3222]_ , \new_[3223]_ , \new_[3224]_ ,
    \new_[3225]_ , \new_[3226]_ , \new_[3227]_ , \new_[3228]_ ,
    \new_[3229]_ , \new_[3230]_ , \new_[3231]_ , \new_[3232]_ ,
    \new_[3233]_ , \new_[3234]_ , \new_[3235]_ , \new_[3236]_ ,
    \new_[3237]_ , \new_[3238]_ , \new_[3239]_ , \new_[3240]_ ,
    \new_[3241]_ , \new_[3242]_ , \new_[3243]_ , \new_[3244]_ ,
    \new_[3245]_ , \new_[3246]_ , \new_[3247]_ , \new_[3248]_ ,
    \new_[3249]_ , \new_[3250]_ , \new_[3251]_ , \new_[3252]_ ,
    \new_[3253]_ , \new_[3254]_ , \new_[3255]_ , \new_[3256]_ ,
    \new_[3257]_ , \new_[3258]_ , \new_[3259]_ , \new_[3260]_ ,
    \new_[3261]_ , \new_[3262]_ , \new_[3263]_ , \new_[3264]_ ,
    \new_[3265]_ , \new_[3266]_ , \new_[3267]_ , \new_[3268]_ ,
    \new_[3269]_ , \new_[3270]_ , \new_[3271]_ , \new_[3272]_ ,
    \new_[3273]_ , \new_[3274]_ , \new_[3275]_ , \new_[3276]_ ,
    \new_[3277]_ , \new_[3278]_ , \new_[3279]_ , \new_[3280]_ ,
    \new_[3281]_ , \new_[3282]_ , \new_[3283]_ , \new_[3284]_ ,
    \new_[3285]_ , \new_[3286]_ , \new_[3287]_ , \new_[3288]_ ,
    \new_[3289]_ , \new_[3290]_ , \new_[3291]_ , \new_[3292]_ ,
    \new_[3293]_ , \new_[3294]_ , \new_[3295]_ , \new_[3296]_ ,
    \new_[3297]_ , \new_[3298]_ , \new_[3299]_ , \new_[3300]_ ,
    \new_[3301]_ , \new_[3302]_ , \new_[3303]_ , \new_[3304]_ ,
    \new_[3305]_ , \new_[3306]_ , \new_[3307]_ , \new_[3308]_ ,
    \new_[3309]_ , \new_[3310]_ , \new_[3311]_ , \new_[3312]_ ,
    \new_[3313]_ , \new_[3314]_ , \new_[3315]_ , \new_[3316]_ ,
    \new_[3317]_ , \new_[3318]_ , \new_[3319]_ , \new_[3320]_ ,
    \new_[3321]_ , \new_[3322]_ , \new_[3323]_ , \new_[3324]_ ,
    \new_[3325]_ , \new_[3326]_ , \new_[3327]_ , \new_[3328]_ ,
    \new_[3329]_ , \new_[3330]_ , \new_[3331]_ , \new_[3332]_ ,
    \new_[3333]_ , \new_[3334]_ , \new_[3335]_ , \new_[3336]_ ,
    \new_[3337]_ , \new_[3338]_ , \new_[3339]_ , \new_[3340]_ ,
    \new_[3341]_ , \new_[3342]_ , \new_[3343]_ , \new_[3344]_ ,
    \new_[3345]_ , \new_[3346]_ , \new_[3347]_ , \new_[3348]_ ,
    \new_[3349]_ , \new_[3350]_ , \new_[3351]_ , \new_[3352]_ ,
    \new_[3353]_ , \new_[3354]_ , \new_[3355]_ , \new_[3356]_ ,
    \new_[3357]_ , \new_[3358]_ , \new_[3359]_ , \new_[3360]_ ,
    \new_[3361]_ , \new_[3362]_ , \new_[3363]_ , \new_[3364]_ ,
    \new_[3365]_ , \new_[3366]_ , \new_[3367]_ , \new_[3368]_ ,
    \new_[3369]_ , \new_[3370]_ , \new_[3371]_ , \new_[3372]_ ,
    \new_[3373]_ , \new_[3374]_ , \new_[3375]_ , \new_[3376]_ ,
    \new_[3377]_ , \new_[3378]_ , \new_[3379]_ , \new_[3380]_ ,
    \new_[3381]_ , \new_[3382]_ , \new_[3383]_ , \new_[3384]_ ,
    \new_[3385]_ , \new_[3386]_ , \new_[3387]_ , \new_[3388]_ ,
    \new_[3389]_ , \new_[3390]_ , \new_[3391]_ , \new_[3392]_ ,
    \new_[3393]_ , \new_[3394]_ , \new_[3395]_ , \new_[3396]_ ,
    \new_[3397]_ , \new_[3398]_ , \new_[3399]_ , \new_[3400]_ ,
    \new_[3401]_ , \new_[3402]_ , \new_[3403]_ , \new_[3404]_ ,
    \new_[3405]_ , \new_[3406]_ , \new_[3407]_ , \new_[3408]_ ,
    \new_[3409]_ , \new_[3410]_ , \new_[3411]_ , \new_[3412]_ ,
    \new_[3413]_ , \new_[3414]_ , \new_[3415]_ , \new_[3416]_ ,
    \new_[3417]_ , \new_[3418]_ , \new_[3419]_ , \new_[3420]_ ,
    \new_[3421]_ , \new_[3422]_ , \new_[3423]_ , \new_[3424]_ ,
    \new_[3425]_ , \new_[3426]_ , \new_[3427]_ , \new_[3428]_ ,
    \new_[3429]_ , \new_[3430]_ , \new_[3431]_ , \new_[3432]_ ,
    \new_[3433]_ , \new_[3434]_ , \new_[3435]_ , \new_[3436]_ ,
    \new_[3437]_ , \new_[3438]_ , \new_[3439]_ , \new_[3440]_ ,
    \new_[3441]_ , \new_[3442]_ , \new_[3443]_ , \new_[3444]_ ,
    \new_[3445]_ , \new_[3446]_ , \new_[3447]_ , \new_[3448]_ ,
    \new_[3449]_ , \new_[3450]_ , \new_[3451]_ , \new_[3452]_ ,
    \new_[3453]_ , \new_[3454]_ , \new_[3455]_ , \new_[3456]_ ,
    \new_[3457]_ , \new_[3458]_ , \new_[3459]_ , \new_[3460]_ ,
    \new_[3461]_ , \new_[3462]_ , \new_[3463]_ , \new_[3464]_ ,
    \new_[3465]_ , \new_[3466]_ , \new_[3467]_ , \new_[3468]_ ,
    \new_[3469]_ , \new_[3470]_ , \new_[3471]_ , \new_[3472]_ ,
    \new_[3473]_ , \new_[3474]_ , \new_[3475]_ , \new_[3476]_ ,
    \new_[3477]_ , \new_[3478]_ , \new_[3479]_ , \new_[3480]_ ,
    \new_[3481]_ , \new_[3482]_ , \new_[3483]_ , \new_[3484]_ ,
    \new_[3485]_ , \new_[3486]_ , \new_[3487]_ , \new_[3488]_ ,
    \new_[3489]_ , \new_[3490]_ , \new_[3491]_ , \new_[3492]_ ,
    \new_[3493]_ , \new_[3494]_ , \new_[3495]_ , \new_[3496]_ ,
    \new_[3497]_ , \new_[3498]_ , \new_[3499]_ , \new_[3500]_ ,
    \new_[3501]_ , \new_[3502]_ , \new_[3503]_ , \new_[3504]_ ,
    \new_[3505]_ , \new_[3506]_ , \new_[3507]_ , \new_[3508]_ ,
    \new_[3509]_ , \new_[3510]_ , \new_[3511]_ , \new_[3512]_ ,
    \new_[3513]_ , \new_[3514]_ , \new_[3515]_ , \new_[3516]_ ,
    \new_[3517]_ , \new_[3518]_ , \new_[3519]_ , \new_[3520]_ ,
    \new_[3521]_ , \new_[3522]_ , \new_[3523]_ , \new_[3524]_ ,
    \new_[3525]_ , \new_[3526]_ , \new_[3527]_ , \new_[3528]_ ,
    \new_[3529]_ , \new_[3530]_ , \new_[3531]_ , \new_[3532]_ ,
    \new_[3533]_ , \new_[3534]_ , \new_[3535]_ , \new_[3536]_ ,
    \new_[3537]_ , \new_[3538]_ , \new_[3539]_ , \new_[3540]_ ,
    \new_[3541]_ , \new_[3542]_ , \new_[3543]_ , \new_[3544]_ ,
    \new_[3545]_ , \new_[3546]_ , \new_[3547]_ , \new_[3548]_ ,
    \new_[3549]_ , \new_[3550]_ , \new_[3551]_ , \new_[3552]_ ,
    \new_[3553]_ , \new_[3554]_ , \new_[3555]_ , \new_[3556]_ ,
    \new_[3557]_ , \new_[3558]_ , \new_[3559]_ , \new_[3560]_ ,
    \new_[3561]_ , \new_[3562]_ , \new_[3563]_ , \new_[3564]_ ,
    \new_[3565]_ , \new_[3566]_ , \new_[3567]_ , \new_[3568]_ ,
    \new_[3569]_ , \new_[3570]_ , \new_[3571]_ , \new_[3572]_ ,
    \new_[3573]_ , \new_[3574]_ , \new_[3575]_ , \new_[3576]_ ,
    \new_[3577]_ , \new_[3578]_ , \new_[3579]_ , \new_[3580]_ ,
    \new_[3581]_ , \new_[3582]_ , \new_[3583]_ , \new_[3584]_ ,
    \new_[3585]_ , \new_[3586]_ , \new_[3587]_ , \new_[3588]_ ,
    \new_[3589]_ , \new_[3590]_ , \new_[3591]_ , \new_[3592]_ ,
    \new_[3593]_ , \new_[3594]_ , \new_[3595]_ , \new_[3596]_ ,
    \new_[3597]_ , \new_[3598]_ , \new_[3599]_ , \new_[3600]_ ,
    \new_[3601]_ , \new_[3602]_ , \new_[3603]_ , \new_[3604]_ ,
    \new_[3605]_ , \new_[3606]_ , \new_[3607]_ , \new_[3608]_ ,
    \new_[3609]_ , \new_[3610]_ , \new_[3611]_ , \new_[3612]_ ,
    \new_[3613]_ , \new_[3614]_ , \new_[3615]_ , \new_[3616]_ ,
    \new_[3617]_ , \new_[3618]_ , \new_[3619]_ , \new_[3620]_ ,
    \new_[3621]_ , \new_[3622]_ , \new_[3623]_ , \new_[3624]_ ,
    \new_[3625]_ , \new_[3626]_ , \new_[3627]_ , \new_[3628]_ ,
    \new_[3629]_ , \new_[3630]_ , \new_[3631]_ , \new_[3632]_ ,
    \new_[3633]_ , \new_[3634]_ , \new_[3635]_ , \new_[3636]_ ,
    \new_[3637]_ , \new_[3638]_ , \new_[3639]_ , \new_[3640]_ ,
    \new_[3641]_ , \new_[3642]_ , \new_[3643]_ , \new_[3644]_ ,
    \new_[3645]_ , \new_[3646]_ , \new_[3647]_ , \new_[3648]_ ,
    \new_[3649]_ , \new_[3650]_ , \new_[3651]_ , \new_[3652]_ ,
    \new_[3653]_ , \new_[3654]_ , \new_[3655]_ , \new_[3656]_ ,
    \new_[3657]_ , \new_[3658]_ , \new_[3659]_ , \new_[3660]_ ,
    \new_[3661]_ , \new_[3662]_ , \new_[3663]_ , \new_[3664]_ ,
    \new_[3665]_ , \new_[3666]_ , \new_[3667]_ , \new_[3668]_ ,
    \new_[3669]_ , \new_[3670]_ , \new_[3671]_ , \new_[3672]_ ,
    \new_[3673]_ , \new_[3674]_ , \new_[3675]_ , \new_[3676]_ ,
    \new_[3677]_ , \new_[3678]_ , \new_[3679]_ , \new_[3680]_ ,
    \new_[3681]_ , \new_[3682]_ , \new_[3683]_ , \new_[3684]_ ,
    \new_[3685]_ , \new_[3686]_ , \new_[3687]_ , \new_[3688]_ ,
    \new_[3689]_ , \new_[3690]_ , \new_[3691]_ , \new_[3692]_ ,
    \new_[3693]_ , \new_[3694]_ , \new_[3695]_ , \new_[3696]_ ,
    \new_[3697]_ , \new_[3698]_ , \new_[3699]_ , \new_[3700]_ ,
    \new_[3701]_ , \new_[3702]_ , \new_[3703]_ , \new_[3704]_ ,
    \new_[3705]_ , \new_[3706]_ , \new_[3707]_ , \new_[3708]_ ,
    \new_[3709]_ , \new_[3710]_ , \new_[3711]_ , \new_[3712]_ ,
    \new_[3713]_ , \new_[3714]_ , \new_[3715]_ , \new_[3716]_ ,
    \new_[3717]_ , \new_[3718]_ , \new_[3719]_ , \new_[3720]_ ,
    \new_[3721]_ , \new_[3722]_ , \new_[3723]_ , \new_[3724]_ ,
    \new_[3725]_ , \new_[3726]_ , \new_[3727]_ , \new_[3728]_ ,
    \new_[3729]_ , \new_[3730]_ , \new_[3731]_ , \new_[3732]_ ,
    \new_[3733]_ , \new_[3734]_ , \new_[3735]_ , \new_[3736]_ ,
    \new_[3737]_ , \new_[3738]_ , \new_[3739]_ , \new_[3740]_ ,
    \new_[3741]_ , \new_[3742]_ , \new_[3743]_ , \new_[3744]_ ,
    \new_[3745]_ , \new_[3746]_ , \new_[3747]_ , \new_[3748]_ ,
    \new_[3749]_ , \new_[3750]_ , \new_[3751]_ , \new_[3752]_ ,
    \new_[3753]_ , \new_[3754]_ , \new_[3755]_ , \new_[3756]_ ,
    \new_[3757]_ , \new_[3758]_ , \new_[3759]_ , \new_[3760]_ ,
    \new_[3761]_ , \new_[3762]_ , \new_[3763]_ , \new_[3764]_ ,
    \new_[3765]_ , \new_[3766]_ , \new_[3767]_ , \new_[3768]_ ,
    \new_[3769]_ , \new_[3770]_ , \new_[3771]_ , \new_[3772]_ ,
    \new_[3776]_ , \new_[3777]_ , \new_[3780]_ , \new_[3783]_ ,
    \new_[3784]_ , \new_[3785]_ , \new_[3789]_ , \new_[3790]_ ,
    \new_[3793]_ , \new_[3796]_ , \new_[3797]_ , \new_[3798]_ ,
    \new_[3799]_ , \new_[3803]_ , \new_[3804]_ , \new_[3807]_ ,
    \new_[3810]_ , \new_[3811]_ , \new_[3812]_ , \new_[3815]_ ,
    \new_[3818]_ , \new_[3819]_ , \new_[3822]_ , \new_[3825]_ ,
    \new_[3826]_ , \new_[3827]_ , \new_[3828]_ , \new_[3829]_ ,
    \new_[3833]_ , \new_[3834]_ , \new_[3837]_ , \new_[3840]_ ,
    \new_[3841]_ , \new_[3842]_ , \new_[3846]_ , \new_[3847]_ ,
    \new_[3850]_ , \new_[3853]_ , \new_[3854]_ , \new_[3855]_ ,
    \new_[3856]_ , \new_[3860]_ , \new_[3861]_ , \new_[3864]_ ,
    \new_[3867]_ , \new_[3868]_ , \new_[3869]_ , \new_[3872]_ ,
    \new_[3875]_ , \new_[3876]_ , \new_[3879]_ , \new_[3882]_ ,
    \new_[3883]_ , \new_[3884]_ , \new_[3885]_ , \new_[3886]_ ,
    \new_[3887]_ , \new_[3891]_ , \new_[3892]_ , \new_[3895]_ ,
    \new_[3898]_ , \new_[3899]_ , \new_[3900]_ , \new_[3904]_ ,
    \new_[3905]_ , \new_[3908]_ , \new_[3911]_ , \new_[3912]_ ,
    \new_[3913]_ , \new_[3914]_ , \new_[3918]_ , \new_[3919]_ ,
    \new_[3922]_ , \new_[3925]_ , \new_[3926]_ , \new_[3927]_ ,
    \new_[3930]_ , \new_[3933]_ , \new_[3934]_ , \new_[3937]_ ,
    \new_[3940]_ , \new_[3941]_ , \new_[3942]_ , \new_[3943]_ ,
    \new_[3944]_ , \new_[3948]_ , \new_[3949]_ , \new_[3952]_ ,
    \new_[3955]_ , \new_[3956]_ , \new_[3957]_ , \new_[3960]_ ,
    \new_[3963]_ , \new_[3964]_ , \new_[3967]_ , \new_[3970]_ ,
    \new_[3971]_ , \new_[3972]_ , \new_[3973]_ , \new_[3977]_ ,
    \new_[3978]_ , \new_[3981]_ , \new_[3984]_ , \new_[3985]_ ,
    \new_[3986]_ , \new_[3989]_ , \new_[3992]_ , \new_[3993]_ ,
    \new_[3996]_ , \new_[3999]_ , \new_[4000]_ , \new_[4001]_ ,
    \new_[4002]_ , \new_[4003]_ , \new_[4004]_ , \new_[4005]_ ,
    \new_[4009]_ , \new_[4010]_ , \new_[4013]_ , \new_[4016]_ ,
    \new_[4017]_ , \new_[4018]_ , \new_[4022]_ , \new_[4023]_ ,
    \new_[4026]_ , \new_[4029]_ , \new_[4030]_ , \new_[4031]_ ,
    \new_[4032]_ , \new_[4036]_ , \new_[4037]_ , \new_[4040]_ ,
    \new_[4043]_ , \new_[4044]_ , \new_[4045]_ , \new_[4048]_ ,
    \new_[4051]_ , \new_[4052]_ , \new_[4055]_ , \new_[4058]_ ,
    \new_[4059]_ , \new_[4060]_ , \new_[4061]_ , \new_[4062]_ ,
    \new_[4066]_ , \new_[4067]_ , \new_[4070]_ , \new_[4073]_ ,
    \new_[4074]_ , \new_[4075]_ , \new_[4078]_ , \new_[4081]_ ,
    \new_[4082]_ , \new_[4085]_ , \new_[4088]_ , \new_[4089]_ ,
    \new_[4090]_ , \new_[4091]_ , \new_[4095]_ , \new_[4096]_ ,
    \new_[4099]_ , \new_[4102]_ , \new_[4103]_ , \new_[4104]_ ,
    \new_[4107]_ , \new_[4110]_ , \new_[4111]_ , \new_[4114]_ ,
    \new_[4117]_ , \new_[4118]_ , \new_[4119]_ , \new_[4120]_ ,
    \new_[4121]_ , \new_[4122]_ , \new_[4126]_ , \new_[4127]_ ,
    \new_[4130]_ , \new_[4133]_ , \new_[4134]_ , \new_[4135]_ ,
    \new_[4139]_ , \new_[4140]_ , \new_[4143]_ , \new_[4146]_ ,
    \new_[4147]_ , \new_[4148]_ , \new_[4149]_ , \new_[4153]_ ,
    \new_[4154]_ , \new_[4157]_ , \new_[4160]_ , \new_[4161]_ ,
    \new_[4162]_ , \new_[4165]_ , \new_[4168]_ , \new_[4169]_ ,
    \new_[4172]_ , \new_[4175]_ , \new_[4176]_ , \new_[4177]_ ,
    \new_[4178]_ , \new_[4179]_ , \new_[4183]_ , \new_[4184]_ ,
    \new_[4187]_ , \new_[4190]_ , \new_[4191]_ , \new_[4192]_ ,
    \new_[4195]_ , \new_[4198]_ , \new_[4199]_ , \new_[4202]_ ,
    \new_[4205]_ , \new_[4206]_ , \new_[4207]_ , \new_[4208]_ ,
    \new_[4212]_ , \new_[4213]_ , \new_[4216]_ , \new_[4219]_ ,
    \new_[4220]_ , \new_[4221]_ , \new_[4224]_ , \new_[4227]_ ,
    \new_[4228]_ , \new_[4231]_ , \new_[4234]_ , \new_[4235]_ ,
    \new_[4236]_ , \new_[4237]_ , \new_[4238]_ , \new_[4239]_ ,
    \new_[4240]_ , \new_[4241]_ , \new_[4245]_ , \new_[4246]_ ,
    \new_[4249]_ , \new_[4252]_ , \new_[4253]_ , \new_[4254]_ ,
    \new_[4258]_ , \new_[4259]_ , \new_[4262]_ , \new_[4265]_ ,
    \new_[4266]_ , \new_[4267]_ , \new_[4268]_ , \new_[4272]_ ,
    \new_[4273]_ , \new_[4276]_ , \new_[4279]_ , \new_[4280]_ ,
    \new_[4281]_ , \new_[4284]_ , \new_[4287]_ , \new_[4288]_ ,
    \new_[4291]_ , \new_[4294]_ , \new_[4295]_ , \new_[4296]_ ,
    \new_[4297]_ , \new_[4298]_ , \new_[4302]_ , \new_[4303]_ ,
    \new_[4306]_ , \new_[4309]_ , \new_[4310]_ , \new_[4311]_ ,
    \new_[4314]_ , \new_[4317]_ , \new_[4318]_ , \new_[4321]_ ,
    \new_[4324]_ , \new_[4325]_ , \new_[4326]_ , \new_[4327]_ ,
    \new_[4331]_ , \new_[4332]_ , \new_[4335]_ , \new_[4338]_ ,
    \new_[4339]_ , \new_[4340]_ , \new_[4343]_ , \new_[4346]_ ,
    \new_[4347]_ , \new_[4350]_ , \new_[4353]_ , \new_[4354]_ ,
    \new_[4355]_ , \new_[4356]_ , \new_[4357]_ , \new_[4358]_ ,
    \new_[4362]_ , \new_[4363]_ , \new_[4366]_ , \new_[4369]_ ,
    \new_[4370]_ , \new_[4371]_ , \new_[4375]_ , \new_[4376]_ ,
    \new_[4379]_ , \new_[4382]_ , \new_[4383]_ , \new_[4384]_ ,
    \new_[4385]_ , \new_[4389]_ , \new_[4390]_ , \new_[4393]_ ,
    \new_[4396]_ , \new_[4397]_ , \new_[4398]_ , \new_[4401]_ ,
    \new_[4404]_ , \new_[4405]_ , \new_[4408]_ , \new_[4411]_ ,
    \new_[4412]_ , \new_[4413]_ , \new_[4414]_ , \new_[4415]_ ,
    \new_[4419]_ , \new_[4420]_ , \new_[4423]_ , \new_[4426]_ ,
    \new_[4427]_ , \new_[4428]_ , \new_[4431]_ , \new_[4434]_ ,
    \new_[4435]_ , \new_[4438]_ , \new_[4441]_ , \new_[4442]_ ,
    \new_[4443]_ , \new_[4444]_ , \new_[4448]_ , \new_[4449]_ ,
    \new_[4452]_ , \new_[4455]_ , \new_[4456]_ , \new_[4457]_ ,
    \new_[4460]_ , \new_[4463]_ , \new_[4464]_ , \new_[4467]_ ,
    \new_[4470]_ , \new_[4471]_ , \new_[4472]_ , \new_[4473]_ ,
    \new_[4474]_ , \new_[4475]_ , \new_[4476]_ , \new_[4480]_ ,
    \new_[4481]_ , \new_[4484]_ , \new_[4487]_ , \new_[4488]_ ,
    \new_[4489]_ , \new_[4493]_ , \new_[4494]_ , \new_[4497]_ ,
    \new_[4500]_ , \new_[4501]_ , \new_[4502]_ , \new_[4503]_ ,
    \new_[4507]_ , \new_[4508]_ , \new_[4511]_ , \new_[4514]_ ,
    \new_[4515]_ , \new_[4516]_ , \new_[4519]_ , \new_[4522]_ ,
    \new_[4523]_ , \new_[4526]_ , \new_[4529]_ , \new_[4530]_ ,
    \new_[4531]_ , \new_[4532]_ , \new_[4533]_ , \new_[4537]_ ,
    \new_[4538]_ , \new_[4541]_ , \new_[4544]_ , \new_[4545]_ ,
    \new_[4546]_ , \new_[4549]_ , \new_[4552]_ , \new_[4553]_ ,
    \new_[4556]_ , \new_[4559]_ , \new_[4560]_ , \new_[4561]_ ,
    \new_[4562]_ , \new_[4566]_ , \new_[4567]_ , \new_[4570]_ ,
    \new_[4573]_ , \new_[4574]_ , \new_[4575]_ , \new_[4578]_ ,
    \new_[4581]_ , \new_[4582]_ , \new_[4585]_ , \new_[4588]_ ,
    \new_[4589]_ , \new_[4590]_ , \new_[4591]_ , \new_[4592]_ ,
    \new_[4593]_ , \new_[4597]_ , \new_[4598]_ , \new_[4601]_ ,
    \new_[4604]_ , \new_[4605]_ , \new_[4606]_ , \new_[4610]_ ,
    \new_[4611]_ , \new_[4614]_ , \new_[4617]_ , \new_[4618]_ ,
    \new_[4619]_ , \new_[4620]_ , \new_[4624]_ , \new_[4625]_ ,
    \new_[4628]_ , \new_[4631]_ , \new_[4632]_ , \new_[4633]_ ,
    \new_[4636]_ , \new_[4639]_ , \new_[4640]_ , \new_[4643]_ ,
    \new_[4646]_ , \new_[4647]_ , \new_[4648]_ , \new_[4649]_ ,
    \new_[4650]_ , \new_[4654]_ , \new_[4655]_ , \new_[4658]_ ,
    \new_[4661]_ , \new_[4662]_ , \new_[4663]_ , \new_[4666]_ ,
    \new_[4669]_ , \new_[4670]_ , \new_[4673]_ , \new_[4676]_ ,
    \new_[4677]_ , \new_[4678]_ , \new_[4679]_ , \new_[4683]_ ,
    \new_[4684]_ , \new_[4687]_ , \new_[4690]_ , \new_[4691]_ ,
    \new_[4692]_ , \new_[4695]_ , \new_[4698]_ , \new_[4699]_ ,
    \new_[4702]_ , \new_[4705]_ , \new_[4706]_ , \new_[4707]_ ,
    \new_[4708]_ , \new_[4709]_ , \new_[4710]_ , \new_[4711]_ ,
    \new_[4712]_ , \new_[4713]_ , \new_[4717]_ , \new_[4718]_ ,
    \new_[4721]_ , \new_[4724]_ , \new_[4725]_ , \new_[4726]_ ,
    \new_[4730]_ , \new_[4731]_ , \new_[4734]_ , \new_[4737]_ ,
    \new_[4738]_ , \new_[4739]_ , \new_[4740]_ , \new_[4744]_ ,
    \new_[4745]_ , \new_[4748]_ , \new_[4751]_ , \new_[4752]_ ,
    \new_[4753]_ , \new_[4756]_ , \new_[4759]_ , \new_[4760]_ ,
    \new_[4763]_ , \new_[4766]_ , \new_[4767]_ , \new_[4768]_ ,
    \new_[4769]_ , \new_[4770]_ , \new_[4774]_ , \new_[4775]_ ,
    \new_[4778]_ , \new_[4781]_ , \new_[4782]_ , \new_[4783]_ ,
    \new_[4786]_ , \new_[4789]_ , \new_[4790]_ , \new_[4793]_ ,
    \new_[4796]_ , \new_[4797]_ , \new_[4798]_ , \new_[4799]_ ,
    \new_[4803]_ , \new_[4804]_ , \new_[4807]_ , \new_[4810]_ ,
    \new_[4811]_ , \new_[4812]_ , \new_[4815]_ , \new_[4818]_ ,
    \new_[4819]_ , \new_[4822]_ , \new_[4825]_ , \new_[4826]_ ,
    \new_[4827]_ , \new_[4828]_ , \new_[4829]_ , \new_[4830]_ ,
    \new_[4834]_ , \new_[4835]_ , \new_[4838]_ , \new_[4841]_ ,
    \new_[4842]_ , \new_[4843]_ , \new_[4847]_ , \new_[4848]_ ,
    \new_[4851]_ , \new_[4854]_ , \new_[4855]_ , \new_[4856]_ ,
    \new_[4857]_ , \new_[4861]_ , \new_[4862]_ , \new_[4865]_ ,
    \new_[4868]_ , \new_[4869]_ , \new_[4870]_ , \new_[4873]_ ,
    \new_[4876]_ , \new_[4877]_ , \new_[4880]_ , \new_[4883]_ ,
    \new_[4884]_ , \new_[4885]_ , \new_[4886]_ , \new_[4887]_ ,
    \new_[4891]_ , \new_[4892]_ , \new_[4895]_ , \new_[4898]_ ,
    \new_[4899]_ , \new_[4900]_ , \new_[4903]_ , \new_[4906]_ ,
    \new_[4907]_ , \new_[4910]_ , \new_[4913]_ , \new_[4914]_ ,
    \new_[4915]_ , \new_[4916]_ , \new_[4920]_ , \new_[4921]_ ,
    \new_[4924]_ , \new_[4927]_ , \new_[4928]_ , \new_[4929]_ ,
    \new_[4932]_ , \new_[4935]_ , \new_[4936]_ , \new_[4939]_ ,
    \new_[4942]_ , \new_[4943]_ , \new_[4944]_ , \new_[4945]_ ,
    \new_[4946]_ , \new_[4947]_ , \new_[4948]_ , \new_[4952]_ ,
    \new_[4953]_ , \new_[4956]_ , \new_[4959]_ , \new_[4960]_ ,
    \new_[4961]_ , \new_[4965]_ , \new_[4966]_ , \new_[4969]_ ,
    \new_[4972]_ , \new_[4973]_ , \new_[4974]_ , \new_[4975]_ ,
    \new_[4979]_ , \new_[4980]_ , \new_[4983]_ , \new_[4986]_ ,
    \new_[4987]_ , \new_[4988]_ , \new_[4991]_ , \new_[4994]_ ,
    \new_[4995]_ , \new_[4998]_ , \new_[5001]_ , \new_[5002]_ ,
    \new_[5003]_ , \new_[5004]_ , \new_[5005]_ , \new_[5009]_ ,
    \new_[5010]_ , \new_[5013]_ , \new_[5016]_ , \new_[5017]_ ,
    \new_[5018]_ , \new_[5021]_ , \new_[5024]_ , \new_[5025]_ ,
    \new_[5028]_ , \new_[5031]_ , \new_[5032]_ , \new_[5033]_ ,
    \new_[5034]_ , \new_[5038]_ , \new_[5039]_ , \new_[5042]_ ,
    \new_[5045]_ , \new_[5046]_ , \new_[5047]_ , \new_[5050]_ ,
    \new_[5053]_ , \new_[5054]_ , \new_[5057]_ , \new_[5060]_ ,
    \new_[5061]_ , \new_[5062]_ , \new_[5063]_ , \new_[5064]_ ,
    \new_[5065]_ , \new_[5069]_ , \new_[5070]_ , \new_[5073]_ ,
    \new_[5076]_ , \new_[5077]_ , \new_[5078]_ , \new_[5082]_ ,
    \new_[5083]_ , \new_[5086]_ , \new_[5089]_ , \new_[5090]_ ,
    \new_[5091]_ , \new_[5092]_ , \new_[5096]_ , \new_[5097]_ ,
    \new_[5100]_ , \new_[5103]_ , \new_[5104]_ , \new_[5105]_ ,
    \new_[5108]_ , \new_[5111]_ , \new_[5112]_ , \new_[5115]_ ,
    \new_[5118]_ , \new_[5119]_ , \new_[5120]_ , \new_[5121]_ ,
    \new_[5122]_ , \new_[5126]_ , \new_[5127]_ , \new_[5130]_ ,
    \new_[5133]_ , \new_[5134]_ , \new_[5135]_ , \new_[5138]_ ,
    \new_[5141]_ , \new_[5142]_ , \new_[5145]_ , \new_[5148]_ ,
    \new_[5149]_ , \new_[5150]_ , \new_[5151]_ , \new_[5155]_ ,
    \new_[5156]_ , \new_[5159]_ , \new_[5162]_ , \new_[5163]_ ,
    \new_[5164]_ , \new_[5167]_ , \new_[5170]_ , \new_[5171]_ ,
    \new_[5174]_ , \new_[5177]_ , \new_[5178]_ , \new_[5179]_ ,
    \new_[5180]_ , \new_[5181]_ , \new_[5182]_ , \new_[5183]_ ,
    \new_[5184]_ , \new_[5188]_ , \new_[5189]_ , \new_[5192]_ ,
    \new_[5195]_ , \new_[5196]_ , \new_[5197]_ , \new_[5201]_ ,
    \new_[5202]_ , \new_[5205]_ , \new_[5208]_ , \new_[5209]_ ,
    \new_[5210]_ , \new_[5211]_ , \new_[5215]_ , \new_[5216]_ ,
    \new_[5219]_ , \new_[5222]_ , \new_[5223]_ , \new_[5224]_ ,
    \new_[5227]_ , \new_[5230]_ , \new_[5231]_ , \new_[5234]_ ,
    \new_[5237]_ , \new_[5238]_ , \new_[5239]_ , \new_[5240]_ ,
    \new_[5241]_ , \new_[5245]_ , \new_[5246]_ , \new_[5249]_ ,
    \new_[5252]_ , \new_[5253]_ , \new_[5254]_ , \new_[5257]_ ,
    \new_[5260]_ , \new_[5261]_ , \new_[5264]_ , \new_[5267]_ ,
    \new_[5268]_ , \new_[5269]_ , \new_[5270]_ , \new_[5274]_ ,
    \new_[5275]_ , \new_[5278]_ , \new_[5281]_ , \new_[5282]_ ,
    \new_[5283]_ , \new_[5286]_ , \new_[5289]_ , \new_[5290]_ ,
    \new_[5293]_ , \new_[5296]_ , \new_[5297]_ , \new_[5298]_ ,
    \new_[5299]_ , \new_[5300]_ , \new_[5301]_ , \new_[5305]_ ,
    \new_[5306]_ , \new_[5309]_ , \new_[5312]_ , \new_[5313]_ ,
    \new_[5314]_ , \new_[5318]_ , \new_[5319]_ , \new_[5322]_ ,
    \new_[5325]_ , \new_[5326]_ , \new_[5327]_ , \new_[5328]_ ,
    \new_[5332]_ , \new_[5333]_ , \new_[5336]_ , \new_[5339]_ ,
    \new_[5340]_ , \new_[5341]_ , \new_[5344]_ , \new_[5347]_ ,
    \new_[5348]_ , \new_[5351]_ , \new_[5354]_ , \new_[5355]_ ,
    \new_[5356]_ , \new_[5357]_ , \new_[5358]_ , \new_[5362]_ ,
    \new_[5363]_ , \new_[5366]_ , \new_[5369]_ , \new_[5370]_ ,
    \new_[5371]_ , \new_[5374]_ , \new_[5377]_ , \new_[5378]_ ,
    \new_[5381]_ , \new_[5384]_ , \new_[5385]_ , \new_[5386]_ ,
    \new_[5387]_ , \new_[5391]_ , \new_[5392]_ , \new_[5395]_ ,
    \new_[5398]_ , \new_[5399]_ , \new_[5400]_ , \new_[5403]_ ,
    \new_[5406]_ , \new_[5407]_ , \new_[5410]_ , \new_[5413]_ ,
    \new_[5414]_ , \new_[5415]_ , \new_[5416]_ , \new_[5417]_ ,
    \new_[5418]_ , \new_[5419]_ , \new_[5423]_ , \new_[5424]_ ,
    \new_[5427]_ , \new_[5430]_ , \new_[5431]_ , \new_[5432]_ ,
    \new_[5436]_ , \new_[5437]_ , \new_[5440]_ , \new_[5443]_ ,
    \new_[5444]_ , \new_[5445]_ , \new_[5446]_ , \new_[5450]_ ,
    \new_[5451]_ , \new_[5454]_ , \new_[5457]_ , \new_[5458]_ ,
    \new_[5459]_ , \new_[5462]_ , \new_[5465]_ , \new_[5466]_ ,
    \new_[5469]_ , \new_[5472]_ , \new_[5473]_ , \new_[5474]_ ,
    \new_[5475]_ , \new_[5476]_ , \new_[5480]_ , \new_[5481]_ ,
    \new_[5484]_ , \new_[5487]_ , \new_[5488]_ , \new_[5489]_ ,
    \new_[5492]_ , \new_[5495]_ , \new_[5496]_ , \new_[5499]_ ,
    \new_[5502]_ , \new_[5503]_ , \new_[5504]_ , \new_[5505]_ ,
    \new_[5509]_ , \new_[5510]_ , \new_[5513]_ , \new_[5516]_ ,
    \new_[5517]_ , \new_[5518]_ , \new_[5521]_ , \new_[5524]_ ,
    \new_[5525]_ , \new_[5528]_ , \new_[5531]_ , \new_[5532]_ ,
    \new_[5533]_ , \new_[5534]_ , \new_[5535]_ , \new_[5536]_ ,
    \new_[5540]_ , \new_[5541]_ , \new_[5544]_ , \new_[5547]_ ,
    \new_[5548]_ , \new_[5549]_ , \new_[5553]_ , \new_[5554]_ ,
    \new_[5557]_ , \new_[5560]_ , \new_[5561]_ , \new_[5562]_ ,
    \new_[5563]_ , \new_[5567]_ , \new_[5568]_ , \new_[5571]_ ,
    \new_[5574]_ , \new_[5575]_ , \new_[5576]_ , \new_[5579]_ ,
    \new_[5582]_ , \new_[5583]_ , \new_[5586]_ , \new_[5589]_ ,
    \new_[5590]_ , \new_[5591]_ , \new_[5592]_ , \new_[5593]_ ,
    \new_[5597]_ , \new_[5598]_ , \new_[5601]_ , \new_[5604]_ ,
    \new_[5605]_ , \new_[5606]_ , \new_[5609]_ , \new_[5612]_ ,
    \new_[5613]_ , \new_[5616]_ , \new_[5619]_ , \new_[5620]_ ,
    \new_[5621]_ , \new_[5622]_ , \new_[5626]_ , \new_[5627]_ ,
    \new_[5630]_ , \new_[5633]_ , \new_[5634]_ , \new_[5635]_ ,
    \new_[5638]_ , \new_[5641]_ , \new_[5642]_ , \new_[5645]_ ,
    \new_[5648]_ , \new_[5649]_ , \new_[5650]_ , \new_[5651]_ ,
    \new_[5652]_ , \new_[5653]_ , \new_[5654]_ , \new_[5655]_ ,
    \new_[5656]_ , \new_[5657]_ , \new_[5661]_ , \new_[5662]_ ,
    \new_[5665]_ , \new_[5668]_ , \new_[5669]_ , \new_[5670]_ ,
    \new_[5674]_ , \new_[5675]_ , \new_[5678]_ , \new_[5681]_ ,
    \new_[5682]_ , \new_[5683]_ , \new_[5684]_ , \new_[5688]_ ,
    \new_[5689]_ , \new_[5692]_ , \new_[5695]_ , \new_[5696]_ ,
    \new_[5697]_ , \new_[5700]_ , \new_[5703]_ , \new_[5704]_ ,
    \new_[5707]_ , \new_[5710]_ , \new_[5711]_ , \new_[5712]_ ,
    \new_[5713]_ , \new_[5714]_ , \new_[5718]_ , \new_[5719]_ ,
    \new_[5722]_ , \new_[5725]_ , \new_[5726]_ , \new_[5727]_ ,
    \new_[5731]_ , \new_[5732]_ , \new_[5735]_ , \new_[5738]_ ,
    \new_[5739]_ , \new_[5740]_ , \new_[5741]_ , \new_[5745]_ ,
    \new_[5746]_ , \new_[5749]_ , \new_[5752]_ , \new_[5753]_ ,
    \new_[5754]_ , \new_[5757]_ , \new_[5760]_ , \new_[5761]_ ,
    \new_[5764]_ , \new_[5767]_ , \new_[5768]_ , \new_[5769]_ ,
    \new_[5770]_ , \new_[5771]_ , \new_[5772]_ , \new_[5776]_ ,
    \new_[5777]_ , \new_[5780]_ , \new_[5783]_ , \new_[5784]_ ,
    \new_[5785]_ , \new_[5789]_ , \new_[5790]_ , \new_[5793]_ ,
    \new_[5796]_ , \new_[5797]_ , \new_[5798]_ , \new_[5799]_ ,
    \new_[5803]_ , \new_[5804]_ , \new_[5807]_ , \new_[5810]_ ,
    \new_[5811]_ , \new_[5812]_ , \new_[5815]_ , \new_[5818]_ ,
    \new_[5819]_ , \new_[5822]_ , \new_[5825]_ , \new_[5826]_ ,
    \new_[5827]_ , \new_[5828]_ , \new_[5829]_ , \new_[5833]_ ,
    \new_[5834]_ , \new_[5837]_ , \new_[5840]_ , \new_[5841]_ ,
    \new_[5842]_ , \new_[5845]_ , \new_[5848]_ , \new_[5849]_ ,
    \new_[5852]_ , \new_[5855]_ , \new_[5856]_ , \new_[5857]_ ,
    \new_[5858]_ , \new_[5862]_ , \new_[5863]_ , \new_[5866]_ ,
    \new_[5869]_ , \new_[5870]_ , \new_[5871]_ , \new_[5874]_ ,
    \new_[5877]_ , \new_[5878]_ , \new_[5881]_ , \new_[5884]_ ,
    \new_[5885]_ , \new_[5886]_ , \new_[5887]_ , \new_[5888]_ ,
    \new_[5889]_ , \new_[5890]_ , \new_[5894]_ , \new_[5895]_ ,
    \new_[5898]_ , \new_[5901]_ , \new_[5902]_ , \new_[5903]_ ,
    \new_[5907]_ , \new_[5908]_ , \new_[5911]_ , \new_[5914]_ ,
    \new_[5915]_ , \new_[5916]_ , \new_[5917]_ , \new_[5921]_ ,
    \new_[5922]_ , \new_[5925]_ , \new_[5928]_ , \new_[5929]_ ,
    \new_[5930]_ , \new_[5933]_ , \new_[5936]_ , \new_[5937]_ ,
    \new_[5940]_ , \new_[5943]_ , \new_[5944]_ , \new_[5945]_ ,
    \new_[5946]_ , \new_[5947]_ , \new_[5951]_ , \new_[5952]_ ,
    \new_[5955]_ , \new_[5958]_ , \new_[5959]_ , \new_[5960]_ ,
    \new_[5963]_ , \new_[5966]_ , \new_[5967]_ , \new_[5970]_ ,
    \new_[5973]_ , \new_[5974]_ , \new_[5975]_ , \new_[5976]_ ,
    \new_[5980]_ , \new_[5981]_ , \new_[5984]_ , \new_[5987]_ ,
    \new_[5988]_ , \new_[5989]_ , \new_[5992]_ , \new_[5995]_ ,
    \new_[5996]_ , \new_[5999]_ , \new_[6002]_ , \new_[6003]_ ,
    \new_[6004]_ , \new_[6005]_ , \new_[6006]_ , \new_[6007]_ ,
    \new_[6011]_ , \new_[6012]_ , \new_[6015]_ , \new_[6018]_ ,
    \new_[6019]_ , \new_[6020]_ , \new_[6024]_ , \new_[6025]_ ,
    \new_[6028]_ , \new_[6031]_ , \new_[6032]_ , \new_[6033]_ ,
    \new_[6034]_ , \new_[6038]_ , \new_[6039]_ , \new_[6042]_ ,
    \new_[6045]_ , \new_[6046]_ , \new_[6047]_ , \new_[6050]_ ,
    \new_[6053]_ , \new_[6054]_ , \new_[6057]_ , \new_[6060]_ ,
    \new_[6061]_ , \new_[6062]_ , \new_[6063]_ , \new_[6064]_ ,
    \new_[6068]_ , \new_[6069]_ , \new_[6072]_ , \new_[6075]_ ,
    \new_[6076]_ , \new_[6077]_ , \new_[6080]_ , \new_[6083]_ ,
    \new_[6084]_ , \new_[6087]_ , \new_[6090]_ , \new_[6091]_ ,
    \new_[6092]_ , \new_[6093]_ , \new_[6097]_ , \new_[6098]_ ,
    \new_[6101]_ , \new_[6104]_ , \new_[6105]_ , \new_[6106]_ ,
    \new_[6109]_ , \new_[6112]_ , \new_[6113]_ , \new_[6116]_ ,
    \new_[6119]_ , \new_[6120]_ , \new_[6121]_ , \new_[6122]_ ,
    \new_[6123]_ , \new_[6124]_ , \new_[6125]_ , \new_[6126]_ ,
    \new_[6130]_ , \new_[6131]_ , \new_[6134]_ , \new_[6137]_ ,
    \new_[6138]_ , \new_[6139]_ , \new_[6143]_ , \new_[6144]_ ,
    \new_[6147]_ , \new_[6150]_ , \new_[6151]_ , \new_[6152]_ ,
    \new_[6153]_ , \new_[6157]_ , \new_[6158]_ , \new_[6161]_ ,
    \new_[6164]_ , \new_[6165]_ , \new_[6166]_ , \new_[6169]_ ,
    \new_[6172]_ , \new_[6173]_ , \new_[6176]_ , \new_[6179]_ ,
    \new_[6180]_ , \new_[6181]_ , \new_[6182]_ , \new_[6183]_ ,
    \new_[6187]_ , \new_[6188]_ , \new_[6191]_ , \new_[6194]_ ,
    \new_[6195]_ , \new_[6196]_ , \new_[6199]_ , \new_[6202]_ ,
    \new_[6203]_ , \new_[6206]_ , \new_[6209]_ , \new_[6210]_ ,
    \new_[6211]_ , \new_[6212]_ , \new_[6216]_ , \new_[6217]_ ,
    \new_[6220]_ , \new_[6223]_ , \new_[6224]_ , \new_[6225]_ ,
    \new_[6228]_ , \new_[6231]_ , \new_[6232]_ , \new_[6235]_ ,
    \new_[6238]_ , \new_[6239]_ , \new_[6240]_ , \new_[6241]_ ,
    \new_[6242]_ , \new_[6243]_ , \new_[6247]_ , \new_[6248]_ ,
    \new_[6251]_ , \new_[6254]_ , \new_[6255]_ , \new_[6256]_ ,
    \new_[6260]_ , \new_[6261]_ , \new_[6264]_ , \new_[6267]_ ,
    \new_[6268]_ , \new_[6269]_ , \new_[6270]_ , \new_[6274]_ ,
    \new_[6275]_ , \new_[6278]_ , \new_[6281]_ , \new_[6282]_ ,
    \new_[6283]_ , \new_[6286]_ , \new_[6289]_ , \new_[6290]_ ,
    \new_[6293]_ , \new_[6296]_ , \new_[6297]_ , \new_[6298]_ ,
    \new_[6299]_ , \new_[6300]_ , \new_[6304]_ , \new_[6305]_ ,
    \new_[6308]_ , \new_[6311]_ , \new_[6312]_ , \new_[6313]_ ,
    \new_[6316]_ , \new_[6319]_ , \new_[6320]_ , \new_[6323]_ ,
    \new_[6326]_ , \new_[6327]_ , \new_[6328]_ , \new_[6329]_ ,
    \new_[6333]_ , \new_[6334]_ , \new_[6337]_ , \new_[6340]_ ,
    \new_[6341]_ , \new_[6342]_ , \new_[6345]_ , \new_[6348]_ ,
    \new_[6349]_ , \new_[6352]_ , \new_[6355]_ , \new_[6356]_ ,
    \new_[6357]_ , \new_[6358]_ , \new_[6359]_ , \new_[6360]_ ,
    \new_[6361]_ , \new_[6365]_ , \new_[6366]_ , \new_[6369]_ ,
    \new_[6372]_ , \new_[6373]_ , \new_[6374]_ , \new_[6378]_ ,
    \new_[6379]_ , \new_[6382]_ , \new_[6385]_ , \new_[6386]_ ,
    \new_[6387]_ , \new_[6388]_ , \new_[6392]_ , \new_[6393]_ ,
    \new_[6396]_ , \new_[6399]_ , \new_[6400]_ , \new_[6401]_ ,
    \new_[6404]_ , \new_[6407]_ , \new_[6408]_ , \new_[6411]_ ,
    \new_[6414]_ , \new_[6415]_ , \new_[6416]_ , \new_[6417]_ ,
    \new_[6418]_ , \new_[6422]_ , \new_[6423]_ , \new_[6426]_ ,
    \new_[6429]_ , \new_[6430]_ , \new_[6431]_ , \new_[6434]_ ,
    \new_[6437]_ , \new_[6438]_ , \new_[6441]_ , \new_[6444]_ ,
    \new_[6445]_ , \new_[6446]_ , \new_[6447]_ , \new_[6451]_ ,
    \new_[6452]_ , \new_[6455]_ , \new_[6458]_ , \new_[6459]_ ,
    \new_[6460]_ , \new_[6463]_ , \new_[6466]_ , \new_[6467]_ ,
    \new_[6470]_ , \new_[6473]_ , \new_[6474]_ , \new_[6475]_ ,
    \new_[6476]_ , \new_[6477]_ , \new_[6478]_ , \new_[6482]_ ,
    \new_[6483]_ , \new_[6486]_ , \new_[6489]_ , \new_[6490]_ ,
    \new_[6491]_ , \new_[6495]_ , \new_[6496]_ , \new_[6499]_ ,
    \new_[6502]_ , \new_[6503]_ , \new_[6504]_ , \new_[6505]_ ,
    \new_[6509]_ , \new_[6510]_ , \new_[6513]_ , \new_[6516]_ ,
    \new_[6517]_ , \new_[6518]_ , \new_[6521]_ , \new_[6524]_ ,
    \new_[6525]_ , \new_[6528]_ , \new_[6531]_ , \new_[6532]_ ,
    \new_[6533]_ , \new_[6534]_ , \new_[6535]_ , \new_[6539]_ ,
    \new_[6540]_ , \new_[6543]_ , \new_[6546]_ , \new_[6547]_ ,
    \new_[6548]_ , \new_[6551]_ , \new_[6554]_ , \new_[6555]_ ,
    \new_[6558]_ , \new_[6561]_ , \new_[6562]_ , \new_[6563]_ ,
    \new_[6564]_ , \new_[6568]_ , \new_[6569]_ , \new_[6572]_ ,
    \new_[6575]_ , \new_[6576]_ , \new_[6577]_ , \new_[6580]_ ,
    \new_[6583]_ , \new_[6584]_ , \new_[6587]_ , \new_[6590]_ ,
    \new_[6591]_ , \new_[6592]_ , \new_[6593]_ , \new_[6594]_ ,
    \new_[6595]_ , \new_[6596]_ , \new_[6597]_ , \new_[6598]_ ,
    \new_[6602]_ , \new_[6603]_ , \new_[6606]_ , \new_[6609]_ ,
    \new_[6610]_ , \new_[6611]_ , \new_[6615]_ , \new_[6616]_ ,
    \new_[6619]_ , \new_[6622]_ , \new_[6623]_ , \new_[6624]_ ,
    \new_[6625]_ , \new_[6629]_ , \new_[6630]_ , \new_[6633]_ ,
    \new_[6636]_ , \new_[6637]_ , \new_[6638]_ , \new_[6641]_ ,
    \new_[6644]_ , \new_[6645]_ , \new_[6648]_ , \new_[6651]_ ,
    \new_[6652]_ , \new_[6653]_ , \new_[6654]_ , \new_[6655]_ ,
    \new_[6659]_ , \new_[6660]_ , \new_[6663]_ , \new_[6666]_ ,
    \new_[6667]_ , \new_[6668]_ , \new_[6671]_ , \new_[6674]_ ,
    \new_[6675]_ , \new_[6678]_ , \new_[6681]_ , \new_[6682]_ ,
    \new_[6683]_ , \new_[6684]_ , \new_[6688]_ , \new_[6689]_ ,
    \new_[6692]_ , \new_[6695]_ , \new_[6696]_ , \new_[6697]_ ,
    \new_[6700]_ , \new_[6703]_ , \new_[6704]_ , \new_[6707]_ ,
    \new_[6710]_ , \new_[6711]_ , \new_[6712]_ , \new_[6713]_ ,
    \new_[6714]_ , \new_[6715]_ , \new_[6719]_ , \new_[6720]_ ,
    \new_[6723]_ , \new_[6726]_ , \new_[6727]_ , \new_[6728]_ ,
    \new_[6732]_ , \new_[6733]_ , \new_[6736]_ , \new_[6739]_ ,
    \new_[6740]_ , \new_[6741]_ , \new_[6742]_ , \new_[6746]_ ,
    \new_[6747]_ , \new_[6750]_ , \new_[6753]_ , \new_[6754]_ ,
    \new_[6755]_ , \new_[6758]_ , \new_[6761]_ , \new_[6762]_ ,
    \new_[6765]_ , \new_[6768]_ , \new_[6769]_ , \new_[6770]_ ,
    \new_[6771]_ , \new_[6772]_ , \new_[6776]_ , \new_[6777]_ ,
    \new_[6780]_ , \new_[6783]_ , \new_[6784]_ , \new_[6785]_ ,
    \new_[6788]_ , \new_[6791]_ , \new_[6792]_ , \new_[6795]_ ,
    \new_[6798]_ , \new_[6799]_ , \new_[6800]_ , \new_[6801]_ ,
    \new_[6805]_ , \new_[6806]_ , \new_[6809]_ , \new_[6812]_ ,
    \new_[6813]_ , \new_[6814]_ , \new_[6817]_ , \new_[6820]_ ,
    \new_[6821]_ , \new_[6824]_ , \new_[6827]_ , \new_[6828]_ ,
    \new_[6829]_ , \new_[6830]_ , \new_[6831]_ , \new_[6832]_ ,
    \new_[6833]_ , \new_[6837]_ , \new_[6838]_ , \new_[6841]_ ,
    \new_[6844]_ , \new_[6845]_ , \new_[6846]_ , \new_[6850]_ ,
    \new_[6851]_ , \new_[6854]_ , \new_[6857]_ , \new_[6858]_ ,
    \new_[6859]_ , \new_[6860]_ , \new_[6864]_ , \new_[6865]_ ,
    \new_[6868]_ , \new_[6871]_ , \new_[6872]_ , \new_[6873]_ ,
    \new_[6876]_ , \new_[6879]_ , \new_[6880]_ , \new_[6883]_ ,
    \new_[6886]_ , \new_[6887]_ , \new_[6888]_ , \new_[6889]_ ,
    \new_[6890]_ , \new_[6894]_ , \new_[6895]_ , \new_[6898]_ ,
    \new_[6901]_ , \new_[6902]_ , \new_[6903]_ , \new_[6906]_ ,
    \new_[6909]_ , \new_[6910]_ , \new_[6913]_ , \new_[6916]_ ,
    \new_[6917]_ , \new_[6918]_ , \new_[6919]_ , \new_[6923]_ ,
    \new_[6924]_ , \new_[6927]_ , \new_[6930]_ , \new_[6931]_ ,
    \new_[6932]_ , \new_[6935]_ , \new_[6938]_ , \new_[6939]_ ,
    \new_[6942]_ , \new_[6945]_ , \new_[6946]_ , \new_[6947]_ ,
    \new_[6948]_ , \new_[6949]_ , \new_[6950]_ , \new_[6954]_ ,
    \new_[6955]_ , \new_[6958]_ , \new_[6961]_ , \new_[6962]_ ,
    \new_[6963]_ , \new_[6967]_ , \new_[6968]_ , \new_[6971]_ ,
    \new_[6974]_ , \new_[6975]_ , \new_[6976]_ , \new_[6977]_ ,
    \new_[6981]_ , \new_[6982]_ , \new_[6985]_ , \new_[6988]_ ,
    \new_[6989]_ , \new_[6990]_ , \new_[6993]_ , \new_[6996]_ ,
    \new_[6997]_ , \new_[7000]_ , \new_[7003]_ , \new_[7004]_ ,
    \new_[7005]_ , \new_[7006]_ , \new_[7007]_ , \new_[7011]_ ,
    \new_[7012]_ , \new_[7015]_ , \new_[7018]_ , \new_[7019]_ ,
    \new_[7020]_ , \new_[7023]_ , \new_[7026]_ , \new_[7027]_ ,
    \new_[7030]_ , \new_[7033]_ , \new_[7034]_ , \new_[7035]_ ,
    \new_[7036]_ , \new_[7040]_ , \new_[7041]_ , \new_[7044]_ ,
    \new_[7047]_ , \new_[7048]_ , \new_[7049]_ , \new_[7052]_ ,
    \new_[7055]_ , \new_[7056]_ , \new_[7059]_ , \new_[7062]_ ,
    \new_[7063]_ , \new_[7064]_ , \new_[7065]_ , \new_[7066]_ ,
    \new_[7067]_ , \new_[7068]_ , \new_[7069]_ , \new_[7073]_ ,
    \new_[7074]_ , \new_[7077]_ , \new_[7080]_ , \new_[7081]_ ,
    \new_[7082]_ , \new_[7086]_ , \new_[7087]_ , \new_[7090]_ ,
    \new_[7093]_ , \new_[7094]_ , \new_[7095]_ , \new_[7096]_ ,
    \new_[7100]_ , \new_[7101]_ , \new_[7104]_ , \new_[7107]_ ,
    \new_[7108]_ , \new_[7109]_ , \new_[7112]_ , \new_[7115]_ ,
    \new_[7116]_ , \new_[7119]_ , \new_[7122]_ , \new_[7123]_ ,
    \new_[7124]_ , \new_[7125]_ , \new_[7126]_ , \new_[7130]_ ,
    \new_[7131]_ , \new_[7134]_ , \new_[7137]_ , \new_[7138]_ ,
    \new_[7139]_ , \new_[7142]_ , \new_[7145]_ , \new_[7146]_ ,
    \new_[7149]_ , \new_[7152]_ , \new_[7153]_ , \new_[7154]_ ,
    \new_[7155]_ , \new_[7159]_ , \new_[7160]_ , \new_[7163]_ ,
    \new_[7166]_ , \new_[7167]_ , \new_[7168]_ , \new_[7171]_ ,
    \new_[7174]_ , \new_[7175]_ , \new_[7178]_ , \new_[7181]_ ,
    \new_[7182]_ , \new_[7183]_ , \new_[7184]_ , \new_[7185]_ ,
    \new_[7186]_ , \new_[7190]_ , \new_[7191]_ , \new_[7194]_ ,
    \new_[7197]_ , \new_[7198]_ , \new_[7199]_ , \new_[7203]_ ,
    \new_[7204]_ , \new_[7207]_ , \new_[7210]_ , \new_[7211]_ ,
    \new_[7212]_ , \new_[7213]_ , \new_[7217]_ , \new_[7218]_ ,
    \new_[7221]_ , \new_[7224]_ , \new_[7225]_ , \new_[7226]_ ,
    \new_[7229]_ , \new_[7232]_ , \new_[7233]_ , \new_[7236]_ ,
    \new_[7239]_ , \new_[7240]_ , \new_[7241]_ , \new_[7242]_ ,
    \new_[7243]_ , \new_[7247]_ , \new_[7248]_ , \new_[7251]_ ,
    \new_[7254]_ , \new_[7255]_ , \new_[7256]_ , \new_[7259]_ ,
    \new_[7262]_ , \new_[7263]_ , \new_[7266]_ , \new_[7269]_ ,
    \new_[7270]_ , \new_[7271]_ , \new_[7272]_ , \new_[7276]_ ,
    \new_[7277]_ , \new_[7280]_ , \new_[7283]_ , \new_[7284]_ ,
    \new_[7285]_ , \new_[7288]_ , \new_[7291]_ , \new_[7292]_ ,
    \new_[7295]_ , \new_[7298]_ , \new_[7299]_ , \new_[7300]_ ,
    \new_[7301]_ , \new_[7302]_ , \new_[7303]_ , \new_[7304]_ ,
    \new_[7308]_ , \new_[7309]_ , \new_[7312]_ , \new_[7315]_ ,
    \new_[7316]_ , \new_[7317]_ , \new_[7321]_ , \new_[7322]_ ,
    \new_[7325]_ , \new_[7328]_ , \new_[7329]_ , \new_[7330]_ ,
    \new_[7331]_ , \new_[7335]_ , \new_[7336]_ , \new_[7339]_ ,
    \new_[7342]_ , \new_[7343]_ , \new_[7344]_ , \new_[7347]_ ,
    \new_[7350]_ , \new_[7351]_ , \new_[7354]_ , \new_[7357]_ ,
    \new_[7358]_ , \new_[7359]_ , \new_[7360]_ , \new_[7361]_ ,
    \new_[7365]_ , \new_[7366]_ , \new_[7369]_ , \new_[7372]_ ,
    \new_[7373]_ , \new_[7374]_ , \new_[7377]_ , \new_[7380]_ ,
    \new_[7381]_ , \new_[7384]_ , \new_[7387]_ , \new_[7388]_ ,
    \new_[7389]_ , \new_[7390]_ , \new_[7394]_ , \new_[7395]_ ,
    \new_[7398]_ , \new_[7401]_ , \new_[7402]_ , \new_[7403]_ ,
    \new_[7406]_ , \new_[7409]_ , \new_[7410]_ , \new_[7413]_ ,
    \new_[7416]_ , \new_[7417]_ , \new_[7418]_ , \new_[7419]_ ,
    \new_[7420]_ , \new_[7421]_ , \new_[7425]_ , \new_[7426]_ ,
    \new_[7429]_ , \new_[7432]_ , \new_[7433]_ , \new_[7434]_ ,
    \new_[7438]_ , \new_[7439]_ , \new_[7442]_ , \new_[7445]_ ,
    \new_[7446]_ , \new_[7447]_ , \new_[7448]_ , \new_[7452]_ ,
    \new_[7453]_ , \new_[7456]_ , \new_[7459]_ , \new_[7460]_ ,
    \new_[7461]_ , \new_[7464]_ , \new_[7467]_ , \new_[7468]_ ,
    \new_[7471]_ , \new_[7474]_ , \new_[7475]_ , \new_[7476]_ ,
    \new_[7477]_ , \new_[7478]_ , \new_[7482]_ , \new_[7483]_ ,
    \new_[7486]_ , \new_[7489]_ , \new_[7490]_ , \new_[7491]_ ,
    \new_[7494]_ , \new_[7497]_ , \new_[7498]_ , \new_[7501]_ ,
    \new_[7504]_ , \new_[7505]_ , \new_[7506]_ , \new_[7507]_ ,
    \new_[7511]_ , \new_[7512]_ , \new_[7515]_ , \new_[7518]_ ,
    \new_[7519]_ , \new_[7520]_ , \new_[7523]_ , \new_[7526]_ ,
    \new_[7527]_ , \new_[7530]_ , \new_[7533]_ , \new_[7534]_ ,
    \new_[7535]_ , \new_[7536]_ , \new_[7537]_ , \new_[7538]_ ,
    \new_[7539]_ , \new_[7540]_ , \new_[7541]_ , \new_[7542]_ ,
    \new_[7543]_ , \new_[7547]_ , \new_[7548]_ , \new_[7551]_ ,
    \new_[7554]_ , \new_[7555]_ , \new_[7556]_ , \new_[7560]_ ,
    \new_[7561]_ , \new_[7564]_ , \new_[7567]_ , \new_[7568]_ ,
    \new_[7569]_ , \new_[7570]_ , \new_[7574]_ , \new_[7575]_ ,
    \new_[7578]_ , \new_[7581]_ , \new_[7582]_ , \new_[7583]_ ,
    \new_[7586]_ , \new_[7589]_ , \new_[7590]_ , \new_[7593]_ ,
    \new_[7596]_ , \new_[7597]_ , \new_[7598]_ , \new_[7599]_ ,
    \new_[7600]_ , \new_[7604]_ , \new_[7605]_ , \new_[7608]_ ,
    \new_[7611]_ , \new_[7612]_ , \new_[7613]_ , \new_[7617]_ ,
    \new_[7618]_ , \new_[7621]_ , \new_[7624]_ , \new_[7625]_ ,
    \new_[7626]_ , \new_[7627]_ , \new_[7631]_ , \new_[7632]_ ,
    \new_[7635]_ , \new_[7638]_ , \new_[7639]_ , \new_[7640]_ ,
    \new_[7643]_ , \new_[7646]_ , \new_[7647]_ , \new_[7650]_ ,
    \new_[7653]_ , \new_[7654]_ , \new_[7655]_ , \new_[7656]_ ,
    \new_[7657]_ , \new_[7658]_ , \new_[7662]_ , \new_[7663]_ ,
    \new_[7666]_ , \new_[7669]_ , \new_[7670]_ , \new_[7671]_ ,
    \new_[7675]_ , \new_[7676]_ , \new_[7679]_ , \new_[7682]_ ,
    \new_[7683]_ , \new_[7684]_ , \new_[7685]_ , \new_[7689]_ ,
    \new_[7690]_ , \new_[7693]_ , \new_[7696]_ , \new_[7697]_ ,
    \new_[7698]_ , \new_[7701]_ , \new_[7704]_ , \new_[7705]_ ,
    \new_[7708]_ , \new_[7711]_ , \new_[7712]_ , \new_[7713]_ ,
    \new_[7714]_ , \new_[7715]_ , \new_[7719]_ , \new_[7720]_ ,
    \new_[7723]_ , \new_[7726]_ , \new_[7727]_ , \new_[7728]_ ,
    \new_[7731]_ , \new_[7734]_ , \new_[7735]_ , \new_[7738]_ ,
    \new_[7741]_ , \new_[7742]_ , \new_[7743]_ , \new_[7744]_ ,
    \new_[7748]_ , \new_[7749]_ , \new_[7752]_ , \new_[7755]_ ,
    \new_[7756]_ , \new_[7757]_ , \new_[7760]_ , \new_[7763]_ ,
    \new_[7764]_ , \new_[7767]_ , \new_[7770]_ , \new_[7771]_ ,
    \new_[7772]_ , \new_[7773]_ , \new_[7774]_ , \new_[7775]_ ,
    \new_[7776]_ , \new_[7780]_ , \new_[7781]_ , \new_[7784]_ ,
    \new_[7787]_ , \new_[7788]_ , \new_[7789]_ , \new_[7793]_ ,
    \new_[7794]_ , \new_[7797]_ , \new_[7800]_ , \new_[7801]_ ,
    \new_[7802]_ , \new_[7803]_ , \new_[7807]_ , \new_[7808]_ ,
    \new_[7811]_ , \new_[7814]_ , \new_[7815]_ , \new_[7816]_ ,
    \new_[7819]_ , \new_[7822]_ , \new_[7823]_ , \new_[7826]_ ,
    \new_[7829]_ , \new_[7830]_ , \new_[7831]_ , \new_[7832]_ ,
    \new_[7833]_ , \new_[7837]_ , \new_[7838]_ , \new_[7841]_ ,
    \new_[7844]_ , \new_[7845]_ , \new_[7846]_ , \new_[7849]_ ,
    \new_[7852]_ , \new_[7853]_ , \new_[7856]_ , \new_[7859]_ ,
    \new_[7860]_ , \new_[7861]_ , \new_[7862]_ , \new_[7866]_ ,
    \new_[7867]_ , \new_[7870]_ , \new_[7873]_ , \new_[7874]_ ,
    \new_[7875]_ , \new_[7878]_ , \new_[7881]_ , \new_[7882]_ ,
    \new_[7885]_ , \new_[7888]_ , \new_[7889]_ , \new_[7890]_ ,
    \new_[7891]_ , \new_[7892]_ , \new_[7893]_ , \new_[7897]_ ,
    \new_[7898]_ , \new_[7901]_ , \new_[7904]_ , \new_[7905]_ ,
    \new_[7906]_ , \new_[7910]_ , \new_[7911]_ , \new_[7914]_ ,
    \new_[7917]_ , \new_[7918]_ , \new_[7919]_ , \new_[7920]_ ,
    \new_[7924]_ , \new_[7925]_ , \new_[7928]_ , \new_[7931]_ ,
    \new_[7932]_ , \new_[7933]_ , \new_[7936]_ , \new_[7939]_ ,
    \new_[7940]_ , \new_[7943]_ , \new_[7946]_ , \new_[7947]_ ,
    \new_[7948]_ , \new_[7949]_ , \new_[7950]_ , \new_[7954]_ ,
    \new_[7955]_ , \new_[7958]_ , \new_[7961]_ , \new_[7962]_ ,
    \new_[7963]_ , \new_[7966]_ , \new_[7969]_ , \new_[7970]_ ,
    \new_[7973]_ , \new_[7976]_ , \new_[7977]_ , \new_[7978]_ ,
    \new_[7979]_ , \new_[7983]_ , \new_[7984]_ , \new_[7987]_ ,
    \new_[7990]_ , \new_[7991]_ , \new_[7992]_ , \new_[7995]_ ,
    \new_[7998]_ , \new_[7999]_ , \new_[8002]_ , \new_[8005]_ ,
    \new_[8006]_ , \new_[8007]_ , \new_[8008]_ , \new_[8009]_ ,
    \new_[8010]_ , \new_[8011]_ , \new_[8012]_ , \new_[8016]_ ,
    \new_[8017]_ , \new_[8020]_ , \new_[8023]_ , \new_[8024]_ ,
    \new_[8025]_ , \new_[8029]_ , \new_[8030]_ , \new_[8033]_ ,
    \new_[8036]_ , \new_[8037]_ , \new_[8038]_ , \new_[8039]_ ,
    \new_[8043]_ , \new_[8044]_ , \new_[8047]_ , \new_[8050]_ ,
    \new_[8051]_ , \new_[8052]_ , \new_[8055]_ , \new_[8058]_ ,
    \new_[8059]_ , \new_[8062]_ , \new_[8065]_ , \new_[8066]_ ,
    \new_[8067]_ , \new_[8068]_ , \new_[8069]_ , \new_[8073]_ ,
    \new_[8074]_ , \new_[8077]_ , \new_[8080]_ , \new_[8081]_ ,
    \new_[8082]_ , \new_[8085]_ , \new_[8088]_ , \new_[8089]_ ,
    \new_[8092]_ , \new_[8095]_ , \new_[8096]_ , \new_[8097]_ ,
    \new_[8098]_ , \new_[8102]_ , \new_[8103]_ , \new_[8106]_ ,
    \new_[8109]_ , \new_[8110]_ , \new_[8111]_ , \new_[8114]_ ,
    \new_[8117]_ , \new_[8118]_ , \new_[8121]_ , \new_[8124]_ ,
    \new_[8125]_ , \new_[8126]_ , \new_[8127]_ , \new_[8128]_ ,
    \new_[8129]_ , \new_[8133]_ , \new_[8134]_ , \new_[8137]_ ,
    \new_[8140]_ , \new_[8141]_ , \new_[8142]_ , \new_[8146]_ ,
    \new_[8147]_ , \new_[8150]_ , \new_[8153]_ , \new_[8154]_ ,
    \new_[8155]_ , \new_[8156]_ , \new_[8160]_ , \new_[8161]_ ,
    \new_[8164]_ , \new_[8167]_ , \new_[8168]_ , \new_[8169]_ ,
    \new_[8172]_ , \new_[8175]_ , \new_[8176]_ , \new_[8179]_ ,
    \new_[8182]_ , \new_[8183]_ , \new_[8184]_ , \new_[8185]_ ,
    \new_[8186]_ , \new_[8190]_ , \new_[8191]_ , \new_[8194]_ ,
    \new_[8197]_ , \new_[8198]_ , \new_[8199]_ , \new_[8202]_ ,
    \new_[8205]_ , \new_[8206]_ , \new_[8209]_ , \new_[8212]_ ,
    \new_[8213]_ , \new_[8214]_ , \new_[8215]_ , \new_[8219]_ ,
    \new_[8220]_ , \new_[8223]_ , \new_[8226]_ , \new_[8227]_ ,
    \new_[8228]_ , \new_[8231]_ , \new_[8234]_ , \new_[8235]_ ,
    \new_[8238]_ , \new_[8241]_ , \new_[8242]_ , \new_[8243]_ ,
    \new_[8244]_ , \new_[8245]_ , \new_[8246]_ , \new_[8247]_ ,
    \new_[8251]_ , \new_[8252]_ , \new_[8255]_ , \new_[8258]_ ,
    \new_[8259]_ , \new_[8260]_ , \new_[8264]_ , \new_[8265]_ ,
    \new_[8268]_ , \new_[8271]_ , \new_[8272]_ , \new_[8273]_ ,
    \new_[8274]_ , \new_[8278]_ , \new_[8279]_ , \new_[8282]_ ,
    \new_[8285]_ , \new_[8286]_ , \new_[8287]_ , \new_[8290]_ ,
    \new_[8293]_ , \new_[8294]_ , \new_[8297]_ , \new_[8300]_ ,
    \new_[8301]_ , \new_[8302]_ , \new_[8303]_ , \new_[8304]_ ,
    \new_[8308]_ , \new_[8309]_ , \new_[8312]_ , \new_[8315]_ ,
    \new_[8316]_ , \new_[8317]_ , \new_[8320]_ , \new_[8323]_ ,
    \new_[8324]_ , \new_[8327]_ , \new_[8330]_ , \new_[8331]_ ,
    \new_[8332]_ , \new_[8333]_ , \new_[8337]_ , \new_[8338]_ ,
    \new_[8341]_ , \new_[8344]_ , \new_[8345]_ , \new_[8346]_ ,
    \new_[8349]_ , \new_[8352]_ , \new_[8353]_ , \new_[8356]_ ,
    \new_[8359]_ , \new_[8360]_ , \new_[8361]_ , \new_[8362]_ ,
    \new_[8363]_ , \new_[8364]_ , \new_[8368]_ , \new_[8369]_ ,
    \new_[8372]_ , \new_[8375]_ , \new_[8376]_ , \new_[8377]_ ,
    \new_[8381]_ , \new_[8382]_ , \new_[8385]_ , \new_[8388]_ ,
    \new_[8389]_ , \new_[8390]_ , \new_[8391]_ , \new_[8395]_ ,
    \new_[8396]_ , \new_[8399]_ , \new_[8402]_ , \new_[8403]_ ,
    \new_[8404]_ , \new_[8407]_ , \new_[8410]_ , \new_[8411]_ ,
    \new_[8414]_ , \new_[8417]_ , \new_[8418]_ , \new_[8419]_ ,
    \new_[8420]_ , \new_[8421]_ , \new_[8425]_ , \new_[8426]_ ,
    \new_[8429]_ , \new_[8432]_ , \new_[8433]_ , \new_[8434]_ ,
    \new_[8437]_ , \new_[8440]_ , \new_[8441]_ , \new_[8444]_ ,
    \new_[8447]_ , \new_[8448]_ , \new_[8449]_ , \new_[8450]_ ,
    \new_[8454]_ , \new_[8455]_ , \new_[8458]_ , \new_[8461]_ ,
    \new_[8462]_ , \new_[8463]_ , \new_[8466]_ , \new_[8469]_ ,
    \new_[8470]_ , \new_[8473]_ , \new_[8476]_ , \new_[8477]_ ,
    \new_[8478]_ , \new_[8479]_ , \new_[8480]_ , \new_[8481]_ ,
    \new_[8482]_ , \new_[8483]_ , \new_[8484]_ , \new_[8488]_ ,
    \new_[8489]_ , \new_[8492]_ , \new_[8495]_ , \new_[8496]_ ,
    \new_[8497]_ , \new_[8501]_ , \new_[8502]_ , \new_[8505]_ ,
    \new_[8508]_ , \new_[8509]_ , \new_[8510]_ , \new_[8511]_ ,
    \new_[8515]_ , \new_[8516]_ , \new_[8519]_ , \new_[8522]_ ,
    \new_[8523]_ , \new_[8524]_ , \new_[8527]_ , \new_[8530]_ ,
    \new_[8531]_ , \new_[8534]_ , \new_[8537]_ , \new_[8538]_ ,
    \new_[8539]_ , \new_[8540]_ , \new_[8541]_ , \new_[8545]_ ,
    \new_[8546]_ , \new_[8549]_ , \new_[8552]_ , \new_[8553]_ ,
    \new_[8554]_ , \new_[8557]_ , \new_[8560]_ , \new_[8561]_ ,
    \new_[8564]_ , \new_[8567]_ , \new_[8568]_ , \new_[8569]_ ,
    \new_[8570]_ , \new_[8574]_ , \new_[8575]_ , \new_[8578]_ ,
    \new_[8581]_ , \new_[8582]_ , \new_[8583]_ , \new_[8586]_ ,
    \new_[8589]_ , \new_[8590]_ , \new_[8593]_ , \new_[8596]_ ,
    \new_[8597]_ , \new_[8598]_ , \new_[8599]_ , \new_[8600]_ ,
    \new_[8601]_ , \new_[8605]_ , \new_[8606]_ , \new_[8609]_ ,
    \new_[8612]_ , \new_[8613]_ , \new_[8614]_ , \new_[8618]_ ,
    \new_[8619]_ , \new_[8622]_ , \new_[8625]_ , \new_[8626]_ ,
    \new_[8627]_ , \new_[8628]_ , \new_[8632]_ , \new_[8633]_ ,
    \new_[8636]_ , \new_[8639]_ , \new_[8640]_ , \new_[8641]_ ,
    \new_[8644]_ , \new_[8647]_ , \new_[8648]_ , \new_[8651]_ ,
    \new_[8654]_ , \new_[8655]_ , \new_[8656]_ , \new_[8657]_ ,
    \new_[8658]_ , \new_[8662]_ , \new_[8663]_ , \new_[8666]_ ,
    \new_[8669]_ , \new_[8670]_ , \new_[8671]_ , \new_[8674]_ ,
    \new_[8677]_ , \new_[8678]_ , \new_[8681]_ , \new_[8684]_ ,
    \new_[8685]_ , \new_[8686]_ , \new_[8687]_ , \new_[8691]_ ,
    \new_[8692]_ , \new_[8695]_ , \new_[8698]_ , \new_[8699]_ ,
    \new_[8700]_ , \new_[8703]_ , \new_[8706]_ , \new_[8707]_ ,
    \new_[8710]_ , \new_[8713]_ , \new_[8714]_ , \new_[8715]_ ,
    \new_[8716]_ , \new_[8717]_ , \new_[8718]_ , \new_[8719]_ ,
    \new_[8723]_ , \new_[8724]_ , \new_[8727]_ , \new_[8730]_ ,
    \new_[8731]_ , \new_[8732]_ , \new_[8736]_ , \new_[8737]_ ,
    \new_[8740]_ , \new_[8743]_ , \new_[8744]_ , \new_[8745]_ ,
    \new_[8746]_ , \new_[8750]_ , \new_[8751]_ , \new_[8754]_ ,
    \new_[8757]_ , \new_[8758]_ , \new_[8759]_ , \new_[8762]_ ,
    \new_[8765]_ , \new_[8766]_ , \new_[8769]_ , \new_[8772]_ ,
    \new_[8773]_ , \new_[8774]_ , \new_[8775]_ , \new_[8776]_ ,
    \new_[8780]_ , \new_[8781]_ , \new_[8784]_ , \new_[8787]_ ,
    \new_[8788]_ , \new_[8789]_ , \new_[8792]_ , \new_[8795]_ ,
    \new_[8796]_ , \new_[8799]_ , \new_[8802]_ , \new_[8803]_ ,
    \new_[8804]_ , \new_[8805]_ , \new_[8809]_ , \new_[8810]_ ,
    \new_[8813]_ , \new_[8816]_ , \new_[8817]_ , \new_[8818]_ ,
    \new_[8821]_ , \new_[8824]_ , \new_[8825]_ , \new_[8828]_ ,
    \new_[8831]_ , \new_[8832]_ , \new_[8833]_ , \new_[8834]_ ,
    \new_[8835]_ , \new_[8836]_ , \new_[8840]_ , \new_[8841]_ ,
    \new_[8844]_ , \new_[8847]_ , \new_[8848]_ , \new_[8849]_ ,
    \new_[8853]_ , \new_[8854]_ , \new_[8857]_ , \new_[8860]_ ,
    \new_[8861]_ , \new_[8862]_ , \new_[8863]_ , \new_[8867]_ ,
    \new_[8868]_ , \new_[8871]_ , \new_[8874]_ , \new_[8875]_ ,
    \new_[8876]_ , \new_[8879]_ , \new_[8882]_ , \new_[8883]_ ,
    \new_[8886]_ , \new_[8889]_ , \new_[8890]_ , \new_[8891]_ ,
    \new_[8892]_ , \new_[8893]_ , \new_[8897]_ , \new_[8898]_ ,
    \new_[8901]_ , \new_[8904]_ , \new_[8905]_ , \new_[8906]_ ,
    \new_[8909]_ , \new_[8912]_ , \new_[8913]_ , \new_[8916]_ ,
    \new_[8919]_ , \new_[8920]_ , \new_[8921]_ , \new_[8922]_ ,
    \new_[8926]_ , \new_[8927]_ , \new_[8930]_ , \new_[8933]_ ,
    \new_[8934]_ , \new_[8935]_ , \new_[8938]_ , \new_[8941]_ ,
    \new_[8942]_ , \new_[8945]_ , \new_[8948]_ , \new_[8949]_ ,
    \new_[8950]_ , \new_[8951]_ , \new_[8952]_ , \new_[8953]_ ,
    \new_[8954]_ , \new_[8955]_ , \new_[8959]_ , \new_[8960]_ ,
    \new_[8963]_ , \new_[8966]_ , \new_[8967]_ , \new_[8968]_ ,
    \new_[8972]_ , \new_[8973]_ , \new_[8976]_ , \new_[8979]_ ,
    \new_[8980]_ , \new_[8981]_ , \new_[8982]_ , \new_[8986]_ ,
    \new_[8987]_ , \new_[8990]_ , \new_[8993]_ , \new_[8994]_ ,
    \new_[8995]_ , \new_[8998]_ , \new_[9001]_ , \new_[9002]_ ,
    \new_[9005]_ , \new_[9008]_ , \new_[9009]_ , \new_[9010]_ ,
    \new_[9011]_ , \new_[9012]_ , \new_[9016]_ , \new_[9017]_ ,
    \new_[9020]_ , \new_[9023]_ , \new_[9024]_ , \new_[9025]_ ,
    \new_[9028]_ , \new_[9031]_ , \new_[9032]_ , \new_[9035]_ ,
    \new_[9038]_ , \new_[9039]_ , \new_[9040]_ , \new_[9041]_ ,
    \new_[9045]_ , \new_[9046]_ , \new_[9049]_ , \new_[9052]_ ,
    \new_[9053]_ , \new_[9054]_ , \new_[9057]_ , \new_[9060]_ ,
    \new_[9061]_ , \new_[9064]_ , \new_[9067]_ , \new_[9068]_ ,
    \new_[9069]_ , \new_[9070]_ , \new_[9071]_ , \new_[9072]_ ,
    \new_[9076]_ , \new_[9077]_ , \new_[9080]_ , \new_[9083]_ ,
    \new_[9084]_ , \new_[9085]_ , \new_[9089]_ , \new_[9090]_ ,
    \new_[9093]_ , \new_[9096]_ , \new_[9097]_ , \new_[9098]_ ,
    \new_[9099]_ , \new_[9103]_ , \new_[9104]_ , \new_[9107]_ ,
    \new_[9110]_ , \new_[9111]_ , \new_[9112]_ , \new_[9115]_ ,
    \new_[9118]_ , \new_[9119]_ , \new_[9122]_ , \new_[9125]_ ,
    \new_[9126]_ , \new_[9127]_ , \new_[9128]_ , \new_[9129]_ ,
    \new_[9133]_ , \new_[9134]_ , \new_[9137]_ , \new_[9140]_ ,
    \new_[9141]_ , \new_[9142]_ , \new_[9145]_ , \new_[9148]_ ,
    \new_[9149]_ , \new_[9152]_ , \new_[9155]_ , \new_[9156]_ ,
    \new_[9157]_ , \new_[9158]_ , \new_[9162]_ , \new_[9163]_ ,
    \new_[9166]_ , \new_[9169]_ , \new_[9170]_ , \new_[9171]_ ,
    \new_[9174]_ , \new_[9177]_ , \new_[9178]_ , \new_[9181]_ ,
    \new_[9184]_ , \new_[9185]_ , \new_[9186]_ , \new_[9187]_ ,
    \new_[9188]_ , \new_[9189]_ , \new_[9190]_ , \new_[9194]_ ,
    \new_[9195]_ , \new_[9198]_ , \new_[9201]_ , \new_[9202]_ ,
    \new_[9203]_ , \new_[9207]_ , \new_[9208]_ , \new_[9211]_ ,
    \new_[9214]_ , \new_[9215]_ , \new_[9216]_ , \new_[9217]_ ,
    \new_[9221]_ , \new_[9222]_ , \new_[9225]_ , \new_[9228]_ ,
    \new_[9229]_ , \new_[9230]_ , \new_[9233]_ , \new_[9236]_ ,
    \new_[9237]_ , \new_[9240]_ , \new_[9243]_ , \new_[9244]_ ,
    \new_[9245]_ , \new_[9246]_ , \new_[9247]_ , \new_[9251]_ ,
    \new_[9252]_ , \new_[9255]_ , \new_[9258]_ , \new_[9259]_ ,
    \new_[9260]_ , \new_[9263]_ , \new_[9266]_ , \new_[9267]_ ,
    \new_[9270]_ , \new_[9273]_ , \new_[9274]_ , \new_[9275]_ ,
    \new_[9276]_ , \new_[9280]_ , \new_[9281]_ , \new_[9284]_ ,
    \new_[9287]_ , \new_[9288]_ , \new_[9289]_ , \new_[9292]_ ,
    \new_[9295]_ , \new_[9296]_ , \new_[9299]_ , \new_[9302]_ ,
    \new_[9303]_ , \new_[9304]_ , \new_[9305]_ , \new_[9306]_ ,
    \new_[9307]_ , \new_[9311]_ , \new_[9312]_ , \new_[9315]_ ,
    \new_[9318]_ , \new_[9319]_ , \new_[9320]_ , \new_[9324]_ ,
    \new_[9325]_ , \new_[9328]_ , \new_[9331]_ , \new_[9332]_ ,
    \new_[9333]_ , \new_[9334]_ , \new_[9338]_ , \new_[9339]_ ,
    \new_[9342]_ , \new_[9345]_ , \new_[9346]_ , \new_[9347]_ ,
    \new_[9350]_ , \new_[9353]_ , \new_[9354]_ , \new_[9357]_ ,
    \new_[9360]_ , \new_[9361]_ , \new_[9362]_ , \new_[9363]_ ,
    \new_[9364]_ , \new_[9368]_ , \new_[9369]_ , \new_[9372]_ ,
    \new_[9375]_ , \new_[9376]_ , \new_[9377]_ , \new_[9380]_ ,
    \new_[9383]_ , \new_[9384]_ , \new_[9387]_ , \new_[9390]_ ,
    \new_[9391]_ , \new_[9392]_ , \new_[9393]_ , \new_[9397]_ ,
    \new_[9398]_ , \new_[9401]_ , \new_[9404]_ , \new_[9405]_ ,
    \new_[9406]_ , \new_[9409]_ , \new_[9412]_ , \new_[9413]_ ,
    \new_[9416]_ , \new_[9419]_ , \new_[9420]_ , \new_[9421]_ ,
    \new_[9422]_ , \new_[9423]_ , \new_[9424]_ , \new_[9425]_ ,
    \new_[9426]_ , \new_[9427]_ , \new_[9428]_ , \new_[9432]_ ,
    \new_[9433]_ , \new_[9436]_ , \new_[9439]_ , \new_[9440]_ ,
    \new_[9441]_ , \new_[9445]_ , \new_[9446]_ , \new_[9449]_ ,
    \new_[9452]_ , \new_[9453]_ , \new_[9454]_ , \new_[9455]_ ,
    \new_[9459]_ , \new_[9460]_ , \new_[9463]_ , \new_[9466]_ ,
    \new_[9467]_ , \new_[9468]_ , \new_[9471]_ , \new_[9474]_ ,
    \new_[9475]_ , \new_[9478]_ , \new_[9481]_ , \new_[9482]_ ,
    \new_[9483]_ , \new_[9484]_ , \new_[9485]_ , \new_[9489]_ ,
    \new_[9490]_ , \new_[9493]_ , \new_[9496]_ , \new_[9497]_ ,
    \new_[9498]_ , \new_[9502]_ , \new_[9503]_ , \new_[9506]_ ,
    \new_[9509]_ , \new_[9510]_ , \new_[9511]_ , \new_[9512]_ ,
    \new_[9516]_ , \new_[9517]_ , \new_[9520]_ , \new_[9523]_ ,
    \new_[9524]_ , \new_[9525]_ , \new_[9528]_ , \new_[9531]_ ,
    \new_[9532]_ , \new_[9535]_ , \new_[9538]_ , \new_[9539]_ ,
    \new_[9540]_ , \new_[9541]_ , \new_[9542]_ , \new_[9543]_ ,
    \new_[9547]_ , \new_[9548]_ , \new_[9551]_ , \new_[9554]_ ,
    \new_[9555]_ , \new_[9556]_ , \new_[9560]_ , \new_[9561]_ ,
    \new_[9564]_ , \new_[9567]_ , \new_[9568]_ , \new_[9569]_ ,
    \new_[9570]_ , \new_[9574]_ , \new_[9575]_ , \new_[9578]_ ,
    \new_[9581]_ , \new_[9582]_ , \new_[9583]_ , \new_[9586]_ ,
    \new_[9589]_ , \new_[9590]_ , \new_[9593]_ , \new_[9596]_ ,
    \new_[9597]_ , \new_[9598]_ , \new_[9599]_ , \new_[9600]_ ,
    \new_[9604]_ , \new_[9605]_ , \new_[9608]_ , \new_[9611]_ ,
    \new_[9612]_ , \new_[9613]_ , \new_[9616]_ , \new_[9619]_ ,
    \new_[9620]_ , \new_[9623]_ , \new_[9626]_ , \new_[9627]_ ,
    \new_[9628]_ , \new_[9629]_ , \new_[9633]_ , \new_[9634]_ ,
    \new_[9637]_ , \new_[9640]_ , \new_[9641]_ , \new_[9642]_ ,
    \new_[9645]_ , \new_[9648]_ , \new_[9649]_ , \new_[9652]_ ,
    \new_[9655]_ , \new_[9656]_ , \new_[9657]_ , \new_[9658]_ ,
    \new_[9659]_ , \new_[9660]_ , \new_[9661]_ , \new_[9665]_ ,
    \new_[9666]_ , \new_[9669]_ , \new_[9672]_ , \new_[9673]_ ,
    \new_[9674]_ , \new_[9678]_ , \new_[9679]_ , \new_[9682]_ ,
    \new_[9685]_ , \new_[9686]_ , \new_[9687]_ , \new_[9688]_ ,
    \new_[9692]_ , \new_[9693]_ , \new_[9696]_ , \new_[9699]_ ,
    \new_[9700]_ , \new_[9701]_ , \new_[9704]_ , \new_[9707]_ ,
    \new_[9708]_ , \new_[9711]_ , \new_[9714]_ , \new_[9715]_ ,
    \new_[9716]_ , \new_[9717]_ , \new_[9718]_ , \new_[9722]_ ,
    \new_[9723]_ , \new_[9726]_ , \new_[9729]_ , \new_[9730]_ ,
    \new_[9731]_ , \new_[9734]_ , \new_[9737]_ , \new_[9738]_ ,
    \new_[9741]_ , \new_[9744]_ , \new_[9745]_ , \new_[9746]_ ,
    \new_[9747]_ , \new_[9751]_ , \new_[9752]_ , \new_[9755]_ ,
    \new_[9758]_ , \new_[9759]_ , \new_[9760]_ , \new_[9763]_ ,
    \new_[9766]_ , \new_[9767]_ , \new_[9770]_ , \new_[9773]_ ,
    \new_[9774]_ , \new_[9775]_ , \new_[9776]_ , \new_[9777]_ ,
    \new_[9778]_ , \new_[9782]_ , \new_[9783]_ , \new_[9786]_ ,
    \new_[9789]_ , \new_[9790]_ , \new_[9791]_ , \new_[9795]_ ,
    \new_[9796]_ , \new_[9799]_ , \new_[9802]_ , \new_[9803]_ ,
    \new_[9804]_ , \new_[9805]_ , \new_[9809]_ , \new_[9810]_ ,
    \new_[9813]_ , \new_[9816]_ , \new_[9817]_ , \new_[9818]_ ,
    \new_[9821]_ , \new_[9824]_ , \new_[9825]_ , \new_[9828]_ ,
    \new_[9831]_ , \new_[9832]_ , \new_[9833]_ , \new_[9834]_ ,
    \new_[9835]_ , \new_[9839]_ , \new_[9840]_ , \new_[9843]_ ,
    \new_[9846]_ , \new_[9847]_ , \new_[9848]_ , \new_[9851]_ ,
    \new_[9854]_ , \new_[9855]_ , \new_[9858]_ , \new_[9861]_ ,
    \new_[9862]_ , \new_[9863]_ , \new_[9864]_ , \new_[9868]_ ,
    \new_[9869]_ , \new_[9872]_ , \new_[9875]_ , \new_[9876]_ ,
    \new_[9877]_ , \new_[9880]_ , \new_[9883]_ , \new_[9884]_ ,
    \new_[9887]_ , \new_[9890]_ , \new_[9891]_ , \new_[9892]_ ,
    \new_[9893]_ , \new_[9894]_ , \new_[9895]_ , \new_[9896]_ ,
    \new_[9897]_ , \new_[9901]_ , \new_[9902]_ , \new_[9905]_ ,
    \new_[9908]_ , \new_[9909]_ , \new_[9910]_ , \new_[9914]_ ,
    \new_[9915]_ , \new_[9918]_ , \new_[9921]_ , \new_[9922]_ ,
    \new_[9923]_ , \new_[9924]_ , \new_[9928]_ , \new_[9929]_ ,
    \new_[9932]_ , \new_[9935]_ , \new_[9936]_ , \new_[9937]_ ,
    \new_[9940]_ , \new_[9943]_ , \new_[9944]_ , \new_[9947]_ ,
    \new_[9950]_ , \new_[9951]_ , \new_[9952]_ , \new_[9953]_ ,
    \new_[9954]_ , \new_[9958]_ , \new_[9959]_ , \new_[9962]_ ,
    \new_[9965]_ , \new_[9966]_ , \new_[9967]_ , \new_[9970]_ ,
    \new_[9973]_ , \new_[9974]_ , \new_[9977]_ , \new_[9980]_ ,
    \new_[9981]_ , \new_[9982]_ , \new_[9983]_ , \new_[9987]_ ,
    \new_[9988]_ , \new_[9991]_ , \new_[9994]_ , \new_[9995]_ ,
    \new_[9996]_ , \new_[9999]_ , \new_[10002]_ , \new_[10003]_ ,
    \new_[10006]_ , \new_[10009]_ , \new_[10010]_ , \new_[10011]_ ,
    \new_[10012]_ , \new_[10013]_ , \new_[10014]_ , \new_[10018]_ ,
    \new_[10019]_ , \new_[10022]_ , \new_[10025]_ , \new_[10026]_ ,
    \new_[10027]_ , \new_[10031]_ , \new_[10032]_ , \new_[10035]_ ,
    \new_[10038]_ , \new_[10039]_ , \new_[10040]_ , \new_[10041]_ ,
    \new_[10045]_ , \new_[10046]_ , \new_[10049]_ , \new_[10052]_ ,
    \new_[10053]_ , \new_[10054]_ , \new_[10057]_ , \new_[10060]_ ,
    \new_[10061]_ , \new_[10064]_ , \new_[10067]_ , \new_[10068]_ ,
    \new_[10069]_ , \new_[10070]_ , \new_[10071]_ , \new_[10075]_ ,
    \new_[10076]_ , \new_[10079]_ , \new_[10082]_ , \new_[10083]_ ,
    \new_[10084]_ , \new_[10087]_ , \new_[10090]_ , \new_[10091]_ ,
    \new_[10094]_ , \new_[10097]_ , \new_[10098]_ , \new_[10099]_ ,
    \new_[10100]_ , \new_[10104]_ , \new_[10105]_ , \new_[10108]_ ,
    \new_[10111]_ , \new_[10112]_ , \new_[10113]_ , \new_[10116]_ ,
    \new_[10119]_ , \new_[10120]_ , \new_[10123]_ , \new_[10126]_ ,
    \new_[10127]_ , \new_[10128]_ , \new_[10129]_ , \new_[10130]_ ,
    \new_[10131]_ , \new_[10132]_ , \new_[10136]_ , \new_[10137]_ ,
    \new_[10140]_ , \new_[10143]_ , \new_[10144]_ , \new_[10145]_ ,
    \new_[10149]_ , \new_[10150]_ , \new_[10153]_ , \new_[10156]_ ,
    \new_[10157]_ , \new_[10158]_ , \new_[10159]_ , \new_[10163]_ ,
    \new_[10164]_ , \new_[10167]_ , \new_[10170]_ , \new_[10171]_ ,
    \new_[10172]_ , \new_[10175]_ , \new_[10178]_ , \new_[10179]_ ,
    \new_[10182]_ , \new_[10185]_ , \new_[10186]_ , \new_[10187]_ ,
    \new_[10188]_ , \new_[10189]_ , \new_[10193]_ , \new_[10194]_ ,
    \new_[10197]_ , \new_[10200]_ , \new_[10201]_ , \new_[10202]_ ,
    \new_[10205]_ , \new_[10208]_ , \new_[10209]_ , \new_[10212]_ ,
    \new_[10215]_ , \new_[10216]_ , \new_[10217]_ , \new_[10218]_ ,
    \new_[10222]_ , \new_[10223]_ , \new_[10226]_ , \new_[10229]_ ,
    \new_[10230]_ , \new_[10231]_ , \new_[10234]_ , \new_[10237]_ ,
    \new_[10238]_ , \new_[10241]_ , \new_[10244]_ , \new_[10245]_ ,
    \new_[10246]_ , \new_[10247]_ , \new_[10248]_ , \new_[10249]_ ,
    \new_[10253]_ , \new_[10254]_ , \new_[10257]_ , \new_[10260]_ ,
    \new_[10261]_ , \new_[10262]_ , \new_[10266]_ , \new_[10267]_ ,
    \new_[10270]_ , \new_[10273]_ , \new_[10274]_ , \new_[10275]_ ,
    \new_[10276]_ , \new_[10280]_ , \new_[10281]_ , \new_[10284]_ ,
    \new_[10287]_ , \new_[10288]_ , \new_[10289]_ , \new_[10292]_ ,
    \new_[10295]_ , \new_[10296]_ , \new_[10299]_ , \new_[10302]_ ,
    \new_[10303]_ , \new_[10304]_ , \new_[10305]_ , \new_[10306]_ ,
    \new_[10310]_ , \new_[10311]_ , \new_[10314]_ , \new_[10317]_ ,
    \new_[10318]_ , \new_[10319]_ , \new_[10322]_ , \new_[10325]_ ,
    \new_[10326]_ , \new_[10329]_ , \new_[10332]_ , \new_[10333]_ ,
    \new_[10334]_ , \new_[10335]_ , \new_[10339]_ , \new_[10340]_ ,
    \new_[10343]_ , \new_[10346]_ , \new_[10347]_ , \new_[10348]_ ,
    \new_[10351]_ , \new_[10354]_ , \new_[10355]_ , \new_[10358]_ ,
    \new_[10361]_ , \new_[10362]_ , \new_[10363]_ , \new_[10364]_ ,
    \new_[10365]_ , \new_[10366]_ , \new_[10367]_ , \new_[10368]_ ,
    \new_[10369]_ , \new_[10373]_ , \new_[10374]_ , \new_[10377]_ ,
    \new_[10380]_ , \new_[10381]_ , \new_[10382]_ , \new_[10386]_ ,
    \new_[10387]_ , \new_[10390]_ , \new_[10393]_ , \new_[10394]_ ,
    \new_[10395]_ , \new_[10396]_ , \new_[10400]_ , \new_[10401]_ ,
    \new_[10404]_ , \new_[10407]_ , \new_[10408]_ , \new_[10409]_ ,
    \new_[10412]_ , \new_[10415]_ , \new_[10416]_ , \new_[10419]_ ,
    \new_[10422]_ , \new_[10423]_ , \new_[10424]_ , \new_[10425]_ ,
    \new_[10426]_ , \new_[10430]_ , \new_[10431]_ , \new_[10434]_ ,
    \new_[10437]_ , \new_[10438]_ , \new_[10439]_ , \new_[10442]_ ,
    \new_[10445]_ , \new_[10446]_ , \new_[10449]_ , \new_[10452]_ ,
    \new_[10453]_ , \new_[10454]_ , \new_[10455]_ , \new_[10459]_ ,
    \new_[10460]_ , \new_[10463]_ , \new_[10466]_ , \new_[10467]_ ,
    \new_[10468]_ , \new_[10471]_ , \new_[10474]_ , \new_[10475]_ ,
    \new_[10478]_ , \new_[10481]_ , \new_[10482]_ , \new_[10483]_ ,
    \new_[10484]_ , \new_[10485]_ , \new_[10486]_ , \new_[10490]_ ,
    \new_[10491]_ , \new_[10494]_ , \new_[10497]_ , \new_[10498]_ ,
    \new_[10499]_ , \new_[10503]_ , \new_[10504]_ , \new_[10507]_ ,
    \new_[10510]_ , \new_[10511]_ , \new_[10512]_ , \new_[10513]_ ,
    \new_[10517]_ , \new_[10518]_ , \new_[10521]_ , \new_[10524]_ ,
    \new_[10525]_ , \new_[10526]_ , \new_[10529]_ , \new_[10532]_ ,
    \new_[10533]_ , \new_[10536]_ , \new_[10539]_ , \new_[10540]_ ,
    \new_[10541]_ , \new_[10542]_ , \new_[10543]_ , \new_[10547]_ ,
    \new_[10548]_ , \new_[10551]_ , \new_[10554]_ , \new_[10555]_ ,
    \new_[10556]_ , \new_[10559]_ , \new_[10562]_ , \new_[10563]_ ,
    \new_[10566]_ , \new_[10569]_ , \new_[10570]_ , \new_[10571]_ ,
    \new_[10572]_ , \new_[10576]_ , \new_[10577]_ , \new_[10580]_ ,
    \new_[10583]_ , \new_[10584]_ , \new_[10585]_ , \new_[10588]_ ,
    \new_[10591]_ , \new_[10592]_ , \new_[10595]_ , \new_[10598]_ ,
    \new_[10599]_ , \new_[10600]_ , \new_[10601]_ , \new_[10602]_ ,
    \new_[10603]_ , \new_[10604]_ , \new_[10608]_ , \new_[10609]_ ,
    \new_[10612]_ , \new_[10615]_ , \new_[10616]_ , \new_[10617]_ ,
    \new_[10621]_ , \new_[10622]_ , \new_[10625]_ , \new_[10628]_ ,
    \new_[10629]_ , \new_[10630]_ , \new_[10631]_ , \new_[10635]_ ,
    \new_[10636]_ , \new_[10639]_ , \new_[10642]_ , \new_[10643]_ ,
    \new_[10644]_ , \new_[10647]_ , \new_[10650]_ , \new_[10651]_ ,
    \new_[10654]_ , \new_[10657]_ , \new_[10658]_ , \new_[10659]_ ,
    \new_[10660]_ , \new_[10661]_ , \new_[10665]_ , \new_[10666]_ ,
    \new_[10669]_ , \new_[10672]_ , \new_[10673]_ , \new_[10674]_ ,
    \new_[10677]_ , \new_[10680]_ , \new_[10681]_ , \new_[10684]_ ,
    \new_[10687]_ , \new_[10688]_ , \new_[10689]_ , \new_[10690]_ ,
    \new_[10694]_ , \new_[10695]_ , \new_[10698]_ , \new_[10701]_ ,
    \new_[10702]_ , \new_[10703]_ , \new_[10706]_ , \new_[10709]_ ,
    \new_[10710]_ , \new_[10713]_ , \new_[10716]_ , \new_[10717]_ ,
    \new_[10718]_ , \new_[10719]_ , \new_[10720]_ , \new_[10721]_ ,
    \new_[10725]_ , \new_[10726]_ , \new_[10729]_ , \new_[10732]_ ,
    \new_[10733]_ , \new_[10734]_ , \new_[10738]_ , \new_[10739]_ ,
    \new_[10742]_ , \new_[10745]_ , \new_[10746]_ , \new_[10747]_ ,
    \new_[10748]_ , \new_[10752]_ , \new_[10753]_ , \new_[10756]_ ,
    \new_[10759]_ , \new_[10760]_ , \new_[10761]_ , \new_[10764]_ ,
    \new_[10767]_ , \new_[10768]_ , \new_[10771]_ , \new_[10774]_ ,
    \new_[10775]_ , \new_[10776]_ , \new_[10777]_ , \new_[10778]_ ,
    \new_[10782]_ , \new_[10783]_ , \new_[10786]_ , \new_[10789]_ ,
    \new_[10790]_ , \new_[10791]_ , \new_[10794]_ , \new_[10797]_ ,
    \new_[10798]_ , \new_[10801]_ , \new_[10804]_ , \new_[10805]_ ,
    \new_[10806]_ , \new_[10807]_ , \new_[10811]_ , \new_[10812]_ ,
    \new_[10815]_ , \new_[10818]_ , \new_[10819]_ , \new_[10820]_ ,
    \new_[10823]_ , \new_[10826]_ , \new_[10827]_ , \new_[10830]_ ,
    \new_[10833]_ , \new_[10834]_ , \new_[10835]_ , \new_[10836]_ ,
    \new_[10837]_ , \new_[10838]_ , \new_[10839]_ , \new_[10840]_ ,
    \new_[10844]_ , \new_[10845]_ , \new_[10848]_ , \new_[10851]_ ,
    \new_[10852]_ , \new_[10853]_ , \new_[10857]_ , \new_[10858]_ ,
    \new_[10861]_ , \new_[10864]_ , \new_[10865]_ , \new_[10866]_ ,
    \new_[10867]_ , \new_[10871]_ , \new_[10872]_ , \new_[10875]_ ,
    \new_[10878]_ , \new_[10879]_ , \new_[10880]_ , \new_[10883]_ ,
    \new_[10886]_ , \new_[10887]_ , \new_[10890]_ , \new_[10893]_ ,
    \new_[10894]_ , \new_[10895]_ , \new_[10896]_ , \new_[10897]_ ,
    \new_[10901]_ , \new_[10902]_ , \new_[10905]_ , \new_[10908]_ ,
    \new_[10909]_ , \new_[10910]_ , \new_[10913]_ , \new_[10916]_ ,
    \new_[10917]_ , \new_[10920]_ , \new_[10923]_ , \new_[10924]_ ,
    \new_[10925]_ , \new_[10926]_ , \new_[10930]_ , \new_[10931]_ ,
    \new_[10934]_ , \new_[10937]_ , \new_[10938]_ , \new_[10939]_ ,
    \new_[10942]_ , \new_[10945]_ , \new_[10946]_ , \new_[10949]_ ,
    \new_[10952]_ , \new_[10953]_ , \new_[10954]_ , \new_[10955]_ ,
    \new_[10956]_ , \new_[10957]_ , \new_[10961]_ , \new_[10962]_ ,
    \new_[10965]_ , \new_[10968]_ , \new_[10969]_ , \new_[10970]_ ,
    \new_[10974]_ , \new_[10975]_ , \new_[10978]_ , \new_[10981]_ ,
    \new_[10982]_ , \new_[10983]_ , \new_[10984]_ , \new_[10988]_ ,
    \new_[10989]_ , \new_[10992]_ , \new_[10995]_ , \new_[10996]_ ,
    \new_[10997]_ , \new_[11000]_ , \new_[11003]_ , \new_[11004]_ ,
    \new_[11007]_ , \new_[11010]_ , \new_[11011]_ , \new_[11012]_ ,
    \new_[11013]_ , \new_[11014]_ , \new_[11018]_ , \new_[11019]_ ,
    \new_[11022]_ , \new_[11025]_ , \new_[11026]_ , \new_[11027]_ ,
    \new_[11030]_ , \new_[11033]_ , \new_[11034]_ , \new_[11037]_ ,
    \new_[11040]_ , \new_[11041]_ , \new_[11042]_ , \new_[11043]_ ,
    \new_[11047]_ , \new_[11048]_ , \new_[11051]_ , \new_[11054]_ ,
    \new_[11055]_ , \new_[11056]_ , \new_[11059]_ , \new_[11062]_ ,
    \new_[11063]_ , \new_[11066]_ , \new_[11069]_ , \new_[11070]_ ,
    \new_[11071]_ , \new_[11072]_ , \new_[11073]_ , \new_[11074]_ ,
    \new_[11075]_ , \new_[11079]_ , \new_[11080]_ , \new_[11083]_ ,
    \new_[11086]_ , \new_[11087]_ , \new_[11088]_ , \new_[11092]_ ,
    \new_[11093]_ , \new_[11096]_ , \new_[11099]_ , \new_[11100]_ ,
    \new_[11101]_ , \new_[11102]_ , \new_[11106]_ , \new_[11107]_ ,
    \new_[11110]_ , \new_[11113]_ , \new_[11114]_ , \new_[11115]_ ,
    \new_[11118]_ , \new_[11121]_ , \new_[11122]_ , \new_[11125]_ ,
    \new_[11128]_ , \new_[11129]_ , \new_[11130]_ , \new_[11131]_ ,
    \new_[11132]_ , \new_[11136]_ , \new_[11137]_ , \new_[11140]_ ,
    \new_[11143]_ , \new_[11144]_ , \new_[11145]_ , \new_[11148]_ ,
    \new_[11151]_ , \new_[11152]_ , \new_[11155]_ , \new_[11158]_ ,
    \new_[11159]_ , \new_[11160]_ , \new_[11161]_ , \new_[11165]_ ,
    \new_[11166]_ , \new_[11169]_ , \new_[11172]_ , \new_[11173]_ ,
    \new_[11174]_ , \new_[11177]_ , \new_[11180]_ , \new_[11181]_ ,
    \new_[11184]_ , \new_[11187]_ , \new_[11188]_ , \new_[11189]_ ,
    \new_[11190]_ , \new_[11191]_ , \new_[11192]_ , \new_[11196]_ ,
    \new_[11197]_ , \new_[11200]_ , \new_[11203]_ , \new_[11204]_ ,
    \new_[11205]_ , \new_[11209]_ , \new_[11210]_ , \new_[11213]_ ,
    \new_[11216]_ , \new_[11217]_ , \new_[11218]_ , \new_[11219]_ ,
    \new_[11223]_ , \new_[11224]_ , \new_[11227]_ , \new_[11230]_ ,
    \new_[11231]_ , \new_[11232]_ , \new_[11235]_ , \new_[11238]_ ,
    \new_[11239]_ , \new_[11242]_ , \new_[11245]_ , \new_[11246]_ ,
    \new_[11247]_ , \new_[11248]_ , \new_[11249]_ , \new_[11253]_ ,
    \new_[11254]_ , \new_[11257]_ , \new_[11260]_ , \new_[11261]_ ,
    \new_[11262]_ , \new_[11265]_ , \new_[11268]_ , \new_[11269]_ ,
    \new_[11272]_ , \new_[11275]_ , \new_[11276]_ , \new_[11277]_ ,
    \new_[11278]_ , \new_[11282]_ , \new_[11283]_ , \new_[11286]_ ,
    \new_[11289]_ , \new_[11290]_ , \new_[11291]_ , \new_[11294]_ ,
    \new_[11297]_ , \new_[11298]_ , \new_[11301]_ , \new_[11304]_ ,
    \new_[11305]_ , \new_[11306]_ , \new_[11307]_ , \new_[11308]_ ,
    \new_[11309]_ , \new_[11310]_ , \new_[11311]_ , \new_[11312]_ ,
    \new_[11313]_ , \new_[11314]_ , \new_[11317]_ , \new_[11320]_ ,
    \new_[11321]_ , \new_[11324]_ , \new_[11327]_ , \new_[11328]_ ,
    \new_[11331]_ , \new_[11334]_ , \new_[11335]_ , \new_[11338]_ ,
    \new_[11341]_ , \new_[11342]_ , \new_[11345]_ , \new_[11348]_ ,
    \new_[11349]_ , \new_[11352]_ , \new_[11355]_ , \new_[11356]_ ,
    \new_[11359]_ , \new_[11362]_ , \new_[11363]_ , \new_[11366]_ ,
    \new_[11369]_ , \new_[11370]_ , \new_[11373]_ , \new_[11376]_ ,
    \new_[11377]_ , \new_[11380]_ , \new_[11383]_ , \new_[11384]_ ,
    \new_[11387]_ , \new_[11390]_ , \new_[11391]_ , \new_[11394]_ ,
    \new_[11397]_ , \new_[11398]_ , \new_[11401]_ , \new_[11404]_ ,
    \new_[11405]_ , \new_[11408]_ , \new_[11411]_ , \new_[11412]_ ,
    \new_[11415]_ , \new_[11418]_ , \new_[11419]_ , \new_[11422]_ ,
    \new_[11425]_ , \new_[11426]_ , \new_[11429]_ , \new_[11432]_ ,
    \new_[11433]_ , \new_[11436]_ , \new_[11439]_ , \new_[11440]_ ,
    \new_[11443]_ , \new_[11446]_ , \new_[11447]_ , \new_[11450]_ ,
    \new_[11453]_ , \new_[11454]_ , \new_[11457]_ , \new_[11460]_ ,
    \new_[11461]_ , \new_[11464]_ , \new_[11467]_ , \new_[11468]_ ,
    \new_[11471]_ , \new_[11474]_ , \new_[11475]_ , \new_[11478]_ ,
    \new_[11481]_ , \new_[11482]_ , \new_[11485]_ , \new_[11488]_ ,
    \new_[11489]_ , \new_[11492]_ , \new_[11496]_ , \new_[11497]_ ,
    \new_[11498]_ , \new_[11501]_ , \new_[11504]_ , \new_[11505]_ ,
    \new_[11508]_ , \new_[11512]_ , \new_[11513]_ , \new_[11514]_ ,
    \new_[11517]_ , \new_[11520]_ , \new_[11521]_ , \new_[11524]_ ,
    \new_[11528]_ , \new_[11529]_ , \new_[11530]_ , \new_[11533]_ ,
    \new_[11536]_ , \new_[11537]_ , \new_[11540]_ , \new_[11544]_ ,
    \new_[11545]_ , \new_[11546]_ , \new_[11549]_ , \new_[11552]_ ,
    \new_[11553]_ , \new_[11556]_ , \new_[11560]_ , \new_[11561]_ ,
    \new_[11562]_ , \new_[11565]_ , \new_[11568]_ , \new_[11569]_ ,
    \new_[11572]_ , \new_[11576]_ , \new_[11577]_ , \new_[11578]_ ,
    \new_[11581]_ , \new_[11584]_ , \new_[11585]_ , \new_[11588]_ ,
    \new_[11592]_ , \new_[11593]_ , \new_[11594]_ , \new_[11597]_ ,
    \new_[11600]_ , \new_[11601]_ , \new_[11604]_ , \new_[11608]_ ,
    \new_[11609]_ , \new_[11610]_ , \new_[11613]_ , \new_[11617]_ ,
    \new_[11618]_ , \new_[11619]_ , \new_[11622]_ , \new_[11626]_ ,
    \new_[11627]_ , \new_[11628]_ , \new_[11631]_ , \new_[11635]_ ,
    \new_[11636]_ , \new_[11637]_ , \new_[11640]_ , \new_[11644]_ ,
    \new_[11645]_ , \new_[11646]_ , \new_[11649]_ , \new_[11653]_ ,
    \new_[11654]_ , \new_[11655]_ , \new_[11658]_ , \new_[11662]_ ,
    \new_[11663]_ , \new_[11664]_ , \new_[11667]_ , \new_[11671]_ ,
    \new_[11672]_ , \new_[11673]_ , \new_[11676]_ , \new_[11680]_ ,
    \new_[11681]_ , \new_[11682]_ , \new_[11685]_ , \new_[11689]_ ,
    \new_[11690]_ , \new_[11691]_ , \new_[11694]_ , \new_[11698]_ ,
    \new_[11699]_ , \new_[11700]_ , \new_[11703]_ , \new_[11707]_ ,
    \new_[11708]_ , \new_[11709]_ , \new_[11712]_ , \new_[11716]_ ,
    \new_[11717]_ , \new_[11718]_ , \new_[11721]_ , \new_[11725]_ ,
    \new_[11726]_ , \new_[11727]_ , \new_[11730]_ , \new_[11734]_ ,
    \new_[11735]_ , \new_[11736]_ , \new_[11739]_ , \new_[11743]_ ,
    \new_[11744]_ , \new_[11745]_ , \new_[11748]_ , \new_[11752]_ ,
    \new_[11753]_ , \new_[11754]_ , \new_[11757]_ , \new_[11761]_ ,
    \new_[11762]_ , \new_[11763]_ , \new_[11766]_ , \new_[11770]_ ,
    \new_[11771]_ , \new_[11772]_ , \new_[11775]_ , \new_[11779]_ ,
    \new_[11780]_ , \new_[11781]_ , \new_[11784]_ , \new_[11788]_ ,
    \new_[11789]_ , \new_[11790]_ , \new_[11793]_ , \new_[11797]_ ,
    \new_[11798]_ , \new_[11799]_ , \new_[11802]_ , \new_[11806]_ ,
    \new_[11807]_ , \new_[11808]_ , \new_[11811]_ , \new_[11815]_ ,
    \new_[11816]_ , \new_[11817]_ , \new_[11820]_ , \new_[11824]_ ,
    \new_[11825]_ , \new_[11826]_ , \new_[11829]_ , \new_[11833]_ ,
    \new_[11834]_ , \new_[11835]_ , \new_[11838]_ , \new_[11842]_ ,
    \new_[11843]_ , \new_[11844]_ , \new_[11847]_ , \new_[11851]_ ,
    \new_[11852]_ , \new_[11853]_ , \new_[11856]_ , \new_[11860]_ ,
    \new_[11861]_ , \new_[11862]_ , \new_[11865]_ , \new_[11869]_ ,
    \new_[11870]_ , \new_[11871]_ , \new_[11874]_ , \new_[11878]_ ,
    \new_[11879]_ , \new_[11880]_ , \new_[11883]_ , \new_[11887]_ ,
    \new_[11888]_ , \new_[11889]_ , \new_[11892]_ , \new_[11896]_ ,
    \new_[11897]_ , \new_[11898]_ , \new_[11901]_ , \new_[11905]_ ,
    \new_[11906]_ , \new_[11907]_ , \new_[11910]_ , \new_[11914]_ ,
    \new_[11915]_ , \new_[11916]_ , \new_[11919]_ , \new_[11923]_ ,
    \new_[11924]_ , \new_[11925]_ , \new_[11928]_ , \new_[11932]_ ,
    \new_[11933]_ , \new_[11934]_ , \new_[11937]_ , \new_[11941]_ ,
    \new_[11942]_ , \new_[11943]_ , \new_[11946]_ , \new_[11950]_ ,
    \new_[11951]_ , \new_[11952]_ , \new_[11955]_ , \new_[11959]_ ,
    \new_[11960]_ , \new_[11961]_ , \new_[11964]_ , \new_[11968]_ ,
    \new_[11969]_ , \new_[11970]_ , \new_[11973]_ , \new_[11977]_ ,
    \new_[11978]_ , \new_[11979]_ , \new_[11982]_ , \new_[11986]_ ,
    \new_[11987]_ , \new_[11988]_ , \new_[11991]_ , \new_[11995]_ ,
    \new_[11996]_ , \new_[11997]_ , \new_[12000]_ , \new_[12004]_ ,
    \new_[12005]_ , \new_[12006]_ , \new_[12009]_ , \new_[12013]_ ,
    \new_[12014]_ , \new_[12015]_ , \new_[12018]_ , \new_[12022]_ ,
    \new_[12023]_ , \new_[12024]_ , \new_[12027]_ , \new_[12031]_ ,
    \new_[12032]_ , \new_[12033]_ , \new_[12036]_ , \new_[12040]_ ,
    \new_[12041]_ , \new_[12042]_ , \new_[12045]_ , \new_[12049]_ ,
    \new_[12050]_ , \new_[12051]_ , \new_[12054]_ , \new_[12058]_ ,
    \new_[12059]_ , \new_[12060]_ , \new_[12063]_ , \new_[12067]_ ,
    \new_[12068]_ , \new_[12069]_ , \new_[12072]_ , \new_[12076]_ ,
    \new_[12077]_ , \new_[12078]_ , \new_[12081]_ , \new_[12085]_ ,
    \new_[12086]_ , \new_[12087]_ , \new_[12090]_ , \new_[12094]_ ,
    \new_[12095]_ , \new_[12096]_ , \new_[12099]_ , \new_[12103]_ ,
    \new_[12104]_ , \new_[12105]_ , \new_[12108]_ , \new_[12112]_ ,
    \new_[12113]_ , \new_[12114]_ , \new_[12117]_ , \new_[12121]_ ,
    \new_[12122]_ , \new_[12123]_ , \new_[12126]_ , \new_[12130]_ ,
    \new_[12131]_ , \new_[12132]_ , \new_[12135]_ , \new_[12139]_ ,
    \new_[12140]_ , \new_[12141]_ , \new_[12144]_ , \new_[12148]_ ,
    \new_[12149]_ , \new_[12150]_ , \new_[12153]_ , \new_[12157]_ ,
    \new_[12158]_ , \new_[12159]_ , \new_[12162]_ , \new_[12166]_ ,
    \new_[12167]_ , \new_[12168]_ , \new_[12171]_ , \new_[12175]_ ,
    \new_[12176]_ , \new_[12177]_ , \new_[12180]_ , \new_[12184]_ ,
    \new_[12185]_ , \new_[12186]_ , \new_[12189]_ , \new_[12193]_ ,
    \new_[12194]_ , \new_[12195]_ , \new_[12198]_ , \new_[12202]_ ,
    \new_[12203]_ , \new_[12204]_ , \new_[12207]_ , \new_[12211]_ ,
    \new_[12212]_ , \new_[12213]_ , \new_[12216]_ , \new_[12220]_ ,
    \new_[12221]_ , \new_[12222]_ , \new_[12225]_ , \new_[12229]_ ,
    \new_[12230]_ , \new_[12231]_ , \new_[12234]_ , \new_[12238]_ ,
    \new_[12239]_ , \new_[12240]_ , \new_[12243]_ , \new_[12247]_ ,
    \new_[12248]_ , \new_[12249]_ , \new_[12252]_ , \new_[12256]_ ,
    \new_[12257]_ , \new_[12258]_ , \new_[12261]_ , \new_[12265]_ ,
    \new_[12266]_ , \new_[12267]_ , \new_[12270]_ , \new_[12274]_ ,
    \new_[12275]_ , \new_[12276]_ , \new_[12279]_ , \new_[12283]_ ,
    \new_[12284]_ , \new_[12285]_ , \new_[12288]_ , \new_[12292]_ ,
    \new_[12293]_ , \new_[12294]_ , \new_[12297]_ , \new_[12301]_ ,
    \new_[12302]_ , \new_[12303]_ , \new_[12306]_ , \new_[12310]_ ,
    \new_[12311]_ , \new_[12312]_ , \new_[12315]_ , \new_[12319]_ ,
    \new_[12320]_ , \new_[12321]_ , \new_[12324]_ , \new_[12328]_ ,
    \new_[12329]_ , \new_[12330]_ , \new_[12333]_ , \new_[12337]_ ,
    \new_[12338]_ , \new_[12339]_ , \new_[12342]_ , \new_[12346]_ ,
    \new_[12347]_ , \new_[12348]_ , \new_[12351]_ , \new_[12355]_ ,
    \new_[12356]_ , \new_[12357]_ , \new_[12360]_ , \new_[12364]_ ,
    \new_[12365]_ , \new_[12366]_ , \new_[12369]_ , \new_[12373]_ ,
    \new_[12374]_ , \new_[12375]_ , \new_[12378]_ , \new_[12382]_ ,
    \new_[12383]_ , \new_[12384]_ , \new_[12387]_ , \new_[12391]_ ,
    \new_[12392]_ , \new_[12393]_ , \new_[12396]_ , \new_[12400]_ ,
    \new_[12401]_ , \new_[12402]_ , \new_[12405]_ , \new_[12409]_ ,
    \new_[12410]_ , \new_[12411]_ , \new_[12414]_ , \new_[12418]_ ,
    \new_[12419]_ , \new_[12420]_ , \new_[12423]_ , \new_[12427]_ ,
    \new_[12428]_ , \new_[12429]_ , \new_[12432]_ , \new_[12436]_ ,
    \new_[12437]_ , \new_[12438]_ , \new_[12441]_ , \new_[12445]_ ,
    \new_[12446]_ , \new_[12447]_ , \new_[12450]_ , \new_[12454]_ ,
    \new_[12455]_ , \new_[12456]_ , \new_[12459]_ , \new_[12463]_ ,
    \new_[12464]_ , \new_[12465]_ , \new_[12468]_ , \new_[12472]_ ,
    \new_[12473]_ , \new_[12474]_ , \new_[12477]_ , \new_[12481]_ ,
    \new_[12482]_ , \new_[12483]_ , \new_[12486]_ , \new_[12490]_ ,
    \new_[12491]_ , \new_[12492]_ , \new_[12495]_ , \new_[12499]_ ,
    \new_[12500]_ , \new_[12501]_ , \new_[12504]_ , \new_[12508]_ ,
    \new_[12509]_ , \new_[12510]_ , \new_[12513]_ , \new_[12517]_ ,
    \new_[12518]_ , \new_[12519]_ , \new_[12522]_ , \new_[12526]_ ,
    \new_[12527]_ , \new_[12528]_ , \new_[12531]_ , \new_[12535]_ ,
    \new_[12536]_ , \new_[12537]_ , \new_[12540]_ , \new_[12544]_ ,
    \new_[12545]_ , \new_[12546]_ , \new_[12549]_ , \new_[12553]_ ,
    \new_[12554]_ , \new_[12555]_ , \new_[12558]_ , \new_[12562]_ ,
    \new_[12563]_ , \new_[12564]_ , \new_[12567]_ , \new_[12571]_ ,
    \new_[12572]_ , \new_[12573]_ , \new_[12576]_ , \new_[12580]_ ,
    \new_[12581]_ , \new_[12582]_ , \new_[12585]_ , \new_[12589]_ ,
    \new_[12590]_ , \new_[12591]_ , \new_[12594]_ , \new_[12598]_ ,
    \new_[12599]_ , \new_[12600]_ , \new_[12603]_ , \new_[12607]_ ,
    \new_[12608]_ , \new_[12609]_ , \new_[12612]_ , \new_[12616]_ ,
    \new_[12617]_ , \new_[12618]_ , \new_[12621]_ , \new_[12625]_ ,
    \new_[12626]_ , \new_[12627]_ , \new_[12630]_ , \new_[12634]_ ,
    \new_[12635]_ , \new_[12636]_ , \new_[12639]_ , \new_[12643]_ ,
    \new_[12644]_ , \new_[12645]_ , \new_[12648]_ , \new_[12652]_ ,
    \new_[12653]_ , \new_[12654]_ , \new_[12657]_ , \new_[12661]_ ,
    \new_[12662]_ , \new_[12663]_ , \new_[12666]_ , \new_[12670]_ ,
    \new_[12671]_ , \new_[12672]_ , \new_[12675]_ , \new_[12679]_ ,
    \new_[12680]_ , \new_[12681]_ , \new_[12684]_ , \new_[12688]_ ,
    \new_[12689]_ , \new_[12690]_ , \new_[12693]_ , \new_[12697]_ ,
    \new_[12698]_ , \new_[12699]_ , \new_[12702]_ , \new_[12706]_ ,
    \new_[12707]_ , \new_[12708]_ , \new_[12711]_ , \new_[12715]_ ,
    \new_[12716]_ , \new_[12717]_ , \new_[12720]_ , \new_[12724]_ ,
    \new_[12725]_ , \new_[12726]_ , \new_[12729]_ , \new_[12733]_ ,
    \new_[12734]_ , \new_[12735]_ , \new_[12738]_ , \new_[12742]_ ,
    \new_[12743]_ , \new_[12744]_ , \new_[12747]_ , \new_[12751]_ ,
    \new_[12752]_ , \new_[12753]_ , \new_[12756]_ , \new_[12760]_ ,
    \new_[12761]_ , \new_[12762]_ , \new_[12765]_ , \new_[12769]_ ,
    \new_[12770]_ , \new_[12771]_ , \new_[12774]_ , \new_[12778]_ ,
    \new_[12779]_ , \new_[12780]_ , \new_[12783]_ , \new_[12787]_ ,
    \new_[12788]_ , \new_[12789]_ , \new_[12792]_ , \new_[12796]_ ,
    \new_[12797]_ , \new_[12798]_ , \new_[12801]_ , \new_[12805]_ ,
    \new_[12806]_ , \new_[12807]_ , \new_[12810]_ , \new_[12814]_ ,
    \new_[12815]_ , \new_[12816]_ , \new_[12819]_ , \new_[12823]_ ,
    \new_[12824]_ , \new_[12825]_ , \new_[12828]_ , \new_[12832]_ ,
    \new_[12833]_ , \new_[12834]_ , \new_[12837]_ , \new_[12841]_ ,
    \new_[12842]_ , \new_[12843]_ , \new_[12846]_ , \new_[12850]_ ,
    \new_[12851]_ , \new_[12852]_ , \new_[12855]_ , \new_[12859]_ ,
    \new_[12860]_ , \new_[12861]_ , \new_[12864]_ , \new_[12868]_ ,
    \new_[12869]_ , \new_[12870]_ , \new_[12873]_ , \new_[12877]_ ,
    \new_[12878]_ , \new_[12879]_ , \new_[12882]_ , \new_[12886]_ ,
    \new_[12887]_ , \new_[12888]_ , \new_[12891]_ , \new_[12895]_ ,
    \new_[12896]_ , \new_[12897]_ , \new_[12900]_ , \new_[12904]_ ,
    \new_[12905]_ , \new_[12906]_ , \new_[12909]_ , \new_[12913]_ ,
    \new_[12914]_ , \new_[12915]_ , \new_[12918]_ , \new_[12922]_ ,
    \new_[12923]_ , \new_[12924]_ , \new_[12927]_ , \new_[12931]_ ,
    \new_[12932]_ , \new_[12933]_ , \new_[12936]_ , \new_[12940]_ ,
    \new_[12941]_ , \new_[12942]_ , \new_[12945]_ , \new_[12949]_ ,
    \new_[12950]_ , \new_[12951]_ , \new_[12954]_ , \new_[12958]_ ,
    \new_[12959]_ , \new_[12960]_ , \new_[12963]_ , \new_[12967]_ ,
    \new_[12968]_ , \new_[12969]_ , \new_[12972]_ , \new_[12976]_ ,
    \new_[12977]_ , \new_[12978]_ , \new_[12981]_ , \new_[12985]_ ,
    \new_[12986]_ , \new_[12987]_ , \new_[12990]_ , \new_[12994]_ ,
    \new_[12995]_ , \new_[12996]_ , \new_[12999]_ , \new_[13003]_ ,
    \new_[13004]_ , \new_[13005]_ , \new_[13008]_ , \new_[13012]_ ,
    \new_[13013]_ , \new_[13014]_ , \new_[13017]_ , \new_[13021]_ ,
    \new_[13022]_ , \new_[13023]_ , \new_[13026]_ , \new_[13030]_ ,
    \new_[13031]_ , \new_[13032]_ , \new_[13035]_ , \new_[13039]_ ,
    \new_[13040]_ , \new_[13041]_ , \new_[13044]_ , \new_[13048]_ ,
    \new_[13049]_ , \new_[13050]_ , \new_[13053]_ , \new_[13057]_ ,
    \new_[13058]_ , \new_[13059]_ , \new_[13062]_ , \new_[13066]_ ,
    \new_[13067]_ , \new_[13068]_ , \new_[13071]_ , \new_[13075]_ ,
    \new_[13076]_ , \new_[13077]_ , \new_[13080]_ , \new_[13084]_ ,
    \new_[13085]_ , \new_[13086]_ , \new_[13089]_ , \new_[13093]_ ,
    \new_[13094]_ , \new_[13095]_ , \new_[13098]_ , \new_[13102]_ ,
    \new_[13103]_ , \new_[13104]_ , \new_[13107]_ , \new_[13111]_ ,
    \new_[13112]_ , \new_[13113]_ , \new_[13116]_ , \new_[13120]_ ,
    \new_[13121]_ , \new_[13122]_ , \new_[13125]_ , \new_[13129]_ ,
    \new_[13130]_ , \new_[13131]_ , \new_[13134]_ , \new_[13138]_ ,
    \new_[13139]_ , \new_[13140]_ , \new_[13143]_ , \new_[13147]_ ,
    \new_[13148]_ , \new_[13149]_ , \new_[13152]_ , \new_[13156]_ ,
    \new_[13157]_ , \new_[13158]_ , \new_[13161]_ , \new_[13165]_ ,
    \new_[13166]_ , \new_[13167]_ , \new_[13170]_ , \new_[13174]_ ,
    \new_[13175]_ , \new_[13176]_ , \new_[13179]_ , \new_[13183]_ ,
    \new_[13184]_ , \new_[13185]_ , \new_[13188]_ , \new_[13192]_ ,
    \new_[13193]_ , \new_[13194]_ , \new_[13197]_ , \new_[13201]_ ,
    \new_[13202]_ , \new_[13203]_ , \new_[13206]_ , \new_[13210]_ ,
    \new_[13211]_ , \new_[13212]_ , \new_[13215]_ , \new_[13219]_ ,
    \new_[13220]_ , \new_[13221]_ , \new_[13224]_ , \new_[13228]_ ,
    \new_[13229]_ , \new_[13230]_ , \new_[13233]_ , \new_[13237]_ ,
    \new_[13238]_ , \new_[13239]_ , \new_[13242]_ , \new_[13246]_ ,
    \new_[13247]_ , \new_[13248]_ , \new_[13251]_ , \new_[13255]_ ,
    \new_[13256]_ , \new_[13257]_ , \new_[13260]_ , \new_[13264]_ ,
    \new_[13265]_ , \new_[13266]_ , \new_[13269]_ , \new_[13273]_ ,
    \new_[13274]_ , \new_[13275]_ , \new_[13278]_ , \new_[13282]_ ,
    \new_[13283]_ , \new_[13284]_ , \new_[13287]_ , \new_[13291]_ ,
    \new_[13292]_ , \new_[13293]_ , \new_[13296]_ , \new_[13300]_ ,
    \new_[13301]_ , \new_[13302]_ , \new_[13305]_ , \new_[13309]_ ,
    \new_[13310]_ , \new_[13311]_ , \new_[13314]_ , \new_[13318]_ ,
    \new_[13319]_ , \new_[13320]_ , \new_[13323]_ , \new_[13327]_ ,
    \new_[13328]_ , \new_[13329]_ , \new_[13332]_ , \new_[13336]_ ,
    \new_[13337]_ , \new_[13338]_ , \new_[13341]_ , \new_[13345]_ ,
    \new_[13346]_ , \new_[13347]_ , \new_[13350]_ , \new_[13354]_ ,
    \new_[13355]_ , \new_[13356]_ , \new_[13359]_ , \new_[13363]_ ,
    \new_[13364]_ , \new_[13365]_ , \new_[13368]_ , \new_[13372]_ ,
    \new_[13373]_ , \new_[13374]_ , \new_[13377]_ , \new_[13381]_ ,
    \new_[13382]_ , \new_[13383]_ , \new_[13386]_ , \new_[13390]_ ,
    \new_[13391]_ , \new_[13392]_ , \new_[13395]_ , \new_[13399]_ ,
    \new_[13400]_ , \new_[13401]_ , \new_[13404]_ , \new_[13408]_ ,
    \new_[13409]_ , \new_[13410]_ , \new_[13413]_ , \new_[13417]_ ,
    \new_[13418]_ , \new_[13419]_ , \new_[13422]_ , \new_[13426]_ ,
    \new_[13427]_ , \new_[13428]_ , \new_[13431]_ , \new_[13435]_ ,
    \new_[13436]_ , \new_[13437]_ , \new_[13440]_ , \new_[13444]_ ,
    \new_[13445]_ , \new_[13446]_ , \new_[13449]_ , \new_[13453]_ ,
    \new_[13454]_ , \new_[13455]_ , \new_[13458]_ , \new_[13462]_ ,
    \new_[13463]_ , \new_[13464]_ , \new_[13467]_ , \new_[13471]_ ,
    \new_[13472]_ , \new_[13473]_ , \new_[13476]_ , \new_[13480]_ ,
    \new_[13481]_ , \new_[13482]_ , \new_[13485]_ , \new_[13489]_ ,
    \new_[13490]_ , \new_[13491]_ , \new_[13494]_ , \new_[13498]_ ,
    \new_[13499]_ , \new_[13500]_ , \new_[13503]_ , \new_[13507]_ ,
    \new_[13508]_ , \new_[13509]_ , \new_[13512]_ , \new_[13516]_ ,
    \new_[13517]_ , \new_[13518]_ , \new_[13521]_ , \new_[13525]_ ,
    \new_[13526]_ , \new_[13527]_ , \new_[13530]_ , \new_[13534]_ ,
    \new_[13535]_ , \new_[13536]_ , \new_[13539]_ , \new_[13543]_ ,
    \new_[13544]_ , \new_[13545]_ , \new_[13548]_ , \new_[13552]_ ,
    \new_[13553]_ , \new_[13554]_ , \new_[13557]_ , \new_[13561]_ ,
    \new_[13562]_ , \new_[13563]_ , \new_[13566]_ , \new_[13570]_ ,
    \new_[13571]_ , \new_[13572]_ , \new_[13575]_ , \new_[13579]_ ,
    \new_[13580]_ , \new_[13581]_ , \new_[13584]_ , \new_[13588]_ ,
    \new_[13589]_ , \new_[13590]_ , \new_[13593]_ , \new_[13597]_ ,
    \new_[13598]_ , \new_[13599]_ , \new_[13602]_ , \new_[13606]_ ,
    \new_[13607]_ , \new_[13608]_ , \new_[13611]_ , \new_[13615]_ ,
    \new_[13616]_ , \new_[13617]_ , \new_[13620]_ , \new_[13624]_ ,
    \new_[13625]_ , \new_[13626]_ , \new_[13629]_ , \new_[13633]_ ,
    \new_[13634]_ , \new_[13635]_ , \new_[13638]_ , \new_[13642]_ ,
    \new_[13643]_ , \new_[13644]_ , \new_[13647]_ , \new_[13651]_ ,
    \new_[13652]_ , \new_[13653]_ , \new_[13656]_ , \new_[13660]_ ,
    \new_[13661]_ , \new_[13662]_ , \new_[13665]_ , \new_[13669]_ ,
    \new_[13670]_ , \new_[13671]_ , \new_[13674]_ , \new_[13678]_ ,
    \new_[13679]_ , \new_[13680]_ , \new_[13683]_ , \new_[13687]_ ,
    \new_[13688]_ , \new_[13689]_ , \new_[13692]_ , \new_[13696]_ ,
    \new_[13697]_ , \new_[13698]_ , \new_[13701]_ , \new_[13705]_ ,
    \new_[13706]_ , \new_[13707]_ , \new_[13710]_ , \new_[13714]_ ,
    \new_[13715]_ , \new_[13716]_ , \new_[13719]_ , \new_[13723]_ ,
    \new_[13724]_ , \new_[13725]_ , \new_[13728]_ , \new_[13732]_ ,
    \new_[13733]_ , \new_[13734]_ , \new_[13737]_ , \new_[13741]_ ,
    \new_[13742]_ , \new_[13743]_ , \new_[13746]_ , \new_[13750]_ ,
    \new_[13751]_ , \new_[13752]_ , \new_[13755]_ , \new_[13759]_ ,
    \new_[13760]_ , \new_[13761]_ , \new_[13764]_ , \new_[13768]_ ,
    \new_[13769]_ , \new_[13770]_ , \new_[13773]_ , \new_[13777]_ ,
    \new_[13778]_ , \new_[13779]_ , \new_[13782]_ , \new_[13786]_ ,
    \new_[13787]_ , \new_[13788]_ , \new_[13791]_ , \new_[13795]_ ,
    \new_[13796]_ , \new_[13797]_ , \new_[13800]_ , \new_[13804]_ ,
    \new_[13805]_ , \new_[13806]_ , \new_[13809]_ , \new_[13813]_ ,
    \new_[13814]_ , \new_[13815]_ , \new_[13818]_ , \new_[13822]_ ,
    \new_[13823]_ , \new_[13824]_ , \new_[13827]_ , \new_[13831]_ ,
    \new_[13832]_ , \new_[13833]_ , \new_[13836]_ , \new_[13840]_ ,
    \new_[13841]_ , \new_[13842]_ , \new_[13845]_ , \new_[13849]_ ,
    \new_[13850]_ , \new_[13851]_ , \new_[13854]_ , \new_[13858]_ ,
    \new_[13859]_ , \new_[13860]_ , \new_[13863]_ , \new_[13867]_ ,
    \new_[13868]_ , \new_[13869]_ , \new_[13872]_ , \new_[13876]_ ,
    \new_[13877]_ , \new_[13878]_ , \new_[13881]_ , \new_[13885]_ ,
    \new_[13886]_ , \new_[13887]_ , \new_[13890]_ , \new_[13894]_ ,
    \new_[13895]_ , \new_[13896]_ , \new_[13899]_ , \new_[13903]_ ,
    \new_[13904]_ , \new_[13905]_ , \new_[13908]_ , \new_[13912]_ ,
    \new_[13913]_ , \new_[13914]_ , \new_[13917]_ , \new_[13921]_ ,
    \new_[13922]_ , \new_[13923]_ , \new_[13926]_ , \new_[13930]_ ,
    \new_[13931]_ , \new_[13932]_ , \new_[13935]_ , \new_[13939]_ ,
    \new_[13940]_ , \new_[13941]_ , \new_[13944]_ , \new_[13948]_ ,
    \new_[13949]_ , \new_[13950]_ , \new_[13953]_ , \new_[13957]_ ,
    \new_[13958]_ , \new_[13959]_ , \new_[13962]_ , \new_[13966]_ ,
    \new_[13967]_ , \new_[13968]_ , \new_[13971]_ , \new_[13975]_ ,
    \new_[13976]_ , \new_[13977]_ , \new_[13980]_ , \new_[13984]_ ,
    \new_[13985]_ , \new_[13986]_ , \new_[13989]_ , \new_[13993]_ ,
    \new_[13994]_ , \new_[13995]_ , \new_[13998]_ , \new_[14002]_ ,
    \new_[14003]_ , \new_[14004]_ , \new_[14007]_ , \new_[14011]_ ,
    \new_[14012]_ , \new_[14013]_ , \new_[14016]_ , \new_[14020]_ ,
    \new_[14021]_ , \new_[14022]_ , \new_[14025]_ , \new_[14029]_ ,
    \new_[14030]_ , \new_[14031]_ , \new_[14034]_ , \new_[14038]_ ,
    \new_[14039]_ , \new_[14040]_ , \new_[14043]_ , \new_[14047]_ ,
    \new_[14048]_ , \new_[14049]_ , \new_[14052]_ , \new_[14056]_ ,
    \new_[14057]_ , \new_[14058]_ , \new_[14061]_ , \new_[14065]_ ,
    \new_[14066]_ , \new_[14067]_ , \new_[14070]_ , \new_[14074]_ ,
    \new_[14075]_ , \new_[14076]_ , \new_[14079]_ , \new_[14083]_ ,
    \new_[14084]_ , \new_[14085]_ , \new_[14088]_ , \new_[14092]_ ,
    \new_[14093]_ , \new_[14094]_ , \new_[14097]_ , \new_[14101]_ ,
    \new_[14102]_ , \new_[14103]_ , \new_[14106]_ , \new_[14110]_ ,
    \new_[14111]_ , \new_[14112]_ , \new_[14115]_ , \new_[14119]_ ,
    \new_[14120]_ , \new_[14121]_ , \new_[14124]_ , \new_[14128]_ ,
    \new_[14129]_ , \new_[14130]_ , \new_[14133]_ , \new_[14137]_ ,
    \new_[14138]_ , \new_[14139]_ , \new_[14142]_ , \new_[14146]_ ,
    \new_[14147]_ , \new_[14148]_ , \new_[14151]_ , \new_[14155]_ ,
    \new_[14156]_ , \new_[14157]_ , \new_[14160]_ , \new_[14164]_ ,
    \new_[14165]_ , \new_[14166]_ , \new_[14169]_ , \new_[14173]_ ,
    \new_[14174]_ , \new_[14175]_ , \new_[14178]_ , \new_[14182]_ ,
    \new_[14183]_ , \new_[14184]_ , \new_[14187]_ , \new_[14191]_ ,
    \new_[14192]_ , \new_[14193]_ , \new_[14196]_ , \new_[14200]_ ,
    \new_[14201]_ , \new_[14202]_ , \new_[14205]_ , \new_[14209]_ ,
    \new_[14210]_ , \new_[14211]_ , \new_[14214]_ , \new_[14218]_ ,
    \new_[14219]_ , \new_[14220]_ , \new_[14223]_ , \new_[14227]_ ,
    \new_[14228]_ , \new_[14229]_ , \new_[14232]_ , \new_[14236]_ ,
    \new_[14237]_ , \new_[14238]_ , \new_[14241]_ , \new_[14245]_ ,
    \new_[14246]_ , \new_[14247]_ , \new_[14250]_ , \new_[14254]_ ,
    \new_[14255]_ , \new_[14256]_ , \new_[14259]_ , \new_[14263]_ ,
    \new_[14264]_ , \new_[14265]_ , \new_[14268]_ , \new_[14272]_ ,
    \new_[14273]_ , \new_[14274]_ , \new_[14277]_ , \new_[14281]_ ,
    \new_[14282]_ , \new_[14283]_ , \new_[14286]_ , \new_[14290]_ ,
    \new_[14291]_ , \new_[14292]_ , \new_[14295]_ , \new_[14299]_ ,
    \new_[14300]_ , \new_[14301]_ , \new_[14304]_ , \new_[14308]_ ,
    \new_[14309]_ , \new_[14310]_ , \new_[14313]_ , \new_[14317]_ ,
    \new_[14318]_ , \new_[14319]_ , \new_[14322]_ , \new_[14326]_ ,
    \new_[14327]_ , \new_[14328]_ , \new_[14331]_ , \new_[14335]_ ,
    \new_[14336]_ , \new_[14337]_ , \new_[14340]_ , \new_[14344]_ ,
    \new_[14345]_ , \new_[14346]_ , \new_[14349]_ , \new_[14353]_ ,
    \new_[14354]_ , \new_[14355]_ , \new_[14358]_ , \new_[14362]_ ,
    \new_[14363]_ , \new_[14364]_ , \new_[14367]_ , \new_[14371]_ ,
    \new_[14372]_ , \new_[14373]_ , \new_[14376]_ , \new_[14380]_ ,
    \new_[14381]_ , \new_[14382]_ , \new_[14385]_ , \new_[14389]_ ,
    \new_[14390]_ , \new_[14391]_ , \new_[14394]_ , \new_[14398]_ ,
    \new_[14399]_ , \new_[14400]_ , \new_[14403]_ , \new_[14407]_ ,
    \new_[14408]_ , \new_[14409]_ , \new_[14412]_ , \new_[14416]_ ,
    \new_[14417]_ , \new_[14418]_ , \new_[14421]_ , \new_[14425]_ ,
    \new_[14426]_ , \new_[14427]_ , \new_[14430]_ , \new_[14434]_ ,
    \new_[14435]_ , \new_[14436]_ , \new_[14439]_ , \new_[14443]_ ,
    \new_[14444]_ , \new_[14445]_ , \new_[14448]_ , \new_[14452]_ ,
    \new_[14453]_ , \new_[14454]_ , \new_[14457]_ , \new_[14461]_ ,
    \new_[14462]_ , \new_[14463]_ , \new_[14466]_ , \new_[14470]_ ,
    \new_[14471]_ , \new_[14472]_ , \new_[14475]_ , \new_[14479]_ ,
    \new_[14480]_ , \new_[14481]_ , \new_[14484]_ , \new_[14488]_ ,
    \new_[14489]_ , \new_[14490]_ , \new_[14493]_ , \new_[14497]_ ,
    \new_[14498]_ , \new_[14499]_ , \new_[14502]_ , \new_[14506]_ ,
    \new_[14507]_ , \new_[14508]_ , \new_[14511]_ , \new_[14515]_ ,
    \new_[14516]_ , \new_[14517]_ , \new_[14520]_ , \new_[14524]_ ,
    \new_[14525]_ , \new_[14526]_ , \new_[14529]_ , \new_[14533]_ ,
    \new_[14534]_ , \new_[14535]_ , \new_[14538]_ , \new_[14542]_ ,
    \new_[14543]_ , \new_[14544]_ , \new_[14547]_ , \new_[14551]_ ,
    \new_[14552]_ , \new_[14553]_ , \new_[14556]_ , \new_[14560]_ ,
    \new_[14561]_ , \new_[14562]_ , \new_[14565]_ , \new_[14569]_ ,
    \new_[14570]_ , \new_[14571]_ , \new_[14574]_ , \new_[14578]_ ,
    \new_[14579]_ , \new_[14580]_ , \new_[14583]_ , \new_[14587]_ ,
    \new_[14588]_ , \new_[14589]_ , \new_[14592]_ , \new_[14596]_ ,
    \new_[14597]_ , \new_[14598]_ , \new_[14601]_ , \new_[14605]_ ,
    \new_[14606]_ , \new_[14607]_ , \new_[14610]_ , \new_[14614]_ ,
    \new_[14615]_ , \new_[14616]_ , \new_[14619]_ , \new_[14623]_ ,
    \new_[14624]_ , \new_[14625]_ , \new_[14628]_ , \new_[14632]_ ,
    \new_[14633]_ , \new_[14634]_ , \new_[14637]_ , \new_[14641]_ ,
    \new_[14642]_ , \new_[14643]_ , \new_[14646]_ , \new_[14650]_ ,
    \new_[14651]_ , \new_[14652]_ , \new_[14655]_ , \new_[14659]_ ,
    \new_[14660]_ , \new_[14661]_ , \new_[14664]_ , \new_[14668]_ ,
    \new_[14669]_ , \new_[14670]_ , \new_[14673]_ , \new_[14677]_ ,
    \new_[14678]_ , \new_[14679]_ , \new_[14682]_ , \new_[14686]_ ,
    \new_[14687]_ , \new_[14688]_ , \new_[14691]_ , \new_[14695]_ ,
    \new_[14696]_ , \new_[14697]_ , \new_[14700]_ , \new_[14704]_ ,
    \new_[14705]_ , \new_[14706]_ , \new_[14709]_ , \new_[14713]_ ,
    \new_[14714]_ , \new_[14715]_ , \new_[14718]_ , \new_[14722]_ ,
    \new_[14723]_ , \new_[14724]_ , \new_[14727]_ , \new_[14731]_ ,
    \new_[14732]_ , \new_[14733]_ , \new_[14736]_ , \new_[14740]_ ,
    \new_[14741]_ , \new_[14742]_ , \new_[14745]_ , \new_[14749]_ ,
    \new_[14750]_ , \new_[14751]_ , \new_[14754]_ , \new_[14758]_ ,
    \new_[14759]_ , \new_[14760]_ , \new_[14763]_ , \new_[14767]_ ,
    \new_[14768]_ , \new_[14769]_ , \new_[14772]_ , \new_[14776]_ ,
    \new_[14777]_ , \new_[14778]_ , \new_[14781]_ , \new_[14785]_ ,
    \new_[14786]_ , \new_[14787]_ , \new_[14790]_ , \new_[14794]_ ,
    \new_[14795]_ , \new_[14796]_ , \new_[14799]_ , \new_[14803]_ ,
    \new_[14804]_ , \new_[14805]_ , \new_[14808]_ , \new_[14812]_ ,
    \new_[14813]_ , \new_[14814]_ , \new_[14817]_ , \new_[14821]_ ,
    \new_[14822]_ , \new_[14823]_ , \new_[14826]_ , \new_[14830]_ ,
    \new_[14831]_ , \new_[14832]_ , \new_[14835]_ , \new_[14839]_ ,
    \new_[14840]_ , \new_[14841]_ , \new_[14844]_ , \new_[14848]_ ,
    \new_[14849]_ , \new_[14850]_ , \new_[14853]_ , \new_[14857]_ ,
    \new_[14858]_ , \new_[14859]_ , \new_[14862]_ , \new_[14866]_ ,
    \new_[14867]_ , \new_[14868]_ , \new_[14871]_ , \new_[14875]_ ,
    \new_[14876]_ , \new_[14877]_ , \new_[14880]_ , \new_[14884]_ ,
    \new_[14885]_ , \new_[14886]_ , \new_[14889]_ , \new_[14893]_ ,
    \new_[14894]_ , \new_[14895]_ , \new_[14898]_ , \new_[14902]_ ,
    \new_[14903]_ , \new_[14904]_ , \new_[14907]_ , \new_[14911]_ ,
    \new_[14912]_ , \new_[14913]_ , \new_[14916]_ , \new_[14920]_ ,
    \new_[14921]_ , \new_[14922]_ , \new_[14925]_ , \new_[14929]_ ,
    \new_[14930]_ , \new_[14931]_ , \new_[14934]_ , \new_[14938]_ ,
    \new_[14939]_ , \new_[14940]_ , \new_[14943]_ , \new_[14947]_ ,
    \new_[14948]_ , \new_[14949]_ , \new_[14952]_ , \new_[14956]_ ,
    \new_[14957]_ , \new_[14958]_ , \new_[14961]_ , \new_[14965]_ ,
    \new_[14966]_ , \new_[14967]_ , \new_[14970]_ , \new_[14974]_ ,
    \new_[14975]_ , \new_[14976]_ , \new_[14979]_ , \new_[14983]_ ,
    \new_[14984]_ , \new_[14985]_ , \new_[14988]_ , \new_[14992]_ ,
    \new_[14993]_ , \new_[14994]_ , \new_[14997]_ , \new_[15001]_ ,
    \new_[15002]_ , \new_[15003]_ , \new_[15006]_ , \new_[15010]_ ,
    \new_[15011]_ , \new_[15012]_ , \new_[15015]_ , \new_[15019]_ ,
    \new_[15020]_ , \new_[15021]_ , \new_[15024]_ , \new_[15028]_ ,
    \new_[15029]_ , \new_[15030]_ , \new_[15033]_ , \new_[15037]_ ,
    \new_[15038]_ , \new_[15039]_ , \new_[15042]_ , \new_[15046]_ ,
    \new_[15047]_ , \new_[15048]_ , \new_[15051]_ , \new_[15055]_ ,
    \new_[15056]_ , \new_[15057]_ , \new_[15060]_ , \new_[15064]_ ,
    \new_[15065]_ , \new_[15066]_ , \new_[15069]_ , \new_[15073]_ ,
    \new_[15074]_ , \new_[15075]_ , \new_[15078]_ , \new_[15082]_ ,
    \new_[15083]_ , \new_[15084]_ , \new_[15087]_ , \new_[15091]_ ,
    \new_[15092]_ , \new_[15093]_ , \new_[15096]_ , \new_[15100]_ ,
    \new_[15101]_ , \new_[15102]_ , \new_[15105]_ , \new_[15109]_ ,
    \new_[15110]_ , \new_[15111]_ , \new_[15114]_ , \new_[15118]_ ,
    \new_[15119]_ , \new_[15120]_ , \new_[15123]_ , \new_[15127]_ ,
    \new_[15128]_ , \new_[15129]_ , \new_[15132]_ , \new_[15136]_ ,
    \new_[15137]_ , \new_[15138]_ , \new_[15141]_ , \new_[15145]_ ,
    \new_[15146]_ , \new_[15147]_ , \new_[15150]_ , \new_[15154]_ ,
    \new_[15155]_ , \new_[15156]_ , \new_[15159]_ , \new_[15163]_ ,
    \new_[15164]_ , \new_[15165]_ , \new_[15168]_ , \new_[15172]_ ,
    \new_[15173]_ , \new_[15174]_ , \new_[15177]_ , \new_[15181]_ ,
    \new_[15182]_ , \new_[15183]_ , \new_[15186]_ , \new_[15190]_ ,
    \new_[15191]_ , \new_[15192]_ , \new_[15195]_ , \new_[15199]_ ,
    \new_[15200]_ , \new_[15201]_ , \new_[15204]_ , \new_[15208]_ ,
    \new_[15209]_ , \new_[15210]_ , \new_[15213]_ , \new_[15217]_ ,
    \new_[15218]_ , \new_[15219]_ , \new_[15222]_ , \new_[15226]_ ,
    \new_[15227]_ , \new_[15228]_ , \new_[15231]_ , \new_[15235]_ ,
    \new_[15236]_ , \new_[15237]_ , \new_[15240]_ , \new_[15244]_ ,
    \new_[15245]_ , \new_[15246]_ , \new_[15249]_ , \new_[15253]_ ,
    \new_[15254]_ , \new_[15255]_ , \new_[15258]_ , \new_[15262]_ ,
    \new_[15263]_ , \new_[15264]_ , \new_[15267]_ , \new_[15271]_ ,
    \new_[15272]_ , \new_[15273]_ , \new_[15276]_ , \new_[15280]_ ,
    \new_[15281]_ , \new_[15282]_ , \new_[15285]_ , \new_[15289]_ ,
    \new_[15290]_ , \new_[15291]_ , \new_[15294]_ , \new_[15298]_ ,
    \new_[15299]_ , \new_[15300]_ , \new_[15303]_ , \new_[15307]_ ,
    \new_[15308]_ , \new_[15309]_ , \new_[15312]_ , \new_[15316]_ ,
    \new_[15317]_ , \new_[15318]_ , \new_[15321]_ , \new_[15325]_ ,
    \new_[15326]_ , \new_[15327]_ , \new_[15330]_ , \new_[15334]_ ,
    \new_[15335]_ , \new_[15336]_ , \new_[15339]_ , \new_[15343]_ ,
    \new_[15344]_ , \new_[15345]_ , \new_[15348]_ , \new_[15352]_ ,
    \new_[15353]_ , \new_[15354]_ , \new_[15357]_ , \new_[15361]_ ,
    \new_[15362]_ , \new_[15363]_ , \new_[15366]_ , \new_[15370]_ ,
    \new_[15371]_ , \new_[15372]_ , \new_[15375]_ , \new_[15379]_ ,
    \new_[15380]_ , \new_[15381]_ , \new_[15384]_ , \new_[15388]_ ,
    \new_[15389]_ , \new_[15390]_ , \new_[15393]_ , \new_[15397]_ ,
    \new_[15398]_ , \new_[15399]_ , \new_[15402]_ , \new_[15406]_ ,
    \new_[15407]_ , \new_[15408]_ , \new_[15411]_ , \new_[15415]_ ,
    \new_[15416]_ , \new_[15417]_ , \new_[15420]_ , \new_[15424]_ ,
    \new_[15425]_ , \new_[15426]_ , \new_[15429]_ , \new_[15433]_ ,
    \new_[15434]_ , \new_[15435]_ , \new_[15438]_ , \new_[15442]_ ,
    \new_[15443]_ , \new_[15444]_ , \new_[15447]_ , \new_[15451]_ ,
    \new_[15452]_ , \new_[15453]_ , \new_[15456]_ , \new_[15460]_ ,
    \new_[15461]_ , \new_[15462]_ , \new_[15465]_ , \new_[15469]_ ,
    \new_[15470]_ , \new_[15471]_ , \new_[15474]_ , \new_[15478]_ ,
    \new_[15479]_ , \new_[15480]_ , \new_[15483]_ , \new_[15487]_ ,
    \new_[15488]_ , \new_[15489]_ , \new_[15492]_ , \new_[15496]_ ,
    \new_[15497]_ , \new_[15498]_ , \new_[15501]_ , \new_[15505]_ ,
    \new_[15506]_ , \new_[15507]_ , \new_[15510]_ , \new_[15514]_ ,
    \new_[15515]_ , \new_[15516]_ , \new_[15519]_ , \new_[15523]_ ,
    \new_[15524]_ , \new_[15525]_ , \new_[15528]_ , \new_[15532]_ ,
    \new_[15533]_ , \new_[15534]_ , \new_[15537]_ , \new_[15541]_ ,
    \new_[15542]_ , \new_[15543]_ , \new_[15546]_ , \new_[15550]_ ,
    \new_[15551]_ , \new_[15552]_ , \new_[15555]_ , \new_[15559]_ ,
    \new_[15560]_ , \new_[15561]_ , \new_[15564]_ , \new_[15568]_ ,
    \new_[15569]_ , \new_[15570]_ , \new_[15573]_ , \new_[15577]_ ,
    \new_[15578]_ , \new_[15579]_ , \new_[15582]_ , \new_[15586]_ ,
    \new_[15587]_ , \new_[15588]_ , \new_[15591]_ , \new_[15595]_ ,
    \new_[15596]_ , \new_[15597]_ , \new_[15600]_ , \new_[15604]_ ,
    \new_[15605]_ , \new_[15606]_ , \new_[15609]_ , \new_[15613]_ ,
    \new_[15614]_ , \new_[15615]_ , \new_[15618]_ , \new_[15622]_ ,
    \new_[15623]_ , \new_[15624]_ , \new_[15627]_ , \new_[15631]_ ,
    \new_[15632]_ , \new_[15633]_ , \new_[15636]_ , \new_[15640]_ ,
    \new_[15641]_ , \new_[15642]_ , \new_[15645]_ , \new_[15649]_ ,
    \new_[15650]_ , \new_[15651]_ , \new_[15654]_ , \new_[15658]_ ,
    \new_[15659]_ , \new_[15660]_ , \new_[15663]_ , \new_[15667]_ ,
    \new_[15668]_ , \new_[15669]_ , \new_[15672]_ , \new_[15676]_ ,
    \new_[15677]_ , \new_[15678]_ , \new_[15681]_ , \new_[15685]_ ,
    \new_[15686]_ , \new_[15687]_ , \new_[15690]_ , \new_[15694]_ ,
    \new_[15695]_ , \new_[15696]_ , \new_[15699]_ , \new_[15703]_ ,
    \new_[15704]_ , \new_[15705]_ , \new_[15708]_ , \new_[15712]_ ,
    \new_[15713]_ , \new_[15714]_ , \new_[15717]_ , \new_[15721]_ ,
    \new_[15722]_ , \new_[15723]_ , \new_[15726]_ , \new_[15730]_ ,
    \new_[15731]_ , \new_[15732]_ , \new_[15735]_ , \new_[15739]_ ,
    \new_[15740]_ , \new_[15741]_ , \new_[15744]_ , \new_[15748]_ ,
    \new_[15749]_ , \new_[15750]_ , \new_[15753]_ , \new_[15757]_ ,
    \new_[15758]_ , \new_[15759]_ , \new_[15762]_ , \new_[15766]_ ,
    \new_[15767]_ , \new_[15768]_ , \new_[15771]_ , \new_[15775]_ ,
    \new_[15776]_ , \new_[15777]_ , \new_[15780]_ , \new_[15784]_ ,
    \new_[15785]_ , \new_[15786]_ , \new_[15789]_ , \new_[15793]_ ,
    \new_[15794]_ , \new_[15795]_ , \new_[15798]_ , \new_[15802]_ ,
    \new_[15803]_ , \new_[15804]_ , \new_[15807]_ , \new_[15811]_ ,
    \new_[15812]_ , \new_[15813]_ , \new_[15816]_ , \new_[15820]_ ,
    \new_[15821]_ , \new_[15822]_ , \new_[15825]_ , \new_[15829]_ ,
    \new_[15830]_ , \new_[15831]_ , \new_[15834]_ , \new_[15838]_ ,
    \new_[15839]_ , \new_[15840]_ , \new_[15843]_ , \new_[15847]_ ,
    \new_[15848]_ , \new_[15849]_ , \new_[15852]_ , \new_[15856]_ ,
    \new_[15857]_ , \new_[15858]_ , \new_[15861]_ , \new_[15865]_ ,
    \new_[15866]_ , \new_[15867]_ , \new_[15870]_ , \new_[15874]_ ,
    \new_[15875]_ , \new_[15876]_ , \new_[15879]_ , \new_[15883]_ ,
    \new_[15884]_ , \new_[15885]_ , \new_[15888]_ , \new_[15892]_ ,
    \new_[15893]_ , \new_[15894]_ , \new_[15897]_ , \new_[15901]_ ,
    \new_[15902]_ , \new_[15903]_ , \new_[15906]_ , \new_[15910]_ ,
    \new_[15911]_ , \new_[15912]_ , \new_[15915]_ , \new_[15919]_ ,
    \new_[15920]_ , \new_[15921]_ , \new_[15924]_ , \new_[15928]_ ,
    \new_[15929]_ , \new_[15930]_ , \new_[15933]_ , \new_[15937]_ ,
    \new_[15938]_ , \new_[15939]_ , \new_[15942]_ , \new_[15946]_ ,
    \new_[15947]_ , \new_[15948]_ , \new_[15951]_ , \new_[15955]_ ,
    \new_[15956]_ , \new_[15957]_ , \new_[15960]_ , \new_[15964]_ ,
    \new_[15965]_ , \new_[15966]_ , \new_[15969]_ , \new_[15973]_ ,
    \new_[15974]_ , \new_[15975]_ , \new_[15978]_ , \new_[15982]_ ,
    \new_[15983]_ , \new_[15984]_ , \new_[15987]_ , \new_[15991]_ ,
    \new_[15992]_ , \new_[15993]_ , \new_[15996]_ , \new_[16000]_ ,
    \new_[16001]_ , \new_[16002]_ , \new_[16005]_ , \new_[16009]_ ,
    \new_[16010]_ , \new_[16011]_ , \new_[16014]_ , \new_[16018]_ ,
    \new_[16019]_ , \new_[16020]_ , \new_[16023]_ , \new_[16027]_ ,
    \new_[16028]_ , \new_[16029]_ , \new_[16032]_ , \new_[16036]_ ,
    \new_[16037]_ , \new_[16038]_ , \new_[16041]_ , \new_[16045]_ ,
    \new_[16046]_ , \new_[16047]_ , \new_[16051]_ , \new_[16052]_ ,
    \new_[16056]_ , \new_[16057]_ , \new_[16058]_ , \new_[16061]_ ,
    \new_[16065]_ , \new_[16066]_ , \new_[16067]_ , \new_[16071]_ ,
    \new_[16072]_ , \new_[16076]_ , \new_[16077]_ , \new_[16078]_ ,
    \new_[16081]_ , \new_[16085]_ , \new_[16086]_ , \new_[16087]_ ,
    \new_[16091]_ , \new_[16092]_ , \new_[16096]_ , \new_[16097]_ ,
    \new_[16098]_ , \new_[16101]_ , \new_[16105]_ , \new_[16106]_ ,
    \new_[16107]_ , \new_[16111]_ , \new_[16112]_ , \new_[16116]_ ,
    \new_[16117]_ , \new_[16118]_ , \new_[16121]_ , \new_[16125]_ ,
    \new_[16126]_ , \new_[16127]_ , \new_[16131]_ , \new_[16132]_ ,
    \new_[16136]_ , \new_[16137]_ , \new_[16138]_ , \new_[16141]_ ,
    \new_[16145]_ , \new_[16146]_ , \new_[16147]_ , \new_[16151]_ ,
    \new_[16152]_ , \new_[16156]_ , \new_[16157]_ , \new_[16158]_ ,
    \new_[16161]_ , \new_[16165]_ , \new_[16166]_ , \new_[16167]_ ,
    \new_[16171]_ , \new_[16172]_ , \new_[16176]_ , \new_[16177]_ ,
    \new_[16178]_ , \new_[16181]_ , \new_[16185]_ , \new_[16186]_ ,
    \new_[16187]_ , \new_[16191]_ , \new_[16192]_ , \new_[16196]_ ,
    \new_[16197]_ , \new_[16198]_ , \new_[16201]_ , \new_[16205]_ ,
    \new_[16206]_ , \new_[16207]_ , \new_[16211]_ , \new_[16212]_ ,
    \new_[16216]_ , \new_[16217]_ , \new_[16218]_ , \new_[16221]_ ,
    \new_[16225]_ , \new_[16226]_ , \new_[16227]_ , \new_[16231]_ ,
    \new_[16232]_ , \new_[16236]_ , \new_[16237]_ , \new_[16238]_ ,
    \new_[16241]_ , \new_[16245]_ , \new_[16246]_ , \new_[16247]_ ,
    \new_[16251]_ , \new_[16252]_ , \new_[16256]_ , \new_[16257]_ ,
    \new_[16258]_ , \new_[16261]_ , \new_[16265]_ , \new_[16266]_ ,
    \new_[16267]_ , \new_[16271]_ , \new_[16272]_ , \new_[16276]_ ,
    \new_[16277]_ , \new_[16278]_ , \new_[16281]_ , \new_[16285]_ ,
    \new_[16286]_ , \new_[16287]_ , \new_[16291]_ , \new_[16292]_ ,
    \new_[16296]_ , \new_[16297]_ , \new_[16298]_ , \new_[16301]_ ,
    \new_[16305]_ , \new_[16306]_ , \new_[16307]_ , \new_[16311]_ ,
    \new_[16312]_ , \new_[16316]_ , \new_[16317]_ , \new_[16318]_ ,
    \new_[16321]_ , \new_[16325]_ , \new_[16326]_ , \new_[16327]_ ,
    \new_[16331]_ , \new_[16332]_ , \new_[16336]_ , \new_[16337]_ ,
    \new_[16338]_ , \new_[16341]_ , \new_[16345]_ , \new_[16346]_ ,
    \new_[16347]_ , \new_[16351]_ , \new_[16352]_ , \new_[16356]_ ,
    \new_[16357]_ , \new_[16358]_ , \new_[16361]_ , \new_[16365]_ ,
    \new_[16366]_ , \new_[16367]_ , \new_[16371]_ , \new_[16372]_ ,
    \new_[16376]_ , \new_[16377]_ , \new_[16378]_ , \new_[16381]_ ,
    \new_[16385]_ , \new_[16386]_ , \new_[16387]_ , \new_[16391]_ ,
    \new_[16392]_ , \new_[16396]_ , \new_[16397]_ , \new_[16398]_ ,
    \new_[16401]_ , \new_[16405]_ , \new_[16406]_ , \new_[16407]_ ,
    \new_[16411]_ , \new_[16412]_ , \new_[16416]_ , \new_[16417]_ ,
    \new_[16418]_ , \new_[16421]_ , \new_[16425]_ , \new_[16426]_ ,
    \new_[16427]_ , \new_[16431]_ , \new_[16432]_ , \new_[16436]_ ,
    \new_[16437]_ , \new_[16438]_ , \new_[16441]_ , \new_[16445]_ ,
    \new_[16446]_ , \new_[16447]_ , \new_[16451]_ , \new_[16452]_ ,
    \new_[16456]_ , \new_[16457]_ , \new_[16458]_ , \new_[16461]_ ,
    \new_[16465]_ , \new_[16466]_ , \new_[16467]_ , \new_[16471]_ ,
    \new_[16472]_ , \new_[16476]_ , \new_[16477]_ , \new_[16478]_ ,
    \new_[16481]_ , \new_[16485]_ , \new_[16486]_ , \new_[16487]_ ,
    \new_[16491]_ , \new_[16492]_ , \new_[16496]_ , \new_[16497]_ ,
    \new_[16498]_ , \new_[16501]_ , \new_[16505]_ , \new_[16506]_ ,
    \new_[16507]_ , \new_[16511]_ , \new_[16512]_ , \new_[16516]_ ,
    \new_[16517]_ , \new_[16518]_ , \new_[16521]_ , \new_[16525]_ ,
    \new_[16526]_ , \new_[16527]_ , \new_[16531]_ , \new_[16532]_ ,
    \new_[16536]_ , \new_[16537]_ , \new_[16538]_ , \new_[16541]_ ,
    \new_[16545]_ , \new_[16546]_ , \new_[16547]_ , \new_[16551]_ ,
    \new_[16552]_ , \new_[16556]_ , \new_[16557]_ , \new_[16558]_ ,
    \new_[16561]_ , \new_[16565]_ , \new_[16566]_ , \new_[16567]_ ,
    \new_[16571]_ , \new_[16572]_ , \new_[16576]_ , \new_[16577]_ ,
    \new_[16578]_ , \new_[16581]_ , \new_[16585]_ , \new_[16586]_ ,
    \new_[16587]_ , \new_[16591]_ , \new_[16592]_ , \new_[16596]_ ,
    \new_[16597]_ , \new_[16598]_ , \new_[16601]_ , \new_[16605]_ ,
    \new_[16606]_ , \new_[16607]_ , \new_[16611]_ , \new_[16612]_ ,
    \new_[16616]_ , \new_[16617]_ , \new_[16618]_ , \new_[16621]_ ,
    \new_[16625]_ , \new_[16626]_ , \new_[16627]_ , \new_[16631]_ ,
    \new_[16632]_ , \new_[16636]_ , \new_[16637]_ , \new_[16638]_ ,
    \new_[16641]_ , \new_[16645]_ , \new_[16646]_ , \new_[16647]_ ,
    \new_[16651]_ , \new_[16652]_ , \new_[16656]_ , \new_[16657]_ ,
    \new_[16658]_ , \new_[16661]_ , \new_[16665]_ , \new_[16666]_ ,
    \new_[16667]_ , \new_[16671]_ , \new_[16672]_ , \new_[16676]_ ,
    \new_[16677]_ , \new_[16678]_ , \new_[16681]_ , \new_[16685]_ ,
    \new_[16686]_ , \new_[16687]_ , \new_[16691]_ , \new_[16692]_ ,
    \new_[16696]_ , \new_[16697]_ , \new_[16698]_ , \new_[16701]_ ,
    \new_[16705]_ , \new_[16706]_ , \new_[16707]_ , \new_[16711]_ ,
    \new_[16712]_ , \new_[16716]_ , \new_[16717]_ , \new_[16718]_ ,
    \new_[16721]_ , \new_[16725]_ , \new_[16726]_ , \new_[16727]_ ,
    \new_[16731]_ , \new_[16732]_ , \new_[16736]_ , \new_[16737]_ ,
    \new_[16738]_ , \new_[16741]_ , \new_[16745]_ , \new_[16746]_ ,
    \new_[16747]_ , \new_[16751]_ , \new_[16752]_ , \new_[16756]_ ,
    \new_[16757]_ , \new_[16758]_ , \new_[16761]_ , \new_[16765]_ ,
    \new_[16766]_ , \new_[16767]_ , \new_[16771]_ , \new_[16772]_ ,
    \new_[16776]_ , \new_[16777]_ , \new_[16778]_ , \new_[16781]_ ,
    \new_[16785]_ , \new_[16786]_ , \new_[16787]_ , \new_[16791]_ ,
    \new_[16792]_ , \new_[16796]_ , \new_[16797]_ , \new_[16798]_ ,
    \new_[16801]_ , \new_[16805]_ , \new_[16806]_ , \new_[16807]_ ,
    \new_[16811]_ , \new_[16812]_ , \new_[16816]_ , \new_[16817]_ ,
    \new_[16818]_ , \new_[16821]_ , \new_[16825]_ , \new_[16826]_ ,
    \new_[16827]_ , \new_[16831]_ , \new_[16832]_ , \new_[16836]_ ,
    \new_[16837]_ , \new_[16838]_ , \new_[16841]_ , \new_[16845]_ ,
    \new_[16846]_ , \new_[16847]_ , \new_[16851]_ , \new_[16852]_ ,
    \new_[16856]_ , \new_[16857]_ , \new_[16858]_ , \new_[16861]_ ,
    \new_[16865]_ , \new_[16866]_ , \new_[16867]_ , \new_[16871]_ ,
    \new_[16872]_ , \new_[16876]_ , \new_[16877]_ , \new_[16878]_ ,
    \new_[16881]_ , \new_[16885]_ , \new_[16886]_ , \new_[16887]_ ,
    \new_[16891]_ , \new_[16892]_ , \new_[16896]_ , \new_[16897]_ ,
    \new_[16898]_ , \new_[16901]_ , \new_[16905]_ , \new_[16906]_ ,
    \new_[16907]_ , \new_[16911]_ , \new_[16912]_ , \new_[16916]_ ,
    \new_[16917]_ , \new_[16918]_ , \new_[16921]_ , \new_[16925]_ ,
    \new_[16926]_ , \new_[16927]_ , \new_[16931]_ , \new_[16932]_ ,
    \new_[16936]_ , \new_[16937]_ , \new_[16938]_ , \new_[16941]_ ,
    \new_[16945]_ , \new_[16946]_ , \new_[16947]_ , \new_[16951]_ ,
    \new_[16952]_ , \new_[16956]_ , \new_[16957]_ , \new_[16958]_ ,
    \new_[16961]_ , \new_[16965]_ , \new_[16966]_ , \new_[16967]_ ,
    \new_[16971]_ , \new_[16972]_ , \new_[16976]_ , \new_[16977]_ ,
    \new_[16978]_ , \new_[16981]_ , \new_[16985]_ , \new_[16986]_ ,
    \new_[16987]_ , \new_[16991]_ , \new_[16992]_ , \new_[16996]_ ,
    \new_[16997]_ , \new_[16998]_ , \new_[17001]_ , \new_[17005]_ ,
    \new_[17006]_ , \new_[17007]_ , \new_[17011]_ , \new_[17012]_ ,
    \new_[17016]_ , \new_[17017]_ , \new_[17018]_ , \new_[17021]_ ,
    \new_[17025]_ , \new_[17026]_ , \new_[17027]_ , \new_[17031]_ ,
    \new_[17032]_ , \new_[17036]_ , \new_[17037]_ , \new_[17038]_ ,
    \new_[17041]_ , \new_[17045]_ , \new_[17046]_ , \new_[17047]_ ,
    \new_[17051]_ , \new_[17052]_ , \new_[17056]_ , \new_[17057]_ ,
    \new_[17058]_ , \new_[17061]_ , \new_[17065]_ , \new_[17066]_ ,
    \new_[17067]_ , \new_[17071]_ , \new_[17072]_ , \new_[17076]_ ,
    \new_[17077]_ , \new_[17078]_ , \new_[17081]_ , \new_[17085]_ ,
    \new_[17086]_ , \new_[17087]_ , \new_[17091]_ , \new_[17092]_ ,
    \new_[17096]_ , \new_[17097]_ , \new_[17098]_ , \new_[17101]_ ,
    \new_[17105]_ , \new_[17106]_ , \new_[17107]_ , \new_[17111]_ ,
    \new_[17112]_ , \new_[17116]_ , \new_[17117]_ , \new_[17118]_ ,
    \new_[17121]_ , \new_[17125]_ , \new_[17126]_ , \new_[17127]_ ,
    \new_[17131]_ , \new_[17132]_ , \new_[17136]_ , \new_[17137]_ ,
    \new_[17138]_ , \new_[17141]_ , \new_[17145]_ , \new_[17146]_ ,
    \new_[17147]_ , \new_[17151]_ , \new_[17152]_ , \new_[17156]_ ,
    \new_[17157]_ , \new_[17158]_ , \new_[17161]_ , \new_[17165]_ ,
    \new_[17166]_ , \new_[17167]_ , \new_[17171]_ , \new_[17172]_ ,
    \new_[17176]_ , \new_[17177]_ , \new_[17178]_ , \new_[17181]_ ,
    \new_[17185]_ , \new_[17186]_ , \new_[17187]_ , \new_[17191]_ ,
    \new_[17192]_ , \new_[17196]_ , \new_[17197]_ , \new_[17198]_ ,
    \new_[17201]_ , \new_[17205]_ , \new_[17206]_ , \new_[17207]_ ,
    \new_[17211]_ , \new_[17212]_ , \new_[17216]_ , \new_[17217]_ ,
    \new_[17218]_ , \new_[17221]_ , \new_[17225]_ , \new_[17226]_ ,
    \new_[17227]_ , \new_[17231]_ , \new_[17232]_ , \new_[17236]_ ,
    \new_[17237]_ , \new_[17238]_ , \new_[17241]_ , \new_[17245]_ ,
    \new_[17246]_ , \new_[17247]_ , \new_[17251]_ , \new_[17252]_ ,
    \new_[17256]_ , \new_[17257]_ , \new_[17258]_ , \new_[17261]_ ,
    \new_[17265]_ , \new_[17266]_ , \new_[17267]_ , \new_[17271]_ ,
    \new_[17272]_ , \new_[17276]_ , \new_[17277]_ , \new_[17278]_ ,
    \new_[17281]_ , \new_[17285]_ , \new_[17286]_ , \new_[17287]_ ,
    \new_[17291]_ , \new_[17292]_ , \new_[17296]_ , \new_[17297]_ ,
    \new_[17298]_ , \new_[17301]_ , \new_[17305]_ , \new_[17306]_ ,
    \new_[17307]_ , \new_[17311]_ , \new_[17312]_ , \new_[17316]_ ,
    \new_[17317]_ , \new_[17318]_ , \new_[17321]_ , \new_[17325]_ ,
    \new_[17326]_ , \new_[17327]_ , \new_[17331]_ , \new_[17332]_ ,
    \new_[17336]_ , \new_[17337]_ , \new_[17338]_ , \new_[17341]_ ,
    \new_[17345]_ , \new_[17346]_ , \new_[17347]_ , \new_[17351]_ ,
    \new_[17352]_ , \new_[17356]_ , \new_[17357]_ , \new_[17358]_ ,
    \new_[17361]_ , \new_[17365]_ , \new_[17366]_ , \new_[17367]_ ,
    \new_[17371]_ , \new_[17372]_ , \new_[17376]_ , \new_[17377]_ ,
    \new_[17378]_ , \new_[17381]_ , \new_[17385]_ , \new_[17386]_ ,
    \new_[17387]_ , \new_[17391]_ , \new_[17392]_ , \new_[17396]_ ,
    \new_[17397]_ , \new_[17398]_ , \new_[17401]_ , \new_[17405]_ ,
    \new_[17406]_ , \new_[17407]_ , \new_[17411]_ , \new_[17412]_ ,
    \new_[17416]_ , \new_[17417]_ , \new_[17418]_ , \new_[17421]_ ,
    \new_[17425]_ , \new_[17426]_ , \new_[17427]_ , \new_[17431]_ ,
    \new_[17432]_ , \new_[17436]_ , \new_[17437]_ , \new_[17438]_ ,
    \new_[17441]_ , \new_[17445]_ , \new_[17446]_ , \new_[17447]_ ,
    \new_[17451]_ , \new_[17452]_ , \new_[17456]_ , \new_[17457]_ ,
    \new_[17458]_ , \new_[17461]_ , \new_[17465]_ , \new_[17466]_ ,
    \new_[17467]_ , \new_[17471]_ , \new_[17472]_ , \new_[17476]_ ,
    \new_[17477]_ , \new_[17478]_ , \new_[17481]_ , \new_[17485]_ ,
    \new_[17486]_ , \new_[17487]_ , \new_[17491]_ , \new_[17492]_ ,
    \new_[17496]_ , \new_[17497]_ , \new_[17498]_ , \new_[17501]_ ,
    \new_[17505]_ , \new_[17506]_ , \new_[17507]_ , \new_[17511]_ ,
    \new_[17512]_ , \new_[17516]_ , \new_[17517]_ , \new_[17518]_ ,
    \new_[17521]_ , \new_[17525]_ , \new_[17526]_ , \new_[17527]_ ,
    \new_[17531]_ , \new_[17532]_ , \new_[17536]_ , \new_[17537]_ ,
    \new_[17538]_ , \new_[17541]_ , \new_[17545]_ , \new_[17546]_ ,
    \new_[17547]_ , \new_[17551]_ , \new_[17552]_ , \new_[17556]_ ,
    \new_[17557]_ , \new_[17558]_ , \new_[17561]_ , \new_[17565]_ ,
    \new_[17566]_ , \new_[17567]_ , \new_[17571]_ , \new_[17572]_ ,
    \new_[17576]_ , \new_[17577]_ , \new_[17578]_ , \new_[17581]_ ,
    \new_[17585]_ , \new_[17586]_ , \new_[17587]_ , \new_[17591]_ ,
    \new_[17592]_ , \new_[17596]_ , \new_[17597]_ , \new_[17598]_ ,
    \new_[17601]_ , \new_[17605]_ , \new_[17606]_ , \new_[17607]_ ,
    \new_[17611]_ , \new_[17612]_ , \new_[17616]_ , \new_[17617]_ ,
    \new_[17618]_ , \new_[17621]_ , \new_[17625]_ , \new_[17626]_ ,
    \new_[17627]_ , \new_[17631]_ , \new_[17632]_ , \new_[17636]_ ,
    \new_[17637]_ , \new_[17638]_ , \new_[17641]_ , \new_[17645]_ ,
    \new_[17646]_ , \new_[17647]_ , \new_[17651]_ , \new_[17652]_ ,
    \new_[17656]_ , \new_[17657]_ , \new_[17658]_ , \new_[17661]_ ,
    \new_[17665]_ , \new_[17666]_ , \new_[17667]_ , \new_[17671]_ ,
    \new_[17672]_ , \new_[17676]_ , \new_[17677]_ , \new_[17678]_ ,
    \new_[17681]_ , \new_[17685]_ , \new_[17686]_ , \new_[17687]_ ,
    \new_[17691]_ , \new_[17692]_ , \new_[17696]_ , \new_[17697]_ ,
    \new_[17698]_ , \new_[17701]_ , \new_[17705]_ , \new_[17706]_ ,
    \new_[17707]_ , \new_[17711]_ , \new_[17712]_ , \new_[17716]_ ,
    \new_[17717]_ , \new_[17718]_ , \new_[17721]_ , \new_[17725]_ ,
    \new_[17726]_ , \new_[17727]_ , \new_[17731]_ , \new_[17732]_ ,
    \new_[17736]_ , \new_[17737]_ , \new_[17738]_ , \new_[17741]_ ,
    \new_[17745]_ , \new_[17746]_ , \new_[17747]_ , \new_[17751]_ ,
    \new_[17752]_ , \new_[17756]_ , \new_[17757]_ , \new_[17758]_ ,
    \new_[17761]_ , \new_[17765]_ , \new_[17766]_ , \new_[17767]_ ,
    \new_[17771]_ , \new_[17772]_ , \new_[17776]_ , \new_[17777]_ ,
    \new_[17778]_ , \new_[17781]_ , \new_[17785]_ , \new_[17786]_ ,
    \new_[17787]_ , \new_[17791]_ , \new_[17792]_ , \new_[17796]_ ,
    \new_[17797]_ , \new_[17798]_ , \new_[17801]_ , \new_[17805]_ ,
    \new_[17806]_ , \new_[17807]_ , \new_[17811]_ , \new_[17812]_ ,
    \new_[17816]_ , \new_[17817]_ , \new_[17818]_ , \new_[17821]_ ,
    \new_[17825]_ , \new_[17826]_ , \new_[17827]_ , \new_[17831]_ ,
    \new_[17832]_ , \new_[17836]_ , \new_[17837]_ , \new_[17838]_ ,
    \new_[17841]_ , \new_[17845]_ , \new_[17846]_ , \new_[17847]_ ,
    \new_[17851]_ , \new_[17852]_ , \new_[17856]_ , \new_[17857]_ ,
    \new_[17858]_ , \new_[17861]_ , \new_[17865]_ , \new_[17866]_ ,
    \new_[17867]_ , \new_[17871]_ , \new_[17872]_ , \new_[17876]_ ,
    \new_[17877]_ , \new_[17878]_ , \new_[17881]_ , \new_[17885]_ ,
    \new_[17886]_ , \new_[17887]_ , \new_[17891]_ , \new_[17892]_ ,
    \new_[17896]_ , \new_[17897]_ , \new_[17898]_ , \new_[17901]_ ,
    \new_[17905]_ , \new_[17906]_ , \new_[17907]_ , \new_[17911]_ ,
    \new_[17912]_ , \new_[17916]_ , \new_[17917]_ , \new_[17918]_ ,
    \new_[17921]_ , \new_[17925]_ , \new_[17926]_ , \new_[17927]_ ,
    \new_[17931]_ , \new_[17932]_ , \new_[17936]_ , \new_[17937]_ ,
    \new_[17938]_ , \new_[17941]_ , \new_[17945]_ , \new_[17946]_ ,
    \new_[17947]_ , \new_[17951]_ , \new_[17952]_ , \new_[17956]_ ,
    \new_[17957]_ , \new_[17958]_ , \new_[17961]_ , \new_[17965]_ ,
    \new_[17966]_ , \new_[17967]_ , \new_[17971]_ , \new_[17972]_ ,
    \new_[17976]_ , \new_[17977]_ , \new_[17978]_ , \new_[17981]_ ,
    \new_[17985]_ , \new_[17986]_ , \new_[17987]_ , \new_[17991]_ ,
    \new_[17992]_ , \new_[17996]_ , \new_[17997]_ , \new_[17998]_ ,
    \new_[18001]_ , \new_[18005]_ , \new_[18006]_ , \new_[18007]_ ,
    \new_[18011]_ , \new_[18012]_ , \new_[18016]_ , \new_[18017]_ ,
    \new_[18018]_ , \new_[18021]_ , \new_[18025]_ , \new_[18026]_ ,
    \new_[18027]_ , \new_[18031]_ , \new_[18032]_ , \new_[18036]_ ,
    \new_[18037]_ , \new_[18038]_ , \new_[18041]_ , \new_[18045]_ ,
    \new_[18046]_ , \new_[18047]_ , \new_[18051]_ , \new_[18052]_ ,
    \new_[18056]_ , \new_[18057]_ , \new_[18058]_ , \new_[18061]_ ,
    \new_[18065]_ , \new_[18066]_ , \new_[18067]_ , \new_[18071]_ ,
    \new_[18072]_ , \new_[18076]_ , \new_[18077]_ , \new_[18078]_ ,
    \new_[18081]_ , \new_[18085]_ , \new_[18086]_ , \new_[18087]_ ,
    \new_[18091]_ , \new_[18092]_ , \new_[18096]_ , \new_[18097]_ ,
    \new_[18098]_ , \new_[18101]_ , \new_[18105]_ , \new_[18106]_ ,
    \new_[18107]_ , \new_[18111]_ , \new_[18112]_ , \new_[18116]_ ,
    \new_[18117]_ , \new_[18118]_ , \new_[18121]_ , \new_[18125]_ ,
    \new_[18126]_ , \new_[18127]_ , \new_[18131]_ , \new_[18132]_ ,
    \new_[18136]_ , \new_[18137]_ , \new_[18138]_ , \new_[18141]_ ,
    \new_[18145]_ , \new_[18146]_ , \new_[18147]_ , \new_[18151]_ ,
    \new_[18152]_ , \new_[18156]_ , \new_[18157]_ , \new_[18158]_ ,
    \new_[18161]_ , \new_[18165]_ , \new_[18166]_ , \new_[18167]_ ,
    \new_[18171]_ , \new_[18172]_ , \new_[18176]_ , \new_[18177]_ ,
    \new_[18178]_ , \new_[18181]_ , \new_[18185]_ , \new_[18186]_ ,
    \new_[18187]_ , \new_[18191]_ , \new_[18192]_ , \new_[18196]_ ,
    \new_[18197]_ , \new_[18198]_ , \new_[18201]_ , \new_[18205]_ ,
    \new_[18206]_ , \new_[18207]_ , \new_[18211]_ , \new_[18212]_ ,
    \new_[18216]_ , \new_[18217]_ , \new_[18218]_ , \new_[18221]_ ,
    \new_[18225]_ , \new_[18226]_ , \new_[18227]_ , \new_[18231]_ ,
    \new_[18232]_ , \new_[18236]_ , \new_[18237]_ , \new_[18238]_ ,
    \new_[18241]_ , \new_[18245]_ , \new_[18246]_ , \new_[18247]_ ,
    \new_[18251]_ , \new_[18252]_ , \new_[18256]_ , \new_[18257]_ ,
    \new_[18258]_ , \new_[18261]_ , \new_[18265]_ , \new_[18266]_ ,
    \new_[18267]_ , \new_[18271]_ , \new_[18272]_ , \new_[18276]_ ,
    \new_[18277]_ , \new_[18278]_ , \new_[18281]_ , \new_[18285]_ ,
    \new_[18286]_ , \new_[18287]_ , \new_[18291]_ , \new_[18292]_ ,
    \new_[18296]_ , \new_[18297]_ , \new_[18298]_ , \new_[18301]_ ,
    \new_[18305]_ , \new_[18306]_ , \new_[18307]_ , \new_[18311]_ ,
    \new_[18312]_ , \new_[18316]_ , \new_[18317]_ , \new_[18318]_ ,
    \new_[18321]_ , \new_[18325]_ , \new_[18326]_ , \new_[18327]_ ,
    \new_[18331]_ , \new_[18332]_ , \new_[18336]_ , \new_[18337]_ ,
    \new_[18338]_ , \new_[18341]_ , \new_[18345]_ , \new_[18346]_ ,
    \new_[18347]_ , \new_[18351]_ , \new_[18352]_ , \new_[18356]_ ,
    \new_[18357]_ , \new_[18358]_ , \new_[18361]_ , \new_[18365]_ ,
    \new_[18366]_ , \new_[18367]_ , \new_[18371]_ , \new_[18372]_ ,
    \new_[18376]_ , \new_[18377]_ , \new_[18378]_ , \new_[18381]_ ,
    \new_[18385]_ , \new_[18386]_ , \new_[18387]_ , \new_[18391]_ ,
    \new_[18392]_ , \new_[18396]_ , \new_[18397]_ , \new_[18398]_ ,
    \new_[18401]_ , \new_[18405]_ , \new_[18406]_ , \new_[18407]_ ,
    \new_[18411]_ , \new_[18412]_ , \new_[18416]_ , \new_[18417]_ ,
    \new_[18418]_ , \new_[18421]_ , \new_[18425]_ , \new_[18426]_ ,
    \new_[18427]_ , \new_[18431]_ , \new_[18432]_ , \new_[18436]_ ,
    \new_[18437]_ , \new_[18438]_ , \new_[18441]_ , \new_[18445]_ ,
    \new_[18446]_ , \new_[18447]_ , \new_[18451]_ , \new_[18452]_ ,
    \new_[18456]_ , \new_[18457]_ , \new_[18458]_ , \new_[18461]_ ,
    \new_[18465]_ , \new_[18466]_ , \new_[18467]_ , \new_[18471]_ ,
    \new_[18472]_ , \new_[18476]_ , \new_[18477]_ , \new_[18478]_ ,
    \new_[18481]_ , \new_[18485]_ , \new_[18486]_ , \new_[18487]_ ,
    \new_[18491]_ , \new_[18492]_ , \new_[18496]_ , \new_[18497]_ ,
    \new_[18498]_ , \new_[18501]_ , \new_[18505]_ , \new_[18506]_ ,
    \new_[18507]_ , \new_[18511]_ , \new_[18512]_ , \new_[18516]_ ,
    \new_[18517]_ , \new_[18518]_ , \new_[18521]_ , \new_[18525]_ ,
    \new_[18526]_ , \new_[18527]_ , \new_[18531]_ , \new_[18532]_ ,
    \new_[18536]_ , \new_[18537]_ , \new_[18538]_ , \new_[18541]_ ,
    \new_[18545]_ , \new_[18546]_ , \new_[18547]_ , \new_[18551]_ ,
    \new_[18552]_ , \new_[18556]_ , \new_[18557]_ , \new_[18558]_ ,
    \new_[18561]_ , \new_[18565]_ , \new_[18566]_ , \new_[18567]_ ,
    \new_[18571]_ , \new_[18572]_ , \new_[18576]_ , \new_[18577]_ ,
    \new_[18578]_ , \new_[18581]_ , \new_[18585]_ , \new_[18586]_ ,
    \new_[18587]_ , \new_[18591]_ , \new_[18592]_ , \new_[18596]_ ,
    \new_[18597]_ , \new_[18598]_ , \new_[18601]_ , \new_[18605]_ ,
    \new_[18606]_ , \new_[18607]_ , \new_[18611]_ , \new_[18612]_ ,
    \new_[18616]_ , \new_[18617]_ , \new_[18618]_ , \new_[18621]_ ,
    \new_[18625]_ , \new_[18626]_ , \new_[18627]_ , \new_[18631]_ ,
    \new_[18632]_ , \new_[18636]_ , \new_[18637]_ , \new_[18638]_ ,
    \new_[18641]_ , \new_[18645]_ , \new_[18646]_ , \new_[18647]_ ,
    \new_[18651]_ , \new_[18652]_ , \new_[18656]_ , \new_[18657]_ ,
    \new_[18658]_ , \new_[18661]_ , \new_[18665]_ , \new_[18666]_ ,
    \new_[18667]_ , \new_[18671]_ , \new_[18672]_ , \new_[18676]_ ,
    \new_[18677]_ , \new_[18678]_ , \new_[18681]_ , \new_[18685]_ ,
    \new_[18686]_ , \new_[18687]_ , \new_[18691]_ , \new_[18692]_ ,
    \new_[18696]_ , \new_[18697]_ , \new_[18698]_ , \new_[18701]_ ,
    \new_[18705]_ , \new_[18706]_ , \new_[18707]_ , \new_[18711]_ ,
    \new_[18712]_ , \new_[18716]_ , \new_[18717]_ , \new_[18718]_ ,
    \new_[18721]_ , \new_[18725]_ , \new_[18726]_ , \new_[18727]_ ,
    \new_[18731]_ , \new_[18732]_ , \new_[18736]_ , \new_[18737]_ ,
    \new_[18738]_ , \new_[18741]_ , \new_[18745]_ , \new_[18746]_ ,
    \new_[18747]_ , \new_[18751]_ , \new_[18752]_ , \new_[18756]_ ,
    \new_[18757]_ , \new_[18758]_ , \new_[18761]_ , \new_[18765]_ ,
    \new_[18766]_ , \new_[18767]_ , \new_[18771]_ , \new_[18772]_ ,
    \new_[18776]_ , \new_[18777]_ , \new_[18778]_ , \new_[18781]_ ,
    \new_[18785]_ , \new_[18786]_ , \new_[18787]_ , \new_[18791]_ ,
    \new_[18792]_ , \new_[18796]_ , \new_[18797]_ , \new_[18798]_ ,
    \new_[18801]_ , \new_[18805]_ , \new_[18806]_ , \new_[18807]_ ,
    \new_[18811]_ , \new_[18812]_ , \new_[18816]_ , \new_[18817]_ ,
    \new_[18818]_ , \new_[18821]_ , \new_[18825]_ , \new_[18826]_ ,
    \new_[18827]_ , \new_[18831]_ , \new_[18832]_ , \new_[18836]_ ,
    \new_[18837]_ , \new_[18838]_ , \new_[18841]_ , \new_[18845]_ ,
    \new_[18846]_ , \new_[18847]_ , \new_[18851]_ , \new_[18852]_ ,
    \new_[18856]_ , \new_[18857]_ , \new_[18858]_ , \new_[18861]_ ,
    \new_[18865]_ , \new_[18866]_ , \new_[18867]_ , \new_[18871]_ ,
    \new_[18872]_ , \new_[18876]_ , \new_[18877]_ , \new_[18878]_ ,
    \new_[18881]_ , \new_[18885]_ , \new_[18886]_ , \new_[18887]_ ,
    \new_[18891]_ , \new_[18892]_ , \new_[18896]_ , \new_[18897]_ ,
    \new_[18898]_ , \new_[18901]_ , \new_[18905]_ , \new_[18906]_ ,
    \new_[18907]_ , \new_[18911]_ , \new_[18912]_ , \new_[18916]_ ,
    \new_[18917]_ , \new_[18918]_ , \new_[18921]_ , \new_[18925]_ ,
    \new_[18926]_ , \new_[18927]_ , \new_[18931]_ , \new_[18932]_ ,
    \new_[18936]_ , \new_[18937]_ , \new_[18938]_ , \new_[18941]_ ,
    \new_[18945]_ , \new_[18946]_ , \new_[18947]_ , \new_[18951]_ ,
    \new_[18952]_ , \new_[18956]_ , \new_[18957]_ , \new_[18958]_ ,
    \new_[18961]_ , \new_[18965]_ , \new_[18966]_ , \new_[18967]_ ,
    \new_[18971]_ , \new_[18972]_ , \new_[18976]_ , \new_[18977]_ ,
    \new_[18978]_ , \new_[18981]_ , \new_[18985]_ , \new_[18986]_ ,
    \new_[18987]_ , \new_[18991]_ , \new_[18992]_ , \new_[18996]_ ,
    \new_[18997]_ , \new_[18998]_ , \new_[19001]_ , \new_[19005]_ ,
    \new_[19006]_ , \new_[19007]_ , \new_[19011]_ , \new_[19012]_ ,
    \new_[19016]_ , \new_[19017]_ , \new_[19018]_ , \new_[19021]_ ,
    \new_[19025]_ , \new_[19026]_ , \new_[19027]_ , \new_[19031]_ ,
    \new_[19032]_ , \new_[19036]_ , \new_[19037]_ , \new_[19038]_ ,
    \new_[19041]_ , \new_[19045]_ , \new_[19046]_ , \new_[19047]_ ,
    \new_[19051]_ , \new_[19052]_ , \new_[19056]_ , \new_[19057]_ ,
    \new_[19058]_ , \new_[19061]_ , \new_[19065]_ , \new_[19066]_ ,
    \new_[19067]_ , \new_[19071]_ , \new_[19072]_ , \new_[19076]_ ,
    \new_[19077]_ , \new_[19078]_ , \new_[19081]_ , \new_[19085]_ ,
    \new_[19086]_ , \new_[19087]_ , \new_[19091]_ , \new_[19092]_ ,
    \new_[19096]_ , \new_[19097]_ , \new_[19098]_ , \new_[19101]_ ,
    \new_[19105]_ , \new_[19106]_ , \new_[19107]_ , \new_[19111]_ ,
    \new_[19112]_ , \new_[19116]_ , \new_[19117]_ , \new_[19118]_ ,
    \new_[19121]_ , \new_[19125]_ , \new_[19126]_ , \new_[19127]_ ,
    \new_[19131]_ , \new_[19132]_ , \new_[19136]_ , \new_[19137]_ ,
    \new_[19138]_ , \new_[19141]_ , \new_[19145]_ , \new_[19146]_ ,
    \new_[19147]_ , \new_[19151]_ , \new_[19152]_ , \new_[19156]_ ,
    \new_[19157]_ , \new_[19158]_ , \new_[19161]_ , \new_[19165]_ ,
    \new_[19166]_ , \new_[19167]_ , \new_[19171]_ , \new_[19172]_ ,
    \new_[19176]_ , \new_[19177]_ , \new_[19178]_ , \new_[19181]_ ,
    \new_[19185]_ , \new_[19186]_ , \new_[19187]_ , \new_[19191]_ ,
    \new_[19192]_ , \new_[19196]_ , \new_[19197]_ , \new_[19198]_ ,
    \new_[19201]_ , \new_[19205]_ , \new_[19206]_ , \new_[19207]_ ,
    \new_[19211]_ , \new_[19212]_ , \new_[19216]_ , \new_[19217]_ ,
    \new_[19218]_ , \new_[19221]_ , \new_[19225]_ , \new_[19226]_ ,
    \new_[19227]_ , \new_[19231]_ , \new_[19232]_ , \new_[19236]_ ,
    \new_[19237]_ , \new_[19238]_ , \new_[19241]_ , \new_[19245]_ ,
    \new_[19246]_ , \new_[19247]_ , \new_[19251]_ , \new_[19252]_ ,
    \new_[19256]_ , \new_[19257]_ , \new_[19258]_ , \new_[19261]_ ,
    \new_[19265]_ , \new_[19266]_ , \new_[19267]_ , \new_[19271]_ ,
    \new_[19272]_ , \new_[19276]_ , \new_[19277]_ , \new_[19278]_ ,
    \new_[19281]_ , \new_[19285]_ , \new_[19286]_ , \new_[19287]_ ,
    \new_[19291]_ , \new_[19292]_ , \new_[19296]_ , \new_[19297]_ ,
    \new_[19298]_ , \new_[19301]_ , \new_[19305]_ , \new_[19306]_ ,
    \new_[19307]_ , \new_[19311]_ , \new_[19312]_ , \new_[19316]_ ,
    \new_[19317]_ , \new_[19318]_ , \new_[19321]_ , \new_[19325]_ ,
    \new_[19326]_ , \new_[19327]_ , \new_[19331]_ , \new_[19332]_ ,
    \new_[19336]_ , \new_[19337]_ , \new_[19338]_ , \new_[19341]_ ,
    \new_[19345]_ , \new_[19346]_ , \new_[19347]_ , \new_[19351]_ ,
    \new_[19352]_ , \new_[19356]_ , \new_[19357]_ , \new_[19358]_ ,
    \new_[19361]_ , \new_[19365]_ , \new_[19366]_ , \new_[19367]_ ,
    \new_[19371]_ , \new_[19372]_ , \new_[19376]_ , \new_[19377]_ ,
    \new_[19378]_ , \new_[19381]_ , \new_[19385]_ , \new_[19386]_ ,
    \new_[19387]_ , \new_[19391]_ , \new_[19392]_ , \new_[19396]_ ,
    \new_[19397]_ , \new_[19398]_ , \new_[19401]_ , \new_[19405]_ ,
    \new_[19406]_ , \new_[19407]_ , \new_[19411]_ , \new_[19412]_ ,
    \new_[19416]_ , \new_[19417]_ , \new_[19418]_ , \new_[19421]_ ,
    \new_[19425]_ , \new_[19426]_ , \new_[19427]_ , \new_[19431]_ ,
    \new_[19432]_ , \new_[19436]_ , \new_[19437]_ , \new_[19438]_ ,
    \new_[19441]_ , \new_[19445]_ , \new_[19446]_ , \new_[19447]_ ,
    \new_[19451]_ , \new_[19452]_ , \new_[19456]_ , \new_[19457]_ ,
    \new_[19458]_ , \new_[19461]_ , \new_[19465]_ , \new_[19466]_ ,
    \new_[19467]_ , \new_[19471]_ , \new_[19472]_ , \new_[19476]_ ,
    \new_[19477]_ , \new_[19478]_ , \new_[19481]_ , \new_[19485]_ ,
    \new_[19486]_ , \new_[19487]_ , \new_[19491]_ , \new_[19492]_ ,
    \new_[19496]_ , \new_[19497]_ , \new_[19498]_ , \new_[19501]_ ,
    \new_[19505]_ , \new_[19506]_ , \new_[19507]_ , \new_[19511]_ ,
    \new_[19512]_ , \new_[19516]_ , \new_[19517]_ , \new_[19518]_ ,
    \new_[19521]_ , \new_[19525]_ , \new_[19526]_ , \new_[19527]_ ,
    \new_[19531]_ , \new_[19532]_ , \new_[19536]_ , \new_[19537]_ ,
    \new_[19538]_ , \new_[19541]_ , \new_[19545]_ , \new_[19546]_ ,
    \new_[19547]_ , \new_[19551]_ , \new_[19552]_ , \new_[19556]_ ,
    \new_[19557]_ , \new_[19558]_ , \new_[19561]_ , \new_[19565]_ ,
    \new_[19566]_ , \new_[19567]_ , \new_[19571]_ , \new_[19572]_ ,
    \new_[19576]_ , \new_[19577]_ , \new_[19578]_ , \new_[19581]_ ,
    \new_[19585]_ , \new_[19586]_ , \new_[19587]_ , \new_[19591]_ ,
    \new_[19592]_ , \new_[19596]_ , \new_[19597]_ , \new_[19598]_ ,
    \new_[19601]_ , \new_[19605]_ , \new_[19606]_ , \new_[19607]_ ,
    \new_[19611]_ , \new_[19612]_ , \new_[19616]_ , \new_[19617]_ ,
    \new_[19618]_ , \new_[19621]_ , \new_[19625]_ , \new_[19626]_ ,
    \new_[19627]_ , \new_[19631]_ , \new_[19632]_ , \new_[19636]_ ,
    \new_[19637]_ , \new_[19638]_ , \new_[19641]_ , \new_[19645]_ ,
    \new_[19646]_ , \new_[19647]_ , \new_[19651]_ , \new_[19652]_ ,
    \new_[19656]_ , \new_[19657]_ , \new_[19658]_ , \new_[19661]_ ,
    \new_[19665]_ , \new_[19666]_ , \new_[19667]_ , \new_[19671]_ ,
    \new_[19672]_ , \new_[19676]_ , \new_[19677]_ , \new_[19678]_ ,
    \new_[19681]_ , \new_[19685]_ , \new_[19686]_ , \new_[19687]_ ,
    \new_[19691]_ , \new_[19692]_ , \new_[19696]_ , \new_[19697]_ ,
    \new_[19698]_ , \new_[19701]_ , \new_[19705]_ , \new_[19706]_ ,
    \new_[19707]_ , \new_[19711]_ , \new_[19712]_ , \new_[19716]_ ,
    \new_[19717]_ , \new_[19718]_ , \new_[19721]_ , \new_[19725]_ ,
    \new_[19726]_ , \new_[19727]_ , \new_[19731]_ , \new_[19732]_ ,
    \new_[19736]_ , \new_[19737]_ , \new_[19738]_ , \new_[19741]_ ,
    \new_[19745]_ , \new_[19746]_ , \new_[19747]_ , \new_[19751]_ ,
    \new_[19752]_ , \new_[19756]_ , \new_[19757]_ , \new_[19758]_ ,
    \new_[19761]_ , \new_[19765]_ , \new_[19766]_ , \new_[19767]_ ,
    \new_[19771]_ , \new_[19772]_ , \new_[19776]_ , \new_[19777]_ ,
    \new_[19778]_ , \new_[19781]_ , \new_[19785]_ , \new_[19786]_ ,
    \new_[19787]_ , \new_[19791]_ , \new_[19792]_ , \new_[19796]_ ,
    \new_[19797]_ , \new_[19798]_ , \new_[19801]_ , \new_[19805]_ ,
    \new_[19806]_ , \new_[19807]_ , \new_[19811]_ , \new_[19812]_ ,
    \new_[19816]_ , \new_[19817]_ , \new_[19818]_ , \new_[19821]_ ,
    \new_[19825]_ , \new_[19826]_ , \new_[19827]_ , \new_[19831]_ ,
    \new_[19832]_ , \new_[19836]_ , \new_[19837]_ , \new_[19838]_ ,
    \new_[19841]_ , \new_[19845]_ , \new_[19846]_ , \new_[19847]_ ,
    \new_[19851]_ , \new_[19852]_ , \new_[19856]_ , \new_[19857]_ ,
    \new_[19858]_ , \new_[19861]_ , \new_[19865]_ , \new_[19866]_ ,
    \new_[19867]_ , \new_[19871]_ , \new_[19872]_ , \new_[19876]_ ,
    \new_[19877]_ , \new_[19878]_ , \new_[19881]_ , \new_[19885]_ ,
    \new_[19886]_ , \new_[19887]_ , \new_[19891]_ , \new_[19892]_ ,
    \new_[19896]_ , \new_[19897]_ , \new_[19898]_ , \new_[19901]_ ,
    \new_[19905]_ , \new_[19906]_ , \new_[19907]_ , \new_[19911]_ ,
    \new_[19912]_ , \new_[19916]_ , \new_[19917]_ , \new_[19918]_ ,
    \new_[19921]_ , \new_[19925]_ , \new_[19926]_ , \new_[19927]_ ,
    \new_[19931]_ , \new_[19932]_ , \new_[19936]_ , \new_[19937]_ ,
    \new_[19938]_ , \new_[19941]_ , \new_[19945]_ , \new_[19946]_ ,
    \new_[19947]_ , \new_[19951]_ , \new_[19952]_ , \new_[19956]_ ,
    \new_[19957]_ , \new_[19958]_ , \new_[19961]_ , \new_[19965]_ ,
    \new_[19966]_ , \new_[19967]_ , \new_[19971]_ , \new_[19972]_ ,
    \new_[19976]_ , \new_[19977]_ , \new_[19978]_ , \new_[19981]_ ,
    \new_[19985]_ , \new_[19986]_ , \new_[19987]_ , \new_[19991]_ ,
    \new_[19992]_ , \new_[19996]_ , \new_[19997]_ , \new_[19998]_ ,
    \new_[20001]_ , \new_[20005]_ , \new_[20006]_ , \new_[20007]_ ,
    \new_[20011]_ , \new_[20012]_ , \new_[20016]_ , \new_[20017]_ ,
    \new_[20018]_ , \new_[20021]_ , \new_[20025]_ , \new_[20026]_ ,
    \new_[20027]_ , \new_[20031]_ , \new_[20032]_ , \new_[20036]_ ,
    \new_[20037]_ , \new_[20038]_ , \new_[20041]_ , \new_[20045]_ ,
    \new_[20046]_ , \new_[20047]_ , \new_[20051]_ , \new_[20052]_ ,
    \new_[20056]_ , \new_[20057]_ , \new_[20058]_ , \new_[20061]_ ,
    \new_[20065]_ , \new_[20066]_ , \new_[20067]_ , \new_[20071]_ ,
    \new_[20072]_ , \new_[20076]_ , \new_[20077]_ , \new_[20078]_ ,
    \new_[20081]_ , \new_[20085]_ , \new_[20086]_ , \new_[20087]_ ,
    \new_[20091]_ , \new_[20092]_ , \new_[20096]_ , \new_[20097]_ ,
    \new_[20098]_ , \new_[20101]_ , \new_[20105]_ , \new_[20106]_ ,
    \new_[20107]_ , \new_[20111]_ , \new_[20112]_ , \new_[20116]_ ,
    \new_[20117]_ , \new_[20118]_ , \new_[20121]_ , \new_[20125]_ ,
    \new_[20126]_ , \new_[20127]_ , \new_[20131]_ , \new_[20132]_ ,
    \new_[20136]_ , \new_[20137]_ , \new_[20138]_ , \new_[20141]_ ,
    \new_[20145]_ , \new_[20146]_ , \new_[20147]_ , \new_[20151]_ ,
    \new_[20152]_ , \new_[20156]_ , \new_[20157]_ , \new_[20158]_ ,
    \new_[20161]_ , \new_[20165]_ , \new_[20166]_ , \new_[20167]_ ,
    \new_[20171]_ , \new_[20172]_ , \new_[20176]_ , \new_[20177]_ ,
    \new_[20178]_ , \new_[20181]_ , \new_[20185]_ , \new_[20186]_ ,
    \new_[20187]_ , \new_[20191]_ , \new_[20192]_ , \new_[20196]_ ,
    \new_[20197]_ , \new_[20198]_ , \new_[20201]_ , \new_[20205]_ ,
    \new_[20206]_ , \new_[20207]_ , \new_[20211]_ , \new_[20212]_ ,
    \new_[20216]_ , \new_[20217]_ , \new_[20218]_ , \new_[20221]_ ,
    \new_[20225]_ , \new_[20226]_ , \new_[20227]_ , \new_[20231]_ ,
    \new_[20232]_ , \new_[20236]_ , \new_[20237]_ , \new_[20238]_ ,
    \new_[20241]_ , \new_[20245]_ , \new_[20246]_ , \new_[20247]_ ,
    \new_[20251]_ , \new_[20252]_ , \new_[20256]_ , \new_[20257]_ ,
    \new_[20258]_ , \new_[20261]_ , \new_[20265]_ , \new_[20266]_ ,
    \new_[20267]_ , \new_[20271]_ , \new_[20272]_ , \new_[20276]_ ,
    \new_[20277]_ , \new_[20278]_ , \new_[20281]_ , \new_[20285]_ ,
    \new_[20286]_ , \new_[20287]_ , \new_[20291]_ , \new_[20292]_ ,
    \new_[20296]_ , \new_[20297]_ , \new_[20298]_ , \new_[20301]_ ,
    \new_[20305]_ , \new_[20306]_ , \new_[20307]_ , \new_[20311]_ ,
    \new_[20312]_ , \new_[20316]_ , \new_[20317]_ , \new_[20318]_ ,
    \new_[20321]_ , \new_[20325]_ , \new_[20326]_ , \new_[20327]_ ,
    \new_[20331]_ , \new_[20332]_ , \new_[20336]_ , \new_[20337]_ ,
    \new_[20338]_ , \new_[20341]_ , \new_[20345]_ , \new_[20346]_ ,
    \new_[20347]_ , \new_[20351]_ , \new_[20352]_ , \new_[20356]_ ,
    \new_[20357]_ , \new_[20358]_ , \new_[20361]_ , \new_[20365]_ ,
    \new_[20366]_ , \new_[20367]_ , \new_[20371]_ , \new_[20372]_ ,
    \new_[20376]_ , \new_[20377]_ , \new_[20378]_ , \new_[20381]_ ,
    \new_[20385]_ , \new_[20386]_ , \new_[20387]_ , \new_[20391]_ ,
    \new_[20392]_ , \new_[20396]_ , \new_[20397]_ , \new_[20398]_ ,
    \new_[20401]_ , \new_[20405]_ , \new_[20406]_ , \new_[20407]_ ,
    \new_[20411]_ , \new_[20412]_ , \new_[20416]_ , \new_[20417]_ ,
    \new_[20418]_ , \new_[20421]_ , \new_[20425]_ , \new_[20426]_ ,
    \new_[20427]_ , \new_[20431]_ , \new_[20432]_ , \new_[20436]_ ,
    \new_[20437]_ , \new_[20438]_ , \new_[20441]_ , \new_[20445]_ ,
    \new_[20446]_ , \new_[20447]_ , \new_[20451]_ , \new_[20452]_ ,
    \new_[20456]_ , \new_[20457]_ , \new_[20458]_ , \new_[20461]_ ,
    \new_[20465]_ , \new_[20466]_ , \new_[20467]_ , \new_[20471]_ ,
    \new_[20472]_ , \new_[20476]_ , \new_[20477]_ , \new_[20478]_ ,
    \new_[20481]_ , \new_[20485]_ , \new_[20486]_ , \new_[20487]_ ,
    \new_[20491]_ , \new_[20492]_ , \new_[20496]_ , \new_[20497]_ ,
    \new_[20498]_ , \new_[20501]_ , \new_[20505]_ , \new_[20506]_ ,
    \new_[20507]_ , \new_[20511]_ , \new_[20512]_ , \new_[20516]_ ,
    \new_[20517]_ , \new_[20518]_ , \new_[20521]_ , \new_[20525]_ ,
    \new_[20526]_ , \new_[20527]_ , \new_[20531]_ , \new_[20532]_ ,
    \new_[20536]_ , \new_[20537]_ , \new_[20538]_ , \new_[20541]_ ,
    \new_[20545]_ , \new_[20546]_ , \new_[20547]_ , \new_[20551]_ ,
    \new_[20552]_ , \new_[20556]_ , \new_[20557]_ , \new_[20558]_ ,
    \new_[20561]_ , \new_[20565]_ , \new_[20566]_ , \new_[20567]_ ,
    \new_[20571]_ , \new_[20572]_ , \new_[20576]_ , \new_[20577]_ ,
    \new_[20578]_ , \new_[20581]_ , \new_[20585]_ , \new_[20586]_ ,
    \new_[20587]_ , \new_[20591]_ , \new_[20592]_ , \new_[20596]_ ,
    \new_[20597]_ , \new_[20598]_ , \new_[20601]_ , \new_[20605]_ ,
    \new_[20606]_ , \new_[20607]_ , \new_[20611]_ , \new_[20612]_ ,
    \new_[20616]_ , \new_[20617]_ , \new_[20618]_ , \new_[20621]_ ,
    \new_[20625]_ , \new_[20626]_ , \new_[20627]_ , \new_[20631]_ ,
    \new_[20632]_ , \new_[20636]_ , \new_[20637]_ , \new_[20638]_ ,
    \new_[20641]_ , \new_[20645]_ , \new_[20646]_ , \new_[20647]_ ,
    \new_[20651]_ , \new_[20652]_ , \new_[20656]_ , \new_[20657]_ ,
    \new_[20658]_ , \new_[20661]_ , \new_[20665]_ , \new_[20666]_ ,
    \new_[20667]_ , \new_[20671]_ , \new_[20672]_ , \new_[20676]_ ,
    \new_[20677]_ , \new_[20678]_ , \new_[20681]_ , \new_[20685]_ ,
    \new_[20686]_ , \new_[20687]_ , \new_[20691]_ , \new_[20692]_ ,
    \new_[20696]_ , \new_[20697]_ , \new_[20698]_ , \new_[20701]_ ,
    \new_[20705]_ , \new_[20706]_ , \new_[20707]_ , \new_[20711]_ ,
    \new_[20712]_ , \new_[20716]_ , \new_[20717]_ , \new_[20718]_ ,
    \new_[20721]_ , \new_[20725]_ , \new_[20726]_ , \new_[20727]_ ,
    \new_[20731]_ , \new_[20732]_ , \new_[20736]_ , \new_[20737]_ ,
    \new_[20738]_ , \new_[20741]_ , \new_[20745]_ , \new_[20746]_ ,
    \new_[20747]_ , \new_[20751]_ , \new_[20752]_ , \new_[20756]_ ,
    \new_[20757]_ , \new_[20758]_ , \new_[20761]_ , \new_[20765]_ ,
    \new_[20766]_ , \new_[20767]_ , \new_[20771]_ , \new_[20772]_ ,
    \new_[20776]_ , \new_[20777]_ , \new_[20778]_ , \new_[20781]_ ,
    \new_[20785]_ , \new_[20786]_ , \new_[20787]_ , \new_[20791]_ ,
    \new_[20792]_ , \new_[20796]_ , \new_[20797]_ , \new_[20798]_ ,
    \new_[20801]_ , \new_[20805]_ , \new_[20806]_ , \new_[20807]_ ,
    \new_[20811]_ , \new_[20812]_ , \new_[20816]_ , \new_[20817]_ ,
    \new_[20818]_ , \new_[20821]_ , \new_[20825]_ , \new_[20826]_ ,
    \new_[20827]_ , \new_[20831]_ , \new_[20832]_ , \new_[20836]_ ,
    \new_[20837]_ , \new_[20838]_ , \new_[20841]_ , \new_[20845]_ ,
    \new_[20846]_ , \new_[20847]_ , \new_[20851]_ , \new_[20852]_ ,
    \new_[20856]_ , \new_[20857]_ , \new_[20858]_ , \new_[20861]_ ,
    \new_[20865]_ , \new_[20866]_ , \new_[20867]_ , \new_[20871]_ ,
    \new_[20872]_ , \new_[20876]_ , \new_[20877]_ , \new_[20878]_ ,
    \new_[20881]_ , \new_[20885]_ , \new_[20886]_ , \new_[20887]_ ,
    \new_[20891]_ , \new_[20892]_ , \new_[20896]_ , \new_[20897]_ ,
    \new_[20898]_ , \new_[20901]_ , \new_[20905]_ , \new_[20906]_ ,
    \new_[20907]_ , \new_[20911]_ , \new_[20912]_ , \new_[20916]_ ,
    \new_[20917]_ , \new_[20918]_ , \new_[20921]_ , \new_[20925]_ ,
    \new_[20926]_ , \new_[20927]_ , \new_[20931]_ , \new_[20932]_ ,
    \new_[20936]_ , \new_[20937]_ , \new_[20938]_ , \new_[20941]_ ,
    \new_[20945]_ , \new_[20946]_ , \new_[20947]_ , \new_[20951]_ ,
    \new_[20952]_ , \new_[20956]_ , \new_[20957]_ , \new_[20958]_ ,
    \new_[20961]_ , \new_[20965]_ , \new_[20966]_ , \new_[20967]_ ,
    \new_[20971]_ , \new_[20972]_ , \new_[20976]_ , \new_[20977]_ ,
    \new_[20978]_ , \new_[20981]_ , \new_[20985]_ , \new_[20986]_ ,
    \new_[20987]_ , \new_[20991]_ , \new_[20992]_ , \new_[20996]_ ,
    \new_[20997]_ , \new_[20998]_ , \new_[21001]_ , \new_[21005]_ ,
    \new_[21006]_ , \new_[21007]_ , \new_[21011]_ , \new_[21012]_ ,
    \new_[21016]_ , \new_[21017]_ , \new_[21018]_ , \new_[21021]_ ,
    \new_[21025]_ , \new_[21026]_ , \new_[21027]_ , \new_[21031]_ ,
    \new_[21032]_ , \new_[21036]_ , \new_[21037]_ , \new_[21038]_ ,
    \new_[21041]_ , \new_[21045]_ , \new_[21046]_ , \new_[21047]_ ,
    \new_[21051]_ , \new_[21052]_ , \new_[21056]_ , \new_[21057]_ ,
    \new_[21058]_ , \new_[21061]_ , \new_[21065]_ , \new_[21066]_ ,
    \new_[21067]_ , \new_[21071]_ , \new_[21072]_ , \new_[21076]_ ,
    \new_[21077]_ , \new_[21078]_ , \new_[21081]_ , \new_[21085]_ ,
    \new_[21086]_ , \new_[21087]_ , \new_[21091]_ , \new_[21092]_ ,
    \new_[21096]_ , \new_[21097]_ , \new_[21098]_ , \new_[21101]_ ,
    \new_[21105]_ , \new_[21106]_ , \new_[21107]_ , \new_[21111]_ ,
    \new_[21112]_ , \new_[21116]_ , \new_[21117]_ , \new_[21118]_ ,
    \new_[21121]_ , \new_[21125]_ , \new_[21126]_ , \new_[21127]_ ,
    \new_[21131]_ , \new_[21132]_ , \new_[21136]_ , \new_[21137]_ ,
    \new_[21138]_ , \new_[21141]_ , \new_[21145]_ , \new_[21146]_ ,
    \new_[21147]_ , \new_[21151]_ , \new_[21152]_ , \new_[21156]_ ,
    \new_[21157]_ , \new_[21158]_ , \new_[21161]_ , \new_[21165]_ ,
    \new_[21166]_ , \new_[21167]_ , \new_[21171]_ , \new_[21172]_ ,
    \new_[21176]_ , \new_[21177]_ , \new_[21178]_ , \new_[21181]_ ,
    \new_[21185]_ , \new_[21186]_ , \new_[21187]_ , \new_[21191]_ ,
    \new_[21192]_ , \new_[21196]_ , \new_[21197]_ , \new_[21198]_ ,
    \new_[21201]_ , \new_[21205]_ , \new_[21206]_ , \new_[21207]_ ,
    \new_[21211]_ , \new_[21212]_ , \new_[21216]_ , \new_[21217]_ ,
    \new_[21218]_ , \new_[21221]_ , \new_[21225]_ , \new_[21226]_ ,
    \new_[21227]_ , \new_[21231]_ , \new_[21232]_ , \new_[21236]_ ,
    \new_[21237]_ , \new_[21238]_ , \new_[21241]_ , \new_[21245]_ ,
    \new_[21246]_ , \new_[21247]_ , \new_[21251]_ , \new_[21252]_ ,
    \new_[21256]_ , \new_[21257]_ , \new_[21258]_ , \new_[21261]_ ,
    \new_[21265]_ , \new_[21266]_ , \new_[21267]_ , \new_[21271]_ ,
    \new_[21272]_ , \new_[21276]_ , \new_[21277]_ , \new_[21278]_ ,
    \new_[21281]_ , \new_[21285]_ , \new_[21286]_ , \new_[21287]_ ,
    \new_[21291]_ , \new_[21292]_ , \new_[21296]_ , \new_[21297]_ ,
    \new_[21298]_ , \new_[21301]_ , \new_[21305]_ , \new_[21306]_ ,
    \new_[21307]_ , \new_[21311]_ , \new_[21312]_ , \new_[21316]_ ,
    \new_[21317]_ , \new_[21318]_ , \new_[21321]_ , \new_[21325]_ ,
    \new_[21326]_ , \new_[21327]_ , \new_[21331]_ , \new_[21332]_ ,
    \new_[21336]_ , \new_[21337]_ , \new_[21338]_ , \new_[21341]_ ,
    \new_[21345]_ , \new_[21346]_ , \new_[21347]_ , \new_[21351]_ ,
    \new_[21352]_ , \new_[21356]_ , \new_[21357]_ , \new_[21358]_ ,
    \new_[21361]_ , \new_[21365]_ , \new_[21366]_ , \new_[21367]_ ,
    \new_[21371]_ , \new_[21372]_ , \new_[21376]_ , \new_[21377]_ ,
    \new_[21378]_ , \new_[21381]_ , \new_[21385]_ , \new_[21386]_ ,
    \new_[21387]_ , \new_[21391]_ , \new_[21392]_ , \new_[21396]_ ,
    \new_[21397]_ , \new_[21398]_ , \new_[21401]_ , \new_[21405]_ ,
    \new_[21406]_ , \new_[21407]_ , \new_[21411]_ , \new_[21412]_ ,
    \new_[21416]_ , \new_[21417]_ , \new_[21418]_ , \new_[21421]_ ,
    \new_[21425]_ , \new_[21426]_ , \new_[21427]_ , \new_[21431]_ ,
    \new_[21432]_ , \new_[21436]_ , \new_[21437]_ , \new_[21438]_ ,
    \new_[21441]_ , \new_[21445]_ , \new_[21446]_ , \new_[21447]_ ,
    \new_[21451]_ , \new_[21452]_ , \new_[21456]_ , \new_[21457]_ ,
    \new_[21458]_ , \new_[21461]_ , \new_[21465]_ , \new_[21466]_ ,
    \new_[21467]_ , \new_[21471]_ , \new_[21472]_ , \new_[21476]_ ,
    \new_[21477]_ , \new_[21478]_ , \new_[21481]_ , \new_[21485]_ ,
    \new_[21486]_ , \new_[21487]_ , \new_[21491]_ , \new_[21492]_ ,
    \new_[21496]_ , \new_[21497]_ , \new_[21498]_ , \new_[21501]_ ,
    \new_[21505]_ , \new_[21506]_ , \new_[21507]_ , \new_[21511]_ ,
    \new_[21512]_ , \new_[21516]_ , \new_[21517]_ , \new_[21518]_ ,
    \new_[21521]_ , \new_[21525]_ , \new_[21526]_ , \new_[21527]_ ,
    \new_[21531]_ , \new_[21532]_ , \new_[21536]_ , \new_[21537]_ ,
    \new_[21538]_ , \new_[21541]_ , \new_[21545]_ , \new_[21546]_ ,
    \new_[21547]_ , \new_[21551]_ , \new_[21552]_ , \new_[21556]_ ,
    \new_[21557]_ , \new_[21558]_ , \new_[21561]_ , \new_[21565]_ ,
    \new_[21566]_ , \new_[21567]_ , \new_[21571]_ , \new_[21572]_ ,
    \new_[21576]_ , \new_[21577]_ , \new_[21578]_ , \new_[21581]_ ,
    \new_[21585]_ , \new_[21586]_ , \new_[21587]_ , \new_[21591]_ ,
    \new_[21592]_ , \new_[21596]_ , \new_[21597]_ , \new_[21598]_ ,
    \new_[21601]_ , \new_[21605]_ , \new_[21606]_ , \new_[21607]_ ,
    \new_[21611]_ , \new_[21612]_ , \new_[21616]_ , \new_[21617]_ ,
    \new_[21618]_ , \new_[21621]_ , \new_[21625]_ , \new_[21626]_ ,
    \new_[21627]_ , \new_[21631]_ , \new_[21632]_ , \new_[21636]_ ,
    \new_[21637]_ , \new_[21638]_ , \new_[21641]_ , \new_[21645]_ ,
    \new_[21646]_ , \new_[21647]_ , \new_[21651]_ , \new_[21652]_ ,
    \new_[21656]_ , \new_[21657]_ , \new_[21658]_ , \new_[21661]_ ,
    \new_[21665]_ , \new_[21666]_ , \new_[21667]_ , \new_[21671]_ ,
    \new_[21672]_ , \new_[21676]_ , \new_[21677]_ , \new_[21678]_ ,
    \new_[21681]_ , \new_[21685]_ , \new_[21686]_ , \new_[21687]_ ,
    \new_[21691]_ , \new_[21692]_ , \new_[21696]_ , \new_[21697]_ ,
    \new_[21698]_ , \new_[21701]_ , \new_[21705]_ , \new_[21706]_ ,
    \new_[21707]_ , \new_[21711]_ , \new_[21712]_ , \new_[21716]_ ,
    \new_[21717]_ , \new_[21718]_ , \new_[21721]_ , \new_[21725]_ ,
    \new_[21726]_ , \new_[21727]_ , \new_[21731]_ , \new_[21732]_ ,
    \new_[21736]_ , \new_[21737]_ , \new_[21738]_ , \new_[21741]_ ,
    \new_[21745]_ , \new_[21746]_ , \new_[21747]_ , \new_[21751]_ ,
    \new_[21752]_ , \new_[21756]_ , \new_[21757]_ , \new_[21758]_ ,
    \new_[21761]_ , \new_[21765]_ , \new_[21766]_ , \new_[21767]_ ,
    \new_[21771]_ , \new_[21772]_ , \new_[21776]_ , \new_[21777]_ ,
    \new_[21778]_ , \new_[21781]_ , \new_[21785]_ , \new_[21786]_ ,
    \new_[21787]_ , \new_[21791]_ , \new_[21792]_ , \new_[21796]_ ,
    \new_[21797]_ , \new_[21798]_ , \new_[21801]_ , \new_[21805]_ ,
    \new_[21806]_ , \new_[21807]_ , \new_[21811]_ , \new_[21812]_ ,
    \new_[21816]_ , \new_[21817]_ , \new_[21818]_ , \new_[21821]_ ,
    \new_[21825]_ , \new_[21826]_ , \new_[21827]_ , \new_[21831]_ ,
    \new_[21832]_ , \new_[21836]_ , \new_[21837]_ , \new_[21838]_ ,
    \new_[21841]_ , \new_[21845]_ , \new_[21846]_ , \new_[21847]_ ,
    \new_[21851]_ , \new_[21852]_ , \new_[21856]_ , \new_[21857]_ ,
    \new_[21858]_ , \new_[21861]_ , \new_[21865]_ , \new_[21866]_ ,
    \new_[21867]_ , \new_[21871]_ , \new_[21872]_ , \new_[21876]_ ,
    \new_[21877]_ , \new_[21878]_ , \new_[21881]_ , \new_[21885]_ ,
    \new_[21886]_ , \new_[21887]_ , \new_[21891]_ , \new_[21892]_ ,
    \new_[21896]_ , \new_[21897]_ , \new_[21898]_ , \new_[21901]_ ,
    \new_[21905]_ , \new_[21906]_ , \new_[21907]_ , \new_[21911]_ ,
    \new_[21912]_ , \new_[21916]_ , \new_[21917]_ , \new_[21918]_ ,
    \new_[21921]_ , \new_[21925]_ , \new_[21926]_ , \new_[21927]_ ,
    \new_[21931]_ , \new_[21932]_ , \new_[21936]_ , \new_[21937]_ ,
    \new_[21938]_ , \new_[21941]_ , \new_[21945]_ , \new_[21946]_ ,
    \new_[21947]_ , \new_[21951]_ , \new_[21952]_ , \new_[21956]_ ,
    \new_[21957]_ , \new_[21958]_ , \new_[21961]_ , \new_[21965]_ ,
    \new_[21966]_ , \new_[21967]_ , \new_[21971]_ , \new_[21972]_ ,
    \new_[21976]_ , \new_[21977]_ , \new_[21978]_ , \new_[21981]_ ,
    \new_[21985]_ , \new_[21986]_ , \new_[21987]_ , \new_[21991]_ ,
    \new_[21992]_ , \new_[21996]_ , \new_[21997]_ , \new_[21998]_ ,
    \new_[22001]_ , \new_[22005]_ , \new_[22006]_ , \new_[22007]_ ,
    \new_[22011]_ , \new_[22012]_ , \new_[22016]_ , \new_[22017]_ ,
    \new_[22018]_ , \new_[22021]_ , \new_[22025]_ , \new_[22026]_ ,
    \new_[22027]_ , \new_[22031]_ , \new_[22032]_ , \new_[22036]_ ,
    \new_[22037]_ , \new_[22038]_ , \new_[22041]_ , \new_[22045]_ ,
    \new_[22046]_ , \new_[22047]_ , \new_[22051]_ , \new_[22052]_ ,
    \new_[22056]_ , \new_[22057]_ , \new_[22058]_ , \new_[22061]_ ,
    \new_[22065]_ , \new_[22066]_ , \new_[22067]_ , \new_[22071]_ ,
    \new_[22072]_ , \new_[22076]_ , \new_[22077]_ , \new_[22078]_ ,
    \new_[22081]_ , \new_[22085]_ , \new_[22086]_ , \new_[22087]_ ,
    \new_[22091]_ , \new_[22092]_ , \new_[22096]_ , \new_[22097]_ ,
    \new_[22098]_ , \new_[22101]_ , \new_[22105]_ , \new_[22106]_ ,
    \new_[22107]_ , \new_[22111]_ , \new_[22112]_ , \new_[22116]_ ,
    \new_[22117]_ , \new_[22118]_ , \new_[22121]_ , \new_[22125]_ ,
    \new_[22126]_ , \new_[22127]_ , \new_[22131]_ , \new_[22132]_ ,
    \new_[22136]_ , \new_[22137]_ , \new_[22138]_ , \new_[22141]_ ,
    \new_[22145]_ , \new_[22146]_ , \new_[22147]_ , \new_[22151]_ ,
    \new_[22152]_ , \new_[22156]_ , \new_[22157]_ , \new_[22158]_ ,
    \new_[22161]_ , \new_[22165]_ , \new_[22166]_ , \new_[22167]_ ,
    \new_[22171]_ , \new_[22172]_ , \new_[22176]_ , \new_[22177]_ ,
    \new_[22178]_ , \new_[22181]_ , \new_[22185]_ , \new_[22186]_ ,
    \new_[22187]_ , \new_[22191]_ , \new_[22192]_ , \new_[22196]_ ,
    \new_[22197]_ , \new_[22198]_ , \new_[22201]_ , \new_[22205]_ ,
    \new_[22206]_ , \new_[22207]_ , \new_[22211]_ , \new_[22212]_ ,
    \new_[22216]_ , \new_[22217]_ , \new_[22218]_ , \new_[22221]_ ,
    \new_[22225]_ , \new_[22226]_ , \new_[22227]_ , \new_[22231]_ ,
    \new_[22232]_ , \new_[22236]_ , \new_[22237]_ , \new_[22238]_ ,
    \new_[22241]_ , \new_[22245]_ , \new_[22246]_ , \new_[22247]_ ,
    \new_[22251]_ , \new_[22252]_ , \new_[22256]_ , \new_[22257]_ ,
    \new_[22258]_ , \new_[22261]_ , \new_[22265]_ , \new_[22266]_ ,
    \new_[22267]_ , \new_[22271]_ , \new_[22272]_ , \new_[22276]_ ,
    \new_[22277]_ , \new_[22278]_ , \new_[22281]_ , \new_[22285]_ ,
    \new_[22286]_ , \new_[22287]_ , \new_[22291]_ , \new_[22292]_ ,
    \new_[22296]_ , \new_[22297]_ , \new_[22298]_ , \new_[22301]_ ,
    \new_[22305]_ , \new_[22306]_ , \new_[22307]_ , \new_[22311]_ ,
    \new_[22312]_ , \new_[22316]_ , \new_[22317]_ , \new_[22318]_ ,
    \new_[22321]_ , \new_[22325]_ , \new_[22326]_ , \new_[22327]_ ,
    \new_[22331]_ , \new_[22332]_ , \new_[22336]_ , \new_[22337]_ ,
    \new_[22338]_ , \new_[22341]_ , \new_[22345]_ , \new_[22346]_ ,
    \new_[22347]_ , \new_[22351]_ , \new_[22352]_ , \new_[22356]_ ,
    \new_[22357]_ , \new_[22358]_ , \new_[22361]_ , \new_[22365]_ ,
    \new_[22366]_ , \new_[22367]_ , \new_[22371]_ , \new_[22372]_ ,
    \new_[22376]_ , \new_[22377]_ , \new_[22378]_ , \new_[22381]_ ,
    \new_[22385]_ , \new_[22386]_ , \new_[22387]_ , \new_[22391]_ ,
    \new_[22392]_ , \new_[22396]_ , \new_[22397]_ , \new_[22398]_ ,
    \new_[22401]_ , \new_[22405]_ , \new_[22406]_ , \new_[22407]_ ,
    \new_[22411]_ , \new_[22412]_ , \new_[22416]_ , \new_[22417]_ ,
    \new_[22418]_ , \new_[22421]_ , \new_[22425]_ , \new_[22426]_ ,
    \new_[22427]_ , \new_[22431]_ , \new_[22432]_ , \new_[22436]_ ,
    \new_[22437]_ , \new_[22438]_ , \new_[22441]_ , \new_[22445]_ ,
    \new_[22446]_ , \new_[22447]_ , \new_[22451]_ , \new_[22452]_ ,
    \new_[22456]_ , \new_[22457]_ , \new_[22458]_ , \new_[22461]_ ,
    \new_[22465]_ , \new_[22466]_ , \new_[22467]_ , \new_[22471]_ ,
    \new_[22472]_ , \new_[22476]_ , \new_[22477]_ , \new_[22478]_ ,
    \new_[22482]_ , \new_[22483]_ , \new_[22487]_ , \new_[22488]_ ,
    \new_[22489]_ , \new_[22493]_ , \new_[22494]_ , \new_[22498]_ ,
    \new_[22499]_ , \new_[22500]_ , \new_[22504]_ , \new_[22505]_ ,
    \new_[22509]_ , \new_[22510]_ , \new_[22511]_ , \new_[22515]_ ,
    \new_[22516]_ , \new_[22520]_ , \new_[22521]_ , \new_[22522]_ ,
    \new_[22526]_ , \new_[22527]_ , \new_[22531]_ , \new_[22532]_ ,
    \new_[22533]_ , \new_[22537]_ , \new_[22538]_ , \new_[22542]_ ,
    \new_[22543]_ , \new_[22544]_ , \new_[22548]_ , \new_[22549]_ ,
    \new_[22553]_ , \new_[22554]_ , \new_[22555]_ , \new_[22559]_ ,
    \new_[22560]_ , \new_[22564]_ , \new_[22565]_ , \new_[22566]_ ,
    \new_[22570]_ , \new_[22571]_ , \new_[22575]_ , \new_[22576]_ ,
    \new_[22577]_ , \new_[22581]_ , \new_[22582]_ , \new_[22586]_ ,
    \new_[22587]_ , \new_[22588]_ , \new_[22592]_ , \new_[22593]_ ,
    \new_[22597]_ , \new_[22598]_ , \new_[22599]_ , \new_[22603]_ ,
    \new_[22604]_ , \new_[22608]_ , \new_[22609]_ , \new_[22610]_ ,
    \new_[22614]_ , \new_[22615]_ , \new_[22619]_ , \new_[22620]_ ,
    \new_[22621]_ , \new_[22625]_ , \new_[22626]_ , \new_[22630]_ ,
    \new_[22631]_ , \new_[22632]_ , \new_[22636]_ , \new_[22637]_ ,
    \new_[22641]_ , \new_[22642]_ , \new_[22643]_ , \new_[22647]_ ,
    \new_[22648]_ , \new_[22652]_ , \new_[22653]_ , \new_[22654]_ ,
    \new_[22658]_ , \new_[22659]_ , \new_[22663]_ , \new_[22664]_ ,
    \new_[22665]_ , \new_[22669]_ , \new_[22670]_ , \new_[22674]_ ,
    \new_[22675]_ , \new_[22676]_ , \new_[22680]_ , \new_[22681]_ ,
    \new_[22685]_ , \new_[22686]_ , \new_[22687]_ , \new_[22691]_ ,
    \new_[22692]_ , \new_[22696]_ , \new_[22697]_ , \new_[22698]_ ,
    \new_[22702]_ , \new_[22703]_ , \new_[22707]_ , \new_[22708]_ ,
    \new_[22709]_ , \new_[22713]_ , \new_[22714]_ , \new_[22718]_ ,
    \new_[22719]_ , \new_[22720]_ , \new_[22724]_ , \new_[22725]_ ,
    \new_[22729]_ , \new_[22730]_ , \new_[22731]_ , \new_[22735]_ ,
    \new_[22736]_ , \new_[22740]_ , \new_[22741]_ , \new_[22742]_ ,
    \new_[22746]_ , \new_[22747]_ , \new_[22751]_ , \new_[22752]_ ,
    \new_[22753]_ , \new_[22757]_ , \new_[22758]_ , \new_[22762]_ ,
    \new_[22763]_ , \new_[22764]_ , \new_[22768]_ , \new_[22769]_ ,
    \new_[22773]_ , \new_[22774]_ , \new_[22775]_ , \new_[22779]_ ,
    \new_[22780]_ , \new_[22784]_ , \new_[22785]_ , \new_[22786]_ ,
    \new_[22790]_ , \new_[22791]_ , \new_[22795]_ , \new_[22796]_ ,
    \new_[22797]_ , \new_[22801]_ , \new_[22802]_ , \new_[22806]_ ,
    \new_[22807]_ , \new_[22808]_ , \new_[22812]_ , \new_[22813]_ ,
    \new_[22817]_ , \new_[22818]_ , \new_[22819]_ , \new_[22823]_ ,
    \new_[22824]_ , \new_[22828]_ , \new_[22829]_ , \new_[22830]_ ,
    \new_[22834]_ , \new_[22835]_ , \new_[22839]_ , \new_[22840]_ ,
    \new_[22841]_ , \new_[22845]_ , \new_[22846]_ , \new_[22850]_ ,
    \new_[22851]_ , \new_[22852]_ , \new_[22856]_ , \new_[22857]_ ,
    \new_[22861]_ , \new_[22862]_ , \new_[22863]_ , \new_[22867]_ ,
    \new_[22868]_ , \new_[22872]_ , \new_[22873]_ , \new_[22874]_ ,
    \new_[22878]_ , \new_[22879]_ , \new_[22883]_ , \new_[22884]_ ,
    \new_[22885]_ , \new_[22889]_ , \new_[22890]_ , \new_[22894]_ ,
    \new_[22895]_ , \new_[22896]_ , \new_[22900]_ , \new_[22901]_ ,
    \new_[22905]_ , \new_[22906]_ , \new_[22907]_ , \new_[22911]_ ,
    \new_[22912]_ , \new_[22916]_ , \new_[22917]_ , \new_[22918]_ ,
    \new_[22922]_ , \new_[22923]_ , \new_[22927]_ , \new_[22928]_ ,
    \new_[22929]_ , \new_[22933]_ , \new_[22934]_ , \new_[22938]_ ,
    \new_[22939]_ , \new_[22940]_ , \new_[22944]_ , \new_[22945]_ ,
    \new_[22949]_ , \new_[22950]_ , \new_[22951]_ , \new_[22955]_ ,
    \new_[22956]_ , \new_[22960]_ , \new_[22961]_ , \new_[22962]_ ,
    \new_[22966]_ , \new_[22967]_ , \new_[22971]_ , \new_[22972]_ ,
    \new_[22973]_ , \new_[22977]_ , \new_[22978]_ , \new_[22982]_ ,
    \new_[22983]_ , \new_[22984]_ , \new_[22988]_ , \new_[22989]_ ,
    \new_[22993]_ , \new_[22994]_ , \new_[22995]_ , \new_[22999]_ ,
    \new_[23000]_ , \new_[23004]_ , \new_[23005]_ , \new_[23006]_ ,
    \new_[23010]_ , \new_[23011]_ , \new_[23015]_ , \new_[23016]_ ,
    \new_[23017]_ , \new_[23021]_ , \new_[23022]_ , \new_[23026]_ ,
    \new_[23027]_ , \new_[23028]_ , \new_[23032]_ , \new_[23033]_ ,
    \new_[23037]_ , \new_[23038]_ , \new_[23039]_ , \new_[23043]_ ,
    \new_[23044]_ , \new_[23048]_ , \new_[23049]_ , \new_[23050]_ ,
    \new_[23054]_ , \new_[23055]_ , \new_[23059]_ , \new_[23060]_ ,
    \new_[23061]_ , \new_[23065]_ , \new_[23066]_ , \new_[23070]_ ,
    \new_[23071]_ , \new_[23072]_ , \new_[23076]_ , \new_[23077]_ ,
    \new_[23081]_ , \new_[23082]_ , \new_[23083]_ , \new_[23087]_ ,
    \new_[23088]_ , \new_[23092]_ , \new_[23093]_ , \new_[23094]_ ,
    \new_[23098]_ , \new_[23099]_ , \new_[23103]_ , \new_[23104]_ ,
    \new_[23105]_ , \new_[23109]_ , \new_[23110]_ , \new_[23114]_ ,
    \new_[23115]_ , \new_[23116]_ , \new_[23120]_ , \new_[23121]_ ,
    \new_[23125]_ , \new_[23126]_ , \new_[23127]_ , \new_[23131]_ ,
    \new_[23132]_ , \new_[23136]_ , \new_[23137]_ , \new_[23138]_ ,
    \new_[23142]_ , \new_[23143]_ , \new_[23147]_ , \new_[23148]_ ,
    \new_[23149]_ , \new_[23153]_ , \new_[23154]_ , \new_[23158]_ ,
    \new_[23159]_ , \new_[23160]_ , \new_[23164]_ , \new_[23165]_ ,
    \new_[23169]_ , \new_[23170]_ , \new_[23171]_ , \new_[23175]_ ,
    \new_[23176]_ , \new_[23180]_ , \new_[23181]_ , \new_[23182]_ ,
    \new_[23186]_ , \new_[23187]_ , \new_[23191]_ , \new_[23192]_ ,
    \new_[23193]_ , \new_[23197]_ , \new_[23198]_ , \new_[23202]_ ,
    \new_[23203]_ , \new_[23204]_ , \new_[23208]_ , \new_[23209]_ ,
    \new_[23213]_ , \new_[23214]_ , \new_[23215]_ , \new_[23219]_ ,
    \new_[23220]_ , \new_[23224]_ , \new_[23225]_ , \new_[23226]_ ,
    \new_[23230]_ , \new_[23231]_ , \new_[23235]_ , \new_[23236]_ ,
    \new_[23237]_ , \new_[23241]_ , \new_[23242]_ , \new_[23246]_ ,
    \new_[23247]_ , \new_[23248]_ , \new_[23252]_ , \new_[23253]_ ,
    \new_[23257]_ , \new_[23258]_ , \new_[23259]_ , \new_[23263]_ ,
    \new_[23264]_ , \new_[23268]_ , \new_[23269]_ , \new_[23270]_ ,
    \new_[23274]_ , \new_[23275]_ , \new_[23279]_ , \new_[23280]_ ,
    \new_[23281]_ , \new_[23285]_ , \new_[23286]_ , \new_[23290]_ ,
    \new_[23291]_ , \new_[23292]_ , \new_[23296]_ , \new_[23297]_ ,
    \new_[23301]_ , \new_[23302]_ , \new_[23303]_ , \new_[23307]_ ,
    \new_[23308]_ , \new_[23312]_ , \new_[23313]_ , \new_[23314]_ ,
    \new_[23318]_ , \new_[23319]_ , \new_[23323]_ , \new_[23324]_ ,
    \new_[23325]_ , \new_[23329]_ , \new_[23330]_ , \new_[23334]_ ,
    \new_[23335]_ , \new_[23336]_ , \new_[23340]_ , \new_[23341]_ ,
    \new_[23345]_ , \new_[23346]_ , \new_[23347]_ , \new_[23351]_ ,
    \new_[23352]_ , \new_[23356]_ , \new_[23357]_ , \new_[23358]_ ,
    \new_[23362]_ , \new_[23363]_ , \new_[23367]_ , \new_[23368]_ ,
    \new_[23369]_ , \new_[23373]_ , \new_[23374]_ , \new_[23378]_ ,
    \new_[23379]_ , \new_[23380]_ , \new_[23384]_ , \new_[23385]_ ,
    \new_[23389]_ , \new_[23390]_ , \new_[23391]_ , \new_[23395]_ ,
    \new_[23396]_ , \new_[23400]_ , \new_[23401]_ , \new_[23402]_ ,
    \new_[23406]_ , \new_[23407]_ , \new_[23411]_ , \new_[23412]_ ,
    \new_[23413]_ , \new_[23417]_ , \new_[23418]_ , \new_[23422]_ ,
    \new_[23423]_ , \new_[23424]_ , \new_[23428]_ , \new_[23429]_ ,
    \new_[23433]_ , \new_[23434]_ , \new_[23435]_ , \new_[23439]_ ,
    \new_[23440]_ , \new_[23444]_ , \new_[23445]_ , \new_[23446]_ ,
    \new_[23450]_ , \new_[23451]_ , \new_[23455]_ , \new_[23456]_ ,
    \new_[23457]_ , \new_[23461]_ , \new_[23462]_ , \new_[23466]_ ,
    \new_[23467]_ , \new_[23468]_ , \new_[23472]_ , \new_[23473]_ ,
    \new_[23477]_ , \new_[23478]_ , \new_[23479]_ , \new_[23483]_ ,
    \new_[23484]_ , \new_[23488]_ , \new_[23489]_ , \new_[23490]_ ,
    \new_[23494]_ , \new_[23495]_ , \new_[23499]_ , \new_[23500]_ ,
    \new_[23501]_ , \new_[23505]_ , \new_[23506]_ , \new_[23510]_ ,
    \new_[23511]_ , \new_[23512]_ , \new_[23516]_ , \new_[23517]_ ,
    \new_[23521]_ , \new_[23522]_ , \new_[23523]_ , \new_[23527]_ ,
    \new_[23528]_ , \new_[23532]_ , \new_[23533]_ , \new_[23534]_ ,
    \new_[23538]_ , \new_[23539]_ , \new_[23543]_ , \new_[23544]_ ,
    \new_[23545]_ , \new_[23549]_ , \new_[23550]_ , \new_[23554]_ ,
    \new_[23555]_ , \new_[23556]_ , \new_[23560]_ , \new_[23561]_ ,
    \new_[23565]_ , \new_[23566]_ , \new_[23567]_ , \new_[23571]_ ,
    \new_[23572]_ , \new_[23576]_ , \new_[23577]_ , \new_[23578]_ ,
    \new_[23582]_ , \new_[23583]_ , \new_[23587]_ , \new_[23588]_ ,
    \new_[23589]_ , \new_[23593]_ , \new_[23594]_ , \new_[23598]_ ,
    \new_[23599]_ , \new_[23600]_ , \new_[23604]_ , \new_[23605]_ ,
    \new_[23609]_ , \new_[23610]_ , \new_[23611]_ , \new_[23615]_ ,
    \new_[23616]_ , \new_[23620]_ , \new_[23621]_ , \new_[23622]_ ,
    \new_[23626]_ , \new_[23627]_ , \new_[23631]_ , \new_[23632]_ ,
    \new_[23633]_ , \new_[23637]_ , \new_[23638]_ , \new_[23642]_ ,
    \new_[23643]_ , \new_[23644]_ , \new_[23648]_ , \new_[23649]_ ,
    \new_[23653]_ , \new_[23654]_ , \new_[23655]_ , \new_[23659]_ ,
    \new_[23660]_ , \new_[23664]_ , \new_[23665]_ , \new_[23666]_ ,
    \new_[23670]_ , \new_[23671]_ , \new_[23675]_ , \new_[23676]_ ,
    \new_[23677]_ , \new_[23681]_ , \new_[23682]_ , \new_[23686]_ ,
    \new_[23687]_ , \new_[23688]_ , \new_[23692]_ , \new_[23693]_ ,
    \new_[23697]_ , \new_[23698]_ , \new_[23699]_ , \new_[23703]_ ,
    \new_[23704]_ , \new_[23708]_ , \new_[23709]_ , \new_[23710]_ ,
    \new_[23714]_ , \new_[23715]_ , \new_[23719]_ , \new_[23720]_ ,
    \new_[23721]_ , \new_[23725]_ , \new_[23726]_ , \new_[23730]_ ,
    \new_[23731]_ , \new_[23732]_ , \new_[23736]_ , \new_[23737]_ ,
    \new_[23741]_ , \new_[23742]_ , \new_[23743]_ , \new_[23747]_ ,
    \new_[23748]_ , \new_[23752]_ , \new_[23753]_ , \new_[23754]_ ,
    \new_[23758]_ , \new_[23759]_ , \new_[23763]_ , \new_[23764]_ ,
    \new_[23765]_ , \new_[23769]_ , \new_[23770]_ , \new_[23774]_ ,
    \new_[23775]_ , \new_[23776]_ , \new_[23780]_ , \new_[23781]_ ,
    \new_[23785]_ , \new_[23786]_ , \new_[23787]_ , \new_[23791]_ ,
    \new_[23792]_ , \new_[23796]_ , \new_[23797]_ , \new_[23798]_ ,
    \new_[23802]_ , \new_[23803]_ , \new_[23807]_ , \new_[23808]_ ,
    \new_[23809]_ , \new_[23813]_ , \new_[23814]_ , \new_[23818]_ ,
    \new_[23819]_ , \new_[23820]_ , \new_[23824]_ , \new_[23825]_ ,
    \new_[23829]_ , \new_[23830]_ , \new_[23831]_ , \new_[23835]_ ,
    \new_[23836]_ , \new_[23840]_ , \new_[23841]_ , \new_[23842]_ ,
    \new_[23846]_ , \new_[23847]_ , \new_[23851]_ , \new_[23852]_ ,
    \new_[23853]_ , \new_[23857]_ , \new_[23858]_ , \new_[23862]_ ,
    \new_[23863]_ , \new_[23864]_ , \new_[23868]_ , \new_[23869]_ ,
    \new_[23873]_ , \new_[23874]_ , \new_[23875]_ , \new_[23879]_ ,
    \new_[23880]_ , \new_[23884]_ , \new_[23885]_ , \new_[23886]_ ,
    \new_[23890]_ , \new_[23891]_ , \new_[23895]_ , \new_[23896]_ ,
    \new_[23897]_ , \new_[23901]_ , \new_[23902]_ , \new_[23906]_ ,
    \new_[23907]_ , \new_[23908]_ , \new_[23912]_ , \new_[23913]_ ,
    \new_[23917]_ , \new_[23918]_ , \new_[23919]_ , \new_[23923]_ ,
    \new_[23924]_ , \new_[23928]_ , \new_[23929]_ , \new_[23930]_ ,
    \new_[23934]_ , \new_[23935]_ , \new_[23939]_ , \new_[23940]_ ,
    \new_[23941]_ , \new_[23945]_ , \new_[23946]_ , \new_[23950]_ ,
    \new_[23951]_ , \new_[23952]_ , \new_[23956]_ , \new_[23957]_ ,
    \new_[23961]_ , \new_[23962]_ , \new_[23963]_ , \new_[23967]_ ,
    \new_[23968]_ , \new_[23972]_ , \new_[23973]_ , \new_[23974]_ ,
    \new_[23978]_ , \new_[23979]_ , \new_[23983]_ , \new_[23984]_ ,
    \new_[23985]_ , \new_[23989]_ , \new_[23990]_ , \new_[23994]_ ,
    \new_[23995]_ , \new_[23996]_ , \new_[24000]_ , \new_[24001]_ ,
    \new_[24005]_ , \new_[24006]_ , \new_[24007]_ , \new_[24011]_ ,
    \new_[24012]_ , \new_[24016]_ , \new_[24017]_ , \new_[24018]_ ,
    \new_[24022]_ , \new_[24023]_ , \new_[24027]_ , \new_[24028]_ ,
    \new_[24029]_ , \new_[24033]_ , \new_[24034]_ , \new_[24038]_ ,
    \new_[24039]_ , \new_[24040]_ , \new_[24044]_ , \new_[24045]_ ,
    \new_[24049]_ , \new_[24050]_ , \new_[24051]_ , \new_[24055]_ ,
    \new_[24056]_ , \new_[24060]_ , \new_[24061]_ , \new_[24062]_ ,
    \new_[24066]_ , \new_[24067]_ , \new_[24071]_ , \new_[24072]_ ,
    \new_[24073]_ , \new_[24077]_ , \new_[24078]_ , \new_[24082]_ ,
    \new_[24083]_ , \new_[24084]_ , \new_[24088]_ , \new_[24089]_ ,
    \new_[24093]_ , \new_[24094]_ , \new_[24095]_ , \new_[24099]_ ,
    \new_[24100]_ , \new_[24104]_ , \new_[24105]_ , \new_[24106]_ ,
    \new_[24110]_ , \new_[24111]_ , \new_[24115]_ , \new_[24116]_ ,
    \new_[24117]_ , \new_[24121]_ , \new_[24122]_ , \new_[24126]_ ,
    \new_[24127]_ , \new_[24128]_ , \new_[24132]_ , \new_[24133]_ ,
    \new_[24137]_ , \new_[24138]_ , \new_[24139]_ , \new_[24143]_ ,
    \new_[24144]_ , \new_[24148]_ , \new_[24149]_ , \new_[24150]_ ,
    \new_[24154]_ , \new_[24155]_ , \new_[24159]_ , \new_[24160]_ ,
    \new_[24161]_ , \new_[24165]_ , \new_[24166]_ , \new_[24170]_ ,
    \new_[24171]_ , \new_[24172]_ , \new_[24176]_ , \new_[24177]_ ,
    \new_[24181]_ , \new_[24182]_ , \new_[24183]_ , \new_[24187]_ ,
    \new_[24188]_ , \new_[24192]_ , \new_[24193]_ , \new_[24194]_ ,
    \new_[24198]_ , \new_[24199]_ , \new_[24203]_ , \new_[24204]_ ,
    \new_[24205]_ , \new_[24209]_ , \new_[24210]_ , \new_[24214]_ ,
    \new_[24215]_ , \new_[24216]_ , \new_[24220]_ , \new_[24221]_ ,
    \new_[24225]_ , \new_[24226]_ , \new_[24227]_ , \new_[24231]_ ,
    \new_[24232]_ , \new_[24236]_ , \new_[24237]_ , \new_[24238]_ ,
    \new_[24242]_ , \new_[24243]_ , \new_[24247]_ , \new_[24248]_ ,
    \new_[24249]_ , \new_[24253]_ , \new_[24254]_ , \new_[24258]_ ,
    \new_[24259]_ , \new_[24260]_ , \new_[24264]_ , \new_[24265]_ ,
    \new_[24269]_ , \new_[24270]_ , \new_[24271]_ , \new_[24275]_ ,
    \new_[24276]_ , \new_[24280]_ , \new_[24281]_ , \new_[24282]_ ,
    \new_[24286]_ , \new_[24287]_ , \new_[24291]_ , \new_[24292]_ ,
    \new_[24293]_ , \new_[24297]_ , \new_[24298]_ , \new_[24302]_ ,
    \new_[24303]_ , \new_[24304]_ , \new_[24308]_ , \new_[24309]_ ,
    \new_[24313]_ , \new_[24314]_ , \new_[24315]_ , \new_[24319]_ ,
    \new_[24320]_ , \new_[24324]_ , \new_[24325]_ , \new_[24326]_ ,
    \new_[24330]_ , \new_[24331]_ , \new_[24335]_ , \new_[24336]_ ,
    \new_[24337]_ , \new_[24341]_ , \new_[24342]_ , \new_[24346]_ ,
    \new_[24347]_ , \new_[24348]_ , \new_[24352]_ , \new_[24353]_ ,
    \new_[24357]_ , \new_[24358]_ , \new_[24359]_ , \new_[24363]_ ,
    \new_[24364]_ , \new_[24368]_ , \new_[24369]_ , \new_[24370]_ ,
    \new_[24374]_ , \new_[24375]_ , \new_[24379]_ , \new_[24380]_ ,
    \new_[24381]_ , \new_[24385]_ , \new_[24386]_ , \new_[24390]_ ,
    \new_[24391]_ , \new_[24392]_ , \new_[24396]_ , \new_[24397]_ ,
    \new_[24401]_ , \new_[24402]_ , \new_[24403]_ , \new_[24407]_ ,
    \new_[24408]_ , \new_[24412]_ , \new_[24413]_ , \new_[24414]_ ,
    \new_[24418]_ , \new_[24419]_ , \new_[24423]_ , \new_[24424]_ ,
    \new_[24425]_ , \new_[24429]_ , \new_[24430]_ , \new_[24434]_ ,
    \new_[24435]_ , \new_[24436]_ , \new_[24440]_ , \new_[24441]_ ,
    \new_[24445]_ , \new_[24446]_ , \new_[24447]_ , \new_[24451]_ ,
    \new_[24452]_ , \new_[24456]_ , \new_[24457]_ , \new_[24458]_ ,
    \new_[24462]_ , \new_[24463]_ , \new_[24467]_ , \new_[24468]_ ,
    \new_[24469]_ , \new_[24473]_ , \new_[24474]_ , \new_[24478]_ ,
    \new_[24479]_ , \new_[24480]_ , \new_[24484]_ , \new_[24485]_ ,
    \new_[24489]_ , \new_[24490]_ , \new_[24491]_ , \new_[24495]_ ,
    \new_[24496]_ , \new_[24500]_ , \new_[24501]_ , \new_[24502]_ ,
    \new_[24506]_ , \new_[24507]_ , \new_[24511]_ , \new_[24512]_ ,
    \new_[24513]_ , \new_[24517]_ , \new_[24518]_ , \new_[24522]_ ,
    \new_[24523]_ , \new_[24524]_ , \new_[24528]_ , \new_[24529]_ ,
    \new_[24533]_ , \new_[24534]_ , \new_[24535]_ , \new_[24539]_ ,
    \new_[24540]_ , \new_[24544]_ , \new_[24545]_ , \new_[24546]_ ,
    \new_[24550]_ , \new_[24551]_ , \new_[24555]_ , \new_[24556]_ ,
    \new_[24557]_ , \new_[24561]_ , \new_[24562]_ , \new_[24566]_ ,
    \new_[24567]_ , \new_[24568]_ , \new_[24572]_ , \new_[24573]_ ,
    \new_[24577]_ , \new_[24578]_ , \new_[24579]_ , \new_[24583]_ ,
    \new_[24584]_ , \new_[24588]_ , \new_[24589]_ , \new_[24590]_ ,
    \new_[24594]_ , \new_[24595]_ , \new_[24599]_ , \new_[24600]_ ,
    \new_[24601]_ , \new_[24605]_ , \new_[24606]_ , \new_[24610]_ ,
    \new_[24611]_ , \new_[24612]_ , \new_[24616]_ , \new_[24617]_ ,
    \new_[24621]_ , \new_[24622]_ , \new_[24623]_ , \new_[24627]_ ,
    \new_[24628]_ , \new_[24632]_ , \new_[24633]_ , \new_[24634]_ ,
    \new_[24638]_ , \new_[24639]_ , \new_[24643]_ , \new_[24644]_ ,
    \new_[24645]_ , \new_[24649]_ , \new_[24650]_ , \new_[24654]_ ,
    \new_[24655]_ , \new_[24656]_ , \new_[24660]_ , \new_[24661]_ ,
    \new_[24665]_ , \new_[24666]_ , \new_[24667]_ , \new_[24671]_ ,
    \new_[24672]_ , \new_[24676]_ , \new_[24677]_ , \new_[24678]_ ,
    \new_[24682]_ , \new_[24683]_ , \new_[24687]_ , \new_[24688]_ ,
    \new_[24689]_ , \new_[24693]_ , \new_[24694]_ , \new_[24698]_ ,
    \new_[24699]_ , \new_[24700]_ , \new_[24704]_ , \new_[24705]_ ,
    \new_[24709]_ , \new_[24710]_ , \new_[24711]_ , \new_[24715]_ ,
    \new_[24716]_ , \new_[24720]_ , \new_[24721]_ , \new_[24722]_ ,
    \new_[24726]_ , \new_[24727]_ , \new_[24731]_ , \new_[24732]_ ,
    \new_[24733]_ , \new_[24737]_ , \new_[24738]_ , \new_[24742]_ ,
    \new_[24743]_ , \new_[24744]_ , \new_[24748]_ , \new_[24749]_ ,
    \new_[24753]_ , \new_[24754]_ , \new_[24755]_ , \new_[24759]_ ,
    \new_[24760]_ , \new_[24764]_ , \new_[24765]_ , \new_[24766]_ ,
    \new_[24770]_ , \new_[24771]_ , \new_[24775]_ , \new_[24776]_ ,
    \new_[24777]_ , \new_[24781]_ , \new_[24782]_ , \new_[24786]_ ,
    \new_[24787]_ , \new_[24788]_ , \new_[24792]_ , \new_[24793]_ ,
    \new_[24797]_ , \new_[24798]_ , \new_[24799]_ , \new_[24803]_ ,
    \new_[24804]_ , \new_[24808]_ , \new_[24809]_ , \new_[24810]_ ,
    \new_[24814]_ , \new_[24815]_ , \new_[24819]_ , \new_[24820]_ ,
    \new_[24821]_ , \new_[24825]_ , \new_[24826]_ , \new_[24830]_ ,
    \new_[24831]_ , \new_[24832]_ , \new_[24836]_ , \new_[24837]_ ,
    \new_[24841]_ , \new_[24842]_ , \new_[24843]_ , \new_[24847]_ ,
    \new_[24848]_ , \new_[24852]_ , \new_[24853]_ , \new_[24854]_ ,
    \new_[24858]_ , \new_[24859]_ , \new_[24863]_ , \new_[24864]_ ,
    \new_[24865]_ , \new_[24869]_ , \new_[24870]_ , \new_[24874]_ ,
    \new_[24875]_ , \new_[24876]_ , \new_[24880]_ , \new_[24881]_ ,
    \new_[24885]_ , \new_[24886]_ , \new_[24887]_ , \new_[24891]_ ,
    \new_[24892]_ , \new_[24896]_ , \new_[24897]_ , \new_[24898]_ ,
    \new_[24902]_ , \new_[24903]_ , \new_[24907]_ , \new_[24908]_ ,
    \new_[24909]_ , \new_[24913]_ , \new_[24914]_ , \new_[24918]_ ,
    \new_[24919]_ , \new_[24920]_ , \new_[24924]_ , \new_[24925]_ ,
    \new_[24929]_ , \new_[24930]_ , \new_[24931]_ , \new_[24935]_ ,
    \new_[24936]_ , \new_[24940]_ , \new_[24941]_ , \new_[24942]_ ,
    \new_[24946]_ , \new_[24947]_ , \new_[24951]_ , \new_[24952]_ ,
    \new_[24953]_ , \new_[24957]_ , \new_[24958]_ , \new_[24962]_ ,
    \new_[24963]_ , \new_[24964]_ , \new_[24968]_ , \new_[24969]_ ,
    \new_[24973]_ , \new_[24974]_ , \new_[24975]_ , \new_[24979]_ ,
    \new_[24980]_ , \new_[24984]_ , \new_[24985]_ , \new_[24986]_ ,
    \new_[24990]_ , \new_[24991]_ , \new_[24995]_ , \new_[24996]_ ,
    \new_[24997]_ , \new_[25001]_ , \new_[25002]_ , \new_[25006]_ ,
    \new_[25007]_ , \new_[25008]_ , \new_[25012]_ , \new_[25013]_ ,
    \new_[25017]_ , \new_[25018]_ , \new_[25019]_ , \new_[25023]_ ,
    \new_[25024]_ , \new_[25028]_ , \new_[25029]_ , \new_[25030]_ ,
    \new_[25034]_ , \new_[25035]_ , \new_[25039]_ , \new_[25040]_ ,
    \new_[25041]_ , \new_[25045]_ , \new_[25046]_ , \new_[25050]_ ,
    \new_[25051]_ , \new_[25052]_ , \new_[25056]_ , \new_[25057]_ ,
    \new_[25061]_ , \new_[25062]_ , \new_[25063]_ , \new_[25067]_ ,
    \new_[25068]_ , \new_[25072]_ , \new_[25073]_ , \new_[25074]_ ,
    \new_[25078]_ , \new_[25079]_ , \new_[25083]_ , \new_[25084]_ ,
    \new_[25085]_ , \new_[25089]_ , \new_[25090]_ , \new_[25094]_ ,
    \new_[25095]_ , \new_[25096]_ , \new_[25100]_ , \new_[25101]_ ,
    \new_[25105]_ , \new_[25106]_ , \new_[25107]_ , \new_[25111]_ ,
    \new_[25112]_ , \new_[25116]_ , \new_[25117]_ , \new_[25118]_ ,
    \new_[25122]_ , \new_[25123]_ , \new_[25127]_ , \new_[25128]_ ,
    \new_[25129]_ , \new_[25133]_ , \new_[25134]_ , \new_[25138]_ ,
    \new_[25139]_ , \new_[25140]_ , \new_[25144]_ , \new_[25145]_ ,
    \new_[25149]_ , \new_[25150]_ , \new_[25151]_ , \new_[25155]_ ,
    \new_[25156]_ , \new_[25160]_ , \new_[25161]_ , \new_[25162]_ ,
    \new_[25166]_ , \new_[25167]_ , \new_[25171]_ , \new_[25172]_ ,
    \new_[25173]_ , \new_[25177]_ , \new_[25178]_ , \new_[25182]_ ,
    \new_[25183]_ , \new_[25184]_ , \new_[25188]_ , \new_[25189]_ ,
    \new_[25193]_ , \new_[25194]_ , \new_[25195]_ , \new_[25199]_ ,
    \new_[25200]_ , \new_[25204]_ , \new_[25205]_ , \new_[25206]_ ,
    \new_[25210]_ , \new_[25211]_ , \new_[25215]_ , \new_[25216]_ ,
    \new_[25217]_ , \new_[25221]_ , \new_[25222]_ , \new_[25226]_ ,
    \new_[25227]_ , \new_[25228]_ , \new_[25232]_ , \new_[25233]_ ,
    \new_[25237]_ , \new_[25238]_ , \new_[25239]_ , \new_[25243]_ ,
    \new_[25244]_ , \new_[25248]_ , \new_[25249]_ , \new_[25250]_ ,
    \new_[25254]_ , \new_[25255]_ , \new_[25259]_ , \new_[25260]_ ,
    \new_[25261]_ , \new_[25265]_ , \new_[25266]_ , \new_[25270]_ ,
    \new_[25271]_ , \new_[25272]_ , \new_[25276]_ , \new_[25277]_ ,
    \new_[25281]_ , \new_[25282]_ , \new_[25283]_ , \new_[25287]_ ,
    \new_[25288]_ , \new_[25292]_ , \new_[25293]_ , \new_[25294]_ ,
    \new_[25298]_ , \new_[25299]_ , \new_[25303]_ , \new_[25304]_ ,
    \new_[25305]_ , \new_[25309]_ , \new_[25310]_ , \new_[25314]_ ,
    \new_[25315]_ , \new_[25316]_ , \new_[25320]_ , \new_[25321]_ ,
    \new_[25325]_ , \new_[25326]_ , \new_[25327]_ , \new_[25331]_ ,
    \new_[25332]_ , \new_[25336]_ , \new_[25337]_ , \new_[25338]_ ,
    \new_[25342]_ , \new_[25343]_ , \new_[25347]_ , \new_[25348]_ ,
    \new_[25349]_ , \new_[25353]_ , \new_[25354]_ , \new_[25358]_ ,
    \new_[25359]_ , \new_[25360]_ , \new_[25364]_ , \new_[25365]_ ,
    \new_[25369]_ , \new_[25370]_ , \new_[25371]_ , \new_[25375]_ ,
    \new_[25376]_ , \new_[25380]_ , \new_[25381]_ , \new_[25382]_ ,
    \new_[25386]_ , \new_[25387]_ , \new_[25391]_ , \new_[25392]_ ,
    \new_[25393]_ , \new_[25397]_ , \new_[25398]_ , \new_[25402]_ ,
    \new_[25403]_ , \new_[25404]_ , \new_[25408]_ , \new_[25409]_ ,
    \new_[25413]_ , \new_[25414]_ , \new_[25415]_ , \new_[25419]_ ,
    \new_[25420]_ , \new_[25424]_ , \new_[25425]_ , \new_[25426]_ ,
    \new_[25430]_ , \new_[25431]_ , \new_[25435]_ , \new_[25436]_ ,
    \new_[25437]_ , \new_[25441]_ , \new_[25442]_ , \new_[25446]_ ,
    \new_[25447]_ , \new_[25448]_ , \new_[25452]_ , \new_[25453]_ ,
    \new_[25457]_ , \new_[25458]_ , \new_[25459]_ , \new_[25463]_ ,
    \new_[25464]_ , \new_[25468]_ , \new_[25469]_ , \new_[25470]_ ,
    \new_[25474]_ , \new_[25475]_ , \new_[25479]_ , \new_[25480]_ ,
    \new_[25481]_ , \new_[25485]_ , \new_[25486]_ , \new_[25490]_ ,
    \new_[25491]_ , \new_[25492]_ , \new_[25496]_ , \new_[25497]_ ,
    \new_[25501]_ , \new_[25502]_ , \new_[25503]_ , \new_[25507]_ ,
    \new_[25508]_ , \new_[25512]_ , \new_[25513]_ , \new_[25514]_ ,
    \new_[25518]_ , \new_[25519]_ , \new_[25523]_ , \new_[25524]_ ,
    \new_[25525]_ , \new_[25529]_ , \new_[25530]_ , \new_[25534]_ ,
    \new_[25535]_ , \new_[25536]_ , \new_[25540]_ , \new_[25541]_ ,
    \new_[25545]_ , \new_[25546]_ , \new_[25547]_ , \new_[25551]_ ,
    \new_[25552]_ , \new_[25556]_ , \new_[25557]_ , \new_[25558]_ ,
    \new_[25562]_ , \new_[25563]_ , \new_[25567]_ , \new_[25568]_ ,
    \new_[25569]_ , \new_[25573]_ , \new_[25574]_ , \new_[25578]_ ,
    \new_[25579]_ , \new_[25580]_ , \new_[25584]_ , \new_[25585]_ ,
    \new_[25589]_ , \new_[25590]_ , \new_[25591]_ , \new_[25595]_ ,
    \new_[25596]_ , \new_[25600]_ , \new_[25601]_ , \new_[25602]_ ,
    \new_[25606]_ , \new_[25607]_ , \new_[25611]_ , \new_[25612]_ ,
    \new_[25613]_ , \new_[25617]_ , \new_[25618]_ , \new_[25622]_ ,
    \new_[25623]_ , \new_[25624]_ , \new_[25628]_ , \new_[25629]_ ,
    \new_[25633]_ , \new_[25634]_ , \new_[25635]_ , \new_[25639]_ ,
    \new_[25640]_ , \new_[25644]_ , \new_[25645]_ , \new_[25646]_ ,
    \new_[25650]_ , \new_[25651]_ , \new_[25655]_ , \new_[25656]_ ,
    \new_[25657]_ , \new_[25661]_ , \new_[25662]_ , \new_[25666]_ ,
    \new_[25667]_ , \new_[25668]_ , \new_[25672]_ , \new_[25673]_ ,
    \new_[25677]_ , \new_[25678]_ , \new_[25679]_ , \new_[25683]_ ,
    \new_[25684]_ , \new_[25688]_ , \new_[25689]_ , \new_[25690]_ ,
    \new_[25694]_ , \new_[25695]_ , \new_[25699]_ , \new_[25700]_ ,
    \new_[25701]_ , \new_[25705]_ , \new_[25706]_ , \new_[25710]_ ,
    \new_[25711]_ , \new_[25712]_ , \new_[25716]_ , \new_[25717]_ ,
    \new_[25721]_ , \new_[25722]_ , \new_[25723]_ , \new_[25727]_ ,
    \new_[25728]_ , \new_[25732]_ , \new_[25733]_ , \new_[25734]_ ,
    \new_[25738]_ , \new_[25739]_ , \new_[25743]_ , \new_[25744]_ ,
    \new_[25745]_ , \new_[25749]_ , \new_[25750]_ , \new_[25754]_ ,
    \new_[25755]_ , \new_[25756]_ , \new_[25760]_ , \new_[25761]_ ,
    \new_[25765]_ , \new_[25766]_ , \new_[25767]_ , \new_[25771]_ ,
    \new_[25772]_ , \new_[25776]_ , \new_[25777]_ , \new_[25778]_ ,
    \new_[25782]_ , \new_[25783]_ , \new_[25787]_ , \new_[25788]_ ,
    \new_[25789]_ , \new_[25793]_ , \new_[25794]_ , \new_[25798]_ ,
    \new_[25799]_ , \new_[25800]_ , \new_[25804]_ , \new_[25805]_ ,
    \new_[25809]_ , \new_[25810]_ , \new_[25811]_ , \new_[25815]_ ,
    \new_[25816]_ , \new_[25820]_ , \new_[25821]_ , \new_[25822]_ ,
    \new_[25826]_ , \new_[25827]_ , \new_[25831]_ , \new_[25832]_ ,
    \new_[25833]_ , \new_[25837]_ , \new_[25838]_ , \new_[25842]_ ,
    \new_[25843]_ , \new_[25844]_ , \new_[25848]_ , \new_[25849]_ ,
    \new_[25853]_ , \new_[25854]_ , \new_[25855]_ , \new_[25859]_ ,
    \new_[25860]_ , \new_[25864]_ , \new_[25865]_ , \new_[25866]_ ,
    \new_[25870]_ , \new_[25871]_ , \new_[25875]_ , \new_[25876]_ ,
    \new_[25877]_ , \new_[25881]_ , \new_[25882]_ , \new_[25886]_ ,
    \new_[25887]_ , \new_[25888]_ , \new_[25892]_ , \new_[25893]_ ,
    \new_[25897]_ , \new_[25898]_ , \new_[25899]_ , \new_[25903]_ ,
    \new_[25904]_ , \new_[25908]_ , \new_[25909]_ , \new_[25910]_ ,
    \new_[25914]_ , \new_[25915]_ , \new_[25919]_ , \new_[25920]_ ,
    \new_[25921]_ , \new_[25925]_ , \new_[25926]_ , \new_[25930]_ ,
    \new_[25931]_ , \new_[25932]_ , \new_[25936]_ , \new_[25937]_ ,
    \new_[25941]_ , \new_[25942]_ , \new_[25943]_ , \new_[25947]_ ,
    \new_[25948]_ , \new_[25952]_ , \new_[25953]_ , \new_[25954]_ ,
    \new_[25958]_ , \new_[25959]_ , \new_[25963]_ , \new_[25964]_ ,
    \new_[25965]_ , \new_[25969]_ , \new_[25970]_ , \new_[25974]_ ,
    \new_[25975]_ , \new_[25976]_ , \new_[25980]_ , \new_[25981]_ ,
    \new_[25985]_ , \new_[25986]_ , \new_[25987]_ , \new_[25991]_ ,
    \new_[25992]_ , \new_[25996]_ , \new_[25997]_ , \new_[25998]_ ,
    \new_[26002]_ , \new_[26003]_ , \new_[26007]_ , \new_[26008]_ ,
    \new_[26009]_ , \new_[26013]_ , \new_[26014]_ , \new_[26018]_ ,
    \new_[26019]_ , \new_[26020]_ , \new_[26024]_ , \new_[26025]_ ,
    \new_[26029]_ , \new_[26030]_ , \new_[26031]_ , \new_[26035]_ ,
    \new_[26036]_ , \new_[26040]_ , \new_[26041]_ , \new_[26042]_ ,
    \new_[26046]_ , \new_[26047]_ , \new_[26051]_ , \new_[26052]_ ,
    \new_[26053]_ , \new_[26057]_ , \new_[26058]_ , \new_[26062]_ ,
    \new_[26063]_ , \new_[26064]_ , \new_[26068]_ , \new_[26069]_ ,
    \new_[26073]_ , \new_[26074]_ , \new_[26075]_ , \new_[26079]_ ,
    \new_[26080]_ , \new_[26084]_ , \new_[26085]_ , \new_[26086]_ ,
    \new_[26090]_ , \new_[26091]_ , \new_[26095]_ , \new_[26096]_ ,
    \new_[26097]_ , \new_[26101]_ , \new_[26102]_ , \new_[26106]_ ,
    \new_[26107]_ , \new_[26108]_ , \new_[26112]_ , \new_[26113]_ ,
    \new_[26117]_ , \new_[26118]_ , \new_[26119]_ , \new_[26123]_ ,
    \new_[26124]_ , \new_[26128]_ , \new_[26129]_ , \new_[26130]_ ,
    \new_[26134]_ , \new_[26135]_ , \new_[26139]_ , \new_[26140]_ ,
    \new_[26141]_ , \new_[26145]_ , \new_[26146]_ , \new_[26150]_ ,
    \new_[26151]_ , \new_[26152]_ , \new_[26156]_ , \new_[26157]_ ,
    \new_[26161]_ , \new_[26162]_ , \new_[26163]_ , \new_[26167]_ ,
    \new_[26168]_ , \new_[26172]_ , \new_[26173]_ , \new_[26174]_ ,
    \new_[26178]_ , \new_[26179]_ , \new_[26183]_ , \new_[26184]_ ,
    \new_[26185]_ , \new_[26189]_ , \new_[26190]_ , \new_[26194]_ ,
    \new_[26195]_ , \new_[26196]_ , \new_[26200]_ , \new_[26201]_ ,
    \new_[26205]_ , \new_[26206]_ , \new_[26207]_ , \new_[26211]_ ,
    \new_[26212]_ , \new_[26216]_ , \new_[26217]_ , \new_[26218]_ ,
    \new_[26222]_ , \new_[26223]_ , \new_[26227]_ , \new_[26228]_ ,
    \new_[26229]_ , \new_[26233]_ , \new_[26234]_ , \new_[26238]_ ,
    \new_[26239]_ , \new_[26240]_ , \new_[26244]_ , \new_[26245]_ ,
    \new_[26249]_ , \new_[26250]_ , \new_[26251]_ , \new_[26255]_ ,
    \new_[26256]_ , \new_[26260]_ , \new_[26261]_ , \new_[26262]_ ,
    \new_[26266]_ , \new_[26267]_ , \new_[26271]_ , \new_[26272]_ ,
    \new_[26273]_ , \new_[26277]_ , \new_[26278]_ , \new_[26282]_ ,
    \new_[26283]_ , \new_[26284]_ , \new_[26288]_ , \new_[26289]_ ,
    \new_[26293]_ , \new_[26294]_ , \new_[26295]_ , \new_[26299]_ ,
    \new_[26300]_ , \new_[26304]_ , \new_[26305]_ , \new_[26306]_ ,
    \new_[26310]_ , \new_[26311]_ , \new_[26315]_ , \new_[26316]_ ,
    \new_[26317]_ , \new_[26321]_ , \new_[26322]_ , \new_[26326]_ ,
    \new_[26327]_ , \new_[26328]_ , \new_[26332]_ , \new_[26333]_ ,
    \new_[26337]_ , \new_[26338]_ , \new_[26339]_ , \new_[26343]_ ,
    \new_[26344]_ , \new_[26348]_ , \new_[26349]_ , \new_[26350]_ ,
    \new_[26354]_ , \new_[26355]_ , \new_[26359]_ , \new_[26360]_ ,
    \new_[26361]_ , \new_[26365]_ , \new_[26366]_ , \new_[26370]_ ,
    \new_[26371]_ , \new_[26372]_ , \new_[26376]_ , \new_[26377]_ ,
    \new_[26381]_ , \new_[26382]_ , \new_[26383]_ , \new_[26387]_ ,
    \new_[26388]_ , \new_[26392]_ , \new_[26393]_ , \new_[26394]_ ,
    \new_[26398]_ , \new_[26399]_ , \new_[26403]_ , \new_[26404]_ ,
    \new_[26405]_ , \new_[26409]_ , \new_[26410]_ , \new_[26414]_ ,
    \new_[26415]_ , \new_[26416]_ , \new_[26420]_ , \new_[26421]_ ,
    \new_[26425]_ , \new_[26426]_ , \new_[26427]_ , \new_[26431]_ ,
    \new_[26432]_ , \new_[26436]_ , \new_[26437]_ , \new_[26438]_ ,
    \new_[26442]_ , \new_[26443]_ , \new_[26447]_ , \new_[26448]_ ,
    \new_[26449]_ , \new_[26453]_ , \new_[26454]_ , \new_[26458]_ ,
    \new_[26459]_ , \new_[26460]_ , \new_[26464]_ , \new_[26465]_ ,
    \new_[26469]_ , \new_[26470]_ , \new_[26471]_ , \new_[26475]_ ,
    \new_[26476]_ , \new_[26480]_ , \new_[26481]_ , \new_[26482]_ ,
    \new_[26486]_ , \new_[26487]_ , \new_[26491]_ , \new_[26492]_ ,
    \new_[26493]_ , \new_[26497]_ , \new_[26498]_ , \new_[26502]_ ,
    \new_[26503]_ , \new_[26504]_ , \new_[26508]_ , \new_[26509]_ ,
    \new_[26513]_ , \new_[26514]_ , \new_[26515]_ , \new_[26519]_ ,
    \new_[26520]_ , \new_[26524]_ , \new_[26525]_ , \new_[26526]_ ,
    \new_[26530]_ , \new_[26531]_ , \new_[26535]_ , \new_[26536]_ ,
    \new_[26537]_ , \new_[26541]_ , \new_[26542]_ , \new_[26546]_ ,
    \new_[26547]_ , \new_[26548]_ , \new_[26552]_ , \new_[26553]_ ,
    \new_[26557]_ , \new_[26558]_ , \new_[26559]_ , \new_[26563]_ ,
    \new_[26564]_ , \new_[26568]_ , \new_[26569]_ , \new_[26570]_ ,
    \new_[26574]_ , \new_[26575]_ , \new_[26579]_ , \new_[26580]_ ,
    \new_[26581]_ , \new_[26585]_ , \new_[26586]_ , \new_[26590]_ ,
    \new_[26591]_ , \new_[26592]_ , \new_[26596]_ , \new_[26597]_ ,
    \new_[26601]_ , \new_[26602]_ , \new_[26603]_ , \new_[26607]_ ,
    \new_[26608]_ , \new_[26612]_ , \new_[26613]_ , \new_[26614]_ ,
    \new_[26618]_ , \new_[26619]_ , \new_[26623]_ , \new_[26624]_ ,
    \new_[26625]_ , \new_[26629]_ , \new_[26630]_ , \new_[26634]_ ,
    \new_[26635]_ , \new_[26636]_ , \new_[26640]_ , \new_[26641]_ ,
    \new_[26645]_ , \new_[26646]_ , \new_[26647]_ , \new_[26651]_ ,
    \new_[26652]_ , \new_[26656]_ , \new_[26657]_ , \new_[26658]_ ,
    \new_[26662]_ , \new_[26663]_ , \new_[26667]_ , \new_[26668]_ ,
    \new_[26669]_ , \new_[26673]_ , \new_[26674]_ , \new_[26678]_ ,
    \new_[26679]_ , \new_[26680]_ , \new_[26684]_ , \new_[26685]_ ,
    \new_[26689]_ , \new_[26690]_ , \new_[26691]_ , \new_[26695]_ ,
    \new_[26696]_ , \new_[26700]_ , \new_[26701]_ , \new_[26702]_ ,
    \new_[26706]_ , \new_[26707]_ , \new_[26711]_ , \new_[26712]_ ,
    \new_[26713]_ , \new_[26717]_ , \new_[26718]_ , \new_[26722]_ ,
    \new_[26723]_ , \new_[26724]_ , \new_[26728]_ , \new_[26729]_ ,
    \new_[26733]_ , \new_[26734]_ , \new_[26735]_ , \new_[26739]_ ,
    \new_[26740]_ , \new_[26744]_ , \new_[26745]_ , \new_[26746]_ ,
    \new_[26750]_ , \new_[26751]_ , \new_[26755]_ , \new_[26756]_ ,
    \new_[26757]_ , \new_[26761]_ , \new_[26762]_ , \new_[26766]_ ,
    \new_[26767]_ , \new_[26768]_ , \new_[26772]_ , \new_[26773]_ ,
    \new_[26777]_ , \new_[26778]_ , \new_[26779]_ , \new_[26783]_ ,
    \new_[26784]_ , \new_[26788]_ , \new_[26789]_ , \new_[26790]_ ,
    \new_[26794]_ , \new_[26795]_ , \new_[26799]_ , \new_[26800]_ ,
    \new_[26801]_ , \new_[26805]_ , \new_[26806]_ , \new_[26810]_ ,
    \new_[26811]_ , \new_[26812]_ , \new_[26816]_ , \new_[26817]_ ,
    \new_[26821]_ , \new_[26822]_ , \new_[26823]_ , \new_[26827]_ ,
    \new_[26828]_ , \new_[26832]_ , \new_[26833]_ , \new_[26834]_ ,
    \new_[26838]_ , \new_[26839]_ , \new_[26843]_ , \new_[26844]_ ,
    \new_[26845]_ , \new_[26849]_ , \new_[26850]_ , \new_[26854]_ ,
    \new_[26855]_ , \new_[26856]_ , \new_[26860]_ , \new_[26861]_ ,
    \new_[26865]_ , \new_[26866]_ , \new_[26867]_ , \new_[26871]_ ,
    \new_[26872]_ , \new_[26876]_ , \new_[26877]_ , \new_[26878]_ ,
    \new_[26882]_ , \new_[26883]_ , \new_[26887]_ , \new_[26888]_ ,
    \new_[26889]_ , \new_[26893]_ , \new_[26894]_ , \new_[26898]_ ,
    \new_[26899]_ , \new_[26900]_ , \new_[26904]_ , \new_[26905]_ ,
    \new_[26909]_ , \new_[26910]_ , \new_[26911]_ , \new_[26915]_ ,
    \new_[26916]_ , \new_[26920]_ , \new_[26921]_ , \new_[26922]_ ,
    \new_[26926]_ , \new_[26927]_ , \new_[26931]_ , \new_[26932]_ ,
    \new_[26933]_ , \new_[26937]_ , \new_[26938]_ , \new_[26942]_ ,
    \new_[26943]_ , \new_[26944]_ , \new_[26948]_ , \new_[26949]_ ,
    \new_[26953]_ , \new_[26954]_ , \new_[26955]_ , \new_[26959]_ ,
    \new_[26960]_ , \new_[26964]_ , \new_[26965]_ , \new_[26966]_ ,
    \new_[26970]_ , \new_[26971]_ , \new_[26975]_ , \new_[26976]_ ,
    \new_[26977]_ , \new_[26981]_ , \new_[26982]_ , \new_[26986]_ ,
    \new_[26987]_ , \new_[26988]_ , \new_[26992]_ , \new_[26993]_ ,
    \new_[26997]_ , \new_[26998]_ , \new_[26999]_ , \new_[27003]_ ,
    \new_[27004]_ , \new_[27008]_ , \new_[27009]_ , \new_[27010]_ ,
    \new_[27014]_ , \new_[27015]_ , \new_[27019]_ , \new_[27020]_ ,
    \new_[27021]_ , \new_[27025]_ , \new_[27026]_ , \new_[27030]_ ,
    \new_[27031]_ , \new_[27032]_ , \new_[27036]_ , \new_[27037]_ ,
    \new_[27041]_ , \new_[27042]_ , \new_[27043]_ , \new_[27047]_ ,
    \new_[27048]_ , \new_[27052]_ , \new_[27053]_ , \new_[27054]_ ,
    \new_[27058]_ , \new_[27059]_ , \new_[27063]_ , \new_[27064]_ ,
    \new_[27065]_ , \new_[27069]_ , \new_[27070]_ , \new_[27074]_ ,
    \new_[27075]_ , \new_[27076]_ , \new_[27080]_ , \new_[27081]_ ,
    \new_[27085]_ , \new_[27086]_ , \new_[27087]_ , \new_[27091]_ ,
    \new_[27092]_ , \new_[27096]_ , \new_[27097]_ , \new_[27098]_ ,
    \new_[27102]_ , \new_[27103]_ , \new_[27107]_ , \new_[27108]_ ,
    \new_[27109]_ , \new_[27113]_ , \new_[27114]_ , \new_[27118]_ ,
    \new_[27119]_ , \new_[27120]_ , \new_[27124]_ , \new_[27125]_ ,
    \new_[27129]_ , \new_[27130]_ , \new_[27131]_ , \new_[27135]_ ,
    \new_[27136]_ , \new_[27140]_ , \new_[27141]_ , \new_[27142]_ ,
    \new_[27146]_ , \new_[27147]_ , \new_[27151]_ , \new_[27152]_ ,
    \new_[27153]_ , \new_[27157]_ , \new_[27158]_ , \new_[27162]_ ,
    \new_[27163]_ , \new_[27164]_ , \new_[27168]_ , \new_[27169]_ ,
    \new_[27173]_ , \new_[27174]_ , \new_[27175]_ , \new_[27179]_ ,
    \new_[27180]_ , \new_[27184]_ , \new_[27185]_ , \new_[27186]_ ,
    \new_[27190]_ , \new_[27191]_ , \new_[27195]_ , \new_[27196]_ ,
    \new_[27197]_ , \new_[27201]_ , \new_[27202]_ , \new_[27206]_ ,
    \new_[27207]_ , \new_[27208]_ , \new_[27212]_ , \new_[27213]_ ,
    \new_[27217]_ , \new_[27218]_ , \new_[27219]_ , \new_[27223]_ ,
    \new_[27224]_ , \new_[27228]_ , \new_[27229]_ , \new_[27230]_ ,
    \new_[27234]_ , \new_[27235]_ , \new_[27239]_ , \new_[27240]_ ,
    \new_[27241]_ , \new_[27245]_ , \new_[27246]_ , \new_[27250]_ ,
    \new_[27251]_ , \new_[27252]_ , \new_[27256]_ , \new_[27257]_ ,
    \new_[27261]_ , \new_[27262]_ , \new_[27263]_ , \new_[27267]_ ,
    \new_[27268]_ , \new_[27272]_ , \new_[27273]_ , \new_[27274]_ ,
    \new_[27278]_ , \new_[27279]_ , \new_[27283]_ , \new_[27284]_ ,
    \new_[27285]_ , \new_[27289]_ , \new_[27290]_ , \new_[27294]_ ,
    \new_[27295]_ , \new_[27296]_ , \new_[27300]_ , \new_[27301]_ ,
    \new_[27305]_ , \new_[27306]_ , \new_[27307]_ , \new_[27311]_ ,
    \new_[27312]_ , \new_[27316]_ , \new_[27317]_ , \new_[27318]_ ,
    \new_[27322]_ , \new_[27323]_ , \new_[27327]_ , \new_[27328]_ ,
    \new_[27329]_ , \new_[27333]_ , \new_[27334]_ , \new_[27338]_ ,
    \new_[27339]_ , \new_[27340]_ , \new_[27344]_ , \new_[27345]_ ,
    \new_[27349]_ , \new_[27350]_ , \new_[27351]_ , \new_[27355]_ ,
    \new_[27356]_ , \new_[27360]_ , \new_[27361]_ , \new_[27362]_ ,
    \new_[27366]_ , \new_[27367]_ , \new_[27371]_ , \new_[27372]_ ,
    \new_[27373]_ , \new_[27377]_ , \new_[27378]_ , \new_[27382]_ ,
    \new_[27383]_ , \new_[27384]_ , \new_[27388]_ , \new_[27389]_ ,
    \new_[27393]_ , \new_[27394]_ , \new_[27395]_ , \new_[27399]_ ,
    \new_[27400]_ , \new_[27404]_ , \new_[27405]_ , \new_[27406]_ ,
    \new_[27410]_ , \new_[27411]_ , \new_[27415]_ , \new_[27416]_ ,
    \new_[27417]_ , \new_[27421]_ , \new_[27422]_ , \new_[27426]_ ,
    \new_[27427]_ , \new_[27428]_ , \new_[27432]_ , \new_[27433]_ ,
    \new_[27437]_ , \new_[27438]_ , \new_[27439]_ , \new_[27443]_ ,
    \new_[27444]_ , \new_[27448]_ , \new_[27449]_ , \new_[27450]_ ,
    \new_[27454]_ , \new_[27455]_ , \new_[27459]_ , \new_[27460]_ ,
    \new_[27461]_ , \new_[27465]_ , \new_[27466]_ , \new_[27470]_ ,
    \new_[27471]_ , \new_[27472]_ , \new_[27476]_ , \new_[27477]_ ,
    \new_[27481]_ , \new_[27482]_ , \new_[27483]_ , \new_[27487]_ ,
    \new_[27488]_ , \new_[27492]_ , \new_[27493]_ , \new_[27494]_ ,
    \new_[27498]_ , \new_[27499]_ , \new_[27503]_ , \new_[27504]_ ,
    \new_[27505]_ , \new_[27509]_ , \new_[27510]_ , \new_[27514]_ ,
    \new_[27515]_ , \new_[27516]_ , \new_[27520]_ , \new_[27521]_ ,
    \new_[27525]_ , \new_[27526]_ , \new_[27527]_ , \new_[27531]_ ,
    \new_[27532]_ , \new_[27536]_ , \new_[27537]_ , \new_[27538]_ ,
    \new_[27542]_ , \new_[27543]_ , \new_[27547]_ , \new_[27548]_ ,
    \new_[27549]_ , \new_[27553]_ , \new_[27554]_ , \new_[27558]_ ,
    \new_[27559]_ , \new_[27560]_ , \new_[27564]_ , \new_[27565]_ ,
    \new_[27569]_ , \new_[27570]_ , \new_[27571]_ , \new_[27575]_ ,
    \new_[27576]_ , \new_[27580]_ , \new_[27581]_ , \new_[27582]_ ,
    \new_[27586]_ , \new_[27587]_ , \new_[27591]_ , \new_[27592]_ ,
    \new_[27593]_ , \new_[27597]_ , \new_[27598]_ , \new_[27602]_ ,
    \new_[27603]_ , \new_[27604]_ , \new_[27608]_ , \new_[27609]_ ,
    \new_[27613]_ , \new_[27614]_ , \new_[27615]_ , \new_[27619]_ ,
    \new_[27620]_ , \new_[27624]_ , \new_[27625]_ , \new_[27626]_ ,
    \new_[27630]_ , \new_[27631]_ , \new_[27635]_ , \new_[27636]_ ,
    \new_[27637]_ , \new_[27641]_ , \new_[27642]_ , \new_[27646]_ ,
    \new_[27647]_ , \new_[27648]_ , \new_[27652]_ , \new_[27653]_ ,
    \new_[27657]_ , \new_[27658]_ , \new_[27659]_ , \new_[27663]_ ,
    \new_[27664]_ , \new_[27668]_ , \new_[27669]_ , \new_[27670]_ ,
    \new_[27674]_ , \new_[27675]_ , \new_[27679]_ , \new_[27680]_ ,
    \new_[27681]_ , \new_[27685]_ , \new_[27686]_ , \new_[27690]_ ,
    \new_[27691]_ , \new_[27692]_ , \new_[27696]_ , \new_[27697]_ ,
    \new_[27701]_ , \new_[27702]_ , \new_[27703]_ , \new_[27707]_ ,
    \new_[27708]_ , \new_[27712]_ , \new_[27713]_ , \new_[27714]_ ,
    \new_[27718]_ , \new_[27719]_ , \new_[27723]_ , \new_[27724]_ ,
    \new_[27725]_ , \new_[27729]_ , \new_[27730]_ , \new_[27734]_ ,
    \new_[27735]_ , \new_[27736]_ , \new_[27740]_ , \new_[27741]_ ,
    \new_[27745]_ , \new_[27746]_ , \new_[27747]_ , \new_[27751]_ ,
    \new_[27752]_ , \new_[27756]_ , \new_[27757]_ , \new_[27758]_ ,
    \new_[27762]_ , \new_[27763]_ , \new_[27767]_ , \new_[27768]_ ,
    \new_[27769]_ , \new_[27773]_ , \new_[27774]_ , \new_[27778]_ ,
    \new_[27779]_ , \new_[27780]_ , \new_[27784]_ , \new_[27785]_ ,
    \new_[27789]_ , \new_[27790]_ , \new_[27791]_ , \new_[27795]_ ,
    \new_[27796]_ , \new_[27800]_ , \new_[27801]_ , \new_[27802]_ ,
    \new_[27806]_ , \new_[27807]_ , \new_[27811]_ , \new_[27812]_ ,
    \new_[27813]_ , \new_[27817]_ , \new_[27818]_ , \new_[27822]_ ,
    \new_[27823]_ , \new_[27824]_ , \new_[27828]_ , \new_[27829]_ ,
    \new_[27833]_ , \new_[27834]_ , \new_[27835]_ , \new_[27839]_ ,
    \new_[27840]_ , \new_[27844]_ , \new_[27845]_ , \new_[27846]_ ,
    \new_[27850]_ , \new_[27851]_ , \new_[27855]_ , \new_[27856]_ ,
    \new_[27857]_ , \new_[27861]_ , \new_[27862]_ , \new_[27866]_ ,
    \new_[27867]_ , \new_[27868]_ , \new_[27872]_ , \new_[27873]_ ,
    \new_[27877]_ , \new_[27878]_ , \new_[27879]_ , \new_[27883]_ ,
    \new_[27884]_ , \new_[27888]_ , \new_[27889]_ , \new_[27890]_ ,
    \new_[27894]_ , \new_[27895]_ , \new_[27899]_ , \new_[27900]_ ,
    \new_[27901]_ , \new_[27905]_ , \new_[27906]_ , \new_[27910]_ ,
    \new_[27911]_ , \new_[27912]_ , \new_[27916]_ , \new_[27917]_ ,
    \new_[27921]_ , \new_[27922]_ , \new_[27923]_ , \new_[27927]_ ,
    \new_[27928]_ , \new_[27932]_ , \new_[27933]_ , \new_[27934]_ ,
    \new_[27938]_ , \new_[27939]_ , \new_[27943]_ , \new_[27944]_ ,
    \new_[27945]_ , \new_[27949]_ , \new_[27950]_ , \new_[27954]_ ,
    \new_[27955]_ , \new_[27956]_ , \new_[27960]_ , \new_[27961]_ ,
    \new_[27965]_ , \new_[27966]_ , \new_[27967]_ , \new_[27971]_ ,
    \new_[27972]_ , \new_[27976]_ , \new_[27977]_ , \new_[27978]_ ,
    \new_[27982]_ , \new_[27983]_ , \new_[27987]_ , \new_[27988]_ ,
    \new_[27989]_ , \new_[27993]_ , \new_[27994]_ , \new_[27998]_ ,
    \new_[27999]_ , \new_[28000]_ , \new_[28004]_ , \new_[28005]_ ,
    \new_[28009]_ , \new_[28010]_ , \new_[28011]_ , \new_[28015]_ ,
    \new_[28016]_ , \new_[28020]_ , \new_[28021]_ , \new_[28022]_ ,
    \new_[28026]_ , \new_[28027]_ , \new_[28031]_ , \new_[28032]_ ,
    \new_[28033]_ , \new_[28037]_ , \new_[28038]_ , \new_[28042]_ ,
    \new_[28043]_ , \new_[28044]_ , \new_[28048]_ , \new_[28049]_ ,
    \new_[28053]_ , \new_[28054]_ , \new_[28055]_ , \new_[28059]_ ,
    \new_[28060]_ , \new_[28064]_ , \new_[28065]_ , \new_[28066]_ ,
    \new_[28070]_ , \new_[28071]_ , \new_[28075]_ , \new_[28076]_ ,
    \new_[28077]_ , \new_[28081]_ , \new_[28082]_ , \new_[28086]_ ,
    \new_[28087]_ , \new_[28088]_ , \new_[28092]_ , \new_[28093]_ ,
    \new_[28097]_ , \new_[28098]_ , \new_[28099]_ , \new_[28103]_ ,
    \new_[28104]_ , \new_[28108]_ , \new_[28109]_ , \new_[28110]_ ,
    \new_[28114]_ , \new_[28115]_ , \new_[28119]_ , \new_[28120]_ ,
    \new_[28121]_ , \new_[28125]_ , \new_[28126]_ , \new_[28130]_ ,
    \new_[28131]_ , \new_[28132]_ , \new_[28136]_ , \new_[28137]_ ,
    \new_[28141]_ , \new_[28142]_ , \new_[28143]_ , \new_[28147]_ ,
    \new_[28148]_ , \new_[28152]_ , \new_[28153]_ , \new_[28154]_ ,
    \new_[28158]_ , \new_[28159]_ , \new_[28163]_ , \new_[28164]_ ,
    \new_[28165]_ , \new_[28169]_ , \new_[28170]_ , \new_[28174]_ ,
    \new_[28175]_ , \new_[28176]_ , \new_[28180]_ , \new_[28181]_ ,
    \new_[28185]_ , \new_[28186]_ , \new_[28187]_ , \new_[28191]_ ,
    \new_[28192]_ , \new_[28196]_ , \new_[28197]_ , \new_[28198]_ ,
    \new_[28202]_ , \new_[28203]_ , \new_[28207]_ , \new_[28208]_ ,
    \new_[28209]_ , \new_[28213]_ , \new_[28214]_ , \new_[28218]_ ,
    \new_[28219]_ , \new_[28220]_ , \new_[28224]_ , \new_[28225]_ ,
    \new_[28229]_ , \new_[28230]_ , \new_[28231]_ , \new_[28235]_ ,
    \new_[28236]_ , \new_[28240]_ , \new_[28241]_ , \new_[28242]_ ,
    \new_[28246]_ , \new_[28247]_ , \new_[28251]_ , \new_[28252]_ ,
    \new_[28253]_ , \new_[28257]_ , \new_[28258]_ , \new_[28262]_ ,
    \new_[28263]_ , \new_[28264]_ , \new_[28268]_ , \new_[28269]_ ,
    \new_[28273]_ , \new_[28274]_ , \new_[28275]_ , \new_[28279]_ ,
    \new_[28280]_ , \new_[28284]_ , \new_[28285]_ , \new_[28286]_ ,
    \new_[28290]_ , \new_[28291]_ , \new_[28295]_ , \new_[28296]_ ,
    \new_[28297]_ , \new_[28301]_ , \new_[28302]_ , \new_[28306]_ ,
    \new_[28307]_ , \new_[28308]_ , \new_[28312]_ , \new_[28313]_ ,
    \new_[28317]_ , \new_[28318]_ , \new_[28319]_ , \new_[28323]_ ,
    \new_[28324]_ , \new_[28328]_ , \new_[28329]_ , \new_[28330]_ ,
    \new_[28334]_ , \new_[28335]_ , \new_[28339]_ , \new_[28340]_ ,
    \new_[28341]_ , \new_[28345]_ , \new_[28346]_ , \new_[28350]_ ,
    \new_[28351]_ , \new_[28352]_ , \new_[28356]_ , \new_[28357]_ ,
    \new_[28361]_ , \new_[28362]_ , \new_[28363]_ , \new_[28367]_ ,
    \new_[28368]_ , \new_[28372]_ , \new_[28373]_ , \new_[28374]_ ,
    \new_[28378]_ , \new_[28379]_ , \new_[28383]_ , \new_[28384]_ ,
    \new_[28385]_ , \new_[28389]_ , \new_[28390]_ , \new_[28394]_ ,
    \new_[28395]_ , \new_[28396]_ , \new_[28400]_ , \new_[28401]_ ,
    \new_[28405]_ , \new_[28406]_ , \new_[28407]_ , \new_[28411]_ ,
    \new_[28412]_ , \new_[28416]_ , \new_[28417]_ , \new_[28418]_ ,
    \new_[28422]_ , \new_[28423]_ , \new_[28427]_ , \new_[28428]_ ,
    \new_[28429]_ , \new_[28433]_ , \new_[28434]_ , \new_[28438]_ ,
    \new_[28439]_ , \new_[28440]_ , \new_[28444]_ , \new_[28445]_ ,
    \new_[28449]_ , \new_[28450]_ , \new_[28451]_ , \new_[28455]_ ,
    \new_[28456]_ , \new_[28460]_ , \new_[28461]_ , \new_[28462]_ ,
    \new_[28466]_ , \new_[28467]_ , \new_[28471]_ , \new_[28472]_ ,
    \new_[28473]_ , \new_[28477]_ , \new_[28478]_ , \new_[28482]_ ,
    \new_[28483]_ , \new_[28484]_ , \new_[28488]_ , \new_[28489]_ ,
    \new_[28493]_ , \new_[28494]_ , \new_[28495]_ , \new_[28499]_ ,
    \new_[28500]_ , \new_[28504]_ , \new_[28505]_ , \new_[28506]_ ,
    \new_[28510]_ , \new_[28511]_ , \new_[28515]_ , \new_[28516]_ ,
    \new_[28517]_ , \new_[28521]_ , \new_[28522]_ , \new_[28526]_ ,
    \new_[28527]_ , \new_[28528]_ , \new_[28532]_ , \new_[28533]_ ,
    \new_[28537]_ , \new_[28538]_ , \new_[28539]_ , \new_[28543]_ ,
    \new_[28544]_ , \new_[28548]_ , \new_[28549]_ , \new_[28550]_ ,
    \new_[28554]_ , \new_[28555]_ , \new_[28559]_ , \new_[28560]_ ,
    \new_[28561]_ , \new_[28565]_ , \new_[28566]_ , \new_[28570]_ ,
    \new_[28571]_ , \new_[28572]_ , \new_[28576]_ , \new_[28577]_ ,
    \new_[28581]_ , \new_[28582]_ , \new_[28583]_ , \new_[28587]_ ,
    \new_[28588]_ , \new_[28592]_ , \new_[28593]_ , \new_[28594]_ ,
    \new_[28598]_ , \new_[28599]_ , \new_[28603]_ , \new_[28604]_ ,
    \new_[28605]_ , \new_[28609]_ , \new_[28610]_ , \new_[28614]_ ,
    \new_[28615]_ , \new_[28616]_ , \new_[28620]_ , \new_[28621]_ ,
    \new_[28625]_ , \new_[28626]_ , \new_[28627]_ , \new_[28631]_ ,
    \new_[28632]_ , \new_[28636]_ , \new_[28637]_ , \new_[28638]_ ,
    \new_[28642]_ , \new_[28643]_ , \new_[28647]_ , \new_[28648]_ ,
    \new_[28649]_ , \new_[28653]_ , \new_[28654]_ , \new_[28658]_ ,
    \new_[28659]_ , \new_[28660]_ , \new_[28664]_ , \new_[28665]_ ,
    \new_[28669]_ , \new_[28670]_ , \new_[28671]_ , \new_[28675]_ ,
    \new_[28676]_ , \new_[28680]_ , \new_[28681]_ , \new_[28682]_ ,
    \new_[28686]_ , \new_[28687]_ , \new_[28691]_ , \new_[28692]_ ,
    \new_[28693]_ , \new_[28697]_ , \new_[28698]_ , \new_[28702]_ ,
    \new_[28703]_ , \new_[28704]_ , \new_[28708]_ , \new_[28709]_ ,
    \new_[28713]_ , \new_[28714]_ , \new_[28715]_ , \new_[28719]_ ,
    \new_[28720]_ , \new_[28724]_ , \new_[28725]_ , \new_[28726]_ ,
    \new_[28730]_ , \new_[28731]_ , \new_[28735]_ , \new_[28736]_ ,
    \new_[28737]_ , \new_[28741]_ , \new_[28742]_ , \new_[28746]_ ,
    \new_[28747]_ , \new_[28748]_ , \new_[28752]_ , \new_[28753]_ ,
    \new_[28757]_ , \new_[28758]_ , \new_[28759]_ , \new_[28763]_ ,
    \new_[28764]_ , \new_[28768]_ , \new_[28769]_ , \new_[28770]_ ,
    \new_[28774]_ , \new_[28775]_ , \new_[28779]_ , \new_[28780]_ ,
    \new_[28781]_ , \new_[28785]_ , \new_[28786]_ , \new_[28790]_ ,
    \new_[28791]_ , \new_[28792]_ , \new_[28796]_ , \new_[28797]_ ,
    \new_[28801]_ , \new_[28802]_ , \new_[28803]_ , \new_[28807]_ ,
    \new_[28808]_ , \new_[28812]_ , \new_[28813]_ , \new_[28814]_ ,
    \new_[28818]_ , \new_[28819]_ , \new_[28823]_ , \new_[28824]_ ,
    \new_[28825]_ , \new_[28829]_ , \new_[28830]_ , \new_[28834]_ ,
    \new_[28835]_ , \new_[28836]_ , \new_[28840]_ , \new_[28841]_ ,
    \new_[28845]_ , \new_[28846]_ , \new_[28847]_ , \new_[28851]_ ,
    \new_[28852]_ , \new_[28856]_ , \new_[28857]_ , \new_[28858]_ ,
    \new_[28862]_ , \new_[28863]_ , \new_[28867]_ , \new_[28868]_ ,
    \new_[28869]_ , \new_[28873]_ , \new_[28874]_ , \new_[28878]_ ,
    \new_[28879]_ , \new_[28880]_ , \new_[28884]_ , \new_[28885]_ ,
    \new_[28889]_ , \new_[28890]_ , \new_[28891]_ , \new_[28895]_ ,
    \new_[28896]_ , \new_[28900]_ , \new_[28901]_ , \new_[28902]_ ,
    \new_[28906]_ , \new_[28907]_ , \new_[28911]_ , \new_[28912]_ ,
    \new_[28913]_ , \new_[28917]_ , \new_[28918]_ , \new_[28922]_ ,
    \new_[28923]_ , \new_[28924]_ , \new_[28928]_ , \new_[28929]_ ,
    \new_[28933]_ , \new_[28934]_ , \new_[28935]_ , \new_[28939]_ ,
    \new_[28940]_ , \new_[28944]_ , \new_[28945]_ , \new_[28946]_ ,
    \new_[28950]_ , \new_[28951]_ , \new_[28955]_ , \new_[28956]_ ,
    \new_[28957]_ , \new_[28961]_ , \new_[28962]_ , \new_[28966]_ ,
    \new_[28967]_ , \new_[28968]_ , \new_[28972]_ , \new_[28973]_ ,
    \new_[28977]_ , \new_[28978]_ , \new_[28979]_ , \new_[28983]_ ,
    \new_[28984]_ , \new_[28988]_ , \new_[28989]_ , \new_[28990]_ ,
    \new_[28994]_ , \new_[28995]_ , \new_[28999]_ , \new_[29000]_ ,
    \new_[29001]_ , \new_[29005]_ , \new_[29006]_ , \new_[29010]_ ,
    \new_[29011]_ , \new_[29012]_ , \new_[29016]_ , \new_[29017]_ ,
    \new_[29021]_ , \new_[29022]_ , \new_[29023]_ , \new_[29027]_ ,
    \new_[29028]_ , \new_[29032]_ , \new_[29033]_ , \new_[29034]_ ,
    \new_[29038]_ , \new_[29039]_ , \new_[29043]_ , \new_[29044]_ ,
    \new_[29045]_ , \new_[29049]_ , \new_[29050]_ , \new_[29054]_ ,
    \new_[29055]_ , \new_[29056]_ , \new_[29060]_ , \new_[29061]_ ,
    \new_[29065]_ , \new_[29066]_ , \new_[29067]_ , \new_[29071]_ ,
    \new_[29072]_ , \new_[29076]_ , \new_[29077]_ , \new_[29078]_ ,
    \new_[29082]_ , \new_[29083]_ , \new_[29087]_ , \new_[29088]_ ,
    \new_[29089]_ , \new_[29093]_ , \new_[29094]_ , \new_[29098]_ ,
    \new_[29099]_ , \new_[29100]_ , \new_[29104]_ , \new_[29105]_ ,
    \new_[29109]_ , \new_[29110]_ , \new_[29111]_ , \new_[29115]_ ,
    \new_[29116]_ , \new_[29120]_ , \new_[29121]_ , \new_[29122]_ ,
    \new_[29126]_ , \new_[29127]_ , \new_[29131]_ , \new_[29132]_ ,
    \new_[29133]_ , \new_[29137]_ , \new_[29138]_ , \new_[29142]_ ,
    \new_[29143]_ , \new_[29144]_ , \new_[29148]_ , \new_[29149]_ ,
    \new_[29153]_ , \new_[29154]_ , \new_[29155]_ , \new_[29159]_ ,
    \new_[29160]_ , \new_[29164]_ , \new_[29165]_ , \new_[29166]_ ,
    \new_[29170]_ , \new_[29171]_ , \new_[29175]_ , \new_[29176]_ ,
    \new_[29177]_ , \new_[29181]_ , \new_[29182]_ , \new_[29186]_ ,
    \new_[29187]_ , \new_[29188]_ , \new_[29192]_ , \new_[29193]_ ,
    \new_[29197]_ , \new_[29198]_ , \new_[29199]_ , \new_[29203]_ ,
    \new_[29204]_ , \new_[29208]_ , \new_[29209]_ , \new_[29210]_ ,
    \new_[29214]_ , \new_[29215]_ , \new_[29219]_ , \new_[29220]_ ,
    \new_[29221]_ , \new_[29225]_ , \new_[29226]_ , \new_[29230]_ ,
    \new_[29231]_ , \new_[29232]_ , \new_[29236]_ , \new_[29237]_ ,
    \new_[29241]_ , \new_[29242]_ , \new_[29243]_ , \new_[29247]_ ,
    \new_[29248]_ , \new_[29252]_ , \new_[29253]_ , \new_[29254]_ ,
    \new_[29258]_ , \new_[29259]_ , \new_[29263]_ , \new_[29264]_ ,
    \new_[29265]_ , \new_[29269]_ , \new_[29270]_ , \new_[29274]_ ,
    \new_[29275]_ , \new_[29276]_ , \new_[29280]_ , \new_[29281]_ ,
    \new_[29285]_ , \new_[29286]_ , \new_[29287]_ , \new_[29291]_ ,
    \new_[29292]_ , \new_[29296]_ , \new_[29297]_ , \new_[29298]_ ,
    \new_[29302]_ , \new_[29303]_ , \new_[29307]_ , \new_[29308]_ ,
    \new_[29309]_ , \new_[29313]_ , \new_[29314]_ , \new_[29318]_ ,
    \new_[29319]_ , \new_[29320]_ , \new_[29324]_ , \new_[29325]_ ,
    \new_[29329]_ , \new_[29330]_ , \new_[29331]_ , \new_[29335]_ ,
    \new_[29336]_ , \new_[29340]_ , \new_[29341]_ , \new_[29342]_ ,
    \new_[29346]_ , \new_[29347]_ , \new_[29351]_ , \new_[29352]_ ,
    \new_[29353]_ , \new_[29357]_ , \new_[29358]_ , \new_[29362]_ ,
    \new_[29363]_ , \new_[29364]_ , \new_[29368]_ , \new_[29369]_ ,
    \new_[29373]_ , \new_[29374]_ , \new_[29375]_ , \new_[29379]_ ,
    \new_[29380]_ , \new_[29384]_ , \new_[29385]_ , \new_[29386]_ ,
    \new_[29390]_ , \new_[29391]_ , \new_[29395]_ , \new_[29396]_ ,
    \new_[29397]_ , \new_[29401]_ , \new_[29402]_ , \new_[29406]_ ,
    \new_[29407]_ , \new_[29408]_ , \new_[29412]_ , \new_[29413]_ ,
    \new_[29417]_ , \new_[29418]_ , \new_[29419]_ , \new_[29423]_ ,
    \new_[29424]_ , \new_[29428]_ , \new_[29429]_ , \new_[29430]_ ,
    \new_[29434]_ , \new_[29435]_ , \new_[29439]_ , \new_[29440]_ ,
    \new_[29441]_ , \new_[29445]_ , \new_[29446]_ , \new_[29450]_ ,
    \new_[29451]_ , \new_[29452]_ , \new_[29456]_ , \new_[29457]_ ,
    \new_[29461]_ , \new_[29462]_ , \new_[29463]_ , \new_[29467]_ ,
    \new_[29468]_ , \new_[29472]_ , \new_[29473]_ , \new_[29474]_ ,
    \new_[29478]_ , \new_[29479]_ , \new_[29483]_ , \new_[29484]_ ,
    \new_[29485]_ , \new_[29489]_ , \new_[29490]_ , \new_[29494]_ ,
    \new_[29495]_ , \new_[29496]_ , \new_[29500]_ , \new_[29501]_ ,
    \new_[29505]_ , \new_[29506]_ , \new_[29507]_ , \new_[29511]_ ,
    \new_[29512]_ , \new_[29516]_ , \new_[29517]_ , \new_[29518]_ ,
    \new_[29522]_ , \new_[29523]_ , \new_[29527]_ , \new_[29528]_ ,
    \new_[29529]_ , \new_[29533]_ , \new_[29534]_ , \new_[29538]_ ,
    \new_[29539]_ , \new_[29540]_ , \new_[29544]_ , \new_[29545]_ ,
    \new_[29549]_ , \new_[29550]_ , \new_[29551]_ , \new_[29555]_ ,
    \new_[29556]_ , \new_[29560]_ , \new_[29561]_ , \new_[29562]_ ,
    \new_[29566]_ , \new_[29567]_ , \new_[29571]_ , \new_[29572]_ ,
    \new_[29573]_ , \new_[29577]_ , \new_[29578]_ , \new_[29582]_ ,
    \new_[29583]_ , \new_[29584]_ , \new_[29588]_ , \new_[29589]_ ,
    \new_[29593]_ , \new_[29594]_ , \new_[29595]_ , \new_[29599]_ ,
    \new_[29600]_ , \new_[29604]_ , \new_[29605]_ , \new_[29606]_ ,
    \new_[29610]_ , \new_[29611]_ , \new_[29615]_ , \new_[29616]_ ,
    \new_[29617]_ , \new_[29621]_ , \new_[29622]_ , \new_[29626]_ ,
    \new_[29627]_ , \new_[29628]_ , \new_[29632]_ , \new_[29633]_ ,
    \new_[29637]_ , \new_[29638]_ , \new_[29639]_ , \new_[29643]_ ,
    \new_[29644]_ , \new_[29648]_ , \new_[29649]_ , \new_[29650]_ ,
    \new_[29654]_ , \new_[29655]_ , \new_[29659]_ , \new_[29660]_ ,
    \new_[29661]_ , \new_[29665]_ , \new_[29666]_ , \new_[29670]_ ,
    \new_[29671]_ , \new_[29672]_ , \new_[29676]_ , \new_[29677]_ ,
    \new_[29681]_ , \new_[29682]_ , \new_[29683]_ , \new_[29687]_ ,
    \new_[29688]_ , \new_[29692]_ , \new_[29693]_ , \new_[29694]_ ,
    \new_[29698]_ , \new_[29699]_ , \new_[29703]_ , \new_[29704]_ ,
    \new_[29705]_ , \new_[29709]_ , \new_[29710]_ , \new_[29714]_ ,
    \new_[29715]_ , \new_[29716]_ , \new_[29720]_ , \new_[29721]_ ,
    \new_[29725]_ , \new_[29726]_ , \new_[29727]_ , \new_[29731]_ ,
    \new_[29732]_ , \new_[29736]_ , \new_[29737]_ , \new_[29738]_ ,
    \new_[29742]_ , \new_[29743]_ , \new_[29747]_ , \new_[29748]_ ,
    \new_[29749]_ , \new_[29753]_ , \new_[29754]_ , \new_[29758]_ ,
    \new_[29759]_ , \new_[29760]_ , \new_[29764]_ , \new_[29765]_ ,
    \new_[29769]_ , \new_[29770]_ , \new_[29771]_ , \new_[29775]_ ,
    \new_[29776]_ , \new_[29780]_ , \new_[29781]_ , \new_[29782]_ ,
    \new_[29786]_ , \new_[29787]_ , \new_[29791]_ , \new_[29792]_ ,
    \new_[29793]_ , \new_[29797]_ , \new_[29798]_ , \new_[29802]_ ,
    \new_[29803]_ , \new_[29804]_ , \new_[29808]_ , \new_[29809]_ ,
    \new_[29813]_ , \new_[29814]_ , \new_[29815]_ , \new_[29819]_ ,
    \new_[29820]_ , \new_[29824]_ , \new_[29825]_ , \new_[29826]_ ,
    \new_[29830]_ , \new_[29831]_ , \new_[29835]_ , \new_[29836]_ ,
    \new_[29837]_ , \new_[29841]_ , \new_[29842]_ , \new_[29846]_ ,
    \new_[29847]_ , \new_[29848]_ , \new_[29852]_ , \new_[29853]_ ,
    \new_[29857]_ , \new_[29858]_ , \new_[29859]_ , \new_[29863]_ ,
    \new_[29864]_ , \new_[29868]_ , \new_[29869]_ , \new_[29870]_ ,
    \new_[29874]_ , \new_[29875]_ , \new_[29879]_ , \new_[29880]_ ,
    \new_[29881]_ , \new_[29885]_ , \new_[29886]_ , \new_[29890]_ ,
    \new_[29891]_ , \new_[29892]_ , \new_[29896]_ , \new_[29897]_ ,
    \new_[29901]_ , \new_[29902]_ , \new_[29903]_ , \new_[29907]_ ,
    \new_[29908]_ , \new_[29912]_ , \new_[29913]_ , \new_[29914]_ ,
    \new_[29918]_ , \new_[29919]_ , \new_[29923]_ , \new_[29924]_ ,
    \new_[29925]_ , \new_[29929]_ , \new_[29930]_ , \new_[29934]_ ,
    \new_[29935]_ , \new_[29936]_ , \new_[29940]_ , \new_[29941]_ ,
    \new_[29945]_ , \new_[29946]_ , \new_[29947]_ , \new_[29951]_ ,
    \new_[29952]_ , \new_[29956]_ , \new_[29957]_ , \new_[29958]_ ,
    \new_[29962]_ , \new_[29963]_ , \new_[29967]_ , \new_[29968]_ ,
    \new_[29969]_ , \new_[29973]_ , \new_[29974]_ , \new_[29978]_ ,
    \new_[29979]_ , \new_[29980]_ , \new_[29984]_ , \new_[29985]_ ,
    \new_[29989]_ , \new_[29990]_ , \new_[29991]_ , \new_[29995]_ ,
    \new_[29996]_ , \new_[30000]_ , \new_[30001]_ , \new_[30002]_ ,
    \new_[30006]_ , \new_[30007]_ , \new_[30011]_ , \new_[30012]_ ,
    \new_[30013]_ , \new_[30017]_ , \new_[30018]_ , \new_[30022]_ ,
    \new_[30023]_ , \new_[30024]_ , \new_[30028]_ , \new_[30029]_ ,
    \new_[30033]_ , \new_[30034]_ , \new_[30035]_ , \new_[30039]_ ,
    \new_[30040]_ , \new_[30044]_ , \new_[30045]_ , \new_[30046]_ ,
    \new_[30050]_ , \new_[30051]_ , \new_[30055]_ , \new_[30056]_ ,
    \new_[30057]_ , \new_[30061]_ , \new_[30062]_ , \new_[30066]_ ,
    \new_[30067]_ , \new_[30068]_ , \new_[30072]_ , \new_[30073]_ ,
    \new_[30077]_ , \new_[30078]_ , \new_[30079]_ , \new_[30083]_ ,
    \new_[30084]_ , \new_[30088]_ , \new_[30089]_ , \new_[30090]_ ,
    \new_[30094]_ , \new_[30095]_ , \new_[30099]_ , \new_[30100]_ ,
    \new_[30101]_ , \new_[30105]_ , \new_[30106]_ , \new_[30110]_ ,
    \new_[30111]_ , \new_[30112]_ , \new_[30116]_ , \new_[30117]_ ,
    \new_[30121]_ , \new_[30122]_ , \new_[30123]_ , \new_[30127]_ ,
    \new_[30128]_ , \new_[30132]_ , \new_[30133]_ , \new_[30134]_ ,
    \new_[30138]_ , \new_[30139]_ , \new_[30143]_ , \new_[30144]_ ,
    \new_[30145]_ , \new_[30149]_ , \new_[30150]_ , \new_[30154]_ ,
    \new_[30155]_ , \new_[30156]_ , \new_[30160]_ , \new_[30161]_ ,
    \new_[30165]_ , \new_[30166]_ , \new_[30167]_ , \new_[30171]_ ,
    \new_[30172]_ , \new_[30176]_ , \new_[30177]_ , \new_[30178]_ ,
    \new_[30182]_ , \new_[30183]_ , \new_[30187]_ , \new_[30188]_ ,
    \new_[30189]_ , \new_[30193]_ , \new_[30194]_ , \new_[30198]_ ,
    \new_[30199]_ , \new_[30200]_ , \new_[30204]_ , \new_[30205]_ ,
    \new_[30209]_ , \new_[30210]_ , \new_[30211]_ , \new_[30215]_ ,
    \new_[30216]_ , \new_[30220]_ , \new_[30221]_ , \new_[30222]_ ,
    \new_[30226]_ , \new_[30227]_ , \new_[30231]_ , \new_[30232]_ ,
    \new_[30233]_ , \new_[30237]_ , \new_[30238]_ , \new_[30242]_ ,
    \new_[30243]_ , \new_[30244]_ , \new_[30248]_ , \new_[30249]_ ,
    \new_[30253]_ , \new_[30254]_ , \new_[30255]_ , \new_[30259]_ ,
    \new_[30260]_ , \new_[30264]_ , \new_[30265]_ , \new_[30266]_ ,
    \new_[30270]_ , \new_[30271]_ , \new_[30275]_ , \new_[30276]_ ,
    \new_[30277]_ , \new_[30281]_ , \new_[30282]_ , \new_[30286]_ ,
    \new_[30287]_ , \new_[30288]_ , \new_[30292]_ , \new_[30293]_ ,
    \new_[30297]_ , \new_[30298]_ , \new_[30299]_ , \new_[30303]_ ,
    \new_[30304]_ , \new_[30308]_ , \new_[30309]_ , \new_[30310]_ ,
    \new_[30314]_ , \new_[30315]_ , \new_[30319]_ , \new_[30320]_ ,
    \new_[30321]_ , \new_[30325]_ , \new_[30326]_ , \new_[30330]_ ,
    \new_[30331]_ , \new_[30332]_ , \new_[30336]_ , \new_[30337]_ ,
    \new_[30341]_ , \new_[30342]_ , \new_[30343]_ , \new_[30347]_ ,
    \new_[30348]_ , \new_[30352]_ , \new_[30353]_ , \new_[30354]_ ,
    \new_[30358]_ , \new_[30359]_ , \new_[30363]_ , \new_[30364]_ ,
    \new_[30365]_ , \new_[30369]_ , \new_[30370]_ , \new_[30374]_ ,
    \new_[30375]_ , \new_[30376]_ , \new_[30380]_ , \new_[30381]_ ,
    \new_[30385]_ , \new_[30386]_ , \new_[30387]_ , \new_[30391]_ ,
    \new_[30392]_ , \new_[30396]_ , \new_[30397]_ , \new_[30398]_ ,
    \new_[30402]_ , \new_[30403]_ , \new_[30407]_ , \new_[30408]_ ,
    \new_[30409]_ , \new_[30413]_ , \new_[30414]_ , \new_[30418]_ ,
    \new_[30419]_ , \new_[30420]_ , \new_[30424]_ , \new_[30425]_ ,
    \new_[30429]_ , \new_[30430]_ , \new_[30431]_ , \new_[30435]_ ,
    \new_[30436]_ , \new_[30440]_ , \new_[30441]_ , \new_[30442]_ ,
    \new_[30446]_ , \new_[30447]_ , \new_[30451]_ , \new_[30452]_ ,
    \new_[30453]_ , \new_[30457]_ , \new_[30458]_ , \new_[30462]_ ,
    \new_[30463]_ , \new_[30464]_ , \new_[30468]_ , \new_[30469]_ ,
    \new_[30473]_ , \new_[30474]_ , \new_[30475]_ , \new_[30479]_ ,
    \new_[30480]_ , \new_[30484]_ , \new_[30485]_ , \new_[30486]_ ,
    \new_[30490]_ , \new_[30491]_ , \new_[30495]_ , \new_[30496]_ ,
    \new_[30497]_ , \new_[30501]_ , \new_[30502]_ , \new_[30506]_ ,
    \new_[30507]_ , \new_[30508]_ , \new_[30512]_ , \new_[30513]_ ,
    \new_[30517]_ , \new_[30518]_ , \new_[30519]_ , \new_[30523]_ ,
    \new_[30524]_ , \new_[30528]_ , \new_[30529]_ , \new_[30530]_ ,
    \new_[30534]_ , \new_[30535]_ , \new_[30539]_ , \new_[30540]_ ,
    \new_[30541]_ , \new_[30545]_ , \new_[30546]_ , \new_[30550]_ ,
    \new_[30551]_ , \new_[30552]_ , \new_[30556]_ , \new_[30557]_ ,
    \new_[30561]_ , \new_[30562]_ , \new_[30563]_ , \new_[30567]_ ,
    \new_[30568]_ , \new_[30572]_ , \new_[30573]_ , \new_[30574]_ ,
    \new_[30578]_ , \new_[30579]_ , \new_[30583]_ , \new_[30584]_ ,
    \new_[30585]_ , \new_[30589]_ , \new_[30590]_ , \new_[30594]_ ,
    \new_[30595]_ , \new_[30596]_ , \new_[30600]_ , \new_[30601]_ ,
    \new_[30605]_ , \new_[30606]_ , \new_[30607]_ , \new_[30611]_ ,
    \new_[30612]_ , \new_[30616]_ , \new_[30617]_ , \new_[30618]_ ,
    \new_[30622]_ , \new_[30623]_ , \new_[30627]_ , \new_[30628]_ ,
    \new_[30629]_ , \new_[30633]_ , \new_[30634]_ , \new_[30638]_ ,
    \new_[30639]_ , \new_[30640]_ , \new_[30644]_ , \new_[30645]_ ,
    \new_[30649]_ , \new_[30650]_ , \new_[30651]_ , \new_[30655]_ ,
    \new_[30656]_ , \new_[30660]_ , \new_[30661]_ , \new_[30662]_ ,
    \new_[30666]_ , \new_[30667]_ , \new_[30671]_ , \new_[30672]_ ,
    \new_[30673]_ , \new_[30677]_ , \new_[30678]_ , \new_[30682]_ ,
    \new_[30683]_ , \new_[30684]_ , \new_[30688]_ , \new_[30689]_ ,
    \new_[30693]_ , \new_[30694]_ , \new_[30695]_ , \new_[30699]_ ,
    \new_[30700]_ , \new_[30704]_ , \new_[30705]_ , \new_[30706]_ ,
    \new_[30710]_ , \new_[30711]_ , \new_[30715]_ , \new_[30716]_ ,
    \new_[30717]_ , \new_[30721]_ , \new_[30722]_ , \new_[30726]_ ,
    \new_[30727]_ , \new_[30728]_ , \new_[30732]_ , \new_[30733]_ ,
    \new_[30737]_ , \new_[30738]_ , \new_[30739]_ , \new_[30743]_ ,
    \new_[30744]_ , \new_[30748]_ , \new_[30749]_ , \new_[30750]_ ,
    \new_[30754]_ , \new_[30755]_ , \new_[30759]_ , \new_[30760]_ ,
    \new_[30761]_ , \new_[30765]_ , \new_[30766]_ , \new_[30770]_ ,
    \new_[30771]_ , \new_[30772]_ , \new_[30776]_ , \new_[30777]_ ,
    \new_[30781]_ , \new_[30782]_ , \new_[30783]_ , \new_[30787]_ ,
    \new_[30788]_ , \new_[30792]_ , \new_[30793]_ , \new_[30794]_ ,
    \new_[30798]_ , \new_[30799]_ , \new_[30803]_ , \new_[30804]_ ,
    \new_[30805]_ , \new_[30809]_ , \new_[30810]_ , \new_[30814]_ ,
    \new_[30815]_ , \new_[30816]_ , \new_[30820]_ , \new_[30821]_ ,
    \new_[30825]_ , \new_[30826]_ , \new_[30827]_ , \new_[30831]_ ,
    \new_[30832]_ , \new_[30836]_ , \new_[30837]_ , \new_[30838]_ ,
    \new_[30842]_ , \new_[30843]_ , \new_[30847]_ , \new_[30848]_ ,
    \new_[30849]_ , \new_[30853]_ , \new_[30854]_ , \new_[30858]_ ,
    \new_[30859]_ , \new_[30860]_ , \new_[30864]_ , \new_[30865]_ ,
    \new_[30869]_ , \new_[30870]_ , \new_[30871]_ , \new_[30875]_ ,
    \new_[30876]_ , \new_[30880]_ , \new_[30881]_ , \new_[30882]_ ,
    \new_[30886]_ , \new_[30887]_ , \new_[30891]_ , \new_[30892]_ ,
    \new_[30893]_ , \new_[30897]_ , \new_[30898]_ , \new_[30902]_ ,
    \new_[30903]_ , \new_[30904]_ , \new_[30908]_ , \new_[30909]_ ,
    \new_[30913]_ , \new_[30914]_ , \new_[30915]_ , \new_[30919]_ ,
    \new_[30920]_ , \new_[30924]_ , \new_[30925]_ , \new_[30926]_ ,
    \new_[30930]_ , \new_[30931]_ , \new_[30935]_ , \new_[30936]_ ,
    \new_[30937]_ , \new_[30941]_ , \new_[30942]_ , \new_[30946]_ ,
    \new_[30947]_ , \new_[30948]_ , \new_[30952]_ , \new_[30953]_ ,
    \new_[30957]_ , \new_[30958]_ , \new_[30959]_ , \new_[30963]_ ,
    \new_[30964]_ , \new_[30968]_ , \new_[30969]_ , \new_[30970]_ ,
    \new_[30974]_ , \new_[30975]_ , \new_[30979]_ , \new_[30980]_ ,
    \new_[30981]_ , \new_[30985]_ , \new_[30986]_ , \new_[30990]_ ,
    \new_[30991]_ , \new_[30992]_ , \new_[30996]_ , \new_[30997]_ ,
    \new_[31001]_ , \new_[31002]_ , \new_[31003]_ , \new_[31007]_ ,
    \new_[31008]_ , \new_[31012]_ , \new_[31013]_ , \new_[31014]_ ,
    \new_[31018]_ , \new_[31019]_ , \new_[31023]_ , \new_[31024]_ ,
    \new_[31025]_ , \new_[31029]_ , \new_[31030]_ , \new_[31034]_ ,
    \new_[31035]_ , \new_[31036]_ , \new_[31040]_ , \new_[31041]_ ,
    \new_[31045]_ , \new_[31046]_ , \new_[31047]_ , \new_[31051]_ ,
    \new_[31052]_ , \new_[31056]_ , \new_[31057]_ , \new_[31058]_ ,
    \new_[31062]_ , \new_[31063]_ , \new_[31067]_ , \new_[31068]_ ,
    \new_[31069]_ , \new_[31073]_ , \new_[31074]_ , \new_[31078]_ ,
    \new_[31079]_ , \new_[31080]_ , \new_[31084]_ , \new_[31085]_ ,
    \new_[31089]_ , \new_[31090]_ , \new_[31091]_ , \new_[31095]_ ,
    \new_[31096]_ , \new_[31100]_ , \new_[31101]_ , \new_[31102]_ ,
    \new_[31106]_ , \new_[31107]_ , \new_[31111]_ , \new_[31112]_ ,
    \new_[31113]_ , \new_[31117]_ , \new_[31118]_ , \new_[31122]_ ,
    \new_[31123]_ , \new_[31124]_ , \new_[31128]_ , \new_[31129]_ ,
    \new_[31133]_ , \new_[31134]_ , \new_[31135]_ , \new_[31139]_ ,
    \new_[31140]_ , \new_[31144]_ , \new_[31145]_ , \new_[31146]_ ,
    \new_[31150]_ , \new_[31151]_ , \new_[31155]_ , \new_[31156]_ ,
    \new_[31157]_ , \new_[31161]_ , \new_[31162]_ , \new_[31166]_ ,
    \new_[31167]_ , \new_[31168]_ , \new_[31172]_ , \new_[31173]_ ,
    \new_[31177]_ , \new_[31178]_ , \new_[31179]_ , \new_[31183]_ ,
    \new_[31184]_ , \new_[31188]_ , \new_[31189]_ , \new_[31190]_ ,
    \new_[31194]_ , \new_[31195]_ , \new_[31199]_ , \new_[31200]_ ,
    \new_[31201]_ , \new_[31205]_ , \new_[31206]_ , \new_[31210]_ ,
    \new_[31211]_ , \new_[31212]_ , \new_[31216]_ , \new_[31217]_ ,
    \new_[31221]_ , \new_[31222]_ , \new_[31223]_ , \new_[31227]_ ,
    \new_[31228]_ , \new_[31232]_ , \new_[31233]_ , \new_[31234]_ ,
    \new_[31238]_ , \new_[31239]_ , \new_[31243]_ , \new_[31244]_ ,
    \new_[31245]_ , \new_[31249]_ , \new_[31250]_ , \new_[31254]_ ,
    \new_[31255]_ , \new_[31256]_ , \new_[31260]_ , \new_[31261]_ ,
    \new_[31265]_ , \new_[31266]_ , \new_[31267]_ , \new_[31271]_ ,
    \new_[31272]_ , \new_[31276]_ , \new_[31277]_ , \new_[31278]_ ,
    \new_[31282]_ , \new_[31283]_ , \new_[31287]_ , \new_[31288]_ ,
    \new_[31289]_ , \new_[31293]_ , \new_[31294]_ , \new_[31298]_ ,
    \new_[31299]_ , \new_[31300]_ , \new_[31304]_ , \new_[31305]_ ,
    \new_[31309]_ , \new_[31310]_ , \new_[31311]_ , \new_[31315]_ ,
    \new_[31316]_ , \new_[31320]_ , \new_[31321]_ , \new_[31322]_ ,
    \new_[31326]_ , \new_[31327]_ , \new_[31331]_ , \new_[31332]_ ,
    \new_[31333]_ , \new_[31337]_ , \new_[31338]_ , \new_[31342]_ ,
    \new_[31343]_ , \new_[31344]_ , \new_[31348]_ , \new_[31349]_ ,
    \new_[31353]_ , \new_[31354]_ , \new_[31355]_ , \new_[31359]_ ,
    \new_[31360]_ , \new_[31364]_ , \new_[31365]_ , \new_[31366]_ ,
    \new_[31370]_ , \new_[31371]_ , \new_[31375]_ , \new_[31376]_ ,
    \new_[31377]_ , \new_[31381]_ , \new_[31382]_ , \new_[31386]_ ,
    \new_[31387]_ , \new_[31388]_ , \new_[31392]_ , \new_[31393]_ ,
    \new_[31397]_ , \new_[31398]_ , \new_[31399]_ , \new_[31403]_ ,
    \new_[31404]_ , \new_[31408]_ , \new_[31409]_ , \new_[31410]_ ,
    \new_[31414]_ , \new_[31415]_ , \new_[31419]_ , \new_[31420]_ ,
    \new_[31421]_ , \new_[31425]_ , \new_[31426]_ , \new_[31430]_ ,
    \new_[31431]_ , \new_[31432]_ , \new_[31436]_ , \new_[31437]_ ,
    \new_[31441]_ , \new_[31442]_ , \new_[31443]_ , \new_[31447]_ ,
    \new_[31448]_ , \new_[31452]_ , \new_[31453]_ , \new_[31454]_ ,
    \new_[31458]_ , \new_[31459]_ , \new_[31463]_ , \new_[31464]_ ,
    \new_[31465]_ , \new_[31469]_ , \new_[31470]_ , \new_[31474]_ ,
    \new_[31475]_ , \new_[31476]_ , \new_[31480]_ , \new_[31481]_ ,
    \new_[31485]_ , \new_[31486]_ , \new_[31487]_ , \new_[31491]_ ,
    \new_[31492]_ , \new_[31496]_ , \new_[31497]_ , \new_[31498]_ ,
    \new_[31502]_ , \new_[31503]_ , \new_[31507]_ , \new_[31508]_ ,
    \new_[31509]_ , \new_[31513]_ , \new_[31514]_ , \new_[31518]_ ,
    \new_[31519]_ , \new_[31520]_ , \new_[31524]_ , \new_[31525]_ ,
    \new_[31529]_ , \new_[31530]_ , \new_[31531]_ , \new_[31535]_ ,
    \new_[31536]_ , \new_[31540]_ , \new_[31541]_ , \new_[31542]_ ,
    \new_[31546]_ , \new_[31547]_ , \new_[31551]_ , \new_[31552]_ ,
    \new_[31553]_ , \new_[31557]_ , \new_[31558]_ , \new_[31562]_ ,
    \new_[31563]_ , \new_[31564]_ , \new_[31568]_ , \new_[31569]_ ,
    \new_[31573]_ , \new_[31574]_ , \new_[31575]_ , \new_[31579]_ ,
    \new_[31580]_ , \new_[31584]_ , \new_[31585]_ , \new_[31586]_ ,
    \new_[31590]_ , \new_[31591]_ , \new_[31595]_ , \new_[31596]_ ,
    \new_[31597]_ , \new_[31601]_ , \new_[31602]_ , \new_[31606]_ ,
    \new_[31607]_ , \new_[31608]_ , \new_[31612]_ , \new_[31613]_ ,
    \new_[31617]_ , \new_[31618]_ , \new_[31619]_ , \new_[31623]_ ,
    \new_[31624]_ , \new_[31628]_ , \new_[31629]_ , \new_[31630]_ ,
    \new_[31634]_ , \new_[31635]_ , \new_[31639]_ , \new_[31640]_ ,
    \new_[31641]_ , \new_[31645]_ , \new_[31646]_ , \new_[31650]_ ,
    \new_[31651]_ , \new_[31652]_ , \new_[31656]_ , \new_[31657]_ ,
    \new_[31661]_ , \new_[31662]_ , \new_[31663]_ , \new_[31667]_ ,
    \new_[31668]_ , \new_[31672]_ , \new_[31673]_ , \new_[31674]_ ,
    \new_[31678]_ , \new_[31679]_ , \new_[31683]_ , \new_[31684]_ ,
    \new_[31685]_ , \new_[31689]_ , \new_[31690]_ , \new_[31694]_ ,
    \new_[31695]_ , \new_[31696]_ , \new_[31700]_ , \new_[31701]_ ,
    \new_[31705]_ , \new_[31706]_ , \new_[31707]_ , \new_[31711]_ ,
    \new_[31712]_ , \new_[31716]_ , \new_[31717]_ , \new_[31718]_ ,
    \new_[31722]_ , \new_[31723]_ , \new_[31727]_ , \new_[31728]_ ,
    \new_[31729]_ , \new_[31733]_ , \new_[31734]_ , \new_[31738]_ ,
    \new_[31739]_ , \new_[31740]_ , \new_[31744]_ , \new_[31745]_ ,
    \new_[31749]_ , \new_[31750]_ , \new_[31751]_ , \new_[31755]_ ,
    \new_[31756]_ , \new_[31760]_ , \new_[31761]_ , \new_[31762]_ ,
    \new_[31766]_ , \new_[31767]_ , \new_[31771]_ , \new_[31772]_ ,
    \new_[31773]_ , \new_[31777]_ , \new_[31778]_ , \new_[31782]_ ,
    \new_[31783]_ , \new_[31784]_ , \new_[31788]_ , \new_[31789]_ ,
    \new_[31793]_ , \new_[31794]_ , \new_[31795]_ , \new_[31799]_ ,
    \new_[31800]_ , \new_[31804]_ , \new_[31805]_ , \new_[31806]_ ,
    \new_[31810]_ , \new_[31811]_ , \new_[31815]_ , \new_[31816]_ ,
    \new_[31817]_ , \new_[31821]_ , \new_[31822]_ , \new_[31826]_ ,
    \new_[31827]_ , \new_[31828]_ , \new_[31832]_ , \new_[31833]_ ,
    \new_[31837]_ , \new_[31838]_ , \new_[31839]_ , \new_[31843]_ ,
    \new_[31844]_ , \new_[31848]_ , \new_[31849]_ , \new_[31850]_ ,
    \new_[31854]_ , \new_[31855]_ , \new_[31859]_ , \new_[31860]_ ,
    \new_[31861]_ , \new_[31865]_ , \new_[31866]_ , \new_[31870]_ ,
    \new_[31871]_ , \new_[31872]_ , \new_[31876]_ , \new_[31877]_ ,
    \new_[31881]_ , \new_[31882]_ , \new_[31883]_ , \new_[31887]_ ,
    \new_[31888]_ , \new_[31892]_ , \new_[31893]_ , \new_[31894]_ ,
    \new_[31898]_ , \new_[31899]_ , \new_[31903]_ , \new_[31904]_ ,
    \new_[31905]_ , \new_[31909]_ , \new_[31910]_ , \new_[31914]_ ,
    \new_[31915]_ , \new_[31916]_ , \new_[31920]_ , \new_[31921]_ ,
    \new_[31925]_ , \new_[31926]_ , \new_[31927]_ , \new_[31931]_ ,
    \new_[31932]_ , \new_[31936]_ , \new_[31937]_ , \new_[31938]_ ,
    \new_[31942]_ , \new_[31943]_ , \new_[31947]_ , \new_[31948]_ ,
    \new_[31949]_ , \new_[31953]_ , \new_[31954]_ , \new_[31958]_ ,
    \new_[31959]_ , \new_[31960]_ , \new_[31964]_ , \new_[31965]_ ,
    \new_[31969]_ , \new_[31970]_ , \new_[31971]_ , \new_[31975]_ ,
    \new_[31976]_ , \new_[31980]_ , \new_[31981]_ , \new_[31982]_ ,
    \new_[31986]_ , \new_[31987]_ , \new_[31991]_ , \new_[31992]_ ,
    \new_[31993]_ , \new_[31997]_ , \new_[31998]_ , \new_[32002]_ ,
    \new_[32003]_ , \new_[32004]_ , \new_[32008]_ , \new_[32009]_ ,
    \new_[32013]_ , \new_[32014]_ , \new_[32015]_ , \new_[32019]_ ,
    \new_[32020]_ , \new_[32024]_ , \new_[32025]_ , \new_[32026]_ ,
    \new_[32030]_ , \new_[32031]_ , \new_[32035]_ , \new_[32036]_ ,
    \new_[32037]_ , \new_[32041]_ , \new_[32042]_ , \new_[32046]_ ,
    \new_[32047]_ , \new_[32048]_ , \new_[32052]_ , \new_[32053]_ ,
    \new_[32057]_ , \new_[32058]_ , \new_[32059]_ , \new_[32063]_ ,
    \new_[32064]_ , \new_[32068]_ , \new_[32069]_ , \new_[32070]_ ,
    \new_[32074]_ , \new_[32075]_ , \new_[32079]_ , \new_[32080]_ ,
    \new_[32081]_ , \new_[32085]_ , \new_[32086]_ , \new_[32090]_ ,
    \new_[32091]_ , \new_[32092]_ , \new_[32096]_ , \new_[32097]_ ,
    \new_[32101]_ , \new_[32102]_ , \new_[32103]_ , \new_[32107]_ ,
    \new_[32108]_ , \new_[32112]_ , \new_[32113]_ , \new_[32114]_ ,
    \new_[32118]_ , \new_[32119]_ , \new_[32123]_ , \new_[32124]_ ,
    \new_[32125]_ , \new_[32129]_ , \new_[32130]_ , \new_[32134]_ ,
    \new_[32135]_ , \new_[32136]_ , \new_[32140]_ , \new_[32141]_ ,
    \new_[32145]_ , \new_[32146]_ , \new_[32147]_ , \new_[32151]_ ,
    \new_[32152]_ , \new_[32156]_ , \new_[32157]_ , \new_[32158]_ ,
    \new_[32162]_ , \new_[32163]_ , \new_[32167]_ , \new_[32168]_ ,
    \new_[32169]_ , \new_[32173]_ , \new_[32174]_ , \new_[32178]_ ,
    \new_[32179]_ , \new_[32180]_ , \new_[32184]_ , \new_[32185]_ ,
    \new_[32189]_ , \new_[32190]_ , \new_[32191]_ , \new_[32195]_ ,
    \new_[32196]_ , \new_[32200]_ , \new_[32201]_ , \new_[32202]_ ,
    \new_[32206]_ , \new_[32207]_ , \new_[32211]_ , \new_[32212]_ ,
    \new_[32213]_ , \new_[32217]_ , \new_[32218]_ , \new_[32222]_ ,
    \new_[32223]_ , \new_[32224]_ , \new_[32228]_ , \new_[32229]_ ,
    \new_[32233]_ , \new_[32234]_ , \new_[32235]_ , \new_[32239]_ ,
    \new_[32240]_ , \new_[32244]_ , \new_[32245]_ , \new_[32246]_ ,
    \new_[32250]_ , \new_[32251]_ , \new_[32255]_ , \new_[32256]_ ,
    \new_[32257]_ , \new_[32261]_ , \new_[32262]_ , \new_[32266]_ ,
    \new_[32267]_ , \new_[32268]_ , \new_[32272]_ , \new_[32273]_ ,
    \new_[32277]_ , \new_[32278]_ , \new_[32279]_ , \new_[32283]_ ,
    \new_[32284]_ , \new_[32288]_ , \new_[32289]_ , \new_[32290]_ ,
    \new_[32294]_ , \new_[32295]_ , \new_[32299]_ , \new_[32300]_ ,
    \new_[32301]_ , \new_[32305]_ , \new_[32306]_ , \new_[32310]_ ,
    \new_[32311]_ , \new_[32312]_ , \new_[32316]_ , \new_[32317]_ ,
    \new_[32321]_ , \new_[32322]_ , \new_[32323]_ , \new_[32327]_ ,
    \new_[32328]_ , \new_[32332]_ , \new_[32333]_ , \new_[32334]_ ,
    \new_[32338]_ , \new_[32339]_ , \new_[32343]_ , \new_[32344]_ ,
    \new_[32345]_ , \new_[32349]_ , \new_[32350]_ , \new_[32354]_ ,
    \new_[32355]_ , \new_[32356]_ , \new_[32360]_ , \new_[32361]_ ,
    \new_[32365]_ , \new_[32366]_ , \new_[32367]_ , \new_[32371]_ ,
    \new_[32372]_ , \new_[32376]_ , \new_[32377]_ , \new_[32378]_ ,
    \new_[32382]_ , \new_[32383]_ , \new_[32387]_ , \new_[32388]_ ,
    \new_[32389]_ , \new_[32393]_ , \new_[32394]_ , \new_[32398]_ ,
    \new_[32399]_ , \new_[32400]_ , \new_[32404]_ , \new_[32405]_ ,
    \new_[32409]_ , \new_[32410]_ , \new_[32411]_ , \new_[32415]_ ,
    \new_[32416]_ , \new_[32420]_ , \new_[32421]_ , \new_[32422]_ ,
    \new_[32426]_ , \new_[32427]_ , \new_[32431]_ , \new_[32432]_ ,
    \new_[32433]_ , \new_[32437]_ , \new_[32438]_ , \new_[32442]_ ,
    \new_[32443]_ , \new_[32444]_ , \new_[32448]_ , \new_[32449]_ ,
    \new_[32453]_ , \new_[32454]_ , \new_[32455]_ , \new_[32459]_ ,
    \new_[32460]_ , \new_[32464]_ , \new_[32465]_ , \new_[32466]_ ,
    \new_[32470]_ , \new_[32471]_ , \new_[32475]_ , \new_[32476]_ ,
    \new_[32477]_ , \new_[32481]_ , \new_[32482]_ , \new_[32486]_ ,
    \new_[32487]_ , \new_[32488]_ , \new_[32492]_ , \new_[32493]_ ,
    \new_[32497]_ , \new_[32498]_ , \new_[32499]_ , \new_[32503]_ ,
    \new_[32504]_ , \new_[32508]_ , \new_[32509]_ , \new_[32510]_ ,
    \new_[32514]_ , \new_[32515]_ , \new_[32519]_ , \new_[32520]_ ,
    \new_[32521]_ , \new_[32525]_ , \new_[32526]_ , \new_[32530]_ ,
    \new_[32531]_ , \new_[32532]_ , \new_[32536]_ , \new_[32537]_ ,
    \new_[32541]_ , \new_[32542]_ , \new_[32543]_ , \new_[32547]_ ,
    \new_[32548]_ , \new_[32552]_ , \new_[32553]_ , \new_[32554]_ ,
    \new_[32558]_ , \new_[32559]_ , \new_[32563]_ , \new_[32564]_ ,
    \new_[32565]_ , \new_[32569]_ , \new_[32570]_ , \new_[32574]_ ,
    \new_[32575]_ , \new_[32576]_ , \new_[32580]_ , \new_[32581]_ ,
    \new_[32585]_ , \new_[32586]_ , \new_[32587]_ , \new_[32591]_ ,
    \new_[32592]_ , \new_[32596]_ , \new_[32597]_ , \new_[32598]_ ,
    \new_[32602]_ , \new_[32603]_ , \new_[32607]_ , \new_[32608]_ ,
    \new_[32609]_ , \new_[32613]_ , \new_[32614]_ , \new_[32618]_ ,
    \new_[32619]_ , \new_[32620]_ , \new_[32624]_ , \new_[32625]_ ,
    \new_[32629]_ , \new_[32630]_ , \new_[32631]_ , \new_[32635]_ ,
    \new_[32636]_ , \new_[32640]_ , \new_[32641]_ , \new_[32642]_ ,
    \new_[32646]_ , \new_[32647]_ , \new_[32651]_ , \new_[32652]_ ,
    \new_[32653]_ , \new_[32657]_ , \new_[32658]_ , \new_[32662]_ ,
    \new_[32663]_ , \new_[32664]_ , \new_[32668]_ , \new_[32669]_ ,
    \new_[32673]_ , \new_[32674]_ , \new_[32675]_ , \new_[32679]_ ,
    \new_[32680]_ , \new_[32684]_ , \new_[32685]_ , \new_[32686]_ ,
    \new_[32690]_ , \new_[32691]_ , \new_[32695]_ , \new_[32696]_ ,
    \new_[32697]_ , \new_[32701]_ , \new_[32702]_ , \new_[32706]_ ,
    \new_[32707]_ , \new_[32708]_ , \new_[32712]_ , \new_[32713]_ ,
    \new_[32717]_ , \new_[32718]_ , \new_[32719]_ , \new_[32723]_ ,
    \new_[32724]_ , \new_[32728]_ , \new_[32729]_ , \new_[32730]_ ,
    \new_[32734]_ , \new_[32735]_ , \new_[32739]_ , \new_[32740]_ ,
    \new_[32741]_ , \new_[32745]_ , \new_[32746]_ , \new_[32750]_ ,
    \new_[32751]_ , \new_[32752]_ , \new_[32756]_ , \new_[32757]_ ,
    \new_[32761]_ , \new_[32762]_ , \new_[32763]_ , \new_[32767]_ ,
    \new_[32768]_ , \new_[32772]_ , \new_[32773]_ , \new_[32774]_ ,
    \new_[32778]_ , \new_[32779]_ , \new_[32783]_ , \new_[32784]_ ,
    \new_[32785]_ , \new_[32789]_ , \new_[32790]_ , \new_[32794]_ ,
    \new_[32795]_ , \new_[32796]_ , \new_[32800]_ , \new_[32801]_ ,
    \new_[32805]_ , \new_[32806]_ , \new_[32807]_ , \new_[32811]_ ,
    \new_[32812]_ , \new_[32816]_ , \new_[32817]_ , \new_[32818]_ ,
    \new_[32822]_ , \new_[32823]_ , \new_[32827]_ , \new_[32828]_ ,
    \new_[32829]_ , \new_[32833]_ , \new_[32834]_ , \new_[32838]_ ,
    \new_[32839]_ , \new_[32840]_ , \new_[32844]_ , \new_[32845]_ ,
    \new_[32849]_ , \new_[32850]_ , \new_[32851]_ , \new_[32855]_ ,
    \new_[32856]_ , \new_[32860]_ , \new_[32861]_ , \new_[32862]_ ,
    \new_[32866]_ , \new_[32867]_ , \new_[32871]_ , \new_[32872]_ ,
    \new_[32873]_ , \new_[32877]_ , \new_[32878]_ , \new_[32882]_ ,
    \new_[32883]_ , \new_[32884]_ , \new_[32888]_ , \new_[32889]_ ,
    \new_[32893]_ , \new_[32894]_ , \new_[32895]_ , \new_[32899]_ ,
    \new_[32900]_ , \new_[32904]_ , \new_[32905]_ , \new_[32906]_ ,
    \new_[32910]_ , \new_[32911]_ , \new_[32915]_ , \new_[32916]_ ,
    \new_[32917]_ , \new_[32921]_ , \new_[32922]_ , \new_[32926]_ ,
    \new_[32927]_ , \new_[32928]_ , \new_[32932]_ , \new_[32933]_ ,
    \new_[32937]_ , \new_[32938]_ , \new_[32939]_ , \new_[32943]_ ,
    \new_[32944]_ , \new_[32948]_ , \new_[32949]_ , \new_[32950]_ ,
    \new_[32954]_ , \new_[32955]_ , \new_[32959]_ , \new_[32960]_ ,
    \new_[32961]_ , \new_[32965]_ , \new_[32966]_ , \new_[32970]_ ,
    \new_[32971]_ , \new_[32972]_ , \new_[32976]_ , \new_[32977]_ ,
    \new_[32981]_ , \new_[32982]_ , \new_[32983]_ , \new_[32987]_ ,
    \new_[32988]_ , \new_[32992]_ , \new_[32993]_ , \new_[32994]_ ,
    \new_[32998]_ , \new_[32999]_ , \new_[33003]_ , \new_[33004]_ ,
    \new_[33005]_ , \new_[33009]_ , \new_[33010]_ , \new_[33014]_ ,
    \new_[33015]_ , \new_[33016]_ , \new_[33020]_ , \new_[33021]_ ,
    \new_[33025]_ , \new_[33026]_ , \new_[33027]_ , \new_[33031]_ ,
    \new_[33032]_ , \new_[33036]_ , \new_[33037]_ , \new_[33038]_ ,
    \new_[33042]_ , \new_[33043]_ , \new_[33047]_ , \new_[33048]_ ,
    \new_[33049]_ , \new_[33053]_ , \new_[33054]_ , \new_[33058]_ ,
    \new_[33059]_ , \new_[33060]_ , \new_[33064]_ , \new_[33065]_ ,
    \new_[33069]_ , \new_[33070]_ , \new_[33071]_ , \new_[33075]_ ,
    \new_[33076]_ , \new_[33080]_ , \new_[33081]_ , \new_[33082]_ ,
    \new_[33086]_ , \new_[33087]_ , \new_[33091]_ , \new_[33092]_ ,
    \new_[33093]_ , \new_[33097]_ , \new_[33098]_ , \new_[33102]_ ,
    \new_[33103]_ , \new_[33104]_ , \new_[33108]_ , \new_[33109]_ ,
    \new_[33113]_ , \new_[33114]_ , \new_[33115]_ , \new_[33119]_ ,
    \new_[33120]_ , \new_[33124]_ , \new_[33125]_ , \new_[33126]_ ,
    \new_[33130]_ , \new_[33131]_ , \new_[33135]_ , \new_[33136]_ ,
    \new_[33137]_ , \new_[33141]_ , \new_[33142]_ , \new_[33146]_ ,
    \new_[33147]_ , \new_[33148]_ , \new_[33152]_ , \new_[33153]_ ,
    \new_[33157]_ , \new_[33158]_ , \new_[33159]_ , \new_[33163]_ ,
    \new_[33164]_ , \new_[33168]_ , \new_[33169]_ , \new_[33170]_ ,
    \new_[33174]_ , \new_[33175]_ , \new_[33179]_ , \new_[33180]_ ,
    \new_[33181]_ , \new_[33185]_ , \new_[33186]_ , \new_[33190]_ ,
    \new_[33191]_ , \new_[33192]_ , \new_[33196]_ , \new_[33197]_ ,
    \new_[33201]_ , \new_[33202]_ , \new_[33203]_ , \new_[33207]_ ,
    \new_[33208]_ , \new_[33212]_ , \new_[33213]_ , \new_[33214]_ ,
    \new_[33218]_ , \new_[33219]_ , \new_[33223]_ , \new_[33224]_ ,
    \new_[33225]_ , \new_[33229]_ , \new_[33230]_ , \new_[33234]_ ,
    \new_[33235]_ , \new_[33236]_ , \new_[33240]_ , \new_[33241]_ ,
    \new_[33245]_ , \new_[33246]_ , \new_[33247]_ , \new_[33251]_ ,
    \new_[33252]_ , \new_[33256]_ , \new_[33257]_ , \new_[33258]_ ,
    \new_[33262]_ , \new_[33263]_ , \new_[33267]_ , \new_[33268]_ ,
    \new_[33269]_ , \new_[33273]_ , \new_[33274]_ , \new_[33278]_ ,
    \new_[33279]_ , \new_[33280]_ , \new_[33284]_ , \new_[33285]_ ,
    \new_[33289]_ , \new_[33290]_ , \new_[33291]_ , \new_[33295]_ ,
    \new_[33296]_ , \new_[33300]_ , \new_[33301]_ , \new_[33302]_ ,
    \new_[33306]_ , \new_[33307]_ , \new_[33311]_ , \new_[33312]_ ,
    \new_[33313]_ , \new_[33317]_ , \new_[33318]_ , \new_[33322]_ ,
    \new_[33323]_ , \new_[33324]_ , \new_[33328]_ , \new_[33329]_ ,
    \new_[33333]_ , \new_[33334]_ , \new_[33335]_ , \new_[33339]_ ,
    \new_[33340]_ , \new_[33344]_ , \new_[33345]_ , \new_[33346]_ ,
    \new_[33350]_ , \new_[33351]_ , \new_[33355]_ , \new_[33356]_ ,
    \new_[33357]_ , \new_[33361]_ , \new_[33362]_ , \new_[33366]_ ,
    \new_[33367]_ , \new_[33368]_ , \new_[33372]_ , \new_[33373]_ ,
    \new_[33377]_ , \new_[33378]_ , \new_[33379]_ , \new_[33383]_ ,
    \new_[33384]_ , \new_[33388]_ , \new_[33389]_ , \new_[33390]_ ,
    \new_[33394]_ , \new_[33395]_ , \new_[33399]_ , \new_[33400]_ ,
    \new_[33401]_ , \new_[33405]_ , \new_[33406]_ , \new_[33410]_ ,
    \new_[33411]_ , \new_[33412]_ , \new_[33416]_ , \new_[33417]_ ,
    \new_[33421]_ , \new_[33422]_ , \new_[33423]_ , \new_[33427]_ ,
    \new_[33428]_ , \new_[33432]_ , \new_[33433]_ , \new_[33434]_ ,
    \new_[33438]_ , \new_[33439]_ , \new_[33443]_ , \new_[33444]_ ,
    \new_[33445]_ , \new_[33449]_ , \new_[33450]_ , \new_[33454]_ ,
    \new_[33455]_ , \new_[33456]_ , \new_[33460]_ , \new_[33461]_ ,
    \new_[33465]_ , \new_[33466]_ , \new_[33467]_ , \new_[33471]_ ,
    \new_[33472]_ , \new_[33476]_ , \new_[33477]_ , \new_[33478]_ ,
    \new_[33482]_ , \new_[33483]_ , \new_[33487]_ , \new_[33488]_ ,
    \new_[33489]_ , \new_[33493]_ , \new_[33494]_ , \new_[33498]_ ,
    \new_[33499]_ , \new_[33500]_ , \new_[33504]_ , \new_[33505]_ ,
    \new_[33509]_ , \new_[33510]_ , \new_[33511]_ , \new_[33515]_ ,
    \new_[33516]_ , \new_[33520]_ , \new_[33521]_ , \new_[33522]_ ,
    \new_[33526]_ , \new_[33527]_ , \new_[33531]_ , \new_[33532]_ ,
    \new_[33533]_ , \new_[33537]_ , \new_[33538]_ , \new_[33542]_ ,
    \new_[33543]_ , \new_[33544]_ , \new_[33548]_ , \new_[33549]_ ,
    \new_[33553]_ , \new_[33554]_ , \new_[33555]_ , \new_[33559]_ ,
    \new_[33560]_ , \new_[33564]_ , \new_[33565]_ , \new_[33566]_ ,
    \new_[33570]_ , \new_[33571]_ , \new_[33575]_ , \new_[33576]_ ,
    \new_[33577]_ , \new_[33581]_ , \new_[33582]_ , \new_[33586]_ ,
    \new_[33587]_ , \new_[33588]_ , \new_[33592]_ , \new_[33593]_ ,
    \new_[33597]_ , \new_[33598]_ , \new_[33599]_ , \new_[33603]_ ,
    \new_[33604]_ , \new_[33608]_ , \new_[33609]_ , \new_[33610]_ ,
    \new_[33614]_ , \new_[33615]_ , \new_[33619]_ , \new_[33620]_ ,
    \new_[33621]_ , \new_[33625]_ , \new_[33626]_ , \new_[33630]_ ,
    \new_[33631]_ , \new_[33632]_ , \new_[33636]_ , \new_[33637]_ ,
    \new_[33641]_ , \new_[33642]_ , \new_[33643]_ , \new_[33647]_ ,
    \new_[33648]_ , \new_[33652]_ , \new_[33653]_ , \new_[33654]_ ,
    \new_[33658]_ , \new_[33659]_ , \new_[33663]_ , \new_[33664]_ ,
    \new_[33665]_ , \new_[33669]_ , \new_[33670]_ , \new_[33674]_ ,
    \new_[33675]_ , \new_[33676]_ , \new_[33680]_ , \new_[33681]_ ,
    \new_[33685]_ , \new_[33686]_ , \new_[33687]_ , \new_[33691]_ ,
    \new_[33692]_ , \new_[33696]_ , \new_[33697]_ , \new_[33698]_ ,
    \new_[33702]_ , \new_[33703]_ , \new_[33707]_ , \new_[33708]_ ,
    \new_[33709]_ , \new_[33713]_ , \new_[33714]_ , \new_[33718]_ ,
    \new_[33719]_ , \new_[33720]_ , \new_[33724]_ , \new_[33725]_ ,
    \new_[33729]_ , \new_[33730]_ , \new_[33731]_ , \new_[33735]_ ,
    \new_[33736]_ , \new_[33740]_ , \new_[33741]_ , \new_[33742]_ ,
    \new_[33746]_ , \new_[33747]_ , \new_[33751]_ , \new_[33752]_ ,
    \new_[33753]_ , \new_[33757]_ , \new_[33758]_ , \new_[33762]_ ,
    \new_[33763]_ , \new_[33764]_ , \new_[33768]_ , \new_[33769]_ ,
    \new_[33773]_ , \new_[33774]_ , \new_[33775]_ , \new_[33779]_ ,
    \new_[33780]_ , \new_[33784]_ , \new_[33785]_ , \new_[33786]_ ,
    \new_[33790]_ , \new_[33791]_ , \new_[33795]_ , \new_[33796]_ ,
    \new_[33797]_ , \new_[33801]_ , \new_[33802]_ , \new_[33806]_ ,
    \new_[33807]_ , \new_[33808]_ , \new_[33812]_ , \new_[33813]_ ,
    \new_[33817]_ , \new_[33818]_ , \new_[33819]_ , \new_[33823]_ ,
    \new_[33824]_ , \new_[33828]_ , \new_[33829]_ , \new_[33830]_ ,
    \new_[33834]_ , \new_[33835]_ , \new_[33839]_ , \new_[33840]_ ,
    \new_[33841]_ , \new_[33845]_ , \new_[33846]_ , \new_[33850]_ ,
    \new_[33851]_ , \new_[33852]_ , \new_[33856]_ , \new_[33857]_ ,
    \new_[33861]_ , \new_[33862]_ , \new_[33863]_ , \new_[33867]_ ,
    \new_[33868]_ , \new_[33872]_ , \new_[33873]_ , \new_[33874]_ ,
    \new_[33878]_ , \new_[33879]_ , \new_[33883]_ , \new_[33884]_ ,
    \new_[33885]_ , \new_[33889]_ , \new_[33890]_ , \new_[33894]_ ,
    \new_[33895]_ , \new_[33896]_ , \new_[33900]_ , \new_[33901]_ ,
    \new_[33905]_ , \new_[33906]_ , \new_[33907]_ , \new_[33911]_ ,
    \new_[33912]_ , \new_[33916]_ , \new_[33917]_ , \new_[33918]_ ,
    \new_[33922]_ , \new_[33923]_ , \new_[33927]_ , \new_[33928]_ ,
    \new_[33929]_ , \new_[33933]_ , \new_[33934]_ , \new_[33938]_ ,
    \new_[33939]_ , \new_[33940]_ , \new_[33944]_ , \new_[33945]_ ,
    \new_[33949]_ , \new_[33950]_ , \new_[33951]_ , \new_[33955]_ ,
    \new_[33956]_ , \new_[33960]_ , \new_[33961]_ , \new_[33962]_ ,
    \new_[33966]_ , \new_[33967]_ , \new_[33971]_ , \new_[33972]_ ,
    \new_[33973]_ , \new_[33977]_ , \new_[33978]_ , \new_[33982]_ ,
    \new_[33983]_ , \new_[33984]_ , \new_[33988]_ , \new_[33989]_ ,
    \new_[33993]_ , \new_[33994]_ , \new_[33995]_ , \new_[33999]_ ,
    \new_[34000]_ , \new_[34004]_ , \new_[34005]_ , \new_[34006]_ ,
    \new_[34010]_ , \new_[34011]_ , \new_[34015]_ , \new_[34016]_ ,
    \new_[34017]_ , \new_[34021]_ , \new_[34022]_ , \new_[34026]_ ,
    \new_[34027]_ , \new_[34028]_ , \new_[34032]_ , \new_[34033]_ ,
    \new_[34037]_ , \new_[34038]_ , \new_[34039]_ , \new_[34043]_ ,
    \new_[34044]_ , \new_[34048]_ , \new_[34049]_ , \new_[34050]_ ,
    \new_[34054]_ , \new_[34055]_ , \new_[34059]_ , \new_[34060]_ ,
    \new_[34061]_ , \new_[34065]_ , \new_[34066]_ , \new_[34070]_ ,
    \new_[34071]_ , \new_[34072]_ , \new_[34076]_ , \new_[34077]_ ,
    \new_[34081]_ , \new_[34082]_ , \new_[34083]_ , \new_[34087]_ ,
    \new_[34088]_ , \new_[34092]_ , \new_[34093]_ , \new_[34094]_ ,
    \new_[34098]_ , \new_[34099]_ , \new_[34103]_ , \new_[34104]_ ,
    \new_[34105]_ , \new_[34109]_ , \new_[34110]_ , \new_[34114]_ ,
    \new_[34115]_ , \new_[34116]_ , \new_[34120]_ , \new_[34121]_ ,
    \new_[34125]_ , \new_[34126]_ , \new_[34127]_ , \new_[34131]_ ,
    \new_[34132]_ , \new_[34136]_ , \new_[34137]_ , \new_[34138]_ ,
    \new_[34142]_ , \new_[34143]_ , \new_[34147]_ , \new_[34148]_ ,
    \new_[34149]_ , \new_[34153]_ , \new_[34154]_ , \new_[34158]_ ,
    \new_[34159]_ , \new_[34160]_ , \new_[34164]_ , \new_[34165]_ ,
    \new_[34169]_ , \new_[34170]_ , \new_[34171]_ , \new_[34175]_ ,
    \new_[34176]_ , \new_[34180]_ , \new_[34181]_ , \new_[34182]_ ,
    \new_[34186]_ , \new_[34187]_ , \new_[34191]_ , \new_[34192]_ ,
    \new_[34193]_ , \new_[34197]_ , \new_[34198]_ , \new_[34202]_ ,
    \new_[34203]_ , \new_[34204]_ , \new_[34208]_ , \new_[34209]_ ,
    \new_[34213]_ , \new_[34214]_ , \new_[34215]_ , \new_[34219]_ ,
    \new_[34220]_ , \new_[34224]_ , \new_[34225]_ , \new_[34226]_ ,
    \new_[34230]_ , \new_[34231]_ , \new_[34235]_ , \new_[34236]_ ,
    \new_[34237]_ , \new_[34241]_ , \new_[34242]_ , \new_[34246]_ ,
    \new_[34247]_ , \new_[34248]_ , \new_[34252]_ , \new_[34253]_ ,
    \new_[34257]_ , \new_[34258]_ , \new_[34259]_ , \new_[34263]_ ,
    \new_[34264]_ , \new_[34268]_ , \new_[34269]_ , \new_[34270]_ ,
    \new_[34274]_ , \new_[34275]_ , \new_[34279]_ , \new_[34280]_ ,
    \new_[34281]_ , \new_[34285]_ , \new_[34286]_ , \new_[34290]_ ,
    \new_[34291]_ , \new_[34292]_ , \new_[34296]_ , \new_[34297]_ ,
    \new_[34301]_ , \new_[34302]_ , \new_[34303]_ , \new_[34307]_ ,
    \new_[34308]_ , \new_[34312]_ , \new_[34313]_ , \new_[34314]_ ,
    \new_[34318]_ , \new_[34319]_ , \new_[34323]_ , \new_[34324]_ ,
    \new_[34325]_ , \new_[34329]_ , \new_[34330]_ , \new_[34334]_ ,
    \new_[34335]_ , \new_[34336]_ , \new_[34340]_ , \new_[34341]_ ,
    \new_[34345]_ , \new_[34346]_ , \new_[34347]_ , \new_[34351]_ ,
    \new_[34352]_ , \new_[34356]_ , \new_[34357]_ , \new_[34358]_ ,
    \new_[34362]_ , \new_[34363]_ , \new_[34367]_ , \new_[34368]_ ,
    \new_[34369]_ , \new_[34373]_ , \new_[34374]_ , \new_[34378]_ ,
    \new_[34379]_ , \new_[34380]_ , \new_[34384]_ , \new_[34385]_ ,
    \new_[34389]_ , \new_[34390]_ , \new_[34391]_ , \new_[34395]_ ,
    \new_[34396]_ , \new_[34400]_ , \new_[34401]_ , \new_[34402]_ ,
    \new_[34406]_ , \new_[34407]_ , \new_[34411]_ , \new_[34412]_ ,
    \new_[34413]_ , \new_[34417]_ , \new_[34418]_ , \new_[34422]_ ,
    \new_[34423]_ , \new_[34424]_ , \new_[34428]_ , \new_[34429]_ ,
    \new_[34433]_ , \new_[34434]_ , \new_[34435]_ , \new_[34439]_ ,
    \new_[34440]_ , \new_[34444]_ , \new_[34445]_ , \new_[34446]_ ,
    \new_[34450]_ , \new_[34451]_ , \new_[34455]_ , \new_[34456]_ ,
    \new_[34457]_ , \new_[34461]_ , \new_[34462]_ , \new_[34466]_ ,
    \new_[34467]_ , \new_[34468]_ , \new_[34472]_ , \new_[34473]_ ,
    \new_[34477]_ , \new_[34478]_ , \new_[34479]_ , \new_[34483]_ ,
    \new_[34484]_ , \new_[34488]_ , \new_[34489]_ , \new_[34490]_ ,
    \new_[34494]_ , \new_[34495]_ , \new_[34499]_ , \new_[34500]_ ,
    \new_[34501]_ , \new_[34505]_ , \new_[34506]_ , \new_[34510]_ ,
    \new_[34511]_ , \new_[34512]_ , \new_[34516]_ , \new_[34517]_ ,
    \new_[34521]_ , \new_[34522]_ , \new_[34523]_ , \new_[34527]_ ,
    \new_[34528]_ , \new_[34532]_ , \new_[34533]_ , \new_[34534]_ ,
    \new_[34538]_ , \new_[34539]_ , \new_[34543]_ , \new_[34544]_ ,
    \new_[34545]_ , \new_[34549]_ , \new_[34550]_ , \new_[34554]_ ,
    \new_[34555]_ , \new_[34556]_ , \new_[34560]_ , \new_[34561]_ ,
    \new_[34565]_ , \new_[34566]_ , \new_[34567]_ , \new_[34571]_ ,
    \new_[34572]_ , \new_[34576]_ , \new_[34577]_ , \new_[34578]_ ,
    \new_[34582]_ , \new_[34583]_ , \new_[34587]_ , \new_[34588]_ ,
    \new_[34589]_ , \new_[34593]_ , \new_[34594]_ , \new_[34598]_ ,
    \new_[34599]_ , \new_[34600]_ , \new_[34604]_ , \new_[34605]_ ,
    \new_[34609]_ , \new_[34610]_ , \new_[34611]_ , \new_[34615]_ ,
    \new_[34616]_ , \new_[34620]_ , \new_[34621]_ , \new_[34622]_ ,
    \new_[34626]_ , \new_[34627]_ , \new_[34631]_ , \new_[34632]_ ,
    \new_[34633]_ , \new_[34637]_ , \new_[34638]_ , \new_[34642]_ ,
    \new_[34643]_ , \new_[34644]_ , \new_[34648]_ , \new_[34649]_ ,
    \new_[34653]_ , \new_[34654]_ , \new_[34655]_ , \new_[34659]_ ,
    \new_[34660]_ , \new_[34664]_ , \new_[34665]_ , \new_[34666]_ ,
    \new_[34670]_ , \new_[34671]_ , \new_[34675]_ , \new_[34676]_ ,
    \new_[34677]_ , \new_[34681]_ , \new_[34682]_ , \new_[34686]_ ,
    \new_[34687]_ , \new_[34688]_ , \new_[34692]_ , \new_[34693]_ ,
    \new_[34697]_ , \new_[34698]_ , \new_[34699]_ , \new_[34703]_ ,
    \new_[34704]_ , \new_[34708]_ , \new_[34709]_ , \new_[34710]_ ,
    \new_[34714]_ , \new_[34715]_ , \new_[34719]_ , \new_[34720]_ ,
    \new_[34721]_ , \new_[34725]_ , \new_[34726]_ , \new_[34730]_ ,
    \new_[34731]_ , \new_[34732]_ , \new_[34736]_ , \new_[34737]_ ,
    \new_[34741]_ , \new_[34742]_ , \new_[34743]_ , \new_[34747]_ ,
    \new_[34748]_ , \new_[34752]_ , \new_[34753]_ , \new_[34754]_ ,
    \new_[34758]_ , \new_[34759]_ , \new_[34763]_ , \new_[34764]_ ,
    \new_[34765]_ , \new_[34769]_ , \new_[34770]_ , \new_[34774]_ ,
    \new_[34775]_ , \new_[34776]_ , \new_[34780]_ , \new_[34781]_ ,
    \new_[34785]_ , \new_[34786]_ , \new_[34787]_ , \new_[34791]_ ,
    \new_[34792]_ , \new_[34796]_ , \new_[34797]_ , \new_[34798]_ ,
    \new_[34802]_ , \new_[34803]_ , \new_[34807]_ , \new_[34808]_ ,
    \new_[34809]_ , \new_[34813]_ , \new_[34814]_ , \new_[34818]_ ,
    \new_[34819]_ , \new_[34820]_ , \new_[34824]_ , \new_[34825]_ ,
    \new_[34829]_ , \new_[34830]_ , \new_[34831]_ , \new_[34835]_ ,
    \new_[34836]_ , \new_[34840]_ , \new_[34841]_ , \new_[34842]_ ,
    \new_[34846]_ , \new_[34847]_ , \new_[34851]_ , \new_[34852]_ ,
    \new_[34853]_ , \new_[34857]_ , \new_[34858]_ , \new_[34862]_ ,
    \new_[34863]_ , \new_[34864]_ , \new_[34868]_ , \new_[34869]_ ,
    \new_[34873]_ , \new_[34874]_ , \new_[34875]_ , \new_[34879]_ ,
    \new_[34880]_ , \new_[34884]_ , \new_[34885]_ , \new_[34886]_ ,
    \new_[34890]_ , \new_[34891]_ , \new_[34895]_ , \new_[34896]_ ,
    \new_[34897]_ , \new_[34901]_ , \new_[34902]_ , \new_[34906]_ ,
    \new_[34907]_ , \new_[34908]_ , \new_[34912]_ , \new_[34913]_ ,
    \new_[34917]_ , \new_[34918]_ , \new_[34919]_ , \new_[34923]_ ,
    \new_[34924]_ , \new_[34928]_ , \new_[34929]_ , \new_[34930]_ ,
    \new_[34934]_ , \new_[34935]_ , \new_[34939]_ , \new_[34940]_ ,
    \new_[34941]_ , \new_[34945]_ , \new_[34946]_ , \new_[34950]_ ,
    \new_[34951]_ , \new_[34952]_ , \new_[34956]_ , \new_[34957]_ ,
    \new_[34961]_ , \new_[34962]_ , \new_[34963]_ , \new_[34967]_ ,
    \new_[34968]_ , \new_[34972]_ , \new_[34973]_ , \new_[34974]_ ,
    \new_[34978]_ , \new_[34979]_ , \new_[34983]_ , \new_[34984]_ ,
    \new_[34985]_ , \new_[34989]_ , \new_[34990]_ , \new_[34994]_ ,
    \new_[34995]_ , \new_[34996]_ , \new_[35000]_ , \new_[35001]_ ,
    \new_[35005]_ , \new_[35006]_ , \new_[35007]_ , \new_[35011]_ ,
    \new_[35012]_ , \new_[35016]_ , \new_[35017]_ , \new_[35018]_ ,
    \new_[35022]_ , \new_[35023]_ , \new_[35027]_ , \new_[35028]_ ,
    \new_[35029]_ , \new_[35033]_ , \new_[35034]_ , \new_[35038]_ ,
    \new_[35039]_ , \new_[35040]_ , \new_[35044]_ , \new_[35045]_ ,
    \new_[35049]_ , \new_[35050]_ , \new_[35051]_ , \new_[35055]_ ,
    \new_[35056]_ , \new_[35060]_ , \new_[35061]_ , \new_[35062]_ ,
    \new_[35066]_ , \new_[35067]_ , \new_[35071]_ , \new_[35072]_ ,
    \new_[35073]_ , \new_[35077]_ , \new_[35078]_ , \new_[35082]_ ,
    \new_[35083]_ , \new_[35084]_ , \new_[35088]_ , \new_[35089]_ ,
    \new_[35093]_ , \new_[35094]_ , \new_[35095]_ , \new_[35099]_ ,
    \new_[35100]_ , \new_[35104]_ , \new_[35105]_ , \new_[35106]_ ,
    \new_[35110]_ , \new_[35111]_ , \new_[35115]_ , \new_[35116]_ ,
    \new_[35117]_ , \new_[35121]_ , \new_[35122]_ , \new_[35126]_ ,
    \new_[35127]_ , \new_[35128]_ , \new_[35132]_ , \new_[35133]_ ,
    \new_[35137]_ , \new_[35138]_ , \new_[35139]_ , \new_[35143]_ ,
    \new_[35144]_ , \new_[35148]_ , \new_[35149]_ , \new_[35150]_ ,
    \new_[35154]_ , \new_[35155]_ , \new_[35159]_ , \new_[35160]_ ,
    \new_[35161]_ , \new_[35165]_ , \new_[35166]_ , \new_[35170]_ ,
    \new_[35171]_ , \new_[35172]_ , \new_[35176]_ , \new_[35177]_ ,
    \new_[35181]_ , \new_[35182]_ , \new_[35183]_ , \new_[35187]_ ,
    \new_[35188]_ , \new_[35192]_ , \new_[35193]_ , \new_[35194]_ ,
    \new_[35198]_ , \new_[35199]_ , \new_[35203]_ , \new_[35204]_ ,
    \new_[35205]_ , \new_[35209]_ , \new_[35210]_ , \new_[35214]_ ,
    \new_[35215]_ , \new_[35216]_ , \new_[35220]_ , \new_[35221]_ ,
    \new_[35225]_ , \new_[35226]_ , \new_[35227]_ , \new_[35231]_ ,
    \new_[35232]_ , \new_[35236]_ , \new_[35237]_ , \new_[35238]_ ,
    \new_[35242]_ , \new_[35243]_ , \new_[35247]_ , \new_[35248]_ ,
    \new_[35249]_ , \new_[35253]_ , \new_[35254]_ , \new_[35258]_ ,
    \new_[35259]_ , \new_[35260]_ , \new_[35264]_ , \new_[35265]_ ,
    \new_[35269]_ , \new_[35270]_ , \new_[35271]_ , \new_[35275]_ ,
    \new_[35276]_ , \new_[35280]_ , \new_[35281]_ , \new_[35282]_ ,
    \new_[35286]_ , \new_[35287]_ , \new_[35291]_ , \new_[35292]_ ,
    \new_[35293]_ , \new_[35297]_ , \new_[35298]_ , \new_[35302]_ ,
    \new_[35303]_ , \new_[35304]_ , \new_[35308]_ , \new_[35309]_ ,
    \new_[35313]_ , \new_[35314]_ , \new_[35315]_ , \new_[35319]_ ,
    \new_[35320]_ , \new_[35324]_ , \new_[35325]_ , \new_[35326]_ ,
    \new_[35330]_ , \new_[35331]_ , \new_[35335]_ , \new_[35336]_ ,
    \new_[35337]_ , \new_[35341]_ , \new_[35342]_ , \new_[35346]_ ,
    \new_[35347]_ , \new_[35348]_ , \new_[35352]_ , \new_[35353]_ ,
    \new_[35357]_ , \new_[35358]_ , \new_[35359]_ , \new_[35363]_ ,
    \new_[35364]_ , \new_[35368]_ , \new_[35369]_ , \new_[35370]_ ,
    \new_[35374]_ , \new_[35375]_ , \new_[35379]_ , \new_[35380]_ ,
    \new_[35381]_ , \new_[35385]_ , \new_[35386]_ , \new_[35390]_ ,
    \new_[35391]_ , \new_[35392]_ , \new_[35396]_ , \new_[35397]_ ,
    \new_[35401]_ , \new_[35402]_ , \new_[35403]_ , \new_[35407]_ ,
    \new_[35408]_ , \new_[35412]_ , \new_[35413]_ , \new_[35414]_ ,
    \new_[35418]_ , \new_[35419]_ , \new_[35423]_ , \new_[35424]_ ,
    \new_[35425]_ , \new_[35429]_ , \new_[35430]_ , \new_[35434]_ ,
    \new_[35435]_ , \new_[35436]_ , \new_[35440]_ , \new_[35441]_ ,
    \new_[35445]_ , \new_[35446]_ , \new_[35447]_ , \new_[35451]_ ,
    \new_[35452]_ , \new_[35456]_ , \new_[35457]_ , \new_[35458]_ ,
    \new_[35462]_ , \new_[35463]_ , \new_[35467]_ , \new_[35468]_ ,
    \new_[35469]_ , \new_[35473]_ , \new_[35474]_ , \new_[35478]_ ,
    \new_[35479]_ , \new_[35480]_ , \new_[35484]_ , \new_[35485]_ ,
    \new_[35489]_ , \new_[35490]_ , \new_[35491]_ , \new_[35495]_ ,
    \new_[35496]_ , \new_[35500]_ , \new_[35501]_ , \new_[35502]_ ,
    \new_[35506]_ , \new_[35507]_ , \new_[35511]_ , \new_[35512]_ ,
    \new_[35513]_ , \new_[35517]_ , \new_[35518]_ , \new_[35522]_ ,
    \new_[35523]_ , \new_[35524]_ , \new_[35528]_ , \new_[35529]_ ,
    \new_[35533]_ , \new_[35534]_ , \new_[35535]_ , \new_[35539]_ ,
    \new_[35540]_ , \new_[35544]_ , \new_[35545]_ , \new_[35546]_ ,
    \new_[35550]_ , \new_[35551]_ , \new_[35555]_ , \new_[35556]_ ,
    \new_[35557]_ , \new_[35561]_ , \new_[35562]_ , \new_[35566]_ ,
    \new_[35567]_ , \new_[35568]_ , \new_[35572]_ , \new_[35573]_ ,
    \new_[35577]_ , \new_[35578]_ , \new_[35579]_ , \new_[35583]_ ,
    \new_[35584]_ , \new_[35588]_ , \new_[35589]_ , \new_[35590]_ ,
    \new_[35594]_ , \new_[35595]_ , \new_[35599]_ , \new_[35600]_ ,
    \new_[35601]_ , \new_[35605]_ , \new_[35606]_ , \new_[35610]_ ,
    \new_[35611]_ , \new_[35612]_ , \new_[35616]_ , \new_[35617]_ ,
    \new_[35621]_ , \new_[35622]_ , \new_[35623]_ , \new_[35627]_ ,
    \new_[35628]_ , \new_[35632]_ , \new_[35633]_ , \new_[35634]_ ,
    \new_[35638]_ , \new_[35639]_ , \new_[35643]_ , \new_[35644]_ ,
    \new_[35645]_ , \new_[35649]_ , \new_[35650]_ , \new_[35654]_ ,
    \new_[35655]_ , \new_[35656]_ , \new_[35660]_ , \new_[35661]_ ,
    \new_[35665]_ , \new_[35666]_ , \new_[35667]_ , \new_[35671]_ ,
    \new_[35672]_ , \new_[35676]_ , \new_[35677]_ , \new_[35678]_ ,
    \new_[35682]_ , \new_[35683]_ , \new_[35687]_ , \new_[35688]_ ,
    \new_[35689]_ , \new_[35693]_ , \new_[35694]_ , \new_[35698]_ ,
    \new_[35699]_ , \new_[35700]_ , \new_[35704]_ , \new_[35705]_ ,
    \new_[35709]_ , \new_[35710]_ , \new_[35711]_ , \new_[35715]_ ,
    \new_[35716]_ , \new_[35720]_ , \new_[35721]_ , \new_[35722]_ ,
    \new_[35726]_ , \new_[35727]_ , \new_[35731]_ , \new_[35732]_ ,
    \new_[35733]_ , \new_[35737]_ , \new_[35738]_ , \new_[35742]_ ,
    \new_[35743]_ , \new_[35744]_ , \new_[35748]_ , \new_[35749]_ ,
    \new_[35753]_ , \new_[35754]_ , \new_[35755]_ , \new_[35759]_ ,
    \new_[35760]_ , \new_[35764]_ , \new_[35765]_ , \new_[35766]_ ,
    \new_[35770]_ , \new_[35771]_ , \new_[35775]_ , \new_[35776]_ ,
    \new_[35777]_ , \new_[35781]_ , \new_[35782]_ , \new_[35786]_ ,
    \new_[35787]_ , \new_[35788]_ , \new_[35792]_ , \new_[35793]_ ,
    \new_[35797]_ , \new_[35798]_ , \new_[35799]_ , \new_[35803]_ ,
    \new_[35804]_ , \new_[35808]_ , \new_[35809]_ , \new_[35810]_ ,
    \new_[35814]_ , \new_[35815]_ , \new_[35819]_ , \new_[35820]_ ,
    \new_[35821]_ , \new_[35825]_ , \new_[35826]_ , \new_[35830]_ ,
    \new_[35831]_ , \new_[35832]_ , \new_[35836]_ , \new_[35837]_ ,
    \new_[35841]_ , \new_[35842]_ , \new_[35843]_ , \new_[35847]_ ,
    \new_[35848]_ , \new_[35852]_ , \new_[35853]_ , \new_[35854]_ ,
    \new_[35858]_ , \new_[35859]_ , \new_[35863]_ , \new_[35864]_ ,
    \new_[35865]_ , \new_[35869]_ , \new_[35870]_ , \new_[35874]_ ,
    \new_[35875]_ , \new_[35876]_ , \new_[35880]_ , \new_[35881]_ ,
    \new_[35885]_ , \new_[35886]_ , \new_[35887]_ , \new_[35891]_ ,
    \new_[35892]_ , \new_[35896]_ , \new_[35897]_ , \new_[35898]_ ,
    \new_[35902]_ , \new_[35903]_ , \new_[35907]_ , \new_[35908]_ ,
    \new_[35909]_ , \new_[35913]_ , \new_[35914]_ , \new_[35918]_ ,
    \new_[35919]_ , \new_[35920]_ , \new_[35924]_ , \new_[35925]_ ,
    \new_[35929]_ , \new_[35930]_ , \new_[35931]_ , \new_[35935]_ ,
    \new_[35936]_ , \new_[35940]_ , \new_[35941]_ , \new_[35942]_ ,
    \new_[35946]_ , \new_[35947]_ , \new_[35951]_ , \new_[35952]_ ,
    \new_[35953]_ , \new_[35957]_ , \new_[35958]_ , \new_[35962]_ ,
    \new_[35963]_ , \new_[35964]_ , \new_[35968]_ , \new_[35969]_ ,
    \new_[35973]_ , \new_[35974]_ , \new_[35975]_ , \new_[35979]_ ,
    \new_[35980]_ , \new_[35984]_ , \new_[35985]_ , \new_[35986]_ ,
    \new_[35990]_ , \new_[35991]_ , \new_[35995]_ , \new_[35996]_ ,
    \new_[35997]_ , \new_[36001]_ , \new_[36002]_ , \new_[36006]_ ,
    \new_[36007]_ , \new_[36008]_ , \new_[36012]_ , \new_[36013]_ ,
    \new_[36017]_ , \new_[36018]_ , \new_[36019]_ , \new_[36023]_ ,
    \new_[36024]_ , \new_[36028]_ , \new_[36029]_ , \new_[36030]_ ,
    \new_[36034]_ , \new_[36035]_ , \new_[36039]_ , \new_[36040]_ ,
    \new_[36041]_ , \new_[36045]_ , \new_[36046]_ , \new_[36050]_ ,
    \new_[36051]_ , \new_[36052]_ , \new_[36056]_ , \new_[36057]_ ,
    \new_[36061]_ , \new_[36062]_ , \new_[36063]_ , \new_[36067]_ ,
    \new_[36068]_ , \new_[36072]_ , \new_[36073]_ , \new_[36074]_ ,
    \new_[36078]_ , \new_[36079]_ , \new_[36083]_ , \new_[36084]_ ,
    \new_[36085]_ , \new_[36089]_ , \new_[36090]_ , \new_[36094]_ ,
    \new_[36095]_ , \new_[36096]_ , \new_[36100]_ , \new_[36101]_ ,
    \new_[36105]_ , \new_[36106]_ , \new_[36107]_ , \new_[36111]_ ,
    \new_[36112]_ , \new_[36116]_ , \new_[36117]_ , \new_[36118]_ ,
    \new_[36122]_ , \new_[36123]_ , \new_[36127]_ , \new_[36128]_ ,
    \new_[36129]_ , \new_[36133]_ , \new_[36134]_ , \new_[36138]_ ,
    \new_[36139]_ , \new_[36140]_ , \new_[36144]_ , \new_[36145]_ ,
    \new_[36149]_ , \new_[36150]_ , \new_[36151]_ , \new_[36155]_ ,
    \new_[36156]_ , \new_[36160]_ , \new_[36161]_ , \new_[36162]_ ,
    \new_[36166]_ , \new_[36167]_ , \new_[36171]_ , \new_[36172]_ ,
    \new_[36173]_ , \new_[36177]_ , \new_[36178]_ , \new_[36182]_ ,
    \new_[36183]_ , \new_[36184]_ , \new_[36188]_ , \new_[36189]_ ,
    \new_[36193]_ , \new_[36194]_ , \new_[36195]_ , \new_[36199]_ ,
    \new_[36200]_ , \new_[36204]_ , \new_[36205]_ , \new_[36206]_ ,
    \new_[36210]_ , \new_[36211]_ , \new_[36215]_ , \new_[36216]_ ,
    \new_[36217]_ , \new_[36221]_ , \new_[36222]_ , \new_[36226]_ ,
    \new_[36227]_ , \new_[36228]_ , \new_[36232]_ , \new_[36233]_ ,
    \new_[36237]_ , \new_[36238]_ , \new_[36239]_ , \new_[36243]_ ,
    \new_[36244]_ , \new_[36248]_ , \new_[36249]_ , \new_[36250]_ ,
    \new_[36254]_ , \new_[36255]_ , \new_[36259]_ , \new_[36260]_ ,
    \new_[36261]_ , \new_[36265]_ , \new_[36266]_ , \new_[36270]_ ,
    \new_[36271]_ , \new_[36272]_ , \new_[36276]_ , \new_[36277]_ ,
    \new_[36281]_ , \new_[36282]_ , \new_[36283]_ , \new_[36287]_ ,
    \new_[36288]_ , \new_[36292]_ , \new_[36293]_ , \new_[36294]_ ,
    \new_[36298]_ , \new_[36299]_ , \new_[36303]_ , \new_[36304]_ ,
    \new_[36305]_ , \new_[36309]_ , \new_[36310]_ , \new_[36314]_ ,
    \new_[36315]_ , \new_[36316]_ , \new_[36320]_ , \new_[36321]_ ,
    \new_[36325]_ , \new_[36326]_ , \new_[36327]_ , \new_[36331]_ ,
    \new_[36332]_ , \new_[36336]_ , \new_[36337]_ , \new_[36338]_ ,
    \new_[36342]_ , \new_[36343]_ , \new_[36347]_ , \new_[36348]_ ,
    \new_[36349]_ , \new_[36353]_ , \new_[36354]_ , \new_[36358]_ ,
    \new_[36359]_ , \new_[36360]_ , \new_[36364]_ , \new_[36365]_ ,
    \new_[36369]_ , \new_[36370]_ , \new_[36371]_ , \new_[36375]_ ,
    \new_[36376]_ , \new_[36380]_ , \new_[36381]_ , \new_[36382]_ ,
    \new_[36386]_ , \new_[36387]_ , \new_[36391]_ , \new_[36392]_ ,
    \new_[36393]_ , \new_[36397]_ , \new_[36398]_ , \new_[36402]_ ,
    \new_[36403]_ , \new_[36404]_ , \new_[36408]_ , \new_[36409]_ ,
    \new_[36413]_ , \new_[36414]_ , \new_[36415]_ , \new_[36419]_ ,
    \new_[36420]_ , \new_[36424]_ , \new_[36425]_ , \new_[36426]_ ,
    \new_[36430]_ , \new_[36431]_ , \new_[36435]_ , \new_[36436]_ ,
    \new_[36437]_ , \new_[36441]_ , \new_[36442]_ , \new_[36446]_ ,
    \new_[36447]_ , \new_[36448]_ , \new_[36452]_ , \new_[36453]_ ,
    \new_[36457]_ , \new_[36458]_ , \new_[36459]_ , \new_[36463]_ ,
    \new_[36464]_ , \new_[36468]_ , \new_[36469]_ , \new_[36470]_ ,
    \new_[36474]_ , \new_[36475]_ , \new_[36479]_ , \new_[36480]_ ,
    \new_[36481]_ , \new_[36485]_ , \new_[36486]_ , \new_[36490]_ ,
    \new_[36491]_ , \new_[36492]_ , \new_[36496]_ , \new_[36497]_ ,
    \new_[36501]_ , \new_[36502]_ , \new_[36503]_ , \new_[36507]_ ,
    \new_[36508]_ , \new_[36512]_ , \new_[36513]_ , \new_[36514]_ ,
    \new_[36518]_ , \new_[36519]_ , \new_[36523]_ , \new_[36524]_ ,
    \new_[36525]_ , \new_[36529]_ , \new_[36530]_ , \new_[36534]_ ,
    \new_[36535]_ , \new_[36536]_ , \new_[36540]_ , \new_[36541]_ ,
    \new_[36545]_ , \new_[36546]_ , \new_[36547]_ , \new_[36551]_ ,
    \new_[36552]_ , \new_[36556]_ , \new_[36557]_ , \new_[36558]_ ,
    \new_[36562]_ , \new_[36563]_ , \new_[36567]_ , \new_[36568]_ ,
    \new_[36569]_ , \new_[36573]_ , \new_[36574]_ , \new_[36578]_ ,
    \new_[36579]_ , \new_[36580]_ , \new_[36584]_ , \new_[36585]_ ,
    \new_[36589]_ , \new_[36590]_ , \new_[36591]_ , \new_[36595]_ ,
    \new_[36596]_ , \new_[36600]_ , \new_[36601]_ , \new_[36602]_ ,
    \new_[36606]_ , \new_[36607]_ , \new_[36611]_ , \new_[36612]_ ,
    \new_[36613]_ , \new_[36617]_ , \new_[36618]_ , \new_[36622]_ ,
    \new_[36623]_ , \new_[36624]_ , \new_[36628]_ , \new_[36629]_ ,
    \new_[36633]_ , \new_[36634]_ , \new_[36635]_ , \new_[36639]_ ,
    \new_[36640]_ , \new_[36644]_ , \new_[36645]_ , \new_[36646]_ ,
    \new_[36650]_ , \new_[36651]_ , \new_[36655]_ , \new_[36656]_ ,
    \new_[36657]_ , \new_[36661]_ , \new_[36662]_ , \new_[36666]_ ,
    \new_[36667]_ , \new_[36668]_ , \new_[36672]_ , \new_[36673]_ ,
    \new_[36677]_ , \new_[36678]_ , \new_[36679]_ , \new_[36683]_ ,
    \new_[36684]_ , \new_[36688]_ , \new_[36689]_ , \new_[36690]_ ,
    \new_[36694]_ , \new_[36695]_ , \new_[36699]_ , \new_[36700]_ ,
    \new_[36701]_ , \new_[36705]_ , \new_[36706]_ , \new_[36710]_ ,
    \new_[36711]_ , \new_[36712]_ , \new_[36716]_ , \new_[36717]_ ,
    \new_[36721]_ , \new_[36722]_ , \new_[36723]_ , \new_[36727]_ ,
    \new_[36728]_ , \new_[36732]_ , \new_[36733]_ , \new_[36734]_ ,
    \new_[36738]_ , \new_[36739]_ , \new_[36743]_ , \new_[36744]_ ,
    \new_[36745]_ , \new_[36749]_ , \new_[36750]_ , \new_[36754]_ ,
    \new_[36755]_ , \new_[36756]_ , \new_[36760]_ , \new_[36761]_ ,
    \new_[36765]_ , \new_[36766]_ , \new_[36767]_ , \new_[36771]_ ,
    \new_[36772]_ , \new_[36776]_ , \new_[36777]_ , \new_[36778]_ ,
    \new_[36782]_ , \new_[36783]_ , \new_[36787]_ , \new_[36788]_ ,
    \new_[36789]_ , \new_[36793]_ , \new_[36794]_ , \new_[36798]_ ,
    \new_[36799]_ , \new_[36800]_ , \new_[36804]_ , \new_[36805]_ ,
    \new_[36809]_ , \new_[36810]_ , \new_[36811]_ , \new_[36815]_ ,
    \new_[36816]_ , \new_[36820]_ , \new_[36821]_ , \new_[36822]_ ,
    \new_[36826]_ , \new_[36827]_ , \new_[36831]_ , \new_[36832]_ ,
    \new_[36833]_ , \new_[36837]_ , \new_[36838]_ , \new_[36842]_ ,
    \new_[36843]_ , \new_[36844]_ , \new_[36848]_ , \new_[36849]_ ,
    \new_[36853]_ , \new_[36854]_ , \new_[36855]_ , \new_[36859]_ ,
    \new_[36860]_ , \new_[36864]_ , \new_[36865]_ , \new_[36866]_ ,
    \new_[36870]_ , \new_[36871]_ , \new_[36875]_ , \new_[36876]_ ,
    \new_[36877]_ , \new_[36881]_ , \new_[36882]_ , \new_[36886]_ ,
    \new_[36887]_ , \new_[36888]_ , \new_[36892]_ , \new_[36893]_ ,
    \new_[36897]_ , \new_[36898]_ , \new_[36899]_ , \new_[36903]_ ,
    \new_[36904]_ , \new_[36908]_ , \new_[36909]_ , \new_[36910]_ ,
    \new_[36914]_ , \new_[36915]_ , \new_[36919]_ , \new_[36920]_ ,
    \new_[36921]_ , \new_[36925]_ , \new_[36926]_ , \new_[36930]_ ,
    \new_[36931]_ , \new_[36932]_ , \new_[36936]_ , \new_[36937]_ ,
    \new_[36941]_ , \new_[36942]_ , \new_[36943]_ , \new_[36947]_ ,
    \new_[36948]_ , \new_[36952]_ , \new_[36953]_ , \new_[36954]_ ,
    \new_[36958]_ , \new_[36959]_ , \new_[36963]_ , \new_[36964]_ ,
    \new_[36965]_ , \new_[36969]_ , \new_[36970]_ , \new_[36974]_ ,
    \new_[36975]_ , \new_[36976]_ , \new_[36980]_ , \new_[36981]_ ,
    \new_[36985]_ , \new_[36986]_ , \new_[36987]_ , \new_[36991]_ ,
    \new_[36992]_ , \new_[36996]_ , \new_[36997]_ , \new_[36998]_ ,
    \new_[37002]_ , \new_[37003]_ , \new_[37007]_ , \new_[37008]_ ,
    \new_[37009]_ , \new_[37013]_ , \new_[37014]_ , \new_[37018]_ ,
    \new_[37019]_ , \new_[37020]_ , \new_[37024]_ , \new_[37025]_ ,
    \new_[37029]_ , \new_[37030]_ , \new_[37031]_ , \new_[37035]_ ,
    \new_[37036]_ , \new_[37040]_ , \new_[37041]_ , \new_[37042]_ ,
    \new_[37046]_ , \new_[37047]_ , \new_[37051]_ , \new_[37052]_ ,
    \new_[37053]_ , \new_[37057]_ , \new_[37058]_ , \new_[37062]_ ,
    \new_[37063]_ , \new_[37064]_ , \new_[37068]_ , \new_[37069]_ ,
    \new_[37073]_ , \new_[37074]_ , \new_[37075]_ , \new_[37079]_ ,
    \new_[37080]_ , \new_[37084]_ , \new_[37085]_ , \new_[37086]_ ,
    \new_[37090]_ , \new_[37091]_ , \new_[37095]_ , \new_[37096]_ ,
    \new_[37097]_ , \new_[37101]_ , \new_[37102]_ , \new_[37106]_ ,
    \new_[37107]_ , \new_[37108]_ , \new_[37112]_ , \new_[37113]_ ,
    \new_[37117]_ , \new_[37118]_ , \new_[37119]_ , \new_[37123]_ ,
    \new_[37124]_ , \new_[37128]_ , \new_[37129]_ , \new_[37130]_ ,
    \new_[37134]_ , \new_[37135]_ , \new_[37139]_ , \new_[37140]_ ,
    \new_[37141]_ , \new_[37145]_ , \new_[37146]_ , \new_[37150]_ ,
    \new_[37151]_ , \new_[37152]_ , \new_[37156]_ , \new_[37157]_ ,
    \new_[37161]_ , \new_[37162]_ , \new_[37163]_ , \new_[37167]_ ,
    \new_[37168]_ , \new_[37172]_ , \new_[37173]_ , \new_[37174]_ ,
    \new_[37178]_ , \new_[37179]_ , \new_[37183]_ , \new_[37184]_ ,
    \new_[37185]_ , \new_[37189]_ , \new_[37190]_ , \new_[37194]_ ,
    \new_[37195]_ , \new_[37196]_ , \new_[37200]_ , \new_[37201]_ ,
    \new_[37205]_ , \new_[37206]_ , \new_[37207]_ , \new_[37211]_ ,
    \new_[37212]_ , \new_[37216]_ , \new_[37217]_ , \new_[37218]_ ,
    \new_[37222]_ , \new_[37223]_ , \new_[37227]_ , \new_[37228]_ ,
    \new_[37229]_ , \new_[37233]_ , \new_[37234]_ , \new_[37238]_ ,
    \new_[37239]_ , \new_[37240]_ , \new_[37244]_ , \new_[37245]_ ,
    \new_[37249]_ , \new_[37250]_ , \new_[37251]_ , \new_[37255]_ ,
    \new_[37256]_ , \new_[37260]_ , \new_[37261]_ , \new_[37262]_ ,
    \new_[37266]_ , \new_[37267]_ , \new_[37271]_ , \new_[37272]_ ,
    \new_[37273]_ , \new_[37277]_ , \new_[37278]_ , \new_[37282]_ ,
    \new_[37283]_ , \new_[37284]_ , \new_[37288]_ , \new_[37289]_ ,
    \new_[37293]_ , \new_[37294]_ , \new_[37295]_ , \new_[37299]_ ,
    \new_[37300]_ , \new_[37304]_ , \new_[37305]_ , \new_[37306]_ ,
    \new_[37310]_ , \new_[37311]_ , \new_[37315]_ , \new_[37316]_ ,
    \new_[37317]_ , \new_[37321]_ , \new_[37322]_ , \new_[37326]_ ,
    \new_[37327]_ , \new_[37328]_ , \new_[37332]_ , \new_[37333]_ ,
    \new_[37337]_ , \new_[37338]_ , \new_[37339]_ , \new_[37343]_ ,
    \new_[37344]_ , \new_[37348]_ , \new_[37349]_ , \new_[37350]_ ,
    \new_[37354]_ , \new_[37355]_ , \new_[37359]_ , \new_[37360]_ ,
    \new_[37361]_ , \new_[37365]_ , \new_[37366]_ , \new_[37370]_ ,
    \new_[37371]_ , \new_[37372]_ , \new_[37376]_ , \new_[37377]_ ,
    \new_[37381]_ , \new_[37382]_ , \new_[37383]_ , \new_[37387]_ ,
    \new_[37388]_ , \new_[37392]_ , \new_[37393]_ , \new_[37394]_ ,
    \new_[37398]_ , \new_[37399]_ , \new_[37403]_ , \new_[37404]_ ,
    \new_[37405]_ , \new_[37409]_ , \new_[37410]_ , \new_[37414]_ ,
    \new_[37415]_ , \new_[37416]_ , \new_[37420]_ , \new_[37421]_ ,
    \new_[37425]_ , \new_[37426]_ , \new_[37427]_ , \new_[37431]_ ,
    \new_[37432]_ , \new_[37436]_ , \new_[37437]_ , \new_[37438]_ ,
    \new_[37442]_ , \new_[37443]_ , \new_[37447]_ , \new_[37448]_ ,
    \new_[37449]_ , \new_[37453]_ , \new_[37454]_ , \new_[37458]_ ,
    \new_[37459]_ , \new_[37460]_ , \new_[37464]_ , \new_[37465]_ ,
    \new_[37469]_ , \new_[37470]_ , \new_[37471]_ , \new_[37475]_ ,
    \new_[37476]_ , \new_[37480]_ , \new_[37481]_ , \new_[37482]_ ,
    \new_[37486]_ , \new_[37487]_ , \new_[37491]_ , \new_[37492]_ ,
    \new_[37493]_ , \new_[37497]_ , \new_[37498]_ , \new_[37502]_ ,
    \new_[37503]_ , \new_[37504]_ , \new_[37508]_ , \new_[37509]_ ,
    \new_[37513]_ , \new_[37514]_ , \new_[37515]_ , \new_[37519]_ ,
    \new_[37520]_ , \new_[37524]_ , \new_[37525]_ , \new_[37526]_ ,
    \new_[37530]_ , \new_[37531]_ , \new_[37535]_ , \new_[37536]_ ,
    \new_[37537]_ , \new_[37541]_ , \new_[37542]_ , \new_[37546]_ ,
    \new_[37547]_ , \new_[37548]_ , \new_[37552]_ , \new_[37553]_ ,
    \new_[37557]_ , \new_[37558]_ , \new_[37559]_ , \new_[37563]_ ,
    \new_[37564]_ , \new_[37568]_ , \new_[37569]_ , \new_[37570]_ ,
    \new_[37574]_ , \new_[37575]_ , \new_[37579]_ , \new_[37580]_ ,
    \new_[37581]_ , \new_[37585]_ , \new_[37586]_ , \new_[37590]_ ,
    \new_[37591]_ , \new_[37592]_ , \new_[37596]_ , \new_[37597]_ ,
    \new_[37601]_ , \new_[37602]_ , \new_[37603]_ , \new_[37607]_ ,
    \new_[37608]_ , \new_[37612]_ , \new_[37613]_ , \new_[37614]_ ,
    \new_[37618]_ , \new_[37619]_ , \new_[37623]_ , \new_[37624]_ ,
    \new_[37625]_ , \new_[37629]_ , \new_[37630]_ , \new_[37634]_ ,
    \new_[37635]_ , \new_[37636]_ , \new_[37640]_ , \new_[37641]_ ,
    \new_[37645]_ , \new_[37646]_ , \new_[37647]_ , \new_[37651]_ ,
    \new_[37652]_ , \new_[37656]_ , \new_[37657]_ , \new_[37658]_ ,
    \new_[37662]_ , \new_[37663]_ , \new_[37667]_ , \new_[37668]_ ,
    \new_[37669]_ , \new_[37673]_ , \new_[37674]_ , \new_[37678]_ ,
    \new_[37679]_ , \new_[37680]_ , \new_[37684]_ , \new_[37685]_ ,
    \new_[37689]_ , \new_[37690]_ , \new_[37691]_ , \new_[37695]_ ,
    \new_[37696]_ , \new_[37700]_ , \new_[37701]_ , \new_[37702]_ ,
    \new_[37706]_ , \new_[37707]_ , \new_[37711]_ , \new_[37712]_ ,
    \new_[37713]_ , \new_[37717]_ , \new_[37718]_ , \new_[37722]_ ,
    \new_[37723]_ , \new_[37724]_ , \new_[37728]_ , \new_[37729]_ ,
    \new_[37733]_ , \new_[37734]_ , \new_[37735]_ , \new_[37739]_ ,
    \new_[37740]_ , \new_[37744]_ , \new_[37745]_ , \new_[37746]_ ,
    \new_[37750]_ , \new_[37751]_ , \new_[37755]_ , \new_[37756]_ ,
    \new_[37757]_ , \new_[37761]_ , \new_[37762]_ , \new_[37766]_ ,
    \new_[37767]_ , \new_[37768]_ , \new_[37772]_ , \new_[37773]_ ,
    \new_[37777]_ , \new_[37778]_ , \new_[37779]_ , \new_[37783]_ ,
    \new_[37784]_ , \new_[37788]_ , \new_[37789]_ , \new_[37790]_ ,
    \new_[37794]_ , \new_[37795]_ , \new_[37799]_ , \new_[37800]_ ,
    \new_[37801]_ , \new_[37805]_ , \new_[37806]_ , \new_[37810]_ ,
    \new_[37811]_ , \new_[37812]_ , \new_[37816]_ , \new_[37817]_ ,
    \new_[37821]_ , \new_[37822]_ , \new_[37823]_ , \new_[37827]_ ,
    \new_[37828]_ , \new_[37832]_ , \new_[37833]_ , \new_[37834]_ ,
    \new_[37838]_ , \new_[37839]_ , \new_[37843]_ , \new_[37844]_ ,
    \new_[37845]_ , \new_[37849]_ , \new_[37850]_ , \new_[37854]_ ,
    \new_[37855]_ , \new_[37856]_ , \new_[37860]_ , \new_[37861]_ ,
    \new_[37865]_ , \new_[37866]_ , \new_[37867]_ , \new_[37871]_ ,
    \new_[37872]_ , \new_[37876]_ , \new_[37877]_ , \new_[37878]_ ,
    \new_[37882]_ , \new_[37883]_ , \new_[37887]_ , \new_[37888]_ ,
    \new_[37889]_ , \new_[37893]_ , \new_[37894]_ , \new_[37898]_ ,
    \new_[37899]_ , \new_[37900]_ , \new_[37904]_ , \new_[37905]_ ,
    \new_[37909]_ , \new_[37910]_ , \new_[37911]_ , \new_[37915]_ ,
    \new_[37916]_ , \new_[37920]_ , \new_[37921]_ , \new_[37922]_ ,
    \new_[37926]_ , \new_[37927]_ , \new_[37931]_ , \new_[37932]_ ,
    \new_[37933]_ , \new_[37937]_ , \new_[37938]_ , \new_[37942]_ ,
    \new_[37943]_ , \new_[37944]_ , \new_[37948]_ , \new_[37949]_ ,
    \new_[37953]_ , \new_[37954]_ , \new_[37955]_ , \new_[37959]_ ,
    \new_[37960]_ , \new_[37964]_ , \new_[37965]_ , \new_[37966]_ ,
    \new_[37970]_ , \new_[37971]_ , \new_[37975]_ , \new_[37976]_ ,
    \new_[37977]_ , \new_[37981]_ , \new_[37982]_ , \new_[37986]_ ,
    \new_[37987]_ , \new_[37988]_ , \new_[37992]_ , \new_[37993]_ ,
    \new_[37997]_ , \new_[37998]_ , \new_[37999]_ , \new_[38003]_ ,
    \new_[38004]_ , \new_[38008]_ , \new_[38009]_ , \new_[38010]_ ,
    \new_[38014]_ , \new_[38015]_ , \new_[38019]_ , \new_[38020]_ ,
    \new_[38021]_ , \new_[38025]_ , \new_[38026]_ , \new_[38030]_ ,
    \new_[38031]_ , \new_[38032]_ , \new_[38036]_ , \new_[38037]_ ,
    \new_[38041]_ , \new_[38042]_ , \new_[38043]_ , \new_[38047]_ ,
    \new_[38048]_ , \new_[38052]_ , \new_[38053]_ , \new_[38054]_ ,
    \new_[38058]_ , \new_[38059]_ , \new_[38063]_ , \new_[38064]_ ,
    \new_[38065]_ , \new_[38069]_ , \new_[38070]_ , \new_[38074]_ ,
    \new_[38075]_ , \new_[38076]_ , \new_[38080]_ , \new_[38081]_ ,
    \new_[38085]_ , \new_[38086]_ , \new_[38087]_ , \new_[38091]_ ,
    \new_[38092]_ , \new_[38096]_ , \new_[38097]_ , \new_[38098]_ ,
    \new_[38102]_ , \new_[38103]_ , \new_[38107]_ , \new_[38108]_ ,
    \new_[38109]_ , \new_[38113]_ , \new_[38114]_ , \new_[38118]_ ,
    \new_[38119]_ , \new_[38120]_ , \new_[38124]_ , \new_[38125]_ ,
    \new_[38129]_ , \new_[38130]_ , \new_[38131]_ , \new_[38135]_ ,
    \new_[38136]_ , \new_[38140]_ , \new_[38141]_ , \new_[38142]_ ,
    \new_[38146]_ , \new_[38147]_ , \new_[38151]_ , \new_[38152]_ ,
    \new_[38153]_ , \new_[38157]_ , \new_[38158]_ , \new_[38162]_ ,
    \new_[38163]_ , \new_[38164]_ , \new_[38168]_ , \new_[38169]_ ,
    \new_[38173]_ , \new_[38174]_ , \new_[38175]_ , \new_[38179]_ ,
    \new_[38180]_ , \new_[38184]_ , \new_[38185]_ , \new_[38186]_ ,
    \new_[38190]_ , \new_[38191]_ , \new_[38195]_ , \new_[38196]_ ,
    \new_[38197]_ , \new_[38201]_ , \new_[38202]_ , \new_[38206]_ ,
    \new_[38207]_ , \new_[38208]_ , \new_[38212]_ , \new_[38213]_ ,
    \new_[38217]_ , \new_[38218]_ , \new_[38219]_ , \new_[38223]_ ,
    \new_[38224]_ , \new_[38228]_ , \new_[38229]_ , \new_[38230]_ ,
    \new_[38234]_ , \new_[38235]_ , \new_[38239]_ , \new_[38240]_ ,
    \new_[38241]_ , \new_[38245]_ , \new_[38246]_ , \new_[38250]_ ,
    \new_[38251]_ , \new_[38252]_ , \new_[38256]_ , \new_[38257]_ ,
    \new_[38261]_ , \new_[38262]_ , \new_[38263]_ , \new_[38267]_ ,
    \new_[38268]_ , \new_[38272]_ , \new_[38273]_ , \new_[38274]_ ,
    \new_[38278]_ , \new_[38279]_ , \new_[38283]_ , \new_[38284]_ ,
    \new_[38285]_ , \new_[38289]_ , \new_[38290]_ , \new_[38294]_ ,
    \new_[38295]_ , \new_[38296]_ , \new_[38300]_ , \new_[38301]_ ,
    \new_[38305]_ , \new_[38306]_ , \new_[38307]_ , \new_[38311]_ ,
    \new_[38312]_ , \new_[38316]_ , \new_[38317]_ , \new_[38318]_ ,
    \new_[38322]_ , \new_[38323]_ , \new_[38327]_ , \new_[38328]_ ,
    \new_[38329]_ , \new_[38333]_ , \new_[38334]_ , \new_[38338]_ ,
    \new_[38339]_ , \new_[38340]_ , \new_[38344]_ , \new_[38345]_ ,
    \new_[38349]_ , \new_[38350]_ , \new_[38351]_ , \new_[38355]_ ,
    \new_[38356]_ , \new_[38360]_ , \new_[38361]_ , \new_[38362]_ ,
    \new_[38366]_ , \new_[38367]_ , \new_[38371]_ , \new_[38372]_ ,
    \new_[38373]_ , \new_[38377]_ , \new_[38378]_ , \new_[38382]_ ,
    \new_[38383]_ , \new_[38384]_ , \new_[38388]_ , \new_[38389]_ ,
    \new_[38393]_ , \new_[38394]_ , \new_[38395]_ , \new_[38399]_ ,
    \new_[38400]_ , \new_[38404]_ , \new_[38405]_ , \new_[38406]_ ,
    \new_[38410]_ , \new_[38411]_ , \new_[38415]_ , \new_[38416]_ ,
    \new_[38417]_ , \new_[38421]_ , \new_[38422]_ , \new_[38426]_ ,
    \new_[38427]_ , \new_[38428]_ , \new_[38432]_ , \new_[38433]_ ,
    \new_[38437]_ , \new_[38438]_ , \new_[38439]_ , \new_[38443]_ ,
    \new_[38444]_ , \new_[38448]_ , \new_[38449]_ , \new_[38450]_ ,
    \new_[38454]_ , \new_[38455]_ , \new_[38459]_ , \new_[38460]_ ,
    \new_[38461]_ , \new_[38465]_ , \new_[38466]_ , \new_[38470]_ ,
    \new_[38471]_ , \new_[38472]_ , \new_[38476]_ , \new_[38477]_ ,
    \new_[38481]_ , \new_[38482]_ , \new_[38483]_ , \new_[38487]_ ,
    \new_[38488]_ , \new_[38492]_ , \new_[38493]_ , \new_[38494]_ ,
    \new_[38498]_ , \new_[38499]_ , \new_[38503]_ , \new_[38504]_ ,
    \new_[38505]_ , \new_[38509]_ , \new_[38510]_ , \new_[38514]_ ,
    \new_[38515]_ , \new_[38516]_ , \new_[38520]_ , \new_[38521]_ ,
    \new_[38525]_ , \new_[38526]_ , \new_[38527]_ , \new_[38531]_ ,
    \new_[38532]_ , \new_[38536]_ , \new_[38537]_ , \new_[38538]_ ,
    \new_[38542]_ , \new_[38543]_ , \new_[38547]_ , \new_[38548]_ ,
    \new_[38549]_ , \new_[38553]_ , \new_[38554]_ , \new_[38558]_ ,
    \new_[38559]_ , \new_[38560]_ , \new_[38564]_ , \new_[38565]_ ,
    \new_[38569]_ , \new_[38570]_ , \new_[38571]_ , \new_[38575]_ ,
    \new_[38576]_ , \new_[38580]_ , \new_[38581]_ , \new_[38582]_ ,
    \new_[38586]_ , \new_[38587]_ , \new_[38591]_ , \new_[38592]_ ,
    \new_[38593]_ , \new_[38597]_ , \new_[38598]_ , \new_[38602]_ ,
    \new_[38603]_ , \new_[38604]_ , \new_[38608]_ , \new_[38609]_ ,
    \new_[38613]_ , \new_[38614]_ , \new_[38615]_ , \new_[38619]_ ,
    \new_[38620]_ , \new_[38624]_ , \new_[38625]_ , \new_[38626]_ ,
    \new_[38630]_ , \new_[38631]_ , \new_[38635]_ , \new_[38636]_ ,
    \new_[38637]_ , \new_[38641]_ , \new_[38642]_ , \new_[38646]_ ,
    \new_[38647]_ , \new_[38648]_ , \new_[38652]_ , \new_[38653]_ ,
    \new_[38657]_ , \new_[38658]_ , \new_[38659]_ , \new_[38663]_ ,
    \new_[38664]_ , \new_[38668]_ , \new_[38669]_ , \new_[38670]_ ,
    \new_[38674]_ , \new_[38675]_ , \new_[38679]_ , \new_[38680]_ ,
    \new_[38681]_ , \new_[38685]_ , \new_[38686]_ , \new_[38690]_ ,
    \new_[38691]_ , \new_[38692]_ , \new_[38696]_ , \new_[38697]_ ,
    \new_[38701]_ , \new_[38702]_ , \new_[38703]_ , \new_[38707]_ ,
    \new_[38708]_ , \new_[38712]_ , \new_[38713]_ , \new_[38714]_ ,
    \new_[38718]_ , \new_[38719]_ , \new_[38723]_ , \new_[38724]_ ,
    \new_[38725]_ , \new_[38729]_ , \new_[38730]_ , \new_[38734]_ ,
    \new_[38735]_ , \new_[38736]_ , \new_[38740]_ , \new_[38741]_ ,
    \new_[38745]_ , \new_[38746]_ , \new_[38747]_ , \new_[38751]_ ,
    \new_[38752]_ , \new_[38756]_ , \new_[38757]_ , \new_[38758]_ ,
    \new_[38762]_ , \new_[38763]_ , \new_[38767]_ , \new_[38768]_ ,
    \new_[38769]_ , \new_[38773]_ , \new_[38774]_ , \new_[38778]_ ,
    \new_[38779]_ , \new_[38780]_ , \new_[38784]_ , \new_[38785]_ ,
    \new_[38789]_ , \new_[38790]_ , \new_[38791]_ , \new_[38795]_ ,
    \new_[38796]_ , \new_[38800]_ , \new_[38801]_ , \new_[38802]_ ,
    \new_[38806]_ , \new_[38807]_ , \new_[38811]_ , \new_[38812]_ ,
    \new_[38813]_ , \new_[38817]_ , \new_[38818]_ , \new_[38822]_ ,
    \new_[38823]_ , \new_[38824]_ , \new_[38828]_ , \new_[38829]_ ,
    \new_[38833]_ , \new_[38834]_ , \new_[38835]_ , \new_[38839]_ ,
    \new_[38840]_ , \new_[38844]_ , \new_[38845]_ , \new_[38846]_ ,
    \new_[38850]_ , \new_[38851]_ , \new_[38855]_ , \new_[38856]_ ,
    \new_[38857]_ , \new_[38861]_ , \new_[38862]_ , \new_[38866]_ ,
    \new_[38867]_ , \new_[38868]_ , \new_[38872]_ , \new_[38873]_ ,
    \new_[38877]_ , \new_[38878]_ , \new_[38879]_ , \new_[38883]_ ,
    \new_[38884]_ , \new_[38888]_ , \new_[38889]_ , \new_[38890]_ ,
    \new_[38894]_ , \new_[38895]_ , \new_[38899]_ , \new_[38900]_ ,
    \new_[38901]_ , \new_[38905]_ , \new_[38906]_ , \new_[38910]_ ,
    \new_[38911]_ , \new_[38912]_ , \new_[38916]_ , \new_[38917]_ ,
    \new_[38921]_ , \new_[38922]_ , \new_[38923]_ , \new_[38927]_ ,
    \new_[38928]_ , \new_[38932]_ , \new_[38933]_ , \new_[38934]_ ,
    \new_[38938]_ , \new_[38939]_ , \new_[38943]_ , \new_[38944]_ ,
    \new_[38945]_ , \new_[38949]_ , \new_[38950]_ , \new_[38954]_ ,
    \new_[38955]_ , \new_[38956]_ , \new_[38960]_ , \new_[38961]_ ,
    \new_[38965]_ , \new_[38966]_ , \new_[38967]_ , \new_[38971]_ ,
    \new_[38972]_ , \new_[38976]_ , \new_[38977]_ , \new_[38978]_ ,
    \new_[38982]_ , \new_[38983]_ , \new_[38987]_ , \new_[38988]_ ,
    \new_[38989]_ , \new_[38993]_ , \new_[38994]_ , \new_[38998]_ ,
    \new_[38999]_ , \new_[39000]_ , \new_[39004]_ , \new_[39005]_ ,
    \new_[39009]_ , \new_[39010]_ , \new_[39011]_ , \new_[39015]_ ,
    \new_[39016]_ , \new_[39020]_ , \new_[39021]_ , \new_[39022]_ ,
    \new_[39026]_ , \new_[39027]_ , \new_[39031]_ , \new_[39032]_ ,
    \new_[39033]_ , \new_[39037]_ , \new_[39038]_ , \new_[39042]_ ,
    \new_[39043]_ , \new_[39044]_ , \new_[39048]_ , \new_[39049]_ ,
    \new_[39053]_ , \new_[39054]_ , \new_[39055]_ , \new_[39059]_ ,
    \new_[39060]_ , \new_[39064]_ , \new_[39065]_ , \new_[39066]_ ,
    \new_[39070]_ , \new_[39071]_ , \new_[39075]_ , \new_[39076]_ ,
    \new_[39077]_ , \new_[39081]_ , \new_[39082]_ , \new_[39086]_ ,
    \new_[39087]_ , \new_[39088]_ , \new_[39092]_ , \new_[39093]_ ,
    \new_[39097]_ , \new_[39098]_ , \new_[39099]_ , \new_[39103]_ ,
    \new_[39104]_ , \new_[39108]_ , \new_[39109]_ , \new_[39110]_ ,
    \new_[39114]_ , \new_[39115]_ , \new_[39119]_ , \new_[39120]_ ,
    \new_[39121]_ , \new_[39125]_ , \new_[39126]_ , \new_[39130]_ ,
    \new_[39131]_ , \new_[39132]_ , \new_[39136]_ , \new_[39137]_ ,
    \new_[39141]_ , \new_[39142]_ , \new_[39143]_ , \new_[39147]_ ,
    \new_[39148]_ , \new_[39152]_ , \new_[39153]_ , \new_[39154]_ ,
    \new_[39158]_ , \new_[39159]_ , \new_[39163]_ , \new_[39164]_ ,
    \new_[39165]_ , \new_[39169]_ , \new_[39170]_ , \new_[39174]_ ,
    \new_[39175]_ , \new_[39176]_ , \new_[39180]_ , \new_[39181]_ ,
    \new_[39185]_ , \new_[39186]_ , \new_[39187]_ , \new_[39191]_ ,
    \new_[39192]_ , \new_[39196]_ , \new_[39197]_ , \new_[39198]_ ,
    \new_[39202]_ , \new_[39203]_ , \new_[39207]_ , \new_[39208]_ ,
    \new_[39209]_ , \new_[39213]_ , \new_[39214]_ , \new_[39218]_ ,
    \new_[39219]_ , \new_[39220]_ , \new_[39224]_ , \new_[39225]_ ,
    \new_[39229]_ , \new_[39230]_ , \new_[39231]_ , \new_[39235]_ ,
    \new_[39236]_ , \new_[39240]_ , \new_[39241]_ , \new_[39242]_ ,
    \new_[39246]_ , \new_[39247]_ , \new_[39251]_ , \new_[39252]_ ,
    \new_[39253]_ , \new_[39257]_ , \new_[39258]_ , \new_[39262]_ ,
    \new_[39263]_ , \new_[39264]_ , \new_[39268]_ , \new_[39269]_ ,
    \new_[39273]_ , \new_[39274]_ , \new_[39275]_ , \new_[39279]_ ,
    \new_[39280]_ , \new_[39284]_ , \new_[39285]_ , \new_[39286]_ ,
    \new_[39290]_ , \new_[39291]_ , \new_[39295]_ , \new_[39296]_ ,
    \new_[39297]_ , \new_[39301]_ , \new_[39302]_ , \new_[39306]_ ,
    \new_[39307]_ , \new_[39308]_ , \new_[39312]_ , \new_[39313]_ ,
    \new_[39317]_ , \new_[39318]_ , \new_[39319]_ , \new_[39323]_ ,
    \new_[39324]_ , \new_[39328]_ , \new_[39329]_ , \new_[39330]_ ,
    \new_[39334]_ , \new_[39335]_ , \new_[39339]_ , \new_[39340]_ ,
    \new_[39341]_ , \new_[39345]_ , \new_[39346]_ , \new_[39350]_ ,
    \new_[39351]_ , \new_[39352]_ , \new_[39356]_ , \new_[39357]_ ,
    \new_[39361]_ , \new_[39362]_ , \new_[39363]_ , \new_[39367]_ ,
    \new_[39368]_ , \new_[39372]_ , \new_[39373]_ , \new_[39374]_ ,
    \new_[39378]_ , \new_[39379]_ , \new_[39383]_ , \new_[39384]_ ,
    \new_[39385]_ , \new_[39389]_ , \new_[39390]_ , \new_[39394]_ ,
    \new_[39395]_ , \new_[39396]_ , \new_[39400]_ , \new_[39401]_ ,
    \new_[39405]_ , \new_[39406]_ , \new_[39407]_ , \new_[39411]_ ,
    \new_[39412]_ , \new_[39416]_ , \new_[39417]_ , \new_[39418]_ ,
    \new_[39422]_ , \new_[39423]_ , \new_[39427]_ , \new_[39428]_ ,
    \new_[39429]_ , \new_[39433]_ , \new_[39434]_ , \new_[39438]_ ,
    \new_[39439]_ , \new_[39440]_ , \new_[39444]_ , \new_[39445]_ ,
    \new_[39449]_ , \new_[39450]_ , \new_[39451]_ , \new_[39455]_ ,
    \new_[39456]_ , \new_[39460]_ , \new_[39461]_ , \new_[39462]_ ,
    \new_[39466]_ , \new_[39467]_ , \new_[39471]_ , \new_[39472]_ ,
    \new_[39473]_ , \new_[39477]_ , \new_[39478]_ , \new_[39482]_ ,
    \new_[39483]_ , \new_[39484]_ , \new_[39488]_ , \new_[39489]_ ,
    \new_[39493]_ , \new_[39494]_ , \new_[39495]_ , \new_[39499]_ ,
    \new_[39500]_ , \new_[39504]_ , \new_[39505]_ , \new_[39506]_ ,
    \new_[39510]_ , \new_[39511]_ , \new_[39515]_ , \new_[39516]_ ,
    \new_[39517]_ , \new_[39521]_ , \new_[39522]_ , \new_[39526]_ ,
    \new_[39527]_ , \new_[39528]_ , \new_[39532]_ , \new_[39533]_ ,
    \new_[39537]_ , \new_[39538]_ , \new_[39539]_ , \new_[39543]_ ,
    \new_[39544]_ , \new_[39548]_ , \new_[39549]_ , \new_[39550]_ ,
    \new_[39554]_ , \new_[39555]_ , \new_[39559]_ , \new_[39560]_ ,
    \new_[39561]_ , \new_[39565]_ , \new_[39566]_ , \new_[39570]_ ,
    \new_[39571]_ , \new_[39572]_ , \new_[39576]_ , \new_[39577]_ ,
    \new_[39581]_ , \new_[39582]_ , \new_[39583]_ , \new_[39587]_ ,
    \new_[39588]_ , \new_[39592]_ , \new_[39593]_ , \new_[39594]_ ,
    \new_[39598]_ , \new_[39599]_ , \new_[39603]_ , \new_[39604]_ ,
    \new_[39605]_ , \new_[39609]_ , \new_[39610]_ , \new_[39614]_ ,
    \new_[39615]_ , \new_[39616]_ , \new_[39620]_ , \new_[39621]_ ,
    \new_[39625]_ , \new_[39626]_ , \new_[39627]_ , \new_[39631]_ ,
    \new_[39632]_ , \new_[39636]_ , \new_[39637]_ , \new_[39638]_ ,
    \new_[39642]_ , \new_[39643]_ , \new_[39647]_ , \new_[39648]_ ,
    \new_[39649]_ , \new_[39653]_ , \new_[39654]_ , \new_[39658]_ ,
    \new_[39659]_ , \new_[39660]_ , \new_[39664]_ , \new_[39665]_ ,
    \new_[39669]_ , \new_[39670]_ , \new_[39671]_ , \new_[39675]_ ,
    \new_[39676]_ , \new_[39680]_ , \new_[39681]_ , \new_[39682]_ ,
    \new_[39686]_ , \new_[39687]_ , \new_[39691]_ , \new_[39692]_ ,
    \new_[39693]_ , \new_[39697]_ , \new_[39698]_ , \new_[39702]_ ,
    \new_[39703]_ , \new_[39704]_ , \new_[39708]_ , \new_[39709]_ ,
    \new_[39713]_ , \new_[39714]_ , \new_[39715]_ , \new_[39719]_ ,
    \new_[39720]_ , \new_[39724]_ , \new_[39725]_ , \new_[39726]_ ,
    \new_[39730]_ , \new_[39731]_ , \new_[39735]_ , \new_[39736]_ ,
    \new_[39737]_ , \new_[39741]_ , \new_[39742]_ , \new_[39746]_ ,
    \new_[39747]_ , \new_[39748]_ , \new_[39752]_ , \new_[39753]_ ,
    \new_[39757]_ , \new_[39758]_ , \new_[39759]_ , \new_[39763]_ ,
    \new_[39764]_ , \new_[39768]_ , \new_[39769]_ , \new_[39770]_ ,
    \new_[39774]_ , \new_[39775]_ , \new_[39779]_ , \new_[39780]_ ,
    \new_[39781]_ , \new_[39785]_ , \new_[39786]_ , \new_[39790]_ ,
    \new_[39791]_ , \new_[39792]_ , \new_[39796]_ , \new_[39797]_ ,
    \new_[39801]_ , \new_[39802]_ , \new_[39803]_ , \new_[39807]_ ,
    \new_[39808]_ , \new_[39812]_ , \new_[39813]_ , \new_[39814]_ ,
    \new_[39818]_ , \new_[39819]_ , \new_[39823]_ , \new_[39824]_ ,
    \new_[39825]_ , \new_[39829]_ , \new_[39830]_ , \new_[39834]_ ,
    \new_[39835]_ , \new_[39836]_ , \new_[39840]_ , \new_[39841]_ ,
    \new_[39845]_ , \new_[39846]_ , \new_[39847]_ , \new_[39851]_ ,
    \new_[39852]_ , \new_[39856]_ , \new_[39857]_ , \new_[39858]_ ,
    \new_[39862]_ , \new_[39863]_ , \new_[39867]_ , \new_[39868]_ ,
    \new_[39869]_ , \new_[39873]_ , \new_[39874]_ , \new_[39878]_ ,
    \new_[39879]_ , \new_[39880]_ , \new_[39884]_ , \new_[39885]_ ,
    \new_[39889]_ , \new_[39890]_ , \new_[39891]_ , \new_[39895]_ ,
    \new_[39896]_ , \new_[39900]_ , \new_[39901]_ , \new_[39902]_ ,
    \new_[39906]_ , \new_[39907]_ , \new_[39911]_ , \new_[39912]_ ,
    \new_[39913]_ , \new_[39917]_ , \new_[39918]_ , \new_[39922]_ ,
    \new_[39923]_ , \new_[39924]_ , \new_[39928]_ , \new_[39929]_ ,
    \new_[39933]_ , \new_[39934]_ , \new_[39935]_ , \new_[39939]_ ,
    \new_[39940]_ , \new_[39944]_ , \new_[39945]_ , \new_[39946]_ ,
    \new_[39950]_ , \new_[39951]_ , \new_[39955]_ , \new_[39956]_ ,
    \new_[39957]_ , \new_[39961]_ , \new_[39962]_ , \new_[39966]_ ,
    \new_[39967]_ , \new_[39968]_ , \new_[39972]_ , \new_[39973]_ ,
    \new_[39977]_ , \new_[39978]_ , \new_[39979]_ , \new_[39983]_ ,
    \new_[39984]_ , \new_[39988]_ , \new_[39989]_ , \new_[39990]_ ,
    \new_[39994]_ , \new_[39995]_ , \new_[39999]_ , \new_[40000]_ ,
    \new_[40001]_ , \new_[40005]_ , \new_[40006]_ , \new_[40010]_ ,
    \new_[40011]_ , \new_[40012]_ , \new_[40016]_ , \new_[40017]_ ,
    \new_[40021]_ , \new_[40022]_ , \new_[40023]_ , \new_[40027]_ ,
    \new_[40028]_ , \new_[40032]_ , \new_[40033]_ , \new_[40034]_ ,
    \new_[40038]_ , \new_[40039]_ , \new_[40043]_ , \new_[40044]_ ,
    \new_[40045]_ , \new_[40049]_ , \new_[40050]_ , \new_[40054]_ ,
    \new_[40055]_ , \new_[40056]_ , \new_[40060]_ , \new_[40061]_ ,
    \new_[40065]_ , \new_[40066]_ , \new_[40067]_ , \new_[40071]_ ,
    \new_[40072]_ , \new_[40076]_ , \new_[40077]_ , \new_[40078]_ ,
    \new_[40082]_ , \new_[40083]_ , \new_[40087]_ , \new_[40088]_ ,
    \new_[40089]_ , \new_[40093]_ , \new_[40094]_ , \new_[40098]_ ,
    \new_[40099]_ , \new_[40100]_ , \new_[40104]_ , \new_[40105]_ ,
    \new_[40109]_ , \new_[40110]_ , \new_[40111]_ , \new_[40115]_ ,
    \new_[40116]_ , \new_[40120]_ , \new_[40121]_ , \new_[40122]_ ,
    \new_[40126]_ , \new_[40127]_ , \new_[40131]_ , \new_[40132]_ ,
    \new_[40133]_ , \new_[40137]_ , \new_[40138]_ , \new_[40142]_ ,
    \new_[40143]_ , \new_[40144]_ , \new_[40148]_ , \new_[40149]_ ,
    \new_[40153]_ , \new_[40154]_ , \new_[40155]_ , \new_[40159]_ ,
    \new_[40160]_ , \new_[40164]_ , \new_[40165]_ , \new_[40166]_ ,
    \new_[40170]_ , \new_[40171]_ , \new_[40175]_ , \new_[40176]_ ,
    \new_[40177]_ , \new_[40181]_ , \new_[40182]_ , \new_[40186]_ ,
    \new_[40187]_ , \new_[40188]_ , \new_[40192]_ , \new_[40193]_ ,
    \new_[40197]_ , \new_[40198]_ , \new_[40199]_ , \new_[40203]_ ,
    \new_[40204]_ , \new_[40208]_ , \new_[40209]_ , \new_[40210]_ ,
    \new_[40214]_ , \new_[40215]_ , \new_[40219]_ , \new_[40220]_ ,
    \new_[40221]_ , \new_[40225]_ , \new_[40226]_ , \new_[40230]_ ,
    \new_[40231]_ , \new_[40232]_ , \new_[40236]_ , \new_[40237]_ ,
    \new_[40241]_ , \new_[40242]_ , \new_[40243]_ , \new_[40247]_ ,
    \new_[40248]_ , \new_[40252]_ , \new_[40253]_ , \new_[40254]_ ,
    \new_[40258]_ , \new_[40259]_ , \new_[40263]_ , \new_[40264]_ ,
    \new_[40265]_ , \new_[40269]_ , \new_[40270]_ , \new_[40274]_ ,
    \new_[40275]_ , \new_[40276]_ , \new_[40280]_ , \new_[40281]_ ,
    \new_[40285]_ , \new_[40286]_ , \new_[40287]_ , \new_[40291]_ ,
    \new_[40292]_ , \new_[40296]_ , \new_[40297]_ , \new_[40298]_ ,
    \new_[40302]_ , \new_[40303]_ , \new_[40307]_ , \new_[40308]_ ,
    \new_[40309]_ , \new_[40313]_ , \new_[40314]_ , \new_[40318]_ ,
    \new_[40319]_ , \new_[40320]_ , \new_[40324]_ , \new_[40325]_ ,
    \new_[40329]_ , \new_[40330]_ , \new_[40331]_ , \new_[40335]_ ,
    \new_[40336]_ , \new_[40340]_ , \new_[40341]_ , \new_[40342]_ ,
    \new_[40346]_ , \new_[40347]_ , \new_[40351]_ , \new_[40352]_ ,
    \new_[40353]_ , \new_[40357]_ , \new_[40358]_ , \new_[40362]_ ,
    \new_[40363]_ , \new_[40364]_ , \new_[40368]_ , \new_[40369]_ ,
    \new_[40373]_ , \new_[40374]_ , \new_[40375]_ , \new_[40379]_ ,
    \new_[40380]_ , \new_[40384]_ , \new_[40385]_ , \new_[40386]_ ,
    \new_[40390]_ , \new_[40391]_ , \new_[40395]_ , \new_[40396]_ ,
    \new_[40397]_ , \new_[40401]_ , \new_[40402]_ , \new_[40406]_ ,
    \new_[40407]_ , \new_[40408]_ , \new_[40412]_ , \new_[40413]_ ,
    \new_[40417]_ , \new_[40418]_ , \new_[40419]_ , \new_[40423]_ ,
    \new_[40424]_ , \new_[40428]_ , \new_[40429]_ , \new_[40430]_ ,
    \new_[40434]_ , \new_[40435]_ , \new_[40439]_ , \new_[40440]_ ,
    \new_[40441]_ , \new_[40445]_ , \new_[40446]_ , \new_[40450]_ ,
    \new_[40451]_ , \new_[40452]_ , \new_[40456]_ , \new_[40457]_ ,
    \new_[40461]_ , \new_[40462]_ , \new_[40463]_ , \new_[40467]_ ,
    \new_[40468]_ , \new_[40472]_ , \new_[40473]_ , \new_[40474]_ ,
    \new_[40478]_ , \new_[40479]_ , \new_[40483]_ , \new_[40484]_ ,
    \new_[40485]_ , \new_[40489]_ , \new_[40490]_ , \new_[40494]_ ,
    \new_[40495]_ , \new_[40496]_ , \new_[40500]_ , \new_[40501]_ ,
    \new_[40505]_ , \new_[40506]_ , \new_[40507]_ , \new_[40511]_ ,
    \new_[40512]_ , \new_[40516]_ , \new_[40517]_ , \new_[40518]_ ,
    \new_[40522]_ , \new_[40523]_ , \new_[40527]_ , \new_[40528]_ ,
    \new_[40529]_ , \new_[40533]_ , \new_[40534]_ , \new_[40538]_ ,
    \new_[40539]_ , \new_[40540]_ , \new_[40544]_ , \new_[40545]_ ,
    \new_[40549]_ , \new_[40550]_ , \new_[40551]_ , \new_[40555]_ ,
    \new_[40556]_ , \new_[40560]_ , \new_[40561]_ , \new_[40562]_ ,
    \new_[40566]_ , \new_[40567]_ , \new_[40571]_ , \new_[40572]_ ,
    \new_[40573]_ , \new_[40577]_ , \new_[40578]_ , \new_[40582]_ ,
    \new_[40583]_ , \new_[40584]_ , \new_[40588]_ , \new_[40589]_ ,
    \new_[40593]_ , \new_[40594]_ , \new_[40595]_ , \new_[40599]_ ,
    \new_[40600]_ , \new_[40604]_ , \new_[40605]_ , \new_[40606]_ ,
    \new_[40610]_ , \new_[40611]_ , \new_[40615]_ , \new_[40616]_ ,
    \new_[40617]_ , \new_[40621]_ , \new_[40622]_ , \new_[40626]_ ,
    \new_[40627]_ , \new_[40628]_ , \new_[40632]_ , \new_[40633]_ ,
    \new_[40637]_ , \new_[40638]_ , \new_[40639]_ , \new_[40643]_ ,
    \new_[40644]_ , \new_[40648]_ , \new_[40649]_ , \new_[40650]_ ,
    \new_[40654]_ , \new_[40655]_ , \new_[40659]_ , \new_[40660]_ ,
    \new_[40661]_ , \new_[40665]_ , \new_[40666]_ , \new_[40670]_ ,
    \new_[40671]_ , \new_[40672]_ , \new_[40676]_ , \new_[40677]_ ,
    \new_[40681]_ , \new_[40682]_ , \new_[40683]_ , \new_[40687]_ ,
    \new_[40688]_ , \new_[40692]_ , \new_[40693]_ , \new_[40694]_ ,
    \new_[40698]_ , \new_[40699]_ , \new_[40703]_ , \new_[40704]_ ,
    \new_[40705]_ , \new_[40709]_ , \new_[40710]_ , \new_[40714]_ ,
    \new_[40715]_ , \new_[40716]_ , \new_[40720]_ , \new_[40721]_ ,
    \new_[40725]_ , \new_[40726]_ , \new_[40727]_ , \new_[40731]_ ,
    \new_[40732]_ , \new_[40736]_ , \new_[40737]_ , \new_[40738]_ ,
    \new_[40742]_ , \new_[40743]_ , \new_[40747]_ , \new_[40748]_ ,
    \new_[40749]_ , \new_[40753]_ , \new_[40754]_ , \new_[40758]_ ,
    \new_[40759]_ , \new_[40760]_ , \new_[40764]_ , \new_[40765]_ ,
    \new_[40769]_ , \new_[40770]_ , \new_[40771]_ , \new_[40775]_ ,
    \new_[40776]_ , \new_[40780]_ , \new_[40781]_ , \new_[40782]_ ,
    \new_[40786]_ , \new_[40787]_ , \new_[40791]_ , \new_[40792]_ ,
    \new_[40793]_ , \new_[40797]_ , \new_[40798]_ , \new_[40802]_ ,
    \new_[40803]_ , \new_[40804]_ , \new_[40808]_ , \new_[40809]_ ,
    \new_[40813]_ , \new_[40814]_ , \new_[40815]_ , \new_[40819]_ ,
    \new_[40820]_ , \new_[40824]_ , \new_[40825]_ , \new_[40826]_ ,
    \new_[40830]_ , \new_[40831]_ , \new_[40835]_ , \new_[40836]_ ,
    \new_[40837]_ , \new_[40841]_ , \new_[40842]_ , \new_[40846]_ ,
    \new_[40847]_ , \new_[40848]_ , \new_[40852]_ , \new_[40853]_ ,
    \new_[40857]_ , \new_[40858]_ , \new_[40859]_ , \new_[40863]_ ,
    \new_[40864]_ , \new_[40868]_ , \new_[40869]_ , \new_[40870]_ ,
    \new_[40874]_ , \new_[40875]_ , \new_[40879]_ , \new_[40880]_ ,
    \new_[40881]_ , \new_[40885]_ , \new_[40886]_ , \new_[40890]_ ,
    \new_[40891]_ , \new_[40892]_ , \new_[40896]_ , \new_[40897]_ ,
    \new_[40901]_ , \new_[40902]_ , \new_[40903]_ , \new_[40907]_ ,
    \new_[40908]_ , \new_[40912]_ , \new_[40913]_ , \new_[40914]_ ,
    \new_[40918]_ , \new_[40919]_ , \new_[40923]_ , \new_[40924]_ ,
    \new_[40925]_ , \new_[40929]_ , \new_[40930]_ , \new_[40934]_ ,
    \new_[40935]_ , \new_[40936]_ , \new_[40940]_ , \new_[40941]_ ,
    \new_[40945]_ , \new_[40946]_ , \new_[40947]_ , \new_[40951]_ ,
    \new_[40952]_ , \new_[40956]_ , \new_[40957]_ , \new_[40958]_ ,
    \new_[40962]_ , \new_[40963]_ , \new_[40967]_ , \new_[40968]_ ,
    \new_[40969]_ , \new_[40973]_ , \new_[40974]_ , \new_[40978]_ ,
    \new_[40979]_ , \new_[40980]_ , \new_[40984]_ , \new_[40985]_ ,
    \new_[40989]_ , \new_[40990]_ , \new_[40991]_ , \new_[40995]_ ,
    \new_[40996]_ , \new_[41000]_ , \new_[41001]_ , \new_[41002]_ ,
    \new_[41006]_ , \new_[41007]_ , \new_[41011]_ , \new_[41012]_ ,
    \new_[41013]_ , \new_[41017]_ , \new_[41018]_ , \new_[41022]_ ,
    \new_[41023]_ , \new_[41024]_ , \new_[41028]_ , \new_[41029]_ ,
    \new_[41033]_ , \new_[41034]_ , \new_[41035]_ , \new_[41039]_ ,
    \new_[41040]_ , \new_[41044]_ , \new_[41045]_ , \new_[41046]_ ,
    \new_[41050]_ , \new_[41051]_ , \new_[41055]_ , \new_[41056]_ ,
    \new_[41057]_ , \new_[41061]_ , \new_[41062]_ , \new_[41066]_ ,
    \new_[41067]_ , \new_[41068]_ , \new_[41072]_ , \new_[41073]_ ,
    \new_[41077]_ , \new_[41078]_ , \new_[41079]_ , \new_[41083]_ ,
    \new_[41084]_ , \new_[41088]_ , \new_[41089]_ , \new_[41090]_ ,
    \new_[41094]_ , \new_[41095]_ , \new_[41099]_ , \new_[41100]_ ,
    \new_[41101]_ , \new_[41105]_ , \new_[41106]_ , \new_[41110]_ ,
    \new_[41111]_ , \new_[41112]_ , \new_[41116]_ , \new_[41117]_ ,
    \new_[41121]_ , \new_[41122]_ , \new_[41123]_ , \new_[41127]_ ,
    \new_[41128]_ , \new_[41132]_ , \new_[41133]_ , \new_[41134]_ ,
    \new_[41138]_ , \new_[41139]_ , \new_[41143]_ , \new_[41144]_ ,
    \new_[41145]_ , \new_[41149]_ , \new_[41150]_ , \new_[41154]_ ,
    \new_[41155]_ , \new_[41156]_ , \new_[41160]_ , \new_[41161]_ ,
    \new_[41165]_ , \new_[41166]_ , \new_[41167]_ , \new_[41171]_ ,
    \new_[41172]_ , \new_[41176]_ , \new_[41177]_ , \new_[41178]_ ,
    \new_[41182]_ , \new_[41183]_ , \new_[41187]_ , \new_[41188]_ ,
    \new_[41189]_ , \new_[41193]_ , \new_[41194]_ , \new_[41198]_ ,
    \new_[41199]_ , \new_[41200]_ , \new_[41204]_ , \new_[41205]_ ,
    \new_[41209]_ , \new_[41210]_ , \new_[41211]_ , \new_[41215]_ ,
    \new_[41216]_ , \new_[41220]_ , \new_[41221]_ , \new_[41222]_ ,
    \new_[41226]_ , \new_[41227]_ , \new_[41231]_ , \new_[41232]_ ,
    \new_[41233]_ , \new_[41237]_ , \new_[41238]_ , \new_[41242]_ ,
    \new_[41243]_ , \new_[41244]_ , \new_[41248]_ , \new_[41249]_ ,
    \new_[41253]_ , \new_[41254]_ , \new_[41255]_ , \new_[41259]_ ,
    \new_[41260]_ , \new_[41264]_ , \new_[41265]_ , \new_[41266]_ ,
    \new_[41270]_ , \new_[41271]_ , \new_[41275]_ , \new_[41276]_ ,
    \new_[41277]_ , \new_[41281]_ , \new_[41282]_ , \new_[41286]_ ,
    \new_[41287]_ , \new_[41288]_ , \new_[41292]_ , \new_[41293]_ ,
    \new_[41297]_ , \new_[41298]_ , \new_[41299]_ , \new_[41303]_ ,
    \new_[41304]_ , \new_[41308]_ , \new_[41309]_ , \new_[41310]_ ,
    \new_[41314]_ , \new_[41315]_ , \new_[41319]_ , \new_[41320]_ ,
    \new_[41321]_ , \new_[41325]_ , \new_[41326]_ , \new_[41329]_ ,
    \new_[41332]_ , \new_[41333]_ , \new_[41334]_ , \new_[41338]_ ,
    \new_[41339]_ , \new_[41343]_ , \new_[41344]_ , \new_[41345]_ ,
    \new_[41349]_ , \new_[41350]_ , \new_[41353]_ , \new_[41356]_ ,
    \new_[41357]_ , \new_[41358]_ , \new_[41362]_ , \new_[41363]_ ,
    \new_[41367]_ , \new_[41368]_ , \new_[41369]_ , \new_[41373]_ ,
    \new_[41374]_ , \new_[41377]_ , \new_[41380]_ , \new_[41381]_ ,
    \new_[41382]_ , \new_[41386]_ , \new_[41387]_ , \new_[41391]_ ,
    \new_[41392]_ , \new_[41393]_ , \new_[41397]_ , \new_[41398]_ ,
    \new_[41401]_ , \new_[41404]_ , \new_[41405]_ , \new_[41406]_ ,
    \new_[41410]_ , \new_[41411]_ , \new_[41415]_ , \new_[41416]_ ,
    \new_[41417]_ , \new_[41421]_ , \new_[41422]_ , \new_[41425]_ ,
    \new_[41428]_ , \new_[41429]_ , \new_[41430]_ , \new_[41434]_ ,
    \new_[41435]_ , \new_[41439]_ , \new_[41440]_ , \new_[41441]_ ,
    \new_[41445]_ , \new_[41446]_ , \new_[41449]_ , \new_[41452]_ ,
    \new_[41453]_ , \new_[41454]_ , \new_[41458]_ , \new_[41459]_ ,
    \new_[41463]_ , \new_[41464]_ , \new_[41465]_ , \new_[41469]_ ,
    \new_[41470]_ , \new_[41473]_ , \new_[41476]_ , \new_[41477]_ ,
    \new_[41478]_ , \new_[41482]_ , \new_[41483]_ , \new_[41487]_ ,
    \new_[41488]_ , \new_[41489]_ , \new_[41493]_ , \new_[41494]_ ,
    \new_[41497]_ , \new_[41500]_ , \new_[41501]_ , \new_[41502]_ ,
    \new_[41506]_ , \new_[41507]_ , \new_[41511]_ , \new_[41512]_ ,
    \new_[41513]_ , \new_[41517]_ , \new_[41518]_ , \new_[41521]_ ,
    \new_[41524]_ , \new_[41525]_ , \new_[41526]_ , \new_[41530]_ ,
    \new_[41531]_ , \new_[41535]_ , \new_[41536]_ , \new_[41537]_ ,
    \new_[41541]_ , \new_[41542]_ , \new_[41545]_ , \new_[41548]_ ,
    \new_[41549]_ , \new_[41550]_ , \new_[41554]_ , \new_[41555]_ ,
    \new_[41559]_ , \new_[41560]_ , \new_[41561]_ , \new_[41565]_ ,
    \new_[41566]_ , \new_[41569]_ , \new_[41572]_ , \new_[41573]_ ,
    \new_[41574]_ , \new_[41578]_ , \new_[41579]_ , \new_[41583]_ ,
    \new_[41584]_ , \new_[41585]_ , \new_[41589]_ , \new_[41590]_ ,
    \new_[41593]_ , \new_[41596]_ , \new_[41597]_ , \new_[41598]_ ,
    \new_[41602]_ , \new_[41603]_ , \new_[41607]_ , \new_[41608]_ ,
    \new_[41609]_ , \new_[41613]_ , \new_[41614]_ , \new_[41617]_ ,
    \new_[41620]_ , \new_[41621]_ , \new_[41622]_ , \new_[41626]_ ,
    \new_[41627]_ , \new_[41631]_ , \new_[41632]_ , \new_[41633]_ ,
    \new_[41637]_ , \new_[41638]_ , \new_[41641]_ , \new_[41644]_ ,
    \new_[41645]_ , \new_[41646]_ , \new_[41650]_ , \new_[41651]_ ,
    \new_[41655]_ , \new_[41656]_ , \new_[41657]_ , \new_[41661]_ ,
    \new_[41662]_ , \new_[41665]_ , \new_[41668]_ , \new_[41669]_ ,
    \new_[41670]_ , \new_[41674]_ , \new_[41675]_ , \new_[41679]_ ,
    \new_[41680]_ , \new_[41681]_ , \new_[41685]_ , \new_[41686]_ ,
    \new_[41689]_ , \new_[41692]_ , \new_[41693]_ , \new_[41694]_ ,
    \new_[41698]_ , \new_[41699]_ , \new_[41703]_ , \new_[41704]_ ,
    \new_[41705]_ , \new_[41709]_ , \new_[41710]_ , \new_[41713]_ ,
    \new_[41716]_ , \new_[41717]_ , \new_[41718]_ , \new_[41722]_ ,
    \new_[41723]_ , \new_[41727]_ , \new_[41728]_ , \new_[41729]_ ,
    \new_[41733]_ , \new_[41734]_ , \new_[41737]_ , \new_[41740]_ ,
    \new_[41741]_ , \new_[41742]_ , \new_[41746]_ , \new_[41747]_ ,
    \new_[41751]_ , \new_[41752]_ , \new_[41753]_ , \new_[41757]_ ,
    \new_[41758]_ , \new_[41761]_ , \new_[41764]_ , \new_[41765]_ ,
    \new_[41766]_ , \new_[41770]_ , \new_[41771]_ , \new_[41775]_ ,
    \new_[41776]_ , \new_[41777]_ , \new_[41781]_ , \new_[41782]_ ,
    \new_[41785]_ , \new_[41788]_ , \new_[41789]_ , \new_[41790]_ ,
    \new_[41794]_ , \new_[41795]_ , \new_[41799]_ , \new_[41800]_ ,
    \new_[41801]_ , \new_[41805]_ , \new_[41806]_ , \new_[41809]_ ,
    \new_[41812]_ , \new_[41813]_ , \new_[41814]_ , \new_[41818]_ ,
    \new_[41819]_ , \new_[41823]_ , \new_[41824]_ , \new_[41825]_ ,
    \new_[41829]_ , \new_[41830]_ , \new_[41833]_ , \new_[41836]_ ,
    \new_[41837]_ , \new_[41838]_ , \new_[41842]_ , \new_[41843]_ ,
    \new_[41847]_ , \new_[41848]_ , \new_[41849]_ , \new_[41853]_ ,
    \new_[41854]_ , \new_[41857]_ , \new_[41860]_ , \new_[41861]_ ,
    \new_[41862]_ , \new_[41866]_ , \new_[41867]_ , \new_[41871]_ ,
    \new_[41872]_ , \new_[41873]_ , \new_[41877]_ , \new_[41878]_ ,
    \new_[41881]_ , \new_[41884]_ , \new_[41885]_ , \new_[41886]_ ,
    \new_[41890]_ , \new_[41891]_ , \new_[41895]_ , \new_[41896]_ ,
    \new_[41897]_ , \new_[41901]_ , \new_[41902]_ , \new_[41905]_ ,
    \new_[41908]_ , \new_[41909]_ , \new_[41910]_ , \new_[41914]_ ,
    \new_[41915]_ , \new_[41919]_ , \new_[41920]_ , \new_[41921]_ ,
    \new_[41925]_ , \new_[41926]_ , \new_[41929]_ , \new_[41932]_ ,
    \new_[41933]_ , \new_[41934]_ , \new_[41938]_ , \new_[41939]_ ,
    \new_[41943]_ , \new_[41944]_ , \new_[41945]_ , \new_[41949]_ ,
    \new_[41950]_ , \new_[41953]_ , \new_[41956]_ , \new_[41957]_ ,
    \new_[41958]_ , \new_[41962]_ , \new_[41963]_ , \new_[41967]_ ,
    \new_[41968]_ , \new_[41969]_ , \new_[41973]_ , \new_[41974]_ ,
    \new_[41977]_ , \new_[41980]_ , \new_[41981]_ , \new_[41982]_ ,
    \new_[41986]_ , \new_[41987]_ , \new_[41991]_ , \new_[41992]_ ,
    \new_[41993]_ , \new_[41997]_ , \new_[41998]_ , \new_[42001]_ ,
    \new_[42004]_ , \new_[42005]_ , \new_[42006]_ , \new_[42010]_ ,
    \new_[42011]_ , \new_[42015]_ , \new_[42016]_ , \new_[42017]_ ,
    \new_[42021]_ , \new_[42022]_ , \new_[42025]_ , \new_[42028]_ ,
    \new_[42029]_ , \new_[42030]_ , \new_[42034]_ , \new_[42035]_ ,
    \new_[42039]_ , \new_[42040]_ , \new_[42041]_ , \new_[42045]_ ,
    \new_[42046]_ , \new_[42049]_ , \new_[42052]_ , \new_[42053]_ ,
    \new_[42054]_ , \new_[42058]_ , \new_[42059]_ , \new_[42063]_ ,
    \new_[42064]_ , \new_[42065]_ , \new_[42069]_ , \new_[42070]_ ,
    \new_[42073]_ , \new_[42076]_ , \new_[42077]_ , \new_[42078]_ ,
    \new_[42082]_ , \new_[42083]_ , \new_[42087]_ , \new_[42088]_ ,
    \new_[42089]_ , \new_[42093]_ , \new_[42094]_ , \new_[42097]_ ,
    \new_[42100]_ , \new_[42101]_ , \new_[42102]_ , \new_[42106]_ ,
    \new_[42107]_ , \new_[42111]_ , \new_[42112]_ , \new_[42113]_ ,
    \new_[42117]_ , \new_[42118]_ , \new_[42121]_ , \new_[42124]_ ,
    \new_[42125]_ , \new_[42126]_ , \new_[42130]_ , \new_[42131]_ ,
    \new_[42135]_ , \new_[42136]_ , \new_[42137]_ , \new_[42141]_ ,
    \new_[42142]_ , \new_[42145]_ , \new_[42148]_ , \new_[42149]_ ,
    \new_[42150]_ , \new_[42154]_ , \new_[42155]_ , \new_[42159]_ ,
    \new_[42160]_ , \new_[42161]_ , \new_[42165]_ , \new_[42166]_ ,
    \new_[42169]_ , \new_[42172]_ , \new_[42173]_ , \new_[42174]_ ,
    \new_[42178]_ , \new_[42179]_ , \new_[42183]_ , \new_[42184]_ ,
    \new_[42185]_ , \new_[42189]_ , \new_[42190]_ , \new_[42193]_ ,
    \new_[42196]_ , \new_[42197]_ , \new_[42198]_ , \new_[42202]_ ,
    \new_[42203]_ , \new_[42207]_ , \new_[42208]_ , \new_[42209]_ ,
    \new_[42213]_ , \new_[42214]_ , \new_[42217]_ , \new_[42220]_ ,
    \new_[42221]_ , \new_[42222]_ , \new_[42226]_ , \new_[42227]_ ,
    \new_[42231]_ , \new_[42232]_ , \new_[42233]_ , \new_[42237]_ ,
    \new_[42238]_ , \new_[42241]_ , \new_[42244]_ , \new_[42245]_ ,
    \new_[42246]_ , \new_[42250]_ , \new_[42251]_ , \new_[42255]_ ,
    \new_[42256]_ , \new_[42257]_ , \new_[42261]_ , \new_[42262]_ ,
    \new_[42265]_ , \new_[42268]_ , \new_[42269]_ , \new_[42270]_ ,
    \new_[42274]_ , \new_[42275]_ , \new_[42279]_ , \new_[42280]_ ,
    \new_[42281]_ , \new_[42285]_ , \new_[42286]_ , \new_[42289]_ ,
    \new_[42292]_ , \new_[42293]_ , \new_[42294]_ , \new_[42298]_ ,
    \new_[42299]_ , \new_[42303]_ , \new_[42304]_ , \new_[42305]_ ,
    \new_[42309]_ , \new_[42310]_ , \new_[42313]_ , \new_[42316]_ ,
    \new_[42317]_ , \new_[42318]_ , \new_[42322]_ , \new_[42323]_ ,
    \new_[42327]_ , \new_[42328]_ , \new_[42329]_ , \new_[42333]_ ,
    \new_[42334]_ , \new_[42337]_ , \new_[42340]_ , \new_[42341]_ ,
    \new_[42342]_ , \new_[42346]_ , \new_[42347]_ , \new_[42351]_ ,
    \new_[42352]_ , \new_[42353]_ , \new_[42357]_ , \new_[42358]_ ,
    \new_[42361]_ , \new_[42364]_ , \new_[42365]_ , \new_[42366]_ ,
    \new_[42370]_ , \new_[42371]_ , \new_[42375]_ , \new_[42376]_ ,
    \new_[42377]_ , \new_[42381]_ , \new_[42382]_ , \new_[42385]_ ,
    \new_[42388]_ , \new_[42389]_ , \new_[42390]_ , \new_[42394]_ ,
    \new_[42395]_ , \new_[42399]_ , \new_[42400]_ , \new_[42401]_ ,
    \new_[42405]_ , \new_[42406]_ , \new_[42409]_ , \new_[42412]_ ,
    \new_[42413]_ , \new_[42414]_ , \new_[42418]_ , \new_[42419]_ ,
    \new_[42423]_ , \new_[42424]_ , \new_[42425]_ , \new_[42429]_ ,
    \new_[42430]_ , \new_[42433]_ , \new_[42436]_ , \new_[42437]_ ,
    \new_[42438]_ , \new_[42442]_ , \new_[42443]_ , \new_[42447]_ ,
    \new_[42448]_ , \new_[42449]_ , \new_[42453]_ , \new_[42454]_ ,
    \new_[42457]_ , \new_[42460]_ , \new_[42461]_ , \new_[42462]_ ,
    \new_[42466]_ , \new_[42467]_ , \new_[42471]_ , \new_[42472]_ ,
    \new_[42473]_ , \new_[42477]_ , \new_[42478]_ , \new_[42481]_ ,
    \new_[42484]_ , \new_[42485]_ , \new_[42486]_ , \new_[42490]_ ,
    \new_[42491]_ , \new_[42495]_ , \new_[42496]_ , \new_[42497]_ ,
    \new_[42501]_ , \new_[42502]_ , \new_[42505]_ , \new_[42508]_ ,
    \new_[42509]_ , \new_[42510]_ , \new_[42514]_ , \new_[42515]_ ,
    \new_[42519]_ , \new_[42520]_ , \new_[42521]_ , \new_[42525]_ ,
    \new_[42526]_ , \new_[42529]_ , \new_[42532]_ , \new_[42533]_ ,
    \new_[42534]_ , \new_[42538]_ , \new_[42539]_ , \new_[42543]_ ,
    \new_[42544]_ , \new_[42545]_ , \new_[42549]_ , \new_[42550]_ ,
    \new_[42553]_ , \new_[42556]_ , \new_[42557]_ , \new_[42558]_ ,
    \new_[42562]_ , \new_[42563]_ , \new_[42567]_ , \new_[42568]_ ,
    \new_[42569]_ , \new_[42573]_ , \new_[42574]_ , \new_[42577]_ ,
    \new_[42580]_ , \new_[42581]_ , \new_[42582]_ , \new_[42586]_ ,
    \new_[42587]_ , \new_[42591]_ , \new_[42592]_ , \new_[42593]_ ,
    \new_[42597]_ , \new_[42598]_ , \new_[42601]_ , \new_[42604]_ ,
    \new_[42605]_ , \new_[42606]_ , \new_[42610]_ , \new_[42611]_ ,
    \new_[42615]_ , \new_[42616]_ , \new_[42617]_ , \new_[42621]_ ,
    \new_[42622]_ , \new_[42625]_ , \new_[42628]_ , \new_[42629]_ ,
    \new_[42630]_ , \new_[42634]_ , \new_[42635]_ , \new_[42639]_ ,
    \new_[42640]_ , \new_[42641]_ , \new_[42645]_ , \new_[42646]_ ,
    \new_[42649]_ , \new_[42652]_ , \new_[42653]_ , \new_[42654]_ ,
    \new_[42658]_ , \new_[42659]_ , \new_[42663]_ , \new_[42664]_ ,
    \new_[42665]_ , \new_[42669]_ , \new_[42670]_ , \new_[42673]_ ,
    \new_[42676]_ , \new_[42677]_ , \new_[42678]_ , \new_[42682]_ ,
    \new_[42683]_ , \new_[42687]_ , \new_[42688]_ , \new_[42689]_ ,
    \new_[42693]_ , \new_[42694]_ , \new_[42697]_ , \new_[42700]_ ,
    \new_[42701]_ , \new_[42702]_ , \new_[42706]_ , \new_[42707]_ ,
    \new_[42711]_ , \new_[42712]_ , \new_[42713]_ , \new_[42717]_ ,
    \new_[42718]_ , \new_[42721]_ , \new_[42724]_ , \new_[42725]_ ,
    \new_[42726]_ , \new_[42730]_ , \new_[42731]_ , \new_[42735]_ ,
    \new_[42736]_ , \new_[42737]_ , \new_[42741]_ , \new_[42742]_ ,
    \new_[42745]_ , \new_[42748]_ , \new_[42749]_ , \new_[42750]_ ,
    \new_[42754]_ , \new_[42755]_ , \new_[42759]_ , \new_[42760]_ ,
    \new_[42761]_ , \new_[42765]_ , \new_[42766]_ , \new_[42769]_ ,
    \new_[42772]_ , \new_[42773]_ , \new_[42774]_ , \new_[42778]_ ,
    \new_[42779]_ , \new_[42783]_ , \new_[42784]_ , \new_[42785]_ ,
    \new_[42789]_ , \new_[42790]_ , \new_[42793]_ , \new_[42796]_ ,
    \new_[42797]_ , \new_[42798]_ , \new_[42802]_ , \new_[42803]_ ,
    \new_[42807]_ , \new_[42808]_ , \new_[42809]_ , \new_[42813]_ ,
    \new_[42814]_ , \new_[42817]_ , \new_[42820]_ , \new_[42821]_ ,
    \new_[42822]_ , \new_[42826]_ , \new_[42827]_ , \new_[42831]_ ,
    \new_[42832]_ , \new_[42833]_ , \new_[42837]_ , \new_[42838]_ ,
    \new_[42841]_ , \new_[42844]_ , \new_[42845]_ , \new_[42846]_ ,
    \new_[42850]_ , \new_[42851]_ , \new_[42855]_ , \new_[42856]_ ,
    \new_[42857]_ , \new_[42861]_ , \new_[42862]_ , \new_[42865]_ ,
    \new_[42868]_ , \new_[42869]_ , \new_[42870]_ , \new_[42874]_ ,
    \new_[42875]_ , \new_[42879]_ , \new_[42880]_ , \new_[42881]_ ,
    \new_[42885]_ , \new_[42886]_ , \new_[42889]_ , \new_[42892]_ ,
    \new_[42893]_ , \new_[42894]_ , \new_[42898]_ , \new_[42899]_ ,
    \new_[42903]_ , \new_[42904]_ , \new_[42905]_ , \new_[42909]_ ,
    \new_[42910]_ , \new_[42913]_ , \new_[42916]_ , \new_[42917]_ ,
    \new_[42918]_ , \new_[42922]_ , \new_[42923]_ , \new_[42927]_ ,
    \new_[42928]_ , \new_[42929]_ , \new_[42933]_ , \new_[42934]_ ,
    \new_[42937]_ , \new_[42940]_ , \new_[42941]_ , \new_[42942]_ ,
    \new_[42946]_ , \new_[42947]_ , \new_[42951]_ , \new_[42952]_ ,
    \new_[42953]_ , \new_[42957]_ , \new_[42958]_ , \new_[42961]_ ,
    \new_[42964]_ , \new_[42965]_ , \new_[42966]_ , \new_[42970]_ ,
    \new_[42971]_ , \new_[42975]_ , \new_[42976]_ , \new_[42977]_ ,
    \new_[42981]_ , \new_[42982]_ , \new_[42985]_ , \new_[42988]_ ,
    \new_[42989]_ , \new_[42990]_ , \new_[42994]_ , \new_[42995]_ ,
    \new_[42999]_ , \new_[43000]_ , \new_[43001]_ , \new_[43005]_ ,
    \new_[43006]_ , \new_[43009]_ , \new_[43012]_ , \new_[43013]_ ,
    \new_[43014]_ , \new_[43018]_ , \new_[43019]_ , \new_[43023]_ ,
    \new_[43024]_ , \new_[43025]_ , \new_[43029]_ , \new_[43030]_ ,
    \new_[43033]_ , \new_[43036]_ , \new_[43037]_ , \new_[43038]_ ,
    \new_[43042]_ , \new_[43043]_ , \new_[43047]_ , \new_[43048]_ ,
    \new_[43049]_ , \new_[43053]_ , \new_[43054]_ , \new_[43057]_ ,
    \new_[43060]_ , \new_[43061]_ , \new_[43062]_ , \new_[43066]_ ,
    \new_[43067]_ , \new_[43071]_ , \new_[43072]_ , \new_[43073]_ ,
    \new_[43077]_ , \new_[43078]_ , \new_[43081]_ , \new_[43084]_ ,
    \new_[43085]_ , \new_[43086]_ , \new_[43090]_ , \new_[43091]_ ,
    \new_[43095]_ , \new_[43096]_ , \new_[43097]_ , \new_[43101]_ ,
    \new_[43102]_ , \new_[43105]_ , \new_[43108]_ , \new_[43109]_ ,
    \new_[43110]_ , \new_[43114]_ , \new_[43115]_ , \new_[43119]_ ,
    \new_[43120]_ , \new_[43121]_ , \new_[43125]_ , \new_[43126]_ ,
    \new_[43129]_ , \new_[43132]_ , \new_[43133]_ , \new_[43134]_ ,
    \new_[43138]_ , \new_[43139]_ , \new_[43143]_ , \new_[43144]_ ,
    \new_[43145]_ , \new_[43149]_ , \new_[43150]_ , \new_[43153]_ ,
    \new_[43156]_ , \new_[43157]_ , \new_[43158]_ , \new_[43162]_ ,
    \new_[43163]_ , \new_[43167]_ , \new_[43168]_ , \new_[43169]_ ,
    \new_[43173]_ , \new_[43174]_ , \new_[43177]_ , \new_[43180]_ ,
    \new_[43181]_ , \new_[43182]_ , \new_[43186]_ , \new_[43187]_ ,
    \new_[43191]_ , \new_[43192]_ , \new_[43193]_ , \new_[43197]_ ,
    \new_[43198]_ , \new_[43201]_ , \new_[43204]_ , \new_[43205]_ ,
    \new_[43206]_ , \new_[43210]_ , \new_[43211]_ , \new_[43215]_ ,
    \new_[43216]_ , \new_[43217]_ , \new_[43221]_ , \new_[43222]_ ,
    \new_[43225]_ , \new_[43228]_ , \new_[43229]_ , \new_[43230]_ ,
    \new_[43234]_ , \new_[43235]_ , \new_[43239]_ , \new_[43240]_ ,
    \new_[43241]_ , \new_[43245]_ , \new_[43246]_ , \new_[43249]_ ,
    \new_[43252]_ , \new_[43253]_ , \new_[43254]_ , \new_[43258]_ ,
    \new_[43259]_ , \new_[43263]_ , \new_[43264]_ , \new_[43265]_ ,
    \new_[43269]_ , \new_[43270]_ , \new_[43273]_ , \new_[43276]_ ,
    \new_[43277]_ , \new_[43278]_ , \new_[43282]_ , \new_[43283]_ ,
    \new_[43287]_ , \new_[43288]_ , \new_[43289]_ , \new_[43293]_ ,
    \new_[43294]_ , \new_[43297]_ , \new_[43300]_ , \new_[43301]_ ,
    \new_[43302]_ , \new_[43306]_ , \new_[43307]_ , \new_[43311]_ ,
    \new_[43312]_ , \new_[43313]_ , \new_[43317]_ , \new_[43318]_ ,
    \new_[43321]_ , \new_[43324]_ , \new_[43325]_ , \new_[43326]_ ,
    \new_[43330]_ , \new_[43331]_ , \new_[43335]_ , \new_[43336]_ ,
    \new_[43337]_ , \new_[43341]_ , \new_[43342]_ , \new_[43345]_ ,
    \new_[43348]_ , \new_[43349]_ , \new_[43350]_ , \new_[43354]_ ,
    \new_[43355]_ , \new_[43359]_ , \new_[43360]_ , \new_[43361]_ ,
    \new_[43365]_ , \new_[43366]_ , \new_[43369]_ , \new_[43372]_ ,
    \new_[43373]_ , \new_[43374]_ , \new_[43378]_ , \new_[43379]_ ,
    \new_[43383]_ , \new_[43384]_ , \new_[43385]_ , \new_[43389]_ ,
    \new_[43390]_ , \new_[43393]_ , \new_[43396]_ , \new_[43397]_ ,
    \new_[43398]_ , \new_[43402]_ , \new_[43403]_ , \new_[43407]_ ,
    \new_[43408]_ , \new_[43409]_ , \new_[43413]_ , \new_[43414]_ ,
    \new_[43417]_ , \new_[43420]_ , \new_[43421]_ , \new_[43422]_ ,
    \new_[43426]_ , \new_[43427]_ , \new_[43431]_ , \new_[43432]_ ,
    \new_[43433]_ , \new_[43437]_ , \new_[43438]_ , \new_[43441]_ ,
    \new_[43444]_ , \new_[43445]_ , \new_[43446]_ , \new_[43450]_ ,
    \new_[43451]_ , \new_[43455]_ , \new_[43456]_ , \new_[43457]_ ,
    \new_[43461]_ , \new_[43462]_ , \new_[43465]_ , \new_[43468]_ ,
    \new_[43469]_ , \new_[43470]_ , \new_[43474]_ , \new_[43475]_ ,
    \new_[43479]_ , \new_[43480]_ , \new_[43481]_ , \new_[43485]_ ,
    \new_[43486]_ , \new_[43489]_ , \new_[43492]_ , \new_[43493]_ ,
    \new_[43494]_ , \new_[43498]_ , \new_[43499]_ , \new_[43503]_ ,
    \new_[43504]_ , \new_[43505]_ , \new_[43509]_ , \new_[43510]_ ,
    \new_[43513]_ , \new_[43516]_ , \new_[43517]_ , \new_[43518]_ ,
    \new_[43522]_ , \new_[43523]_ , \new_[43527]_ , \new_[43528]_ ,
    \new_[43529]_ , \new_[43533]_ , \new_[43534]_ , \new_[43537]_ ,
    \new_[43540]_ , \new_[43541]_ , \new_[43542]_ , \new_[43546]_ ,
    \new_[43547]_ , \new_[43551]_ , \new_[43552]_ , \new_[43553]_ ,
    \new_[43557]_ , \new_[43558]_ , \new_[43561]_ , \new_[43564]_ ,
    \new_[43565]_ , \new_[43566]_ , \new_[43570]_ , \new_[43571]_ ,
    \new_[43575]_ , \new_[43576]_ , \new_[43577]_ , \new_[43581]_ ,
    \new_[43582]_ , \new_[43585]_ , \new_[43588]_ , \new_[43589]_ ,
    \new_[43590]_ , \new_[43594]_ , \new_[43595]_ , \new_[43599]_ ,
    \new_[43600]_ , \new_[43601]_ , \new_[43605]_ , \new_[43606]_ ,
    \new_[43609]_ , \new_[43612]_ , \new_[43613]_ , \new_[43614]_ ,
    \new_[43618]_ , \new_[43619]_ , \new_[43623]_ , \new_[43624]_ ,
    \new_[43625]_ , \new_[43629]_ , \new_[43630]_ , \new_[43633]_ ,
    \new_[43636]_ , \new_[43637]_ , \new_[43638]_ , \new_[43642]_ ,
    \new_[43643]_ , \new_[43647]_ , \new_[43648]_ , \new_[43649]_ ,
    \new_[43653]_ , \new_[43654]_ , \new_[43657]_ , \new_[43660]_ ,
    \new_[43661]_ , \new_[43662]_ , \new_[43666]_ , \new_[43667]_ ,
    \new_[43671]_ , \new_[43672]_ , \new_[43673]_ , \new_[43677]_ ,
    \new_[43678]_ , \new_[43681]_ , \new_[43684]_ , \new_[43685]_ ,
    \new_[43686]_ , \new_[43690]_ , \new_[43691]_ , \new_[43695]_ ,
    \new_[43696]_ , \new_[43697]_ , \new_[43701]_ , \new_[43702]_ ,
    \new_[43705]_ , \new_[43708]_ , \new_[43709]_ , \new_[43710]_ ,
    \new_[43714]_ , \new_[43715]_ , \new_[43719]_ , \new_[43720]_ ,
    \new_[43721]_ , \new_[43725]_ , \new_[43726]_ , \new_[43729]_ ,
    \new_[43732]_ , \new_[43733]_ , \new_[43734]_ , \new_[43738]_ ,
    \new_[43739]_ , \new_[43743]_ , \new_[43744]_ , \new_[43745]_ ,
    \new_[43749]_ , \new_[43750]_ , \new_[43753]_ , \new_[43756]_ ,
    \new_[43757]_ , \new_[43758]_ , \new_[43762]_ , \new_[43763]_ ,
    \new_[43767]_ , \new_[43768]_ , \new_[43769]_ , \new_[43773]_ ,
    \new_[43774]_ , \new_[43777]_ , \new_[43780]_ , \new_[43781]_ ,
    \new_[43782]_ , \new_[43786]_ , \new_[43787]_ , \new_[43791]_ ,
    \new_[43792]_ , \new_[43793]_ , \new_[43797]_ , \new_[43798]_ ,
    \new_[43801]_ , \new_[43804]_ , \new_[43805]_ , \new_[43806]_ ,
    \new_[43810]_ , \new_[43811]_ , \new_[43815]_ , \new_[43816]_ ,
    \new_[43817]_ , \new_[43821]_ , \new_[43822]_ , \new_[43825]_ ,
    \new_[43828]_ , \new_[43829]_ , \new_[43830]_ , \new_[43834]_ ,
    \new_[43835]_ , \new_[43839]_ , \new_[43840]_ , \new_[43841]_ ,
    \new_[43845]_ , \new_[43846]_ , \new_[43849]_ , \new_[43852]_ ,
    \new_[43853]_ , \new_[43854]_ , \new_[43858]_ , \new_[43859]_ ,
    \new_[43863]_ , \new_[43864]_ , \new_[43865]_ , \new_[43869]_ ,
    \new_[43870]_ , \new_[43873]_ , \new_[43876]_ , \new_[43877]_ ,
    \new_[43878]_ , \new_[43882]_ , \new_[43883]_ , \new_[43887]_ ,
    \new_[43888]_ , \new_[43889]_ , \new_[43893]_ , \new_[43894]_ ,
    \new_[43897]_ , \new_[43900]_ , \new_[43901]_ , \new_[43902]_ ,
    \new_[43906]_ , \new_[43907]_ , \new_[43911]_ , \new_[43912]_ ,
    \new_[43913]_ , \new_[43917]_ , \new_[43918]_ , \new_[43921]_ ,
    \new_[43924]_ , \new_[43925]_ , \new_[43926]_ , \new_[43930]_ ,
    \new_[43931]_ , \new_[43935]_ , \new_[43936]_ , \new_[43937]_ ,
    \new_[43941]_ , \new_[43942]_ , \new_[43945]_ , \new_[43948]_ ,
    \new_[43949]_ , \new_[43950]_ , \new_[43954]_ , \new_[43955]_ ,
    \new_[43959]_ , \new_[43960]_ , \new_[43961]_ , \new_[43965]_ ,
    \new_[43966]_ , \new_[43969]_ , \new_[43972]_ , \new_[43973]_ ,
    \new_[43974]_ , \new_[43978]_ , \new_[43979]_ , \new_[43983]_ ,
    \new_[43984]_ , \new_[43985]_ , \new_[43989]_ , \new_[43990]_ ,
    \new_[43993]_ , \new_[43996]_ , \new_[43997]_ , \new_[43998]_ ,
    \new_[44002]_ , \new_[44003]_ , \new_[44007]_ , \new_[44008]_ ,
    \new_[44009]_ , \new_[44013]_ , \new_[44014]_ , \new_[44017]_ ,
    \new_[44020]_ , \new_[44021]_ , \new_[44022]_ , \new_[44026]_ ,
    \new_[44027]_ , \new_[44031]_ , \new_[44032]_ , \new_[44033]_ ,
    \new_[44037]_ , \new_[44038]_ , \new_[44041]_ , \new_[44044]_ ,
    \new_[44045]_ , \new_[44046]_ , \new_[44050]_ , \new_[44051]_ ,
    \new_[44055]_ , \new_[44056]_ , \new_[44057]_ , \new_[44061]_ ,
    \new_[44062]_ , \new_[44065]_ , \new_[44068]_ , \new_[44069]_ ,
    \new_[44070]_ , \new_[44074]_ , \new_[44075]_ , \new_[44079]_ ,
    \new_[44080]_ , \new_[44081]_ , \new_[44085]_ , \new_[44086]_ ,
    \new_[44089]_ , \new_[44092]_ , \new_[44093]_ , \new_[44094]_ ,
    \new_[44098]_ , \new_[44099]_ , \new_[44103]_ , \new_[44104]_ ,
    \new_[44105]_ , \new_[44109]_ , \new_[44110]_ , \new_[44113]_ ,
    \new_[44116]_ , \new_[44117]_ , \new_[44118]_ , \new_[44122]_ ,
    \new_[44123]_ , \new_[44127]_ , \new_[44128]_ , \new_[44129]_ ,
    \new_[44133]_ , \new_[44134]_ , \new_[44137]_ , \new_[44140]_ ,
    \new_[44141]_ , \new_[44142]_ , \new_[44146]_ , \new_[44147]_ ,
    \new_[44151]_ , \new_[44152]_ , \new_[44153]_ , \new_[44157]_ ,
    \new_[44158]_ , \new_[44161]_ , \new_[44164]_ , \new_[44165]_ ,
    \new_[44166]_ , \new_[44170]_ , \new_[44171]_ , \new_[44175]_ ,
    \new_[44176]_ , \new_[44177]_ , \new_[44181]_ , \new_[44182]_ ,
    \new_[44185]_ , \new_[44188]_ , \new_[44189]_ , \new_[44190]_ ,
    \new_[44194]_ , \new_[44195]_ , \new_[44199]_ , \new_[44200]_ ,
    \new_[44201]_ , \new_[44205]_ , \new_[44206]_ , \new_[44209]_ ,
    \new_[44212]_ , \new_[44213]_ , \new_[44214]_ , \new_[44218]_ ,
    \new_[44219]_ , \new_[44223]_ , \new_[44224]_ , \new_[44225]_ ,
    \new_[44229]_ , \new_[44230]_ , \new_[44233]_ , \new_[44236]_ ,
    \new_[44237]_ , \new_[44238]_ , \new_[44242]_ , \new_[44243]_ ,
    \new_[44247]_ , \new_[44248]_ , \new_[44249]_ , \new_[44253]_ ,
    \new_[44254]_ , \new_[44257]_ , \new_[44260]_ , \new_[44261]_ ,
    \new_[44262]_ , \new_[44266]_ , \new_[44267]_ , \new_[44271]_ ,
    \new_[44272]_ , \new_[44273]_ , \new_[44277]_ , \new_[44278]_ ,
    \new_[44281]_ , \new_[44284]_ , \new_[44285]_ , \new_[44286]_ ,
    \new_[44290]_ , \new_[44291]_ , \new_[44295]_ , \new_[44296]_ ,
    \new_[44297]_ , \new_[44301]_ , \new_[44302]_ , \new_[44305]_ ,
    \new_[44308]_ , \new_[44309]_ , \new_[44310]_ , \new_[44314]_ ,
    \new_[44315]_ , \new_[44319]_ , \new_[44320]_ , \new_[44321]_ ,
    \new_[44325]_ , \new_[44326]_ , \new_[44329]_ , \new_[44332]_ ,
    \new_[44333]_ , \new_[44334]_ , \new_[44338]_ , \new_[44339]_ ,
    \new_[44343]_ , \new_[44344]_ , \new_[44345]_ , \new_[44349]_ ,
    \new_[44350]_ , \new_[44353]_ , \new_[44356]_ , \new_[44357]_ ,
    \new_[44358]_ , \new_[44362]_ , \new_[44363]_ , \new_[44367]_ ,
    \new_[44368]_ , \new_[44369]_ , \new_[44373]_ , \new_[44374]_ ,
    \new_[44377]_ , \new_[44380]_ , \new_[44381]_ , \new_[44382]_ ,
    \new_[44386]_ , \new_[44387]_ , \new_[44391]_ , \new_[44392]_ ,
    \new_[44393]_ , \new_[44397]_ , \new_[44398]_ , \new_[44401]_ ,
    \new_[44404]_ , \new_[44405]_ , \new_[44406]_ , \new_[44410]_ ,
    \new_[44411]_ , \new_[44415]_ , \new_[44416]_ , \new_[44417]_ ,
    \new_[44421]_ , \new_[44422]_ , \new_[44425]_ , \new_[44428]_ ,
    \new_[44429]_ , \new_[44430]_ , \new_[44434]_ , \new_[44435]_ ,
    \new_[44439]_ , \new_[44440]_ , \new_[44441]_ , \new_[44445]_ ,
    \new_[44446]_ , \new_[44449]_ , \new_[44452]_ , \new_[44453]_ ,
    \new_[44454]_ , \new_[44458]_ , \new_[44459]_ , \new_[44463]_ ,
    \new_[44464]_ , \new_[44465]_ , \new_[44469]_ , \new_[44470]_ ,
    \new_[44473]_ , \new_[44476]_ , \new_[44477]_ , \new_[44478]_ ,
    \new_[44482]_ , \new_[44483]_ , \new_[44487]_ , \new_[44488]_ ,
    \new_[44489]_ , \new_[44493]_ , \new_[44494]_ , \new_[44497]_ ,
    \new_[44500]_ , \new_[44501]_ , \new_[44502]_ , \new_[44506]_ ,
    \new_[44507]_ , \new_[44511]_ , \new_[44512]_ , \new_[44513]_ ,
    \new_[44517]_ , \new_[44518]_ , \new_[44521]_ , \new_[44524]_ ,
    \new_[44525]_ , \new_[44526]_ , \new_[44530]_ , \new_[44531]_ ,
    \new_[44535]_ , \new_[44536]_ , \new_[44537]_ , \new_[44541]_ ,
    \new_[44542]_ , \new_[44545]_ , \new_[44548]_ , \new_[44549]_ ,
    \new_[44550]_ , \new_[44554]_ , \new_[44555]_ , \new_[44559]_ ,
    \new_[44560]_ , \new_[44561]_ , \new_[44565]_ , \new_[44566]_ ,
    \new_[44569]_ , \new_[44572]_ , \new_[44573]_ , \new_[44574]_ ,
    \new_[44578]_ , \new_[44579]_ , \new_[44583]_ , \new_[44584]_ ,
    \new_[44585]_ , \new_[44589]_ , \new_[44590]_ , \new_[44593]_ ,
    \new_[44596]_ , \new_[44597]_ , \new_[44598]_ , \new_[44602]_ ,
    \new_[44603]_ , \new_[44607]_ , \new_[44608]_ , \new_[44609]_ ,
    \new_[44613]_ , \new_[44614]_ , \new_[44617]_ , \new_[44620]_ ,
    \new_[44621]_ , \new_[44622]_ , \new_[44626]_ , \new_[44627]_ ,
    \new_[44631]_ , \new_[44632]_ , \new_[44633]_ , \new_[44637]_ ,
    \new_[44638]_ , \new_[44641]_ , \new_[44644]_ , \new_[44645]_ ,
    \new_[44646]_ , \new_[44650]_ , \new_[44651]_ , \new_[44655]_ ,
    \new_[44656]_ , \new_[44657]_ , \new_[44661]_ , \new_[44662]_ ,
    \new_[44665]_ , \new_[44668]_ , \new_[44669]_ , \new_[44670]_ ,
    \new_[44674]_ , \new_[44675]_ , \new_[44679]_ , \new_[44680]_ ,
    \new_[44681]_ , \new_[44685]_ , \new_[44686]_ , \new_[44689]_ ,
    \new_[44692]_ , \new_[44693]_ , \new_[44694]_ , \new_[44698]_ ,
    \new_[44699]_ , \new_[44703]_ , \new_[44704]_ , \new_[44705]_ ,
    \new_[44709]_ , \new_[44710]_ , \new_[44713]_ , \new_[44716]_ ,
    \new_[44717]_ , \new_[44718]_ , \new_[44722]_ , \new_[44723]_ ,
    \new_[44727]_ , \new_[44728]_ , \new_[44729]_ , \new_[44733]_ ,
    \new_[44734]_ , \new_[44737]_ , \new_[44740]_ , \new_[44741]_ ,
    \new_[44742]_ , \new_[44746]_ , \new_[44747]_ , \new_[44751]_ ,
    \new_[44752]_ , \new_[44753]_ , \new_[44757]_ , \new_[44758]_ ,
    \new_[44761]_ , \new_[44764]_ , \new_[44765]_ , \new_[44766]_ ,
    \new_[44770]_ , \new_[44771]_ , \new_[44775]_ , \new_[44776]_ ,
    \new_[44777]_ , \new_[44781]_ , \new_[44782]_ , \new_[44785]_ ,
    \new_[44788]_ , \new_[44789]_ , \new_[44790]_ , \new_[44794]_ ,
    \new_[44795]_ , \new_[44799]_ , \new_[44800]_ , \new_[44801]_ ,
    \new_[44805]_ , \new_[44806]_ , \new_[44809]_ , \new_[44812]_ ,
    \new_[44813]_ , \new_[44814]_ , \new_[44818]_ , \new_[44819]_ ,
    \new_[44823]_ , \new_[44824]_ , \new_[44825]_ , \new_[44829]_ ,
    \new_[44830]_ , \new_[44833]_ , \new_[44836]_ , \new_[44837]_ ,
    \new_[44838]_ , \new_[44842]_ , \new_[44843]_ , \new_[44847]_ ,
    \new_[44848]_ , \new_[44849]_ , \new_[44853]_ , \new_[44854]_ ,
    \new_[44857]_ , \new_[44860]_ , \new_[44861]_ , \new_[44862]_ ,
    \new_[44866]_ , \new_[44867]_ , \new_[44871]_ , \new_[44872]_ ,
    \new_[44873]_ , \new_[44877]_ , \new_[44878]_ , \new_[44881]_ ,
    \new_[44884]_ , \new_[44885]_ , \new_[44886]_ , \new_[44890]_ ,
    \new_[44891]_ , \new_[44895]_ , \new_[44896]_ , \new_[44897]_ ,
    \new_[44901]_ , \new_[44902]_ , \new_[44905]_ , \new_[44908]_ ,
    \new_[44909]_ , \new_[44910]_ , \new_[44914]_ , \new_[44915]_ ,
    \new_[44919]_ , \new_[44920]_ , \new_[44921]_ , \new_[44925]_ ,
    \new_[44926]_ , \new_[44929]_ , \new_[44932]_ , \new_[44933]_ ,
    \new_[44934]_ , \new_[44938]_ , \new_[44939]_ , \new_[44943]_ ,
    \new_[44944]_ , \new_[44945]_ , \new_[44949]_ , \new_[44950]_ ,
    \new_[44953]_ , \new_[44956]_ , \new_[44957]_ , \new_[44958]_ ,
    \new_[44962]_ , \new_[44963]_ , \new_[44967]_ , \new_[44968]_ ,
    \new_[44969]_ , \new_[44973]_ , \new_[44974]_ , \new_[44977]_ ,
    \new_[44980]_ , \new_[44981]_ , \new_[44982]_ , \new_[44986]_ ,
    \new_[44987]_ , \new_[44991]_ , \new_[44992]_ , \new_[44993]_ ,
    \new_[44997]_ , \new_[44998]_ , \new_[45001]_ , \new_[45004]_ ,
    \new_[45005]_ , \new_[45006]_ , \new_[45010]_ , \new_[45011]_ ,
    \new_[45015]_ , \new_[45016]_ , \new_[45017]_ , \new_[45021]_ ,
    \new_[45022]_ , \new_[45025]_ , \new_[45028]_ , \new_[45029]_ ,
    \new_[45030]_ , \new_[45034]_ , \new_[45035]_ , \new_[45039]_ ,
    \new_[45040]_ , \new_[45041]_ , \new_[45045]_ , \new_[45046]_ ,
    \new_[45049]_ , \new_[45052]_ , \new_[45053]_ , \new_[45054]_ ,
    \new_[45058]_ , \new_[45059]_ , \new_[45063]_ , \new_[45064]_ ,
    \new_[45065]_ , \new_[45069]_ , \new_[45070]_ , \new_[45073]_ ,
    \new_[45076]_ , \new_[45077]_ , \new_[45078]_ , \new_[45082]_ ,
    \new_[45083]_ , \new_[45087]_ , \new_[45088]_ , \new_[45089]_ ,
    \new_[45093]_ , \new_[45094]_ , \new_[45097]_ , \new_[45100]_ ,
    \new_[45101]_ , \new_[45102]_ , \new_[45106]_ , \new_[45107]_ ,
    \new_[45111]_ , \new_[45112]_ , \new_[45113]_ , \new_[45117]_ ,
    \new_[45118]_ , \new_[45121]_ , \new_[45124]_ , \new_[45125]_ ,
    \new_[45126]_ , \new_[45130]_ , \new_[45131]_ , \new_[45135]_ ,
    \new_[45136]_ , \new_[45137]_ , \new_[45141]_ , \new_[45142]_ ,
    \new_[45145]_ , \new_[45148]_ , \new_[45149]_ , \new_[45150]_ ,
    \new_[45154]_ , \new_[45155]_ , \new_[45159]_ , \new_[45160]_ ,
    \new_[45161]_ , \new_[45165]_ , \new_[45166]_ , \new_[45169]_ ,
    \new_[45172]_ , \new_[45173]_ , \new_[45174]_ , \new_[45178]_ ,
    \new_[45179]_ , \new_[45183]_ , \new_[45184]_ , \new_[45185]_ ,
    \new_[45189]_ , \new_[45190]_ , \new_[45193]_ , \new_[45196]_ ,
    \new_[45197]_ , \new_[45198]_ , \new_[45202]_ , \new_[45203]_ ,
    \new_[45207]_ , \new_[45208]_ , \new_[45209]_ , \new_[45213]_ ,
    \new_[45214]_ , \new_[45217]_ , \new_[45220]_ , \new_[45221]_ ,
    \new_[45222]_ , \new_[45226]_ , \new_[45227]_ , \new_[45231]_ ,
    \new_[45232]_ , \new_[45233]_ , \new_[45237]_ , \new_[45238]_ ,
    \new_[45241]_ , \new_[45244]_ , \new_[45245]_ , \new_[45246]_ ,
    \new_[45250]_ , \new_[45251]_ , \new_[45255]_ , \new_[45256]_ ,
    \new_[45257]_ , \new_[45261]_ , \new_[45262]_ , \new_[45265]_ ,
    \new_[45268]_ , \new_[45269]_ , \new_[45270]_ , \new_[45274]_ ,
    \new_[45275]_ , \new_[45279]_ , \new_[45280]_ , \new_[45281]_ ,
    \new_[45285]_ , \new_[45286]_ , \new_[45289]_ , \new_[45292]_ ,
    \new_[45293]_ , \new_[45294]_ , \new_[45298]_ , \new_[45299]_ ,
    \new_[45303]_ , \new_[45304]_ , \new_[45305]_ , \new_[45309]_ ,
    \new_[45310]_ , \new_[45313]_ , \new_[45316]_ , \new_[45317]_ ,
    \new_[45318]_ , \new_[45322]_ , \new_[45323]_ , \new_[45327]_ ,
    \new_[45328]_ , \new_[45329]_ , \new_[45333]_ , \new_[45334]_ ,
    \new_[45337]_ , \new_[45340]_ , \new_[45341]_ , \new_[45342]_ ,
    \new_[45346]_ , \new_[45347]_ , \new_[45351]_ , \new_[45352]_ ,
    \new_[45353]_ , \new_[45357]_ , \new_[45358]_ , \new_[45361]_ ,
    \new_[45364]_ , \new_[45365]_ , \new_[45366]_ , \new_[45370]_ ,
    \new_[45371]_ , \new_[45375]_ , \new_[45376]_ , \new_[45377]_ ,
    \new_[45381]_ , \new_[45382]_ , \new_[45385]_ , \new_[45388]_ ,
    \new_[45389]_ , \new_[45390]_ , \new_[45394]_ , \new_[45395]_ ,
    \new_[45399]_ , \new_[45400]_ , \new_[45401]_ , \new_[45405]_ ,
    \new_[45406]_ , \new_[45409]_ , \new_[45412]_ , \new_[45413]_ ,
    \new_[45414]_ , \new_[45418]_ , \new_[45419]_ , \new_[45423]_ ,
    \new_[45424]_ , \new_[45425]_ , \new_[45429]_ , \new_[45430]_ ,
    \new_[45433]_ , \new_[45436]_ , \new_[45437]_ , \new_[45438]_ ,
    \new_[45442]_ , \new_[45443]_ , \new_[45447]_ , \new_[45448]_ ,
    \new_[45449]_ , \new_[45453]_ , \new_[45454]_ , \new_[45457]_ ,
    \new_[45460]_ , \new_[45461]_ , \new_[45462]_ , \new_[45466]_ ,
    \new_[45467]_ , \new_[45471]_ , \new_[45472]_ , \new_[45473]_ ,
    \new_[45477]_ , \new_[45478]_ , \new_[45481]_ , \new_[45484]_ ,
    \new_[45485]_ , \new_[45486]_ , \new_[45490]_ , \new_[45491]_ ,
    \new_[45495]_ , \new_[45496]_ , \new_[45497]_ , \new_[45501]_ ,
    \new_[45502]_ , \new_[45505]_ , \new_[45508]_ , \new_[45509]_ ,
    \new_[45510]_ , \new_[45514]_ , \new_[45515]_ , \new_[45519]_ ,
    \new_[45520]_ , \new_[45521]_ , \new_[45525]_ , \new_[45526]_ ,
    \new_[45529]_ , \new_[45532]_ , \new_[45533]_ , \new_[45534]_ ,
    \new_[45538]_ , \new_[45539]_ , \new_[45543]_ , \new_[45544]_ ,
    \new_[45545]_ , \new_[45549]_ , \new_[45550]_ , \new_[45553]_ ,
    \new_[45556]_ , \new_[45557]_ , \new_[45558]_ , \new_[45562]_ ,
    \new_[45563]_ , \new_[45567]_ , \new_[45568]_ , \new_[45569]_ ,
    \new_[45573]_ , \new_[45574]_ , \new_[45577]_ , \new_[45580]_ ,
    \new_[45581]_ , \new_[45582]_ , \new_[45586]_ , \new_[45587]_ ,
    \new_[45591]_ , \new_[45592]_ , \new_[45593]_ , \new_[45597]_ ,
    \new_[45598]_ , \new_[45601]_ , \new_[45604]_ , \new_[45605]_ ,
    \new_[45606]_ , \new_[45610]_ , \new_[45611]_ , \new_[45615]_ ,
    \new_[45616]_ , \new_[45617]_ , \new_[45621]_ , \new_[45622]_ ,
    \new_[45625]_ , \new_[45628]_ , \new_[45629]_ , \new_[45630]_ ,
    \new_[45634]_ , \new_[45635]_ , \new_[45639]_ , \new_[45640]_ ,
    \new_[45641]_ , \new_[45645]_ , \new_[45646]_ , \new_[45649]_ ,
    \new_[45652]_ , \new_[45653]_ , \new_[45654]_ , \new_[45658]_ ,
    \new_[45659]_ , \new_[45663]_ , \new_[45664]_ , \new_[45665]_ ,
    \new_[45669]_ , \new_[45670]_ , \new_[45673]_ , \new_[45676]_ ,
    \new_[45677]_ , \new_[45678]_ , \new_[45682]_ , \new_[45683]_ ,
    \new_[45687]_ , \new_[45688]_ , \new_[45689]_ , \new_[45693]_ ,
    \new_[45694]_ , \new_[45697]_ , \new_[45700]_ , \new_[45701]_ ,
    \new_[45702]_ , \new_[45706]_ , \new_[45707]_ , \new_[45711]_ ,
    \new_[45712]_ , \new_[45713]_ , \new_[45717]_ , \new_[45718]_ ,
    \new_[45721]_ , \new_[45724]_ , \new_[45725]_ , \new_[45726]_ ,
    \new_[45730]_ , \new_[45731]_ , \new_[45735]_ , \new_[45736]_ ,
    \new_[45737]_ , \new_[45741]_ , \new_[45742]_ , \new_[45745]_ ,
    \new_[45748]_ , \new_[45749]_ , \new_[45750]_ , \new_[45754]_ ,
    \new_[45755]_ , \new_[45759]_ , \new_[45760]_ , \new_[45761]_ ,
    \new_[45765]_ , \new_[45766]_ , \new_[45769]_ , \new_[45772]_ ,
    \new_[45773]_ , \new_[45774]_ , \new_[45778]_ , \new_[45779]_ ,
    \new_[45783]_ , \new_[45784]_ , \new_[45785]_ , \new_[45789]_ ,
    \new_[45790]_ , \new_[45793]_ , \new_[45796]_ , \new_[45797]_ ,
    \new_[45798]_ , \new_[45802]_ , \new_[45803]_ , \new_[45807]_ ,
    \new_[45808]_ , \new_[45809]_ , \new_[45813]_ , \new_[45814]_ ,
    \new_[45817]_ , \new_[45820]_ , \new_[45821]_ , \new_[45822]_ ,
    \new_[45826]_ , \new_[45827]_ , \new_[45831]_ , \new_[45832]_ ,
    \new_[45833]_ , \new_[45837]_ , \new_[45838]_ , \new_[45841]_ ,
    \new_[45844]_ , \new_[45845]_ , \new_[45846]_ , \new_[45850]_ ,
    \new_[45851]_ , \new_[45855]_ , \new_[45856]_ , \new_[45857]_ ,
    \new_[45861]_ , \new_[45862]_ , \new_[45865]_ , \new_[45868]_ ,
    \new_[45869]_ , \new_[45870]_ , \new_[45874]_ , \new_[45875]_ ,
    \new_[45879]_ , \new_[45880]_ , \new_[45881]_ , \new_[45885]_ ,
    \new_[45886]_ , \new_[45889]_ , \new_[45892]_ , \new_[45893]_ ,
    \new_[45894]_ , \new_[45898]_ , \new_[45899]_ , \new_[45903]_ ,
    \new_[45904]_ , \new_[45905]_ , \new_[45909]_ , \new_[45910]_ ,
    \new_[45913]_ , \new_[45916]_ , \new_[45917]_ , \new_[45918]_ ,
    \new_[45922]_ , \new_[45923]_ , \new_[45927]_ , \new_[45928]_ ,
    \new_[45929]_ , \new_[45933]_ , \new_[45934]_ , \new_[45937]_ ,
    \new_[45940]_ , \new_[45941]_ , \new_[45942]_ , \new_[45946]_ ,
    \new_[45947]_ , \new_[45951]_ , \new_[45952]_ , \new_[45953]_ ,
    \new_[45957]_ , \new_[45958]_ , \new_[45961]_ , \new_[45964]_ ,
    \new_[45965]_ , \new_[45966]_ , \new_[45970]_ , \new_[45971]_ ,
    \new_[45975]_ , \new_[45976]_ , \new_[45977]_ , \new_[45981]_ ,
    \new_[45982]_ , \new_[45985]_ , \new_[45988]_ , \new_[45989]_ ,
    \new_[45990]_ , \new_[45994]_ , \new_[45995]_ , \new_[45999]_ ,
    \new_[46000]_ , \new_[46001]_ , \new_[46005]_ , \new_[46006]_ ,
    \new_[46009]_ , \new_[46012]_ , \new_[46013]_ , \new_[46014]_ ,
    \new_[46018]_ , \new_[46019]_ , \new_[46023]_ , \new_[46024]_ ,
    \new_[46025]_ , \new_[46029]_ , \new_[46030]_ , \new_[46033]_ ,
    \new_[46036]_ , \new_[46037]_ , \new_[46038]_ , \new_[46042]_ ,
    \new_[46043]_ , \new_[46047]_ , \new_[46048]_ , \new_[46049]_ ,
    \new_[46053]_ , \new_[46054]_ , \new_[46057]_ , \new_[46060]_ ,
    \new_[46061]_ , \new_[46062]_ , \new_[46066]_ , \new_[46067]_ ,
    \new_[46071]_ , \new_[46072]_ , \new_[46073]_ , \new_[46077]_ ,
    \new_[46078]_ , \new_[46081]_ , \new_[46084]_ , \new_[46085]_ ,
    \new_[46086]_ , \new_[46090]_ , \new_[46091]_ , \new_[46095]_ ,
    \new_[46096]_ , \new_[46097]_ , \new_[46101]_ , \new_[46102]_ ,
    \new_[46105]_ , \new_[46108]_ , \new_[46109]_ , \new_[46110]_ ,
    \new_[46114]_ , \new_[46115]_ , \new_[46119]_ , \new_[46120]_ ,
    \new_[46121]_ , \new_[46125]_ , \new_[46126]_ , \new_[46129]_ ,
    \new_[46132]_ , \new_[46133]_ , \new_[46134]_ , \new_[46138]_ ,
    \new_[46139]_ , \new_[46143]_ , \new_[46144]_ , \new_[46145]_ ,
    \new_[46149]_ , \new_[46150]_ , \new_[46153]_ , \new_[46156]_ ,
    \new_[46157]_ , \new_[46158]_ , \new_[46162]_ , \new_[46163]_ ,
    \new_[46167]_ , \new_[46168]_ , \new_[46169]_ , \new_[46173]_ ,
    \new_[46174]_ , \new_[46177]_ , \new_[46180]_ , \new_[46181]_ ,
    \new_[46182]_ , \new_[46186]_ , \new_[46187]_ , \new_[46191]_ ,
    \new_[46192]_ , \new_[46193]_ , \new_[46197]_ , \new_[46198]_ ,
    \new_[46201]_ , \new_[46204]_ , \new_[46205]_ , \new_[46206]_ ,
    \new_[46210]_ , \new_[46211]_ , \new_[46215]_ , \new_[46216]_ ,
    \new_[46217]_ , \new_[46221]_ , \new_[46222]_ , \new_[46225]_ ,
    \new_[46228]_ , \new_[46229]_ , \new_[46230]_ , \new_[46234]_ ,
    \new_[46235]_ , \new_[46239]_ , \new_[46240]_ , \new_[46241]_ ,
    \new_[46245]_ , \new_[46246]_ , \new_[46249]_ , \new_[46252]_ ,
    \new_[46253]_ , \new_[46254]_ , \new_[46258]_ , \new_[46259]_ ,
    \new_[46263]_ , \new_[46264]_ , \new_[46265]_ , \new_[46269]_ ,
    \new_[46270]_ , \new_[46273]_ , \new_[46276]_ , \new_[46277]_ ,
    \new_[46278]_ , \new_[46282]_ , \new_[46283]_ , \new_[46287]_ ,
    \new_[46288]_ , \new_[46289]_ , \new_[46293]_ , \new_[46294]_ ,
    \new_[46297]_ , \new_[46300]_ , \new_[46301]_ , \new_[46302]_ ,
    \new_[46306]_ , \new_[46307]_ , \new_[46311]_ , \new_[46312]_ ,
    \new_[46313]_ , \new_[46317]_ , \new_[46318]_ , \new_[46321]_ ,
    \new_[46324]_ , \new_[46325]_ , \new_[46326]_ , \new_[46330]_ ,
    \new_[46331]_ , \new_[46335]_ , \new_[46336]_ , \new_[46337]_ ,
    \new_[46341]_ , \new_[46342]_ , \new_[46345]_ , \new_[46348]_ ,
    \new_[46349]_ , \new_[46350]_ , \new_[46354]_ , \new_[46355]_ ,
    \new_[46359]_ , \new_[46360]_ , \new_[46361]_ , \new_[46365]_ ,
    \new_[46366]_ , \new_[46369]_ , \new_[46372]_ , \new_[46373]_ ,
    \new_[46374]_ , \new_[46378]_ , \new_[46379]_ , \new_[46383]_ ,
    \new_[46384]_ , \new_[46385]_ , \new_[46389]_ , \new_[46390]_ ,
    \new_[46393]_ , \new_[46396]_ , \new_[46397]_ , \new_[46398]_ ,
    \new_[46402]_ , \new_[46403]_ , \new_[46407]_ , \new_[46408]_ ,
    \new_[46409]_ , \new_[46413]_ , \new_[46414]_ , \new_[46417]_ ,
    \new_[46420]_ , \new_[46421]_ , \new_[46422]_ , \new_[46426]_ ,
    \new_[46427]_ , \new_[46431]_ , \new_[46432]_ , \new_[46433]_ ,
    \new_[46437]_ , \new_[46438]_ , \new_[46441]_ , \new_[46444]_ ,
    \new_[46445]_ , \new_[46446]_ , \new_[46450]_ , \new_[46451]_ ,
    \new_[46455]_ , \new_[46456]_ , \new_[46457]_ , \new_[46461]_ ,
    \new_[46462]_ , \new_[46465]_ , \new_[46468]_ , \new_[46469]_ ,
    \new_[46470]_ , \new_[46474]_ , \new_[46475]_ , \new_[46479]_ ,
    \new_[46480]_ , \new_[46481]_ , \new_[46485]_ , \new_[46486]_ ,
    \new_[46489]_ , \new_[46492]_ , \new_[46493]_ , \new_[46494]_ ,
    \new_[46498]_ , \new_[46499]_ , \new_[46503]_ , \new_[46504]_ ,
    \new_[46505]_ , \new_[46509]_ , \new_[46510]_ , \new_[46513]_ ,
    \new_[46516]_ , \new_[46517]_ , \new_[46518]_ , \new_[46522]_ ,
    \new_[46523]_ , \new_[46527]_ , \new_[46528]_ , \new_[46529]_ ,
    \new_[46533]_ , \new_[46534]_ , \new_[46537]_ , \new_[46540]_ ,
    \new_[46541]_ , \new_[46542]_ , \new_[46546]_ , \new_[46547]_ ,
    \new_[46551]_ , \new_[46552]_ , \new_[46553]_ , \new_[46557]_ ,
    \new_[46558]_ , \new_[46561]_ , \new_[46564]_ , \new_[46565]_ ,
    \new_[46566]_ , \new_[46570]_ , \new_[46571]_ , \new_[46575]_ ,
    \new_[46576]_ , \new_[46577]_ , \new_[46581]_ , \new_[46582]_ ,
    \new_[46585]_ , \new_[46588]_ , \new_[46589]_ , \new_[46590]_ ,
    \new_[46594]_ , \new_[46595]_ , \new_[46599]_ , \new_[46600]_ ,
    \new_[46601]_ , \new_[46605]_ , \new_[46606]_ , \new_[46609]_ ,
    \new_[46612]_ , \new_[46613]_ , \new_[46614]_ , \new_[46618]_ ,
    \new_[46619]_ , \new_[46623]_ , \new_[46624]_ , \new_[46625]_ ,
    \new_[46629]_ , \new_[46630]_ , \new_[46633]_ , \new_[46636]_ ,
    \new_[46637]_ , \new_[46638]_ , \new_[46642]_ , \new_[46643]_ ,
    \new_[46647]_ , \new_[46648]_ , \new_[46649]_ , \new_[46653]_ ,
    \new_[46654]_ , \new_[46657]_ , \new_[46660]_ , \new_[46661]_ ,
    \new_[46662]_ , \new_[46666]_ , \new_[46667]_ , \new_[46671]_ ,
    \new_[46672]_ , \new_[46673]_ , \new_[46677]_ , \new_[46678]_ ,
    \new_[46681]_ , \new_[46684]_ , \new_[46685]_ , \new_[46686]_ ,
    \new_[46690]_ , \new_[46691]_ , \new_[46695]_ , \new_[46696]_ ,
    \new_[46697]_ , \new_[46701]_ , \new_[46702]_ , \new_[46705]_ ,
    \new_[46708]_ , \new_[46709]_ , \new_[46710]_ , \new_[46714]_ ,
    \new_[46715]_ , \new_[46719]_ , \new_[46720]_ , \new_[46721]_ ,
    \new_[46725]_ , \new_[46726]_ , \new_[46729]_ , \new_[46732]_ ,
    \new_[46733]_ , \new_[46734]_ , \new_[46738]_ , \new_[46739]_ ,
    \new_[46743]_ , \new_[46744]_ , \new_[46745]_ , \new_[46749]_ ,
    \new_[46750]_ , \new_[46753]_ , \new_[46756]_ , \new_[46757]_ ,
    \new_[46758]_ , \new_[46762]_ , \new_[46763]_ , \new_[46767]_ ,
    \new_[46768]_ , \new_[46769]_ , \new_[46773]_ , \new_[46774]_ ,
    \new_[46777]_ , \new_[46780]_ , \new_[46781]_ , \new_[46782]_ ,
    \new_[46786]_ , \new_[46787]_ , \new_[46791]_ , \new_[46792]_ ,
    \new_[46793]_ , \new_[46797]_ , \new_[46798]_ , \new_[46801]_ ,
    \new_[46804]_ , \new_[46805]_ , \new_[46806]_ , \new_[46810]_ ,
    \new_[46811]_ , \new_[46815]_ , \new_[46816]_ , \new_[46817]_ ,
    \new_[46821]_ , \new_[46822]_ , \new_[46825]_ , \new_[46828]_ ,
    \new_[46829]_ , \new_[46830]_ , \new_[46834]_ , \new_[46835]_ ,
    \new_[46839]_ , \new_[46840]_ , \new_[46841]_ , \new_[46845]_ ,
    \new_[46846]_ , \new_[46849]_ , \new_[46852]_ , \new_[46853]_ ,
    \new_[46854]_ , \new_[46858]_ , \new_[46859]_ , \new_[46863]_ ,
    \new_[46864]_ , \new_[46865]_ , \new_[46869]_ , \new_[46870]_ ,
    \new_[46873]_ , \new_[46876]_ , \new_[46877]_ , \new_[46878]_ ,
    \new_[46882]_ , \new_[46883]_ , \new_[46887]_ , \new_[46888]_ ,
    \new_[46889]_ , \new_[46893]_ , \new_[46894]_ , \new_[46897]_ ,
    \new_[46900]_ , \new_[46901]_ , \new_[46902]_ , \new_[46906]_ ,
    \new_[46907]_ , \new_[46911]_ , \new_[46912]_ , \new_[46913]_ ,
    \new_[46917]_ , \new_[46918]_ , \new_[46921]_ , \new_[46924]_ ,
    \new_[46925]_ , \new_[46926]_ , \new_[46930]_ , \new_[46931]_ ,
    \new_[46935]_ , \new_[46936]_ , \new_[46937]_ , \new_[46941]_ ,
    \new_[46942]_ , \new_[46945]_ , \new_[46948]_ , \new_[46949]_ ,
    \new_[46950]_ , \new_[46954]_ , \new_[46955]_ , \new_[46959]_ ,
    \new_[46960]_ , \new_[46961]_ , \new_[46965]_ , \new_[46966]_ ,
    \new_[46969]_ , \new_[46972]_ , \new_[46973]_ , \new_[46974]_ ,
    \new_[46978]_ , \new_[46979]_ , \new_[46983]_ , \new_[46984]_ ,
    \new_[46985]_ , \new_[46989]_ , \new_[46990]_ , \new_[46993]_ ,
    \new_[46996]_ , \new_[46997]_ , \new_[46998]_ , \new_[47002]_ ,
    \new_[47003]_ , \new_[47007]_ , \new_[47008]_ , \new_[47009]_ ,
    \new_[47013]_ , \new_[47014]_ , \new_[47017]_ , \new_[47020]_ ,
    \new_[47021]_ , \new_[47022]_ , \new_[47026]_ , \new_[47027]_ ,
    \new_[47031]_ , \new_[47032]_ , \new_[47033]_ , \new_[47037]_ ,
    \new_[47038]_ , \new_[47041]_ , \new_[47044]_ , \new_[47045]_ ,
    \new_[47046]_ , \new_[47050]_ , \new_[47051]_ , \new_[47055]_ ,
    \new_[47056]_ , \new_[47057]_ , \new_[47061]_ , \new_[47062]_ ,
    \new_[47065]_ , \new_[47068]_ , \new_[47069]_ , \new_[47070]_ ,
    \new_[47074]_ , \new_[47075]_ , \new_[47079]_ , \new_[47080]_ ,
    \new_[47081]_ , \new_[47085]_ , \new_[47086]_ , \new_[47089]_ ,
    \new_[47092]_ , \new_[47093]_ , \new_[47094]_ , \new_[47098]_ ,
    \new_[47099]_ , \new_[47103]_ , \new_[47104]_ , \new_[47105]_ ,
    \new_[47109]_ , \new_[47110]_ , \new_[47113]_ , \new_[47116]_ ,
    \new_[47117]_ , \new_[47118]_ , \new_[47122]_ , \new_[47123]_ ,
    \new_[47127]_ , \new_[47128]_ , \new_[47129]_ , \new_[47133]_ ,
    \new_[47134]_ , \new_[47137]_ , \new_[47140]_ , \new_[47141]_ ,
    \new_[47142]_ , \new_[47146]_ , \new_[47147]_ , \new_[47151]_ ,
    \new_[47152]_ , \new_[47153]_ , \new_[47157]_ , \new_[47158]_ ,
    \new_[47161]_ , \new_[47164]_ , \new_[47165]_ , \new_[47166]_ ,
    \new_[47170]_ , \new_[47171]_ , \new_[47175]_ , \new_[47176]_ ,
    \new_[47177]_ , \new_[47181]_ , \new_[47182]_ , \new_[47185]_ ,
    \new_[47188]_ , \new_[47189]_ , \new_[47190]_ , \new_[47194]_ ,
    \new_[47195]_ , \new_[47199]_ , \new_[47200]_ , \new_[47201]_ ,
    \new_[47205]_ , \new_[47206]_ , \new_[47209]_ , \new_[47212]_ ,
    \new_[47213]_ , \new_[47214]_ , \new_[47218]_ , \new_[47219]_ ,
    \new_[47223]_ , \new_[47224]_ , \new_[47225]_ , \new_[47229]_ ,
    \new_[47230]_ , \new_[47233]_ , \new_[47236]_ , \new_[47237]_ ,
    \new_[47238]_ , \new_[47242]_ , \new_[47243]_ , \new_[47247]_ ,
    \new_[47248]_ , \new_[47249]_ , \new_[47253]_ , \new_[47254]_ ,
    \new_[47257]_ , \new_[47260]_ , \new_[47261]_ , \new_[47262]_ ,
    \new_[47266]_ , \new_[47267]_ , \new_[47271]_ , \new_[47272]_ ,
    \new_[47273]_ , \new_[47277]_ , \new_[47278]_ , \new_[47281]_ ,
    \new_[47284]_ , \new_[47285]_ , \new_[47286]_ , \new_[47290]_ ,
    \new_[47291]_ , \new_[47295]_ , \new_[47296]_ , \new_[47297]_ ,
    \new_[47301]_ , \new_[47302]_ , \new_[47305]_ , \new_[47308]_ ,
    \new_[47309]_ , \new_[47310]_ , \new_[47314]_ , \new_[47315]_ ,
    \new_[47319]_ , \new_[47320]_ , \new_[47321]_ , \new_[47325]_ ,
    \new_[47326]_ , \new_[47329]_ , \new_[47332]_ , \new_[47333]_ ,
    \new_[47334]_ , \new_[47338]_ , \new_[47339]_ , \new_[47343]_ ,
    \new_[47344]_ , \new_[47345]_ , \new_[47349]_ , \new_[47350]_ ,
    \new_[47353]_ , \new_[47356]_ , \new_[47357]_ , \new_[47358]_ ,
    \new_[47362]_ , \new_[47363]_ , \new_[47367]_ , \new_[47368]_ ,
    \new_[47369]_ , \new_[47373]_ , \new_[47374]_ , \new_[47377]_ ,
    \new_[47380]_ , \new_[47381]_ , \new_[47382]_ , \new_[47386]_ ,
    \new_[47387]_ , \new_[47391]_ , \new_[47392]_ , \new_[47393]_ ,
    \new_[47397]_ , \new_[47398]_ , \new_[47401]_ , \new_[47404]_ ,
    \new_[47405]_ , \new_[47406]_ , \new_[47410]_ , \new_[47411]_ ,
    \new_[47415]_ , \new_[47416]_ , \new_[47417]_ , \new_[47421]_ ,
    \new_[47422]_ , \new_[47425]_ , \new_[47428]_ , \new_[47429]_ ,
    \new_[47430]_ , \new_[47434]_ , \new_[47435]_ , \new_[47439]_ ,
    \new_[47440]_ , \new_[47441]_ , \new_[47445]_ , \new_[47446]_ ,
    \new_[47449]_ , \new_[47452]_ , \new_[47453]_ , \new_[47454]_ ,
    \new_[47458]_ , \new_[47459]_ , \new_[47463]_ , \new_[47464]_ ,
    \new_[47465]_ , \new_[47469]_ , \new_[47470]_ , \new_[47473]_ ,
    \new_[47476]_ , \new_[47477]_ , \new_[47478]_ , \new_[47482]_ ,
    \new_[47483]_ , \new_[47487]_ , \new_[47488]_ , \new_[47489]_ ,
    \new_[47493]_ , \new_[47494]_ , \new_[47497]_ , \new_[47500]_ ,
    \new_[47501]_ , \new_[47502]_ , \new_[47506]_ , \new_[47507]_ ,
    \new_[47511]_ , \new_[47512]_ , \new_[47513]_ , \new_[47517]_ ,
    \new_[47518]_ , \new_[47521]_ , \new_[47524]_ , \new_[47525]_ ,
    \new_[47526]_ , \new_[47530]_ , \new_[47531]_ , \new_[47535]_ ,
    \new_[47536]_ , \new_[47537]_ , \new_[47541]_ , \new_[47542]_ ,
    \new_[47545]_ , \new_[47548]_ , \new_[47549]_ , \new_[47550]_ ,
    \new_[47554]_ , \new_[47555]_ , \new_[47559]_ , \new_[47560]_ ,
    \new_[47561]_ , \new_[47565]_ , \new_[47566]_ , \new_[47569]_ ,
    \new_[47572]_ , \new_[47573]_ , \new_[47574]_ , \new_[47578]_ ,
    \new_[47579]_ , \new_[47583]_ , \new_[47584]_ , \new_[47585]_ ,
    \new_[47589]_ , \new_[47590]_ , \new_[47593]_ , \new_[47596]_ ,
    \new_[47597]_ , \new_[47598]_ , \new_[47602]_ , \new_[47603]_ ,
    \new_[47607]_ , \new_[47608]_ , \new_[47609]_ , \new_[47613]_ ,
    \new_[47614]_ , \new_[47617]_ , \new_[47620]_ , \new_[47621]_ ,
    \new_[47622]_ , \new_[47626]_ , \new_[47627]_ , \new_[47631]_ ,
    \new_[47632]_ , \new_[47633]_ , \new_[47637]_ , \new_[47638]_ ,
    \new_[47641]_ , \new_[47644]_ , \new_[47645]_ , \new_[47646]_ ,
    \new_[47650]_ , \new_[47651]_ , \new_[47655]_ , \new_[47656]_ ,
    \new_[47657]_ , \new_[47661]_ , \new_[47662]_ , \new_[47665]_ ,
    \new_[47668]_ , \new_[47669]_ , \new_[47670]_ , \new_[47674]_ ,
    \new_[47675]_ , \new_[47679]_ , \new_[47680]_ , \new_[47681]_ ,
    \new_[47685]_ , \new_[47686]_ , \new_[47689]_ , \new_[47692]_ ,
    \new_[47693]_ , \new_[47694]_ , \new_[47698]_ , \new_[47699]_ ,
    \new_[47703]_ , \new_[47704]_ , \new_[47705]_ , \new_[47709]_ ,
    \new_[47710]_ , \new_[47713]_ , \new_[47716]_ , \new_[47717]_ ,
    \new_[47718]_ , \new_[47722]_ , \new_[47723]_ , \new_[47727]_ ,
    \new_[47728]_ , \new_[47729]_ , \new_[47733]_ , \new_[47734]_ ,
    \new_[47737]_ , \new_[47740]_ , \new_[47741]_ , \new_[47742]_ ,
    \new_[47746]_ , \new_[47747]_ , \new_[47751]_ , \new_[47752]_ ,
    \new_[47753]_ , \new_[47757]_ , \new_[47758]_ , \new_[47761]_ ,
    \new_[47764]_ , \new_[47765]_ , \new_[47766]_ , \new_[47770]_ ,
    \new_[47771]_ , \new_[47775]_ , \new_[47776]_ , \new_[47777]_ ,
    \new_[47781]_ , \new_[47782]_ , \new_[47785]_ , \new_[47788]_ ,
    \new_[47789]_ , \new_[47790]_ , \new_[47794]_ , \new_[47795]_ ,
    \new_[47799]_ , \new_[47800]_ , \new_[47801]_ , \new_[47805]_ ,
    \new_[47806]_ , \new_[47809]_ , \new_[47812]_ , \new_[47813]_ ,
    \new_[47814]_ , \new_[47818]_ , \new_[47819]_ , \new_[47823]_ ,
    \new_[47824]_ , \new_[47825]_ , \new_[47829]_ , \new_[47830]_ ,
    \new_[47833]_ , \new_[47836]_ , \new_[47837]_ , \new_[47838]_ ,
    \new_[47842]_ , \new_[47843]_ , \new_[47847]_ , \new_[47848]_ ,
    \new_[47849]_ , \new_[47853]_ , \new_[47854]_ , \new_[47857]_ ,
    \new_[47860]_ , \new_[47861]_ , \new_[47862]_ , \new_[47866]_ ,
    \new_[47867]_ , \new_[47871]_ , \new_[47872]_ , \new_[47873]_ ,
    \new_[47877]_ , \new_[47878]_ , \new_[47881]_ , \new_[47884]_ ,
    \new_[47885]_ , \new_[47886]_ , \new_[47890]_ , \new_[47891]_ ,
    \new_[47895]_ , \new_[47896]_ , \new_[47897]_ , \new_[47901]_ ,
    \new_[47902]_ , \new_[47905]_ , \new_[47908]_ , \new_[47909]_ ,
    \new_[47910]_ , \new_[47914]_ , \new_[47915]_ , \new_[47919]_ ,
    \new_[47920]_ , \new_[47921]_ , \new_[47925]_ , \new_[47926]_ ,
    \new_[47929]_ , \new_[47932]_ , \new_[47933]_ , \new_[47934]_ ,
    \new_[47938]_ , \new_[47939]_ , \new_[47943]_ , \new_[47944]_ ,
    \new_[47945]_ , \new_[47949]_ , \new_[47950]_ , \new_[47953]_ ,
    \new_[47956]_ , \new_[47957]_ , \new_[47958]_ , \new_[47962]_ ,
    \new_[47963]_ , \new_[47967]_ , \new_[47968]_ , \new_[47969]_ ,
    \new_[47973]_ , \new_[47974]_ , \new_[47977]_ , \new_[47980]_ ,
    \new_[47981]_ , \new_[47982]_ , \new_[47986]_ , \new_[47987]_ ,
    \new_[47991]_ , \new_[47992]_ , \new_[47993]_ , \new_[47997]_ ,
    \new_[47998]_ , \new_[48001]_ , \new_[48004]_ , \new_[48005]_ ,
    \new_[48006]_ , \new_[48010]_ , \new_[48011]_ , \new_[48015]_ ,
    \new_[48016]_ , \new_[48017]_ , \new_[48021]_ , \new_[48022]_ ,
    \new_[48025]_ , \new_[48028]_ , \new_[48029]_ , \new_[48030]_ ,
    \new_[48034]_ , \new_[48035]_ , \new_[48039]_ , \new_[48040]_ ,
    \new_[48041]_ , \new_[48045]_ , \new_[48046]_ , \new_[48049]_ ,
    \new_[48052]_ , \new_[48053]_ , \new_[48054]_ , \new_[48058]_ ,
    \new_[48059]_ , \new_[48063]_ , \new_[48064]_ , \new_[48065]_ ,
    \new_[48069]_ , \new_[48070]_ , \new_[48073]_ , \new_[48076]_ ,
    \new_[48077]_ , \new_[48078]_ , \new_[48082]_ , \new_[48083]_ ,
    \new_[48087]_ , \new_[48088]_ , \new_[48089]_ , \new_[48093]_ ,
    \new_[48094]_ , \new_[48097]_ , \new_[48100]_ , \new_[48101]_ ,
    \new_[48102]_ , \new_[48106]_ , \new_[48107]_ , \new_[48111]_ ,
    \new_[48112]_ , \new_[48113]_ , \new_[48117]_ , \new_[48118]_ ,
    \new_[48121]_ , \new_[48124]_ , \new_[48125]_ , \new_[48126]_ ,
    \new_[48130]_ , \new_[48131]_ , \new_[48135]_ , \new_[48136]_ ,
    \new_[48137]_ , \new_[48141]_ , \new_[48142]_ , \new_[48145]_ ,
    \new_[48148]_ , \new_[48149]_ , \new_[48150]_ , \new_[48154]_ ,
    \new_[48155]_ , \new_[48159]_ , \new_[48160]_ , \new_[48161]_ ,
    \new_[48165]_ , \new_[48166]_ , \new_[48169]_ , \new_[48172]_ ,
    \new_[48173]_ , \new_[48174]_ , \new_[48178]_ , \new_[48179]_ ,
    \new_[48183]_ , \new_[48184]_ , \new_[48185]_ , \new_[48189]_ ,
    \new_[48190]_ , \new_[48193]_ , \new_[48196]_ , \new_[48197]_ ,
    \new_[48198]_ , \new_[48202]_ , \new_[48203]_ , \new_[48207]_ ,
    \new_[48208]_ , \new_[48209]_ , \new_[48213]_ , \new_[48214]_ ,
    \new_[48217]_ , \new_[48220]_ , \new_[48221]_ , \new_[48222]_ ,
    \new_[48226]_ , \new_[48227]_ , \new_[48231]_ , \new_[48232]_ ,
    \new_[48233]_ , \new_[48237]_ , \new_[48238]_ , \new_[48241]_ ,
    \new_[48244]_ , \new_[48245]_ , \new_[48246]_ , \new_[48250]_ ,
    \new_[48251]_ , \new_[48255]_ , \new_[48256]_ , \new_[48257]_ ,
    \new_[48261]_ , \new_[48262]_ , \new_[48265]_ , \new_[48268]_ ,
    \new_[48269]_ , \new_[48270]_ , \new_[48274]_ , \new_[48275]_ ,
    \new_[48279]_ , \new_[48280]_ , \new_[48281]_ , \new_[48285]_ ,
    \new_[48286]_ , \new_[48289]_ , \new_[48292]_ , \new_[48293]_ ,
    \new_[48294]_ , \new_[48298]_ , \new_[48299]_ , \new_[48303]_ ,
    \new_[48304]_ , \new_[48305]_ , \new_[48309]_ , \new_[48310]_ ,
    \new_[48313]_ , \new_[48316]_ , \new_[48317]_ , \new_[48318]_ ,
    \new_[48322]_ , \new_[48323]_ , \new_[48327]_ , \new_[48328]_ ,
    \new_[48329]_ , \new_[48333]_ , \new_[48334]_ , \new_[48337]_ ,
    \new_[48340]_ , \new_[48341]_ , \new_[48342]_ , \new_[48346]_ ,
    \new_[48347]_ , \new_[48351]_ , \new_[48352]_ , \new_[48353]_ ,
    \new_[48357]_ , \new_[48358]_ , \new_[48361]_ , \new_[48364]_ ,
    \new_[48365]_ , \new_[48366]_ , \new_[48370]_ , \new_[48371]_ ,
    \new_[48375]_ , \new_[48376]_ , \new_[48377]_ , \new_[48381]_ ,
    \new_[48382]_ , \new_[48385]_ , \new_[48388]_ , \new_[48389]_ ,
    \new_[48390]_ , \new_[48394]_ , \new_[48395]_ , \new_[48399]_ ,
    \new_[48400]_ , \new_[48401]_ , \new_[48405]_ , \new_[48406]_ ,
    \new_[48409]_ , \new_[48412]_ , \new_[48413]_ , \new_[48414]_ ,
    \new_[48418]_ , \new_[48419]_ , \new_[48423]_ , \new_[48424]_ ,
    \new_[48425]_ , \new_[48429]_ , \new_[48430]_ , \new_[48433]_ ,
    \new_[48436]_ , \new_[48437]_ , \new_[48438]_ , \new_[48442]_ ,
    \new_[48443]_ , \new_[48447]_ , \new_[48448]_ , \new_[48449]_ ,
    \new_[48453]_ , \new_[48454]_ , \new_[48457]_ , \new_[48460]_ ,
    \new_[48461]_ , \new_[48462]_ , \new_[48466]_ , \new_[48467]_ ,
    \new_[48471]_ , \new_[48472]_ , \new_[48473]_ , \new_[48477]_ ,
    \new_[48478]_ , \new_[48481]_ , \new_[48484]_ , \new_[48485]_ ,
    \new_[48486]_ , \new_[48490]_ , \new_[48491]_ , \new_[48495]_ ,
    \new_[48496]_ , \new_[48497]_ , \new_[48501]_ , \new_[48502]_ ,
    \new_[48505]_ , \new_[48508]_ , \new_[48509]_ , \new_[48510]_ ,
    \new_[48514]_ , \new_[48515]_ , \new_[48519]_ , \new_[48520]_ ,
    \new_[48521]_ , \new_[48525]_ , \new_[48526]_ , \new_[48529]_ ,
    \new_[48532]_ , \new_[48533]_ , \new_[48534]_ , \new_[48538]_ ,
    \new_[48539]_ , \new_[48543]_ , \new_[48544]_ , \new_[48545]_ ,
    \new_[48549]_ , \new_[48550]_ , \new_[48553]_ , \new_[48556]_ ,
    \new_[48557]_ , \new_[48558]_ , \new_[48562]_ , \new_[48563]_ ,
    \new_[48567]_ , \new_[48568]_ , \new_[48569]_ , \new_[48573]_ ,
    \new_[48574]_ , \new_[48577]_ , \new_[48580]_ , \new_[48581]_ ,
    \new_[48582]_ , \new_[48586]_ , \new_[48587]_ , \new_[48591]_ ,
    \new_[48592]_ , \new_[48593]_ , \new_[48597]_ , \new_[48598]_ ,
    \new_[48601]_ , \new_[48604]_ , \new_[48605]_ , \new_[48606]_ ,
    \new_[48610]_ , \new_[48611]_ , \new_[48615]_ , \new_[48616]_ ,
    \new_[48617]_ , \new_[48621]_ , \new_[48622]_ , \new_[48625]_ ,
    \new_[48628]_ , \new_[48629]_ , \new_[48630]_ , \new_[48634]_ ,
    \new_[48635]_ , \new_[48639]_ , \new_[48640]_ , \new_[48641]_ ,
    \new_[48645]_ , \new_[48646]_ , \new_[48649]_ , \new_[48652]_ ,
    \new_[48653]_ , \new_[48654]_ , \new_[48658]_ , \new_[48659]_ ,
    \new_[48663]_ , \new_[48664]_ , \new_[48665]_ , \new_[48669]_ ,
    \new_[48670]_ , \new_[48673]_ , \new_[48676]_ , \new_[48677]_ ,
    \new_[48678]_ , \new_[48682]_ , \new_[48683]_ , \new_[48687]_ ,
    \new_[48688]_ , \new_[48689]_ , \new_[48693]_ , \new_[48694]_ ,
    \new_[48697]_ , \new_[48700]_ , \new_[48701]_ , \new_[48702]_ ,
    \new_[48706]_ , \new_[48707]_ , \new_[48711]_ , \new_[48712]_ ,
    \new_[48713]_ , \new_[48717]_ , \new_[48718]_ , \new_[48721]_ ,
    \new_[48724]_ , \new_[48725]_ , \new_[48726]_ , \new_[48730]_ ,
    \new_[48731]_ , \new_[48735]_ , \new_[48736]_ , \new_[48737]_ ,
    \new_[48741]_ , \new_[48742]_ , \new_[48745]_ , \new_[48748]_ ,
    \new_[48749]_ , \new_[48750]_ , \new_[48754]_ , \new_[48755]_ ,
    \new_[48759]_ , \new_[48760]_ , \new_[48761]_ , \new_[48765]_ ,
    \new_[48766]_ , \new_[48769]_ , \new_[48772]_ , \new_[48773]_ ,
    \new_[48774]_ , \new_[48778]_ , \new_[48779]_ , \new_[48783]_ ,
    \new_[48784]_ , \new_[48785]_ , \new_[48789]_ , \new_[48790]_ ,
    \new_[48793]_ , \new_[48796]_ , \new_[48797]_ , \new_[48798]_ ,
    \new_[48802]_ , \new_[48803]_ , \new_[48807]_ , \new_[48808]_ ,
    \new_[48809]_ , \new_[48813]_ , \new_[48814]_ , \new_[48817]_ ,
    \new_[48820]_ , \new_[48821]_ , \new_[48822]_ , \new_[48826]_ ,
    \new_[48827]_ , \new_[48831]_ , \new_[48832]_ , \new_[48833]_ ,
    \new_[48837]_ , \new_[48838]_ , \new_[48841]_ , \new_[48844]_ ,
    \new_[48845]_ , \new_[48846]_ , \new_[48850]_ , \new_[48851]_ ,
    \new_[48855]_ , \new_[48856]_ , \new_[48857]_ , \new_[48861]_ ,
    \new_[48862]_ , \new_[48865]_ , \new_[48868]_ , \new_[48869]_ ,
    \new_[48870]_ , \new_[48874]_ , \new_[48875]_ , \new_[48879]_ ,
    \new_[48880]_ , \new_[48881]_ , \new_[48885]_ , \new_[48886]_ ,
    \new_[48889]_ , \new_[48892]_ , \new_[48893]_ , \new_[48894]_ ,
    \new_[48898]_ , \new_[48899]_ , \new_[48903]_ , \new_[48904]_ ,
    \new_[48905]_ , \new_[48909]_ , \new_[48910]_ , \new_[48913]_ ,
    \new_[48916]_ , \new_[48917]_ , \new_[48918]_ , \new_[48922]_ ,
    \new_[48923]_ , \new_[48927]_ , \new_[48928]_ , \new_[48929]_ ,
    \new_[48933]_ , \new_[48934]_ , \new_[48937]_ , \new_[48940]_ ,
    \new_[48941]_ , \new_[48942]_ , \new_[48946]_ , \new_[48947]_ ,
    \new_[48951]_ , \new_[48952]_ , \new_[48953]_ , \new_[48957]_ ,
    \new_[48958]_ , \new_[48961]_ , \new_[48964]_ , \new_[48965]_ ,
    \new_[48966]_ , \new_[48970]_ , \new_[48971]_ , \new_[48975]_ ,
    \new_[48976]_ , \new_[48977]_ , \new_[48981]_ , \new_[48982]_ ,
    \new_[48985]_ , \new_[48988]_ , \new_[48989]_ , \new_[48990]_ ,
    \new_[48994]_ , \new_[48995]_ , \new_[48999]_ , \new_[49000]_ ,
    \new_[49001]_ , \new_[49005]_ , \new_[49006]_ , \new_[49009]_ ,
    \new_[49012]_ , \new_[49013]_ , \new_[49014]_ , \new_[49018]_ ,
    \new_[49019]_ , \new_[49023]_ , \new_[49024]_ , \new_[49025]_ ,
    \new_[49029]_ , \new_[49030]_ , \new_[49033]_ , \new_[49036]_ ,
    \new_[49037]_ , \new_[49038]_ , \new_[49042]_ , \new_[49043]_ ,
    \new_[49047]_ , \new_[49048]_ , \new_[49049]_ , \new_[49053]_ ,
    \new_[49054]_ , \new_[49057]_ , \new_[49060]_ , \new_[49061]_ ,
    \new_[49062]_ , \new_[49066]_ , \new_[49067]_ , \new_[49071]_ ,
    \new_[49072]_ , \new_[49073]_ , \new_[49077]_ , \new_[49078]_ ,
    \new_[49081]_ , \new_[49084]_ , \new_[49085]_ , \new_[49086]_ ,
    \new_[49090]_ , \new_[49091]_ , \new_[49095]_ , \new_[49096]_ ,
    \new_[49097]_ , \new_[49101]_ , \new_[49102]_ , \new_[49105]_ ,
    \new_[49108]_ , \new_[49109]_ , \new_[49110]_ , \new_[49114]_ ,
    \new_[49115]_ , \new_[49119]_ , \new_[49120]_ , \new_[49121]_ ,
    \new_[49125]_ , \new_[49126]_ , \new_[49129]_ , \new_[49132]_ ,
    \new_[49133]_ , \new_[49134]_ , \new_[49138]_ , \new_[49139]_ ,
    \new_[49143]_ , \new_[49144]_ , \new_[49145]_ , \new_[49149]_ ,
    \new_[49150]_ , \new_[49153]_ , \new_[49156]_ , \new_[49157]_ ,
    \new_[49158]_ , \new_[49162]_ , \new_[49163]_ , \new_[49167]_ ,
    \new_[49168]_ , \new_[49169]_ , \new_[49173]_ , \new_[49174]_ ,
    \new_[49177]_ , \new_[49180]_ , \new_[49181]_ , \new_[49182]_ ,
    \new_[49186]_ , \new_[49187]_ , \new_[49191]_ , \new_[49192]_ ,
    \new_[49193]_ , \new_[49197]_ , \new_[49198]_ , \new_[49201]_ ,
    \new_[49204]_ , \new_[49205]_ , \new_[49206]_ , \new_[49210]_ ,
    \new_[49211]_ , \new_[49215]_ , \new_[49216]_ , \new_[49217]_ ,
    \new_[49221]_ , \new_[49222]_ , \new_[49225]_ , \new_[49228]_ ,
    \new_[49229]_ , \new_[49230]_ , \new_[49234]_ , \new_[49235]_ ,
    \new_[49239]_ , \new_[49240]_ , \new_[49241]_ , \new_[49245]_ ,
    \new_[49246]_ , \new_[49249]_ , \new_[49252]_ , \new_[49253]_ ,
    \new_[49254]_ , \new_[49258]_ , \new_[49259]_ , \new_[49263]_ ,
    \new_[49264]_ , \new_[49265]_ , \new_[49269]_ , \new_[49270]_ ,
    \new_[49273]_ , \new_[49276]_ , \new_[49277]_ , \new_[49278]_ ,
    \new_[49282]_ , \new_[49283]_ , \new_[49287]_ , \new_[49288]_ ,
    \new_[49289]_ , \new_[49293]_ , \new_[49294]_ , \new_[49297]_ ,
    \new_[49300]_ , \new_[49301]_ , \new_[49302]_ , \new_[49306]_ ,
    \new_[49307]_ , \new_[49311]_ , \new_[49312]_ , \new_[49313]_ ,
    \new_[49317]_ , \new_[49318]_ , \new_[49321]_ , \new_[49324]_ ,
    \new_[49325]_ , \new_[49326]_ , \new_[49330]_ , \new_[49331]_ ,
    \new_[49335]_ , \new_[49336]_ , \new_[49337]_ , \new_[49341]_ ,
    \new_[49342]_ , \new_[49345]_ , \new_[49348]_ , \new_[49349]_ ,
    \new_[49350]_ , \new_[49354]_ , \new_[49355]_ , \new_[49359]_ ,
    \new_[49360]_ , \new_[49361]_ , \new_[49365]_ , \new_[49366]_ ,
    \new_[49369]_ , \new_[49372]_ , \new_[49373]_ , \new_[49374]_ ,
    \new_[49378]_ , \new_[49379]_ , \new_[49383]_ , \new_[49384]_ ,
    \new_[49385]_ , \new_[49389]_ , \new_[49390]_ , \new_[49393]_ ,
    \new_[49396]_ , \new_[49397]_ , \new_[49398]_ , \new_[49402]_ ,
    \new_[49403]_ , \new_[49407]_ , \new_[49408]_ , \new_[49409]_ ,
    \new_[49413]_ , \new_[49414]_ , \new_[49417]_ , \new_[49420]_ ,
    \new_[49421]_ , \new_[49422]_ , \new_[49426]_ , \new_[49427]_ ,
    \new_[49431]_ , \new_[49432]_ , \new_[49433]_ , \new_[49437]_ ,
    \new_[49438]_ , \new_[49441]_ , \new_[49444]_ , \new_[49445]_ ,
    \new_[49446]_ , \new_[49450]_ , \new_[49451]_ , \new_[49455]_ ,
    \new_[49456]_ , \new_[49457]_ , \new_[49461]_ , \new_[49462]_ ,
    \new_[49465]_ , \new_[49468]_ , \new_[49469]_ , \new_[49470]_ ,
    \new_[49474]_ , \new_[49475]_ , \new_[49479]_ , \new_[49480]_ ,
    \new_[49481]_ , \new_[49485]_ , \new_[49486]_ , \new_[49489]_ ,
    \new_[49492]_ , \new_[49493]_ , \new_[49494]_ , \new_[49498]_ ,
    \new_[49499]_ , \new_[49503]_ , \new_[49504]_ , \new_[49505]_ ,
    \new_[49509]_ , \new_[49510]_ , \new_[49513]_ , \new_[49516]_ ,
    \new_[49517]_ , \new_[49518]_ , \new_[49522]_ , \new_[49523]_ ,
    \new_[49527]_ , \new_[49528]_ , \new_[49529]_ , \new_[49533]_ ,
    \new_[49534]_ , \new_[49537]_ , \new_[49540]_ , \new_[49541]_ ,
    \new_[49542]_ , \new_[49546]_ , \new_[49547]_ , \new_[49551]_ ,
    \new_[49552]_ , \new_[49553]_ , \new_[49557]_ , \new_[49558]_ ,
    \new_[49561]_ , \new_[49564]_ , \new_[49565]_ , \new_[49566]_ ,
    \new_[49570]_ , \new_[49571]_ , \new_[49575]_ , \new_[49576]_ ,
    \new_[49577]_ , \new_[49581]_ , \new_[49582]_ , \new_[49585]_ ,
    \new_[49588]_ , \new_[49589]_ , \new_[49590]_ , \new_[49594]_ ,
    \new_[49595]_ , \new_[49599]_ , \new_[49600]_ , \new_[49601]_ ,
    \new_[49605]_ , \new_[49606]_ , \new_[49609]_ , \new_[49612]_ ,
    \new_[49613]_ , \new_[49614]_ , \new_[49618]_ , \new_[49619]_ ,
    \new_[49623]_ , \new_[49624]_ , \new_[49625]_ , \new_[49629]_ ,
    \new_[49630]_ , \new_[49633]_ , \new_[49636]_ , \new_[49637]_ ,
    \new_[49638]_ , \new_[49642]_ , \new_[49643]_ , \new_[49647]_ ,
    \new_[49648]_ , \new_[49649]_ , \new_[49653]_ , \new_[49654]_ ,
    \new_[49657]_ , \new_[49660]_ , \new_[49661]_ , \new_[49662]_ ,
    \new_[49666]_ , \new_[49667]_ , \new_[49671]_ , \new_[49672]_ ,
    \new_[49673]_ , \new_[49677]_ , \new_[49678]_ , \new_[49681]_ ,
    \new_[49684]_ , \new_[49685]_ , \new_[49686]_ , \new_[49690]_ ,
    \new_[49691]_ , \new_[49695]_ , \new_[49696]_ , \new_[49697]_ ,
    \new_[49701]_ , \new_[49702]_ , \new_[49705]_ , \new_[49708]_ ,
    \new_[49709]_ , \new_[49710]_ , \new_[49714]_ , \new_[49715]_ ,
    \new_[49719]_ , \new_[49720]_ , \new_[49721]_ , \new_[49725]_ ,
    \new_[49726]_ , \new_[49729]_ , \new_[49732]_ , \new_[49733]_ ,
    \new_[49734]_ , \new_[49738]_ , \new_[49739]_ , \new_[49743]_ ,
    \new_[49744]_ , \new_[49745]_ , \new_[49749]_ , \new_[49750]_ ,
    \new_[49753]_ , \new_[49756]_ , \new_[49757]_ , \new_[49758]_ ,
    \new_[49762]_ , \new_[49763]_ , \new_[49767]_ , \new_[49768]_ ,
    \new_[49769]_ , \new_[49773]_ , \new_[49774]_ , \new_[49777]_ ,
    \new_[49780]_ , \new_[49781]_ , \new_[49782]_ , \new_[49786]_ ,
    \new_[49787]_ , \new_[49791]_ , \new_[49792]_ , \new_[49793]_ ,
    \new_[49797]_ , \new_[49798]_ , \new_[49801]_ , \new_[49804]_ ,
    \new_[49805]_ , \new_[49806]_ , \new_[49810]_ , \new_[49811]_ ,
    \new_[49815]_ , \new_[49816]_ , \new_[49817]_ , \new_[49821]_ ,
    \new_[49822]_ , \new_[49825]_ , \new_[49828]_ , \new_[49829]_ ,
    \new_[49830]_ , \new_[49834]_ , \new_[49835]_ , \new_[49839]_ ,
    \new_[49840]_ , \new_[49841]_ , \new_[49845]_ , \new_[49846]_ ,
    \new_[49849]_ , \new_[49852]_ , \new_[49853]_ , \new_[49854]_ ,
    \new_[49858]_ , \new_[49859]_ , \new_[49863]_ , \new_[49864]_ ,
    \new_[49865]_ , \new_[49869]_ , \new_[49870]_ , \new_[49873]_ ,
    \new_[49876]_ , \new_[49877]_ , \new_[49878]_ , \new_[49882]_ ,
    \new_[49883]_ , \new_[49887]_ , \new_[49888]_ , \new_[49889]_ ,
    \new_[49893]_ , \new_[49894]_ , \new_[49897]_ , \new_[49900]_ ,
    \new_[49901]_ , \new_[49902]_ , \new_[49906]_ , \new_[49907]_ ,
    \new_[49911]_ , \new_[49912]_ , \new_[49913]_ , \new_[49917]_ ,
    \new_[49918]_ , \new_[49921]_ , \new_[49924]_ , \new_[49925]_ ,
    \new_[49926]_ , \new_[49930]_ , \new_[49931]_ , \new_[49935]_ ,
    \new_[49936]_ , \new_[49937]_ , \new_[49941]_ , \new_[49942]_ ,
    \new_[49945]_ , \new_[49948]_ , \new_[49949]_ , \new_[49950]_ ,
    \new_[49954]_ , \new_[49955]_ , \new_[49959]_ , \new_[49960]_ ,
    \new_[49961]_ , \new_[49965]_ , \new_[49966]_ , \new_[49969]_ ,
    \new_[49972]_ , \new_[49973]_ , \new_[49974]_ , \new_[49978]_ ,
    \new_[49979]_ , \new_[49983]_ , \new_[49984]_ , \new_[49985]_ ,
    \new_[49989]_ , \new_[49990]_ , \new_[49993]_ , \new_[49996]_ ,
    \new_[49997]_ , \new_[49998]_ , \new_[50002]_ , \new_[50003]_ ,
    \new_[50007]_ , \new_[50008]_ , \new_[50009]_ , \new_[50013]_ ,
    \new_[50014]_ , \new_[50017]_ , \new_[50020]_ , \new_[50021]_ ,
    \new_[50022]_ , \new_[50026]_ , \new_[50027]_ , \new_[50031]_ ,
    \new_[50032]_ , \new_[50033]_ , \new_[50037]_ , \new_[50038]_ ,
    \new_[50041]_ , \new_[50044]_ , \new_[50045]_ , \new_[50046]_ ,
    \new_[50050]_ , \new_[50051]_ , \new_[50055]_ , \new_[50056]_ ,
    \new_[50057]_ , \new_[50061]_ , \new_[50062]_ , \new_[50065]_ ,
    \new_[50068]_ , \new_[50069]_ , \new_[50070]_ , \new_[50074]_ ,
    \new_[50075]_ , \new_[50079]_ , \new_[50080]_ , \new_[50081]_ ,
    \new_[50085]_ , \new_[50086]_ , \new_[50089]_ , \new_[50092]_ ,
    \new_[50093]_ , \new_[50094]_ , \new_[50098]_ , \new_[50099]_ ,
    \new_[50103]_ , \new_[50104]_ , \new_[50105]_ , \new_[50109]_ ,
    \new_[50110]_ , \new_[50113]_ , \new_[50116]_ , \new_[50117]_ ,
    \new_[50118]_ , \new_[50122]_ , \new_[50123]_ , \new_[50127]_ ,
    \new_[50128]_ , \new_[50129]_ , \new_[50133]_ , \new_[50134]_ ,
    \new_[50137]_ , \new_[50140]_ , \new_[50141]_ , \new_[50142]_ ,
    \new_[50146]_ , \new_[50147]_ , \new_[50151]_ , \new_[50152]_ ,
    \new_[50153]_ , \new_[50157]_ , \new_[50158]_ , \new_[50161]_ ,
    \new_[50164]_ , \new_[50165]_ , \new_[50166]_ , \new_[50170]_ ,
    \new_[50171]_ , \new_[50175]_ , \new_[50176]_ , \new_[50177]_ ,
    \new_[50181]_ , \new_[50182]_ , \new_[50185]_ , \new_[50188]_ ,
    \new_[50189]_ , \new_[50190]_ , \new_[50194]_ , \new_[50195]_ ,
    \new_[50199]_ , \new_[50200]_ , \new_[50201]_ , \new_[50205]_ ,
    \new_[50206]_ , \new_[50209]_ , \new_[50212]_ , \new_[50213]_ ,
    \new_[50214]_ , \new_[50218]_ , \new_[50219]_ , \new_[50223]_ ,
    \new_[50224]_ , \new_[50225]_ , \new_[50229]_ , \new_[50230]_ ,
    \new_[50233]_ , \new_[50236]_ , \new_[50237]_ , \new_[50238]_ ,
    \new_[50242]_ , \new_[50243]_ , \new_[50247]_ , \new_[50248]_ ,
    \new_[50249]_ , \new_[50253]_ , \new_[50254]_ , \new_[50257]_ ,
    \new_[50260]_ , \new_[50261]_ , \new_[50262]_ , \new_[50266]_ ,
    \new_[50267]_ , \new_[50271]_ , \new_[50272]_ , \new_[50273]_ ,
    \new_[50277]_ , \new_[50278]_ , \new_[50281]_ , \new_[50284]_ ,
    \new_[50285]_ , \new_[50286]_ , \new_[50290]_ , \new_[50291]_ ,
    \new_[50295]_ , \new_[50296]_ , \new_[50297]_ , \new_[50301]_ ,
    \new_[50302]_ , \new_[50305]_ , \new_[50308]_ , \new_[50309]_ ,
    \new_[50310]_ , \new_[50314]_ , \new_[50315]_ , \new_[50319]_ ,
    \new_[50320]_ , \new_[50321]_ , \new_[50325]_ , \new_[50326]_ ,
    \new_[50329]_ , \new_[50332]_ , \new_[50333]_ , \new_[50334]_ ,
    \new_[50338]_ , \new_[50339]_ , \new_[50343]_ , \new_[50344]_ ,
    \new_[50345]_ , \new_[50349]_ , \new_[50350]_ , \new_[50353]_ ,
    \new_[50356]_ , \new_[50357]_ , \new_[50358]_ , \new_[50362]_ ,
    \new_[50363]_ , \new_[50367]_ , \new_[50368]_ , \new_[50369]_ ,
    \new_[50373]_ , \new_[50374]_ , \new_[50377]_ , \new_[50380]_ ,
    \new_[50381]_ , \new_[50382]_ , \new_[50386]_ , \new_[50387]_ ,
    \new_[50391]_ , \new_[50392]_ , \new_[50393]_ , \new_[50397]_ ,
    \new_[50398]_ , \new_[50401]_ , \new_[50404]_ , \new_[50405]_ ,
    \new_[50406]_ , \new_[50410]_ , \new_[50411]_ , \new_[50415]_ ,
    \new_[50416]_ , \new_[50417]_ , \new_[50421]_ , \new_[50422]_ ,
    \new_[50425]_ , \new_[50428]_ , \new_[50429]_ , \new_[50430]_ ,
    \new_[50434]_ , \new_[50435]_ , \new_[50439]_ , \new_[50440]_ ,
    \new_[50441]_ , \new_[50445]_ , \new_[50446]_ , \new_[50449]_ ,
    \new_[50452]_ , \new_[50453]_ , \new_[50454]_ , \new_[50458]_ ,
    \new_[50459]_ , \new_[50463]_ , \new_[50464]_ , \new_[50465]_ ,
    \new_[50469]_ , \new_[50470]_ , \new_[50473]_ , \new_[50476]_ ,
    \new_[50477]_ , \new_[50478]_ , \new_[50482]_ , \new_[50483]_ ,
    \new_[50487]_ , \new_[50488]_ , \new_[50489]_ , \new_[50493]_ ,
    \new_[50494]_ , \new_[50497]_ , \new_[50500]_ , \new_[50501]_ ,
    \new_[50502]_ , \new_[50506]_ , \new_[50507]_ , \new_[50511]_ ,
    \new_[50512]_ , \new_[50513]_ , \new_[50517]_ , \new_[50518]_ ,
    \new_[50521]_ , \new_[50524]_ , \new_[50525]_ , \new_[50526]_ ,
    \new_[50530]_ , \new_[50531]_ , \new_[50535]_ , \new_[50536]_ ,
    \new_[50537]_ , \new_[50541]_ , \new_[50542]_ , \new_[50545]_ ,
    \new_[50548]_ , \new_[50549]_ , \new_[50550]_ , \new_[50554]_ ,
    \new_[50555]_ , \new_[50559]_ , \new_[50560]_ , \new_[50561]_ ,
    \new_[50565]_ , \new_[50566]_ , \new_[50569]_ , \new_[50572]_ ,
    \new_[50573]_ , \new_[50574]_ , \new_[50578]_ , \new_[50579]_ ,
    \new_[50583]_ , \new_[50584]_ , \new_[50585]_ , \new_[50589]_ ,
    \new_[50590]_ , \new_[50593]_ , \new_[50596]_ , \new_[50597]_ ,
    \new_[50598]_ , \new_[50602]_ , \new_[50603]_ , \new_[50607]_ ,
    \new_[50608]_ , \new_[50609]_ , \new_[50613]_ , \new_[50614]_ ,
    \new_[50617]_ , \new_[50620]_ , \new_[50621]_ , \new_[50622]_ ,
    \new_[50626]_ , \new_[50627]_ , \new_[50631]_ , \new_[50632]_ ,
    \new_[50633]_ , \new_[50637]_ , \new_[50638]_ , \new_[50641]_ ,
    \new_[50644]_ , \new_[50645]_ , \new_[50646]_ , \new_[50650]_ ,
    \new_[50651]_ , \new_[50655]_ , \new_[50656]_ , \new_[50657]_ ,
    \new_[50661]_ , \new_[50662]_ , \new_[50665]_ , \new_[50668]_ ,
    \new_[50669]_ , \new_[50670]_ , \new_[50674]_ , \new_[50675]_ ,
    \new_[50679]_ , \new_[50680]_ , \new_[50681]_ , \new_[50685]_ ,
    \new_[50686]_ , \new_[50689]_ , \new_[50692]_ , \new_[50693]_ ,
    \new_[50694]_ , \new_[50698]_ , \new_[50699]_ , \new_[50703]_ ,
    \new_[50704]_ , \new_[50705]_ , \new_[50709]_ , \new_[50710]_ ,
    \new_[50713]_ , \new_[50716]_ , \new_[50717]_ , \new_[50718]_ ,
    \new_[50722]_ , \new_[50723]_ , \new_[50727]_ , \new_[50728]_ ,
    \new_[50729]_ , \new_[50733]_ , \new_[50734]_ , \new_[50737]_ ,
    \new_[50740]_ , \new_[50741]_ , \new_[50742]_ , \new_[50746]_ ,
    \new_[50747]_ , \new_[50751]_ , \new_[50752]_ , \new_[50753]_ ,
    \new_[50757]_ , \new_[50758]_ , \new_[50761]_ , \new_[50764]_ ,
    \new_[50765]_ , \new_[50766]_ , \new_[50770]_ , \new_[50771]_ ,
    \new_[50775]_ , \new_[50776]_ , \new_[50777]_ , \new_[50781]_ ,
    \new_[50782]_ , \new_[50785]_ , \new_[50788]_ , \new_[50789]_ ,
    \new_[50790]_ , \new_[50794]_ , \new_[50795]_ , \new_[50799]_ ,
    \new_[50800]_ , \new_[50801]_ , \new_[50805]_ , \new_[50806]_ ,
    \new_[50809]_ , \new_[50812]_ , \new_[50813]_ , \new_[50814]_ ,
    \new_[50818]_ , \new_[50819]_ , \new_[50823]_ , \new_[50824]_ ,
    \new_[50825]_ , \new_[50829]_ , \new_[50830]_ , \new_[50833]_ ,
    \new_[50836]_ , \new_[50837]_ , \new_[50838]_ , \new_[50842]_ ,
    \new_[50843]_ , \new_[50847]_ , \new_[50848]_ , \new_[50849]_ ,
    \new_[50853]_ , \new_[50854]_ , \new_[50857]_ , \new_[50860]_ ,
    \new_[50861]_ , \new_[50862]_ , \new_[50866]_ , \new_[50867]_ ,
    \new_[50871]_ , \new_[50872]_ , \new_[50873]_ , \new_[50877]_ ,
    \new_[50878]_ , \new_[50881]_ , \new_[50884]_ , \new_[50885]_ ,
    \new_[50886]_ , \new_[50890]_ , \new_[50891]_ , \new_[50895]_ ,
    \new_[50896]_ , \new_[50897]_ , \new_[50901]_ , \new_[50902]_ ,
    \new_[50905]_ , \new_[50908]_ , \new_[50909]_ , \new_[50910]_ ,
    \new_[50914]_ , \new_[50915]_ , \new_[50919]_ , \new_[50920]_ ,
    \new_[50921]_ , \new_[50925]_ , \new_[50926]_ , \new_[50929]_ ,
    \new_[50932]_ , \new_[50933]_ , \new_[50934]_ , \new_[50938]_ ,
    \new_[50939]_ , \new_[50943]_ , \new_[50944]_ , \new_[50945]_ ,
    \new_[50949]_ , \new_[50950]_ , \new_[50953]_ , \new_[50956]_ ,
    \new_[50957]_ , \new_[50958]_ , \new_[50962]_ , \new_[50963]_ ,
    \new_[50967]_ , \new_[50968]_ , \new_[50969]_ , \new_[50973]_ ,
    \new_[50974]_ , \new_[50977]_ , \new_[50980]_ , \new_[50981]_ ,
    \new_[50982]_ , \new_[50986]_ , \new_[50987]_ , \new_[50991]_ ,
    \new_[50992]_ , \new_[50993]_ , \new_[50997]_ , \new_[50998]_ ,
    \new_[51001]_ , \new_[51004]_ , \new_[51005]_ , \new_[51006]_ ,
    \new_[51010]_ , \new_[51011]_ , \new_[51015]_ , \new_[51016]_ ,
    \new_[51017]_ , \new_[51021]_ , \new_[51022]_ , \new_[51025]_ ,
    \new_[51028]_ , \new_[51029]_ , \new_[51030]_ , \new_[51034]_ ,
    \new_[51035]_ , \new_[51039]_ , \new_[51040]_ , \new_[51041]_ ,
    \new_[51045]_ , \new_[51046]_ , \new_[51049]_ , \new_[51052]_ ,
    \new_[51053]_ , \new_[51054]_ , \new_[51058]_ , \new_[51059]_ ,
    \new_[51063]_ , \new_[51064]_ , \new_[51065]_ , \new_[51069]_ ,
    \new_[51070]_ , \new_[51073]_ , \new_[51076]_ , \new_[51077]_ ,
    \new_[51078]_ , \new_[51082]_ , \new_[51083]_ , \new_[51087]_ ,
    \new_[51088]_ , \new_[51089]_ , \new_[51093]_ , \new_[51094]_ ,
    \new_[51097]_ , \new_[51100]_ , \new_[51101]_ , \new_[51102]_ ,
    \new_[51106]_ , \new_[51107]_ , \new_[51111]_ , \new_[51112]_ ,
    \new_[51113]_ , \new_[51117]_ , \new_[51118]_ , \new_[51121]_ ,
    \new_[51124]_ , \new_[51125]_ , \new_[51126]_ , \new_[51130]_ ,
    \new_[51131]_ , \new_[51135]_ , \new_[51136]_ , \new_[51137]_ ,
    \new_[51141]_ , \new_[51142]_ , \new_[51145]_ , \new_[51148]_ ,
    \new_[51149]_ , \new_[51150]_ , \new_[51154]_ , \new_[51155]_ ,
    \new_[51159]_ , \new_[51160]_ , \new_[51161]_ , \new_[51165]_ ,
    \new_[51166]_ , \new_[51169]_ , \new_[51172]_ , \new_[51173]_ ,
    \new_[51174]_ , \new_[51178]_ , \new_[51179]_ , \new_[51183]_ ,
    \new_[51184]_ , \new_[51185]_ , \new_[51189]_ , \new_[51190]_ ,
    \new_[51193]_ , \new_[51196]_ , \new_[51197]_ , \new_[51198]_ ,
    \new_[51202]_ , \new_[51203]_ , \new_[51207]_ , \new_[51208]_ ,
    \new_[51209]_ , \new_[51213]_ , \new_[51214]_ , \new_[51217]_ ,
    \new_[51220]_ , \new_[51221]_ , \new_[51222]_ , \new_[51226]_ ,
    \new_[51227]_ , \new_[51231]_ , \new_[51232]_ , \new_[51233]_ ,
    \new_[51237]_ , \new_[51238]_ , \new_[51241]_ , \new_[51244]_ ,
    \new_[51245]_ , \new_[51246]_ , \new_[51250]_ , \new_[51251]_ ,
    \new_[51255]_ , \new_[51256]_ , \new_[51257]_ , \new_[51261]_ ,
    \new_[51262]_ , \new_[51265]_ , \new_[51268]_ , \new_[51269]_ ,
    \new_[51270]_ , \new_[51274]_ , \new_[51275]_ , \new_[51279]_ ,
    \new_[51280]_ , \new_[51281]_ , \new_[51285]_ , \new_[51286]_ ,
    \new_[51289]_ , \new_[51292]_ , \new_[51293]_ , \new_[51294]_ ,
    \new_[51298]_ , \new_[51299]_ , \new_[51303]_ , \new_[51304]_ ,
    \new_[51305]_ , \new_[51309]_ , \new_[51310]_ , \new_[51313]_ ,
    \new_[51316]_ , \new_[51317]_ , \new_[51318]_ , \new_[51322]_ ,
    \new_[51323]_ , \new_[51327]_ , \new_[51328]_ , \new_[51329]_ ,
    \new_[51333]_ , \new_[51334]_ , \new_[51337]_ , \new_[51340]_ ,
    \new_[51341]_ , \new_[51342]_ , \new_[51346]_ , \new_[51347]_ ,
    \new_[51351]_ , \new_[51352]_ , \new_[51353]_ , \new_[51357]_ ,
    \new_[51358]_ , \new_[51361]_ , \new_[51364]_ , \new_[51365]_ ,
    \new_[51366]_ , \new_[51370]_ , \new_[51371]_ , \new_[51375]_ ,
    \new_[51376]_ , \new_[51377]_ , \new_[51381]_ , \new_[51382]_ ,
    \new_[51385]_ , \new_[51388]_ , \new_[51389]_ , \new_[51390]_ ,
    \new_[51394]_ , \new_[51395]_ , \new_[51399]_ , \new_[51400]_ ,
    \new_[51401]_ , \new_[51405]_ , \new_[51406]_ , \new_[51409]_ ,
    \new_[51412]_ , \new_[51413]_ , \new_[51414]_ , \new_[51418]_ ,
    \new_[51419]_ , \new_[51423]_ , \new_[51424]_ , \new_[51425]_ ,
    \new_[51429]_ , \new_[51430]_ , \new_[51433]_ , \new_[51436]_ ,
    \new_[51437]_ , \new_[51438]_ , \new_[51442]_ , \new_[51443]_ ,
    \new_[51447]_ , \new_[51448]_ , \new_[51449]_ , \new_[51453]_ ,
    \new_[51454]_ , \new_[51457]_ , \new_[51460]_ , \new_[51461]_ ,
    \new_[51462]_ , \new_[51466]_ , \new_[51467]_ , \new_[51471]_ ,
    \new_[51472]_ , \new_[51473]_ , \new_[51477]_ , \new_[51478]_ ,
    \new_[51481]_ , \new_[51484]_ , \new_[51485]_ , \new_[51486]_ ,
    \new_[51490]_ , \new_[51491]_ , \new_[51495]_ , \new_[51496]_ ,
    \new_[51497]_ , \new_[51501]_ , \new_[51502]_ , \new_[51505]_ ,
    \new_[51508]_ , \new_[51509]_ , \new_[51510]_ , \new_[51514]_ ,
    \new_[51515]_ , \new_[51519]_ , \new_[51520]_ , \new_[51521]_ ,
    \new_[51525]_ , \new_[51526]_ , \new_[51529]_ , \new_[51532]_ ,
    \new_[51533]_ , \new_[51534]_ , \new_[51538]_ , \new_[51539]_ ,
    \new_[51543]_ , \new_[51544]_ , \new_[51545]_ , \new_[51549]_ ,
    \new_[51550]_ , \new_[51553]_ , \new_[51556]_ , \new_[51557]_ ,
    \new_[51558]_ , \new_[51562]_ , \new_[51563]_ , \new_[51567]_ ,
    \new_[51568]_ , \new_[51569]_ , \new_[51573]_ , \new_[51574]_ ,
    \new_[51577]_ , \new_[51580]_ , \new_[51581]_ , \new_[51582]_ ,
    \new_[51586]_ , \new_[51587]_ , \new_[51591]_ , \new_[51592]_ ,
    \new_[51593]_ , \new_[51597]_ , \new_[51598]_ , \new_[51601]_ ,
    \new_[51604]_ , \new_[51605]_ , \new_[51606]_ , \new_[51610]_ ,
    \new_[51611]_ , \new_[51615]_ , \new_[51616]_ , \new_[51617]_ ,
    \new_[51621]_ , \new_[51622]_ , \new_[51625]_ , \new_[51628]_ ,
    \new_[51629]_ , \new_[51630]_ , \new_[51634]_ , \new_[51635]_ ,
    \new_[51639]_ , \new_[51640]_ , \new_[51641]_ , \new_[51645]_ ,
    \new_[51646]_ , \new_[51649]_ , \new_[51652]_ , \new_[51653]_ ,
    \new_[51654]_ , \new_[51658]_ , \new_[51659]_ , \new_[51663]_ ,
    \new_[51664]_ , \new_[51665]_ , \new_[51669]_ , \new_[51670]_ ,
    \new_[51673]_ , \new_[51676]_ , \new_[51677]_ , \new_[51678]_ ,
    \new_[51682]_ , \new_[51683]_ , \new_[51687]_ , \new_[51688]_ ,
    \new_[51689]_ , \new_[51693]_ , \new_[51694]_ , \new_[51697]_ ,
    \new_[51700]_ , \new_[51701]_ , \new_[51702]_ , \new_[51706]_ ,
    \new_[51707]_ , \new_[51711]_ , \new_[51712]_ , \new_[51713]_ ,
    \new_[51717]_ , \new_[51718]_ , \new_[51721]_ , \new_[51724]_ ,
    \new_[51725]_ , \new_[51726]_ , \new_[51730]_ , \new_[51731]_ ,
    \new_[51735]_ , \new_[51736]_ , \new_[51737]_ , \new_[51741]_ ,
    \new_[51742]_ , \new_[51745]_ , \new_[51748]_ , \new_[51749]_ ,
    \new_[51750]_ , \new_[51754]_ , \new_[51755]_ , \new_[51759]_ ,
    \new_[51760]_ , \new_[51761]_ , \new_[51765]_ , \new_[51766]_ ,
    \new_[51769]_ , \new_[51772]_ , \new_[51773]_ , \new_[51774]_ ,
    \new_[51778]_ , \new_[51779]_ , \new_[51783]_ , \new_[51784]_ ,
    \new_[51785]_ , \new_[51789]_ , \new_[51790]_ , \new_[51793]_ ,
    \new_[51796]_ , \new_[51797]_ , \new_[51798]_ , \new_[51802]_ ,
    \new_[51803]_ , \new_[51807]_ , \new_[51808]_ , \new_[51809]_ ,
    \new_[51813]_ , \new_[51814]_ , \new_[51817]_ , \new_[51820]_ ,
    \new_[51821]_ , \new_[51822]_ , \new_[51826]_ , \new_[51827]_ ,
    \new_[51831]_ , \new_[51832]_ , \new_[51833]_ , \new_[51837]_ ,
    \new_[51838]_ , \new_[51841]_ , \new_[51844]_ , \new_[51845]_ ,
    \new_[51846]_ , \new_[51850]_ , \new_[51851]_ , \new_[51855]_ ,
    \new_[51856]_ , \new_[51857]_ , \new_[51861]_ , \new_[51862]_ ,
    \new_[51865]_ , \new_[51868]_ , \new_[51869]_ , \new_[51870]_ ,
    \new_[51874]_ , \new_[51875]_ , \new_[51879]_ , \new_[51880]_ ,
    \new_[51881]_ , \new_[51885]_ , \new_[51886]_ , \new_[51889]_ ,
    \new_[51892]_ , \new_[51893]_ , \new_[51894]_ , \new_[51898]_ ,
    \new_[51899]_ , \new_[51903]_ , \new_[51904]_ , \new_[51905]_ ,
    \new_[51909]_ , \new_[51910]_ , \new_[51913]_ , \new_[51916]_ ,
    \new_[51917]_ , \new_[51918]_ , \new_[51922]_ , \new_[51923]_ ,
    \new_[51927]_ , \new_[51928]_ , \new_[51929]_ , \new_[51933]_ ,
    \new_[51934]_ , \new_[51937]_ , \new_[51940]_ , \new_[51941]_ ,
    \new_[51942]_ , \new_[51946]_ , \new_[51947]_ , \new_[51951]_ ,
    \new_[51952]_ , \new_[51953]_ , \new_[51957]_ , \new_[51958]_ ,
    \new_[51961]_ , \new_[51964]_ , \new_[51965]_ , \new_[51966]_ ,
    \new_[51970]_ , \new_[51971]_ , \new_[51975]_ , \new_[51976]_ ,
    \new_[51977]_ , \new_[51981]_ , \new_[51982]_ , \new_[51985]_ ,
    \new_[51988]_ , \new_[51989]_ , \new_[51990]_ , \new_[51994]_ ,
    \new_[51995]_ , \new_[51999]_ , \new_[52000]_ , \new_[52001]_ ,
    \new_[52005]_ , \new_[52006]_ , \new_[52009]_ , \new_[52012]_ ,
    \new_[52013]_ , \new_[52014]_ , \new_[52018]_ , \new_[52019]_ ,
    \new_[52023]_ , \new_[52024]_ , \new_[52025]_ , \new_[52029]_ ,
    \new_[52030]_ , \new_[52033]_ , \new_[52036]_ , \new_[52037]_ ,
    \new_[52038]_ , \new_[52042]_ , \new_[52043]_ , \new_[52047]_ ,
    \new_[52048]_ , \new_[52049]_ , \new_[52053]_ , \new_[52054]_ ,
    \new_[52057]_ , \new_[52060]_ , \new_[52061]_ , \new_[52062]_ ,
    \new_[52066]_ , \new_[52067]_ , \new_[52071]_ , \new_[52072]_ ,
    \new_[52073]_ , \new_[52077]_ , \new_[52078]_ , \new_[52081]_ ,
    \new_[52084]_ , \new_[52085]_ , \new_[52086]_ , \new_[52090]_ ,
    \new_[52091]_ , \new_[52095]_ , \new_[52096]_ , \new_[52097]_ ,
    \new_[52101]_ , \new_[52102]_ , \new_[52105]_ , \new_[52108]_ ,
    \new_[52109]_ , \new_[52110]_ , \new_[52114]_ , \new_[52115]_ ,
    \new_[52119]_ , \new_[52120]_ , \new_[52121]_ , \new_[52125]_ ,
    \new_[52126]_ , \new_[52129]_ , \new_[52132]_ , \new_[52133]_ ,
    \new_[52134]_ , \new_[52138]_ , \new_[52139]_ , \new_[52143]_ ,
    \new_[52144]_ , \new_[52145]_ , \new_[52149]_ , \new_[52150]_ ,
    \new_[52153]_ , \new_[52156]_ , \new_[52157]_ , \new_[52158]_ ,
    \new_[52162]_ , \new_[52163]_ , \new_[52167]_ , \new_[52168]_ ,
    \new_[52169]_ , \new_[52173]_ , \new_[52174]_ , \new_[52177]_ ,
    \new_[52180]_ , \new_[52181]_ , \new_[52182]_ , \new_[52186]_ ,
    \new_[52187]_ , \new_[52191]_ , \new_[52192]_ , \new_[52193]_ ,
    \new_[52197]_ , \new_[52198]_ , \new_[52201]_ , \new_[52204]_ ,
    \new_[52205]_ , \new_[52206]_ , \new_[52210]_ , \new_[52211]_ ,
    \new_[52215]_ , \new_[52216]_ , \new_[52217]_ , \new_[52221]_ ,
    \new_[52222]_ , \new_[52225]_ , \new_[52228]_ , \new_[52229]_ ,
    \new_[52230]_ , \new_[52234]_ , \new_[52235]_ , \new_[52239]_ ,
    \new_[52240]_ , \new_[52241]_ , \new_[52245]_ , \new_[52246]_ ,
    \new_[52249]_ , \new_[52252]_ , \new_[52253]_ , \new_[52254]_ ,
    \new_[52258]_ , \new_[52259]_ , \new_[52263]_ , \new_[52264]_ ,
    \new_[52265]_ , \new_[52269]_ , \new_[52270]_ , \new_[52273]_ ,
    \new_[52276]_ , \new_[52277]_ , \new_[52278]_ , \new_[52282]_ ,
    \new_[52283]_ , \new_[52287]_ , \new_[52288]_ , \new_[52289]_ ,
    \new_[52293]_ , \new_[52294]_ , \new_[52297]_ , \new_[52300]_ ,
    \new_[52301]_ , \new_[52302]_ , \new_[52306]_ , \new_[52307]_ ,
    \new_[52311]_ , \new_[52312]_ , \new_[52313]_ , \new_[52317]_ ,
    \new_[52318]_ , \new_[52321]_ , \new_[52324]_ , \new_[52325]_ ,
    \new_[52326]_ , \new_[52330]_ , \new_[52331]_ , \new_[52335]_ ,
    \new_[52336]_ , \new_[52337]_ , \new_[52341]_ , \new_[52342]_ ,
    \new_[52345]_ , \new_[52348]_ , \new_[52349]_ , \new_[52350]_ ,
    \new_[52354]_ , \new_[52355]_ , \new_[52359]_ , \new_[52360]_ ,
    \new_[52361]_ , \new_[52365]_ , \new_[52366]_ , \new_[52369]_ ,
    \new_[52372]_ , \new_[52373]_ , \new_[52374]_ , \new_[52378]_ ,
    \new_[52379]_ , \new_[52383]_ , \new_[52384]_ , \new_[52385]_ ,
    \new_[52389]_ , \new_[52390]_ , \new_[52393]_ , \new_[52396]_ ,
    \new_[52397]_ , \new_[52398]_ , \new_[52402]_ , \new_[52403]_ ,
    \new_[52407]_ , \new_[52408]_ , \new_[52409]_ , \new_[52413]_ ,
    \new_[52414]_ , \new_[52417]_ , \new_[52420]_ , \new_[52421]_ ,
    \new_[52422]_ , \new_[52426]_ , \new_[52427]_ , \new_[52431]_ ,
    \new_[52432]_ , \new_[52433]_ , \new_[52437]_ , \new_[52438]_ ,
    \new_[52441]_ , \new_[52444]_ , \new_[52445]_ , \new_[52446]_ ,
    \new_[52450]_ , \new_[52451]_ , \new_[52455]_ , \new_[52456]_ ,
    \new_[52457]_ , \new_[52461]_ , \new_[52462]_ , \new_[52465]_ ,
    \new_[52468]_ , \new_[52469]_ , \new_[52470]_ , \new_[52474]_ ,
    \new_[52475]_ , \new_[52479]_ , \new_[52480]_ , \new_[52481]_ ,
    \new_[52485]_ , \new_[52486]_ , \new_[52489]_ , \new_[52492]_ ,
    \new_[52493]_ , \new_[52494]_ , \new_[52498]_ , \new_[52499]_ ,
    \new_[52503]_ , \new_[52504]_ , \new_[52505]_ , \new_[52509]_ ,
    \new_[52510]_ , \new_[52513]_ , \new_[52516]_ , \new_[52517]_ ,
    \new_[52518]_ , \new_[52522]_ , \new_[52523]_ , \new_[52527]_ ,
    \new_[52528]_ , \new_[52529]_ , \new_[52533]_ , \new_[52534]_ ,
    \new_[52537]_ , \new_[52540]_ , \new_[52541]_ , \new_[52542]_ ,
    \new_[52546]_ , \new_[52547]_ , \new_[52551]_ , \new_[52552]_ ,
    \new_[52553]_ , \new_[52557]_ , \new_[52558]_ , \new_[52561]_ ,
    \new_[52564]_ , \new_[52565]_ , \new_[52566]_ , \new_[52570]_ ,
    \new_[52571]_ , \new_[52575]_ , \new_[52576]_ , \new_[52577]_ ,
    \new_[52581]_ , \new_[52582]_ , \new_[52585]_ , \new_[52588]_ ,
    \new_[52589]_ , \new_[52590]_ , \new_[52594]_ , \new_[52595]_ ,
    \new_[52599]_ , \new_[52600]_ , \new_[52601]_ , \new_[52605]_ ,
    \new_[52606]_ , \new_[52609]_ , \new_[52612]_ , \new_[52613]_ ,
    \new_[52614]_ , \new_[52618]_ , \new_[52619]_ , \new_[52623]_ ,
    \new_[52624]_ , \new_[52625]_ , \new_[52629]_ , \new_[52630]_ ,
    \new_[52633]_ , \new_[52636]_ , \new_[52637]_ , \new_[52638]_ ,
    \new_[52642]_ , \new_[52643]_ , \new_[52647]_ , \new_[52648]_ ,
    \new_[52649]_ , \new_[52653]_ , \new_[52654]_ , \new_[52657]_ ,
    \new_[52660]_ , \new_[52661]_ , \new_[52662]_ , \new_[52666]_ ,
    \new_[52667]_ , \new_[52671]_ , \new_[52672]_ , \new_[52673]_ ,
    \new_[52677]_ , \new_[52678]_ , \new_[52681]_ , \new_[52684]_ ,
    \new_[52685]_ , \new_[52686]_ , \new_[52690]_ , \new_[52691]_ ,
    \new_[52695]_ , \new_[52696]_ , \new_[52697]_ , \new_[52701]_ ,
    \new_[52702]_ , \new_[52705]_ , \new_[52708]_ , \new_[52709]_ ,
    \new_[52710]_ , \new_[52714]_ , \new_[52715]_ , \new_[52719]_ ,
    \new_[52720]_ , \new_[52721]_ , \new_[52725]_ , \new_[52726]_ ,
    \new_[52729]_ , \new_[52732]_ , \new_[52733]_ , \new_[52734]_ ,
    \new_[52738]_ , \new_[52739]_ , \new_[52743]_ , \new_[52744]_ ,
    \new_[52745]_ , \new_[52749]_ , \new_[52750]_ , \new_[52753]_ ,
    \new_[52756]_ , \new_[52757]_ , \new_[52758]_ , \new_[52762]_ ,
    \new_[52763]_ , \new_[52767]_ , \new_[52768]_ , \new_[52769]_ ,
    \new_[52773]_ , \new_[52774]_ , \new_[52777]_ , \new_[52780]_ ,
    \new_[52781]_ , \new_[52782]_ , \new_[52786]_ , \new_[52787]_ ,
    \new_[52791]_ , \new_[52792]_ , \new_[52793]_ , \new_[52797]_ ,
    \new_[52798]_ , \new_[52801]_ , \new_[52804]_ , \new_[52805]_ ,
    \new_[52806]_ , \new_[52810]_ , \new_[52811]_ , \new_[52815]_ ,
    \new_[52816]_ , \new_[52817]_ , \new_[52821]_ , \new_[52822]_ ,
    \new_[52825]_ , \new_[52828]_ , \new_[52829]_ , \new_[52830]_ ,
    \new_[52834]_ , \new_[52835]_ , \new_[52839]_ , \new_[52840]_ ,
    \new_[52841]_ , \new_[52845]_ , \new_[52846]_ , \new_[52849]_ ,
    \new_[52852]_ , \new_[52853]_ , \new_[52854]_ , \new_[52858]_ ,
    \new_[52859]_ , \new_[52863]_ , \new_[52864]_ , \new_[52865]_ ,
    \new_[52869]_ , \new_[52870]_ , \new_[52873]_ , \new_[52876]_ ,
    \new_[52877]_ , \new_[52878]_ , \new_[52882]_ , \new_[52883]_ ,
    \new_[52887]_ , \new_[52888]_ , \new_[52889]_ , \new_[52893]_ ,
    \new_[52894]_ , \new_[52897]_ , \new_[52900]_ , \new_[52901]_ ,
    \new_[52902]_ , \new_[52906]_ , \new_[52907]_ , \new_[52911]_ ,
    \new_[52912]_ , \new_[52913]_ , \new_[52917]_ , \new_[52918]_ ,
    \new_[52921]_ , \new_[52924]_ , \new_[52925]_ , \new_[52926]_ ,
    \new_[52930]_ , \new_[52931]_ , \new_[52935]_ , \new_[52936]_ ,
    \new_[52937]_ , \new_[52941]_ , \new_[52942]_ , \new_[52945]_ ,
    \new_[52948]_ , \new_[52949]_ , \new_[52950]_ , \new_[52954]_ ,
    \new_[52955]_ , \new_[52959]_ , \new_[52960]_ , \new_[52961]_ ,
    \new_[52965]_ , \new_[52966]_ , \new_[52969]_ , \new_[52972]_ ,
    \new_[52973]_ , \new_[52974]_ , \new_[52978]_ , \new_[52979]_ ,
    \new_[52983]_ , \new_[52984]_ , \new_[52985]_ , \new_[52989]_ ,
    \new_[52990]_ , \new_[52993]_ , \new_[52996]_ , \new_[52997]_ ,
    \new_[52998]_ , \new_[53002]_ , \new_[53003]_ , \new_[53007]_ ,
    \new_[53008]_ , \new_[53009]_ , \new_[53013]_ , \new_[53014]_ ,
    \new_[53017]_ , \new_[53020]_ , \new_[53021]_ , \new_[53022]_ ,
    \new_[53026]_ , \new_[53027]_ , \new_[53031]_ , \new_[53032]_ ,
    \new_[53033]_ , \new_[53037]_ , \new_[53038]_ , \new_[53041]_ ,
    \new_[53044]_ , \new_[53045]_ , \new_[53046]_ , \new_[53050]_ ,
    \new_[53051]_ , \new_[53055]_ , \new_[53056]_ , \new_[53057]_ ,
    \new_[53061]_ , \new_[53062]_ , \new_[53065]_ , \new_[53068]_ ,
    \new_[53069]_ , \new_[53070]_ , \new_[53074]_ , \new_[53075]_ ,
    \new_[53079]_ , \new_[53080]_ , \new_[53081]_ , \new_[53085]_ ,
    \new_[53086]_ , \new_[53089]_ , \new_[53092]_ , \new_[53093]_ ,
    \new_[53094]_ , \new_[53098]_ , \new_[53099]_ , \new_[53103]_ ,
    \new_[53104]_ , \new_[53105]_ , \new_[53109]_ , \new_[53110]_ ,
    \new_[53113]_ , \new_[53116]_ , \new_[53117]_ , \new_[53118]_ ,
    \new_[53122]_ , \new_[53123]_ , \new_[53127]_ , \new_[53128]_ ,
    \new_[53129]_ , \new_[53133]_ , \new_[53134]_ , \new_[53137]_ ,
    \new_[53140]_ , \new_[53141]_ , \new_[53142]_ , \new_[53146]_ ,
    \new_[53147]_ , \new_[53151]_ , \new_[53152]_ , \new_[53153]_ ,
    \new_[53157]_ , \new_[53158]_ , \new_[53161]_ , \new_[53164]_ ,
    \new_[53165]_ , \new_[53166]_ , \new_[53170]_ , \new_[53171]_ ,
    \new_[53175]_ , \new_[53176]_ , \new_[53177]_ , \new_[53181]_ ,
    \new_[53182]_ , \new_[53185]_ , \new_[53188]_ , \new_[53189]_ ,
    \new_[53190]_ , \new_[53194]_ , \new_[53195]_ , \new_[53199]_ ,
    \new_[53200]_ , \new_[53201]_ , \new_[53205]_ , \new_[53206]_ ,
    \new_[53209]_ , \new_[53212]_ , \new_[53213]_ , \new_[53214]_ ,
    \new_[53218]_ , \new_[53219]_ , \new_[53223]_ , \new_[53224]_ ,
    \new_[53225]_ , \new_[53229]_ , \new_[53230]_ , \new_[53233]_ ,
    \new_[53236]_ , \new_[53237]_ , \new_[53238]_ , \new_[53242]_ ,
    \new_[53243]_ , \new_[53247]_ , \new_[53248]_ , \new_[53249]_ ,
    \new_[53253]_ , \new_[53254]_ , \new_[53257]_ , \new_[53260]_ ,
    \new_[53261]_ , \new_[53262]_ , \new_[53266]_ , \new_[53267]_ ,
    \new_[53271]_ , \new_[53272]_ , \new_[53273]_ , \new_[53277]_ ,
    \new_[53278]_ , \new_[53281]_ , \new_[53284]_ , \new_[53285]_ ,
    \new_[53286]_ , \new_[53290]_ , \new_[53291]_ , \new_[53295]_ ,
    \new_[53296]_ , \new_[53297]_ , \new_[53301]_ , \new_[53302]_ ,
    \new_[53305]_ , \new_[53308]_ , \new_[53309]_ , \new_[53310]_ ,
    \new_[53314]_ , \new_[53315]_ , \new_[53319]_ , \new_[53320]_ ,
    \new_[53321]_ , \new_[53325]_ , \new_[53326]_ , \new_[53329]_ ,
    \new_[53332]_ , \new_[53333]_ , \new_[53334]_ , \new_[53338]_ ,
    \new_[53339]_ , \new_[53343]_ , \new_[53344]_ , \new_[53345]_ ,
    \new_[53349]_ , \new_[53350]_ , \new_[53353]_ , \new_[53356]_ ,
    \new_[53357]_ , \new_[53358]_ , \new_[53362]_ , \new_[53363]_ ,
    \new_[53367]_ , \new_[53368]_ , \new_[53369]_ , \new_[53373]_ ,
    \new_[53374]_ , \new_[53377]_ , \new_[53380]_ , \new_[53381]_ ,
    \new_[53382]_ , \new_[53386]_ , \new_[53387]_ , \new_[53391]_ ,
    \new_[53392]_ , \new_[53393]_ , \new_[53397]_ , \new_[53398]_ ,
    \new_[53401]_ , \new_[53404]_ , \new_[53405]_ , \new_[53406]_ ,
    \new_[53410]_ , \new_[53411]_ , \new_[53415]_ , \new_[53416]_ ,
    \new_[53417]_ , \new_[53421]_ , \new_[53422]_ , \new_[53425]_ ,
    \new_[53428]_ , \new_[53429]_ , \new_[53430]_ , \new_[53434]_ ,
    \new_[53435]_ , \new_[53439]_ , \new_[53440]_ , \new_[53441]_ ,
    \new_[53445]_ , \new_[53446]_ , \new_[53449]_ , \new_[53452]_ ,
    \new_[53453]_ , \new_[53454]_ , \new_[53458]_ , \new_[53459]_ ,
    \new_[53463]_ , \new_[53464]_ , \new_[53465]_ , \new_[53469]_ ,
    \new_[53470]_ , \new_[53473]_ , \new_[53476]_ , \new_[53477]_ ,
    \new_[53478]_ , \new_[53482]_ , \new_[53483]_ , \new_[53487]_ ,
    \new_[53488]_ , \new_[53489]_ , \new_[53493]_ , \new_[53494]_ ,
    \new_[53497]_ , \new_[53500]_ , \new_[53501]_ , \new_[53502]_ ,
    \new_[53506]_ , \new_[53507]_ , \new_[53511]_ , \new_[53512]_ ,
    \new_[53513]_ , \new_[53517]_ , \new_[53518]_ , \new_[53521]_ ,
    \new_[53524]_ , \new_[53525]_ , \new_[53526]_ , \new_[53530]_ ,
    \new_[53531]_ , \new_[53535]_ , \new_[53536]_ , \new_[53537]_ ,
    \new_[53541]_ , \new_[53542]_ , \new_[53545]_ , \new_[53548]_ ,
    \new_[53549]_ , \new_[53550]_ , \new_[53554]_ , \new_[53555]_ ,
    \new_[53559]_ , \new_[53560]_ , \new_[53561]_ , \new_[53565]_ ,
    \new_[53566]_ , \new_[53569]_ , \new_[53572]_ , \new_[53573]_ ,
    \new_[53574]_ , \new_[53578]_ , \new_[53579]_ , \new_[53583]_ ,
    \new_[53584]_ , \new_[53585]_ , \new_[53589]_ , \new_[53590]_ ,
    \new_[53593]_ , \new_[53596]_ , \new_[53597]_ , \new_[53598]_ ,
    \new_[53602]_ , \new_[53603]_ , \new_[53607]_ , \new_[53608]_ ,
    \new_[53609]_ , \new_[53613]_ , \new_[53614]_ , \new_[53617]_ ,
    \new_[53620]_ , \new_[53621]_ , \new_[53622]_ , \new_[53626]_ ,
    \new_[53627]_ , \new_[53631]_ , \new_[53632]_ , \new_[53633]_ ,
    \new_[53637]_ , \new_[53638]_ , \new_[53641]_ , \new_[53644]_ ,
    \new_[53645]_ , \new_[53646]_ , \new_[53650]_ , \new_[53651]_ ,
    \new_[53655]_ , \new_[53656]_ , \new_[53657]_ , \new_[53661]_ ,
    \new_[53662]_ , \new_[53665]_ , \new_[53668]_ , \new_[53669]_ ,
    \new_[53670]_ , \new_[53674]_ , \new_[53675]_ , \new_[53679]_ ,
    \new_[53680]_ , \new_[53681]_ , \new_[53685]_ , \new_[53686]_ ,
    \new_[53689]_ , \new_[53692]_ , \new_[53693]_ , \new_[53694]_ ,
    \new_[53698]_ , \new_[53699]_ , \new_[53703]_ , \new_[53704]_ ,
    \new_[53705]_ , \new_[53709]_ , \new_[53710]_ , \new_[53713]_ ,
    \new_[53716]_ , \new_[53717]_ , \new_[53718]_ , \new_[53722]_ ,
    \new_[53723]_ , \new_[53727]_ , \new_[53728]_ , \new_[53729]_ ,
    \new_[53733]_ , \new_[53734]_ , \new_[53737]_ , \new_[53740]_ ,
    \new_[53741]_ , \new_[53742]_ , \new_[53746]_ , \new_[53747]_ ,
    \new_[53751]_ , \new_[53752]_ , \new_[53753]_ , \new_[53757]_ ,
    \new_[53758]_ , \new_[53761]_ , \new_[53764]_ , \new_[53765]_ ,
    \new_[53766]_ , \new_[53770]_ , \new_[53771]_ , \new_[53775]_ ,
    \new_[53776]_ , \new_[53777]_ , \new_[53781]_ , \new_[53782]_ ,
    \new_[53785]_ , \new_[53788]_ , \new_[53789]_ , \new_[53790]_ ,
    \new_[53794]_ , \new_[53795]_ , \new_[53799]_ , \new_[53800]_ ,
    \new_[53801]_ , \new_[53805]_ , \new_[53806]_ , \new_[53809]_ ,
    \new_[53812]_ , \new_[53813]_ , \new_[53814]_ , \new_[53818]_ ,
    \new_[53819]_ , \new_[53823]_ , \new_[53824]_ , \new_[53825]_ ,
    \new_[53829]_ , \new_[53830]_ , \new_[53833]_ , \new_[53836]_ ,
    \new_[53837]_ , \new_[53838]_ , \new_[53842]_ , \new_[53843]_ ,
    \new_[53847]_ , \new_[53848]_ , \new_[53849]_ , \new_[53853]_ ,
    \new_[53854]_ , \new_[53857]_ , \new_[53860]_ , \new_[53861]_ ,
    \new_[53862]_ , \new_[53866]_ , \new_[53867]_ , \new_[53871]_ ,
    \new_[53872]_ , \new_[53873]_ , \new_[53877]_ , \new_[53878]_ ,
    \new_[53881]_ , \new_[53884]_ , \new_[53885]_ , \new_[53886]_ ,
    \new_[53890]_ , \new_[53891]_ , \new_[53895]_ , \new_[53896]_ ,
    \new_[53897]_ , \new_[53901]_ , \new_[53902]_ , \new_[53905]_ ,
    \new_[53908]_ , \new_[53909]_ , \new_[53910]_ , \new_[53914]_ ,
    \new_[53915]_ , \new_[53919]_ , \new_[53920]_ , \new_[53921]_ ,
    \new_[53925]_ , \new_[53926]_ , \new_[53929]_ , \new_[53932]_ ,
    \new_[53933]_ , \new_[53934]_ , \new_[53938]_ , \new_[53939]_ ,
    \new_[53943]_ , \new_[53944]_ , \new_[53945]_ , \new_[53949]_ ,
    \new_[53950]_ , \new_[53953]_ , \new_[53956]_ , \new_[53957]_ ,
    \new_[53958]_ , \new_[53962]_ , \new_[53963]_ , \new_[53967]_ ,
    \new_[53968]_ , \new_[53969]_ , \new_[53973]_ , \new_[53974]_ ,
    \new_[53977]_ , \new_[53980]_ , \new_[53981]_ , \new_[53982]_ ,
    \new_[53986]_ , \new_[53987]_ , \new_[53991]_ , \new_[53992]_ ,
    \new_[53993]_ , \new_[53997]_ , \new_[53998]_ , \new_[54001]_ ,
    \new_[54004]_ , \new_[54005]_ , \new_[54006]_ , \new_[54010]_ ,
    \new_[54011]_ , \new_[54015]_ , \new_[54016]_ , \new_[54017]_ ,
    \new_[54021]_ , \new_[54022]_ , \new_[54025]_ , \new_[54028]_ ,
    \new_[54029]_ , \new_[54030]_ , \new_[54034]_ , \new_[54035]_ ,
    \new_[54039]_ , \new_[54040]_ , \new_[54041]_ , \new_[54045]_ ,
    \new_[54046]_ , \new_[54049]_ , \new_[54052]_ , \new_[54053]_ ,
    \new_[54054]_ , \new_[54058]_ , \new_[54059]_ , \new_[54063]_ ,
    \new_[54064]_ , \new_[54065]_ , \new_[54069]_ , \new_[54070]_ ,
    \new_[54073]_ , \new_[54076]_ , \new_[54077]_ , \new_[54078]_ ,
    \new_[54082]_ , \new_[54083]_ , \new_[54087]_ , \new_[54088]_ ,
    \new_[54089]_ , \new_[54093]_ , \new_[54094]_ , \new_[54097]_ ,
    \new_[54100]_ , \new_[54101]_ , \new_[54102]_ , \new_[54106]_ ,
    \new_[54107]_ , \new_[54111]_ , \new_[54112]_ , \new_[54113]_ ,
    \new_[54117]_ , \new_[54118]_ , \new_[54121]_ , \new_[54124]_ ,
    \new_[54125]_ , \new_[54126]_ , \new_[54130]_ , \new_[54131]_ ,
    \new_[54135]_ , \new_[54136]_ , \new_[54137]_ , \new_[54141]_ ,
    \new_[54142]_ , \new_[54145]_ , \new_[54148]_ , \new_[54149]_ ,
    \new_[54150]_ , \new_[54154]_ , \new_[54155]_ , \new_[54159]_ ,
    \new_[54160]_ , \new_[54161]_ , \new_[54165]_ , \new_[54166]_ ,
    \new_[54169]_ , \new_[54172]_ , \new_[54173]_ , \new_[54174]_ ,
    \new_[54178]_ , \new_[54179]_ , \new_[54183]_ , \new_[54184]_ ,
    \new_[54185]_ , \new_[54189]_ , \new_[54190]_ , \new_[54193]_ ,
    \new_[54196]_ , \new_[54197]_ , \new_[54198]_ , \new_[54202]_ ,
    \new_[54203]_ , \new_[54207]_ , \new_[54208]_ , \new_[54209]_ ,
    \new_[54213]_ , \new_[54214]_ , \new_[54217]_ , \new_[54220]_ ,
    \new_[54221]_ , \new_[54222]_ , \new_[54226]_ , \new_[54227]_ ,
    \new_[54231]_ , \new_[54232]_ , \new_[54233]_ , \new_[54237]_ ,
    \new_[54238]_ , \new_[54241]_ , \new_[54244]_ , \new_[54245]_ ,
    \new_[54246]_ , \new_[54250]_ , \new_[54251]_ , \new_[54255]_ ,
    \new_[54256]_ , \new_[54257]_ , \new_[54261]_ , \new_[54262]_ ,
    \new_[54265]_ , \new_[54268]_ , \new_[54269]_ , \new_[54270]_ ,
    \new_[54274]_ , \new_[54275]_ , \new_[54279]_ , \new_[54280]_ ,
    \new_[54281]_ , \new_[54285]_ , \new_[54286]_ , \new_[54289]_ ,
    \new_[54292]_ , \new_[54293]_ , \new_[54294]_ , \new_[54298]_ ,
    \new_[54299]_ , \new_[54303]_ , \new_[54304]_ , \new_[54305]_ ,
    \new_[54309]_ , \new_[54310]_ , \new_[54313]_ , \new_[54316]_ ,
    \new_[54317]_ , \new_[54318]_ , \new_[54322]_ , \new_[54323]_ ,
    \new_[54327]_ , \new_[54328]_ , \new_[54329]_ , \new_[54333]_ ,
    \new_[54334]_ , \new_[54337]_ , \new_[54340]_ , \new_[54341]_ ,
    \new_[54342]_ , \new_[54346]_ , \new_[54347]_ , \new_[54351]_ ,
    \new_[54352]_ , \new_[54353]_ , \new_[54357]_ , \new_[54358]_ ,
    \new_[54361]_ , \new_[54364]_ , \new_[54365]_ , \new_[54366]_ ,
    \new_[54370]_ , \new_[54371]_ , \new_[54375]_ , \new_[54376]_ ,
    \new_[54377]_ , \new_[54381]_ , \new_[54382]_ , \new_[54385]_ ,
    \new_[54388]_ , \new_[54389]_ , \new_[54390]_ , \new_[54394]_ ,
    \new_[54395]_ , \new_[54399]_ , \new_[54400]_ , \new_[54401]_ ,
    \new_[54405]_ , \new_[54406]_ , \new_[54409]_ , \new_[54412]_ ,
    \new_[54413]_ , \new_[54414]_ , \new_[54418]_ , \new_[54419]_ ,
    \new_[54423]_ , \new_[54424]_ , \new_[54425]_ , \new_[54429]_ ,
    \new_[54430]_ , \new_[54433]_ , \new_[54436]_ , \new_[54437]_ ,
    \new_[54438]_ , \new_[54442]_ , \new_[54443]_ , \new_[54447]_ ,
    \new_[54448]_ , \new_[54449]_ , \new_[54453]_ , \new_[54454]_ ,
    \new_[54457]_ , \new_[54460]_ , \new_[54461]_ , \new_[54462]_ ,
    \new_[54466]_ , \new_[54467]_ , \new_[54471]_ , \new_[54472]_ ,
    \new_[54473]_ , \new_[54477]_ , \new_[54478]_ , \new_[54481]_ ,
    \new_[54484]_ , \new_[54485]_ , \new_[54486]_ , \new_[54490]_ ,
    \new_[54491]_ , \new_[54495]_ , \new_[54496]_ , \new_[54497]_ ,
    \new_[54501]_ , \new_[54502]_ , \new_[54505]_ , \new_[54508]_ ,
    \new_[54509]_ , \new_[54510]_ , \new_[54514]_ , \new_[54515]_ ,
    \new_[54519]_ , \new_[54520]_ , \new_[54521]_ , \new_[54525]_ ,
    \new_[54526]_ , \new_[54529]_ , \new_[54532]_ , \new_[54533]_ ,
    \new_[54534]_ , \new_[54538]_ , \new_[54539]_ , \new_[54543]_ ,
    \new_[54544]_ , \new_[54545]_ , \new_[54549]_ , \new_[54550]_ ,
    \new_[54553]_ , \new_[54556]_ , \new_[54557]_ , \new_[54558]_ ,
    \new_[54562]_ , \new_[54563]_ , \new_[54567]_ , \new_[54568]_ ,
    \new_[54569]_ , \new_[54573]_ , \new_[54574]_ , \new_[54577]_ ,
    \new_[54580]_ , \new_[54581]_ , \new_[54582]_ , \new_[54586]_ ,
    \new_[54587]_ , \new_[54591]_ , \new_[54592]_ , \new_[54593]_ ,
    \new_[54597]_ , \new_[54598]_ , \new_[54601]_ , \new_[54604]_ ,
    \new_[54605]_ , \new_[54606]_ , \new_[54610]_ , \new_[54611]_ ,
    \new_[54615]_ , \new_[54616]_ , \new_[54617]_ , \new_[54621]_ ,
    \new_[54622]_ , \new_[54625]_ , \new_[54628]_ , \new_[54629]_ ,
    \new_[54630]_ , \new_[54634]_ , \new_[54635]_ , \new_[54639]_ ,
    \new_[54640]_ , \new_[54641]_ , \new_[54645]_ , \new_[54646]_ ,
    \new_[54649]_ , \new_[54652]_ , \new_[54653]_ , \new_[54654]_ ,
    \new_[54658]_ , \new_[54659]_ , \new_[54663]_ , \new_[54664]_ ,
    \new_[54665]_ , \new_[54669]_ , \new_[54670]_ , \new_[54673]_ ,
    \new_[54676]_ , \new_[54677]_ , \new_[54678]_ , \new_[54682]_ ,
    \new_[54683]_ , \new_[54687]_ , \new_[54688]_ , \new_[54689]_ ,
    \new_[54693]_ , \new_[54694]_ , \new_[54697]_ , \new_[54700]_ ,
    \new_[54701]_ , \new_[54702]_ , \new_[54706]_ , \new_[54707]_ ,
    \new_[54711]_ , \new_[54712]_ , \new_[54713]_ , \new_[54717]_ ,
    \new_[54718]_ , \new_[54721]_ , \new_[54724]_ , \new_[54725]_ ,
    \new_[54726]_ , \new_[54730]_ , \new_[54731]_ , \new_[54735]_ ,
    \new_[54736]_ , \new_[54737]_ , \new_[54741]_ , \new_[54742]_ ,
    \new_[54745]_ , \new_[54748]_ , \new_[54749]_ , \new_[54750]_ ,
    \new_[54754]_ , \new_[54755]_ , \new_[54759]_ , \new_[54760]_ ,
    \new_[54761]_ , \new_[54765]_ , \new_[54766]_ , \new_[54769]_ ,
    \new_[54772]_ , \new_[54773]_ , \new_[54774]_ , \new_[54778]_ ,
    \new_[54779]_ , \new_[54783]_ , \new_[54784]_ , \new_[54785]_ ,
    \new_[54789]_ , \new_[54790]_ , \new_[54793]_ , \new_[54796]_ ,
    \new_[54797]_ , \new_[54798]_ , \new_[54802]_ , \new_[54803]_ ,
    \new_[54807]_ , \new_[54808]_ , \new_[54809]_ , \new_[54813]_ ,
    \new_[54814]_ , \new_[54817]_ , \new_[54820]_ , \new_[54821]_ ,
    \new_[54822]_ , \new_[54826]_ , \new_[54827]_ , \new_[54831]_ ,
    \new_[54832]_ , \new_[54833]_ , \new_[54837]_ , \new_[54838]_ ,
    \new_[54841]_ , \new_[54844]_ , \new_[54845]_ , \new_[54846]_ ,
    \new_[54850]_ , \new_[54851]_ , \new_[54855]_ , \new_[54856]_ ,
    \new_[54857]_ , \new_[54861]_ , \new_[54862]_ , \new_[54865]_ ,
    \new_[54868]_ , \new_[54869]_ , \new_[54870]_ , \new_[54874]_ ,
    \new_[54875]_ , \new_[54879]_ , \new_[54880]_ , \new_[54881]_ ,
    \new_[54885]_ , \new_[54886]_ , \new_[54889]_ , \new_[54892]_ ,
    \new_[54893]_ , \new_[54894]_ , \new_[54898]_ , \new_[54899]_ ,
    \new_[54903]_ , \new_[54904]_ , \new_[54905]_ , \new_[54909]_ ,
    \new_[54910]_ , \new_[54913]_ , \new_[54916]_ , \new_[54917]_ ,
    \new_[54918]_ , \new_[54922]_ , \new_[54923]_ , \new_[54927]_ ,
    \new_[54928]_ , \new_[54929]_ , \new_[54933]_ , \new_[54934]_ ,
    \new_[54937]_ , \new_[54940]_ , \new_[54941]_ , \new_[54942]_ ,
    \new_[54946]_ , \new_[54947]_ , \new_[54951]_ , \new_[54952]_ ,
    \new_[54953]_ , \new_[54957]_ , \new_[54958]_ , \new_[54961]_ ,
    \new_[54964]_ , \new_[54965]_ , \new_[54966]_ , \new_[54970]_ ,
    \new_[54971]_ , \new_[54975]_ , \new_[54976]_ , \new_[54977]_ ,
    \new_[54981]_ , \new_[54982]_ , \new_[54985]_ , \new_[54988]_ ,
    \new_[54989]_ , \new_[54990]_ , \new_[54994]_ , \new_[54995]_ ,
    \new_[54999]_ , \new_[55000]_ , \new_[55001]_ , \new_[55005]_ ,
    \new_[55006]_ , \new_[55009]_ , \new_[55012]_ , \new_[55013]_ ,
    \new_[55014]_ , \new_[55018]_ , \new_[55019]_ , \new_[55023]_ ,
    \new_[55024]_ , \new_[55025]_ , \new_[55029]_ , \new_[55030]_ ,
    \new_[55033]_ , \new_[55036]_ , \new_[55037]_ , \new_[55038]_ ,
    \new_[55042]_ , \new_[55043]_ , \new_[55047]_ , \new_[55048]_ ,
    \new_[55049]_ , \new_[55053]_ , \new_[55054]_ , \new_[55057]_ ,
    \new_[55060]_ , \new_[55061]_ , \new_[55062]_ , \new_[55066]_ ,
    \new_[55067]_ , \new_[55071]_ , \new_[55072]_ , \new_[55073]_ ,
    \new_[55077]_ , \new_[55078]_ , \new_[55081]_ , \new_[55084]_ ,
    \new_[55085]_ , \new_[55086]_ , \new_[55090]_ , \new_[55091]_ ,
    \new_[55095]_ , \new_[55096]_ , \new_[55097]_ , \new_[55101]_ ,
    \new_[55102]_ , \new_[55105]_ , \new_[55108]_ , \new_[55109]_ ,
    \new_[55110]_ , \new_[55114]_ , \new_[55115]_ , \new_[55119]_ ,
    \new_[55120]_ , \new_[55121]_ , \new_[55125]_ , \new_[55126]_ ,
    \new_[55129]_ , \new_[55132]_ , \new_[55133]_ , \new_[55134]_ ,
    \new_[55138]_ , \new_[55139]_ , \new_[55143]_ , \new_[55144]_ ,
    \new_[55145]_ , \new_[55149]_ , \new_[55150]_ , \new_[55153]_ ,
    \new_[55156]_ , \new_[55157]_ , \new_[55158]_ , \new_[55162]_ ,
    \new_[55163]_ , \new_[55167]_ , \new_[55168]_ , \new_[55169]_ ,
    \new_[55173]_ , \new_[55174]_ , \new_[55177]_ , \new_[55180]_ ,
    \new_[55181]_ , \new_[55182]_ , \new_[55186]_ , \new_[55187]_ ,
    \new_[55191]_ , \new_[55192]_ , \new_[55193]_ , \new_[55197]_ ,
    \new_[55198]_ , \new_[55201]_ , \new_[55204]_ , \new_[55205]_ ,
    \new_[55206]_ , \new_[55210]_ , \new_[55211]_ , \new_[55215]_ ,
    \new_[55216]_ , \new_[55217]_ , \new_[55221]_ , \new_[55222]_ ,
    \new_[55225]_ , \new_[55228]_ , \new_[55229]_ , \new_[55230]_ ,
    \new_[55234]_ , \new_[55235]_ , \new_[55239]_ , \new_[55240]_ ,
    \new_[55241]_ , \new_[55245]_ , \new_[55246]_ , \new_[55249]_ ,
    \new_[55252]_ , \new_[55253]_ , \new_[55254]_ , \new_[55258]_ ,
    \new_[55259]_ , \new_[55263]_ , \new_[55264]_ , \new_[55265]_ ,
    \new_[55269]_ , \new_[55270]_ , \new_[55273]_ , \new_[55276]_ ,
    \new_[55277]_ , \new_[55278]_ , \new_[55282]_ , \new_[55283]_ ,
    \new_[55287]_ , \new_[55288]_ , \new_[55289]_ , \new_[55293]_ ,
    \new_[55294]_ , \new_[55297]_ , \new_[55300]_ , \new_[55301]_ ,
    \new_[55302]_ , \new_[55306]_ , \new_[55307]_ , \new_[55311]_ ,
    \new_[55312]_ , \new_[55313]_ , \new_[55317]_ , \new_[55318]_ ,
    \new_[55321]_ , \new_[55324]_ , \new_[55325]_ , \new_[55326]_ ,
    \new_[55330]_ , \new_[55331]_ , \new_[55335]_ , \new_[55336]_ ,
    \new_[55337]_ , \new_[55341]_ , \new_[55342]_ , \new_[55345]_ ,
    \new_[55348]_ , \new_[55349]_ , \new_[55350]_ , \new_[55354]_ ,
    \new_[55355]_ , \new_[55359]_ , \new_[55360]_ , \new_[55361]_ ,
    \new_[55365]_ , \new_[55366]_ , \new_[55369]_ , \new_[55372]_ ,
    \new_[55373]_ , \new_[55374]_ , \new_[55378]_ , \new_[55379]_ ,
    \new_[55383]_ , \new_[55384]_ , \new_[55385]_ , \new_[55389]_ ,
    \new_[55390]_ , \new_[55393]_ , \new_[55396]_ , \new_[55397]_ ,
    \new_[55398]_ , \new_[55402]_ , \new_[55403]_ , \new_[55407]_ ,
    \new_[55408]_ , \new_[55409]_ , \new_[55413]_ , \new_[55414]_ ,
    \new_[55417]_ , \new_[55420]_ , \new_[55421]_ , \new_[55422]_ ,
    \new_[55426]_ , \new_[55427]_ , \new_[55431]_ , \new_[55432]_ ,
    \new_[55433]_ , \new_[55437]_ , \new_[55438]_ , \new_[55441]_ ,
    \new_[55444]_ , \new_[55445]_ , \new_[55446]_ , \new_[55450]_ ,
    \new_[55451]_ , \new_[55455]_ , \new_[55456]_ , \new_[55457]_ ,
    \new_[55461]_ , \new_[55462]_ , \new_[55465]_ , \new_[55468]_ ,
    \new_[55469]_ , \new_[55470]_ , \new_[55474]_ , \new_[55475]_ ,
    \new_[55479]_ , \new_[55480]_ , \new_[55481]_ , \new_[55485]_ ,
    \new_[55486]_ , \new_[55489]_ , \new_[55492]_ , \new_[55493]_ ,
    \new_[55494]_ , \new_[55498]_ , \new_[55499]_ , \new_[55503]_ ,
    \new_[55504]_ , \new_[55505]_ , \new_[55509]_ , \new_[55510]_ ,
    \new_[55513]_ , \new_[55516]_ , \new_[55517]_ , \new_[55518]_ ,
    \new_[55522]_ , \new_[55523]_ , \new_[55527]_ , \new_[55528]_ ,
    \new_[55529]_ , \new_[55533]_ , \new_[55534]_ , \new_[55537]_ ,
    \new_[55540]_ , \new_[55541]_ , \new_[55542]_ , \new_[55546]_ ,
    \new_[55547]_ , \new_[55551]_ , \new_[55552]_ , \new_[55553]_ ,
    \new_[55557]_ , \new_[55558]_ , \new_[55561]_ , \new_[55564]_ ,
    \new_[55565]_ , \new_[55566]_ , \new_[55570]_ , \new_[55571]_ ,
    \new_[55575]_ , \new_[55576]_ , \new_[55577]_ , \new_[55581]_ ,
    \new_[55582]_ , \new_[55585]_ , \new_[55588]_ , \new_[55589]_ ,
    \new_[55590]_ , \new_[55594]_ , \new_[55595]_ , \new_[55599]_ ,
    \new_[55600]_ , \new_[55601]_ , \new_[55605]_ , \new_[55606]_ ,
    \new_[55609]_ , \new_[55612]_ , \new_[55613]_ , \new_[55614]_ ,
    \new_[55618]_ , \new_[55619]_ , \new_[55623]_ , \new_[55624]_ ,
    \new_[55625]_ , \new_[55629]_ , \new_[55630]_ , \new_[55633]_ ,
    \new_[55636]_ , \new_[55637]_ , \new_[55638]_ , \new_[55642]_ ,
    \new_[55643]_ , \new_[55647]_ , \new_[55648]_ , \new_[55649]_ ,
    \new_[55653]_ , \new_[55654]_ , \new_[55657]_ , \new_[55660]_ ,
    \new_[55661]_ , \new_[55662]_ , \new_[55666]_ , \new_[55667]_ ,
    \new_[55671]_ , \new_[55672]_ , \new_[55673]_ , \new_[55677]_ ,
    \new_[55678]_ , \new_[55681]_ , \new_[55684]_ , \new_[55685]_ ,
    \new_[55686]_ , \new_[55690]_ , \new_[55691]_ , \new_[55695]_ ,
    \new_[55696]_ , \new_[55697]_ , \new_[55701]_ , \new_[55702]_ ,
    \new_[55705]_ , \new_[55708]_ , \new_[55709]_ , \new_[55710]_ ,
    \new_[55714]_ , \new_[55715]_ , \new_[55719]_ , \new_[55720]_ ,
    \new_[55721]_ , \new_[55725]_ , \new_[55726]_ , \new_[55729]_ ,
    \new_[55732]_ , \new_[55733]_ , \new_[55734]_ , \new_[55738]_ ,
    \new_[55739]_ , \new_[55743]_ , \new_[55744]_ , \new_[55745]_ ,
    \new_[55749]_ , \new_[55750]_ , \new_[55753]_ , \new_[55756]_ ,
    \new_[55757]_ , \new_[55758]_ , \new_[55762]_ , \new_[55763]_ ,
    \new_[55767]_ , \new_[55768]_ , \new_[55769]_ , \new_[55773]_ ,
    \new_[55774]_ , \new_[55777]_ , \new_[55780]_ , \new_[55781]_ ,
    \new_[55782]_ , \new_[55786]_ , \new_[55787]_ , \new_[55791]_ ,
    \new_[55792]_ , \new_[55793]_ , \new_[55797]_ , \new_[55798]_ ,
    \new_[55801]_ , \new_[55804]_ , \new_[55805]_ , \new_[55806]_ ,
    \new_[55810]_ , \new_[55811]_ , \new_[55815]_ , \new_[55816]_ ,
    \new_[55817]_ , \new_[55821]_ , \new_[55822]_ , \new_[55825]_ ,
    \new_[55828]_ , \new_[55829]_ , \new_[55830]_ , \new_[55834]_ ,
    \new_[55835]_ , \new_[55839]_ , \new_[55840]_ , \new_[55841]_ ,
    \new_[55845]_ , \new_[55846]_ , \new_[55849]_ , \new_[55852]_ ,
    \new_[55853]_ , \new_[55854]_ , \new_[55858]_ , \new_[55859]_ ,
    \new_[55863]_ , \new_[55864]_ , \new_[55865]_ , \new_[55869]_ ,
    \new_[55870]_ , \new_[55873]_ , \new_[55876]_ , \new_[55877]_ ,
    \new_[55878]_ , \new_[55882]_ , \new_[55883]_ , \new_[55887]_ ,
    \new_[55888]_ , \new_[55889]_ , \new_[55893]_ , \new_[55894]_ ,
    \new_[55897]_ , \new_[55900]_ , \new_[55901]_ , \new_[55902]_ ,
    \new_[55906]_ , \new_[55907]_ , \new_[55911]_ , \new_[55912]_ ,
    \new_[55913]_ , \new_[55917]_ , \new_[55918]_ , \new_[55921]_ ,
    \new_[55924]_ , \new_[55925]_ , \new_[55926]_ , \new_[55930]_ ,
    \new_[55931]_ , \new_[55935]_ , \new_[55936]_ , \new_[55937]_ ,
    \new_[55941]_ , \new_[55942]_ , \new_[55945]_ , \new_[55948]_ ,
    \new_[55949]_ , \new_[55950]_ , \new_[55954]_ , \new_[55955]_ ,
    \new_[55959]_ , \new_[55960]_ , \new_[55961]_ , \new_[55965]_ ,
    \new_[55966]_ , \new_[55969]_ , \new_[55972]_ , \new_[55973]_ ,
    \new_[55974]_ , \new_[55978]_ , \new_[55979]_ , \new_[55983]_ ,
    \new_[55984]_ , \new_[55985]_ , \new_[55989]_ , \new_[55990]_ ,
    \new_[55993]_ , \new_[55996]_ , \new_[55997]_ , \new_[55998]_ ,
    \new_[56002]_ , \new_[56003]_ , \new_[56007]_ , \new_[56008]_ ,
    \new_[56009]_ , \new_[56013]_ , \new_[56014]_ , \new_[56017]_ ,
    \new_[56020]_ , \new_[56021]_ , \new_[56022]_ , \new_[56026]_ ,
    \new_[56027]_ , \new_[56031]_ , \new_[56032]_ , \new_[56033]_ ,
    \new_[56037]_ , \new_[56038]_ , \new_[56041]_ , \new_[56044]_ ,
    \new_[56045]_ , \new_[56046]_ , \new_[56050]_ , \new_[56051]_ ,
    \new_[56055]_ , \new_[56056]_ , \new_[56057]_ , \new_[56061]_ ,
    \new_[56062]_ , \new_[56065]_ , \new_[56068]_ , \new_[56069]_ ,
    \new_[56070]_ , \new_[56074]_ , \new_[56075]_ , \new_[56079]_ ,
    \new_[56080]_ , \new_[56081]_ , \new_[56085]_ , \new_[56086]_ ,
    \new_[56089]_ , \new_[56092]_ , \new_[56093]_ , \new_[56094]_ ,
    \new_[56098]_ , \new_[56099]_ , \new_[56103]_ , \new_[56104]_ ,
    \new_[56105]_ , \new_[56109]_ , \new_[56110]_ , \new_[56113]_ ,
    \new_[56116]_ , \new_[56117]_ , \new_[56118]_ , \new_[56122]_ ,
    \new_[56123]_ , \new_[56127]_ , \new_[56128]_ , \new_[56129]_ ,
    \new_[56133]_ , \new_[56134]_ , \new_[56137]_ , \new_[56140]_ ,
    \new_[56141]_ , \new_[56142]_ , \new_[56146]_ , \new_[56147]_ ,
    \new_[56151]_ , \new_[56152]_ , \new_[56153]_ , \new_[56157]_ ,
    \new_[56158]_ , \new_[56161]_ , \new_[56164]_ , \new_[56165]_ ,
    \new_[56166]_ , \new_[56170]_ , \new_[56171]_ , \new_[56175]_ ,
    \new_[56176]_ , \new_[56177]_ , \new_[56181]_ , \new_[56182]_ ,
    \new_[56185]_ , \new_[56188]_ , \new_[56189]_ , \new_[56190]_ ,
    \new_[56194]_ , \new_[56195]_ , \new_[56199]_ , \new_[56200]_ ,
    \new_[56201]_ , \new_[56205]_ , \new_[56206]_ , \new_[56209]_ ,
    \new_[56212]_ , \new_[56213]_ , \new_[56214]_ , \new_[56218]_ ,
    \new_[56219]_ , \new_[56223]_ , \new_[56224]_ , \new_[56225]_ ,
    \new_[56229]_ , \new_[56230]_ , \new_[56233]_ , \new_[56236]_ ,
    \new_[56237]_ , \new_[56238]_ , \new_[56242]_ , \new_[56243]_ ,
    \new_[56247]_ , \new_[56248]_ , \new_[56249]_ , \new_[56253]_ ,
    \new_[56254]_ , \new_[56257]_ , \new_[56260]_ , \new_[56261]_ ,
    \new_[56262]_ , \new_[56266]_ , \new_[56267]_ , \new_[56271]_ ,
    \new_[56272]_ , \new_[56273]_ , \new_[56277]_ , \new_[56278]_ ,
    \new_[56281]_ , \new_[56284]_ , \new_[56285]_ , \new_[56286]_ ,
    \new_[56290]_ , \new_[56291]_ , \new_[56295]_ , \new_[56296]_ ,
    \new_[56297]_ , \new_[56301]_ , \new_[56302]_ , \new_[56305]_ ,
    \new_[56308]_ , \new_[56309]_ , \new_[56310]_ , \new_[56314]_ ,
    \new_[56315]_ , \new_[56319]_ , \new_[56320]_ , \new_[56321]_ ,
    \new_[56325]_ , \new_[56326]_ , \new_[56329]_ , \new_[56332]_ ,
    \new_[56333]_ , \new_[56334]_ , \new_[56338]_ , \new_[56339]_ ,
    \new_[56343]_ , \new_[56344]_ , \new_[56345]_ , \new_[56349]_ ,
    \new_[56350]_ , \new_[56353]_ , \new_[56356]_ , \new_[56357]_ ,
    \new_[56358]_ , \new_[56362]_ , \new_[56363]_ , \new_[56367]_ ,
    \new_[56368]_ , \new_[56369]_ , \new_[56373]_ , \new_[56374]_ ,
    \new_[56377]_ , \new_[56380]_ , \new_[56381]_ , \new_[56382]_ ,
    \new_[56386]_ , \new_[56387]_ , \new_[56391]_ , \new_[56392]_ ,
    \new_[56393]_ , \new_[56397]_ , \new_[56398]_ , \new_[56401]_ ,
    \new_[56404]_ , \new_[56405]_ , \new_[56406]_ , \new_[56410]_ ,
    \new_[56411]_ , \new_[56415]_ , \new_[56416]_ , \new_[56417]_ ,
    \new_[56421]_ , \new_[56422]_ , \new_[56425]_ , \new_[56428]_ ,
    \new_[56429]_ , \new_[56430]_ , \new_[56434]_ , \new_[56435]_ ,
    \new_[56439]_ , \new_[56440]_ , \new_[56441]_ , \new_[56445]_ ,
    \new_[56446]_ , \new_[56449]_ , \new_[56452]_ , \new_[56453]_ ,
    \new_[56454]_ , \new_[56458]_ , \new_[56459]_ , \new_[56463]_ ,
    \new_[56464]_ , \new_[56465]_ , \new_[56469]_ , \new_[56470]_ ,
    \new_[56473]_ , \new_[56476]_ , \new_[56477]_ , \new_[56478]_ ,
    \new_[56482]_ , \new_[56483]_ , \new_[56487]_ , \new_[56488]_ ,
    \new_[56489]_ , \new_[56493]_ , \new_[56494]_ , \new_[56497]_ ,
    \new_[56500]_ , \new_[56501]_ , \new_[56502]_ , \new_[56506]_ ,
    \new_[56507]_ , \new_[56511]_ , \new_[56512]_ , \new_[56513]_ ,
    \new_[56517]_ , \new_[56518]_ , \new_[56521]_ , \new_[56524]_ ,
    \new_[56525]_ , \new_[56526]_ , \new_[56530]_ , \new_[56531]_ ,
    \new_[56535]_ , \new_[56536]_ , \new_[56537]_ , \new_[56541]_ ,
    \new_[56542]_ , \new_[56545]_ , \new_[56548]_ , \new_[56549]_ ,
    \new_[56550]_ , \new_[56554]_ , \new_[56555]_ , \new_[56559]_ ,
    \new_[56560]_ , \new_[56561]_ , \new_[56565]_ , \new_[56566]_ ,
    \new_[56569]_ , \new_[56572]_ , \new_[56573]_ , \new_[56574]_ ,
    \new_[56578]_ , \new_[56579]_ , \new_[56583]_ , \new_[56584]_ ,
    \new_[56585]_ , \new_[56589]_ , \new_[56590]_ , \new_[56593]_ ,
    \new_[56596]_ , \new_[56597]_ , \new_[56598]_ , \new_[56602]_ ,
    \new_[56603]_ , \new_[56607]_ , \new_[56608]_ , \new_[56609]_ ,
    \new_[56613]_ , \new_[56614]_ , \new_[56617]_ , \new_[56620]_ ,
    \new_[56621]_ , \new_[56622]_ , \new_[56626]_ , \new_[56627]_ ,
    \new_[56631]_ , \new_[56632]_ , \new_[56633]_ , \new_[56637]_ ,
    \new_[56638]_ , \new_[56641]_ , \new_[56644]_ , \new_[56645]_ ,
    \new_[56646]_ , \new_[56650]_ , \new_[56651]_ , \new_[56655]_ ,
    \new_[56656]_ , \new_[56657]_ , \new_[56661]_ , \new_[56662]_ ,
    \new_[56665]_ , \new_[56668]_ , \new_[56669]_ , \new_[56670]_ ,
    \new_[56674]_ , \new_[56675]_ , \new_[56679]_ , \new_[56680]_ ,
    \new_[56681]_ , \new_[56685]_ , \new_[56686]_ , \new_[56689]_ ,
    \new_[56692]_ , \new_[56693]_ , \new_[56694]_ , \new_[56698]_ ,
    \new_[56699]_ , \new_[56703]_ , \new_[56704]_ , \new_[56705]_ ,
    \new_[56709]_ , \new_[56710]_ , \new_[56713]_ , \new_[56716]_ ,
    \new_[56717]_ , \new_[56718]_ , \new_[56722]_ , \new_[56723]_ ,
    \new_[56727]_ , \new_[56728]_ , \new_[56729]_ , \new_[56733]_ ,
    \new_[56734]_ , \new_[56737]_ , \new_[56740]_ , \new_[56741]_ ,
    \new_[56742]_ , \new_[56746]_ , \new_[56747]_ , \new_[56751]_ ,
    \new_[56752]_ , \new_[56753]_ , \new_[56757]_ , \new_[56758]_ ,
    \new_[56761]_ , \new_[56764]_ , \new_[56765]_ , \new_[56766]_ ,
    \new_[56770]_ , \new_[56771]_ , \new_[56775]_ , \new_[56776]_ ,
    \new_[56777]_ , \new_[56781]_ , \new_[56782]_ , \new_[56785]_ ,
    \new_[56788]_ , \new_[56789]_ , \new_[56790]_ , \new_[56794]_ ,
    \new_[56795]_ , \new_[56799]_ , \new_[56800]_ , \new_[56801]_ ,
    \new_[56805]_ , \new_[56806]_ , \new_[56809]_ , \new_[56812]_ ,
    \new_[56813]_ , \new_[56814]_ , \new_[56818]_ , \new_[56819]_ ,
    \new_[56823]_ , \new_[56824]_ , \new_[56825]_ , \new_[56829]_ ,
    \new_[56830]_ , \new_[56833]_ , \new_[56836]_ , \new_[56837]_ ,
    \new_[56838]_ , \new_[56842]_ , \new_[56843]_ , \new_[56847]_ ,
    \new_[56848]_ , \new_[56849]_ , \new_[56853]_ , \new_[56854]_ ,
    \new_[56857]_ , \new_[56860]_ , \new_[56861]_ , \new_[56862]_ ,
    \new_[56866]_ , \new_[56867]_ , \new_[56871]_ , \new_[56872]_ ,
    \new_[56873]_ , \new_[56877]_ , \new_[56878]_ , \new_[56881]_ ,
    \new_[56884]_ , \new_[56885]_ , \new_[56886]_ , \new_[56890]_ ,
    \new_[56891]_ , \new_[56895]_ , \new_[56896]_ , \new_[56897]_ ,
    \new_[56901]_ , \new_[56902]_ , \new_[56905]_ , \new_[56908]_ ,
    \new_[56909]_ , \new_[56910]_ , \new_[56914]_ , \new_[56915]_ ,
    \new_[56919]_ , \new_[56920]_ , \new_[56921]_ , \new_[56925]_ ,
    \new_[56926]_ , \new_[56929]_ , \new_[56932]_ , \new_[56933]_ ,
    \new_[56934]_ , \new_[56938]_ , \new_[56939]_ , \new_[56943]_ ,
    \new_[56944]_ , \new_[56945]_ , \new_[56949]_ , \new_[56950]_ ,
    \new_[56953]_ , \new_[56956]_ , \new_[56957]_ , \new_[56958]_ ,
    \new_[56962]_ , \new_[56963]_ , \new_[56967]_ , \new_[56968]_ ,
    \new_[56969]_ , \new_[56973]_ , \new_[56974]_ , \new_[56977]_ ,
    \new_[56980]_ , \new_[56981]_ , \new_[56982]_ , \new_[56986]_ ,
    \new_[56987]_ , \new_[56991]_ , \new_[56992]_ , \new_[56993]_ ,
    \new_[56997]_ , \new_[56998]_ , \new_[57001]_ , \new_[57004]_ ,
    \new_[57005]_ , \new_[57006]_ , \new_[57010]_ , \new_[57011]_ ,
    \new_[57015]_ , \new_[57016]_ , \new_[57017]_ , \new_[57021]_ ,
    \new_[57022]_ , \new_[57025]_ , \new_[57028]_ , \new_[57029]_ ,
    \new_[57030]_ , \new_[57034]_ , \new_[57035]_ , \new_[57039]_ ,
    \new_[57040]_ , \new_[57041]_ , \new_[57045]_ , \new_[57046]_ ,
    \new_[57049]_ , \new_[57052]_ , \new_[57053]_ , \new_[57054]_ ,
    \new_[57058]_ , \new_[57059]_ , \new_[57063]_ , \new_[57064]_ ,
    \new_[57065]_ , \new_[57069]_ , \new_[57070]_ , \new_[57073]_ ,
    \new_[57076]_ , \new_[57077]_ , \new_[57078]_ , \new_[57082]_ ,
    \new_[57083]_ , \new_[57087]_ , \new_[57088]_ , \new_[57089]_ ,
    \new_[57093]_ , \new_[57094]_ , \new_[57097]_ , \new_[57100]_ ,
    \new_[57101]_ , \new_[57102]_ , \new_[57106]_ , \new_[57107]_ ,
    \new_[57111]_ , \new_[57112]_ , \new_[57113]_ , \new_[57117]_ ,
    \new_[57118]_ , \new_[57121]_ , \new_[57124]_ , \new_[57125]_ ,
    \new_[57126]_ , \new_[57130]_ , \new_[57131]_ , \new_[57135]_ ,
    \new_[57136]_ , \new_[57137]_ , \new_[57141]_ , \new_[57142]_ ,
    \new_[57145]_ , \new_[57148]_ , \new_[57149]_ , \new_[57150]_ ,
    \new_[57154]_ , \new_[57155]_ , \new_[57159]_ , \new_[57160]_ ,
    \new_[57161]_ , \new_[57165]_ , \new_[57166]_ , \new_[57169]_ ,
    \new_[57172]_ , \new_[57173]_ , \new_[57174]_ , \new_[57178]_ ,
    \new_[57179]_ , \new_[57183]_ , \new_[57184]_ , \new_[57185]_ ,
    \new_[57189]_ , \new_[57190]_ , \new_[57193]_ , \new_[57196]_ ,
    \new_[57197]_ , \new_[57198]_ , \new_[57202]_ , \new_[57203]_ ,
    \new_[57207]_ , \new_[57208]_ , \new_[57209]_ , \new_[57213]_ ,
    \new_[57214]_ , \new_[57217]_ , \new_[57220]_ , \new_[57221]_ ,
    \new_[57222]_ , \new_[57226]_ , \new_[57227]_ , \new_[57231]_ ,
    \new_[57232]_ , \new_[57233]_ , \new_[57237]_ , \new_[57238]_ ,
    \new_[57241]_ , \new_[57244]_ , \new_[57245]_ , \new_[57246]_ ,
    \new_[57250]_ , \new_[57251]_ , \new_[57255]_ , \new_[57256]_ ,
    \new_[57257]_ , \new_[57261]_ , \new_[57262]_ , \new_[57265]_ ,
    \new_[57268]_ , \new_[57269]_ , \new_[57270]_ , \new_[57274]_ ,
    \new_[57275]_ , \new_[57279]_ , \new_[57280]_ , \new_[57281]_ ,
    \new_[57285]_ , \new_[57286]_ , \new_[57289]_ , \new_[57292]_ ,
    \new_[57293]_ , \new_[57294]_ , \new_[57298]_ , \new_[57299]_ ,
    \new_[57303]_ , \new_[57304]_ , \new_[57305]_ , \new_[57309]_ ,
    \new_[57310]_ , \new_[57313]_ , \new_[57316]_ , \new_[57317]_ ,
    \new_[57318]_ , \new_[57322]_ , \new_[57323]_ , \new_[57327]_ ,
    \new_[57328]_ , \new_[57329]_ , \new_[57333]_ , \new_[57334]_ ,
    \new_[57337]_ , \new_[57340]_ , \new_[57341]_ , \new_[57342]_ ,
    \new_[57346]_ , \new_[57347]_ , \new_[57351]_ , \new_[57352]_ ,
    \new_[57353]_ , \new_[57357]_ , \new_[57358]_ , \new_[57361]_ ,
    \new_[57364]_ , \new_[57365]_ , \new_[57366]_ , \new_[57370]_ ,
    \new_[57371]_ , \new_[57375]_ , \new_[57376]_ , \new_[57377]_ ,
    \new_[57381]_ , \new_[57382]_ , \new_[57385]_ , \new_[57388]_ ,
    \new_[57389]_ , \new_[57390]_ , \new_[57394]_ , \new_[57395]_ ,
    \new_[57399]_ , \new_[57400]_ , \new_[57401]_ , \new_[57405]_ ,
    \new_[57406]_ , \new_[57409]_ , \new_[57412]_ , \new_[57413]_ ,
    \new_[57414]_ , \new_[57418]_ , \new_[57419]_ , \new_[57423]_ ,
    \new_[57424]_ , \new_[57425]_ , \new_[57429]_ , \new_[57430]_ ,
    \new_[57433]_ , \new_[57436]_ , \new_[57437]_ , \new_[57438]_ ,
    \new_[57442]_ , \new_[57443]_ , \new_[57447]_ , \new_[57448]_ ,
    \new_[57449]_ , \new_[57453]_ , \new_[57454]_ , \new_[57457]_ ,
    \new_[57460]_ , \new_[57461]_ , \new_[57462]_ , \new_[57466]_ ,
    \new_[57467]_ , \new_[57471]_ , \new_[57472]_ , \new_[57473]_ ,
    \new_[57477]_ , \new_[57478]_ , \new_[57481]_ , \new_[57484]_ ,
    \new_[57485]_ , \new_[57486]_ , \new_[57490]_ , \new_[57491]_ ,
    \new_[57495]_ , \new_[57496]_ , \new_[57497]_ , \new_[57501]_ ,
    \new_[57502]_ , \new_[57505]_ , \new_[57508]_ , \new_[57509]_ ,
    \new_[57510]_ , \new_[57514]_ , \new_[57515]_ , \new_[57519]_ ,
    \new_[57520]_ , \new_[57521]_ , \new_[57525]_ , \new_[57526]_ ,
    \new_[57529]_ , \new_[57532]_ , \new_[57533]_ , \new_[57534]_ ,
    \new_[57538]_ , \new_[57539]_ , \new_[57543]_ , \new_[57544]_ ,
    \new_[57545]_ , \new_[57549]_ , \new_[57550]_ , \new_[57553]_ ,
    \new_[57556]_ , \new_[57557]_ , \new_[57558]_ , \new_[57562]_ ,
    \new_[57563]_ , \new_[57567]_ , \new_[57568]_ , \new_[57569]_ ,
    \new_[57573]_ , \new_[57574]_ , \new_[57577]_ , \new_[57580]_ ,
    \new_[57581]_ , \new_[57582]_ , \new_[57586]_ , \new_[57587]_ ,
    \new_[57591]_ , \new_[57592]_ , \new_[57593]_ , \new_[57597]_ ,
    \new_[57598]_ , \new_[57601]_ , \new_[57604]_ , \new_[57605]_ ,
    \new_[57606]_ , \new_[57610]_ , \new_[57611]_ , \new_[57615]_ ,
    \new_[57616]_ , \new_[57617]_ , \new_[57621]_ , \new_[57622]_ ,
    \new_[57625]_ , \new_[57628]_ , \new_[57629]_ , \new_[57630]_ ,
    \new_[57634]_ , \new_[57635]_ , \new_[57639]_ , \new_[57640]_ ,
    \new_[57641]_ , \new_[57645]_ , \new_[57646]_ , \new_[57649]_ ,
    \new_[57652]_ , \new_[57653]_ , \new_[57654]_ , \new_[57658]_ ,
    \new_[57659]_ , \new_[57663]_ , \new_[57664]_ , \new_[57665]_ ,
    \new_[57669]_ , \new_[57670]_ , \new_[57673]_ , \new_[57676]_ ,
    \new_[57677]_ , \new_[57678]_ , \new_[57682]_ , \new_[57683]_ ,
    \new_[57687]_ , \new_[57688]_ , \new_[57689]_ , \new_[57693]_ ,
    \new_[57694]_ , \new_[57697]_ , \new_[57700]_ , \new_[57701]_ ,
    \new_[57702]_ , \new_[57706]_ , \new_[57707]_ , \new_[57711]_ ,
    \new_[57712]_ , \new_[57713]_ , \new_[57717]_ , \new_[57718]_ ,
    \new_[57721]_ , \new_[57724]_ , \new_[57725]_ , \new_[57726]_ ,
    \new_[57730]_ , \new_[57731]_ , \new_[57735]_ , \new_[57736]_ ,
    \new_[57737]_ , \new_[57741]_ , \new_[57742]_ , \new_[57745]_ ,
    \new_[57748]_ , \new_[57749]_ , \new_[57750]_ , \new_[57754]_ ,
    \new_[57755]_ , \new_[57759]_ , \new_[57760]_ , \new_[57761]_ ,
    \new_[57765]_ , \new_[57766]_ , \new_[57769]_ , \new_[57772]_ ,
    \new_[57773]_ , \new_[57774]_ , \new_[57778]_ , \new_[57779]_ ,
    \new_[57783]_ , \new_[57784]_ , \new_[57785]_ , \new_[57789]_ ,
    \new_[57790]_ , \new_[57793]_ , \new_[57796]_ , \new_[57797]_ ,
    \new_[57798]_ , \new_[57802]_ , \new_[57803]_ , \new_[57807]_ ,
    \new_[57808]_ , \new_[57809]_ , \new_[57813]_ , \new_[57814]_ ,
    \new_[57817]_ , \new_[57820]_ , \new_[57821]_ , \new_[57822]_ ,
    \new_[57826]_ , \new_[57827]_ , \new_[57831]_ , \new_[57832]_ ,
    \new_[57833]_ , \new_[57837]_ , \new_[57838]_ , \new_[57841]_ ,
    \new_[57844]_ , \new_[57845]_ , \new_[57846]_ , \new_[57850]_ ,
    \new_[57851]_ , \new_[57855]_ , \new_[57856]_ , \new_[57857]_ ,
    \new_[57861]_ , \new_[57862]_ , \new_[57865]_ , \new_[57868]_ ,
    \new_[57869]_ , \new_[57870]_ , \new_[57874]_ , \new_[57875]_ ,
    \new_[57879]_ , \new_[57880]_ , \new_[57881]_ , \new_[57885]_ ,
    \new_[57886]_ , \new_[57889]_ , \new_[57892]_ , \new_[57893]_ ,
    \new_[57894]_ , \new_[57898]_ , \new_[57899]_ , \new_[57903]_ ,
    \new_[57904]_ , \new_[57905]_ , \new_[57909]_ , \new_[57910]_ ,
    \new_[57913]_ , \new_[57916]_ , \new_[57917]_ , \new_[57918]_ ,
    \new_[57922]_ , \new_[57923]_ , \new_[57927]_ , \new_[57928]_ ,
    \new_[57929]_ , \new_[57933]_ , \new_[57934]_ , \new_[57937]_ ,
    \new_[57940]_ , \new_[57941]_ , \new_[57942]_ , \new_[57946]_ ,
    \new_[57947]_ , \new_[57951]_ , \new_[57952]_ , \new_[57953]_ ,
    \new_[57957]_ , \new_[57958]_ , \new_[57961]_ , \new_[57964]_ ,
    \new_[57965]_ , \new_[57966]_ , \new_[57970]_ , \new_[57971]_ ,
    \new_[57975]_ , \new_[57976]_ , \new_[57977]_ , \new_[57981]_ ,
    \new_[57982]_ , \new_[57985]_ , \new_[57988]_ , \new_[57989]_ ,
    \new_[57990]_ , \new_[57994]_ , \new_[57995]_ , \new_[57999]_ ,
    \new_[58000]_ , \new_[58001]_ , \new_[58005]_ , \new_[58006]_ ,
    \new_[58009]_ , \new_[58012]_ , \new_[58013]_ , \new_[58014]_ ,
    \new_[58018]_ , \new_[58019]_ , \new_[58023]_ , \new_[58024]_ ,
    \new_[58025]_ , \new_[58029]_ , \new_[58030]_ , \new_[58033]_ ,
    \new_[58036]_ , \new_[58037]_ , \new_[58038]_ , \new_[58042]_ ,
    \new_[58043]_ , \new_[58047]_ , \new_[58048]_ , \new_[58049]_ ,
    \new_[58053]_ , \new_[58054]_ , \new_[58057]_ , \new_[58060]_ ,
    \new_[58061]_ , \new_[58062]_ , \new_[58066]_ , \new_[58067]_ ,
    \new_[58071]_ , \new_[58072]_ , \new_[58073]_ , \new_[58077]_ ,
    \new_[58078]_ , \new_[58081]_ , \new_[58084]_ , \new_[58085]_ ,
    \new_[58086]_ , \new_[58090]_ , \new_[58091]_ , \new_[58095]_ ,
    \new_[58096]_ , \new_[58097]_ , \new_[58101]_ , \new_[58102]_ ,
    \new_[58105]_ , \new_[58108]_ , \new_[58109]_ , \new_[58110]_ ,
    \new_[58114]_ , \new_[58115]_ , \new_[58119]_ , \new_[58120]_ ,
    \new_[58121]_ , \new_[58125]_ , \new_[58126]_ , \new_[58129]_ ,
    \new_[58132]_ , \new_[58133]_ , \new_[58134]_ , \new_[58138]_ ,
    \new_[58139]_ , \new_[58143]_ , \new_[58144]_ , \new_[58145]_ ,
    \new_[58149]_ , \new_[58150]_ , \new_[58153]_ , \new_[58156]_ ,
    \new_[58157]_ , \new_[58158]_ , \new_[58162]_ , \new_[58163]_ ,
    \new_[58167]_ , \new_[58168]_ , \new_[58169]_ , \new_[58173]_ ,
    \new_[58174]_ , \new_[58177]_ , \new_[58180]_ , \new_[58181]_ ,
    \new_[58182]_ , \new_[58186]_ , \new_[58187]_ , \new_[58191]_ ,
    \new_[58192]_ , \new_[58193]_ , \new_[58197]_ , \new_[58198]_ ,
    \new_[58201]_ , \new_[58204]_ , \new_[58205]_ , \new_[58206]_ ,
    \new_[58210]_ , \new_[58211]_ , \new_[58215]_ , \new_[58216]_ ,
    \new_[58217]_ , \new_[58221]_ , \new_[58222]_ , \new_[58225]_ ,
    \new_[58228]_ , \new_[58229]_ , \new_[58230]_ , \new_[58234]_ ,
    \new_[58235]_ , \new_[58239]_ , \new_[58240]_ , \new_[58241]_ ,
    \new_[58245]_ , \new_[58246]_ , \new_[58249]_ , \new_[58252]_ ,
    \new_[58253]_ , \new_[58254]_ , \new_[58258]_ , \new_[58259]_ ,
    \new_[58263]_ , \new_[58264]_ , \new_[58265]_ , \new_[58269]_ ,
    \new_[58270]_ , \new_[58273]_ , \new_[58276]_ , \new_[58277]_ ,
    \new_[58278]_ , \new_[58282]_ , \new_[58283]_ , \new_[58287]_ ,
    \new_[58288]_ , \new_[58289]_ , \new_[58293]_ , \new_[58294]_ ,
    \new_[58297]_ , \new_[58300]_ , \new_[58301]_ , \new_[58302]_ ,
    \new_[58306]_ , \new_[58307]_ , \new_[58311]_ , \new_[58312]_ ,
    \new_[58313]_ , \new_[58317]_ , \new_[58318]_ , \new_[58321]_ ,
    \new_[58324]_ , \new_[58325]_ , \new_[58326]_ , \new_[58330]_ ,
    \new_[58331]_ , \new_[58335]_ , \new_[58336]_ , \new_[58337]_ ,
    \new_[58341]_ , \new_[58342]_ , \new_[58345]_ , \new_[58348]_ ,
    \new_[58349]_ , \new_[58350]_ , \new_[58354]_ , \new_[58355]_ ,
    \new_[58359]_ , \new_[58360]_ , \new_[58361]_ , \new_[58365]_ ,
    \new_[58366]_ , \new_[58369]_ , \new_[58372]_ , \new_[58373]_ ,
    \new_[58374]_ , \new_[58378]_ , \new_[58379]_ , \new_[58383]_ ,
    \new_[58384]_ , \new_[58385]_ , \new_[58389]_ , \new_[58390]_ ,
    \new_[58393]_ , \new_[58396]_ , \new_[58397]_ , \new_[58398]_ ,
    \new_[58402]_ , \new_[58403]_ , \new_[58407]_ , \new_[58408]_ ,
    \new_[58409]_ , \new_[58413]_ , \new_[58414]_ , \new_[58417]_ ,
    \new_[58420]_ , \new_[58421]_ , \new_[58422]_ , \new_[58426]_ ,
    \new_[58427]_ , \new_[58431]_ , \new_[58432]_ , \new_[58433]_ ,
    \new_[58437]_ , \new_[58438]_ , \new_[58441]_ , \new_[58444]_ ,
    \new_[58445]_ , \new_[58446]_ , \new_[58450]_ , \new_[58451]_ ,
    \new_[58455]_ , \new_[58456]_ , \new_[58457]_ , \new_[58461]_ ,
    \new_[58462]_ , \new_[58465]_ , \new_[58468]_ , \new_[58469]_ ,
    \new_[58470]_ , \new_[58474]_ , \new_[58475]_ , \new_[58479]_ ,
    \new_[58480]_ , \new_[58481]_ , \new_[58485]_ , \new_[58486]_ ,
    \new_[58489]_ , \new_[58492]_ , \new_[58493]_ , \new_[58494]_ ,
    \new_[58498]_ , \new_[58499]_ , \new_[58503]_ , \new_[58504]_ ,
    \new_[58505]_ , \new_[58509]_ , \new_[58510]_ , \new_[58513]_ ,
    \new_[58516]_ , \new_[58517]_ , \new_[58518]_ , \new_[58522]_ ,
    \new_[58523]_ , \new_[58527]_ , \new_[58528]_ , \new_[58529]_ ,
    \new_[58533]_ , \new_[58534]_ , \new_[58537]_ , \new_[58540]_ ,
    \new_[58541]_ , \new_[58542]_ , \new_[58546]_ , \new_[58547]_ ,
    \new_[58551]_ , \new_[58552]_ , \new_[58553]_ , \new_[58557]_ ,
    \new_[58558]_ , \new_[58561]_ , \new_[58564]_ , \new_[58565]_ ,
    \new_[58566]_ , \new_[58570]_ , \new_[58571]_ , \new_[58575]_ ,
    \new_[58576]_ , \new_[58577]_ , \new_[58581]_ , \new_[58582]_ ,
    \new_[58585]_ , \new_[58588]_ , \new_[58589]_ , \new_[58590]_ ,
    \new_[58594]_ , \new_[58595]_ , \new_[58599]_ , \new_[58600]_ ,
    \new_[58601]_ , \new_[58605]_ , \new_[58606]_ , \new_[58609]_ ,
    \new_[58612]_ , \new_[58613]_ , \new_[58614]_ , \new_[58618]_ ,
    \new_[58619]_ , \new_[58623]_ , \new_[58624]_ , \new_[58625]_ ,
    \new_[58629]_ , \new_[58630]_ , \new_[58633]_ , \new_[58636]_ ,
    \new_[58637]_ , \new_[58638]_ , \new_[58642]_ , \new_[58643]_ ,
    \new_[58647]_ , \new_[58648]_ , \new_[58649]_ , \new_[58653]_ ,
    \new_[58654]_ , \new_[58657]_ , \new_[58660]_ , \new_[58661]_ ,
    \new_[58662]_ , \new_[58666]_ , \new_[58667]_ , \new_[58671]_ ,
    \new_[58672]_ , \new_[58673]_ , \new_[58677]_ , \new_[58678]_ ,
    \new_[58681]_ , \new_[58684]_ , \new_[58685]_ , \new_[58686]_ ,
    \new_[58690]_ , \new_[58691]_ , \new_[58695]_ , \new_[58696]_ ,
    \new_[58697]_ , \new_[58701]_ , \new_[58702]_ , \new_[58705]_ ,
    \new_[58708]_ , \new_[58709]_ , \new_[58710]_ , \new_[58714]_ ,
    \new_[58715]_ , \new_[58719]_ , \new_[58720]_ , \new_[58721]_ ,
    \new_[58725]_ , \new_[58726]_ , \new_[58729]_ , \new_[58732]_ ,
    \new_[58733]_ , \new_[58734]_ , \new_[58738]_ , \new_[58739]_ ,
    \new_[58743]_ , \new_[58744]_ , \new_[58745]_ , \new_[58749]_ ,
    \new_[58750]_ , \new_[58753]_ , \new_[58756]_ , \new_[58757]_ ,
    \new_[58758]_ , \new_[58762]_ , \new_[58763]_ , \new_[58767]_ ,
    \new_[58768]_ , \new_[58769]_ , \new_[58773]_ , \new_[58774]_ ,
    \new_[58777]_ , \new_[58780]_ , \new_[58781]_ , \new_[58782]_ ,
    \new_[58786]_ , \new_[58787]_ , \new_[58791]_ , \new_[58792]_ ,
    \new_[58793]_ , \new_[58797]_ , \new_[58798]_ , \new_[58801]_ ,
    \new_[58804]_ , \new_[58805]_ , \new_[58806]_ , \new_[58810]_ ,
    \new_[58811]_ , \new_[58815]_ , \new_[58816]_ , \new_[58817]_ ,
    \new_[58821]_ , \new_[58822]_ , \new_[58825]_ , \new_[58828]_ ,
    \new_[58829]_ , \new_[58830]_ , \new_[58834]_ , \new_[58835]_ ,
    \new_[58839]_ , \new_[58840]_ , \new_[58841]_ , \new_[58845]_ ,
    \new_[58846]_ , \new_[58849]_ , \new_[58852]_ , \new_[58853]_ ,
    \new_[58854]_ , \new_[58858]_ , \new_[58859]_ , \new_[58863]_ ,
    \new_[58864]_ , \new_[58865]_ , \new_[58869]_ , \new_[58870]_ ,
    \new_[58873]_ , \new_[58876]_ , \new_[58877]_ , \new_[58878]_ ,
    \new_[58882]_ , \new_[58883]_ , \new_[58887]_ , \new_[58888]_ ,
    \new_[58889]_ , \new_[58893]_ , \new_[58894]_ , \new_[58897]_ ,
    \new_[58900]_ , \new_[58901]_ , \new_[58902]_ , \new_[58906]_ ,
    \new_[58907]_ , \new_[58911]_ , \new_[58912]_ , \new_[58913]_ ,
    \new_[58917]_ , \new_[58918]_ , \new_[58921]_ , \new_[58924]_ ,
    \new_[58925]_ , \new_[58926]_ , \new_[58930]_ , \new_[58931]_ ,
    \new_[58935]_ , \new_[58936]_ , \new_[58937]_ , \new_[58941]_ ,
    \new_[58942]_ , \new_[58945]_ , \new_[58948]_ , \new_[58949]_ ,
    \new_[58950]_ , \new_[58954]_ , \new_[58955]_ , \new_[58959]_ ,
    \new_[58960]_ , \new_[58961]_ , \new_[58965]_ , \new_[58966]_ ,
    \new_[58969]_ , \new_[58972]_ , \new_[58973]_ , \new_[58974]_ ,
    \new_[58978]_ , \new_[58979]_ , \new_[58983]_ , \new_[58984]_ ,
    \new_[58985]_ , \new_[58989]_ , \new_[58990]_ , \new_[58993]_ ,
    \new_[58996]_ , \new_[58997]_ , \new_[58998]_ , \new_[59002]_ ,
    \new_[59003]_ , \new_[59007]_ , \new_[59008]_ , \new_[59009]_ ,
    \new_[59013]_ , \new_[59014]_ , \new_[59017]_ , \new_[59020]_ ,
    \new_[59021]_ , \new_[59022]_ , \new_[59026]_ , \new_[59027]_ ,
    \new_[59031]_ , \new_[59032]_ , \new_[59033]_ , \new_[59037]_ ,
    \new_[59038]_ , \new_[59041]_ , \new_[59044]_ , \new_[59045]_ ,
    \new_[59046]_ , \new_[59050]_ , \new_[59051]_ , \new_[59055]_ ,
    \new_[59056]_ , \new_[59057]_ , \new_[59061]_ , \new_[59062]_ ,
    \new_[59065]_ , \new_[59068]_ , \new_[59069]_ , \new_[59070]_ ,
    \new_[59074]_ , \new_[59075]_ , \new_[59079]_ , \new_[59080]_ ,
    \new_[59081]_ , \new_[59085]_ , \new_[59086]_ , \new_[59089]_ ,
    \new_[59092]_ , \new_[59093]_ , \new_[59094]_ , \new_[59098]_ ,
    \new_[59099]_ , \new_[59103]_ , \new_[59104]_ , \new_[59105]_ ,
    \new_[59109]_ , \new_[59110]_ , \new_[59113]_ , \new_[59116]_ ,
    \new_[59117]_ , \new_[59118]_ , \new_[59122]_ , \new_[59123]_ ,
    \new_[59127]_ , \new_[59128]_ , \new_[59129]_ , \new_[59133]_ ,
    \new_[59134]_ , \new_[59137]_ , \new_[59140]_ , \new_[59141]_ ,
    \new_[59142]_ , \new_[59146]_ , \new_[59147]_ , \new_[59151]_ ,
    \new_[59152]_ , \new_[59153]_ , \new_[59157]_ , \new_[59158]_ ,
    \new_[59161]_ , \new_[59164]_ , \new_[59165]_ , \new_[59166]_ ,
    \new_[59170]_ , \new_[59171]_ , \new_[59175]_ , \new_[59176]_ ,
    \new_[59177]_ , \new_[59181]_ , \new_[59182]_ , \new_[59185]_ ,
    \new_[59188]_ , \new_[59189]_ , \new_[59190]_ , \new_[59194]_ ,
    \new_[59195]_ , \new_[59199]_ , \new_[59200]_ , \new_[59201]_ ,
    \new_[59205]_ , \new_[59206]_ , \new_[59209]_ , \new_[59212]_ ,
    \new_[59213]_ , \new_[59214]_ , \new_[59218]_ , \new_[59219]_ ,
    \new_[59223]_ , \new_[59224]_ , \new_[59225]_ , \new_[59229]_ ,
    \new_[59230]_ , \new_[59233]_ , \new_[59236]_ , \new_[59237]_ ,
    \new_[59238]_ , \new_[59242]_ , \new_[59243]_ , \new_[59247]_ ,
    \new_[59248]_ , \new_[59249]_ , \new_[59253]_ , \new_[59254]_ ,
    \new_[59257]_ , \new_[59260]_ , \new_[59261]_ , \new_[59262]_ ,
    \new_[59266]_ , \new_[59267]_ , \new_[59271]_ , \new_[59272]_ ,
    \new_[59273]_ , \new_[59277]_ , \new_[59278]_ , \new_[59281]_ ,
    \new_[59284]_ , \new_[59285]_ , \new_[59286]_ , \new_[59290]_ ,
    \new_[59291]_ , \new_[59295]_ , \new_[59296]_ , \new_[59297]_ ,
    \new_[59301]_ , \new_[59302]_ , \new_[59305]_ , \new_[59308]_ ,
    \new_[59309]_ , \new_[59310]_ , \new_[59314]_ , \new_[59315]_ ,
    \new_[59319]_ , \new_[59320]_ , \new_[59321]_ , \new_[59325]_ ,
    \new_[59326]_ , \new_[59329]_ , \new_[59332]_ , \new_[59333]_ ,
    \new_[59334]_ , \new_[59338]_ , \new_[59339]_ , \new_[59343]_ ,
    \new_[59344]_ , \new_[59345]_ , \new_[59349]_ , \new_[59350]_ ,
    \new_[59353]_ , \new_[59356]_ , \new_[59357]_ , \new_[59358]_ ,
    \new_[59362]_ , \new_[59363]_ , \new_[59367]_ , \new_[59368]_ ,
    \new_[59369]_ , \new_[59373]_ , \new_[59374]_ , \new_[59377]_ ,
    \new_[59380]_ , \new_[59381]_ , \new_[59382]_ , \new_[59386]_ ,
    \new_[59387]_ , \new_[59391]_ , \new_[59392]_ , \new_[59393]_ ,
    \new_[59397]_ , \new_[59398]_ , \new_[59401]_ , \new_[59404]_ ,
    \new_[59405]_ , \new_[59406]_ , \new_[59410]_ , \new_[59411]_ ,
    \new_[59415]_ , \new_[59416]_ , \new_[59417]_ , \new_[59421]_ ,
    \new_[59422]_ , \new_[59425]_ , \new_[59428]_ , \new_[59429]_ ,
    \new_[59430]_ , \new_[59434]_ , \new_[59435]_ , \new_[59439]_ ,
    \new_[59440]_ , \new_[59441]_ , \new_[59445]_ , \new_[59446]_ ,
    \new_[59449]_ , \new_[59452]_ , \new_[59453]_ , \new_[59454]_ ,
    \new_[59458]_ , \new_[59459]_ , \new_[59463]_ , \new_[59464]_ ,
    \new_[59465]_ , \new_[59469]_ , \new_[59470]_ , \new_[59473]_ ,
    \new_[59476]_ , \new_[59477]_ , \new_[59478]_ , \new_[59482]_ ,
    \new_[59483]_ , \new_[59487]_ , \new_[59488]_ , \new_[59489]_ ,
    \new_[59493]_ , \new_[59494]_ , \new_[59497]_ , \new_[59500]_ ,
    \new_[59501]_ , \new_[59502]_ , \new_[59506]_ , \new_[59507]_ ,
    \new_[59511]_ , \new_[59512]_ , \new_[59513]_ , \new_[59517]_ ,
    \new_[59518]_ , \new_[59521]_ , \new_[59524]_ , \new_[59525]_ ,
    \new_[59526]_ , \new_[59530]_ , \new_[59531]_ , \new_[59535]_ ,
    \new_[59536]_ , \new_[59537]_ , \new_[59541]_ , \new_[59542]_ ,
    \new_[59545]_ , \new_[59548]_ , \new_[59549]_ , \new_[59550]_ ,
    \new_[59554]_ , \new_[59555]_ , \new_[59559]_ , \new_[59560]_ ,
    \new_[59561]_ , \new_[59565]_ , \new_[59566]_ , \new_[59569]_ ,
    \new_[59572]_ , \new_[59573]_ , \new_[59574]_ , \new_[59578]_ ,
    \new_[59579]_ , \new_[59583]_ , \new_[59584]_ , \new_[59585]_ ,
    \new_[59589]_ , \new_[59590]_ , \new_[59593]_ , \new_[59596]_ ,
    \new_[59597]_ , \new_[59598]_ , \new_[59602]_ , \new_[59603]_ ,
    \new_[59607]_ , \new_[59608]_ , \new_[59609]_ , \new_[59613]_ ,
    \new_[59614]_ , \new_[59617]_ , \new_[59620]_ , \new_[59621]_ ,
    \new_[59622]_ , \new_[59626]_ , \new_[59627]_ , \new_[59631]_ ,
    \new_[59632]_ , \new_[59633]_ , \new_[59637]_ , \new_[59638]_ ,
    \new_[59641]_ , \new_[59644]_ , \new_[59645]_ , \new_[59646]_ ,
    \new_[59650]_ , \new_[59651]_ , \new_[59655]_ , \new_[59656]_ ,
    \new_[59657]_ , \new_[59661]_ , \new_[59662]_ , \new_[59665]_ ,
    \new_[59668]_ , \new_[59669]_ , \new_[59670]_ , \new_[59674]_ ,
    \new_[59675]_ , \new_[59679]_ , \new_[59680]_ , \new_[59681]_ ,
    \new_[59685]_ , \new_[59686]_ , \new_[59689]_ , \new_[59692]_ ,
    \new_[59693]_ , \new_[59694]_ , \new_[59698]_ , \new_[59699]_ ,
    \new_[59703]_ , \new_[59704]_ , \new_[59705]_ , \new_[59709]_ ,
    \new_[59710]_ , \new_[59713]_ , \new_[59716]_ , \new_[59717]_ ,
    \new_[59718]_ , \new_[59722]_ , \new_[59723]_ , \new_[59727]_ ,
    \new_[59728]_ , \new_[59729]_ , \new_[59733]_ , \new_[59734]_ ,
    \new_[59737]_ , \new_[59740]_ , \new_[59741]_ , \new_[59742]_ ,
    \new_[59746]_ , \new_[59747]_ , \new_[59751]_ , \new_[59752]_ ,
    \new_[59753]_ , \new_[59757]_ , \new_[59758]_ , \new_[59761]_ ,
    \new_[59764]_ , \new_[59765]_ , \new_[59766]_ , \new_[59770]_ ,
    \new_[59771]_ , \new_[59775]_ , \new_[59776]_ , \new_[59777]_ ,
    \new_[59781]_ , \new_[59782]_ , \new_[59785]_ , \new_[59788]_ ,
    \new_[59789]_ , \new_[59790]_ , \new_[59794]_ , \new_[59795]_ ,
    \new_[59799]_ , \new_[59800]_ , \new_[59801]_ , \new_[59805]_ ,
    \new_[59806]_ , \new_[59809]_ , \new_[59812]_ , \new_[59813]_ ,
    \new_[59814]_ , \new_[59818]_ , \new_[59819]_ , \new_[59823]_ ,
    \new_[59824]_ , \new_[59825]_ , \new_[59829]_ , \new_[59830]_ ,
    \new_[59833]_ , \new_[59836]_ , \new_[59837]_ , \new_[59838]_ ,
    \new_[59842]_ , \new_[59843]_ , \new_[59847]_ , \new_[59848]_ ,
    \new_[59849]_ , \new_[59853]_ , \new_[59854]_ , \new_[59857]_ ,
    \new_[59860]_ , \new_[59861]_ , \new_[59862]_ , \new_[59866]_ ,
    \new_[59867]_ , \new_[59871]_ , \new_[59872]_ , \new_[59873]_ ,
    \new_[59877]_ , \new_[59878]_ , \new_[59881]_ , \new_[59884]_ ,
    \new_[59885]_ , \new_[59886]_ , \new_[59890]_ , \new_[59891]_ ,
    \new_[59895]_ , \new_[59896]_ , \new_[59897]_ , \new_[59901]_ ,
    \new_[59902]_ , \new_[59905]_ , \new_[59908]_ , \new_[59909]_ ,
    \new_[59910]_ , \new_[59914]_ , \new_[59915]_ , \new_[59919]_ ,
    \new_[59920]_ , \new_[59921]_ , \new_[59925]_ , \new_[59926]_ ,
    \new_[59929]_ , \new_[59932]_ , \new_[59933]_ , \new_[59934]_ ,
    \new_[59938]_ , \new_[59939]_ , \new_[59943]_ , \new_[59944]_ ,
    \new_[59945]_ , \new_[59949]_ , \new_[59950]_ , \new_[59953]_ ,
    \new_[59956]_ , \new_[59957]_ , \new_[59958]_ , \new_[59962]_ ,
    \new_[59963]_ , \new_[59967]_ , \new_[59968]_ , \new_[59969]_ ,
    \new_[59973]_ , \new_[59974]_ , \new_[59977]_ , \new_[59980]_ ,
    \new_[59981]_ , \new_[59982]_ , \new_[59986]_ , \new_[59987]_ ,
    \new_[59991]_ , \new_[59992]_ , \new_[59993]_ , \new_[59997]_ ,
    \new_[59998]_ , \new_[60001]_ , \new_[60004]_ , \new_[60005]_ ,
    \new_[60006]_ , \new_[60010]_ , \new_[60011]_ , \new_[60015]_ ,
    \new_[60016]_ , \new_[60017]_ , \new_[60021]_ , \new_[60022]_ ,
    \new_[60025]_ , \new_[60028]_ , \new_[60029]_ , \new_[60030]_ ,
    \new_[60034]_ , \new_[60035]_ , \new_[60039]_ , \new_[60040]_ ,
    \new_[60041]_ , \new_[60045]_ , \new_[60046]_ , \new_[60049]_ ,
    \new_[60052]_ , \new_[60053]_ , \new_[60054]_ , \new_[60058]_ ,
    \new_[60059]_ , \new_[60063]_ , \new_[60064]_ , \new_[60065]_ ,
    \new_[60069]_ , \new_[60070]_ , \new_[60073]_ , \new_[60076]_ ,
    \new_[60077]_ , \new_[60078]_ , \new_[60082]_ , \new_[60083]_ ,
    \new_[60087]_ , \new_[60088]_ , \new_[60089]_ , \new_[60093]_ ,
    \new_[60094]_ , \new_[60097]_ , \new_[60100]_ , \new_[60101]_ ,
    \new_[60102]_ , \new_[60106]_ , \new_[60107]_ , \new_[60111]_ ,
    \new_[60112]_ , \new_[60113]_ , \new_[60117]_ , \new_[60118]_ ,
    \new_[60121]_ , \new_[60124]_ , \new_[60125]_ , \new_[60126]_ ,
    \new_[60130]_ , \new_[60131]_ , \new_[60135]_ , \new_[60136]_ ,
    \new_[60137]_ , \new_[60141]_ , \new_[60142]_ , \new_[60145]_ ,
    \new_[60148]_ , \new_[60149]_ , \new_[60150]_ , \new_[60154]_ ,
    \new_[60155]_ , \new_[60159]_ , \new_[60160]_ , \new_[60161]_ ,
    \new_[60165]_ , \new_[60166]_ , \new_[60169]_ , \new_[60172]_ ,
    \new_[60173]_ , \new_[60174]_ , \new_[60178]_ , \new_[60179]_ ,
    \new_[60183]_ , \new_[60184]_ , \new_[60185]_ , \new_[60189]_ ,
    \new_[60190]_ , \new_[60193]_ , \new_[60196]_ , \new_[60197]_ ,
    \new_[60198]_ , \new_[60202]_ , \new_[60203]_ , \new_[60207]_ ,
    \new_[60208]_ , \new_[60209]_ , \new_[60213]_ , \new_[60214]_ ,
    \new_[60217]_ , \new_[60220]_ , \new_[60221]_ , \new_[60222]_ ,
    \new_[60226]_ , \new_[60227]_ , \new_[60231]_ , \new_[60232]_ ,
    \new_[60233]_ , \new_[60237]_ , \new_[60238]_ , \new_[60241]_ ,
    \new_[60244]_ , \new_[60245]_ , \new_[60246]_ , \new_[60250]_ ,
    \new_[60251]_ , \new_[60255]_ , \new_[60256]_ , \new_[60257]_ ,
    \new_[60261]_ , \new_[60262]_ , \new_[60265]_ , \new_[60268]_ ,
    \new_[60269]_ , \new_[60270]_ , \new_[60274]_ , \new_[60275]_ ,
    \new_[60279]_ , \new_[60280]_ , \new_[60281]_ , \new_[60285]_ ,
    \new_[60286]_ , \new_[60289]_ , \new_[60292]_ , \new_[60293]_ ,
    \new_[60294]_ , \new_[60298]_ , \new_[60299]_ , \new_[60303]_ ,
    \new_[60304]_ , \new_[60305]_ , \new_[60309]_ , \new_[60310]_ ,
    \new_[60313]_ , \new_[60316]_ , \new_[60317]_ , \new_[60318]_ ,
    \new_[60322]_ , \new_[60323]_ , \new_[60327]_ , \new_[60328]_ ,
    \new_[60329]_ , \new_[60333]_ , \new_[60334]_ , \new_[60337]_ ,
    \new_[60340]_ , \new_[60341]_ , \new_[60342]_ , \new_[60346]_ ,
    \new_[60347]_ , \new_[60351]_ , \new_[60352]_ , \new_[60353]_ ,
    \new_[60357]_ , \new_[60358]_ , \new_[60361]_ , \new_[60364]_ ,
    \new_[60365]_ , \new_[60366]_ , \new_[60370]_ , \new_[60371]_ ,
    \new_[60375]_ , \new_[60376]_ , \new_[60377]_ , \new_[60381]_ ,
    \new_[60382]_ , \new_[60385]_ , \new_[60388]_ , \new_[60389]_ ,
    \new_[60390]_ , \new_[60394]_ , \new_[60395]_ , \new_[60399]_ ,
    \new_[60400]_ , \new_[60401]_ , \new_[60405]_ , \new_[60406]_ ,
    \new_[60409]_ , \new_[60412]_ , \new_[60413]_ , \new_[60414]_ ,
    \new_[60418]_ , \new_[60419]_ , \new_[60423]_ , \new_[60424]_ ,
    \new_[60425]_ , \new_[60429]_ , \new_[60430]_ , \new_[60433]_ ,
    \new_[60436]_ , \new_[60437]_ , \new_[60438]_ , \new_[60442]_ ,
    \new_[60443]_ , \new_[60447]_ , \new_[60448]_ , \new_[60449]_ ,
    \new_[60453]_ , \new_[60454]_ , \new_[60457]_ , \new_[60460]_ ,
    \new_[60461]_ , \new_[60462]_ , \new_[60466]_ , \new_[60467]_ ,
    \new_[60471]_ , \new_[60472]_ , \new_[60473]_ , \new_[60477]_ ,
    \new_[60478]_ , \new_[60481]_ , \new_[60484]_ , \new_[60485]_ ,
    \new_[60486]_ , \new_[60490]_ , \new_[60491]_ , \new_[60495]_ ,
    \new_[60496]_ , \new_[60497]_ , \new_[60501]_ , \new_[60502]_ ,
    \new_[60505]_ , \new_[60508]_ , \new_[60509]_ , \new_[60510]_ ,
    \new_[60514]_ , \new_[60515]_ , \new_[60519]_ , \new_[60520]_ ,
    \new_[60521]_ , \new_[60525]_ , \new_[60526]_ , \new_[60529]_ ,
    \new_[60532]_ , \new_[60533]_ , \new_[60534]_ , \new_[60538]_ ,
    \new_[60539]_ , \new_[60543]_ , \new_[60544]_ , \new_[60545]_ ,
    \new_[60549]_ , \new_[60550]_ , \new_[60553]_ , \new_[60556]_ ,
    \new_[60557]_ , \new_[60558]_ , \new_[60562]_ , \new_[60563]_ ,
    \new_[60567]_ , \new_[60568]_ , \new_[60569]_ , \new_[60573]_ ,
    \new_[60574]_ , \new_[60577]_ , \new_[60580]_ , \new_[60581]_ ,
    \new_[60582]_ , \new_[60586]_ , \new_[60587]_ , \new_[60591]_ ,
    \new_[60592]_ , \new_[60593]_ , \new_[60597]_ , \new_[60598]_ ,
    \new_[60601]_ , \new_[60604]_ , \new_[60605]_ , \new_[60606]_ ,
    \new_[60610]_ , \new_[60611]_ , \new_[60615]_ , \new_[60616]_ ,
    \new_[60617]_ , \new_[60621]_ , \new_[60622]_ , \new_[60625]_ ,
    \new_[60628]_ , \new_[60629]_ , \new_[60630]_ , \new_[60634]_ ,
    \new_[60635]_ , \new_[60639]_ , \new_[60640]_ , \new_[60641]_ ,
    \new_[60645]_ , \new_[60646]_ , \new_[60649]_ , \new_[60652]_ ,
    \new_[60653]_ , \new_[60654]_ , \new_[60658]_ , \new_[60659]_ ,
    \new_[60663]_ , \new_[60664]_ , \new_[60665]_ , \new_[60669]_ ,
    \new_[60670]_ , \new_[60673]_ , \new_[60676]_ , \new_[60677]_ ,
    \new_[60678]_ , \new_[60682]_ , \new_[60683]_ , \new_[60687]_ ,
    \new_[60688]_ , \new_[60689]_ , \new_[60693]_ , \new_[60694]_ ,
    \new_[60697]_ , \new_[60700]_ , \new_[60701]_ , \new_[60702]_ ,
    \new_[60706]_ , \new_[60707]_ , \new_[60711]_ , \new_[60712]_ ,
    \new_[60713]_ , \new_[60717]_ , \new_[60718]_ , \new_[60721]_ ,
    \new_[60724]_ , \new_[60725]_ , \new_[60726]_ , \new_[60730]_ ,
    \new_[60731]_ , \new_[60735]_ , \new_[60736]_ , \new_[60737]_ ,
    \new_[60741]_ , \new_[60742]_ , \new_[60745]_ , \new_[60748]_ ,
    \new_[60749]_ , \new_[60750]_ , \new_[60754]_ , \new_[60755]_ ,
    \new_[60759]_ , \new_[60760]_ , \new_[60761]_ , \new_[60765]_ ,
    \new_[60766]_ , \new_[60769]_ , \new_[60772]_ , \new_[60773]_ ,
    \new_[60774]_ , \new_[60778]_ , \new_[60779]_ , \new_[60783]_ ,
    \new_[60784]_ , \new_[60785]_ , \new_[60789]_ , \new_[60790]_ ,
    \new_[60793]_ , \new_[60796]_ , \new_[60797]_ , \new_[60798]_ ,
    \new_[60802]_ , \new_[60803]_ , \new_[60807]_ , \new_[60808]_ ,
    \new_[60809]_ , \new_[60813]_ , \new_[60814]_ , \new_[60817]_ ,
    \new_[60820]_ , \new_[60821]_ , \new_[60822]_ , \new_[60826]_ ,
    \new_[60827]_ , \new_[60831]_ , \new_[60832]_ , \new_[60833]_ ,
    \new_[60837]_ , \new_[60838]_ , \new_[60841]_ , \new_[60844]_ ,
    \new_[60845]_ , \new_[60846]_ , \new_[60850]_ , \new_[60851]_ ,
    \new_[60855]_ , \new_[60856]_ , \new_[60857]_ , \new_[60861]_ ,
    \new_[60862]_ , \new_[60865]_ , \new_[60868]_ , \new_[60869]_ ,
    \new_[60870]_ , \new_[60874]_ , \new_[60875]_ , \new_[60879]_ ,
    \new_[60880]_ , \new_[60881]_ , \new_[60885]_ , \new_[60886]_ ,
    \new_[60889]_ , \new_[60892]_ , \new_[60893]_ , \new_[60894]_ ,
    \new_[60898]_ , \new_[60899]_ , \new_[60903]_ , \new_[60904]_ ,
    \new_[60905]_ , \new_[60909]_ , \new_[60910]_ , \new_[60913]_ ,
    \new_[60916]_ , \new_[60917]_ , \new_[60918]_ , \new_[60922]_ ,
    \new_[60923]_ , \new_[60927]_ , \new_[60928]_ , \new_[60929]_ ,
    \new_[60933]_ , \new_[60934]_ , \new_[60937]_ , \new_[60940]_ ,
    \new_[60941]_ , \new_[60942]_ , \new_[60946]_ , \new_[60947]_ ,
    \new_[60951]_ , \new_[60952]_ , \new_[60953]_ , \new_[60957]_ ,
    \new_[60958]_ , \new_[60961]_ , \new_[60964]_ , \new_[60965]_ ,
    \new_[60966]_ , \new_[60970]_ , \new_[60971]_ , \new_[60975]_ ,
    \new_[60976]_ , \new_[60977]_ , \new_[60981]_ , \new_[60982]_ ,
    \new_[60985]_ , \new_[60988]_ , \new_[60989]_ , \new_[60990]_ ,
    \new_[60994]_ , \new_[60995]_ , \new_[60999]_ , \new_[61000]_ ,
    \new_[61001]_ , \new_[61005]_ , \new_[61006]_ , \new_[61009]_ ,
    \new_[61012]_ , \new_[61013]_ , \new_[61014]_ , \new_[61018]_ ,
    \new_[61019]_ , \new_[61023]_ , \new_[61024]_ , \new_[61025]_ ,
    \new_[61029]_ , \new_[61030]_ , \new_[61033]_ , \new_[61036]_ ,
    \new_[61037]_ , \new_[61038]_ , \new_[61042]_ , \new_[61043]_ ,
    \new_[61047]_ , \new_[61048]_ , \new_[61049]_ , \new_[61053]_ ,
    \new_[61054]_ , \new_[61057]_ , \new_[61060]_ , \new_[61061]_ ,
    \new_[61062]_ , \new_[61066]_ , \new_[61067]_ , \new_[61071]_ ,
    \new_[61072]_ , \new_[61073]_ , \new_[61077]_ , \new_[61078]_ ,
    \new_[61081]_ , \new_[61084]_ , \new_[61085]_ , \new_[61086]_ ,
    \new_[61090]_ , \new_[61091]_ , \new_[61095]_ , \new_[61096]_ ,
    \new_[61097]_ , \new_[61101]_ , \new_[61102]_ , \new_[61105]_ ,
    \new_[61108]_ , \new_[61109]_ , \new_[61110]_ , \new_[61114]_ ,
    \new_[61115]_ , \new_[61119]_ , \new_[61120]_ , \new_[61121]_ ,
    \new_[61125]_ , \new_[61126]_ , \new_[61129]_ , \new_[61132]_ ,
    \new_[61133]_ , \new_[61134]_ , \new_[61138]_ , \new_[61139]_ ,
    \new_[61143]_ , \new_[61144]_ , \new_[61145]_ , \new_[61149]_ ,
    \new_[61150]_ , \new_[61153]_ , \new_[61156]_ , \new_[61157]_ ,
    \new_[61158]_ , \new_[61162]_ , \new_[61163]_ , \new_[61167]_ ,
    \new_[61168]_ , \new_[61169]_ , \new_[61173]_ , \new_[61174]_ ,
    \new_[61177]_ , \new_[61180]_ , \new_[61181]_ , \new_[61182]_ ,
    \new_[61186]_ , \new_[61187]_ , \new_[61191]_ , \new_[61192]_ ,
    \new_[61193]_ , \new_[61197]_ , \new_[61198]_ , \new_[61201]_ ,
    \new_[61204]_ , \new_[61205]_ , \new_[61206]_ , \new_[61210]_ ,
    \new_[61211]_ , \new_[61215]_ , \new_[61216]_ , \new_[61217]_ ,
    \new_[61221]_ , \new_[61222]_ , \new_[61225]_ , \new_[61228]_ ,
    \new_[61229]_ , \new_[61230]_ , \new_[61234]_ , \new_[61235]_ ,
    \new_[61239]_ , \new_[61240]_ , \new_[61241]_ , \new_[61245]_ ,
    \new_[61246]_ , \new_[61249]_ , \new_[61252]_ , \new_[61253]_ ,
    \new_[61254]_ , \new_[61258]_ , \new_[61259]_ , \new_[61263]_ ,
    \new_[61264]_ , \new_[61265]_ , \new_[61269]_ , \new_[61270]_ ,
    \new_[61273]_ , \new_[61276]_ , \new_[61277]_ , \new_[61278]_ ,
    \new_[61282]_ , \new_[61283]_ , \new_[61287]_ , \new_[61288]_ ,
    \new_[61289]_ , \new_[61293]_ , \new_[61294]_ , \new_[61297]_ ,
    \new_[61300]_ , \new_[61301]_ , \new_[61302]_ , \new_[61306]_ ,
    \new_[61307]_ , \new_[61311]_ , \new_[61312]_ , \new_[61313]_ ,
    \new_[61317]_ , \new_[61318]_ , \new_[61321]_ , \new_[61324]_ ,
    \new_[61325]_ , \new_[61326]_ , \new_[61330]_ , \new_[61331]_ ,
    \new_[61335]_ , \new_[61336]_ , \new_[61337]_ , \new_[61341]_ ,
    \new_[61342]_ , \new_[61345]_ , \new_[61348]_ , \new_[61349]_ ,
    \new_[61350]_ , \new_[61354]_ , \new_[61355]_ , \new_[61359]_ ,
    \new_[61360]_ , \new_[61361]_ , \new_[61365]_ , \new_[61366]_ ,
    \new_[61369]_ , \new_[61372]_ , \new_[61373]_ , \new_[61374]_ ,
    \new_[61378]_ , \new_[61379]_ , \new_[61383]_ , \new_[61384]_ ,
    \new_[61385]_ , \new_[61389]_ , \new_[61390]_ , \new_[61393]_ ,
    \new_[61396]_ , \new_[61397]_ , \new_[61398]_ , \new_[61402]_ ,
    \new_[61403]_ , \new_[61407]_ , \new_[61408]_ , \new_[61409]_ ,
    \new_[61413]_ , \new_[61414]_ , \new_[61417]_ , \new_[61420]_ ,
    \new_[61421]_ , \new_[61422]_ , \new_[61426]_ , \new_[61427]_ ,
    \new_[61431]_ , \new_[61432]_ , \new_[61433]_ , \new_[61437]_ ,
    \new_[61438]_ , \new_[61441]_ , \new_[61444]_ , \new_[61445]_ ,
    \new_[61446]_ , \new_[61450]_ , \new_[61451]_ , \new_[61455]_ ,
    \new_[61456]_ , \new_[61457]_ , \new_[61461]_ , \new_[61462]_ ,
    \new_[61465]_ , \new_[61468]_ , \new_[61469]_ , \new_[61470]_ ,
    \new_[61474]_ , \new_[61475]_ , \new_[61479]_ , \new_[61480]_ ,
    \new_[61481]_ , \new_[61485]_ , \new_[61486]_ , \new_[61489]_ ,
    \new_[61492]_ , \new_[61493]_ , \new_[61494]_ , \new_[61498]_ ,
    \new_[61499]_ , \new_[61503]_ , \new_[61504]_ , \new_[61505]_ ,
    \new_[61509]_ , \new_[61510]_ , \new_[61513]_ , \new_[61516]_ ,
    \new_[61517]_ , \new_[61518]_ , \new_[61522]_ , \new_[61523]_ ,
    \new_[61527]_ , \new_[61528]_ , \new_[61529]_ , \new_[61533]_ ,
    \new_[61534]_ , \new_[61537]_ , \new_[61540]_ , \new_[61541]_ ,
    \new_[61542]_ , \new_[61546]_ , \new_[61547]_ , \new_[61551]_ ,
    \new_[61552]_ , \new_[61553]_ , \new_[61557]_ , \new_[61558]_ ,
    \new_[61561]_ , \new_[61564]_ , \new_[61565]_ , \new_[61566]_ ,
    \new_[61570]_ , \new_[61571]_ , \new_[61575]_ , \new_[61576]_ ,
    \new_[61577]_ , \new_[61581]_ , \new_[61582]_ , \new_[61585]_ ,
    \new_[61588]_ , \new_[61589]_ , \new_[61590]_ , \new_[61594]_ ,
    \new_[61595]_ , \new_[61599]_ , \new_[61600]_ , \new_[61601]_ ,
    \new_[61605]_ , \new_[61606]_ , \new_[61609]_ , \new_[61612]_ ,
    \new_[61613]_ , \new_[61614]_ , \new_[61618]_ , \new_[61619]_ ,
    \new_[61623]_ , \new_[61624]_ , \new_[61625]_ , \new_[61629]_ ,
    \new_[61630]_ , \new_[61633]_ , \new_[61636]_ , \new_[61637]_ ,
    \new_[61638]_ , \new_[61642]_ , \new_[61643]_ , \new_[61647]_ ,
    \new_[61648]_ , \new_[61649]_ , \new_[61653]_ , \new_[61654]_ ,
    \new_[61657]_ , \new_[61660]_ , \new_[61661]_ , \new_[61662]_ ,
    \new_[61666]_ , \new_[61667]_ , \new_[61671]_ , \new_[61672]_ ,
    \new_[61673]_ , \new_[61677]_ , \new_[61678]_ , \new_[61681]_ ,
    \new_[61684]_ , \new_[61685]_ , \new_[61686]_ , \new_[61690]_ ,
    \new_[61691]_ , \new_[61695]_ , \new_[61696]_ , \new_[61697]_ ,
    \new_[61701]_ , \new_[61702]_ , \new_[61705]_ , \new_[61708]_ ,
    \new_[61709]_ , \new_[61710]_ , \new_[61714]_ , \new_[61715]_ ,
    \new_[61719]_ , \new_[61720]_ , \new_[61721]_ , \new_[61725]_ ,
    \new_[61726]_ , \new_[61729]_ , \new_[61732]_ , \new_[61733]_ ,
    \new_[61734]_ , \new_[61738]_ , \new_[61739]_ , \new_[61743]_ ,
    \new_[61744]_ , \new_[61745]_ , \new_[61749]_ , \new_[61750]_ ,
    \new_[61753]_ , \new_[61756]_ , \new_[61757]_ , \new_[61758]_ ,
    \new_[61762]_ , \new_[61763]_ , \new_[61767]_ , \new_[61768]_ ,
    \new_[61769]_ , \new_[61773]_ , \new_[61774]_ , \new_[61777]_ ,
    \new_[61780]_ , \new_[61781]_ , \new_[61782]_ , \new_[61786]_ ,
    \new_[61787]_ , \new_[61791]_ , \new_[61792]_ , \new_[61793]_ ,
    \new_[61797]_ , \new_[61798]_ , \new_[61801]_ , \new_[61804]_ ,
    \new_[61805]_ , \new_[61806]_ , \new_[61810]_ , \new_[61811]_ ,
    \new_[61815]_ , \new_[61816]_ , \new_[61817]_ , \new_[61821]_ ,
    \new_[61822]_ , \new_[61825]_ , \new_[61828]_ , \new_[61829]_ ,
    \new_[61830]_ , \new_[61834]_ , \new_[61835]_ , \new_[61839]_ ,
    \new_[61840]_ , \new_[61841]_ , \new_[61845]_ , \new_[61846]_ ,
    \new_[61849]_ , \new_[61852]_ , \new_[61853]_ , \new_[61854]_ ,
    \new_[61858]_ , \new_[61859]_ , \new_[61863]_ , \new_[61864]_ ,
    \new_[61865]_ , \new_[61869]_ , \new_[61870]_ , \new_[61873]_ ,
    \new_[61876]_ , \new_[61877]_ , \new_[61878]_ , \new_[61882]_ ,
    \new_[61883]_ , \new_[61887]_ , \new_[61888]_ , \new_[61889]_ ,
    \new_[61893]_ , \new_[61894]_ , \new_[61897]_ , \new_[61900]_ ,
    \new_[61901]_ , \new_[61902]_ , \new_[61906]_ , \new_[61907]_ ,
    \new_[61911]_ , \new_[61912]_ , \new_[61913]_ , \new_[61917]_ ,
    \new_[61918]_ , \new_[61921]_ , \new_[61924]_ , \new_[61925]_ ,
    \new_[61926]_ , \new_[61930]_ , \new_[61931]_ , \new_[61935]_ ,
    \new_[61936]_ , \new_[61937]_ , \new_[61941]_ , \new_[61942]_ ,
    \new_[61945]_ , \new_[61948]_ , \new_[61949]_ , \new_[61950]_ ,
    \new_[61954]_ , \new_[61955]_ , \new_[61959]_ , \new_[61960]_ ,
    \new_[61961]_ , \new_[61965]_ , \new_[61966]_ , \new_[61969]_ ,
    \new_[61972]_ , \new_[61973]_ , \new_[61974]_ , \new_[61978]_ ,
    \new_[61979]_ , \new_[61983]_ , \new_[61984]_ , \new_[61985]_ ,
    \new_[61989]_ , \new_[61990]_ , \new_[61993]_ , \new_[61996]_ ,
    \new_[61997]_ , \new_[61998]_ , \new_[62002]_ , \new_[62003]_ ,
    \new_[62007]_ , \new_[62008]_ , \new_[62009]_ , \new_[62013]_ ,
    \new_[62014]_ , \new_[62017]_ , \new_[62020]_ , \new_[62021]_ ,
    \new_[62022]_ , \new_[62026]_ , \new_[62027]_ , \new_[62031]_ ,
    \new_[62032]_ , \new_[62033]_ , \new_[62037]_ , \new_[62038]_ ,
    \new_[62041]_ , \new_[62044]_ , \new_[62045]_ , \new_[62046]_ ,
    \new_[62050]_ , \new_[62051]_ , \new_[62055]_ , \new_[62056]_ ,
    \new_[62057]_ , \new_[62061]_ , \new_[62062]_ , \new_[62065]_ ,
    \new_[62068]_ , \new_[62069]_ , \new_[62070]_ , \new_[62074]_ ,
    \new_[62075]_ , \new_[62079]_ , \new_[62080]_ , \new_[62081]_ ,
    \new_[62085]_ , \new_[62086]_ , \new_[62089]_ , \new_[62092]_ ,
    \new_[62093]_ , \new_[62094]_ , \new_[62098]_ , \new_[62099]_ ,
    \new_[62103]_ , \new_[62104]_ , \new_[62105]_ , \new_[62109]_ ,
    \new_[62110]_ , \new_[62113]_ , \new_[62116]_ , \new_[62117]_ ,
    \new_[62118]_ , \new_[62122]_ , \new_[62123]_ , \new_[62127]_ ,
    \new_[62128]_ , \new_[62129]_ , \new_[62133]_ , \new_[62134]_ ,
    \new_[62137]_ , \new_[62140]_ , \new_[62141]_ , \new_[62142]_ ,
    \new_[62146]_ , \new_[62147]_ , \new_[62151]_ , \new_[62152]_ ,
    \new_[62153]_ , \new_[62157]_ , \new_[62158]_ , \new_[62161]_ ,
    \new_[62164]_ , \new_[62165]_ , \new_[62166]_ , \new_[62170]_ ,
    \new_[62171]_ , \new_[62175]_ , \new_[62176]_ , \new_[62177]_ ,
    \new_[62181]_ , \new_[62182]_ , \new_[62185]_ , \new_[62188]_ ,
    \new_[62189]_ , \new_[62190]_ , \new_[62194]_ , \new_[62195]_ ,
    \new_[62199]_ , \new_[62200]_ , \new_[62201]_ , \new_[62205]_ ,
    \new_[62206]_ , \new_[62209]_ , \new_[62212]_ , \new_[62213]_ ,
    \new_[62214]_ , \new_[62218]_ , \new_[62219]_ , \new_[62223]_ ,
    \new_[62224]_ , \new_[62225]_ , \new_[62229]_ , \new_[62230]_ ,
    \new_[62233]_ , \new_[62236]_ , \new_[62237]_ , \new_[62238]_ ,
    \new_[62242]_ , \new_[62243]_ , \new_[62247]_ , \new_[62248]_ ,
    \new_[62249]_ , \new_[62253]_ , \new_[62254]_ , \new_[62257]_ ,
    \new_[62260]_ , \new_[62261]_ , \new_[62262]_ , \new_[62266]_ ,
    \new_[62267]_ , \new_[62271]_ , \new_[62272]_ , \new_[62273]_ ,
    \new_[62277]_ , \new_[62278]_ , \new_[62281]_ , \new_[62284]_ ,
    \new_[62285]_ , \new_[62286]_ , \new_[62290]_ , \new_[62291]_ ,
    \new_[62295]_ , \new_[62296]_ , \new_[62297]_ , \new_[62301]_ ,
    \new_[62302]_ , \new_[62305]_ , \new_[62308]_ , \new_[62309]_ ,
    \new_[62310]_ , \new_[62314]_ , \new_[62315]_ , \new_[62319]_ ,
    \new_[62320]_ , \new_[62321]_ , \new_[62325]_ , \new_[62326]_ ,
    \new_[62329]_ , \new_[62332]_ , \new_[62333]_ , \new_[62334]_ ,
    \new_[62338]_ , \new_[62339]_ , \new_[62343]_ , \new_[62344]_ ,
    \new_[62345]_ , \new_[62349]_ , \new_[62350]_ , \new_[62353]_ ,
    \new_[62356]_ , \new_[62357]_ , \new_[62358]_ , \new_[62362]_ ,
    \new_[62363]_ , \new_[62367]_ , \new_[62368]_ , \new_[62369]_ ,
    \new_[62373]_ , \new_[62374]_ , \new_[62377]_ , \new_[62380]_ ,
    \new_[62381]_ , \new_[62382]_ , \new_[62386]_ , \new_[62387]_ ,
    \new_[62391]_ , \new_[62392]_ , \new_[62393]_ , \new_[62397]_ ,
    \new_[62398]_ , \new_[62401]_ , \new_[62404]_ , \new_[62405]_ ,
    \new_[62406]_ , \new_[62410]_ , \new_[62411]_ , \new_[62415]_ ,
    \new_[62416]_ , \new_[62417]_ , \new_[62421]_ , \new_[62422]_ ,
    \new_[62425]_ , \new_[62428]_ , \new_[62429]_ , \new_[62430]_ ,
    \new_[62434]_ , \new_[62435]_ , \new_[62439]_ , \new_[62440]_ ,
    \new_[62441]_ , \new_[62445]_ , \new_[62446]_ , \new_[62449]_ ,
    \new_[62452]_ , \new_[62453]_ , \new_[62454]_ , \new_[62458]_ ,
    \new_[62459]_ , \new_[62463]_ , \new_[62464]_ , \new_[62465]_ ,
    \new_[62469]_ , \new_[62470]_ , \new_[62473]_ , \new_[62476]_ ,
    \new_[62477]_ , \new_[62478]_ , \new_[62482]_ , \new_[62483]_ ,
    \new_[62487]_ , \new_[62488]_ , \new_[62489]_ , \new_[62493]_ ,
    \new_[62494]_ , \new_[62497]_ , \new_[62500]_ , \new_[62501]_ ,
    \new_[62502]_ , \new_[62506]_ , \new_[62507]_ , \new_[62511]_ ,
    \new_[62512]_ , \new_[62513]_ , \new_[62517]_ , \new_[62518]_ ,
    \new_[62521]_ , \new_[62524]_ , \new_[62525]_ , \new_[62526]_ ,
    \new_[62530]_ , \new_[62531]_ , \new_[62535]_ , \new_[62536]_ ,
    \new_[62537]_ , \new_[62541]_ , \new_[62542]_ , \new_[62545]_ ,
    \new_[62548]_ , \new_[62549]_ , \new_[62550]_ , \new_[62554]_ ,
    \new_[62555]_ , \new_[62559]_ , \new_[62560]_ , \new_[62561]_ ,
    \new_[62565]_ , \new_[62566]_ , \new_[62569]_ , \new_[62572]_ ,
    \new_[62573]_ , \new_[62574]_ , \new_[62578]_ , \new_[62579]_ ,
    \new_[62583]_ , \new_[62584]_ , \new_[62585]_ , \new_[62589]_ ,
    \new_[62590]_ , \new_[62593]_ , \new_[62596]_ , \new_[62597]_ ,
    \new_[62598]_ , \new_[62602]_ , \new_[62603]_ , \new_[62607]_ ,
    \new_[62608]_ , \new_[62609]_ , \new_[62613]_ , \new_[62614]_ ,
    \new_[62617]_ , \new_[62620]_ , \new_[62621]_ , \new_[62622]_ ,
    \new_[62626]_ , \new_[62627]_ , \new_[62631]_ , \new_[62632]_ ,
    \new_[62633]_ , \new_[62637]_ , \new_[62638]_ , \new_[62641]_ ,
    \new_[62644]_ , \new_[62645]_ , \new_[62646]_ , \new_[62650]_ ,
    \new_[62651]_ , \new_[62655]_ , \new_[62656]_ , \new_[62657]_ ,
    \new_[62661]_ , \new_[62662]_ , \new_[62665]_ , \new_[62668]_ ,
    \new_[62669]_ , \new_[62670]_ , \new_[62674]_ , \new_[62675]_ ,
    \new_[62679]_ , \new_[62680]_ , \new_[62681]_ , \new_[62685]_ ,
    \new_[62686]_ , \new_[62689]_ , \new_[62692]_ , \new_[62693]_ ,
    \new_[62694]_ , \new_[62698]_ , \new_[62699]_ , \new_[62703]_ ,
    \new_[62704]_ , \new_[62705]_ , \new_[62709]_ , \new_[62710]_ ,
    \new_[62713]_ , \new_[62716]_ , \new_[62717]_ , \new_[62718]_ ,
    \new_[62722]_ , \new_[62723]_ , \new_[62727]_ , \new_[62728]_ ,
    \new_[62729]_ , \new_[62733]_ , \new_[62734]_ , \new_[62737]_ ,
    \new_[62740]_ , \new_[62741]_ , \new_[62742]_ , \new_[62746]_ ,
    \new_[62747]_ , \new_[62751]_ , \new_[62752]_ , \new_[62753]_ ,
    \new_[62757]_ , \new_[62758]_ , \new_[62761]_ , \new_[62764]_ ,
    \new_[62765]_ , \new_[62766]_ , \new_[62770]_ , \new_[62771]_ ,
    \new_[62775]_ , \new_[62776]_ , \new_[62777]_ , \new_[62781]_ ,
    \new_[62782]_ , \new_[62785]_ , \new_[62788]_ , \new_[62789]_ ,
    \new_[62790]_ , \new_[62794]_ , \new_[62795]_ , \new_[62799]_ ,
    \new_[62800]_ , \new_[62801]_ , \new_[62805]_ , \new_[62806]_ ,
    \new_[62809]_ , \new_[62812]_ , \new_[62813]_ , \new_[62814]_ ,
    \new_[62818]_ , \new_[62819]_ , \new_[62823]_ , \new_[62824]_ ,
    \new_[62825]_ , \new_[62829]_ , \new_[62830]_ , \new_[62833]_ ,
    \new_[62836]_ , \new_[62837]_ , \new_[62838]_ , \new_[62842]_ ,
    \new_[62843]_ , \new_[62847]_ , \new_[62848]_ , \new_[62849]_ ,
    \new_[62853]_ , \new_[62854]_ , \new_[62857]_ , \new_[62860]_ ,
    \new_[62861]_ , \new_[62862]_ , \new_[62866]_ , \new_[62867]_ ,
    \new_[62871]_ , \new_[62872]_ , \new_[62873]_ , \new_[62877]_ ,
    \new_[62878]_ , \new_[62881]_ , \new_[62884]_ , \new_[62885]_ ,
    \new_[62886]_ , \new_[62890]_ , \new_[62891]_ , \new_[62895]_ ,
    \new_[62896]_ , \new_[62897]_ , \new_[62901]_ , \new_[62902]_ ,
    \new_[62905]_ , \new_[62908]_ , \new_[62909]_ , \new_[62910]_ ,
    \new_[62914]_ , \new_[62915]_ , \new_[62919]_ , \new_[62920]_ ,
    \new_[62921]_ , \new_[62925]_ , \new_[62926]_ , \new_[62929]_ ,
    \new_[62932]_ , \new_[62933]_ , \new_[62934]_ , \new_[62938]_ ,
    \new_[62939]_ , \new_[62943]_ , \new_[62944]_ , \new_[62945]_ ,
    \new_[62949]_ , \new_[62950]_ , \new_[62953]_ , \new_[62956]_ ,
    \new_[62957]_ , \new_[62958]_ , \new_[62962]_ , \new_[62963]_ ,
    \new_[62967]_ , \new_[62968]_ , \new_[62969]_ , \new_[62973]_ ,
    \new_[62974]_ , \new_[62977]_ , \new_[62980]_ , \new_[62981]_ ,
    \new_[62982]_ , \new_[62986]_ , \new_[62987]_ , \new_[62991]_ ,
    \new_[62992]_ , \new_[62993]_ , \new_[62997]_ , \new_[62998]_ ,
    \new_[63001]_ , \new_[63004]_ , \new_[63005]_ , \new_[63006]_ ,
    \new_[63010]_ , \new_[63011]_ , \new_[63015]_ , \new_[63016]_ ,
    \new_[63017]_ , \new_[63021]_ , \new_[63022]_ , \new_[63025]_ ,
    \new_[63028]_ , \new_[63029]_ , \new_[63030]_ , \new_[63034]_ ,
    \new_[63035]_ , \new_[63039]_ , \new_[63040]_ , \new_[63041]_ ,
    \new_[63045]_ , \new_[63046]_ , \new_[63049]_ , \new_[63052]_ ,
    \new_[63053]_ , \new_[63054]_ , \new_[63058]_ , \new_[63059]_ ,
    \new_[63063]_ , \new_[63064]_ , \new_[63065]_ , \new_[63069]_ ,
    \new_[63070]_ , \new_[63073]_ , \new_[63076]_ , \new_[63077]_ ,
    \new_[63078]_ , \new_[63082]_ , \new_[63083]_ , \new_[63087]_ ,
    \new_[63088]_ , \new_[63089]_ , \new_[63093]_ , \new_[63094]_ ,
    \new_[63097]_ , \new_[63100]_ , \new_[63101]_ , \new_[63102]_ ,
    \new_[63106]_ , \new_[63107]_ , \new_[63111]_ , \new_[63112]_ ,
    \new_[63113]_ , \new_[63117]_ , \new_[63118]_ , \new_[63121]_ ,
    \new_[63124]_ , \new_[63125]_ , \new_[63126]_ , \new_[63130]_ ,
    \new_[63131]_ , \new_[63135]_ , \new_[63136]_ , \new_[63137]_ ,
    \new_[63141]_ , \new_[63142]_ , \new_[63145]_ , \new_[63148]_ ,
    \new_[63149]_ , \new_[63150]_ , \new_[63154]_ , \new_[63155]_ ,
    \new_[63159]_ , \new_[63160]_ , \new_[63161]_ , \new_[63165]_ ,
    \new_[63166]_ , \new_[63169]_ , \new_[63172]_ , \new_[63173]_ ,
    \new_[63174]_ , \new_[63178]_ , \new_[63179]_ , \new_[63183]_ ,
    \new_[63184]_ , \new_[63185]_ , \new_[63189]_ , \new_[63190]_ ,
    \new_[63193]_ , \new_[63196]_ , \new_[63197]_ , \new_[63198]_ ,
    \new_[63202]_ , \new_[63203]_ , \new_[63207]_ , \new_[63208]_ ,
    \new_[63209]_ , \new_[63213]_ , \new_[63214]_ , \new_[63217]_ ,
    \new_[63220]_ , \new_[63221]_ , \new_[63222]_ , \new_[63226]_ ,
    \new_[63227]_ , \new_[63231]_ , \new_[63232]_ , \new_[63233]_ ,
    \new_[63237]_ , \new_[63238]_ , \new_[63241]_ , \new_[63244]_ ,
    \new_[63245]_ , \new_[63246]_ , \new_[63250]_ , \new_[63251]_ ,
    \new_[63255]_ , \new_[63256]_ , \new_[63257]_ , \new_[63261]_ ,
    \new_[63262]_ , \new_[63265]_ , \new_[63268]_ , \new_[63269]_ ,
    \new_[63270]_ , \new_[63274]_ , \new_[63275]_ , \new_[63279]_ ,
    \new_[63280]_ , \new_[63281]_ , \new_[63285]_ , \new_[63286]_ ,
    \new_[63289]_ , \new_[63292]_ , \new_[63293]_ , \new_[63294]_ ,
    \new_[63298]_ , \new_[63299]_ , \new_[63303]_ , \new_[63304]_ ,
    \new_[63305]_ , \new_[63309]_ , \new_[63310]_ , \new_[63313]_ ,
    \new_[63316]_ , \new_[63317]_ , \new_[63318]_ , \new_[63322]_ ,
    \new_[63323]_ , \new_[63327]_ , \new_[63328]_ , \new_[63329]_ ,
    \new_[63333]_ , \new_[63334]_ , \new_[63337]_ , \new_[63340]_ ,
    \new_[63341]_ , \new_[63342]_ , \new_[63346]_ , \new_[63347]_ ,
    \new_[63351]_ , \new_[63352]_ , \new_[63353]_ , \new_[63357]_ ,
    \new_[63358]_ , \new_[63361]_ , \new_[63364]_ , \new_[63365]_ ,
    \new_[63366]_ , \new_[63370]_ , \new_[63371]_ , \new_[63375]_ ,
    \new_[63376]_ , \new_[63377]_ , \new_[63381]_ , \new_[63382]_ ,
    \new_[63385]_ , \new_[63388]_ , \new_[63389]_ , \new_[63390]_ ,
    \new_[63394]_ , \new_[63395]_ , \new_[63399]_ , \new_[63400]_ ,
    \new_[63401]_ , \new_[63405]_ , \new_[63406]_ , \new_[63409]_ ,
    \new_[63412]_ , \new_[63413]_ , \new_[63414]_ , \new_[63418]_ ,
    \new_[63419]_ , \new_[63423]_ , \new_[63424]_ , \new_[63425]_ ,
    \new_[63429]_ , \new_[63430]_ , \new_[63433]_ , \new_[63436]_ ,
    \new_[63437]_ , \new_[63438]_ , \new_[63442]_ , \new_[63443]_ ,
    \new_[63447]_ , \new_[63448]_ , \new_[63449]_ , \new_[63453]_ ,
    \new_[63454]_ , \new_[63457]_ , \new_[63460]_ , \new_[63461]_ ,
    \new_[63462]_ , \new_[63466]_ , \new_[63467]_ , \new_[63471]_ ,
    \new_[63472]_ , \new_[63473]_ , \new_[63477]_ , \new_[63478]_ ,
    \new_[63481]_ , \new_[63484]_ , \new_[63485]_ , \new_[63486]_ ,
    \new_[63490]_ , \new_[63491]_ , \new_[63495]_ , \new_[63496]_ ,
    \new_[63497]_ , \new_[63501]_ , \new_[63502]_ , \new_[63505]_ ,
    \new_[63508]_ , \new_[63509]_ , \new_[63510]_ , \new_[63514]_ ,
    \new_[63515]_ , \new_[63519]_ , \new_[63520]_ , \new_[63521]_ ,
    \new_[63525]_ , \new_[63526]_ , \new_[63529]_ , \new_[63532]_ ,
    \new_[63533]_ , \new_[63534]_ , \new_[63538]_ , \new_[63539]_ ,
    \new_[63543]_ , \new_[63544]_ , \new_[63545]_ , \new_[63549]_ ,
    \new_[63550]_ , \new_[63553]_ , \new_[63556]_ , \new_[63557]_ ,
    \new_[63558]_ , \new_[63562]_ , \new_[63563]_ , \new_[63567]_ ,
    \new_[63568]_ , \new_[63569]_ , \new_[63573]_ , \new_[63574]_ ,
    \new_[63577]_ , \new_[63580]_ , \new_[63581]_ , \new_[63582]_ ,
    \new_[63586]_ , \new_[63587]_ , \new_[63591]_ , \new_[63592]_ ,
    \new_[63593]_ , \new_[63597]_ , \new_[63598]_ , \new_[63601]_ ,
    \new_[63604]_ , \new_[63605]_ , \new_[63606]_ , \new_[63610]_ ,
    \new_[63611]_ , \new_[63615]_ , \new_[63616]_ , \new_[63617]_ ,
    \new_[63621]_ , \new_[63622]_ , \new_[63625]_ , \new_[63628]_ ,
    \new_[63629]_ , \new_[63630]_ , \new_[63634]_ , \new_[63635]_ ,
    \new_[63639]_ , \new_[63640]_ , \new_[63641]_ , \new_[63645]_ ,
    \new_[63646]_ , \new_[63649]_ , \new_[63652]_ , \new_[63653]_ ,
    \new_[63654]_ , \new_[63658]_ , \new_[63659]_ , \new_[63663]_ ,
    \new_[63664]_ , \new_[63665]_ , \new_[63669]_ , \new_[63670]_ ,
    \new_[63673]_ , \new_[63676]_ , \new_[63677]_ , \new_[63678]_ ,
    \new_[63682]_ , \new_[63683]_ , \new_[63687]_ , \new_[63688]_ ,
    \new_[63689]_ , \new_[63693]_ , \new_[63694]_ , \new_[63697]_ ,
    \new_[63700]_ , \new_[63701]_ , \new_[63702]_ , \new_[63706]_ ,
    \new_[63707]_ , \new_[63711]_ , \new_[63712]_ , \new_[63713]_ ,
    \new_[63717]_ , \new_[63718]_ , \new_[63721]_ , \new_[63724]_ ,
    \new_[63725]_ , \new_[63726]_ , \new_[63730]_ , \new_[63731]_ ,
    \new_[63735]_ , \new_[63736]_ , \new_[63737]_ , \new_[63741]_ ,
    \new_[63742]_ , \new_[63745]_ , \new_[63748]_ , \new_[63749]_ ,
    \new_[63750]_ , \new_[63754]_ , \new_[63755]_ , \new_[63759]_ ,
    \new_[63760]_ , \new_[63761]_ , \new_[63765]_ , \new_[63766]_ ,
    \new_[63769]_ , \new_[63772]_ , \new_[63773]_ , \new_[63774]_ ,
    \new_[63778]_ , \new_[63779]_ , \new_[63783]_ , \new_[63784]_ ,
    \new_[63785]_ , \new_[63789]_ , \new_[63790]_ , \new_[63793]_ ,
    \new_[63796]_ , \new_[63797]_ , \new_[63798]_ , \new_[63802]_ ,
    \new_[63803]_ , \new_[63807]_ , \new_[63808]_ , \new_[63809]_ ,
    \new_[63813]_ , \new_[63814]_ , \new_[63817]_ , \new_[63820]_ ,
    \new_[63821]_ , \new_[63822]_ , \new_[63826]_ , \new_[63827]_ ,
    \new_[63831]_ , \new_[63832]_ , \new_[63833]_ , \new_[63837]_ ,
    \new_[63838]_ , \new_[63841]_ , \new_[63844]_ , \new_[63845]_ ,
    \new_[63846]_ , \new_[63850]_ , \new_[63851]_ , \new_[63855]_ ,
    \new_[63856]_ , \new_[63857]_ , \new_[63861]_ , \new_[63862]_ ,
    \new_[63865]_ , \new_[63868]_ , \new_[63869]_ , \new_[63870]_ ,
    \new_[63874]_ , \new_[63875]_ , \new_[63879]_ , \new_[63880]_ ,
    \new_[63881]_ , \new_[63885]_ , \new_[63886]_ , \new_[63889]_ ,
    \new_[63892]_ , \new_[63893]_ , \new_[63894]_ , \new_[63898]_ ,
    \new_[63899]_ , \new_[63903]_ , \new_[63904]_ , \new_[63905]_ ,
    \new_[63909]_ , \new_[63910]_ , \new_[63913]_ , \new_[63916]_ ,
    \new_[63917]_ , \new_[63918]_ , \new_[63922]_ , \new_[63923]_ ,
    \new_[63927]_ , \new_[63928]_ , \new_[63929]_ , \new_[63933]_ ,
    \new_[63934]_ , \new_[63937]_ , \new_[63940]_ , \new_[63941]_ ,
    \new_[63942]_ , \new_[63946]_ , \new_[63947]_ , \new_[63951]_ ,
    \new_[63952]_ , \new_[63953]_ , \new_[63957]_ , \new_[63958]_ ,
    \new_[63961]_ , \new_[63964]_ , \new_[63965]_ , \new_[63966]_ ,
    \new_[63970]_ , \new_[63971]_ , \new_[63975]_ , \new_[63976]_ ,
    \new_[63977]_ , \new_[63981]_ , \new_[63982]_ , \new_[63985]_ ,
    \new_[63988]_ , \new_[63989]_ , \new_[63990]_ , \new_[63994]_ ,
    \new_[63995]_ , \new_[63999]_ , \new_[64000]_ , \new_[64001]_ ,
    \new_[64005]_ , \new_[64006]_ , \new_[64009]_ , \new_[64012]_ ,
    \new_[64013]_ , \new_[64014]_ , \new_[64018]_ , \new_[64019]_ ,
    \new_[64023]_ , \new_[64024]_ , \new_[64025]_ , \new_[64029]_ ,
    \new_[64030]_ , \new_[64033]_ , \new_[64036]_ , \new_[64037]_ ,
    \new_[64038]_ , \new_[64042]_ , \new_[64043]_ , \new_[64047]_ ,
    \new_[64048]_ , \new_[64049]_ , \new_[64053]_ , \new_[64054]_ ,
    \new_[64057]_ , \new_[64060]_ , \new_[64061]_ , \new_[64062]_ ,
    \new_[64066]_ , \new_[64067]_ , \new_[64071]_ , \new_[64072]_ ,
    \new_[64073]_ , \new_[64077]_ , \new_[64078]_ , \new_[64081]_ ,
    \new_[64084]_ , \new_[64085]_ , \new_[64086]_ , \new_[64090]_ ,
    \new_[64091]_ , \new_[64095]_ , \new_[64096]_ , \new_[64097]_ ,
    \new_[64101]_ , \new_[64102]_ , \new_[64105]_ , \new_[64108]_ ,
    \new_[64109]_ , \new_[64110]_ , \new_[64114]_ , \new_[64115]_ ,
    \new_[64119]_ , \new_[64120]_ , \new_[64121]_ , \new_[64125]_ ,
    \new_[64126]_ , \new_[64129]_ , \new_[64132]_ , \new_[64133]_ ,
    \new_[64134]_ , \new_[64138]_ , \new_[64139]_ , \new_[64143]_ ,
    \new_[64144]_ , \new_[64145]_ , \new_[64149]_ , \new_[64150]_ ,
    \new_[64153]_ , \new_[64156]_ , \new_[64157]_ , \new_[64158]_ ,
    \new_[64162]_ , \new_[64163]_ , \new_[64167]_ , \new_[64168]_ ,
    \new_[64169]_ , \new_[64173]_ , \new_[64174]_ , \new_[64177]_ ,
    \new_[64180]_ , \new_[64181]_ , \new_[64182]_ , \new_[64186]_ ,
    \new_[64187]_ , \new_[64191]_ , \new_[64192]_ , \new_[64193]_ ,
    \new_[64197]_ , \new_[64198]_ , \new_[64201]_ , \new_[64204]_ ,
    \new_[64205]_ , \new_[64206]_ , \new_[64210]_ , \new_[64211]_ ,
    \new_[64215]_ , \new_[64216]_ , \new_[64217]_ , \new_[64221]_ ,
    \new_[64222]_ , \new_[64225]_ , \new_[64228]_ , \new_[64229]_ ,
    \new_[64230]_ , \new_[64234]_ , \new_[64235]_ , \new_[64239]_ ,
    \new_[64240]_ , \new_[64241]_ , \new_[64245]_ , \new_[64246]_ ,
    \new_[64249]_ , \new_[64252]_ , \new_[64253]_ , \new_[64254]_ ,
    \new_[64258]_ , \new_[64259]_ , \new_[64263]_ , \new_[64264]_ ,
    \new_[64265]_ , \new_[64269]_ , \new_[64270]_ , \new_[64273]_ ,
    \new_[64276]_ , \new_[64277]_ , \new_[64278]_ , \new_[64282]_ ,
    \new_[64283]_ , \new_[64287]_ , \new_[64288]_ , \new_[64289]_ ,
    \new_[64293]_ , \new_[64294]_ , \new_[64297]_ , \new_[64300]_ ,
    \new_[64301]_ , \new_[64302]_ , \new_[64306]_ , \new_[64307]_ ,
    \new_[64311]_ , \new_[64312]_ , \new_[64313]_ , \new_[64317]_ ,
    \new_[64318]_ , \new_[64321]_ , \new_[64324]_ , \new_[64325]_ ,
    \new_[64326]_ , \new_[64330]_ , \new_[64331]_ , \new_[64335]_ ,
    \new_[64336]_ , \new_[64337]_ , \new_[64341]_ , \new_[64342]_ ,
    \new_[64345]_ , \new_[64348]_ , \new_[64349]_ , \new_[64350]_ ,
    \new_[64354]_ , \new_[64355]_ , \new_[64359]_ , \new_[64360]_ ,
    \new_[64361]_ , \new_[64365]_ , \new_[64366]_ , \new_[64369]_ ,
    \new_[64372]_ , \new_[64373]_ , \new_[64374]_ , \new_[64378]_ ,
    \new_[64379]_ , \new_[64383]_ , \new_[64384]_ , \new_[64385]_ ,
    \new_[64389]_ , \new_[64390]_ , \new_[64393]_ , \new_[64396]_ ,
    \new_[64397]_ , \new_[64398]_ , \new_[64402]_ , \new_[64403]_ ,
    \new_[64407]_ , \new_[64408]_ , \new_[64409]_ , \new_[64413]_ ,
    \new_[64414]_ , \new_[64417]_ , \new_[64420]_ , \new_[64421]_ ,
    \new_[64422]_ , \new_[64426]_ , \new_[64427]_ , \new_[64431]_ ,
    \new_[64432]_ , \new_[64433]_ , \new_[64437]_ , \new_[64438]_ ,
    \new_[64441]_ , \new_[64444]_ , \new_[64445]_ , \new_[64446]_ ,
    \new_[64450]_ , \new_[64451]_ , \new_[64455]_ , \new_[64456]_ ,
    \new_[64457]_ , \new_[64461]_ , \new_[64462]_ , \new_[64465]_ ,
    \new_[64468]_ , \new_[64469]_ , \new_[64470]_ , \new_[64474]_ ,
    \new_[64475]_ , \new_[64479]_ , \new_[64480]_ , \new_[64481]_ ,
    \new_[64485]_ , \new_[64486]_ , \new_[64489]_ , \new_[64492]_ ,
    \new_[64493]_ , \new_[64494]_ , \new_[64498]_ , \new_[64499]_ ,
    \new_[64503]_ , \new_[64504]_ , \new_[64505]_ , \new_[64509]_ ,
    \new_[64510]_ , \new_[64513]_ , \new_[64516]_ , \new_[64517]_ ,
    \new_[64518]_ , \new_[64522]_ , \new_[64523]_ , \new_[64527]_ ,
    \new_[64528]_ , \new_[64529]_ , \new_[64533]_ , \new_[64534]_ ,
    \new_[64537]_ , \new_[64540]_ , \new_[64541]_ , \new_[64542]_ ,
    \new_[64546]_ , \new_[64547]_ , \new_[64551]_ , \new_[64552]_ ,
    \new_[64553]_ , \new_[64557]_ , \new_[64558]_ , \new_[64561]_ ,
    \new_[64564]_ , \new_[64565]_ , \new_[64566]_ , \new_[64570]_ ,
    \new_[64571]_ , \new_[64575]_ , \new_[64576]_ , \new_[64577]_ ,
    \new_[64581]_ , \new_[64582]_ , \new_[64585]_ , \new_[64588]_ ,
    \new_[64589]_ , \new_[64590]_ , \new_[64594]_ , \new_[64595]_ ,
    \new_[64599]_ , \new_[64600]_ , \new_[64601]_ , \new_[64605]_ ,
    \new_[64606]_ , \new_[64609]_ , \new_[64612]_ , \new_[64613]_ ,
    \new_[64614]_ , \new_[64618]_ , \new_[64619]_ , \new_[64623]_ ,
    \new_[64624]_ , \new_[64625]_ , \new_[64629]_ , \new_[64630]_ ,
    \new_[64633]_ , \new_[64636]_ , \new_[64637]_ , \new_[64638]_ ,
    \new_[64642]_ , \new_[64643]_ , \new_[64646]_ , \new_[64649]_ ,
    \new_[64650]_ , \new_[64651]_ , \new_[64655]_ , \new_[64656]_ ,
    \new_[64659]_ , \new_[64662]_ , \new_[64663]_ , \new_[64664]_ ,
    \new_[64668]_ , \new_[64669]_ , \new_[64672]_ , \new_[64675]_ ,
    \new_[64676]_ , \new_[64677]_ , \new_[64681]_ , \new_[64682]_ ,
    \new_[64685]_ , \new_[64688]_ , \new_[64689]_ , \new_[64690]_ ,
    \new_[64694]_ , \new_[64695]_ , \new_[64698]_ , \new_[64701]_ ,
    \new_[64702]_ , \new_[64703]_ , \new_[64707]_ , \new_[64708]_ ,
    \new_[64711]_ , \new_[64714]_ , \new_[64715]_ , \new_[64716]_ ,
    \new_[64720]_ , \new_[64721]_ , \new_[64724]_ , \new_[64727]_ ,
    \new_[64728]_ , \new_[64729]_ , \new_[64733]_ , \new_[64734]_ ,
    \new_[64737]_ , \new_[64740]_ , \new_[64741]_ , \new_[64742]_ ,
    \new_[64746]_ , \new_[64747]_ , \new_[64750]_ , \new_[64753]_ ,
    \new_[64754]_ , \new_[64755]_ , \new_[64759]_ , \new_[64760]_ ,
    \new_[64763]_ , \new_[64766]_ , \new_[64767]_ , \new_[64768]_ ,
    \new_[64772]_ , \new_[64773]_ , \new_[64776]_ , \new_[64779]_ ,
    \new_[64780]_ , \new_[64781]_ , \new_[64785]_ , \new_[64786]_ ,
    \new_[64789]_ , \new_[64792]_ , \new_[64793]_ , \new_[64794]_ ,
    \new_[64798]_ , \new_[64799]_ , \new_[64802]_ , \new_[64805]_ ,
    \new_[64806]_ , \new_[64807]_ , \new_[64811]_ , \new_[64812]_ ,
    \new_[64815]_ , \new_[64818]_ , \new_[64819]_ , \new_[64820]_ ,
    \new_[64824]_ , \new_[64825]_ , \new_[64828]_ , \new_[64831]_ ,
    \new_[64832]_ , \new_[64833]_ , \new_[64837]_ , \new_[64838]_ ,
    \new_[64841]_ , \new_[64844]_ , \new_[64845]_ , \new_[64846]_ ,
    \new_[64850]_ , \new_[64851]_ , \new_[64854]_ , \new_[64857]_ ,
    \new_[64858]_ , \new_[64859]_ , \new_[64863]_ , \new_[64864]_ ,
    \new_[64867]_ , \new_[64870]_ , \new_[64871]_ , \new_[64872]_ ,
    \new_[64876]_ , \new_[64877]_ , \new_[64880]_ , \new_[64883]_ ,
    \new_[64884]_ , \new_[64885]_ , \new_[64889]_ , \new_[64890]_ ,
    \new_[64893]_ , \new_[64896]_ , \new_[64897]_ , \new_[64898]_ ,
    \new_[64902]_ , \new_[64903]_ , \new_[64906]_ , \new_[64909]_ ,
    \new_[64910]_ , \new_[64911]_ , \new_[64915]_ , \new_[64916]_ ,
    \new_[64919]_ , \new_[64922]_ , \new_[64923]_ , \new_[64924]_ ,
    \new_[64928]_ , \new_[64929]_ , \new_[64932]_ , \new_[64935]_ ,
    \new_[64936]_ , \new_[64937]_ , \new_[64941]_ , \new_[64942]_ ,
    \new_[64945]_ , \new_[64948]_ , \new_[64949]_ , \new_[64950]_ ,
    \new_[64954]_ , \new_[64955]_ , \new_[64958]_ , \new_[64961]_ ,
    \new_[64962]_ , \new_[64963]_ , \new_[64967]_ , \new_[64968]_ ,
    \new_[64971]_ , \new_[64974]_ , \new_[64975]_ , \new_[64976]_ ,
    \new_[64980]_ , \new_[64981]_ , \new_[64984]_ , \new_[64987]_ ,
    \new_[64988]_ , \new_[64989]_ , \new_[64993]_ , \new_[64994]_ ,
    \new_[64997]_ , \new_[65000]_ , \new_[65001]_ , \new_[65002]_ ,
    \new_[65006]_ , \new_[65007]_ , \new_[65010]_ , \new_[65013]_ ,
    \new_[65014]_ , \new_[65015]_ , \new_[65019]_ , \new_[65020]_ ,
    \new_[65023]_ , \new_[65026]_ , \new_[65027]_ , \new_[65028]_ ,
    \new_[65032]_ , \new_[65033]_ , \new_[65036]_ , \new_[65039]_ ,
    \new_[65040]_ , \new_[65041]_ , \new_[65045]_ , \new_[65046]_ ,
    \new_[65049]_ , \new_[65052]_ , \new_[65053]_ , \new_[65054]_ ,
    \new_[65058]_ , \new_[65059]_ , \new_[65062]_ , \new_[65065]_ ,
    \new_[65066]_ , \new_[65067]_ , \new_[65071]_ , \new_[65072]_ ,
    \new_[65075]_ , \new_[65078]_ , \new_[65079]_ , \new_[65080]_ ,
    \new_[65084]_ , \new_[65085]_ , \new_[65088]_ , \new_[65091]_ ,
    \new_[65092]_ , \new_[65093]_ , \new_[65097]_ , \new_[65098]_ ,
    \new_[65101]_ , \new_[65104]_ , \new_[65105]_ , \new_[65106]_ ,
    \new_[65110]_ , \new_[65111]_ , \new_[65114]_ , \new_[65117]_ ,
    \new_[65118]_ , \new_[65119]_ , \new_[65123]_ , \new_[65124]_ ,
    \new_[65127]_ , \new_[65130]_ , \new_[65131]_ , \new_[65132]_ ,
    \new_[65136]_ , \new_[65137]_ , \new_[65140]_ , \new_[65143]_ ,
    \new_[65144]_ , \new_[65145]_ , \new_[65149]_ , \new_[65150]_ ,
    \new_[65153]_ , \new_[65156]_ , \new_[65157]_ , \new_[65158]_ ,
    \new_[65162]_ , \new_[65163]_ , \new_[65166]_ , \new_[65169]_ ,
    \new_[65170]_ , \new_[65171]_ , \new_[65175]_ , \new_[65176]_ ,
    \new_[65179]_ , \new_[65182]_ , \new_[65183]_ , \new_[65184]_ ,
    \new_[65188]_ , \new_[65189]_ , \new_[65192]_ , \new_[65195]_ ,
    \new_[65196]_ , \new_[65197]_ , \new_[65201]_ , \new_[65202]_ ,
    \new_[65205]_ , \new_[65208]_ , \new_[65209]_ , \new_[65210]_ ,
    \new_[65214]_ , \new_[65215]_ , \new_[65218]_ , \new_[65221]_ ,
    \new_[65222]_ , \new_[65223]_ , \new_[65227]_ , \new_[65228]_ ,
    \new_[65231]_ , \new_[65234]_ , \new_[65235]_ , \new_[65236]_ ,
    \new_[65240]_ , \new_[65241]_ , \new_[65244]_ , \new_[65247]_ ,
    \new_[65248]_ , \new_[65249]_ , \new_[65253]_ , \new_[65254]_ ,
    \new_[65257]_ , \new_[65260]_ , \new_[65261]_ , \new_[65262]_ ,
    \new_[65266]_ , \new_[65267]_ , \new_[65270]_ , \new_[65273]_ ,
    \new_[65274]_ , \new_[65275]_ , \new_[65279]_ , \new_[65280]_ ,
    \new_[65283]_ , \new_[65286]_ , \new_[65287]_ , \new_[65288]_ ,
    \new_[65292]_ , \new_[65293]_ , \new_[65296]_ , \new_[65299]_ ,
    \new_[65300]_ , \new_[65301]_ , \new_[65305]_ , \new_[65306]_ ,
    \new_[65309]_ , \new_[65312]_ , \new_[65313]_ , \new_[65314]_ ,
    \new_[65318]_ , \new_[65319]_ , \new_[65322]_ , \new_[65325]_ ,
    \new_[65326]_ , \new_[65327]_ , \new_[65331]_ , \new_[65332]_ ,
    \new_[65335]_ , \new_[65338]_ , \new_[65339]_ , \new_[65340]_ ,
    \new_[65344]_ , \new_[65345]_ , \new_[65348]_ , \new_[65351]_ ,
    \new_[65352]_ , \new_[65353]_ , \new_[65357]_ , \new_[65358]_ ,
    \new_[65361]_ , \new_[65364]_ , \new_[65365]_ , \new_[65366]_ ,
    \new_[65370]_ , \new_[65371]_ , \new_[65374]_ , \new_[65377]_ ,
    \new_[65378]_ , \new_[65379]_ , \new_[65383]_ , \new_[65384]_ ,
    \new_[65387]_ , \new_[65390]_ , \new_[65391]_ , \new_[65392]_ ,
    \new_[65396]_ , \new_[65397]_ , \new_[65400]_ , \new_[65403]_ ,
    \new_[65404]_ , \new_[65405]_ , \new_[65409]_ , \new_[65410]_ ,
    \new_[65413]_ , \new_[65416]_ , \new_[65417]_ , \new_[65418]_ ,
    \new_[65422]_ , \new_[65423]_ , \new_[65426]_ , \new_[65429]_ ,
    \new_[65430]_ , \new_[65431]_ , \new_[65435]_ , \new_[65436]_ ,
    \new_[65439]_ , \new_[65442]_ , \new_[65443]_ , \new_[65444]_ ,
    \new_[65448]_ , \new_[65449]_ , \new_[65452]_ , \new_[65455]_ ,
    \new_[65456]_ , \new_[65457]_ , \new_[65461]_ , \new_[65462]_ ,
    \new_[65465]_ , \new_[65468]_ , \new_[65469]_ , \new_[65470]_ ,
    \new_[65474]_ , \new_[65475]_ , \new_[65478]_ , \new_[65481]_ ,
    \new_[65482]_ , \new_[65483]_ , \new_[65487]_ , \new_[65488]_ ,
    \new_[65491]_ , \new_[65494]_ , \new_[65495]_ , \new_[65496]_ ,
    \new_[65500]_ , \new_[65501]_ , \new_[65504]_ , \new_[65507]_ ,
    \new_[65508]_ , \new_[65509]_ , \new_[65513]_ , \new_[65514]_ ,
    \new_[65517]_ , \new_[65520]_ , \new_[65521]_ , \new_[65522]_ ,
    \new_[65526]_ , \new_[65527]_ , \new_[65530]_ , \new_[65533]_ ,
    \new_[65534]_ , \new_[65535]_ , \new_[65539]_ , \new_[65540]_ ,
    \new_[65543]_ , \new_[65546]_ , \new_[65547]_ , \new_[65548]_ ,
    \new_[65552]_ , \new_[65553]_ , \new_[65556]_ , \new_[65559]_ ,
    \new_[65560]_ , \new_[65561]_ , \new_[65565]_ , \new_[65566]_ ,
    \new_[65569]_ , \new_[65572]_ , \new_[65573]_ , \new_[65574]_ ,
    \new_[65578]_ , \new_[65579]_ , \new_[65582]_ , \new_[65585]_ ,
    \new_[65586]_ , \new_[65587]_ , \new_[65591]_ , \new_[65592]_ ,
    \new_[65595]_ , \new_[65598]_ , \new_[65599]_ , \new_[65600]_ ,
    \new_[65604]_ , \new_[65605]_ , \new_[65608]_ , \new_[65611]_ ,
    \new_[65612]_ , \new_[65613]_ , \new_[65617]_ , \new_[65618]_ ,
    \new_[65621]_ , \new_[65624]_ , \new_[65625]_ , \new_[65626]_ ,
    \new_[65630]_ , \new_[65631]_ , \new_[65634]_ , \new_[65637]_ ,
    \new_[65638]_ , \new_[65639]_ , \new_[65643]_ , \new_[65644]_ ,
    \new_[65647]_ , \new_[65650]_ , \new_[65651]_ , \new_[65652]_ ,
    \new_[65656]_ , \new_[65657]_ , \new_[65660]_ , \new_[65663]_ ,
    \new_[65664]_ , \new_[65665]_ , \new_[65669]_ , \new_[65670]_ ,
    \new_[65673]_ , \new_[65676]_ , \new_[65677]_ , \new_[65678]_ ,
    \new_[65682]_ , \new_[65683]_ , \new_[65686]_ , \new_[65689]_ ,
    \new_[65690]_ , \new_[65691]_ , \new_[65695]_ , \new_[65696]_ ,
    \new_[65699]_ , \new_[65702]_ , \new_[65703]_ , \new_[65704]_ ,
    \new_[65708]_ , \new_[65709]_ , \new_[65712]_ , \new_[65715]_ ,
    \new_[65716]_ , \new_[65717]_ , \new_[65721]_ , \new_[65722]_ ,
    \new_[65725]_ , \new_[65728]_ , \new_[65729]_ , \new_[65730]_ ,
    \new_[65734]_ , \new_[65735]_ , \new_[65738]_ , \new_[65741]_ ,
    \new_[65742]_ , \new_[65743]_ , \new_[65747]_ , \new_[65748]_ ,
    \new_[65751]_ , \new_[65754]_ , \new_[65755]_ , \new_[65756]_ ,
    \new_[65760]_ , \new_[65761]_ , \new_[65764]_ , \new_[65767]_ ,
    \new_[65768]_ , \new_[65769]_ , \new_[65773]_ , \new_[65774]_ ,
    \new_[65777]_ , \new_[65780]_ , \new_[65781]_ , \new_[65782]_ ,
    \new_[65786]_ , \new_[65787]_ , \new_[65790]_ , \new_[65793]_ ,
    \new_[65794]_ , \new_[65795]_ , \new_[65799]_ , \new_[65800]_ ,
    \new_[65803]_ , \new_[65806]_ , \new_[65807]_ , \new_[65808]_ ,
    \new_[65812]_ , \new_[65813]_ , \new_[65816]_ , \new_[65819]_ ,
    \new_[65820]_ , \new_[65821]_ , \new_[65825]_ , \new_[65826]_ ,
    \new_[65829]_ , \new_[65832]_ , \new_[65833]_ , \new_[65834]_ ,
    \new_[65838]_ , \new_[65839]_ , \new_[65842]_ , \new_[65845]_ ,
    \new_[65846]_ , \new_[65847]_ , \new_[65851]_ , \new_[65852]_ ,
    \new_[65855]_ , \new_[65858]_ , \new_[65859]_ , \new_[65860]_ ,
    \new_[65864]_ , \new_[65865]_ , \new_[65868]_ , \new_[65871]_ ,
    \new_[65872]_ , \new_[65873]_ , \new_[65877]_ , \new_[65878]_ ,
    \new_[65881]_ , \new_[65884]_ , \new_[65885]_ , \new_[65886]_ ,
    \new_[65890]_ , \new_[65891]_ , \new_[65894]_ , \new_[65897]_ ,
    \new_[65898]_ , \new_[65899]_ , \new_[65903]_ , \new_[65904]_ ,
    \new_[65907]_ , \new_[65910]_ , \new_[65911]_ , \new_[65912]_ ,
    \new_[65916]_ , \new_[65917]_ , \new_[65920]_ , \new_[65923]_ ,
    \new_[65924]_ , \new_[65925]_ , \new_[65929]_ , \new_[65930]_ ,
    \new_[65933]_ , \new_[65936]_ , \new_[65937]_ , \new_[65938]_ ,
    \new_[65942]_ , \new_[65943]_ , \new_[65946]_ , \new_[65949]_ ,
    \new_[65950]_ , \new_[65951]_ , \new_[65955]_ , \new_[65956]_ ,
    \new_[65959]_ , \new_[65962]_ , \new_[65963]_ , \new_[65964]_ ,
    \new_[65968]_ , \new_[65969]_ , \new_[65972]_ , \new_[65975]_ ,
    \new_[65976]_ , \new_[65977]_ , \new_[65981]_ , \new_[65982]_ ,
    \new_[65985]_ , \new_[65988]_ , \new_[65989]_ , \new_[65990]_ ,
    \new_[65994]_ , \new_[65995]_ , \new_[65998]_ , \new_[66001]_ ,
    \new_[66002]_ , \new_[66003]_ , \new_[66007]_ , \new_[66008]_ ,
    \new_[66011]_ , \new_[66014]_ , \new_[66015]_ , \new_[66016]_ ,
    \new_[66020]_ , \new_[66021]_ , \new_[66024]_ , \new_[66027]_ ,
    \new_[66028]_ , \new_[66029]_ , \new_[66033]_ , \new_[66034]_ ,
    \new_[66037]_ , \new_[66040]_ , \new_[66041]_ , \new_[66042]_ ,
    \new_[66046]_ , \new_[66047]_ , \new_[66050]_ , \new_[66053]_ ,
    \new_[66054]_ , \new_[66055]_ , \new_[66059]_ , \new_[66060]_ ,
    \new_[66063]_ , \new_[66066]_ , \new_[66067]_ , \new_[66068]_ ,
    \new_[66072]_ , \new_[66073]_ , \new_[66076]_ , \new_[66079]_ ,
    \new_[66080]_ , \new_[66081]_ , \new_[66085]_ , \new_[66086]_ ,
    \new_[66089]_ , \new_[66092]_ , \new_[66093]_ , \new_[66094]_ ,
    \new_[66098]_ , \new_[66099]_ , \new_[66102]_ , \new_[66105]_ ,
    \new_[66106]_ , \new_[66107]_ , \new_[66111]_ , \new_[66112]_ ,
    \new_[66115]_ , \new_[66118]_ , \new_[66119]_ , \new_[66120]_ ,
    \new_[66124]_ , \new_[66125]_ , \new_[66128]_ , \new_[66131]_ ,
    \new_[66132]_ , \new_[66133]_ , \new_[66137]_ , \new_[66138]_ ,
    \new_[66141]_ , \new_[66144]_ , \new_[66145]_ , \new_[66146]_ ,
    \new_[66150]_ , \new_[66151]_ , \new_[66154]_ , \new_[66157]_ ,
    \new_[66158]_ , \new_[66159]_ , \new_[66163]_ , \new_[66164]_ ,
    \new_[66167]_ , \new_[66170]_ , \new_[66171]_ , \new_[66172]_ ,
    \new_[66176]_ , \new_[66177]_ , \new_[66180]_ , \new_[66183]_ ,
    \new_[66184]_ , \new_[66185]_ , \new_[66189]_ , \new_[66190]_ ,
    \new_[66193]_ , \new_[66196]_ , \new_[66197]_ , \new_[66198]_ ,
    \new_[66202]_ , \new_[66203]_ , \new_[66206]_ , \new_[66209]_ ,
    \new_[66210]_ , \new_[66211]_ , \new_[66215]_ , \new_[66216]_ ,
    \new_[66219]_ , \new_[66222]_ , \new_[66223]_ , \new_[66224]_ ,
    \new_[66228]_ , \new_[66229]_ , \new_[66232]_ , \new_[66235]_ ,
    \new_[66236]_ , \new_[66237]_ , \new_[66241]_ , \new_[66242]_ ,
    \new_[66245]_ , \new_[66248]_ , \new_[66249]_ , \new_[66250]_ ,
    \new_[66254]_ , \new_[66255]_ , \new_[66258]_ , \new_[66261]_ ,
    \new_[66262]_ , \new_[66263]_ , \new_[66267]_ , \new_[66268]_ ,
    \new_[66271]_ , \new_[66274]_ , \new_[66275]_ , \new_[66276]_ ,
    \new_[66280]_ , \new_[66281]_ , \new_[66284]_ , \new_[66287]_ ,
    \new_[66288]_ , \new_[66289]_ , \new_[66293]_ , \new_[66294]_ ,
    \new_[66297]_ , \new_[66300]_ , \new_[66301]_ , \new_[66302]_ ,
    \new_[66306]_ , \new_[66307]_ , \new_[66310]_ , \new_[66313]_ ,
    \new_[66314]_ , \new_[66315]_ , \new_[66319]_ , \new_[66320]_ ,
    \new_[66323]_ , \new_[66326]_ , \new_[66327]_ , \new_[66328]_ ,
    \new_[66332]_ , \new_[66333]_ , \new_[66336]_ , \new_[66339]_ ,
    \new_[66340]_ , \new_[66341]_ , \new_[66345]_ , \new_[66346]_ ,
    \new_[66349]_ , \new_[66352]_ , \new_[66353]_ , \new_[66354]_ ,
    \new_[66358]_ , \new_[66359]_ , \new_[66362]_ , \new_[66365]_ ,
    \new_[66366]_ , \new_[66367]_ , \new_[66371]_ , \new_[66372]_ ,
    \new_[66375]_ , \new_[66378]_ , \new_[66379]_ , \new_[66380]_ ,
    \new_[66384]_ , \new_[66385]_ , \new_[66388]_ , \new_[66391]_ ,
    \new_[66392]_ , \new_[66393]_ , \new_[66397]_ , \new_[66398]_ ,
    \new_[66401]_ , \new_[66404]_ , \new_[66405]_ , \new_[66406]_ ,
    \new_[66410]_ , \new_[66411]_ , \new_[66414]_ , \new_[66417]_ ,
    \new_[66418]_ , \new_[66419]_ , \new_[66423]_ , \new_[66424]_ ,
    \new_[66427]_ , \new_[66430]_ , \new_[66431]_ , \new_[66432]_ ,
    \new_[66436]_ , \new_[66437]_ , \new_[66440]_ , \new_[66443]_ ,
    \new_[66444]_ , \new_[66445]_ , \new_[66449]_ , \new_[66450]_ ,
    \new_[66453]_ , \new_[66456]_ , \new_[66457]_ , \new_[66458]_ ,
    \new_[66462]_ , \new_[66463]_ , \new_[66466]_ , \new_[66469]_ ,
    \new_[66470]_ , \new_[66471]_ , \new_[66475]_ , \new_[66476]_ ,
    \new_[66479]_ , \new_[66482]_ , \new_[66483]_ , \new_[66484]_ ,
    \new_[66488]_ , \new_[66489]_ , \new_[66492]_ , \new_[66495]_ ,
    \new_[66496]_ , \new_[66497]_ , \new_[66501]_ , \new_[66502]_ ,
    \new_[66505]_ , \new_[66508]_ , \new_[66509]_ , \new_[66510]_ ,
    \new_[66514]_ , \new_[66515]_ , \new_[66518]_ , \new_[66521]_ ,
    \new_[66522]_ , \new_[66523]_ , \new_[66527]_ , \new_[66528]_ ,
    \new_[66531]_ , \new_[66534]_ , \new_[66535]_ , \new_[66536]_ ,
    \new_[66540]_ , \new_[66541]_ , \new_[66544]_ , \new_[66547]_ ,
    \new_[66548]_ , \new_[66549]_ , \new_[66553]_ , \new_[66554]_ ,
    \new_[66557]_ , \new_[66560]_ , \new_[66561]_ , \new_[66562]_ ,
    \new_[66566]_ , \new_[66567]_ , \new_[66570]_ , \new_[66573]_ ,
    \new_[66574]_ , \new_[66575]_ , \new_[66579]_ , \new_[66580]_ ,
    \new_[66583]_ , \new_[66586]_ , \new_[66587]_ , \new_[66588]_ ,
    \new_[66592]_ , \new_[66593]_ , \new_[66596]_ , \new_[66599]_ ,
    \new_[66600]_ , \new_[66601]_ , \new_[66605]_ , \new_[66606]_ ,
    \new_[66609]_ , \new_[66612]_ , \new_[66613]_ , \new_[66614]_ ,
    \new_[66618]_ , \new_[66619]_ , \new_[66622]_ , \new_[66625]_ ,
    \new_[66626]_ , \new_[66627]_ , \new_[66631]_ , \new_[66632]_ ,
    \new_[66635]_ , \new_[66638]_ , \new_[66639]_ , \new_[66640]_ ,
    \new_[66644]_ , \new_[66645]_ , \new_[66648]_ , \new_[66651]_ ,
    \new_[66652]_ , \new_[66653]_ , \new_[66657]_ , \new_[66658]_ ,
    \new_[66661]_ , \new_[66664]_ , \new_[66665]_ , \new_[66666]_ ,
    \new_[66670]_ , \new_[66671]_ , \new_[66674]_ , \new_[66677]_ ,
    \new_[66678]_ , \new_[66679]_ , \new_[66683]_ , \new_[66684]_ ,
    \new_[66687]_ , \new_[66690]_ , \new_[66691]_ , \new_[66692]_ ,
    \new_[66696]_ , \new_[66697]_ , \new_[66700]_ , \new_[66703]_ ,
    \new_[66704]_ , \new_[66705]_ , \new_[66709]_ , \new_[66710]_ ,
    \new_[66713]_ , \new_[66716]_ , \new_[66717]_ , \new_[66718]_ ,
    \new_[66722]_ , \new_[66723]_ , \new_[66726]_ , \new_[66729]_ ,
    \new_[66730]_ , \new_[66731]_ , \new_[66735]_ , \new_[66736]_ ,
    \new_[66739]_ , \new_[66742]_ , \new_[66743]_ , \new_[66744]_ ,
    \new_[66748]_ , \new_[66749]_ , \new_[66752]_ , \new_[66755]_ ,
    \new_[66756]_ , \new_[66757]_ , \new_[66761]_ , \new_[66762]_ ,
    \new_[66765]_ , \new_[66768]_ , \new_[66769]_ , \new_[66770]_ ,
    \new_[66774]_ , \new_[66775]_ , \new_[66778]_ , \new_[66781]_ ,
    \new_[66782]_ , \new_[66783]_ , \new_[66787]_ , \new_[66788]_ ,
    \new_[66791]_ , \new_[66794]_ , \new_[66795]_ , \new_[66796]_ ,
    \new_[66800]_ , \new_[66801]_ , \new_[66804]_ , \new_[66807]_ ,
    \new_[66808]_ , \new_[66809]_ , \new_[66813]_ , \new_[66814]_ ,
    \new_[66817]_ , \new_[66820]_ , \new_[66821]_ , \new_[66822]_ ,
    \new_[66826]_ , \new_[66827]_ , \new_[66830]_ , \new_[66833]_ ,
    \new_[66834]_ , \new_[66835]_ , \new_[66839]_ , \new_[66840]_ ,
    \new_[66843]_ , \new_[66846]_ , \new_[66847]_ , \new_[66848]_ ,
    \new_[66852]_ , \new_[66853]_ , \new_[66856]_ , \new_[66859]_ ,
    \new_[66860]_ , \new_[66861]_ , \new_[66865]_ , \new_[66866]_ ,
    \new_[66869]_ , \new_[66872]_ , \new_[66873]_ , \new_[66874]_ ,
    \new_[66878]_ , \new_[66879]_ , \new_[66882]_ , \new_[66885]_ ,
    \new_[66886]_ , \new_[66887]_ , \new_[66891]_ , \new_[66892]_ ,
    \new_[66895]_ , \new_[66898]_ , \new_[66899]_ , \new_[66900]_ ,
    \new_[66904]_ , \new_[66905]_ , \new_[66908]_ , \new_[66911]_ ,
    \new_[66912]_ , \new_[66913]_ , \new_[66917]_ , \new_[66918]_ ,
    \new_[66921]_ , \new_[66924]_ , \new_[66925]_ , \new_[66926]_ ,
    \new_[66930]_ , \new_[66931]_ , \new_[66934]_ , \new_[66937]_ ,
    \new_[66938]_ , \new_[66939]_ , \new_[66943]_ , \new_[66944]_ ,
    \new_[66947]_ , \new_[66950]_ , \new_[66951]_ , \new_[66952]_ ,
    \new_[66956]_ , \new_[66957]_ , \new_[66960]_ , \new_[66963]_ ,
    \new_[66964]_ , \new_[66965]_ , \new_[66969]_ , \new_[66970]_ ,
    \new_[66973]_ , \new_[66976]_ , \new_[66977]_ , \new_[66978]_ ,
    \new_[66982]_ , \new_[66983]_ , \new_[66986]_ , \new_[66989]_ ,
    \new_[66990]_ , \new_[66991]_ , \new_[66995]_ , \new_[66996]_ ,
    \new_[66999]_ , \new_[67002]_ , \new_[67003]_ , \new_[67004]_ ,
    \new_[67008]_ , \new_[67009]_ , \new_[67012]_ , \new_[67015]_ ,
    \new_[67016]_ , \new_[67017]_ , \new_[67021]_ , \new_[67022]_ ,
    \new_[67025]_ , \new_[67028]_ , \new_[67029]_ , \new_[67030]_ ,
    \new_[67034]_ , \new_[67035]_ , \new_[67038]_ , \new_[67041]_ ,
    \new_[67042]_ , \new_[67043]_ , \new_[67047]_ , \new_[67048]_ ,
    \new_[67051]_ , \new_[67054]_ , \new_[67055]_ , \new_[67056]_ ,
    \new_[67060]_ , \new_[67061]_ , \new_[67064]_ , \new_[67067]_ ,
    \new_[67068]_ , \new_[67069]_ , \new_[67073]_ , \new_[67074]_ ,
    \new_[67077]_ , \new_[67080]_ , \new_[67081]_ , \new_[67082]_ ,
    \new_[67086]_ , \new_[67087]_ , \new_[67090]_ , \new_[67093]_ ,
    \new_[67094]_ , \new_[67095]_ , \new_[67099]_ , \new_[67100]_ ,
    \new_[67103]_ , \new_[67106]_ , \new_[67107]_ , \new_[67108]_ ,
    \new_[67112]_ , \new_[67113]_ , \new_[67116]_ , \new_[67119]_ ,
    \new_[67120]_ , \new_[67121]_ , \new_[67125]_ , \new_[67126]_ ,
    \new_[67129]_ , \new_[67132]_ , \new_[67133]_ , \new_[67134]_ ,
    \new_[67138]_ , \new_[67139]_ , \new_[67142]_ , \new_[67145]_ ,
    \new_[67146]_ , \new_[67147]_ , \new_[67151]_ , \new_[67152]_ ,
    \new_[67155]_ , \new_[67158]_ , \new_[67159]_ , \new_[67160]_ ,
    \new_[67164]_ , \new_[67165]_ , \new_[67168]_ , \new_[67171]_ ,
    \new_[67172]_ , \new_[67173]_ , \new_[67177]_ , \new_[67178]_ ,
    \new_[67181]_ , \new_[67184]_ , \new_[67185]_ , \new_[67186]_ ,
    \new_[67190]_ , \new_[67191]_ , \new_[67194]_ , \new_[67197]_ ,
    \new_[67198]_ , \new_[67199]_ , \new_[67203]_ , \new_[67204]_ ,
    \new_[67207]_ , \new_[67210]_ , \new_[67211]_ , \new_[67212]_ ,
    \new_[67216]_ , \new_[67217]_ , \new_[67220]_ , \new_[67223]_ ,
    \new_[67224]_ , \new_[67225]_ , \new_[67229]_ , \new_[67230]_ ,
    \new_[67233]_ , \new_[67236]_ , \new_[67237]_ , \new_[67238]_ ,
    \new_[67242]_ , \new_[67243]_ , \new_[67246]_ , \new_[67249]_ ,
    \new_[67250]_ , \new_[67251]_ , \new_[67255]_ , \new_[67256]_ ,
    \new_[67259]_ , \new_[67262]_ , \new_[67263]_ , \new_[67264]_ ,
    \new_[67268]_ , \new_[67269]_ , \new_[67272]_ , \new_[67275]_ ,
    \new_[67276]_ , \new_[67277]_ , \new_[67281]_ , \new_[67282]_ ,
    \new_[67285]_ , \new_[67288]_ , \new_[67289]_ , \new_[67290]_ ,
    \new_[67294]_ , \new_[67295]_ , \new_[67298]_ , \new_[67301]_ ,
    \new_[67302]_ , \new_[67303]_ , \new_[67307]_ , \new_[67308]_ ,
    \new_[67311]_ , \new_[67314]_ , \new_[67315]_ , \new_[67316]_ ,
    \new_[67320]_ , \new_[67321]_ , \new_[67324]_ , \new_[67327]_ ,
    \new_[67328]_ , \new_[67329]_ , \new_[67333]_ , \new_[67334]_ ,
    \new_[67337]_ , \new_[67340]_ , \new_[67341]_ , \new_[67342]_ ,
    \new_[67346]_ , \new_[67347]_ , \new_[67350]_ , \new_[67353]_ ,
    \new_[67354]_ , \new_[67355]_ , \new_[67359]_ , \new_[67360]_ ,
    \new_[67363]_ , \new_[67366]_ , \new_[67367]_ , \new_[67368]_ ,
    \new_[67372]_ , \new_[67373]_ , \new_[67376]_ , \new_[67379]_ ,
    \new_[67380]_ , \new_[67381]_ , \new_[67385]_ , \new_[67386]_ ,
    \new_[67389]_ , \new_[67392]_ , \new_[67393]_ , \new_[67394]_ ,
    \new_[67398]_ , \new_[67399]_ , \new_[67402]_ , \new_[67405]_ ,
    \new_[67406]_ , \new_[67407]_ , \new_[67411]_ , \new_[67412]_ ,
    \new_[67415]_ , \new_[67418]_ , \new_[67419]_ , \new_[67420]_ ,
    \new_[67424]_ , \new_[67425]_ , \new_[67428]_ , \new_[67431]_ ,
    \new_[67432]_ , \new_[67433]_ , \new_[67437]_ , \new_[67438]_ ,
    \new_[67441]_ , \new_[67444]_ , \new_[67445]_ , \new_[67446]_ ,
    \new_[67450]_ , \new_[67451]_ , \new_[67454]_ , \new_[67457]_ ,
    \new_[67458]_ , \new_[67459]_ , \new_[67463]_ , \new_[67464]_ ,
    \new_[67467]_ , \new_[67470]_ , \new_[67471]_ , \new_[67472]_ ,
    \new_[67476]_ , \new_[67477]_ , \new_[67480]_ , \new_[67483]_ ,
    \new_[67484]_ , \new_[67485]_ , \new_[67489]_ , \new_[67490]_ ,
    \new_[67493]_ , \new_[67496]_ , \new_[67497]_ , \new_[67498]_ ,
    \new_[67502]_ , \new_[67503]_ , \new_[67506]_ , \new_[67509]_ ,
    \new_[67510]_ , \new_[67511]_ , \new_[67515]_ , \new_[67516]_ ,
    \new_[67519]_ , \new_[67522]_ , \new_[67523]_ , \new_[67524]_ ,
    \new_[67528]_ , \new_[67529]_ , \new_[67532]_ , \new_[67535]_ ,
    \new_[67536]_ , \new_[67537]_ , \new_[67541]_ , \new_[67542]_ ,
    \new_[67545]_ , \new_[67548]_ , \new_[67549]_ , \new_[67550]_ ,
    \new_[67554]_ , \new_[67555]_ , \new_[67558]_ , \new_[67561]_ ,
    \new_[67562]_ , \new_[67563]_ , \new_[67567]_ , \new_[67568]_ ,
    \new_[67571]_ , \new_[67574]_ , \new_[67575]_ , \new_[67576]_ ,
    \new_[67580]_ , \new_[67581]_ , \new_[67584]_ , \new_[67587]_ ,
    \new_[67588]_ , \new_[67589]_ , \new_[67593]_ , \new_[67594]_ ,
    \new_[67597]_ , \new_[67600]_ , \new_[67601]_ , \new_[67602]_ ,
    \new_[67606]_ , \new_[67607]_ , \new_[67610]_ , \new_[67613]_ ,
    \new_[67614]_ , \new_[67615]_ , \new_[67619]_ , \new_[67620]_ ,
    \new_[67623]_ , \new_[67626]_ , \new_[67627]_ , \new_[67628]_ ,
    \new_[67632]_ , \new_[67633]_ , \new_[67636]_ , \new_[67639]_ ,
    \new_[67640]_ , \new_[67641]_ , \new_[67645]_ , \new_[67646]_ ,
    \new_[67649]_ , \new_[67652]_ , \new_[67653]_ , \new_[67654]_ ,
    \new_[67658]_ , \new_[67659]_ , \new_[67662]_ , \new_[67665]_ ,
    \new_[67666]_ , \new_[67667]_ , \new_[67671]_ , \new_[67672]_ ,
    \new_[67675]_ , \new_[67678]_ , \new_[67679]_ , \new_[67680]_ ,
    \new_[67684]_ , \new_[67685]_ , \new_[67688]_ , \new_[67691]_ ,
    \new_[67692]_ , \new_[67693]_ , \new_[67697]_ , \new_[67698]_ ,
    \new_[67701]_ , \new_[67704]_ , \new_[67705]_ , \new_[67706]_ ,
    \new_[67710]_ , \new_[67711]_ , \new_[67714]_ , \new_[67717]_ ,
    \new_[67718]_ , \new_[67719]_ , \new_[67723]_ , \new_[67724]_ ,
    \new_[67727]_ , \new_[67730]_ , \new_[67731]_ , \new_[67732]_ ,
    \new_[67736]_ , \new_[67737]_ , \new_[67740]_ , \new_[67743]_ ,
    \new_[67744]_ , \new_[67745]_ , \new_[67749]_ , \new_[67750]_ ,
    \new_[67753]_ , \new_[67756]_ , \new_[67757]_ , \new_[67758]_ ,
    \new_[67762]_ , \new_[67763]_ , \new_[67766]_ , \new_[67769]_ ,
    \new_[67770]_ , \new_[67771]_ , \new_[67775]_ , \new_[67776]_ ,
    \new_[67779]_ , \new_[67782]_ , \new_[67783]_ , \new_[67784]_ ,
    \new_[67788]_ , \new_[67789]_ , \new_[67792]_ , \new_[67795]_ ,
    \new_[67796]_ , \new_[67797]_ , \new_[67801]_ , \new_[67802]_ ,
    \new_[67805]_ , \new_[67808]_ , \new_[67809]_ , \new_[67810]_ ,
    \new_[67814]_ , \new_[67815]_ , \new_[67818]_ , \new_[67821]_ ,
    \new_[67822]_ , \new_[67823]_ , \new_[67827]_ , \new_[67828]_ ,
    \new_[67831]_ , \new_[67834]_ , \new_[67835]_ , \new_[67836]_ ,
    \new_[67840]_ , \new_[67841]_ , \new_[67844]_ , \new_[67847]_ ,
    \new_[67848]_ , \new_[67849]_ , \new_[67853]_ , \new_[67854]_ ,
    \new_[67857]_ , \new_[67860]_ , \new_[67861]_ , \new_[67862]_ ,
    \new_[67866]_ , \new_[67867]_ , \new_[67870]_ , \new_[67873]_ ,
    \new_[67874]_ , \new_[67875]_ , \new_[67879]_ , \new_[67880]_ ,
    \new_[67883]_ , \new_[67886]_ , \new_[67887]_ , \new_[67888]_ ,
    \new_[67892]_ , \new_[67893]_ , \new_[67896]_ , \new_[67899]_ ,
    \new_[67900]_ , \new_[67901]_ , \new_[67905]_ , \new_[67906]_ ,
    \new_[67909]_ , \new_[67912]_ , \new_[67913]_ , \new_[67914]_ ,
    \new_[67918]_ , \new_[67919]_ , \new_[67922]_ , \new_[67925]_ ,
    \new_[67926]_ , \new_[67927]_ , \new_[67931]_ , \new_[67932]_ ,
    \new_[67935]_ , \new_[67938]_ , \new_[67939]_ , \new_[67940]_ ,
    \new_[67944]_ , \new_[67945]_ , \new_[67948]_ , \new_[67951]_ ,
    \new_[67952]_ , \new_[67953]_ , \new_[67957]_ , \new_[67958]_ ,
    \new_[67961]_ , \new_[67964]_ , \new_[67965]_ , \new_[67966]_ ,
    \new_[67970]_ , \new_[67971]_ , \new_[67974]_ , \new_[67977]_ ,
    \new_[67978]_ , \new_[67979]_ , \new_[67983]_ , \new_[67984]_ ,
    \new_[67987]_ , \new_[67990]_ , \new_[67991]_ , \new_[67992]_ ,
    \new_[67996]_ , \new_[67997]_ , \new_[68000]_ , \new_[68003]_ ,
    \new_[68004]_ , \new_[68005]_ , \new_[68009]_ , \new_[68010]_ ,
    \new_[68013]_ , \new_[68016]_ , \new_[68017]_ , \new_[68018]_ ,
    \new_[68022]_ , \new_[68023]_ , \new_[68026]_ , \new_[68029]_ ,
    \new_[68030]_ , \new_[68031]_ , \new_[68035]_ , \new_[68036]_ ,
    \new_[68039]_ , \new_[68042]_ , \new_[68043]_ , \new_[68044]_ ,
    \new_[68048]_ , \new_[68049]_ , \new_[68052]_ , \new_[68055]_ ,
    \new_[68056]_ , \new_[68057]_ , \new_[68061]_ , \new_[68062]_ ,
    \new_[68065]_ , \new_[68068]_ , \new_[68069]_ , \new_[68070]_ ,
    \new_[68074]_ , \new_[68075]_ , \new_[68078]_ , \new_[68081]_ ,
    \new_[68082]_ , \new_[68083]_ , \new_[68087]_ , \new_[68088]_ ,
    \new_[68091]_ , \new_[68094]_ , \new_[68095]_ , \new_[68096]_ ,
    \new_[68100]_ , \new_[68101]_ , \new_[68104]_ , \new_[68107]_ ,
    \new_[68108]_ , \new_[68109]_ , \new_[68113]_ , \new_[68114]_ ,
    \new_[68117]_ , \new_[68120]_ , \new_[68121]_ , \new_[68122]_ ,
    \new_[68126]_ , \new_[68127]_ , \new_[68130]_ , \new_[68133]_ ,
    \new_[68134]_ , \new_[68135]_ , \new_[68139]_ , \new_[68140]_ ,
    \new_[68143]_ , \new_[68146]_ , \new_[68147]_ , \new_[68148]_ ,
    \new_[68152]_ , \new_[68153]_ , \new_[68156]_ , \new_[68159]_ ,
    \new_[68160]_ , \new_[68161]_ , \new_[68165]_ , \new_[68166]_ ,
    \new_[68169]_ , \new_[68172]_ , \new_[68173]_ , \new_[68174]_ ,
    \new_[68178]_ , \new_[68179]_ , \new_[68182]_ , \new_[68185]_ ,
    \new_[68186]_ , \new_[68187]_ , \new_[68191]_ , \new_[68192]_ ,
    \new_[68195]_ , \new_[68198]_ , \new_[68199]_ , \new_[68200]_ ,
    \new_[68204]_ , \new_[68205]_ , \new_[68208]_ , \new_[68211]_ ,
    \new_[68212]_ , \new_[68213]_ , \new_[68217]_ , \new_[68218]_ ,
    \new_[68221]_ , \new_[68224]_ , \new_[68225]_ , \new_[68226]_ ,
    \new_[68230]_ , \new_[68231]_ , \new_[68234]_ , \new_[68237]_ ,
    \new_[68238]_ , \new_[68239]_ , \new_[68243]_ , \new_[68244]_ ,
    \new_[68247]_ , \new_[68250]_ , \new_[68251]_ , \new_[68252]_ ,
    \new_[68256]_ , \new_[68257]_ , \new_[68260]_ , \new_[68263]_ ,
    \new_[68264]_ , \new_[68265]_ , \new_[68269]_ , \new_[68270]_ ,
    \new_[68273]_ , \new_[68276]_ , \new_[68277]_ , \new_[68278]_ ,
    \new_[68282]_ , \new_[68283]_ , \new_[68286]_ , \new_[68289]_ ,
    \new_[68290]_ , \new_[68291]_ , \new_[68295]_ , \new_[68296]_ ,
    \new_[68299]_ , \new_[68302]_ , \new_[68303]_ , \new_[68304]_ ,
    \new_[68308]_ , \new_[68309]_ , \new_[68312]_ , \new_[68315]_ ,
    \new_[68316]_ , \new_[68317]_ , \new_[68321]_ , \new_[68322]_ ,
    \new_[68325]_ , \new_[68328]_ , \new_[68329]_ , \new_[68330]_ ,
    \new_[68334]_ , \new_[68335]_ , \new_[68338]_ , \new_[68341]_ ,
    \new_[68342]_ , \new_[68343]_ , \new_[68347]_ , \new_[68348]_ ,
    \new_[68351]_ , \new_[68354]_ , \new_[68355]_ , \new_[68356]_ ,
    \new_[68360]_ , \new_[68361]_ , \new_[68364]_ , \new_[68367]_ ,
    \new_[68368]_ , \new_[68369]_ , \new_[68373]_ , \new_[68374]_ ,
    \new_[68377]_ , \new_[68380]_ , \new_[68381]_ , \new_[68382]_ ,
    \new_[68386]_ , \new_[68387]_ , \new_[68390]_ , \new_[68393]_ ,
    \new_[68394]_ , \new_[68395]_ , \new_[68399]_ , \new_[68400]_ ,
    \new_[68403]_ , \new_[68406]_ , \new_[68407]_ , \new_[68408]_ ,
    \new_[68412]_ , \new_[68413]_ , \new_[68416]_ , \new_[68419]_ ,
    \new_[68420]_ , \new_[68421]_ , \new_[68425]_ , \new_[68426]_ ,
    \new_[68429]_ , \new_[68432]_ , \new_[68433]_ , \new_[68434]_ ,
    \new_[68438]_ , \new_[68439]_ , \new_[68442]_ , \new_[68445]_ ,
    \new_[68446]_ , \new_[68447]_ , \new_[68451]_ , \new_[68452]_ ,
    \new_[68455]_ , \new_[68458]_ , \new_[68459]_ , \new_[68460]_ ,
    \new_[68464]_ , \new_[68465]_ , \new_[68468]_ , \new_[68471]_ ,
    \new_[68472]_ , \new_[68473]_ , \new_[68477]_ , \new_[68478]_ ,
    \new_[68481]_ , \new_[68484]_ , \new_[68485]_ , \new_[68486]_ ,
    \new_[68490]_ , \new_[68491]_ , \new_[68494]_ , \new_[68497]_ ,
    \new_[68498]_ , \new_[68499]_ , \new_[68503]_ , \new_[68504]_ ,
    \new_[68507]_ , \new_[68510]_ , \new_[68511]_ , \new_[68512]_ ,
    \new_[68516]_ , \new_[68517]_ , \new_[68520]_ , \new_[68523]_ ,
    \new_[68524]_ , \new_[68525]_ , \new_[68529]_ , \new_[68530]_ ,
    \new_[68533]_ , \new_[68536]_ , \new_[68537]_ , \new_[68538]_ ,
    \new_[68542]_ , \new_[68543]_ , \new_[68546]_ , \new_[68549]_ ,
    \new_[68550]_ , \new_[68551]_ , \new_[68555]_ , \new_[68556]_ ,
    \new_[68559]_ , \new_[68562]_ , \new_[68563]_ , \new_[68564]_ ,
    \new_[68568]_ , \new_[68569]_ , \new_[68572]_ , \new_[68575]_ ,
    \new_[68576]_ , \new_[68577]_ , \new_[68581]_ , \new_[68582]_ ,
    \new_[68585]_ , \new_[68588]_ , \new_[68589]_ , \new_[68590]_ ,
    \new_[68594]_ , \new_[68595]_ , \new_[68598]_ , \new_[68601]_ ,
    \new_[68602]_ , \new_[68603]_ , \new_[68607]_ , \new_[68608]_ ,
    \new_[68611]_ , \new_[68614]_ , \new_[68615]_ , \new_[68616]_ ,
    \new_[68620]_ , \new_[68621]_ , \new_[68624]_ , \new_[68627]_ ,
    \new_[68628]_ , \new_[68629]_ , \new_[68633]_ , \new_[68634]_ ,
    \new_[68637]_ , \new_[68640]_ , \new_[68641]_ , \new_[68642]_ ,
    \new_[68646]_ , \new_[68647]_ , \new_[68650]_ , \new_[68653]_ ,
    \new_[68654]_ , \new_[68655]_ , \new_[68659]_ , \new_[68660]_ ,
    \new_[68663]_ , \new_[68666]_ , \new_[68667]_ , \new_[68668]_ ,
    \new_[68672]_ , \new_[68673]_ , \new_[68676]_ , \new_[68679]_ ,
    \new_[68680]_ , \new_[68681]_ , \new_[68685]_ , \new_[68686]_ ,
    \new_[68689]_ , \new_[68692]_ , \new_[68693]_ , \new_[68694]_ ,
    \new_[68698]_ , \new_[68699]_ , \new_[68702]_ , \new_[68705]_ ,
    \new_[68706]_ , \new_[68707]_ , \new_[68711]_ , \new_[68712]_ ,
    \new_[68715]_ , \new_[68718]_ , \new_[68719]_ , \new_[68720]_ ,
    \new_[68724]_ , \new_[68725]_ , \new_[68728]_ , \new_[68731]_ ,
    \new_[68732]_ , \new_[68733]_ , \new_[68737]_ , \new_[68738]_ ,
    \new_[68741]_ , \new_[68744]_ , \new_[68745]_ , \new_[68746]_ ,
    \new_[68750]_ , \new_[68751]_ , \new_[68754]_ , \new_[68757]_ ,
    \new_[68758]_ , \new_[68759]_ , \new_[68763]_ , \new_[68764]_ ,
    \new_[68767]_ , \new_[68770]_ , \new_[68771]_ , \new_[68772]_ ,
    \new_[68776]_ , \new_[68777]_ , \new_[68780]_ , \new_[68783]_ ,
    \new_[68784]_ , \new_[68785]_ , \new_[68789]_ , \new_[68790]_ ,
    \new_[68793]_ , \new_[68796]_ , \new_[68797]_ , \new_[68798]_ ,
    \new_[68802]_ , \new_[68803]_ , \new_[68806]_ , \new_[68809]_ ,
    \new_[68810]_ , \new_[68811]_ , \new_[68815]_ , \new_[68816]_ ,
    \new_[68819]_ , \new_[68822]_ , \new_[68823]_ , \new_[68824]_ ,
    \new_[68828]_ , \new_[68829]_ , \new_[68832]_ , \new_[68835]_ ,
    \new_[68836]_ , \new_[68837]_ , \new_[68841]_ , \new_[68842]_ ,
    \new_[68845]_ , \new_[68848]_ , \new_[68849]_ , \new_[68850]_ ,
    \new_[68854]_ , \new_[68855]_ , \new_[68858]_ , \new_[68861]_ ,
    \new_[68862]_ , \new_[68863]_ , \new_[68867]_ , \new_[68868]_ ,
    \new_[68871]_ , \new_[68874]_ , \new_[68875]_ , \new_[68876]_ ,
    \new_[68880]_ , \new_[68881]_ , \new_[68884]_ , \new_[68887]_ ,
    \new_[68888]_ , \new_[68889]_ , \new_[68893]_ , \new_[68894]_ ,
    \new_[68897]_ , \new_[68900]_ , \new_[68901]_ , \new_[68902]_ ,
    \new_[68906]_ , \new_[68907]_ , \new_[68910]_ , \new_[68913]_ ,
    \new_[68914]_ , \new_[68915]_ , \new_[68919]_ , \new_[68920]_ ,
    \new_[68923]_ , \new_[68926]_ , \new_[68927]_ , \new_[68928]_ ,
    \new_[68932]_ , \new_[68933]_ , \new_[68936]_ , \new_[68939]_ ,
    \new_[68940]_ , \new_[68941]_ , \new_[68945]_ , \new_[68946]_ ,
    \new_[68949]_ , \new_[68952]_ , \new_[68953]_ , \new_[68954]_ ,
    \new_[68958]_ , \new_[68959]_ , \new_[68962]_ , \new_[68965]_ ,
    \new_[68966]_ , \new_[68967]_ , \new_[68971]_ , \new_[68972]_ ,
    \new_[68975]_ , \new_[68978]_ , \new_[68979]_ , \new_[68980]_ ,
    \new_[68984]_ , \new_[68985]_ , \new_[68988]_ , \new_[68991]_ ,
    \new_[68992]_ , \new_[68993]_ , \new_[68997]_ , \new_[68998]_ ,
    \new_[69001]_ , \new_[69004]_ , \new_[69005]_ , \new_[69006]_ ,
    \new_[69010]_ , \new_[69011]_ , \new_[69014]_ , \new_[69017]_ ,
    \new_[69018]_ , \new_[69019]_ , \new_[69023]_ , \new_[69024]_ ,
    \new_[69027]_ , \new_[69030]_ , \new_[69031]_ , \new_[69032]_ ,
    \new_[69036]_ , \new_[69037]_ , \new_[69040]_ , \new_[69043]_ ,
    \new_[69044]_ , \new_[69045]_ , \new_[69049]_ , \new_[69050]_ ,
    \new_[69053]_ , \new_[69056]_ , \new_[69057]_ , \new_[69058]_ ,
    \new_[69062]_ , \new_[69063]_ , \new_[69066]_ , \new_[69069]_ ,
    \new_[69070]_ , \new_[69071]_ , \new_[69075]_ , \new_[69076]_ ,
    \new_[69079]_ , \new_[69082]_ , \new_[69083]_ , \new_[69084]_ ,
    \new_[69088]_ , \new_[69089]_ , \new_[69092]_ , \new_[69095]_ ,
    \new_[69096]_ , \new_[69097]_ , \new_[69101]_ , \new_[69102]_ ,
    \new_[69105]_ , \new_[69108]_ , \new_[69109]_ , \new_[69110]_ ,
    \new_[69114]_ , \new_[69115]_ , \new_[69118]_ , \new_[69121]_ ,
    \new_[69122]_ , \new_[69123]_ , \new_[69127]_ , \new_[69128]_ ,
    \new_[69131]_ , \new_[69134]_ , \new_[69135]_ , \new_[69136]_ ,
    \new_[69140]_ , \new_[69141]_ , \new_[69144]_ , \new_[69147]_ ,
    \new_[69148]_ , \new_[69149]_ , \new_[69153]_ , \new_[69154]_ ,
    \new_[69157]_ , \new_[69160]_ , \new_[69161]_ , \new_[69162]_ ,
    \new_[69166]_ , \new_[69167]_ , \new_[69170]_ , \new_[69173]_ ,
    \new_[69174]_ , \new_[69175]_ , \new_[69179]_ , \new_[69180]_ ,
    \new_[69183]_ , \new_[69186]_ , \new_[69187]_ , \new_[69188]_ ,
    \new_[69192]_ , \new_[69193]_ , \new_[69196]_ , \new_[69199]_ ,
    \new_[69200]_ , \new_[69201]_ , \new_[69205]_ , \new_[69206]_ ,
    \new_[69209]_ , \new_[69212]_ , \new_[69213]_ , \new_[69214]_ ,
    \new_[69218]_ , \new_[69219]_ , \new_[69222]_ , \new_[69225]_ ,
    \new_[69226]_ , \new_[69227]_ , \new_[69231]_ , \new_[69232]_ ,
    \new_[69235]_ , \new_[69238]_ , \new_[69239]_ , \new_[69240]_ ,
    \new_[69244]_ , \new_[69245]_ , \new_[69248]_ , \new_[69251]_ ,
    \new_[69252]_ , \new_[69253]_ , \new_[69257]_ , \new_[69258]_ ,
    \new_[69261]_ , \new_[69264]_ , \new_[69265]_ , \new_[69266]_ ,
    \new_[69270]_ , \new_[69271]_ , \new_[69274]_ , \new_[69277]_ ,
    \new_[69278]_ , \new_[69279]_ , \new_[69283]_ , \new_[69284]_ ,
    \new_[69287]_ , \new_[69290]_ , \new_[69291]_ , \new_[69292]_ ,
    \new_[69296]_ , \new_[69297]_ , \new_[69300]_ , \new_[69303]_ ,
    \new_[69304]_ , \new_[69305]_ , \new_[69309]_ , \new_[69310]_ ,
    \new_[69313]_ , \new_[69316]_ , \new_[69317]_ , \new_[69318]_ ,
    \new_[69322]_ , \new_[69323]_ , \new_[69326]_ , \new_[69329]_ ,
    \new_[69330]_ , \new_[69331]_ , \new_[69335]_ , \new_[69336]_ ,
    \new_[69339]_ , \new_[69342]_ , \new_[69343]_ , \new_[69344]_ ,
    \new_[69348]_ , \new_[69349]_ , \new_[69352]_ , \new_[69355]_ ,
    \new_[69356]_ , \new_[69357]_ , \new_[69361]_ , \new_[69362]_ ,
    \new_[69365]_ , \new_[69368]_ , \new_[69369]_ , \new_[69370]_ ,
    \new_[69374]_ , \new_[69375]_ , \new_[69378]_ , \new_[69381]_ ,
    \new_[69382]_ , \new_[69383]_ , \new_[69387]_ , \new_[69388]_ ,
    \new_[69391]_ , \new_[69394]_ , \new_[69395]_ , \new_[69396]_ ,
    \new_[69400]_ , \new_[69401]_ , \new_[69404]_ , \new_[69407]_ ,
    \new_[69408]_ , \new_[69409]_ , \new_[69413]_ , \new_[69414]_ ,
    \new_[69417]_ , \new_[69420]_ , \new_[69421]_ , \new_[69422]_ ,
    \new_[69426]_ , \new_[69427]_ , \new_[69430]_ , \new_[69433]_ ,
    \new_[69434]_ , \new_[69435]_ , \new_[69439]_ , \new_[69440]_ ,
    \new_[69443]_ , \new_[69446]_ , \new_[69447]_ , \new_[69448]_ ,
    \new_[69452]_ , \new_[69453]_ , \new_[69456]_ , \new_[69459]_ ,
    \new_[69460]_ , \new_[69461]_ , \new_[69465]_ , \new_[69466]_ ,
    \new_[69469]_ , \new_[69472]_ , \new_[69473]_ , \new_[69474]_ ,
    \new_[69478]_ , \new_[69479]_ , \new_[69482]_ , \new_[69485]_ ,
    \new_[69486]_ , \new_[69487]_ , \new_[69491]_ , \new_[69492]_ ,
    \new_[69495]_ , \new_[69498]_ , \new_[69499]_ , \new_[69500]_ ,
    \new_[69504]_ , \new_[69505]_ , \new_[69508]_ , \new_[69511]_ ,
    \new_[69512]_ , \new_[69513]_ , \new_[69517]_ , \new_[69518]_ ,
    \new_[69521]_ , \new_[69524]_ , \new_[69525]_ , \new_[69526]_ ,
    \new_[69530]_ , \new_[69531]_ , \new_[69534]_ , \new_[69537]_ ,
    \new_[69538]_ , \new_[69539]_ , \new_[69543]_ , \new_[69544]_ ,
    \new_[69547]_ , \new_[69550]_ , \new_[69551]_ , \new_[69552]_ ,
    \new_[69556]_ , \new_[69557]_ , \new_[69560]_ , \new_[69563]_ ,
    \new_[69564]_ , \new_[69565]_ , \new_[69569]_ , \new_[69570]_ ,
    \new_[69573]_ , \new_[69576]_ , \new_[69577]_ , \new_[69578]_ ,
    \new_[69582]_ , \new_[69583]_ , \new_[69586]_ , \new_[69589]_ ,
    \new_[69590]_ , \new_[69591]_ , \new_[69595]_ , \new_[69596]_ ,
    \new_[69599]_ , \new_[69602]_ , \new_[69603]_ , \new_[69604]_ ,
    \new_[69608]_ , \new_[69609]_ , \new_[69612]_ , \new_[69615]_ ,
    \new_[69616]_ , \new_[69617]_ , \new_[69621]_ , \new_[69622]_ ,
    \new_[69625]_ , \new_[69628]_ , \new_[69629]_ , \new_[69630]_ ,
    \new_[69634]_ , \new_[69635]_ , \new_[69638]_ , \new_[69641]_ ,
    \new_[69642]_ , \new_[69643]_ , \new_[69647]_ , \new_[69648]_ ,
    \new_[69651]_ , \new_[69654]_ , \new_[69655]_ , \new_[69656]_ ,
    \new_[69660]_ , \new_[69661]_ , \new_[69664]_ , \new_[69667]_ ,
    \new_[69668]_ , \new_[69669]_ , \new_[69673]_ , \new_[69674]_ ,
    \new_[69677]_ , \new_[69680]_ , \new_[69681]_ , \new_[69682]_ ,
    \new_[69686]_ , \new_[69687]_ , \new_[69690]_ , \new_[69693]_ ,
    \new_[69694]_ , \new_[69695]_ , \new_[69699]_ , \new_[69700]_ ,
    \new_[69703]_ , \new_[69706]_ , \new_[69707]_ , \new_[69708]_ ,
    \new_[69712]_ , \new_[69713]_ , \new_[69716]_ , \new_[69719]_ ,
    \new_[69720]_ , \new_[69721]_ , \new_[69725]_ , \new_[69726]_ ,
    \new_[69729]_ , \new_[69732]_ , \new_[69733]_ , \new_[69734]_ ,
    \new_[69738]_ , \new_[69739]_ , \new_[69742]_ , \new_[69745]_ ,
    \new_[69746]_ , \new_[69747]_ , \new_[69751]_ , \new_[69752]_ ,
    \new_[69755]_ , \new_[69758]_ , \new_[69759]_ , \new_[69760]_ ,
    \new_[69764]_ , \new_[69765]_ , \new_[69768]_ , \new_[69771]_ ,
    \new_[69772]_ , \new_[69773]_ , \new_[69777]_ , \new_[69778]_ ,
    \new_[69781]_ , \new_[69784]_ , \new_[69785]_ , \new_[69786]_ ,
    \new_[69790]_ , \new_[69791]_ , \new_[69794]_ , \new_[69797]_ ,
    \new_[69798]_ , \new_[69799]_ , \new_[69803]_ , \new_[69804]_ ,
    \new_[69807]_ , \new_[69810]_ , \new_[69811]_ , \new_[69812]_ ,
    \new_[69816]_ , \new_[69817]_ , \new_[69820]_ , \new_[69823]_ ,
    \new_[69824]_ , \new_[69825]_ , \new_[69829]_ , \new_[69830]_ ,
    \new_[69833]_ , \new_[69836]_ , \new_[69837]_ , \new_[69838]_ ,
    \new_[69842]_ , \new_[69843]_ , \new_[69846]_ , \new_[69849]_ ,
    \new_[69850]_ , \new_[69851]_ , \new_[69855]_ , \new_[69856]_ ,
    \new_[69859]_ , \new_[69862]_ , \new_[69863]_ , \new_[69864]_ ,
    \new_[69868]_ , \new_[69869]_ , \new_[69872]_ , \new_[69875]_ ,
    \new_[69876]_ , \new_[69877]_ , \new_[69881]_ , \new_[69882]_ ,
    \new_[69885]_ , \new_[69888]_ , \new_[69889]_ , \new_[69890]_ ,
    \new_[69894]_ , \new_[69895]_ , \new_[69898]_ , \new_[69901]_ ,
    \new_[69902]_ , \new_[69903]_ , \new_[69907]_ , \new_[69908]_ ,
    \new_[69911]_ , \new_[69914]_ , \new_[69915]_ , \new_[69916]_ ,
    \new_[69920]_ , \new_[69921]_ , \new_[69924]_ , \new_[69927]_ ,
    \new_[69928]_ , \new_[69929]_ , \new_[69933]_ , \new_[69934]_ ,
    \new_[69937]_ , \new_[69940]_ , \new_[69941]_ , \new_[69942]_ ,
    \new_[69946]_ , \new_[69947]_ , \new_[69950]_ , \new_[69953]_ ,
    \new_[69954]_ , \new_[69955]_ , \new_[69959]_ , \new_[69960]_ ,
    \new_[69963]_ , \new_[69966]_ , \new_[69967]_ , \new_[69968]_ ,
    \new_[69972]_ , \new_[69973]_ , \new_[69976]_ , \new_[69979]_ ,
    \new_[69980]_ , \new_[69981]_ , \new_[69985]_ , \new_[69986]_ ,
    \new_[69989]_ , \new_[69992]_ , \new_[69993]_ , \new_[69994]_ ,
    \new_[69998]_ , \new_[69999]_ , \new_[70002]_ , \new_[70005]_ ,
    \new_[70006]_ , \new_[70007]_ , \new_[70011]_ , \new_[70012]_ ,
    \new_[70015]_ , \new_[70018]_ , \new_[70019]_ , \new_[70020]_ ,
    \new_[70024]_ , \new_[70025]_ , \new_[70028]_ , \new_[70031]_ ,
    \new_[70032]_ , \new_[70033]_ , \new_[70037]_ , \new_[70038]_ ,
    \new_[70041]_ , \new_[70044]_ , \new_[70045]_ , \new_[70046]_ ,
    \new_[70050]_ , \new_[70051]_ , \new_[70054]_ , \new_[70057]_ ,
    \new_[70058]_ , \new_[70059]_ , \new_[70063]_ , \new_[70064]_ ,
    \new_[70067]_ , \new_[70070]_ , \new_[70071]_ , \new_[70072]_ ,
    \new_[70076]_ , \new_[70077]_ , \new_[70080]_ , \new_[70083]_ ,
    \new_[70084]_ , \new_[70085]_ , \new_[70089]_ , \new_[70090]_ ,
    \new_[70093]_ , \new_[70096]_ , \new_[70097]_ , \new_[70098]_ ,
    \new_[70102]_ , \new_[70103]_ , \new_[70106]_ , \new_[70109]_ ,
    \new_[70110]_ , \new_[70111]_ , \new_[70115]_ , \new_[70116]_ ,
    \new_[70119]_ , \new_[70122]_ , \new_[70123]_ , \new_[70124]_ ,
    \new_[70128]_ , \new_[70129]_ , \new_[70132]_ , \new_[70135]_ ,
    \new_[70136]_ , \new_[70137]_ , \new_[70141]_ , \new_[70142]_ ,
    \new_[70145]_ , \new_[70148]_ , \new_[70149]_ , \new_[70150]_ ,
    \new_[70154]_ , \new_[70155]_ , \new_[70158]_ , \new_[70161]_ ,
    \new_[70162]_ , \new_[70163]_ , \new_[70167]_ , \new_[70168]_ ,
    \new_[70171]_ , \new_[70174]_ , \new_[70175]_ , \new_[70176]_ ,
    \new_[70180]_ , \new_[70181]_ , \new_[70184]_ , \new_[70187]_ ,
    \new_[70188]_ , \new_[70189]_ , \new_[70193]_ , \new_[70194]_ ,
    \new_[70197]_ , \new_[70200]_ , \new_[70201]_ , \new_[70202]_ ,
    \new_[70206]_ , \new_[70207]_ , \new_[70210]_ , \new_[70213]_ ,
    \new_[70214]_ , \new_[70215]_ , \new_[70219]_ , \new_[70220]_ ,
    \new_[70223]_ , \new_[70226]_ , \new_[70227]_ , \new_[70228]_ ,
    \new_[70232]_ , \new_[70233]_ , \new_[70236]_ , \new_[70239]_ ,
    \new_[70240]_ , \new_[70241]_ , \new_[70245]_ , \new_[70246]_ ,
    \new_[70249]_ , \new_[70252]_ , \new_[70253]_ , \new_[70254]_ ,
    \new_[70258]_ , \new_[70259]_ , \new_[70262]_ , \new_[70265]_ ,
    \new_[70266]_ , \new_[70267]_ , \new_[70271]_ , \new_[70272]_ ,
    \new_[70275]_ , \new_[70278]_ , \new_[70279]_ , \new_[70280]_ ,
    \new_[70284]_ , \new_[70285]_ , \new_[70288]_ , \new_[70291]_ ,
    \new_[70292]_ , \new_[70293]_ , \new_[70297]_ , \new_[70298]_ ,
    \new_[70301]_ , \new_[70304]_ , \new_[70305]_ , \new_[70306]_ ,
    \new_[70310]_ , \new_[70311]_ , \new_[70314]_ , \new_[70317]_ ,
    \new_[70318]_ , \new_[70319]_ , \new_[70323]_ , \new_[70324]_ ,
    \new_[70327]_ , \new_[70330]_ , \new_[70331]_ , \new_[70332]_ ,
    \new_[70336]_ , \new_[70337]_ , \new_[70340]_ , \new_[70343]_ ,
    \new_[70344]_ , \new_[70345]_ , \new_[70349]_ , \new_[70350]_ ,
    \new_[70353]_ , \new_[70356]_ , \new_[70357]_ , \new_[70358]_ ,
    \new_[70362]_ , \new_[70363]_ , \new_[70366]_ , \new_[70369]_ ,
    \new_[70370]_ , \new_[70371]_ , \new_[70375]_ , \new_[70376]_ ,
    \new_[70379]_ , \new_[70382]_ , \new_[70383]_ , \new_[70384]_ ,
    \new_[70388]_ , \new_[70389]_ , \new_[70392]_ , \new_[70395]_ ,
    \new_[70396]_ , \new_[70397]_ , \new_[70401]_ , \new_[70402]_ ,
    \new_[70405]_ , \new_[70408]_ , \new_[70409]_ , \new_[70410]_ ,
    \new_[70414]_ , \new_[70415]_ , \new_[70418]_ , \new_[70421]_ ,
    \new_[70422]_ , \new_[70423]_ , \new_[70427]_ , \new_[70428]_ ,
    \new_[70431]_ , \new_[70434]_ , \new_[70435]_ , \new_[70436]_ ,
    \new_[70440]_ , \new_[70441]_ , \new_[70444]_ , \new_[70447]_ ,
    \new_[70448]_ , \new_[70449]_ , \new_[70453]_ , \new_[70454]_ ,
    \new_[70457]_ , \new_[70460]_ , \new_[70461]_ , \new_[70462]_ ,
    \new_[70466]_ , \new_[70467]_ , \new_[70470]_ , \new_[70473]_ ,
    \new_[70474]_ , \new_[70475]_ , \new_[70479]_ , \new_[70480]_ ,
    \new_[70483]_ , \new_[70486]_ , \new_[70487]_ , \new_[70488]_ ,
    \new_[70492]_ , \new_[70493]_ , \new_[70496]_ , \new_[70499]_ ,
    \new_[70500]_ , \new_[70501]_ , \new_[70505]_ , \new_[70506]_ ,
    \new_[70509]_ , \new_[70512]_ , \new_[70513]_ , \new_[70514]_ ,
    \new_[70518]_ , \new_[70519]_ , \new_[70522]_ , \new_[70525]_ ,
    \new_[70526]_ , \new_[70527]_ , \new_[70531]_ , \new_[70532]_ ,
    \new_[70535]_ , \new_[70538]_ , \new_[70539]_ , \new_[70540]_ ,
    \new_[70544]_ , \new_[70545]_ , \new_[70548]_ , \new_[70551]_ ,
    \new_[70552]_ , \new_[70553]_ , \new_[70557]_ , \new_[70558]_ ,
    \new_[70561]_ , \new_[70564]_ , \new_[70565]_ , \new_[70566]_ ,
    \new_[70570]_ , \new_[70571]_ , \new_[70574]_ , \new_[70577]_ ,
    \new_[70578]_ , \new_[70579]_ , \new_[70583]_ , \new_[70584]_ ,
    \new_[70587]_ , \new_[70590]_ , \new_[70591]_ , \new_[70592]_ ,
    \new_[70596]_ , \new_[70597]_ , \new_[70600]_ , \new_[70603]_ ,
    \new_[70604]_ , \new_[70605]_ , \new_[70609]_ , \new_[70610]_ ,
    \new_[70613]_ , \new_[70616]_ , \new_[70617]_ , \new_[70618]_ ,
    \new_[70622]_ , \new_[70623]_ , \new_[70626]_ , \new_[70629]_ ,
    \new_[70630]_ , \new_[70631]_ , \new_[70635]_ , \new_[70636]_ ,
    \new_[70639]_ , \new_[70642]_ , \new_[70643]_ , \new_[70644]_ ,
    \new_[70648]_ , \new_[70649]_ , \new_[70652]_ , \new_[70655]_ ,
    \new_[70656]_ , \new_[70657]_ , \new_[70661]_ , \new_[70662]_ ,
    \new_[70665]_ , \new_[70668]_ , \new_[70669]_ , \new_[70670]_ ,
    \new_[70674]_ , \new_[70675]_ , \new_[70678]_ , \new_[70681]_ ,
    \new_[70682]_ , \new_[70683]_ , \new_[70687]_ , \new_[70688]_ ,
    \new_[70691]_ , \new_[70694]_ , \new_[70695]_ , \new_[70696]_ ,
    \new_[70700]_ , \new_[70701]_ , \new_[70704]_ , \new_[70707]_ ,
    \new_[70708]_ , \new_[70709]_ , \new_[70713]_ , \new_[70714]_ ,
    \new_[70717]_ , \new_[70720]_ , \new_[70721]_ , \new_[70722]_ ,
    \new_[70726]_ , \new_[70727]_ , \new_[70730]_ , \new_[70733]_ ,
    \new_[70734]_ , \new_[70735]_ , \new_[70739]_ , \new_[70740]_ ,
    \new_[70743]_ , \new_[70746]_ , \new_[70747]_ , \new_[70748]_ ,
    \new_[70752]_ , \new_[70753]_ , \new_[70756]_ , \new_[70759]_ ,
    \new_[70760]_ , \new_[70761]_ , \new_[70765]_ , \new_[70766]_ ,
    \new_[70769]_ , \new_[70772]_ , \new_[70773]_ , \new_[70774]_ ,
    \new_[70778]_ , \new_[70779]_ , \new_[70782]_ , \new_[70785]_ ,
    \new_[70786]_ , \new_[70787]_ , \new_[70791]_ , \new_[70792]_ ,
    \new_[70795]_ , \new_[70798]_ , \new_[70799]_ , \new_[70800]_ ,
    \new_[70804]_ , \new_[70805]_ , \new_[70808]_ , \new_[70811]_ ,
    \new_[70812]_ , \new_[70813]_ , \new_[70817]_ , \new_[70818]_ ,
    \new_[70821]_ , \new_[70824]_ , \new_[70825]_ , \new_[70826]_ ,
    \new_[70830]_ , \new_[70831]_ , \new_[70834]_ , \new_[70837]_ ,
    \new_[70838]_ , \new_[70839]_ , \new_[70843]_ , \new_[70844]_ ,
    \new_[70847]_ , \new_[70850]_ , \new_[70851]_ , \new_[70852]_ ,
    \new_[70856]_ , \new_[70857]_ , \new_[70860]_ , \new_[70863]_ ,
    \new_[70864]_ , \new_[70865]_ , \new_[70869]_ , \new_[70870]_ ,
    \new_[70873]_ , \new_[70876]_ , \new_[70877]_ , \new_[70878]_ ,
    \new_[70882]_ , \new_[70883]_ , \new_[70886]_ , \new_[70889]_ ,
    \new_[70890]_ , \new_[70891]_ , \new_[70895]_ , \new_[70896]_ ,
    \new_[70899]_ , \new_[70902]_ , \new_[70903]_ , \new_[70904]_ ,
    \new_[70908]_ , \new_[70909]_ , \new_[70912]_ , \new_[70915]_ ,
    \new_[70916]_ , \new_[70917]_ , \new_[70921]_ , \new_[70922]_ ,
    \new_[70925]_ , \new_[70928]_ , \new_[70929]_ , \new_[70930]_ ,
    \new_[70934]_ , \new_[70935]_ , \new_[70938]_ , \new_[70941]_ ,
    \new_[70942]_ , \new_[70943]_ , \new_[70947]_ , \new_[70948]_ ,
    \new_[70951]_ , \new_[70954]_ , \new_[70955]_ , \new_[70956]_ ,
    \new_[70960]_ , \new_[70961]_ , \new_[70964]_ , \new_[70967]_ ,
    \new_[70968]_ , \new_[70969]_ , \new_[70973]_ , \new_[70974]_ ,
    \new_[70977]_ , \new_[70980]_ , \new_[70981]_ , \new_[70982]_ ,
    \new_[70986]_ , \new_[70987]_ , \new_[70990]_ , \new_[70993]_ ,
    \new_[70994]_ , \new_[70995]_ , \new_[70999]_ , \new_[71000]_ ,
    \new_[71003]_ , \new_[71006]_ , \new_[71007]_ , \new_[71008]_ ,
    \new_[71012]_ , \new_[71013]_ , \new_[71016]_ , \new_[71019]_ ,
    \new_[71020]_ , \new_[71021]_ , \new_[71025]_ , \new_[71026]_ ,
    \new_[71029]_ , \new_[71032]_ , \new_[71033]_ , \new_[71034]_ ,
    \new_[71038]_ , \new_[71039]_ , \new_[71042]_ , \new_[71045]_ ,
    \new_[71046]_ , \new_[71047]_ , \new_[71051]_ , \new_[71052]_ ,
    \new_[71055]_ , \new_[71058]_ , \new_[71059]_ , \new_[71060]_ ,
    \new_[71064]_ , \new_[71065]_ , \new_[71068]_ , \new_[71071]_ ,
    \new_[71072]_ , \new_[71073]_ , \new_[71077]_ , \new_[71078]_ ,
    \new_[71081]_ , \new_[71084]_ , \new_[71085]_ , \new_[71086]_ ,
    \new_[71090]_ , \new_[71091]_ , \new_[71094]_ , \new_[71097]_ ,
    \new_[71098]_ , \new_[71099]_ , \new_[71103]_ , \new_[71104]_ ,
    \new_[71107]_ , \new_[71110]_ , \new_[71111]_ , \new_[71112]_ ,
    \new_[71116]_ , \new_[71117]_ , \new_[71120]_ , \new_[71123]_ ,
    \new_[71124]_ , \new_[71125]_ , \new_[71129]_ , \new_[71130]_ ,
    \new_[71133]_ , \new_[71136]_ , \new_[71137]_ , \new_[71138]_ ,
    \new_[71142]_ , \new_[71143]_ , \new_[71146]_ , \new_[71149]_ ,
    \new_[71150]_ , \new_[71151]_ , \new_[71155]_ , \new_[71156]_ ,
    \new_[71159]_ , \new_[71162]_ , \new_[71163]_ , \new_[71164]_ ,
    \new_[71168]_ , \new_[71169]_ , \new_[71172]_ , \new_[71175]_ ,
    \new_[71176]_ , \new_[71177]_ , \new_[71181]_ , \new_[71182]_ ,
    \new_[71185]_ , \new_[71188]_ , \new_[71189]_ , \new_[71190]_ ,
    \new_[71194]_ , \new_[71195]_ , \new_[71198]_ , \new_[71201]_ ,
    \new_[71202]_ , \new_[71203]_ , \new_[71207]_ , \new_[71208]_ ,
    \new_[71211]_ , \new_[71214]_ , \new_[71215]_ , \new_[71216]_ ,
    \new_[71220]_ , \new_[71221]_ , \new_[71224]_ , \new_[71227]_ ,
    \new_[71228]_ , \new_[71229]_ , \new_[71233]_ , \new_[71234]_ ,
    \new_[71237]_ , \new_[71240]_ , \new_[71241]_ , \new_[71242]_ ,
    \new_[71246]_ , \new_[71247]_ , \new_[71250]_ , \new_[71253]_ ,
    \new_[71254]_ , \new_[71255]_ , \new_[71259]_ , \new_[71260]_ ,
    \new_[71263]_ , \new_[71266]_ , \new_[71267]_ , \new_[71268]_ ,
    \new_[71272]_ , \new_[71273]_ , \new_[71276]_ , \new_[71279]_ ,
    \new_[71280]_ , \new_[71281]_ , \new_[71285]_ , \new_[71286]_ ,
    \new_[71289]_ , \new_[71292]_ , \new_[71293]_ , \new_[71294]_ ,
    \new_[71298]_ , \new_[71299]_ , \new_[71302]_ , \new_[71305]_ ,
    \new_[71306]_ , \new_[71307]_ , \new_[71311]_ , \new_[71312]_ ,
    \new_[71315]_ , \new_[71318]_ , \new_[71319]_ , \new_[71320]_ ,
    \new_[71324]_ , \new_[71325]_ , \new_[71328]_ , \new_[71331]_ ,
    \new_[71332]_ , \new_[71333]_ , \new_[71337]_ , \new_[71338]_ ,
    \new_[71341]_ , \new_[71344]_ , \new_[71345]_ , \new_[71346]_ ,
    \new_[71350]_ , \new_[71351]_ , \new_[71354]_ , \new_[71357]_ ,
    \new_[71358]_ , \new_[71359]_ , \new_[71363]_ , \new_[71364]_ ,
    \new_[71367]_ , \new_[71370]_ , \new_[71371]_ , \new_[71372]_ ,
    \new_[71376]_ , \new_[71377]_ , \new_[71380]_ , \new_[71383]_ ,
    \new_[71384]_ , \new_[71385]_ , \new_[71389]_ , \new_[71390]_ ,
    \new_[71393]_ , \new_[71396]_ , \new_[71397]_ , \new_[71398]_ ,
    \new_[71402]_ , \new_[71403]_ , \new_[71406]_ , \new_[71409]_ ,
    \new_[71410]_ , \new_[71411]_ , \new_[71415]_ , \new_[71416]_ ,
    \new_[71419]_ , \new_[71422]_ , \new_[71423]_ , \new_[71424]_ ,
    \new_[71428]_ , \new_[71429]_ , \new_[71432]_ , \new_[71435]_ ,
    \new_[71436]_ , \new_[71437]_ , \new_[71441]_ , \new_[71442]_ ,
    \new_[71445]_ , \new_[71448]_ , \new_[71449]_ , \new_[71450]_ ,
    \new_[71454]_ , \new_[71455]_ , \new_[71458]_ , \new_[71461]_ ,
    \new_[71462]_ , \new_[71463]_ , \new_[71467]_ , \new_[71468]_ ,
    \new_[71471]_ , \new_[71474]_ , \new_[71475]_ , \new_[71476]_ ,
    \new_[71480]_ , \new_[71481]_ , \new_[71484]_ , \new_[71487]_ ,
    \new_[71488]_ , \new_[71489]_ , \new_[71493]_ , \new_[71494]_ ,
    \new_[71497]_ , \new_[71500]_ , \new_[71501]_ , \new_[71502]_ ,
    \new_[71506]_ , \new_[71507]_ , \new_[71510]_ , \new_[71513]_ ,
    \new_[71514]_ , \new_[71515]_ , \new_[71519]_ , \new_[71520]_ ,
    \new_[71523]_ , \new_[71526]_ , \new_[71527]_ , \new_[71528]_ ,
    \new_[71532]_ , \new_[71533]_ , \new_[71536]_ , \new_[71539]_ ,
    \new_[71540]_ , \new_[71541]_ , \new_[71545]_ , \new_[71546]_ ,
    \new_[71549]_ , \new_[71552]_ , \new_[71553]_ , \new_[71554]_ ,
    \new_[71558]_ , \new_[71559]_ , \new_[71562]_ , \new_[71565]_ ,
    \new_[71566]_ , \new_[71567]_ , \new_[71571]_ , \new_[71572]_ ,
    \new_[71575]_ , \new_[71578]_ , \new_[71579]_ , \new_[71580]_ ,
    \new_[71584]_ , \new_[71585]_ , \new_[71588]_ , \new_[71591]_ ,
    \new_[71592]_ , \new_[71593]_ , \new_[71597]_ , \new_[71598]_ ,
    \new_[71601]_ , \new_[71604]_ , \new_[71605]_ , \new_[71606]_ ,
    \new_[71610]_ , \new_[71611]_ , \new_[71614]_ , \new_[71617]_ ,
    \new_[71618]_ , \new_[71619]_ , \new_[71623]_ , \new_[71624]_ ,
    \new_[71627]_ , \new_[71630]_ , \new_[71631]_ , \new_[71632]_ ,
    \new_[71636]_ , \new_[71637]_ , \new_[71640]_ , \new_[71643]_ ,
    \new_[71644]_ , \new_[71645]_ , \new_[71649]_ , \new_[71650]_ ,
    \new_[71653]_ , \new_[71656]_ , \new_[71657]_ , \new_[71658]_ ,
    \new_[71662]_ , \new_[71663]_ , \new_[71666]_ , \new_[71669]_ ,
    \new_[71670]_ , \new_[71671]_ , \new_[71675]_ , \new_[71676]_ ,
    \new_[71679]_ , \new_[71682]_ , \new_[71683]_ , \new_[71684]_ ,
    \new_[71688]_ , \new_[71689]_ , \new_[71692]_ , \new_[71695]_ ,
    \new_[71696]_ , \new_[71697]_ , \new_[71701]_ , \new_[71702]_ ,
    \new_[71705]_ , \new_[71708]_ , \new_[71709]_ , \new_[71710]_ ,
    \new_[71714]_ , \new_[71715]_ , \new_[71718]_ , \new_[71721]_ ,
    \new_[71722]_ , \new_[71723]_ , \new_[71727]_ , \new_[71728]_ ,
    \new_[71731]_ , \new_[71734]_ , \new_[71735]_ , \new_[71736]_ ,
    \new_[71740]_ , \new_[71741]_ , \new_[71744]_ , \new_[71747]_ ,
    \new_[71748]_ , \new_[71749]_ , \new_[71753]_ , \new_[71754]_ ,
    \new_[71757]_ , \new_[71760]_ , \new_[71761]_ , \new_[71762]_ ,
    \new_[71766]_ , \new_[71767]_ , \new_[71770]_ , \new_[71773]_ ,
    \new_[71774]_ , \new_[71775]_ , \new_[71779]_ , \new_[71780]_ ,
    \new_[71783]_ , \new_[71786]_ , \new_[71787]_ , \new_[71788]_ ,
    \new_[71792]_ , \new_[71793]_ , \new_[71796]_ , \new_[71799]_ ,
    \new_[71800]_ , \new_[71801]_ , \new_[71805]_ , \new_[71806]_ ,
    \new_[71809]_ , \new_[71812]_ , \new_[71813]_ , \new_[71814]_ ,
    \new_[71818]_ , \new_[71819]_ , \new_[71822]_ , \new_[71825]_ ,
    \new_[71826]_ , \new_[71827]_ , \new_[71831]_ , \new_[71832]_ ,
    \new_[71835]_ , \new_[71838]_ , \new_[71839]_ , \new_[71840]_ ,
    \new_[71844]_ , \new_[71845]_ , \new_[71848]_ , \new_[71851]_ ,
    \new_[71852]_ , \new_[71853]_ , \new_[71857]_ , \new_[71858]_ ,
    \new_[71861]_ , \new_[71864]_ , \new_[71865]_ , \new_[71866]_ ,
    \new_[71870]_ , \new_[71871]_ , \new_[71874]_ , \new_[71877]_ ,
    \new_[71878]_ , \new_[71879]_ , \new_[71883]_ , \new_[71884]_ ,
    \new_[71887]_ , \new_[71890]_ , \new_[71891]_ , \new_[71892]_ ,
    \new_[71896]_ , \new_[71897]_ , \new_[71900]_ , \new_[71903]_ ,
    \new_[71904]_ , \new_[71905]_ , \new_[71909]_ , \new_[71910]_ ,
    \new_[71913]_ , \new_[71916]_ , \new_[71917]_ , \new_[71918]_ ,
    \new_[71922]_ , \new_[71923]_ , \new_[71926]_ , \new_[71929]_ ,
    \new_[71930]_ , \new_[71931]_ , \new_[71935]_ , \new_[71936]_ ,
    \new_[71939]_ , \new_[71942]_ , \new_[71943]_ , \new_[71944]_ ,
    \new_[71948]_ , \new_[71949]_ , \new_[71952]_ , \new_[71955]_ ,
    \new_[71956]_ , \new_[71957]_ , \new_[71961]_ , \new_[71962]_ ,
    \new_[71965]_ , \new_[71968]_ , \new_[71969]_ , \new_[71970]_ ,
    \new_[71974]_ , \new_[71975]_ , \new_[71978]_ , \new_[71981]_ ,
    \new_[71982]_ , \new_[71983]_ , \new_[71987]_ , \new_[71988]_ ,
    \new_[71991]_ , \new_[71994]_ , \new_[71995]_ , \new_[71996]_ ,
    \new_[72000]_ , \new_[72001]_ , \new_[72004]_ , \new_[72007]_ ,
    \new_[72008]_ , \new_[72009]_ , \new_[72013]_ , \new_[72014]_ ,
    \new_[72017]_ , \new_[72020]_ , \new_[72021]_ , \new_[72022]_ ,
    \new_[72026]_ , \new_[72027]_ , \new_[72030]_ , \new_[72033]_ ,
    \new_[72034]_ , \new_[72035]_ , \new_[72039]_ , \new_[72040]_ ,
    \new_[72043]_ , \new_[72046]_ , \new_[72047]_ , \new_[72048]_ ,
    \new_[72052]_ , \new_[72053]_ , \new_[72056]_ , \new_[72059]_ ,
    \new_[72060]_ , \new_[72061]_ , \new_[72065]_ , \new_[72066]_ ,
    \new_[72069]_ , \new_[72072]_ , \new_[72073]_ , \new_[72074]_ ,
    \new_[72078]_ , \new_[72079]_ , \new_[72082]_ , \new_[72085]_ ,
    \new_[72086]_ , \new_[72087]_ , \new_[72091]_ , \new_[72092]_ ,
    \new_[72095]_ , \new_[72098]_ , \new_[72099]_ , \new_[72100]_ ,
    \new_[72104]_ , \new_[72105]_ , \new_[72108]_ , \new_[72111]_ ,
    \new_[72112]_ , \new_[72113]_ , \new_[72117]_ , \new_[72118]_ ,
    \new_[72121]_ , \new_[72124]_ , \new_[72125]_ , \new_[72126]_ ,
    \new_[72130]_ , \new_[72131]_ , \new_[72134]_ , \new_[72137]_ ,
    \new_[72138]_ , \new_[72139]_ , \new_[72143]_ , \new_[72144]_ ,
    \new_[72147]_ , \new_[72150]_ , \new_[72151]_ , \new_[72152]_ ,
    \new_[72156]_ , \new_[72157]_ , \new_[72160]_ , \new_[72163]_ ,
    \new_[72164]_ , \new_[72165]_ , \new_[72169]_ , \new_[72170]_ ,
    \new_[72173]_ , \new_[72176]_ , \new_[72177]_ , \new_[72178]_ ,
    \new_[72182]_ , \new_[72183]_ , \new_[72186]_ , \new_[72189]_ ,
    \new_[72190]_ , \new_[72191]_ , \new_[72195]_ , \new_[72196]_ ,
    \new_[72199]_ , \new_[72202]_ , \new_[72203]_ , \new_[72204]_ ,
    \new_[72208]_ , \new_[72209]_ , \new_[72212]_ , \new_[72215]_ ,
    \new_[72216]_ , \new_[72217]_ , \new_[72221]_ , \new_[72222]_ ,
    \new_[72225]_ , \new_[72228]_ , \new_[72229]_ , \new_[72230]_ ,
    \new_[72234]_ , \new_[72235]_ , \new_[72238]_ , \new_[72241]_ ,
    \new_[72242]_ , \new_[72243]_ , \new_[72247]_ , \new_[72248]_ ,
    \new_[72251]_ , \new_[72254]_ , \new_[72255]_ , \new_[72256]_ ,
    \new_[72260]_ , \new_[72261]_ , \new_[72264]_ , \new_[72267]_ ,
    \new_[72268]_ , \new_[72269]_ , \new_[72273]_ , \new_[72274]_ ,
    \new_[72277]_ , \new_[72280]_ , \new_[72281]_ , \new_[72282]_ ,
    \new_[72286]_ , \new_[72287]_ , \new_[72290]_ , \new_[72293]_ ,
    \new_[72294]_ , \new_[72295]_ , \new_[72299]_ , \new_[72300]_ ,
    \new_[72303]_ , \new_[72306]_ , \new_[72307]_ , \new_[72308]_ ,
    \new_[72312]_ , \new_[72313]_ , \new_[72316]_ , \new_[72319]_ ,
    \new_[72320]_ , \new_[72321]_ , \new_[72325]_ , \new_[72326]_ ,
    \new_[72329]_ , \new_[72332]_ , \new_[72333]_ , \new_[72334]_ ,
    \new_[72338]_ , \new_[72339]_ , \new_[72342]_ , \new_[72345]_ ,
    \new_[72346]_ , \new_[72347]_ , \new_[72351]_ , \new_[72352]_ ,
    \new_[72355]_ , \new_[72358]_ , \new_[72359]_ , \new_[72360]_ ,
    \new_[72364]_ , \new_[72365]_ , \new_[72368]_ , \new_[72371]_ ,
    \new_[72372]_ , \new_[72373]_ , \new_[72377]_ , \new_[72378]_ ,
    \new_[72381]_ , \new_[72384]_ , \new_[72385]_ , \new_[72386]_ ,
    \new_[72390]_ , \new_[72391]_ , \new_[72394]_ , \new_[72397]_ ,
    \new_[72398]_ , \new_[72399]_ , \new_[72403]_ , \new_[72404]_ ,
    \new_[72407]_ , \new_[72410]_ , \new_[72411]_ , \new_[72412]_ ,
    \new_[72416]_ , \new_[72417]_ , \new_[72420]_ , \new_[72423]_ ,
    \new_[72424]_ , \new_[72425]_ , \new_[72429]_ , \new_[72430]_ ,
    \new_[72433]_ , \new_[72436]_ , \new_[72437]_ , \new_[72438]_ ,
    \new_[72442]_ , \new_[72443]_ , \new_[72446]_ , \new_[72449]_ ,
    \new_[72450]_ , \new_[72451]_ , \new_[72455]_ , \new_[72456]_ ,
    \new_[72459]_ , \new_[72462]_ , \new_[72463]_ , \new_[72464]_ ,
    \new_[72468]_ , \new_[72469]_ , \new_[72472]_ , \new_[72475]_ ,
    \new_[72476]_ , \new_[72477]_ , \new_[72481]_ , \new_[72482]_ ,
    \new_[72485]_ , \new_[72488]_ , \new_[72489]_ , \new_[72490]_ ,
    \new_[72494]_ , \new_[72495]_ , \new_[72498]_ , \new_[72501]_ ,
    \new_[72502]_ , \new_[72503]_ , \new_[72507]_ , \new_[72508]_ ,
    \new_[72511]_ , \new_[72514]_ , \new_[72515]_ , \new_[72516]_ ,
    \new_[72520]_ , \new_[72521]_ , \new_[72524]_ , \new_[72527]_ ,
    \new_[72528]_ , \new_[72529]_ , \new_[72533]_ , \new_[72534]_ ,
    \new_[72537]_ , \new_[72540]_ , \new_[72541]_ , \new_[72542]_ ,
    \new_[72546]_ , \new_[72547]_ , \new_[72550]_ , \new_[72553]_ ,
    \new_[72554]_ , \new_[72555]_ , \new_[72559]_ , \new_[72560]_ ,
    \new_[72563]_ , \new_[72566]_ , \new_[72567]_ , \new_[72568]_ ,
    \new_[72572]_ , \new_[72573]_ , \new_[72576]_ , \new_[72579]_ ,
    \new_[72580]_ , \new_[72581]_ , \new_[72585]_ , \new_[72586]_ ,
    \new_[72589]_ , \new_[72592]_ , \new_[72593]_ , \new_[72594]_ ,
    \new_[72598]_ , \new_[72599]_ , \new_[72602]_ , \new_[72605]_ ,
    \new_[72606]_ , \new_[72607]_ , \new_[72611]_ , \new_[72612]_ ,
    \new_[72615]_ , \new_[72618]_ , \new_[72619]_ , \new_[72620]_ ,
    \new_[72624]_ , \new_[72625]_ , \new_[72628]_ , \new_[72631]_ ,
    \new_[72632]_ , \new_[72633]_ , \new_[72637]_ , \new_[72638]_ ,
    \new_[72641]_ , \new_[72644]_ , \new_[72645]_ , \new_[72646]_ ,
    \new_[72650]_ , \new_[72651]_ , \new_[72654]_ , \new_[72657]_ ,
    \new_[72658]_ , \new_[72659]_ , \new_[72663]_ , \new_[72664]_ ,
    \new_[72667]_ , \new_[72670]_ , \new_[72671]_ , \new_[72672]_ ,
    \new_[72676]_ , \new_[72677]_ , \new_[72680]_ , \new_[72683]_ ,
    \new_[72684]_ , \new_[72685]_ , \new_[72689]_ , \new_[72690]_ ,
    \new_[72693]_ , \new_[72696]_ , \new_[72697]_ , \new_[72698]_ ,
    \new_[72702]_ , \new_[72703]_ , \new_[72706]_ , \new_[72709]_ ,
    \new_[72710]_ , \new_[72711]_ , \new_[72715]_ , \new_[72716]_ ,
    \new_[72719]_ , \new_[72722]_ , \new_[72723]_ , \new_[72724]_ ,
    \new_[72728]_ , \new_[72729]_ , \new_[72732]_ , \new_[72735]_ ,
    \new_[72736]_ , \new_[72737]_ , \new_[72741]_ , \new_[72742]_ ,
    \new_[72745]_ , \new_[72748]_ , \new_[72749]_ , \new_[72750]_ ,
    \new_[72754]_ , \new_[72755]_ , \new_[72758]_ , \new_[72761]_ ,
    \new_[72762]_ , \new_[72763]_ , \new_[72767]_ , \new_[72768]_ ,
    \new_[72771]_ , \new_[72774]_ , \new_[72775]_ , \new_[72776]_ ,
    \new_[72780]_ , \new_[72781]_ , \new_[72784]_ , \new_[72787]_ ,
    \new_[72788]_ , \new_[72789]_ , \new_[72793]_ , \new_[72794]_ ,
    \new_[72797]_ , \new_[72800]_ , \new_[72801]_ , \new_[72802]_ ,
    \new_[72806]_ , \new_[72807]_ , \new_[72810]_ , \new_[72813]_ ,
    \new_[72814]_ , \new_[72815]_ , \new_[72819]_ , \new_[72820]_ ,
    \new_[72823]_ , \new_[72826]_ , \new_[72827]_ , \new_[72828]_ ,
    \new_[72832]_ , \new_[72833]_ , \new_[72836]_ , \new_[72839]_ ,
    \new_[72840]_ , \new_[72841]_ , \new_[72845]_ , \new_[72846]_ ,
    \new_[72849]_ , \new_[72852]_ , \new_[72853]_ , \new_[72854]_ ,
    \new_[72858]_ , \new_[72859]_ , \new_[72862]_ , \new_[72865]_ ,
    \new_[72866]_ , \new_[72867]_ , \new_[72871]_ , \new_[72872]_ ,
    \new_[72875]_ , \new_[72878]_ , \new_[72879]_ , \new_[72880]_ ,
    \new_[72884]_ , \new_[72885]_ , \new_[72888]_ , \new_[72891]_ ,
    \new_[72892]_ , \new_[72893]_ , \new_[72897]_ , \new_[72898]_ ,
    \new_[72901]_ , \new_[72904]_ , \new_[72905]_ , \new_[72906]_ ,
    \new_[72910]_ , \new_[72911]_ , \new_[72914]_ , \new_[72917]_ ,
    \new_[72918]_ , \new_[72919]_ , \new_[72923]_ , \new_[72924]_ ,
    \new_[72927]_ , \new_[72930]_ , \new_[72931]_ , \new_[72932]_ ,
    \new_[72936]_ , \new_[72937]_ , \new_[72940]_ , \new_[72943]_ ,
    \new_[72944]_ , \new_[72945]_ , \new_[72949]_ , \new_[72950]_ ,
    \new_[72953]_ , \new_[72956]_ , \new_[72957]_ , \new_[72958]_ ,
    \new_[72962]_ , \new_[72963]_ , \new_[72966]_ , \new_[72969]_ ,
    \new_[72970]_ , \new_[72971]_ , \new_[72975]_ , \new_[72976]_ ,
    \new_[72979]_ , \new_[72982]_ , \new_[72983]_ , \new_[72984]_ ,
    \new_[72988]_ , \new_[72989]_ , \new_[72992]_ , \new_[72995]_ ,
    \new_[72996]_ , \new_[72997]_ , \new_[73001]_ , \new_[73002]_ ,
    \new_[73005]_ , \new_[73008]_ , \new_[73009]_ , \new_[73010]_ ,
    \new_[73014]_ , \new_[73015]_ , \new_[73018]_ , \new_[73021]_ ,
    \new_[73022]_ , \new_[73023]_ , \new_[73027]_ , \new_[73028]_ ,
    \new_[73031]_ , \new_[73034]_ , \new_[73035]_ , \new_[73036]_ ,
    \new_[73040]_ , \new_[73041]_ , \new_[73044]_ , \new_[73047]_ ,
    \new_[73048]_ , \new_[73049]_ , \new_[73053]_ , \new_[73054]_ ,
    \new_[73057]_ , \new_[73060]_ , \new_[73061]_ , \new_[73062]_ ,
    \new_[73066]_ , \new_[73067]_ , \new_[73070]_ , \new_[73073]_ ,
    \new_[73074]_ , \new_[73075]_ , \new_[73079]_ , \new_[73080]_ ,
    \new_[73083]_ , \new_[73086]_ , \new_[73087]_ , \new_[73088]_ ,
    \new_[73092]_ , \new_[73093]_ , \new_[73096]_ , \new_[73099]_ ,
    \new_[73100]_ , \new_[73101]_ , \new_[73105]_ , \new_[73106]_ ,
    \new_[73109]_ , \new_[73112]_ , \new_[73113]_ , \new_[73114]_ ,
    \new_[73118]_ , \new_[73119]_ , \new_[73122]_ , \new_[73125]_ ,
    \new_[73126]_ , \new_[73127]_ , \new_[73131]_ , \new_[73132]_ ,
    \new_[73135]_ , \new_[73138]_ , \new_[73139]_ , \new_[73140]_ ,
    \new_[73144]_ , \new_[73145]_ , \new_[73148]_ , \new_[73151]_ ,
    \new_[73152]_ , \new_[73153]_ , \new_[73157]_ , \new_[73158]_ ,
    \new_[73161]_ , \new_[73164]_ , \new_[73165]_ , \new_[73166]_ ,
    \new_[73170]_ , \new_[73171]_ , \new_[73174]_ , \new_[73177]_ ,
    \new_[73178]_ , \new_[73179]_ , \new_[73183]_ , \new_[73184]_ ,
    \new_[73187]_ , \new_[73190]_ , \new_[73191]_ , \new_[73192]_ ,
    \new_[73196]_ , \new_[73197]_ , \new_[73200]_ , \new_[73203]_ ,
    \new_[73204]_ , \new_[73205]_ , \new_[73209]_ , \new_[73210]_ ,
    \new_[73213]_ , \new_[73216]_ , \new_[73217]_ , \new_[73218]_ ,
    \new_[73222]_ , \new_[73223]_ , \new_[73226]_ , \new_[73229]_ ,
    \new_[73230]_ , \new_[73231]_ , \new_[73235]_ , \new_[73236]_ ,
    \new_[73239]_ , \new_[73242]_ , \new_[73243]_ , \new_[73244]_ ,
    \new_[73248]_ , \new_[73249]_ , \new_[73252]_ , \new_[73255]_ ,
    \new_[73256]_ , \new_[73257]_ , \new_[73261]_ , \new_[73262]_ ,
    \new_[73265]_ , \new_[73268]_ , \new_[73269]_ , \new_[73270]_ ,
    \new_[73274]_ , \new_[73275]_ , \new_[73278]_ , \new_[73281]_ ,
    \new_[73282]_ , \new_[73283]_ , \new_[73287]_ , \new_[73288]_ ,
    \new_[73291]_ , \new_[73294]_ , \new_[73295]_ , \new_[73296]_ ,
    \new_[73300]_ , \new_[73301]_ , \new_[73304]_ , \new_[73307]_ ,
    \new_[73308]_ , \new_[73309]_ , \new_[73313]_ , \new_[73314]_ ,
    \new_[73317]_ , \new_[73320]_ , \new_[73321]_ , \new_[73322]_ ,
    \new_[73326]_ , \new_[73327]_ , \new_[73330]_ , \new_[73333]_ ,
    \new_[73334]_ , \new_[73335]_ , \new_[73339]_ , \new_[73340]_ ,
    \new_[73343]_ , \new_[73346]_ , \new_[73347]_ , \new_[73348]_ ,
    \new_[73352]_ , \new_[73353]_ , \new_[73356]_ , \new_[73359]_ ,
    \new_[73360]_ , \new_[73361]_ , \new_[73365]_ , \new_[73366]_ ,
    \new_[73369]_ , \new_[73372]_ , \new_[73373]_ , \new_[73374]_ ,
    \new_[73378]_ , \new_[73379]_ , \new_[73382]_ , \new_[73385]_ ,
    \new_[73386]_ , \new_[73387]_ , \new_[73391]_ , \new_[73392]_ ,
    \new_[73395]_ , \new_[73398]_ , \new_[73399]_ , \new_[73400]_ ,
    \new_[73404]_ , \new_[73405]_ , \new_[73408]_ , \new_[73411]_ ,
    \new_[73412]_ , \new_[73413]_ , \new_[73417]_ , \new_[73418]_ ,
    \new_[73421]_ , \new_[73424]_ , \new_[73425]_ , \new_[73426]_ ,
    \new_[73430]_ , \new_[73431]_ , \new_[73434]_ , \new_[73437]_ ,
    \new_[73438]_ , \new_[73439]_ , \new_[73443]_ , \new_[73444]_ ,
    \new_[73447]_ , \new_[73450]_ , \new_[73451]_ , \new_[73452]_ ,
    \new_[73456]_ , \new_[73457]_ , \new_[73460]_ , \new_[73463]_ ,
    \new_[73464]_ , \new_[73465]_ , \new_[73469]_ , \new_[73470]_ ,
    \new_[73473]_ , \new_[73476]_ , \new_[73477]_ , \new_[73478]_ ,
    \new_[73482]_ , \new_[73483]_ , \new_[73486]_ , \new_[73489]_ ,
    \new_[73490]_ , \new_[73491]_ , \new_[73495]_ , \new_[73496]_ ,
    \new_[73499]_ , \new_[73502]_ , \new_[73503]_ , \new_[73504]_ ,
    \new_[73508]_ , \new_[73509]_ , \new_[73512]_ , \new_[73515]_ ,
    \new_[73516]_ , \new_[73517]_ , \new_[73521]_ , \new_[73522]_ ,
    \new_[73525]_ , \new_[73528]_ , \new_[73529]_ , \new_[73530]_ ,
    \new_[73534]_ , \new_[73535]_ , \new_[73538]_ , \new_[73541]_ ,
    \new_[73542]_ , \new_[73543]_ , \new_[73547]_ , \new_[73548]_ ,
    \new_[73551]_ , \new_[73554]_ , \new_[73555]_ , \new_[73556]_ ,
    \new_[73560]_ , \new_[73561]_ , \new_[73564]_ , \new_[73567]_ ,
    \new_[73568]_ , \new_[73569]_ , \new_[73573]_ , \new_[73574]_ ,
    \new_[73577]_ , \new_[73580]_ , \new_[73581]_ , \new_[73582]_ ,
    \new_[73586]_ , \new_[73587]_ , \new_[73590]_ , \new_[73593]_ ,
    \new_[73594]_ , \new_[73595]_ , \new_[73599]_ , \new_[73600]_ ,
    \new_[73603]_ , \new_[73606]_ , \new_[73607]_ , \new_[73608]_ ,
    \new_[73612]_ , \new_[73613]_ , \new_[73616]_ , \new_[73619]_ ,
    \new_[73620]_ , \new_[73621]_ , \new_[73625]_ , \new_[73626]_ ,
    \new_[73629]_ , \new_[73632]_ , \new_[73633]_ , \new_[73634]_ ,
    \new_[73638]_ , \new_[73639]_ , \new_[73642]_ , \new_[73645]_ ,
    \new_[73646]_ , \new_[73647]_ , \new_[73651]_ , \new_[73652]_ ,
    \new_[73655]_ , \new_[73658]_ , \new_[73659]_ , \new_[73660]_ ,
    \new_[73664]_ , \new_[73665]_ , \new_[73668]_ , \new_[73671]_ ,
    \new_[73672]_ , \new_[73673]_ , \new_[73677]_ , \new_[73678]_ ,
    \new_[73681]_ , \new_[73684]_ , \new_[73685]_ , \new_[73686]_ ,
    \new_[73690]_ , \new_[73691]_ , \new_[73694]_ , \new_[73697]_ ,
    \new_[73698]_ , \new_[73699]_ , \new_[73703]_ , \new_[73704]_ ,
    \new_[73707]_ , \new_[73710]_ , \new_[73711]_ , \new_[73712]_ ,
    \new_[73716]_ , \new_[73717]_ , \new_[73720]_ , \new_[73723]_ ,
    \new_[73724]_ , \new_[73725]_ , \new_[73729]_ , \new_[73730]_ ,
    \new_[73733]_ , \new_[73736]_ , \new_[73737]_ , \new_[73738]_ ,
    \new_[73742]_ , \new_[73743]_ , \new_[73746]_ , \new_[73749]_ ,
    \new_[73750]_ , \new_[73751]_ , \new_[73755]_ , \new_[73756]_ ,
    \new_[73759]_ , \new_[73762]_ , \new_[73763]_ , \new_[73764]_ ,
    \new_[73768]_ , \new_[73769]_ , \new_[73772]_ , \new_[73775]_ ,
    \new_[73776]_ , \new_[73777]_ , \new_[73781]_ , \new_[73782]_ ,
    \new_[73785]_ , \new_[73788]_ , \new_[73789]_ , \new_[73790]_ ,
    \new_[73794]_ , \new_[73795]_ , \new_[73798]_ , \new_[73801]_ ,
    \new_[73802]_ , \new_[73803]_ , \new_[73807]_ , \new_[73808]_ ,
    \new_[73811]_ , \new_[73814]_ , \new_[73815]_ , \new_[73816]_ ,
    \new_[73820]_ , \new_[73821]_ , \new_[73824]_ , \new_[73827]_ ,
    \new_[73828]_ , \new_[73829]_ , \new_[73833]_ , \new_[73834]_ ,
    \new_[73837]_ , \new_[73840]_ , \new_[73841]_ , \new_[73842]_ ,
    \new_[73846]_ , \new_[73847]_ , \new_[73850]_ , \new_[73853]_ ,
    \new_[73854]_ , \new_[73855]_ , \new_[73859]_ , \new_[73860]_ ,
    \new_[73863]_ , \new_[73866]_ , \new_[73867]_ , \new_[73868]_ ,
    \new_[73872]_ , \new_[73873]_ , \new_[73876]_ , \new_[73879]_ ,
    \new_[73880]_ , \new_[73881]_ , \new_[73885]_ , \new_[73886]_ ,
    \new_[73889]_ , \new_[73892]_ , \new_[73893]_ , \new_[73894]_ ,
    \new_[73898]_ , \new_[73899]_ , \new_[73902]_ , \new_[73905]_ ,
    \new_[73906]_ , \new_[73907]_ , \new_[73911]_ , \new_[73912]_ ,
    \new_[73915]_ , \new_[73918]_ , \new_[73919]_ , \new_[73920]_ ,
    \new_[73924]_ , \new_[73925]_ , \new_[73928]_ , \new_[73931]_ ,
    \new_[73932]_ , \new_[73933]_ , \new_[73937]_ , \new_[73938]_ ,
    \new_[73941]_ , \new_[73944]_ , \new_[73945]_ , \new_[73946]_ ,
    \new_[73950]_ , \new_[73951]_ , \new_[73954]_ , \new_[73957]_ ,
    \new_[73958]_ , \new_[73959]_ , \new_[73963]_ , \new_[73964]_ ,
    \new_[73967]_ , \new_[73970]_ , \new_[73971]_ , \new_[73972]_ ,
    \new_[73976]_ , \new_[73977]_ , \new_[73980]_ , \new_[73983]_ ,
    \new_[73984]_ , \new_[73985]_ , \new_[73989]_ , \new_[73990]_ ,
    \new_[73993]_ , \new_[73996]_ , \new_[73997]_ , \new_[73998]_ ,
    \new_[74002]_ , \new_[74003]_ , \new_[74006]_ , \new_[74009]_ ,
    \new_[74010]_ , \new_[74011]_ , \new_[74015]_ , \new_[74016]_ ,
    \new_[74019]_ , \new_[74022]_ , \new_[74023]_ , \new_[74024]_ ,
    \new_[74028]_ , \new_[74029]_ , \new_[74032]_ , \new_[74035]_ ,
    \new_[74036]_ , \new_[74037]_ , \new_[74041]_ , \new_[74042]_ ,
    \new_[74045]_ , \new_[74048]_ , \new_[74049]_ , \new_[74050]_ ,
    \new_[74054]_ , \new_[74055]_ , \new_[74058]_ , \new_[74061]_ ,
    \new_[74062]_ , \new_[74063]_ , \new_[74067]_ , \new_[74068]_ ,
    \new_[74071]_ , \new_[74074]_ , \new_[74075]_ , \new_[74076]_ ,
    \new_[74080]_ , \new_[74081]_ , \new_[74084]_ , \new_[74087]_ ,
    \new_[74088]_ , \new_[74089]_ , \new_[74093]_ , \new_[74094]_ ,
    \new_[74097]_ , \new_[74100]_ , \new_[74101]_ , \new_[74102]_ ,
    \new_[74106]_ , \new_[74107]_ , \new_[74110]_ , \new_[74113]_ ,
    \new_[74114]_ , \new_[74115]_ , \new_[74119]_ , \new_[74120]_ ,
    \new_[74123]_ , \new_[74126]_ , \new_[74127]_ , \new_[74128]_ ,
    \new_[74132]_ , \new_[74133]_ , \new_[74136]_ , \new_[74139]_ ,
    \new_[74140]_ , \new_[74141]_ , \new_[74145]_ , \new_[74146]_ ,
    \new_[74149]_ , \new_[74152]_ , \new_[74153]_ , \new_[74154]_ ,
    \new_[74158]_ , \new_[74159]_ , \new_[74162]_ , \new_[74165]_ ,
    \new_[74166]_ , \new_[74167]_ , \new_[74171]_ , \new_[74172]_ ,
    \new_[74175]_ , \new_[74178]_ , \new_[74179]_ , \new_[74180]_ ,
    \new_[74184]_ , \new_[74185]_ , \new_[74188]_ , \new_[74191]_ ,
    \new_[74192]_ , \new_[74193]_ , \new_[74197]_ , \new_[74198]_ ,
    \new_[74201]_ , \new_[74204]_ , \new_[74205]_ , \new_[74206]_ ,
    \new_[74210]_ , \new_[74211]_ , \new_[74214]_ , \new_[74217]_ ,
    \new_[74218]_ , \new_[74219]_ , \new_[74223]_ , \new_[74224]_ ,
    \new_[74227]_ , \new_[74230]_ , \new_[74231]_ , \new_[74232]_ ,
    \new_[74236]_ , \new_[74237]_ , \new_[74240]_ , \new_[74243]_ ,
    \new_[74244]_ , \new_[74245]_ , \new_[74249]_ , \new_[74250]_ ,
    \new_[74253]_ , \new_[74256]_ , \new_[74257]_ , \new_[74258]_ ,
    \new_[74262]_ , \new_[74263]_ , \new_[74266]_ , \new_[74269]_ ,
    \new_[74270]_ , \new_[74271]_ , \new_[74275]_ , \new_[74276]_ ,
    \new_[74279]_ , \new_[74282]_ , \new_[74283]_ , \new_[74284]_ ,
    \new_[74288]_ , \new_[74289]_ , \new_[74292]_ , \new_[74295]_ ,
    \new_[74296]_ , \new_[74297]_ , \new_[74301]_ , \new_[74302]_ ,
    \new_[74305]_ , \new_[74308]_ , \new_[74309]_ , \new_[74310]_ ,
    \new_[74314]_ , \new_[74315]_ , \new_[74318]_ , \new_[74321]_ ,
    \new_[74322]_ , \new_[74323]_ , \new_[74327]_ , \new_[74328]_ ,
    \new_[74331]_ , \new_[74334]_ , \new_[74335]_ , \new_[74336]_ ,
    \new_[74340]_ , \new_[74341]_ , \new_[74344]_ , \new_[74347]_ ,
    \new_[74348]_ , \new_[74349]_ , \new_[74353]_ , \new_[74354]_ ,
    \new_[74357]_ , \new_[74360]_ , \new_[74361]_ , \new_[74362]_ ,
    \new_[74366]_ , \new_[74367]_ , \new_[74370]_ , \new_[74373]_ ,
    \new_[74374]_ , \new_[74375]_ , \new_[74379]_ , \new_[74380]_ ,
    \new_[74383]_ , \new_[74386]_ , \new_[74387]_ , \new_[74388]_ ,
    \new_[74392]_ , \new_[74393]_ , \new_[74396]_ , \new_[74399]_ ,
    \new_[74400]_ , \new_[74401]_ , \new_[74405]_ , \new_[74406]_ ,
    \new_[74409]_ , \new_[74412]_ , \new_[74413]_ , \new_[74414]_ ,
    \new_[74418]_ , \new_[74419]_ , \new_[74422]_ , \new_[74425]_ ,
    \new_[74426]_ , \new_[74427]_ , \new_[74431]_ , \new_[74432]_ ,
    \new_[74435]_ , \new_[74438]_ , \new_[74439]_ , \new_[74440]_ ,
    \new_[74444]_ , \new_[74445]_ , \new_[74448]_ , \new_[74451]_ ,
    \new_[74452]_ , \new_[74453]_ , \new_[74457]_ , \new_[74458]_ ,
    \new_[74461]_ , \new_[74464]_ , \new_[74465]_ , \new_[74466]_ ,
    \new_[74470]_ , \new_[74471]_ , \new_[74474]_ , \new_[74477]_ ,
    \new_[74478]_ , \new_[74479]_ , \new_[74483]_ , \new_[74484]_ ,
    \new_[74487]_ , \new_[74490]_ , \new_[74491]_ , \new_[74492]_ ,
    \new_[74496]_ , \new_[74497]_ , \new_[74500]_ , \new_[74503]_ ,
    \new_[74504]_ , \new_[74505]_ , \new_[74509]_ , \new_[74510]_ ,
    \new_[74513]_ , \new_[74516]_ , \new_[74517]_ , \new_[74518]_ ,
    \new_[74522]_ , \new_[74523]_ , \new_[74526]_ , \new_[74529]_ ,
    \new_[74530]_ , \new_[74531]_ , \new_[74535]_ , \new_[74536]_ ,
    \new_[74539]_ , \new_[74542]_ , \new_[74543]_ , \new_[74544]_ ,
    \new_[74548]_ , \new_[74549]_ , \new_[74552]_ , \new_[74555]_ ,
    \new_[74556]_ , \new_[74557]_ , \new_[74561]_ , \new_[74562]_ ,
    \new_[74565]_ , \new_[74568]_ , \new_[74569]_ , \new_[74570]_ ,
    \new_[74574]_ , \new_[74575]_ , \new_[74578]_ , \new_[74581]_ ,
    \new_[74582]_ , \new_[74583]_ , \new_[74587]_ , \new_[74588]_ ,
    \new_[74591]_ , \new_[74594]_ , \new_[74595]_ , \new_[74596]_ ,
    \new_[74600]_ , \new_[74601]_ , \new_[74604]_ , \new_[74607]_ ,
    \new_[74608]_ , \new_[74609]_ , \new_[74613]_ , \new_[74614]_ ,
    \new_[74617]_ , \new_[74620]_ , \new_[74621]_ , \new_[74622]_ ,
    \new_[74626]_ , \new_[74627]_ , \new_[74630]_ , \new_[74633]_ ,
    \new_[74634]_ , \new_[74635]_ , \new_[74639]_ , \new_[74640]_ ,
    \new_[74643]_ , \new_[74646]_ , \new_[74647]_ , \new_[74648]_ ,
    \new_[74652]_ , \new_[74653]_ , \new_[74656]_ , \new_[74659]_ ,
    \new_[74660]_ , \new_[74661]_ , \new_[74665]_ , \new_[74666]_ ,
    \new_[74669]_ , \new_[74672]_ , \new_[74673]_ , \new_[74674]_ ,
    \new_[74678]_ , \new_[74679]_ , \new_[74682]_ , \new_[74685]_ ,
    \new_[74686]_ , \new_[74687]_ , \new_[74691]_ , \new_[74692]_ ,
    \new_[74695]_ , \new_[74698]_ , \new_[74699]_ , \new_[74700]_ ,
    \new_[74704]_ , \new_[74705]_ , \new_[74708]_ , \new_[74711]_ ,
    \new_[74712]_ , \new_[74713]_ , \new_[74717]_ , \new_[74718]_ ,
    \new_[74721]_ , \new_[74724]_ , \new_[74725]_ , \new_[74726]_ ,
    \new_[74730]_ , \new_[74731]_ , \new_[74734]_ , \new_[74737]_ ,
    \new_[74738]_ , \new_[74739]_ , \new_[74743]_ , \new_[74744]_ ,
    \new_[74747]_ , \new_[74750]_ , \new_[74751]_ , \new_[74752]_ ,
    \new_[74756]_ , \new_[74757]_ , \new_[74760]_ , \new_[74763]_ ,
    \new_[74764]_ , \new_[74765]_ , \new_[74769]_ , \new_[74770]_ ,
    \new_[74773]_ , \new_[74776]_ , \new_[74777]_ , \new_[74778]_ ,
    \new_[74782]_ , \new_[74783]_ , \new_[74786]_ , \new_[74789]_ ,
    \new_[74790]_ , \new_[74791]_ , \new_[74795]_ , \new_[74796]_ ,
    \new_[74799]_ , \new_[74802]_ , \new_[74803]_ , \new_[74804]_ ,
    \new_[74808]_ , \new_[74809]_ , \new_[74812]_ , \new_[74815]_ ,
    \new_[74816]_ , \new_[74817]_ , \new_[74821]_ , \new_[74822]_ ,
    \new_[74825]_ , \new_[74828]_ , \new_[74829]_ , \new_[74830]_ ,
    \new_[74834]_ , \new_[74835]_ , \new_[74838]_ , \new_[74841]_ ,
    \new_[74842]_ , \new_[74843]_ , \new_[74847]_ , \new_[74848]_ ,
    \new_[74851]_ , \new_[74854]_ , \new_[74855]_ , \new_[74856]_ ,
    \new_[74860]_ , \new_[74861]_ , \new_[74864]_ , \new_[74867]_ ,
    \new_[74868]_ , \new_[74869]_ , \new_[74873]_ , \new_[74874]_ ,
    \new_[74877]_ , \new_[74880]_ , \new_[74881]_ , \new_[74882]_ ,
    \new_[74886]_ , \new_[74887]_ , \new_[74890]_ , \new_[74893]_ ,
    \new_[74894]_ , \new_[74895]_ , \new_[74899]_ , \new_[74900]_ ,
    \new_[74903]_ , \new_[74906]_ , \new_[74907]_ , \new_[74908]_ ,
    \new_[74912]_ , \new_[74913]_ , \new_[74916]_ , \new_[74919]_ ,
    \new_[74920]_ , \new_[74921]_ , \new_[74925]_ , \new_[74926]_ ,
    \new_[74929]_ , \new_[74932]_ , \new_[74933]_ , \new_[74934]_ ,
    \new_[74938]_ , \new_[74939]_ , \new_[74942]_ , \new_[74945]_ ,
    \new_[74946]_ , \new_[74947]_ , \new_[74951]_ , \new_[74952]_ ,
    \new_[74955]_ , \new_[74958]_ , \new_[74959]_ , \new_[74960]_ ,
    \new_[74964]_ , \new_[74965]_ , \new_[74968]_ , \new_[74971]_ ,
    \new_[74972]_ , \new_[74973]_ , \new_[74977]_ , \new_[74978]_ ,
    \new_[74981]_ , \new_[74984]_ , \new_[74985]_ , \new_[74986]_ ,
    \new_[74990]_ , \new_[74991]_ , \new_[74994]_ , \new_[74997]_ ,
    \new_[74998]_ , \new_[74999]_ , \new_[75003]_ , \new_[75004]_ ,
    \new_[75007]_ , \new_[75010]_ , \new_[75011]_ , \new_[75012]_ ,
    \new_[75016]_ , \new_[75017]_ , \new_[75020]_ , \new_[75023]_ ,
    \new_[75024]_ , \new_[75025]_ , \new_[75029]_ , \new_[75030]_ ,
    \new_[75033]_ , \new_[75036]_ , \new_[75037]_ , \new_[75038]_ ,
    \new_[75042]_ , \new_[75043]_ , \new_[75046]_ , \new_[75049]_ ,
    \new_[75050]_ , \new_[75051]_ , \new_[75055]_ , \new_[75056]_ ,
    \new_[75059]_ , \new_[75062]_ , \new_[75063]_ , \new_[75064]_ ,
    \new_[75068]_ , \new_[75069]_ , \new_[75072]_ , \new_[75075]_ ,
    \new_[75076]_ , \new_[75077]_ , \new_[75081]_ , \new_[75082]_ ,
    \new_[75085]_ , \new_[75088]_ , \new_[75089]_ , \new_[75090]_ ,
    \new_[75094]_ , \new_[75095]_ , \new_[75098]_ , \new_[75101]_ ,
    \new_[75102]_ , \new_[75103]_ , \new_[75107]_ , \new_[75108]_ ,
    \new_[75111]_ , \new_[75114]_ , \new_[75115]_ , \new_[75116]_ ,
    \new_[75120]_ , \new_[75121]_ , \new_[75124]_ , \new_[75127]_ ,
    \new_[75128]_ , \new_[75129]_ , \new_[75133]_ , \new_[75134]_ ,
    \new_[75137]_ , \new_[75140]_ , \new_[75141]_ , \new_[75142]_ ,
    \new_[75146]_ , \new_[75147]_ , \new_[75150]_ , \new_[75153]_ ,
    \new_[75154]_ , \new_[75155]_ , \new_[75159]_ , \new_[75160]_ ,
    \new_[75163]_ , \new_[75166]_ , \new_[75167]_ , \new_[75168]_ ,
    \new_[75172]_ , \new_[75173]_ , \new_[75176]_ , \new_[75179]_ ,
    \new_[75180]_ , \new_[75181]_ , \new_[75185]_ , \new_[75186]_ ,
    \new_[75189]_ , \new_[75192]_ , \new_[75193]_ , \new_[75194]_ ,
    \new_[75198]_ , \new_[75199]_ , \new_[75202]_ , \new_[75205]_ ,
    \new_[75206]_ , \new_[75207]_ , \new_[75211]_ , \new_[75212]_ ,
    \new_[75215]_ , \new_[75218]_ , \new_[75219]_ , \new_[75220]_ ,
    \new_[75224]_ , \new_[75225]_ , \new_[75228]_ , \new_[75231]_ ,
    \new_[75232]_ , \new_[75233]_ , \new_[75237]_ , \new_[75238]_ ,
    \new_[75241]_ , \new_[75244]_ , \new_[75245]_ , \new_[75246]_ ,
    \new_[75250]_ , \new_[75251]_ , \new_[75254]_ , \new_[75257]_ ,
    \new_[75258]_ , \new_[75259]_ , \new_[75263]_ , \new_[75264]_ ,
    \new_[75267]_ , \new_[75270]_ , \new_[75271]_ , \new_[75272]_ ,
    \new_[75276]_ , \new_[75277]_ , \new_[75280]_ , \new_[75283]_ ,
    \new_[75284]_ , \new_[75285]_ , \new_[75289]_ , \new_[75290]_ ,
    \new_[75293]_ , \new_[75296]_ , \new_[75297]_ , \new_[75298]_ ,
    \new_[75302]_ , \new_[75303]_ , \new_[75306]_ , \new_[75309]_ ,
    \new_[75310]_ , \new_[75311]_ , \new_[75315]_ , \new_[75316]_ ,
    \new_[75319]_ , \new_[75322]_ , \new_[75323]_ , \new_[75324]_ ,
    \new_[75328]_ , \new_[75329]_ , \new_[75332]_ , \new_[75335]_ ,
    \new_[75336]_ , \new_[75337]_ , \new_[75341]_ , \new_[75342]_ ,
    \new_[75345]_ , \new_[75348]_ , \new_[75349]_ , \new_[75350]_ ,
    \new_[75354]_ , \new_[75355]_ , \new_[75358]_ , \new_[75361]_ ,
    \new_[75362]_ , \new_[75363]_ , \new_[75367]_ , \new_[75368]_ ,
    \new_[75371]_ , \new_[75374]_ , \new_[75375]_ , \new_[75376]_ ,
    \new_[75380]_ , \new_[75381]_ , \new_[75384]_ , \new_[75387]_ ,
    \new_[75388]_ , \new_[75389]_ , \new_[75393]_ , \new_[75394]_ ,
    \new_[75397]_ , \new_[75400]_ , \new_[75401]_ , \new_[75402]_ ,
    \new_[75406]_ , \new_[75407]_ , \new_[75410]_ , \new_[75413]_ ,
    \new_[75414]_ , \new_[75415]_ , \new_[75419]_ , \new_[75420]_ ,
    \new_[75423]_ , \new_[75426]_ , \new_[75427]_ , \new_[75428]_ ,
    \new_[75432]_ , \new_[75433]_ , \new_[75436]_ , \new_[75439]_ ,
    \new_[75440]_ , \new_[75441]_ , \new_[75445]_ , \new_[75446]_ ,
    \new_[75449]_ , \new_[75452]_ , \new_[75453]_ , \new_[75454]_ ,
    \new_[75458]_ , \new_[75459]_ , \new_[75462]_ , \new_[75465]_ ,
    \new_[75466]_ , \new_[75467]_ , \new_[75471]_ , \new_[75472]_ ,
    \new_[75475]_ , \new_[75478]_ , \new_[75479]_ , \new_[75480]_ ,
    \new_[75484]_ , \new_[75485]_ , \new_[75488]_ , \new_[75491]_ ,
    \new_[75492]_ , \new_[75493]_ , \new_[75497]_ , \new_[75498]_ ,
    \new_[75501]_ , \new_[75504]_ , \new_[75505]_ , \new_[75506]_ ,
    \new_[75510]_ , \new_[75511]_ , \new_[75514]_ , \new_[75517]_ ,
    \new_[75518]_ , \new_[75519]_ , \new_[75523]_ , \new_[75524]_ ,
    \new_[75527]_ , \new_[75530]_ , \new_[75531]_ , \new_[75532]_ ,
    \new_[75536]_ , \new_[75537]_ , \new_[75540]_ , \new_[75543]_ ,
    \new_[75544]_ , \new_[75545]_ , \new_[75549]_ , \new_[75550]_ ,
    \new_[75553]_ , \new_[75556]_ , \new_[75557]_ , \new_[75558]_ ,
    \new_[75562]_ , \new_[75563]_ , \new_[75566]_ , \new_[75569]_ ,
    \new_[75570]_ , \new_[75571]_ , \new_[75575]_ , \new_[75576]_ ,
    \new_[75579]_ , \new_[75582]_ , \new_[75583]_ , \new_[75584]_ ,
    \new_[75588]_ , \new_[75589]_ , \new_[75592]_ , \new_[75595]_ ,
    \new_[75596]_ , \new_[75597]_ , \new_[75601]_ , \new_[75602]_ ,
    \new_[75605]_ , \new_[75608]_ , \new_[75609]_ , \new_[75610]_ ,
    \new_[75614]_ , \new_[75615]_ , \new_[75618]_ , \new_[75621]_ ,
    \new_[75622]_ , \new_[75623]_ , \new_[75627]_ , \new_[75628]_ ,
    \new_[75631]_ , \new_[75634]_ , \new_[75635]_ , \new_[75636]_ ,
    \new_[75640]_ , \new_[75641]_ , \new_[75644]_ , \new_[75647]_ ,
    \new_[75648]_ , \new_[75649]_ , \new_[75653]_ , \new_[75654]_ ,
    \new_[75657]_ , \new_[75660]_ , \new_[75661]_ , \new_[75662]_ ,
    \new_[75666]_ , \new_[75667]_ , \new_[75670]_ , \new_[75673]_ ,
    \new_[75674]_ , \new_[75675]_ , \new_[75679]_ , \new_[75680]_ ,
    \new_[75683]_ , \new_[75686]_ , \new_[75687]_ , \new_[75688]_ ,
    \new_[75692]_ , \new_[75693]_ , \new_[75696]_ , \new_[75699]_ ,
    \new_[75700]_ , \new_[75701]_ , \new_[75705]_ , \new_[75706]_ ,
    \new_[75709]_ , \new_[75712]_ , \new_[75713]_ , \new_[75714]_ ,
    \new_[75718]_ , \new_[75719]_ , \new_[75722]_ , \new_[75725]_ ,
    \new_[75726]_ , \new_[75727]_ , \new_[75731]_ , \new_[75732]_ ,
    \new_[75735]_ , \new_[75738]_ , \new_[75739]_ , \new_[75740]_ ,
    \new_[75744]_ , \new_[75745]_ , \new_[75748]_ , \new_[75751]_ ,
    \new_[75752]_ , \new_[75753]_ , \new_[75757]_ , \new_[75758]_ ,
    \new_[75761]_ , \new_[75764]_ , \new_[75765]_ , \new_[75766]_ ,
    \new_[75770]_ , \new_[75771]_ , \new_[75774]_ , \new_[75777]_ ,
    \new_[75778]_ , \new_[75779]_ , \new_[75783]_ , \new_[75784]_ ,
    \new_[75787]_ , \new_[75790]_ , \new_[75791]_ , \new_[75792]_ ,
    \new_[75796]_ , \new_[75797]_ , \new_[75800]_ , \new_[75803]_ ,
    \new_[75804]_ , \new_[75805]_ , \new_[75809]_ , \new_[75810]_ ,
    \new_[75813]_ , \new_[75816]_ , \new_[75817]_ , \new_[75818]_ ,
    \new_[75822]_ , \new_[75823]_ , \new_[75826]_ , \new_[75829]_ ,
    \new_[75830]_ , \new_[75831]_ , \new_[75835]_ , \new_[75836]_ ,
    \new_[75839]_ , \new_[75842]_ , \new_[75843]_ , \new_[75844]_ ,
    \new_[75848]_ , \new_[75849]_ , \new_[75852]_ , \new_[75855]_ ,
    \new_[75856]_ , \new_[75857]_ , \new_[75861]_ , \new_[75862]_ ,
    \new_[75865]_ , \new_[75868]_ , \new_[75869]_ , \new_[75870]_ ,
    \new_[75874]_ , \new_[75875]_ , \new_[75878]_ , \new_[75881]_ ,
    \new_[75882]_ , \new_[75883]_ , \new_[75887]_ , \new_[75888]_ ,
    \new_[75891]_ , \new_[75894]_ , \new_[75895]_ , \new_[75896]_ ,
    \new_[75900]_ , \new_[75901]_ , \new_[75904]_ , \new_[75907]_ ,
    \new_[75908]_ , \new_[75909]_ , \new_[75913]_ , \new_[75914]_ ,
    \new_[75917]_ , \new_[75920]_ , \new_[75921]_ , \new_[75922]_ ,
    \new_[75926]_ , \new_[75927]_ , \new_[75930]_ , \new_[75933]_ ,
    \new_[75934]_ , \new_[75935]_ , \new_[75939]_ , \new_[75940]_ ,
    \new_[75943]_ , \new_[75946]_ , \new_[75947]_ , \new_[75948]_ ,
    \new_[75952]_ , \new_[75953]_ , \new_[75956]_ , \new_[75959]_ ,
    \new_[75960]_ , \new_[75961]_ , \new_[75965]_ , \new_[75966]_ ,
    \new_[75969]_ , \new_[75972]_ , \new_[75973]_ , \new_[75974]_ ,
    \new_[75978]_ , \new_[75979]_ , \new_[75982]_ , \new_[75985]_ ,
    \new_[75986]_ , \new_[75987]_ , \new_[75991]_ , \new_[75992]_ ,
    \new_[75995]_ , \new_[75998]_ , \new_[75999]_ , \new_[76000]_ ,
    \new_[76004]_ , \new_[76005]_ , \new_[76008]_ , \new_[76011]_ ,
    \new_[76012]_ , \new_[76013]_ , \new_[76017]_ , \new_[76018]_ ,
    \new_[76021]_ , \new_[76024]_ , \new_[76025]_ , \new_[76026]_ ,
    \new_[76030]_ , \new_[76031]_ , \new_[76034]_ , \new_[76037]_ ,
    \new_[76038]_ , \new_[76039]_ , \new_[76043]_ , \new_[76044]_ ,
    \new_[76047]_ , \new_[76050]_ , \new_[76051]_ , \new_[76052]_ ,
    \new_[76056]_ , \new_[76057]_ , \new_[76060]_ , \new_[76063]_ ,
    \new_[76064]_ , \new_[76065]_ , \new_[76069]_ , \new_[76070]_ ,
    \new_[76073]_ , \new_[76076]_ , \new_[76077]_ , \new_[76078]_ ,
    \new_[76082]_ , \new_[76083]_ , \new_[76086]_ , \new_[76089]_ ,
    \new_[76090]_ , \new_[76091]_ , \new_[76095]_ , \new_[76096]_ ,
    \new_[76099]_ , \new_[76102]_ , \new_[76103]_ , \new_[76104]_ ,
    \new_[76108]_ , \new_[76109]_ , \new_[76112]_ , \new_[76115]_ ,
    \new_[76116]_ , \new_[76117]_ , \new_[76121]_ , \new_[76122]_ ,
    \new_[76125]_ , \new_[76128]_ , \new_[76129]_ , \new_[76130]_ ,
    \new_[76134]_ , \new_[76135]_ , \new_[76138]_ , \new_[76141]_ ,
    \new_[76142]_ , \new_[76143]_ , \new_[76147]_ , \new_[76148]_ ,
    \new_[76151]_ , \new_[76154]_ , \new_[76155]_ , \new_[76156]_ ,
    \new_[76160]_ , \new_[76161]_ , \new_[76164]_ , \new_[76167]_ ,
    \new_[76168]_ , \new_[76169]_ , \new_[76173]_ , \new_[76174]_ ,
    \new_[76177]_ , \new_[76180]_ , \new_[76181]_ , \new_[76182]_ ,
    \new_[76186]_ , \new_[76187]_ , \new_[76190]_ , \new_[76193]_ ,
    \new_[76194]_ , \new_[76195]_ , \new_[76199]_ , \new_[76200]_ ,
    \new_[76203]_ , \new_[76206]_ , \new_[76207]_ , \new_[76208]_ ,
    \new_[76212]_ , \new_[76213]_ , \new_[76216]_ , \new_[76219]_ ,
    \new_[76220]_ , \new_[76221]_ , \new_[76225]_ , \new_[76226]_ ,
    \new_[76229]_ , \new_[76232]_ , \new_[76233]_ , \new_[76234]_ ,
    \new_[76238]_ , \new_[76239]_ , \new_[76242]_ , \new_[76245]_ ,
    \new_[76246]_ , \new_[76247]_ , \new_[76251]_ , \new_[76252]_ ,
    \new_[76255]_ , \new_[76258]_ , \new_[76259]_ , \new_[76260]_ ,
    \new_[76264]_ , \new_[76265]_ , \new_[76268]_ , \new_[76271]_ ,
    \new_[76272]_ , \new_[76273]_ , \new_[76277]_ , \new_[76278]_ ,
    \new_[76281]_ , \new_[76284]_ , \new_[76285]_ , \new_[76286]_ ,
    \new_[76290]_ , \new_[76291]_ , \new_[76294]_ , \new_[76297]_ ,
    \new_[76298]_ , \new_[76299]_ , \new_[76303]_ , \new_[76304]_ ,
    \new_[76307]_ , \new_[76310]_ , \new_[76311]_ , \new_[76312]_ ,
    \new_[76316]_ , \new_[76317]_ , \new_[76320]_ , \new_[76323]_ ,
    \new_[76324]_ , \new_[76325]_ , \new_[76329]_ , \new_[76330]_ ,
    \new_[76333]_ , \new_[76336]_ , \new_[76337]_ , \new_[76338]_ ,
    \new_[76342]_ , \new_[76343]_ , \new_[76346]_ , \new_[76349]_ ,
    \new_[76350]_ , \new_[76351]_ , \new_[76355]_ , \new_[76356]_ ,
    \new_[76359]_ , \new_[76362]_ , \new_[76363]_ , \new_[76364]_ ,
    \new_[76368]_ , \new_[76369]_ , \new_[76372]_ , \new_[76375]_ ,
    \new_[76376]_ , \new_[76377]_ , \new_[76381]_ , \new_[76382]_ ,
    \new_[76385]_ , \new_[76388]_ , \new_[76389]_ , \new_[76390]_ ,
    \new_[76394]_ , \new_[76395]_ , \new_[76398]_ , \new_[76401]_ ,
    \new_[76402]_ , \new_[76403]_ , \new_[76407]_ , \new_[76408]_ ,
    \new_[76411]_ , \new_[76414]_ , \new_[76415]_ , \new_[76416]_ ,
    \new_[76420]_ , \new_[76421]_ , \new_[76424]_ , \new_[76427]_ ,
    \new_[76428]_ , \new_[76429]_ , \new_[76433]_ , \new_[76434]_ ,
    \new_[76437]_ , \new_[76440]_ , \new_[76441]_ , \new_[76442]_ ,
    \new_[76446]_ , \new_[76447]_ , \new_[76450]_ , \new_[76453]_ ,
    \new_[76454]_ , \new_[76455]_ , \new_[76459]_ , \new_[76460]_ ,
    \new_[76463]_ , \new_[76466]_ , \new_[76467]_ , \new_[76468]_ ,
    \new_[76472]_ , \new_[76473]_ , \new_[76476]_ , \new_[76479]_ ,
    \new_[76480]_ , \new_[76481]_ , \new_[76485]_ , \new_[76486]_ ,
    \new_[76489]_ , \new_[76492]_ , \new_[76493]_ , \new_[76494]_ ,
    \new_[76498]_ , \new_[76499]_ , \new_[76502]_ , \new_[76505]_ ,
    \new_[76506]_ , \new_[76507]_ , \new_[76511]_ , \new_[76512]_ ,
    \new_[76515]_ , \new_[76518]_ , \new_[76519]_ , \new_[76520]_ ,
    \new_[76524]_ , \new_[76525]_ , \new_[76528]_ , \new_[76531]_ ,
    \new_[76532]_ , \new_[76533]_ , \new_[76537]_ , \new_[76538]_ ,
    \new_[76541]_ , \new_[76544]_ , \new_[76545]_ , \new_[76546]_ ,
    \new_[76550]_ , \new_[76551]_ , \new_[76554]_ , \new_[76557]_ ,
    \new_[76558]_ , \new_[76559]_ , \new_[76563]_ , \new_[76564]_ ,
    \new_[76567]_ , \new_[76570]_ , \new_[76571]_ , \new_[76572]_ ,
    \new_[76576]_ , \new_[76577]_ , \new_[76580]_ , \new_[76583]_ ,
    \new_[76584]_ , \new_[76585]_ , \new_[76589]_ , \new_[76590]_ ,
    \new_[76593]_ , \new_[76596]_ , \new_[76597]_ , \new_[76598]_ ,
    \new_[76602]_ , \new_[76603]_ , \new_[76606]_ , \new_[76609]_ ,
    \new_[76610]_ , \new_[76611]_ , \new_[76615]_ , \new_[76616]_ ,
    \new_[76619]_ , \new_[76622]_ , \new_[76623]_ , \new_[76624]_ ,
    \new_[76628]_ , \new_[76629]_ , \new_[76632]_ , \new_[76635]_ ,
    \new_[76636]_ , \new_[76637]_ , \new_[76641]_ , \new_[76642]_ ,
    \new_[76645]_ , \new_[76648]_ , \new_[76649]_ , \new_[76650]_ ,
    \new_[76654]_ , \new_[76655]_ , \new_[76658]_ , \new_[76661]_ ,
    \new_[76662]_ , \new_[76663]_ , \new_[76667]_ , \new_[76668]_ ,
    \new_[76671]_ , \new_[76674]_ , \new_[76675]_ , \new_[76676]_ ,
    \new_[76680]_ , \new_[76681]_ , \new_[76684]_ , \new_[76687]_ ,
    \new_[76688]_ , \new_[76689]_ , \new_[76693]_ , \new_[76694]_ ,
    \new_[76697]_ , \new_[76700]_ , \new_[76701]_ , \new_[76702]_ ,
    \new_[76706]_ , \new_[76707]_ , \new_[76710]_ , \new_[76713]_ ,
    \new_[76714]_ , \new_[76715]_ , \new_[76719]_ , \new_[76720]_ ,
    \new_[76723]_ , \new_[76726]_ , \new_[76727]_ , \new_[76728]_ ,
    \new_[76732]_ , \new_[76733]_ , \new_[76736]_ , \new_[76739]_ ,
    \new_[76740]_ , \new_[76741]_ , \new_[76745]_ , \new_[76746]_ ,
    \new_[76749]_ , \new_[76752]_ , \new_[76753]_ , \new_[76754]_ ,
    \new_[76758]_ , \new_[76759]_ , \new_[76762]_ , \new_[76765]_ ,
    \new_[76766]_ , \new_[76767]_ , \new_[76771]_ , \new_[76772]_ ,
    \new_[76775]_ , \new_[76778]_ , \new_[76779]_ , \new_[76780]_ ,
    \new_[76784]_ , \new_[76785]_ , \new_[76788]_ , \new_[76791]_ ,
    \new_[76792]_ , \new_[76793]_ , \new_[76797]_ , \new_[76798]_ ,
    \new_[76801]_ , \new_[76804]_ , \new_[76805]_ , \new_[76806]_ ,
    \new_[76810]_ , \new_[76811]_ , \new_[76814]_ , \new_[76817]_ ,
    \new_[76818]_ , \new_[76819]_ , \new_[76823]_ , \new_[76824]_ ,
    \new_[76827]_ , \new_[76830]_ , \new_[76831]_ , \new_[76832]_ ,
    \new_[76836]_ , \new_[76837]_ , \new_[76840]_ , \new_[76843]_ ,
    \new_[76844]_ , \new_[76845]_ , \new_[76849]_ , \new_[76850]_ ,
    \new_[76853]_ , \new_[76856]_ , \new_[76857]_ , \new_[76858]_ ,
    \new_[76862]_ , \new_[76863]_ , \new_[76866]_ , \new_[76869]_ ,
    \new_[76870]_ , \new_[76871]_ , \new_[76875]_ , \new_[76876]_ ,
    \new_[76879]_ , \new_[76882]_ , \new_[76883]_ , \new_[76884]_ ,
    \new_[76888]_ , \new_[76889]_ , \new_[76892]_ , \new_[76895]_ ,
    \new_[76896]_ , \new_[76897]_ , \new_[76901]_ , \new_[76902]_ ,
    \new_[76905]_ , \new_[76908]_ , \new_[76909]_ , \new_[76910]_ ,
    \new_[76914]_ , \new_[76915]_ , \new_[76918]_ , \new_[76921]_ ,
    \new_[76922]_ , \new_[76923]_ , \new_[76927]_ , \new_[76928]_ ,
    \new_[76931]_ , \new_[76934]_ , \new_[76935]_ , \new_[76936]_ ,
    \new_[76940]_ , \new_[76941]_ , \new_[76944]_ , \new_[76947]_ ,
    \new_[76948]_ , \new_[76949]_ , \new_[76953]_ , \new_[76954]_ ,
    \new_[76957]_ , \new_[76960]_ , \new_[76961]_ , \new_[76962]_ ,
    \new_[76966]_ , \new_[76967]_ , \new_[76970]_ , \new_[76973]_ ,
    \new_[76974]_ , \new_[76975]_ , \new_[76979]_ , \new_[76980]_ ,
    \new_[76983]_ , \new_[76986]_ , \new_[76987]_ , \new_[76988]_ ,
    \new_[76992]_ , \new_[76993]_ , \new_[76996]_ , \new_[76999]_ ,
    \new_[77000]_ , \new_[77001]_ , \new_[77005]_ , \new_[77006]_ ,
    \new_[77009]_ , \new_[77012]_ , \new_[77013]_ , \new_[77014]_ ,
    \new_[77018]_ , \new_[77019]_ , \new_[77022]_ , \new_[77025]_ ,
    \new_[77026]_ , \new_[77027]_ , \new_[77031]_ , \new_[77032]_ ,
    \new_[77035]_ , \new_[77038]_ , \new_[77039]_ , \new_[77040]_ ,
    \new_[77044]_ , \new_[77045]_ , \new_[77048]_ , \new_[77051]_ ,
    \new_[77052]_ , \new_[77053]_ , \new_[77057]_ , \new_[77058]_ ,
    \new_[77061]_ , \new_[77064]_ , \new_[77065]_ , \new_[77066]_ ,
    \new_[77070]_ , \new_[77071]_ , \new_[77074]_ , \new_[77077]_ ,
    \new_[77078]_ , \new_[77079]_ , \new_[77083]_ , \new_[77084]_ ,
    \new_[77087]_ , \new_[77090]_ , \new_[77091]_ , \new_[77092]_ ,
    \new_[77096]_ , \new_[77097]_ , \new_[77100]_ , \new_[77103]_ ,
    \new_[77104]_ , \new_[77105]_ , \new_[77109]_ , \new_[77110]_ ,
    \new_[77113]_ , \new_[77116]_ , \new_[77117]_ , \new_[77118]_ ,
    \new_[77122]_ , \new_[77123]_ , \new_[77126]_ , \new_[77129]_ ,
    \new_[77130]_ , \new_[77131]_ , \new_[77135]_ , \new_[77136]_ ,
    \new_[77139]_ , \new_[77142]_ , \new_[77143]_ , \new_[77144]_ ,
    \new_[77148]_ , \new_[77149]_ , \new_[77152]_ , \new_[77155]_ ,
    \new_[77156]_ , \new_[77157]_ , \new_[77161]_ , \new_[77162]_ ,
    \new_[77165]_ , \new_[77168]_ , \new_[77169]_ , \new_[77170]_ ,
    \new_[77174]_ , \new_[77175]_ , \new_[77178]_ , \new_[77181]_ ,
    \new_[77182]_ , \new_[77183]_ , \new_[77187]_ , \new_[77188]_ ,
    \new_[77191]_ , \new_[77194]_ , \new_[77195]_ , \new_[77196]_ ,
    \new_[77200]_ , \new_[77201]_ , \new_[77204]_ , \new_[77207]_ ,
    \new_[77208]_ , \new_[77209]_ , \new_[77213]_ , \new_[77214]_ ,
    \new_[77217]_ , \new_[77220]_ , \new_[77221]_ , \new_[77222]_ ,
    \new_[77226]_ , \new_[77227]_ , \new_[77230]_ , \new_[77233]_ ,
    \new_[77234]_ , \new_[77235]_ , \new_[77239]_ , \new_[77240]_ ,
    \new_[77243]_ , \new_[77246]_ , \new_[77247]_ , \new_[77248]_ ,
    \new_[77252]_ , \new_[77253]_ , \new_[77256]_ , \new_[77259]_ ,
    \new_[77260]_ , \new_[77261]_ , \new_[77265]_ , \new_[77266]_ ,
    \new_[77269]_ , \new_[77272]_ , \new_[77273]_ , \new_[77274]_ ,
    \new_[77278]_ , \new_[77279]_ , \new_[77282]_ , \new_[77285]_ ,
    \new_[77286]_ , \new_[77287]_ , \new_[77291]_ , \new_[77292]_ ,
    \new_[77295]_ , \new_[77298]_ , \new_[77299]_ , \new_[77300]_ ,
    \new_[77304]_ , \new_[77305]_ , \new_[77308]_ , \new_[77311]_ ,
    \new_[77312]_ , \new_[77313]_ , \new_[77317]_ , \new_[77318]_ ,
    \new_[77321]_ , \new_[77324]_ , \new_[77325]_ , \new_[77326]_ ,
    \new_[77330]_ , \new_[77331]_ , \new_[77334]_ , \new_[77337]_ ,
    \new_[77338]_ , \new_[77339]_ , \new_[77343]_ , \new_[77344]_ ,
    \new_[77347]_ , \new_[77350]_ , \new_[77351]_ , \new_[77352]_ ,
    \new_[77356]_ , \new_[77357]_ , \new_[77360]_ , \new_[77363]_ ,
    \new_[77364]_ , \new_[77365]_ , \new_[77369]_ , \new_[77370]_ ,
    \new_[77373]_ , \new_[77376]_ , \new_[77377]_ , \new_[77378]_ ,
    \new_[77382]_ , \new_[77383]_ , \new_[77386]_ , \new_[77389]_ ,
    \new_[77390]_ , \new_[77391]_ , \new_[77395]_ , \new_[77396]_ ,
    \new_[77399]_ , \new_[77402]_ , \new_[77403]_ , \new_[77404]_ ,
    \new_[77408]_ , \new_[77409]_ , \new_[77412]_ , \new_[77415]_ ,
    \new_[77416]_ , \new_[77417]_ , \new_[77421]_ , \new_[77422]_ ,
    \new_[77425]_ , \new_[77428]_ , \new_[77429]_ , \new_[77430]_ ,
    \new_[77434]_ , \new_[77435]_ , \new_[77438]_ , \new_[77441]_ ,
    \new_[77442]_ , \new_[77443]_ , \new_[77447]_ , \new_[77448]_ ,
    \new_[77451]_ , \new_[77454]_ , \new_[77455]_ , \new_[77456]_ ,
    \new_[77460]_ , \new_[77461]_ , \new_[77464]_ , \new_[77467]_ ,
    \new_[77468]_ , \new_[77469]_ , \new_[77473]_ , \new_[77474]_ ,
    \new_[77477]_ , \new_[77480]_ , \new_[77481]_ , \new_[77482]_ ,
    \new_[77486]_ , \new_[77487]_ , \new_[77490]_ , \new_[77493]_ ,
    \new_[77494]_ , \new_[77495]_ , \new_[77499]_ , \new_[77500]_ ,
    \new_[77503]_ , \new_[77506]_ , \new_[77507]_ , \new_[77508]_ ,
    \new_[77512]_ , \new_[77513]_ , \new_[77516]_ , \new_[77519]_ ,
    \new_[77520]_ , \new_[77521]_ , \new_[77525]_ , \new_[77526]_ ,
    \new_[77529]_ , \new_[77532]_ , \new_[77533]_ , \new_[77534]_ ,
    \new_[77538]_ , \new_[77539]_ , \new_[77542]_ , \new_[77545]_ ,
    \new_[77546]_ , \new_[77547]_ , \new_[77551]_ , \new_[77552]_ ,
    \new_[77555]_ , \new_[77558]_ , \new_[77559]_ , \new_[77560]_ ,
    \new_[77564]_ , \new_[77565]_ , \new_[77568]_ , \new_[77571]_ ,
    \new_[77572]_ , \new_[77573]_ , \new_[77577]_ , \new_[77578]_ ,
    \new_[77581]_ , \new_[77584]_ , \new_[77585]_ , \new_[77586]_ ,
    \new_[77590]_ , \new_[77591]_ , \new_[77594]_ , \new_[77597]_ ,
    \new_[77598]_ , \new_[77599]_ , \new_[77603]_ , \new_[77604]_ ,
    \new_[77607]_ , \new_[77610]_ , \new_[77611]_ , \new_[77612]_ ,
    \new_[77616]_ , \new_[77617]_ , \new_[77620]_ , \new_[77623]_ ,
    \new_[77624]_ , \new_[77625]_ , \new_[77629]_ , \new_[77630]_ ,
    \new_[77633]_ , \new_[77636]_ , \new_[77637]_ , \new_[77638]_ ,
    \new_[77642]_ , \new_[77643]_ , \new_[77646]_ , \new_[77649]_ ,
    \new_[77650]_ , \new_[77651]_ , \new_[77655]_ , \new_[77656]_ ,
    \new_[77659]_ , \new_[77662]_ , \new_[77663]_ , \new_[77664]_ ,
    \new_[77668]_ , \new_[77669]_ , \new_[77672]_ , \new_[77675]_ ,
    \new_[77676]_ , \new_[77677]_ , \new_[77681]_ , \new_[77682]_ ,
    \new_[77685]_ , \new_[77688]_ , \new_[77689]_ , \new_[77690]_ ,
    \new_[77694]_ , \new_[77695]_ , \new_[77698]_ , \new_[77701]_ ,
    \new_[77702]_ , \new_[77703]_ , \new_[77707]_ , \new_[77708]_ ,
    \new_[77711]_ , \new_[77714]_ , \new_[77715]_ , \new_[77716]_ ,
    \new_[77720]_ , \new_[77721]_ , \new_[77724]_ , \new_[77727]_ ,
    \new_[77728]_ , \new_[77729]_ , \new_[77733]_ , \new_[77734]_ ,
    \new_[77737]_ , \new_[77740]_ , \new_[77741]_ , \new_[77742]_ ,
    \new_[77746]_ , \new_[77747]_ , \new_[77750]_ , \new_[77753]_ ,
    \new_[77754]_ , \new_[77755]_ , \new_[77759]_ , \new_[77760]_ ,
    \new_[77763]_ , \new_[77766]_ , \new_[77767]_ , \new_[77768]_ ,
    \new_[77772]_ , \new_[77773]_ , \new_[77776]_ , \new_[77779]_ ,
    \new_[77780]_ , \new_[77781]_ , \new_[77785]_ , \new_[77786]_ ,
    \new_[77789]_ , \new_[77792]_ , \new_[77793]_ , \new_[77794]_ ,
    \new_[77798]_ , \new_[77799]_ , \new_[77802]_ , \new_[77805]_ ,
    \new_[77806]_ , \new_[77807]_ , \new_[77811]_ , \new_[77812]_ ,
    \new_[77815]_ , \new_[77818]_ , \new_[77819]_ , \new_[77820]_ ,
    \new_[77824]_ , \new_[77825]_ , \new_[77828]_ , \new_[77831]_ ,
    \new_[77832]_ , \new_[77833]_ , \new_[77837]_ , \new_[77838]_ ,
    \new_[77841]_ , \new_[77844]_ , \new_[77845]_ , \new_[77846]_ ,
    \new_[77850]_ , \new_[77851]_ , \new_[77854]_ , \new_[77857]_ ,
    \new_[77858]_ , \new_[77859]_ , \new_[77863]_ , \new_[77864]_ ,
    \new_[77867]_ , \new_[77870]_ , \new_[77871]_ , \new_[77872]_ ,
    \new_[77876]_ , \new_[77877]_ , \new_[77880]_ , \new_[77883]_ ,
    \new_[77884]_ , \new_[77885]_ , \new_[77889]_ , \new_[77890]_ ,
    \new_[77893]_ , \new_[77896]_ , \new_[77897]_ , \new_[77898]_ ,
    \new_[77902]_ , \new_[77903]_ , \new_[77906]_ , \new_[77909]_ ,
    \new_[77910]_ , \new_[77911]_ , \new_[77915]_ , \new_[77916]_ ,
    \new_[77919]_ , \new_[77922]_ , \new_[77923]_ , \new_[77924]_ ,
    \new_[77928]_ , \new_[77929]_ , \new_[77932]_ , \new_[77935]_ ,
    \new_[77936]_ , \new_[77937]_ , \new_[77941]_ , \new_[77942]_ ,
    \new_[77945]_ , \new_[77948]_ , \new_[77949]_ , \new_[77950]_ ,
    \new_[77954]_ , \new_[77955]_ , \new_[77958]_ , \new_[77961]_ ,
    \new_[77962]_ , \new_[77963]_ , \new_[77967]_ , \new_[77968]_ ,
    \new_[77971]_ , \new_[77974]_ , \new_[77975]_ , \new_[77976]_ ,
    \new_[77980]_ , \new_[77981]_ , \new_[77984]_ , \new_[77987]_ ,
    \new_[77988]_ , \new_[77989]_ , \new_[77993]_ , \new_[77994]_ ,
    \new_[77997]_ , \new_[78000]_ , \new_[78001]_ , \new_[78002]_ ,
    \new_[78006]_ , \new_[78007]_ , \new_[78010]_ , \new_[78013]_ ,
    \new_[78014]_ , \new_[78015]_ , \new_[78019]_ , \new_[78020]_ ,
    \new_[78023]_ , \new_[78026]_ , \new_[78027]_ , \new_[78028]_ ,
    \new_[78032]_ , \new_[78033]_ , \new_[78036]_ , \new_[78039]_ ,
    \new_[78040]_ , \new_[78041]_ , \new_[78045]_ , \new_[78046]_ ,
    \new_[78049]_ , \new_[78052]_ , \new_[78053]_ , \new_[78054]_ ,
    \new_[78058]_ , \new_[78059]_ , \new_[78062]_ , \new_[78065]_ ,
    \new_[78066]_ , \new_[78067]_ , \new_[78071]_ , \new_[78072]_ ,
    \new_[78075]_ , \new_[78078]_ , \new_[78079]_ , \new_[78080]_ ,
    \new_[78084]_ , \new_[78085]_ , \new_[78088]_ , \new_[78091]_ ,
    \new_[78092]_ , \new_[78093]_ , \new_[78097]_ , \new_[78098]_ ,
    \new_[78101]_ , \new_[78104]_ , \new_[78105]_ , \new_[78106]_ ,
    \new_[78110]_ , \new_[78111]_ , \new_[78114]_ , \new_[78117]_ ,
    \new_[78118]_ , \new_[78119]_ , \new_[78123]_ , \new_[78124]_ ,
    \new_[78127]_ , \new_[78130]_ , \new_[78131]_ , \new_[78132]_ ,
    \new_[78136]_ , \new_[78137]_ , \new_[78140]_ , \new_[78143]_ ,
    \new_[78144]_ , \new_[78145]_ , \new_[78149]_ , \new_[78150]_ ,
    \new_[78153]_ , \new_[78156]_ , \new_[78157]_ , \new_[78158]_ ,
    \new_[78162]_ , \new_[78163]_ , \new_[78166]_ , \new_[78169]_ ,
    \new_[78170]_ , \new_[78171]_ , \new_[78175]_ , \new_[78176]_ ,
    \new_[78179]_ , \new_[78182]_ , \new_[78183]_ , \new_[78184]_ ,
    \new_[78188]_ , \new_[78189]_ , \new_[78192]_ , \new_[78195]_ ,
    \new_[78196]_ , \new_[78197]_ , \new_[78201]_ , \new_[78202]_ ,
    \new_[78205]_ , \new_[78208]_ , \new_[78209]_ , \new_[78210]_ ,
    \new_[78214]_ , \new_[78215]_ , \new_[78218]_ , \new_[78221]_ ,
    \new_[78222]_ , \new_[78223]_ , \new_[78227]_ , \new_[78228]_ ,
    \new_[78231]_ , \new_[78234]_ , \new_[78235]_ , \new_[78236]_ ,
    \new_[78240]_ , \new_[78241]_ , \new_[78244]_ , \new_[78247]_ ,
    \new_[78248]_ , \new_[78249]_ , \new_[78253]_ , \new_[78254]_ ,
    \new_[78257]_ , \new_[78260]_ , \new_[78261]_ , \new_[78262]_ ,
    \new_[78266]_ , \new_[78267]_ , \new_[78270]_ , \new_[78273]_ ,
    \new_[78274]_ , \new_[78275]_ , \new_[78279]_ , \new_[78280]_ ,
    \new_[78283]_ , \new_[78286]_ , \new_[78287]_ , \new_[78288]_ ,
    \new_[78292]_ , \new_[78293]_ , \new_[78296]_ , \new_[78299]_ ,
    \new_[78300]_ , \new_[78301]_ , \new_[78305]_ , \new_[78306]_ ,
    \new_[78309]_ , \new_[78312]_ , \new_[78313]_ , \new_[78314]_ ,
    \new_[78318]_ , \new_[78319]_ , \new_[78322]_ , \new_[78325]_ ,
    \new_[78326]_ , \new_[78327]_ , \new_[78331]_ , \new_[78332]_ ,
    \new_[78335]_ , \new_[78338]_ , \new_[78339]_ , \new_[78340]_ ,
    \new_[78344]_ , \new_[78345]_ , \new_[78348]_ , \new_[78351]_ ,
    \new_[78352]_ , \new_[78353]_ , \new_[78357]_ , \new_[78358]_ ,
    \new_[78361]_ , \new_[78364]_ , \new_[78365]_ , \new_[78366]_ ,
    \new_[78370]_ , \new_[78371]_ , \new_[78374]_ , \new_[78377]_ ,
    \new_[78378]_ , \new_[78379]_ , \new_[78383]_ , \new_[78384]_ ,
    \new_[78387]_ , \new_[78390]_ , \new_[78391]_ , \new_[78392]_ ,
    \new_[78396]_ , \new_[78397]_ , \new_[78400]_ , \new_[78403]_ ,
    \new_[78404]_ , \new_[78405]_ , \new_[78409]_ , \new_[78410]_ ,
    \new_[78413]_ , \new_[78416]_ , \new_[78417]_ , \new_[78418]_ ,
    \new_[78422]_ , \new_[78423]_ , \new_[78426]_ , \new_[78429]_ ,
    \new_[78430]_ , \new_[78431]_ , \new_[78435]_ , \new_[78436]_ ,
    \new_[78439]_ , \new_[78442]_ , \new_[78443]_ , \new_[78444]_ ,
    \new_[78448]_ , \new_[78449]_ , \new_[78452]_ , \new_[78455]_ ,
    \new_[78456]_ , \new_[78457]_ , \new_[78461]_ , \new_[78462]_ ,
    \new_[78465]_ , \new_[78468]_ , \new_[78469]_ , \new_[78470]_ ,
    \new_[78474]_ , \new_[78475]_ , \new_[78478]_ , \new_[78481]_ ,
    \new_[78482]_ , \new_[78483]_ , \new_[78487]_ , \new_[78488]_ ,
    \new_[78491]_ , \new_[78494]_ , \new_[78495]_ , \new_[78496]_ ,
    \new_[78500]_ , \new_[78501]_ , \new_[78504]_ , \new_[78507]_ ,
    \new_[78508]_ , \new_[78509]_ , \new_[78513]_ , \new_[78514]_ ,
    \new_[78517]_ , \new_[78520]_ , \new_[78521]_ , \new_[78522]_ ,
    \new_[78526]_ , \new_[78527]_ , \new_[78530]_ , \new_[78533]_ ,
    \new_[78534]_ , \new_[78535]_ , \new_[78539]_ , \new_[78540]_ ,
    \new_[78543]_ , \new_[78546]_ , \new_[78547]_ , \new_[78548]_ ,
    \new_[78552]_ , \new_[78553]_ , \new_[78556]_ , \new_[78559]_ ,
    \new_[78560]_ , \new_[78561]_ , \new_[78565]_ , \new_[78566]_ ,
    \new_[78569]_ , \new_[78572]_ , \new_[78573]_ , \new_[78574]_ ,
    \new_[78578]_ , \new_[78579]_ , \new_[78582]_ , \new_[78585]_ ,
    \new_[78586]_ , \new_[78587]_ , \new_[78591]_ , \new_[78592]_ ,
    \new_[78595]_ , \new_[78598]_ , \new_[78599]_ , \new_[78600]_ ,
    \new_[78604]_ , \new_[78605]_ , \new_[78608]_ , \new_[78611]_ ,
    \new_[78612]_ , \new_[78613]_ , \new_[78617]_ , \new_[78618]_ ,
    \new_[78621]_ , \new_[78624]_ , \new_[78625]_ , \new_[78626]_ ,
    \new_[78630]_ , \new_[78631]_ , \new_[78634]_ , \new_[78637]_ ,
    \new_[78638]_ , \new_[78639]_ , \new_[78643]_ , \new_[78644]_ ,
    \new_[78647]_ , \new_[78650]_ , \new_[78651]_ , \new_[78652]_ ,
    \new_[78656]_ , \new_[78657]_ , \new_[78660]_ , \new_[78663]_ ,
    \new_[78664]_ , \new_[78665]_ , \new_[78669]_ , \new_[78670]_ ,
    \new_[78673]_ , \new_[78676]_ , \new_[78677]_ , \new_[78678]_ ,
    \new_[78682]_ , \new_[78683]_ , \new_[78686]_ , \new_[78689]_ ,
    \new_[78690]_ , \new_[78691]_ , \new_[78695]_ , \new_[78696]_ ,
    \new_[78699]_ , \new_[78702]_ , \new_[78703]_ , \new_[78704]_ ,
    \new_[78708]_ , \new_[78709]_ , \new_[78712]_ , \new_[78715]_ ,
    \new_[78716]_ , \new_[78717]_ , \new_[78721]_ , \new_[78722]_ ,
    \new_[78725]_ , \new_[78728]_ , \new_[78729]_ , \new_[78730]_ ,
    \new_[78734]_ , \new_[78735]_ , \new_[78738]_ , \new_[78741]_ ,
    \new_[78742]_ , \new_[78743]_ , \new_[78747]_ , \new_[78748]_ ,
    \new_[78751]_ , \new_[78754]_ , \new_[78755]_ , \new_[78756]_ ,
    \new_[78760]_ , \new_[78761]_ , \new_[78764]_ , \new_[78767]_ ,
    \new_[78768]_ , \new_[78769]_ , \new_[78773]_ , \new_[78774]_ ,
    \new_[78777]_ , \new_[78780]_ , \new_[78781]_ , \new_[78782]_ ,
    \new_[78786]_ , \new_[78787]_ , \new_[78790]_ , \new_[78793]_ ,
    \new_[78794]_ , \new_[78795]_ , \new_[78799]_ , \new_[78800]_ ,
    \new_[78803]_ , \new_[78806]_ , \new_[78807]_ , \new_[78808]_ ,
    \new_[78812]_ , \new_[78813]_ , \new_[78816]_ , \new_[78819]_ ,
    \new_[78820]_ , \new_[78821]_ , \new_[78825]_ , \new_[78826]_ ,
    \new_[78829]_ , \new_[78832]_ , \new_[78833]_ , \new_[78834]_ ,
    \new_[78838]_ , \new_[78839]_ , \new_[78842]_ , \new_[78845]_ ,
    \new_[78846]_ , \new_[78847]_ , \new_[78851]_ , \new_[78852]_ ,
    \new_[78855]_ , \new_[78858]_ , \new_[78859]_ , \new_[78860]_ ,
    \new_[78864]_ , \new_[78865]_ , \new_[78868]_ , \new_[78871]_ ,
    \new_[78872]_ , \new_[78873]_ , \new_[78877]_ , \new_[78878]_ ,
    \new_[78881]_ , \new_[78884]_ , \new_[78885]_ , \new_[78886]_ ,
    \new_[78890]_ , \new_[78891]_ , \new_[78894]_ , \new_[78897]_ ,
    \new_[78898]_ , \new_[78899]_ , \new_[78903]_ , \new_[78904]_ ,
    \new_[78907]_ , \new_[78910]_ , \new_[78911]_ , \new_[78912]_ ,
    \new_[78916]_ , \new_[78917]_ , \new_[78920]_ , \new_[78923]_ ,
    \new_[78924]_ , \new_[78925]_ , \new_[78929]_ , \new_[78930]_ ,
    \new_[78933]_ , \new_[78936]_ , \new_[78937]_ , \new_[78938]_ ,
    \new_[78942]_ , \new_[78943]_ , \new_[78946]_ , \new_[78949]_ ,
    \new_[78950]_ , \new_[78951]_ , \new_[78955]_ , \new_[78956]_ ,
    \new_[78959]_ , \new_[78962]_ , \new_[78963]_ , \new_[78964]_ ,
    \new_[78968]_ , \new_[78969]_ , \new_[78972]_ , \new_[78975]_ ,
    \new_[78976]_ , \new_[78977]_ , \new_[78981]_ , \new_[78982]_ ,
    \new_[78985]_ , \new_[78988]_ , \new_[78989]_ , \new_[78990]_ ,
    \new_[78994]_ , \new_[78995]_ , \new_[78998]_ , \new_[79001]_ ,
    \new_[79002]_ , \new_[79003]_ , \new_[79007]_ , \new_[79008]_ ,
    \new_[79011]_ , \new_[79014]_ , \new_[79015]_ , \new_[79016]_ ,
    \new_[79020]_ , \new_[79021]_ , \new_[79024]_ , \new_[79027]_ ,
    \new_[79028]_ , \new_[79029]_ , \new_[79033]_ , \new_[79034]_ ,
    \new_[79037]_ , \new_[79040]_ , \new_[79041]_ , \new_[79042]_ ,
    \new_[79046]_ , \new_[79047]_ , \new_[79050]_ , \new_[79053]_ ,
    \new_[79054]_ , \new_[79055]_ , \new_[79059]_ , \new_[79060]_ ,
    \new_[79063]_ , \new_[79066]_ , \new_[79067]_ , \new_[79068]_ ,
    \new_[79072]_ , \new_[79073]_ , \new_[79076]_ , \new_[79079]_ ,
    \new_[79080]_ , \new_[79081]_ , \new_[79085]_ , \new_[79086]_ ,
    \new_[79089]_ , \new_[79092]_ , \new_[79093]_ , \new_[79094]_ ,
    \new_[79098]_ , \new_[79099]_ , \new_[79102]_ , \new_[79105]_ ,
    \new_[79106]_ , \new_[79107]_ , \new_[79111]_ , \new_[79112]_ ,
    \new_[79115]_ , \new_[79118]_ , \new_[79119]_ , \new_[79120]_ ,
    \new_[79124]_ , \new_[79125]_ , \new_[79128]_ , \new_[79131]_ ,
    \new_[79132]_ , \new_[79133]_ , \new_[79137]_ , \new_[79138]_ ,
    \new_[79141]_ , \new_[79144]_ , \new_[79145]_ , \new_[79146]_ ,
    \new_[79150]_ , \new_[79151]_ , \new_[79154]_ , \new_[79157]_ ,
    \new_[79158]_ , \new_[79159]_ , \new_[79163]_ , \new_[79164]_ ,
    \new_[79167]_ , \new_[79170]_ , \new_[79171]_ , \new_[79172]_ ,
    \new_[79176]_ , \new_[79177]_ , \new_[79180]_ , \new_[79183]_ ,
    \new_[79184]_ , \new_[79185]_ , \new_[79189]_ , \new_[79190]_ ,
    \new_[79193]_ , \new_[79196]_ , \new_[79197]_ , \new_[79198]_ ,
    \new_[79202]_ , \new_[79203]_ , \new_[79206]_ , \new_[79209]_ ,
    \new_[79210]_ , \new_[79211]_ , \new_[79215]_ , \new_[79216]_ ,
    \new_[79219]_ , \new_[79222]_ , \new_[79223]_ , \new_[79224]_ ,
    \new_[79228]_ , \new_[79229]_ , \new_[79232]_ , \new_[79235]_ ,
    \new_[79236]_ , \new_[79237]_ , \new_[79241]_ , \new_[79242]_ ,
    \new_[79245]_ , \new_[79248]_ , \new_[79249]_ , \new_[79250]_ ,
    \new_[79254]_ , \new_[79255]_ , \new_[79258]_ , \new_[79261]_ ,
    \new_[79262]_ , \new_[79263]_ , \new_[79267]_ , \new_[79268]_ ,
    \new_[79271]_ , \new_[79274]_ , \new_[79275]_ , \new_[79276]_ ,
    \new_[79280]_ , \new_[79281]_ , \new_[79284]_ , \new_[79287]_ ,
    \new_[79288]_ , \new_[79289]_ , \new_[79293]_ , \new_[79294]_ ,
    \new_[79297]_ , \new_[79300]_ , \new_[79301]_ , \new_[79302]_ ,
    \new_[79306]_ , \new_[79307]_ , \new_[79310]_ , \new_[79313]_ ,
    \new_[79314]_ , \new_[79315]_ , \new_[79319]_ , \new_[79320]_ ,
    \new_[79323]_ , \new_[79326]_ , \new_[79327]_ , \new_[79328]_ ,
    \new_[79332]_ , \new_[79333]_ , \new_[79336]_ , \new_[79339]_ ,
    \new_[79340]_ , \new_[79341]_ , \new_[79345]_ , \new_[79346]_ ,
    \new_[79349]_ , \new_[79352]_ , \new_[79353]_ , \new_[79354]_ ,
    \new_[79358]_ , \new_[79359]_ , \new_[79362]_ , \new_[79365]_ ,
    \new_[79366]_ , \new_[79367]_ , \new_[79371]_ , \new_[79372]_ ,
    \new_[79375]_ , \new_[79378]_ , \new_[79379]_ , \new_[79380]_ ,
    \new_[79384]_ , \new_[79385]_ , \new_[79388]_ , \new_[79391]_ ,
    \new_[79392]_ , \new_[79393]_ , \new_[79397]_ , \new_[79398]_ ,
    \new_[79401]_ , \new_[79404]_ , \new_[79405]_ , \new_[79406]_ ,
    \new_[79410]_ , \new_[79411]_ , \new_[79414]_ , \new_[79417]_ ,
    \new_[79418]_ , \new_[79419]_ , \new_[79423]_ , \new_[79424]_ ,
    \new_[79427]_ , \new_[79430]_ , \new_[79431]_ , \new_[79432]_ ,
    \new_[79436]_ , \new_[79437]_ , \new_[79440]_ , \new_[79443]_ ,
    \new_[79444]_ , \new_[79445]_ , \new_[79449]_ , \new_[79450]_ ,
    \new_[79453]_ , \new_[79456]_ , \new_[79457]_ , \new_[79458]_ ,
    \new_[79462]_ , \new_[79463]_ , \new_[79466]_ , \new_[79469]_ ,
    \new_[79470]_ , \new_[79471]_ , \new_[79475]_ , \new_[79476]_ ,
    \new_[79479]_ , \new_[79482]_ , \new_[79483]_ , \new_[79484]_ ,
    \new_[79488]_ , \new_[79489]_ , \new_[79492]_ , \new_[79495]_ ,
    \new_[79496]_ , \new_[79497]_ , \new_[79501]_ , \new_[79502]_ ,
    \new_[79505]_ , \new_[79508]_ , \new_[79509]_ , \new_[79510]_ ,
    \new_[79514]_ , \new_[79515]_ , \new_[79518]_ , \new_[79521]_ ,
    \new_[79522]_ , \new_[79523]_ , \new_[79527]_ , \new_[79528]_ ,
    \new_[79531]_ , \new_[79534]_ , \new_[79535]_ , \new_[79536]_ ,
    \new_[79540]_ , \new_[79541]_ , \new_[79544]_ , \new_[79547]_ ,
    \new_[79548]_ , \new_[79549]_ , \new_[79553]_ , \new_[79554]_ ,
    \new_[79557]_ , \new_[79560]_ , \new_[79561]_ , \new_[79562]_ ,
    \new_[79566]_ , \new_[79567]_ , \new_[79570]_ , \new_[79573]_ ,
    \new_[79574]_ , \new_[79575]_ , \new_[79579]_ , \new_[79580]_ ,
    \new_[79583]_ , \new_[79586]_ , \new_[79587]_ , \new_[79588]_ ,
    \new_[79592]_ , \new_[79593]_ , \new_[79596]_ , \new_[79599]_ ,
    \new_[79600]_ , \new_[79601]_ , \new_[79605]_ , \new_[79606]_ ,
    \new_[79609]_ , \new_[79612]_ , \new_[79613]_ , \new_[79614]_ ,
    \new_[79618]_ , \new_[79619]_ , \new_[79622]_ , \new_[79625]_ ,
    \new_[79626]_ , \new_[79627]_ , \new_[79631]_ , \new_[79632]_ ,
    \new_[79635]_ , \new_[79638]_ , \new_[79639]_ , \new_[79640]_ ,
    \new_[79644]_ , \new_[79645]_ , \new_[79648]_ , \new_[79651]_ ,
    \new_[79652]_ , \new_[79653]_ , \new_[79657]_ , \new_[79658]_ ,
    \new_[79661]_ , \new_[79664]_ , \new_[79665]_ , \new_[79666]_ ,
    \new_[79670]_ , \new_[79671]_ , \new_[79674]_ , \new_[79677]_ ,
    \new_[79678]_ , \new_[79679]_ , \new_[79683]_ , \new_[79684]_ ,
    \new_[79687]_ , \new_[79690]_ , \new_[79691]_ , \new_[79692]_ ,
    \new_[79696]_ , \new_[79697]_ , \new_[79700]_ , \new_[79703]_ ,
    \new_[79704]_ , \new_[79705]_ , \new_[79709]_ , \new_[79710]_ ,
    \new_[79713]_ , \new_[79716]_ , \new_[79717]_ , \new_[79718]_ ,
    \new_[79722]_ , \new_[79723]_ , \new_[79726]_ , \new_[79729]_ ,
    \new_[79730]_ , \new_[79731]_ , \new_[79735]_ , \new_[79736]_ ,
    \new_[79739]_ , \new_[79742]_ , \new_[79743]_ , \new_[79744]_ ,
    \new_[79748]_ , \new_[79749]_ , \new_[79752]_ , \new_[79755]_ ,
    \new_[79756]_ , \new_[79757]_ , \new_[79761]_ , \new_[79762]_ ,
    \new_[79765]_ , \new_[79768]_ , \new_[79769]_ , \new_[79770]_ ,
    \new_[79774]_ , \new_[79775]_ , \new_[79778]_ , \new_[79781]_ ,
    \new_[79782]_ , \new_[79783]_ , \new_[79787]_ , \new_[79788]_ ,
    \new_[79791]_ , \new_[79794]_ , \new_[79795]_ , \new_[79796]_ ,
    \new_[79800]_ , \new_[79801]_ , \new_[79804]_ , \new_[79807]_ ,
    \new_[79808]_ , \new_[79809]_ , \new_[79813]_ , \new_[79814]_ ,
    \new_[79817]_ , \new_[79820]_ , \new_[79821]_ , \new_[79822]_ ,
    \new_[79826]_ , \new_[79827]_ , \new_[79830]_ , \new_[79833]_ ,
    \new_[79834]_ , \new_[79835]_ , \new_[79839]_ , \new_[79840]_ ,
    \new_[79843]_ , \new_[79846]_ , \new_[79847]_ , \new_[79848]_ ,
    \new_[79852]_ , \new_[79853]_ , \new_[79856]_ , \new_[79859]_ ,
    \new_[79860]_ , \new_[79861]_ , \new_[79865]_ , \new_[79866]_ ,
    \new_[79869]_ , \new_[79872]_ , \new_[79873]_ , \new_[79874]_ ,
    \new_[79878]_ , \new_[79879]_ , \new_[79882]_ , \new_[79885]_ ,
    \new_[79886]_ , \new_[79887]_ , \new_[79891]_ , \new_[79892]_ ,
    \new_[79895]_ , \new_[79898]_ , \new_[79899]_ , \new_[79900]_ ,
    \new_[79904]_ , \new_[79905]_ , \new_[79908]_ , \new_[79911]_ ,
    \new_[79912]_ , \new_[79913]_ , \new_[79917]_ , \new_[79918]_ ,
    \new_[79921]_ , \new_[79924]_ , \new_[79925]_ , \new_[79926]_ ,
    \new_[79930]_ , \new_[79931]_ , \new_[79934]_ , \new_[79937]_ ,
    \new_[79938]_ , \new_[79939]_ , \new_[79943]_ , \new_[79944]_ ,
    \new_[79947]_ , \new_[79950]_ , \new_[79951]_ , \new_[79952]_ ,
    \new_[79956]_ , \new_[79957]_ , \new_[79960]_ , \new_[79963]_ ,
    \new_[79964]_ , \new_[79965]_ , \new_[79969]_ , \new_[79970]_ ,
    \new_[79973]_ , \new_[79976]_ , \new_[79977]_ , \new_[79978]_ ,
    \new_[79982]_ , \new_[79983]_ , \new_[79986]_ , \new_[79989]_ ,
    \new_[79990]_ , \new_[79991]_ , \new_[79995]_ , \new_[79996]_ ,
    \new_[79999]_ , \new_[80002]_ , \new_[80003]_ , \new_[80004]_ ,
    \new_[80008]_ , \new_[80009]_ , \new_[80012]_ , \new_[80015]_ ,
    \new_[80016]_ , \new_[80017]_ , \new_[80021]_ , \new_[80022]_ ,
    \new_[80025]_ , \new_[80028]_ , \new_[80029]_ , \new_[80030]_ ,
    \new_[80034]_ , \new_[80035]_ , \new_[80038]_ , \new_[80041]_ ,
    \new_[80042]_ , \new_[80043]_ , \new_[80047]_ , \new_[80048]_ ,
    \new_[80051]_ , \new_[80054]_ , \new_[80055]_ , \new_[80056]_ ,
    \new_[80060]_ , \new_[80061]_ , \new_[80064]_ , \new_[80067]_ ,
    \new_[80068]_ , \new_[80069]_ , \new_[80073]_ , \new_[80074]_ ,
    \new_[80077]_ , \new_[80080]_ , \new_[80081]_ , \new_[80082]_ ,
    \new_[80086]_ , \new_[80087]_ , \new_[80090]_ , \new_[80093]_ ,
    \new_[80094]_ , \new_[80095]_ , \new_[80099]_ , \new_[80100]_ ,
    \new_[80103]_ , \new_[80106]_ , \new_[80107]_ , \new_[80108]_ ,
    \new_[80112]_ , \new_[80113]_ , \new_[80116]_ , \new_[80119]_ ,
    \new_[80120]_ , \new_[80121]_ , \new_[80125]_ , \new_[80126]_ ,
    \new_[80129]_ , \new_[80132]_ , \new_[80133]_ , \new_[80134]_ ,
    \new_[80138]_ , \new_[80139]_ , \new_[80142]_ , \new_[80145]_ ,
    \new_[80146]_ , \new_[80147]_ , \new_[80151]_ , \new_[80152]_ ,
    \new_[80155]_ , \new_[80158]_ , \new_[80159]_ , \new_[80160]_ ,
    \new_[80164]_ , \new_[80165]_ , \new_[80168]_ , \new_[80171]_ ,
    \new_[80172]_ , \new_[80173]_ , \new_[80177]_ , \new_[80178]_ ,
    \new_[80181]_ , \new_[80184]_ , \new_[80185]_ , \new_[80186]_ ,
    \new_[80190]_ , \new_[80191]_ , \new_[80194]_ , \new_[80197]_ ,
    \new_[80198]_ , \new_[80199]_ , \new_[80203]_ , \new_[80204]_ ,
    \new_[80207]_ , \new_[80210]_ , \new_[80211]_ , \new_[80212]_ ,
    \new_[80216]_ , \new_[80217]_ , \new_[80220]_ , \new_[80223]_ ,
    \new_[80224]_ , \new_[80225]_ , \new_[80229]_ , \new_[80230]_ ,
    \new_[80233]_ , \new_[80236]_ , \new_[80237]_ , \new_[80238]_ ,
    \new_[80242]_ , \new_[80243]_ , \new_[80246]_ , \new_[80249]_ ,
    \new_[80250]_ , \new_[80251]_ , \new_[80255]_ , \new_[80256]_ ,
    \new_[80259]_ , \new_[80262]_ , \new_[80263]_ , \new_[80264]_ ,
    \new_[80268]_ , \new_[80269]_ , \new_[80272]_ , \new_[80275]_ ,
    \new_[80276]_ , \new_[80277]_ , \new_[80281]_ , \new_[80282]_ ,
    \new_[80285]_ , \new_[80288]_ , \new_[80289]_ , \new_[80290]_ ,
    \new_[80294]_ , \new_[80295]_ , \new_[80298]_ , \new_[80301]_ ,
    \new_[80302]_ , \new_[80303]_ , \new_[80307]_ , \new_[80308]_ ,
    \new_[80311]_ , \new_[80314]_ , \new_[80315]_ , \new_[80316]_ ,
    \new_[80320]_ , \new_[80321]_ , \new_[80324]_ , \new_[80327]_ ,
    \new_[80328]_ , \new_[80329]_ , \new_[80333]_ , \new_[80334]_ ,
    \new_[80337]_ , \new_[80340]_ , \new_[80341]_ , \new_[80342]_ ,
    \new_[80346]_ , \new_[80347]_ , \new_[80350]_ , \new_[80353]_ ,
    \new_[80354]_ , \new_[80355]_ , \new_[80359]_ , \new_[80360]_ ,
    \new_[80363]_ , \new_[80366]_ , \new_[80367]_ , \new_[80368]_ ,
    \new_[80372]_ , \new_[80373]_ , \new_[80376]_ , \new_[80379]_ ,
    \new_[80380]_ , \new_[80381]_ , \new_[80385]_ , \new_[80386]_ ,
    \new_[80389]_ , \new_[80392]_ , \new_[80393]_ , \new_[80394]_ ,
    \new_[80398]_ , \new_[80399]_ , \new_[80402]_ , \new_[80405]_ ,
    \new_[80406]_ , \new_[80407]_ , \new_[80411]_ , \new_[80412]_ ,
    \new_[80415]_ , \new_[80418]_ , \new_[80419]_ , \new_[80420]_ ,
    \new_[80424]_ , \new_[80425]_ , \new_[80428]_ , \new_[80431]_ ,
    \new_[80432]_ , \new_[80433]_ , \new_[80437]_ , \new_[80438]_ ,
    \new_[80441]_ , \new_[80444]_ , \new_[80445]_ , \new_[80446]_ ,
    \new_[80450]_ , \new_[80451]_ , \new_[80454]_ , \new_[80457]_ ,
    \new_[80458]_ , \new_[80459]_ , \new_[80463]_ , \new_[80464]_ ,
    \new_[80467]_ , \new_[80470]_ , \new_[80471]_ , \new_[80472]_ ,
    \new_[80476]_ , \new_[80477]_ , \new_[80480]_ , \new_[80483]_ ,
    \new_[80484]_ , \new_[80485]_ , \new_[80489]_ , \new_[80490]_ ,
    \new_[80493]_ , \new_[80496]_ , \new_[80497]_ , \new_[80498]_ ,
    \new_[80502]_ , \new_[80503]_ , \new_[80506]_ , \new_[80509]_ ,
    \new_[80510]_ , \new_[80511]_ , \new_[80515]_ , \new_[80516]_ ,
    \new_[80519]_ , \new_[80522]_ , \new_[80523]_ , \new_[80524]_ ,
    \new_[80528]_ , \new_[80529]_ , \new_[80532]_ , \new_[80535]_ ,
    \new_[80536]_ , \new_[80537]_ , \new_[80541]_ , \new_[80542]_ ,
    \new_[80545]_ , \new_[80548]_ , \new_[80549]_ , \new_[80550]_ ,
    \new_[80554]_ , \new_[80555]_ , \new_[80558]_ , \new_[80561]_ ,
    \new_[80562]_ , \new_[80563]_ , \new_[80567]_ , \new_[80568]_ ,
    \new_[80571]_ , \new_[80574]_ , \new_[80575]_ , \new_[80576]_ ,
    \new_[80580]_ , \new_[80581]_ , \new_[80584]_ , \new_[80587]_ ,
    \new_[80588]_ , \new_[80589]_ , \new_[80593]_ , \new_[80594]_ ,
    \new_[80597]_ , \new_[80600]_ , \new_[80601]_ , \new_[80602]_ ,
    \new_[80606]_ , \new_[80607]_ , \new_[80610]_ , \new_[80613]_ ,
    \new_[80614]_ , \new_[80615]_ , \new_[80619]_ , \new_[80620]_ ,
    \new_[80623]_ , \new_[80626]_ , \new_[80627]_ , \new_[80628]_ ,
    \new_[80632]_ , \new_[80633]_ , \new_[80636]_ , \new_[80639]_ ,
    \new_[80640]_ , \new_[80641]_ , \new_[80645]_ , \new_[80646]_ ,
    \new_[80649]_ , \new_[80652]_ , \new_[80653]_ , \new_[80654]_ ,
    \new_[80658]_ , \new_[80659]_ , \new_[80662]_ , \new_[80665]_ ,
    \new_[80666]_ , \new_[80667]_ , \new_[80671]_ , \new_[80672]_ ,
    \new_[80675]_ , \new_[80678]_ , \new_[80679]_ , \new_[80680]_ ,
    \new_[80684]_ , \new_[80685]_ , \new_[80688]_ , \new_[80691]_ ,
    \new_[80692]_ , \new_[80693]_ , \new_[80697]_ , \new_[80698]_ ,
    \new_[80701]_ , \new_[80704]_ , \new_[80705]_ , \new_[80706]_ ,
    \new_[80710]_ , \new_[80711]_ , \new_[80714]_ , \new_[80717]_ ,
    \new_[80718]_ , \new_[80719]_ , \new_[80723]_ , \new_[80724]_ ,
    \new_[80727]_ , \new_[80730]_ , \new_[80731]_ , \new_[80732]_ ,
    \new_[80736]_ , \new_[80737]_ , \new_[80740]_ , \new_[80743]_ ,
    \new_[80744]_ , \new_[80745]_ , \new_[80749]_ , \new_[80750]_ ,
    \new_[80753]_ , \new_[80756]_ , \new_[80757]_ , \new_[80758]_ ,
    \new_[80762]_ , \new_[80763]_ , \new_[80766]_ , \new_[80769]_ ,
    \new_[80770]_ , \new_[80771]_ , \new_[80775]_ , \new_[80776]_ ,
    \new_[80779]_ , \new_[80782]_ , \new_[80783]_ , \new_[80784]_ ,
    \new_[80788]_ , \new_[80789]_ , \new_[80792]_ , \new_[80795]_ ,
    \new_[80796]_ , \new_[80797]_ , \new_[80801]_ , \new_[80802]_ ,
    \new_[80805]_ , \new_[80808]_ , \new_[80809]_ , \new_[80810]_ ,
    \new_[80814]_ , \new_[80815]_ , \new_[80818]_ , \new_[80821]_ ,
    \new_[80822]_ , \new_[80823]_ , \new_[80827]_ , \new_[80828]_ ,
    \new_[80831]_ , \new_[80834]_ , \new_[80835]_ , \new_[80836]_ ,
    \new_[80840]_ , \new_[80841]_ , \new_[80844]_ , \new_[80847]_ ,
    \new_[80848]_ , \new_[80849]_ , \new_[80853]_ , \new_[80854]_ ,
    \new_[80857]_ , \new_[80860]_ , \new_[80861]_ , \new_[80862]_ ,
    \new_[80866]_ , \new_[80867]_ , \new_[80870]_ , \new_[80873]_ ,
    \new_[80874]_ , \new_[80875]_ , \new_[80879]_ , \new_[80880]_ ,
    \new_[80883]_ , \new_[80886]_ , \new_[80887]_ , \new_[80888]_ ,
    \new_[80892]_ , \new_[80893]_ , \new_[80896]_ , \new_[80899]_ ,
    \new_[80900]_ , \new_[80901]_ , \new_[80905]_ , \new_[80906]_ ,
    \new_[80909]_ , \new_[80912]_ , \new_[80913]_ , \new_[80914]_ ,
    \new_[80918]_ , \new_[80919]_ , \new_[80922]_ , \new_[80925]_ ,
    \new_[80926]_ , \new_[80927]_ , \new_[80931]_ , \new_[80932]_ ,
    \new_[80935]_ , \new_[80938]_ , \new_[80939]_ , \new_[80940]_ ,
    \new_[80944]_ , \new_[80945]_ , \new_[80948]_ , \new_[80951]_ ,
    \new_[80952]_ , \new_[80953]_ , \new_[80957]_ , \new_[80958]_ ,
    \new_[80961]_ , \new_[80964]_ , \new_[80965]_ , \new_[80966]_ ,
    \new_[80970]_ , \new_[80971]_ , \new_[80974]_ , \new_[80977]_ ,
    \new_[80978]_ , \new_[80979]_ , \new_[80983]_ , \new_[80984]_ ,
    \new_[80987]_ , \new_[80990]_ , \new_[80991]_ , \new_[80992]_ ,
    \new_[80996]_ , \new_[80997]_ , \new_[81000]_ , \new_[81003]_ ,
    \new_[81004]_ , \new_[81005]_ , \new_[81009]_ , \new_[81010]_ ,
    \new_[81013]_ , \new_[81016]_ , \new_[81017]_ , \new_[81018]_ ,
    \new_[81022]_ , \new_[81023]_ , \new_[81026]_ , \new_[81029]_ ,
    \new_[81030]_ , \new_[81031]_ , \new_[81035]_ , \new_[81036]_ ,
    \new_[81039]_ , \new_[81042]_ , \new_[81043]_ , \new_[81044]_ ,
    \new_[81048]_ , \new_[81049]_ , \new_[81052]_ , \new_[81055]_ ,
    \new_[81056]_ , \new_[81057]_ , \new_[81061]_ , \new_[81062]_ ,
    \new_[81065]_ , \new_[81068]_ , \new_[81069]_ , \new_[81070]_ ,
    \new_[81074]_ , \new_[81075]_ , \new_[81078]_ , \new_[81081]_ ,
    \new_[81082]_ , \new_[81083]_ , \new_[81087]_ , \new_[81088]_ ,
    \new_[81091]_ , \new_[81094]_ , \new_[81095]_ , \new_[81096]_ ,
    \new_[81100]_ , \new_[81101]_ , \new_[81104]_ , \new_[81107]_ ,
    \new_[81108]_ , \new_[81109]_ , \new_[81113]_ , \new_[81114]_ ,
    \new_[81117]_ , \new_[81120]_ , \new_[81121]_ , \new_[81122]_ ,
    \new_[81126]_ , \new_[81127]_ , \new_[81130]_ , \new_[81133]_ ,
    \new_[81134]_ , \new_[81135]_ , \new_[81139]_ , \new_[81140]_ ,
    \new_[81143]_ , \new_[81146]_ , \new_[81147]_ , \new_[81148]_ ,
    \new_[81152]_ , \new_[81153]_ , \new_[81156]_ , \new_[81159]_ ,
    \new_[81160]_ , \new_[81161]_ , \new_[81165]_ , \new_[81166]_ ,
    \new_[81169]_ , \new_[81172]_ , \new_[81173]_ , \new_[81174]_ ,
    \new_[81178]_ , \new_[81179]_ , \new_[81182]_ , \new_[81185]_ ,
    \new_[81186]_ , \new_[81187]_ , \new_[81191]_ , \new_[81192]_ ,
    \new_[81195]_ , \new_[81198]_ , \new_[81199]_ , \new_[81200]_ ,
    \new_[81204]_ , \new_[81205]_ , \new_[81208]_ , \new_[81211]_ ,
    \new_[81212]_ , \new_[81213]_ , \new_[81217]_ , \new_[81218]_ ,
    \new_[81221]_ , \new_[81224]_ , \new_[81225]_ , \new_[81226]_ ,
    \new_[81230]_ , \new_[81231]_ , \new_[81234]_ , \new_[81237]_ ,
    \new_[81238]_ , \new_[81239]_ , \new_[81243]_ , \new_[81244]_ ,
    \new_[81247]_ , \new_[81250]_ , \new_[81251]_ , \new_[81252]_ ,
    \new_[81256]_ , \new_[81257]_ , \new_[81260]_ , \new_[81263]_ ,
    \new_[81264]_ , \new_[81265]_ , \new_[81269]_ , \new_[81270]_ ,
    \new_[81273]_ , \new_[81276]_ , \new_[81277]_ , \new_[81278]_ ,
    \new_[81282]_ , \new_[81283]_ , \new_[81286]_ , \new_[81289]_ ,
    \new_[81290]_ , \new_[81291]_ , \new_[81295]_ , \new_[81296]_ ,
    \new_[81299]_ , \new_[81302]_ , \new_[81303]_ , \new_[81304]_ ,
    \new_[81308]_ , \new_[81309]_ , \new_[81312]_ , \new_[81315]_ ,
    \new_[81316]_ , \new_[81317]_ , \new_[81321]_ , \new_[81322]_ ,
    \new_[81325]_ , \new_[81328]_ , \new_[81329]_ , \new_[81330]_ ,
    \new_[81334]_ , \new_[81335]_ , \new_[81338]_ , \new_[81341]_ ,
    \new_[81342]_ , \new_[81343]_ , \new_[81347]_ , \new_[81348]_ ,
    \new_[81351]_ , \new_[81354]_ , \new_[81355]_ , \new_[81356]_ ,
    \new_[81360]_ , \new_[81361]_ , \new_[81364]_ , \new_[81367]_ ,
    \new_[81368]_ , \new_[81369]_ , \new_[81373]_ , \new_[81374]_ ,
    \new_[81377]_ , \new_[81380]_ , \new_[81381]_ , \new_[81382]_ ,
    \new_[81386]_ , \new_[81387]_ , \new_[81390]_ , \new_[81393]_ ,
    \new_[81394]_ , \new_[81395]_ , \new_[81399]_ , \new_[81400]_ ,
    \new_[81403]_ , \new_[81406]_ , \new_[81407]_ , \new_[81408]_ ,
    \new_[81412]_ , \new_[81413]_ , \new_[81416]_ , \new_[81419]_ ,
    \new_[81420]_ , \new_[81421]_ , \new_[81425]_ , \new_[81426]_ ,
    \new_[81429]_ , \new_[81432]_ , \new_[81433]_ , \new_[81434]_ ,
    \new_[81438]_ , \new_[81439]_ , \new_[81442]_ , \new_[81445]_ ,
    \new_[81446]_ , \new_[81447]_ , \new_[81451]_ , \new_[81452]_ ,
    \new_[81455]_ , \new_[81458]_ , \new_[81459]_ , \new_[81460]_ ,
    \new_[81464]_ , \new_[81465]_ , \new_[81468]_ , \new_[81471]_ ,
    \new_[81472]_ , \new_[81473]_ , \new_[81477]_ , \new_[81478]_ ,
    \new_[81481]_ , \new_[81484]_ , \new_[81485]_ , \new_[81486]_ ,
    \new_[81490]_ , \new_[81491]_ , \new_[81494]_ , \new_[81497]_ ,
    \new_[81498]_ , \new_[81499]_ , \new_[81503]_ , \new_[81504]_ ,
    \new_[81507]_ , \new_[81510]_ , \new_[81511]_ , \new_[81512]_ ,
    \new_[81516]_ , \new_[81517]_ , \new_[81520]_ , \new_[81523]_ ,
    \new_[81524]_ , \new_[81525]_ , \new_[81529]_ , \new_[81530]_ ,
    \new_[81533]_ , \new_[81536]_ , \new_[81537]_ , \new_[81538]_ ,
    \new_[81542]_ , \new_[81543]_ , \new_[81546]_ , \new_[81549]_ ,
    \new_[81550]_ , \new_[81551]_ , \new_[81555]_ , \new_[81556]_ ,
    \new_[81559]_ , \new_[81562]_ , \new_[81563]_ , \new_[81564]_ ,
    \new_[81568]_ , \new_[81569]_ , \new_[81572]_ , \new_[81575]_ ,
    \new_[81576]_ , \new_[81577]_ , \new_[81581]_ , \new_[81582]_ ,
    \new_[81585]_ , \new_[81588]_ , \new_[81589]_ , \new_[81590]_ ,
    \new_[81594]_ , \new_[81595]_ , \new_[81598]_ , \new_[81601]_ ,
    \new_[81602]_ , \new_[81603]_ , \new_[81607]_ , \new_[81608]_ ,
    \new_[81611]_ , \new_[81614]_ , \new_[81615]_ , \new_[81616]_ ,
    \new_[81620]_ , \new_[81621]_ , \new_[81624]_ , \new_[81627]_ ,
    \new_[81628]_ , \new_[81629]_ , \new_[81633]_ , \new_[81634]_ ,
    \new_[81637]_ , \new_[81640]_ , \new_[81641]_ , \new_[81642]_ ,
    \new_[81646]_ , \new_[81647]_ , \new_[81650]_ , \new_[81653]_ ,
    \new_[81654]_ , \new_[81655]_ , \new_[81659]_ , \new_[81660]_ ,
    \new_[81663]_ , \new_[81666]_ , \new_[81667]_ , \new_[81668]_ ,
    \new_[81672]_ , \new_[81673]_ , \new_[81676]_ , \new_[81679]_ ,
    \new_[81680]_ , \new_[81681]_ , \new_[81685]_ , \new_[81686]_ ,
    \new_[81689]_ , \new_[81692]_ , \new_[81693]_ , \new_[81694]_ ,
    \new_[81698]_ , \new_[81699]_ , \new_[81702]_ , \new_[81705]_ ,
    \new_[81706]_ , \new_[81707]_ , \new_[81711]_ , \new_[81712]_ ,
    \new_[81715]_ , \new_[81718]_ , \new_[81719]_ , \new_[81720]_ ,
    \new_[81724]_ , \new_[81725]_ , \new_[81728]_ , \new_[81731]_ ,
    \new_[81732]_ , \new_[81733]_ , \new_[81737]_ , \new_[81738]_ ,
    \new_[81741]_ , \new_[81744]_ , \new_[81745]_ , \new_[81746]_ ,
    \new_[81750]_ , \new_[81751]_ , \new_[81754]_ , \new_[81757]_ ,
    \new_[81758]_ , \new_[81759]_ , \new_[81763]_ , \new_[81764]_ ,
    \new_[81767]_ , \new_[81770]_ , \new_[81771]_ , \new_[81772]_ ,
    \new_[81776]_ , \new_[81777]_ , \new_[81780]_ , \new_[81783]_ ,
    \new_[81784]_ , \new_[81785]_ , \new_[81789]_ , \new_[81790]_ ,
    \new_[81793]_ , \new_[81796]_ , \new_[81797]_ , \new_[81798]_ ,
    \new_[81802]_ , \new_[81803]_ , \new_[81806]_ , \new_[81809]_ ,
    \new_[81810]_ , \new_[81811]_ , \new_[81815]_ , \new_[81816]_ ,
    \new_[81819]_ , \new_[81822]_ , \new_[81823]_ , \new_[81824]_ ,
    \new_[81828]_ , \new_[81829]_ , \new_[81832]_ , \new_[81835]_ ,
    \new_[81836]_ , \new_[81837]_ , \new_[81841]_ , \new_[81842]_ ,
    \new_[81845]_ , \new_[81848]_ , \new_[81849]_ , \new_[81850]_ ,
    \new_[81854]_ , \new_[81855]_ , \new_[81858]_ , \new_[81861]_ ,
    \new_[81862]_ , \new_[81863]_ , \new_[81867]_ , \new_[81868]_ ,
    \new_[81871]_ , \new_[81874]_ , \new_[81875]_ , \new_[81876]_ ,
    \new_[81880]_ , \new_[81881]_ , \new_[81884]_ , \new_[81887]_ ,
    \new_[81888]_ , \new_[81889]_ , \new_[81893]_ , \new_[81894]_ ,
    \new_[81897]_ , \new_[81900]_ , \new_[81901]_ , \new_[81902]_ ,
    \new_[81906]_ , \new_[81907]_ , \new_[81910]_ , \new_[81913]_ ,
    \new_[81914]_ , \new_[81915]_ , \new_[81919]_ , \new_[81920]_ ,
    \new_[81923]_ , \new_[81926]_ , \new_[81927]_ , \new_[81928]_ ,
    \new_[81932]_ , \new_[81933]_ , \new_[81936]_ , \new_[81939]_ ,
    \new_[81940]_ , \new_[81941]_ , \new_[81945]_ , \new_[81946]_ ,
    \new_[81949]_ , \new_[81952]_ , \new_[81953]_ , \new_[81954]_ ,
    \new_[81958]_ , \new_[81959]_ , \new_[81962]_ , \new_[81965]_ ,
    \new_[81966]_ , \new_[81967]_ , \new_[81971]_ , \new_[81972]_ ,
    \new_[81975]_ , \new_[81978]_ , \new_[81979]_ , \new_[81980]_ ,
    \new_[81984]_ , \new_[81985]_ , \new_[81988]_ , \new_[81991]_ ,
    \new_[81992]_ , \new_[81993]_ , \new_[81997]_ , \new_[81998]_ ,
    \new_[82001]_ , \new_[82004]_ , \new_[82005]_ , \new_[82006]_ ,
    \new_[82010]_ , \new_[82011]_ , \new_[82014]_ , \new_[82017]_ ,
    \new_[82018]_ , \new_[82019]_ , \new_[82023]_ , \new_[82024]_ ,
    \new_[82027]_ , \new_[82030]_ , \new_[82031]_ , \new_[82032]_ ,
    \new_[82036]_ , \new_[82037]_ , \new_[82040]_ , \new_[82043]_ ,
    \new_[82044]_ , \new_[82045]_ , \new_[82049]_ , \new_[82050]_ ,
    \new_[82053]_ , \new_[82056]_ , \new_[82057]_ , \new_[82058]_ ,
    \new_[82062]_ , \new_[82063]_ , \new_[82066]_ , \new_[82069]_ ,
    \new_[82070]_ , \new_[82071]_ , \new_[82075]_ , \new_[82076]_ ,
    \new_[82079]_ , \new_[82082]_ , \new_[82083]_ , \new_[82084]_ ,
    \new_[82088]_ , \new_[82089]_ , \new_[82092]_ , \new_[82095]_ ,
    \new_[82096]_ , \new_[82097]_ , \new_[82101]_ , \new_[82102]_ ,
    \new_[82105]_ , \new_[82108]_ , \new_[82109]_ , \new_[82110]_ ,
    \new_[82114]_ , \new_[82115]_ , \new_[82118]_ , \new_[82121]_ ,
    \new_[82122]_ , \new_[82123]_ , \new_[82127]_ , \new_[82128]_ ,
    \new_[82131]_ , \new_[82134]_ , \new_[82135]_ , \new_[82136]_ ,
    \new_[82140]_ , \new_[82141]_ , \new_[82144]_ , \new_[82147]_ ,
    \new_[82148]_ , \new_[82149]_ , \new_[82153]_ , \new_[82154]_ ,
    \new_[82157]_ , \new_[82160]_ , \new_[82161]_ , \new_[82162]_ ,
    \new_[82166]_ , \new_[82167]_ , \new_[82170]_ , \new_[82173]_ ,
    \new_[82174]_ , \new_[82175]_ , \new_[82179]_ , \new_[82180]_ ,
    \new_[82183]_ , \new_[82186]_ , \new_[82187]_ , \new_[82188]_ ,
    \new_[82192]_ , \new_[82193]_ , \new_[82196]_ , \new_[82199]_ ,
    \new_[82200]_ , \new_[82201]_ , \new_[82205]_ , \new_[82206]_ ,
    \new_[82209]_ , \new_[82212]_ , \new_[82213]_ , \new_[82214]_ ,
    \new_[82218]_ , \new_[82219]_ , \new_[82222]_ , \new_[82225]_ ,
    \new_[82226]_ , \new_[82227]_ , \new_[82231]_ , \new_[82232]_ ,
    \new_[82235]_ , \new_[82238]_ , \new_[82239]_ , \new_[82240]_ ,
    \new_[82244]_ , \new_[82245]_ , \new_[82248]_ , \new_[82251]_ ,
    \new_[82252]_ , \new_[82253]_ , \new_[82257]_ , \new_[82258]_ ,
    \new_[82261]_ , \new_[82264]_ , \new_[82265]_ , \new_[82266]_ ,
    \new_[82270]_ , \new_[82271]_ , \new_[82274]_ , \new_[82277]_ ,
    \new_[82278]_ , \new_[82279]_ , \new_[82283]_ , \new_[82284]_ ,
    \new_[82287]_ , \new_[82290]_ , \new_[82291]_ , \new_[82292]_ ,
    \new_[82296]_ , \new_[82297]_ , \new_[82300]_ , \new_[82303]_ ,
    \new_[82304]_ , \new_[82305]_ , \new_[82309]_ , \new_[82310]_ ,
    \new_[82313]_ , \new_[82316]_ , \new_[82317]_ , \new_[82318]_ ,
    \new_[82322]_ , \new_[82323]_ , \new_[82326]_ , \new_[82329]_ ,
    \new_[82330]_ , \new_[82331]_ , \new_[82335]_ , \new_[82336]_ ,
    \new_[82339]_ , \new_[82342]_ , \new_[82343]_ , \new_[82344]_ ,
    \new_[82348]_ , \new_[82349]_ , \new_[82352]_ , \new_[82355]_ ,
    \new_[82356]_ , \new_[82357]_ , \new_[82361]_ , \new_[82362]_ ,
    \new_[82365]_ , \new_[82368]_ , \new_[82369]_ , \new_[82370]_ ,
    \new_[82374]_ , \new_[82375]_ , \new_[82378]_ , \new_[82381]_ ,
    \new_[82382]_ , \new_[82383]_ , \new_[82387]_ , \new_[82388]_ ,
    \new_[82391]_ , \new_[82394]_ , \new_[82395]_ , \new_[82396]_ ,
    \new_[82400]_ , \new_[82401]_ , \new_[82404]_ , \new_[82407]_ ,
    \new_[82408]_ , \new_[82409]_ , \new_[82413]_ , \new_[82414]_ ,
    \new_[82417]_ , \new_[82420]_ , \new_[82421]_ , \new_[82422]_ ,
    \new_[82426]_ , \new_[82427]_ , \new_[82430]_ , \new_[82433]_ ,
    \new_[82434]_ , \new_[82435]_ , \new_[82439]_ , \new_[82440]_ ,
    \new_[82443]_ , \new_[82446]_ , \new_[82447]_ , \new_[82448]_ ,
    \new_[82452]_ , \new_[82453]_ , \new_[82456]_ , \new_[82459]_ ,
    \new_[82460]_ , \new_[82461]_ , \new_[82465]_ , \new_[82466]_ ,
    \new_[82469]_ , \new_[82472]_ , \new_[82473]_ , \new_[82474]_ ,
    \new_[82478]_ , \new_[82479]_ , \new_[82482]_ , \new_[82485]_ ,
    \new_[82486]_ , \new_[82487]_ , \new_[82491]_ , \new_[82492]_ ,
    \new_[82495]_ , \new_[82498]_ , \new_[82499]_ , \new_[82500]_ ,
    \new_[82504]_ , \new_[82505]_ , \new_[82508]_ , \new_[82511]_ ,
    \new_[82512]_ , \new_[82513]_ , \new_[82517]_ , \new_[82518]_ ,
    \new_[82521]_ , \new_[82524]_ , \new_[82525]_ , \new_[82526]_ ,
    \new_[82530]_ , \new_[82531]_ , \new_[82534]_ , \new_[82537]_ ,
    \new_[82538]_ , \new_[82539]_ , \new_[82543]_ , \new_[82544]_ ,
    \new_[82547]_ , \new_[82550]_ , \new_[82551]_ , \new_[82552]_ ,
    \new_[82556]_ , \new_[82557]_ , \new_[82560]_ , \new_[82563]_ ,
    \new_[82564]_ , \new_[82565]_ , \new_[82569]_ , \new_[82570]_ ,
    \new_[82573]_ , \new_[82576]_ , \new_[82577]_ , \new_[82578]_ ,
    \new_[82582]_ , \new_[82583]_ , \new_[82586]_ , \new_[82589]_ ,
    \new_[82590]_ , \new_[82591]_ , \new_[82595]_ , \new_[82596]_ ,
    \new_[82599]_ , \new_[82602]_ , \new_[82603]_ , \new_[82604]_ ,
    \new_[82608]_ , \new_[82609]_ , \new_[82612]_ , \new_[82615]_ ,
    \new_[82616]_ , \new_[82617]_ , \new_[82621]_ , \new_[82622]_ ,
    \new_[82625]_ , \new_[82628]_ , \new_[82629]_ , \new_[82630]_ ,
    \new_[82634]_ , \new_[82635]_ , \new_[82638]_ , \new_[82641]_ ,
    \new_[82642]_ , \new_[82643]_ , \new_[82647]_ , \new_[82648]_ ,
    \new_[82651]_ , \new_[82654]_ , \new_[82655]_ , \new_[82656]_ ,
    \new_[82660]_ , \new_[82661]_ , \new_[82664]_ , \new_[82667]_ ,
    \new_[82668]_ , \new_[82669]_ , \new_[82673]_ , \new_[82674]_ ,
    \new_[82677]_ , \new_[82680]_ , \new_[82681]_ , \new_[82682]_ ,
    \new_[82686]_ , \new_[82687]_ , \new_[82690]_ , \new_[82693]_ ,
    \new_[82694]_ , \new_[82695]_ , \new_[82699]_ , \new_[82700]_ ,
    \new_[82703]_ , \new_[82706]_ , \new_[82707]_ , \new_[82708]_ ,
    \new_[82712]_ , \new_[82713]_ , \new_[82716]_ , \new_[82719]_ ,
    \new_[82720]_ , \new_[82721]_ , \new_[82725]_ , \new_[82726]_ ,
    \new_[82729]_ , \new_[82732]_ , \new_[82733]_ , \new_[82734]_ ,
    \new_[82738]_ , \new_[82739]_ , \new_[82742]_ , \new_[82745]_ ,
    \new_[82746]_ , \new_[82747]_ , \new_[82751]_ , \new_[82752]_ ,
    \new_[82755]_ , \new_[82758]_ , \new_[82759]_ , \new_[82760]_ ,
    \new_[82764]_ , \new_[82765]_ , \new_[82768]_ , \new_[82771]_ ,
    \new_[82772]_ , \new_[82773]_ , \new_[82777]_ , \new_[82778]_ ,
    \new_[82781]_ , \new_[82784]_ , \new_[82785]_ , \new_[82786]_ ,
    \new_[82790]_ , \new_[82791]_ , \new_[82794]_ , \new_[82797]_ ,
    \new_[82798]_ , \new_[82799]_ , \new_[82803]_ , \new_[82804]_ ,
    \new_[82807]_ , \new_[82810]_ , \new_[82811]_ , \new_[82812]_ ,
    \new_[82816]_ , \new_[82817]_ , \new_[82820]_ , \new_[82823]_ ,
    \new_[82824]_ , \new_[82825]_ , \new_[82829]_ , \new_[82830]_ ,
    \new_[82833]_ , \new_[82836]_ , \new_[82837]_ , \new_[82838]_ ,
    \new_[82842]_ , \new_[82843]_ , \new_[82846]_ , \new_[82849]_ ,
    \new_[82850]_ , \new_[82851]_ , \new_[82855]_ , \new_[82856]_ ,
    \new_[82859]_ , \new_[82862]_ , \new_[82863]_ , \new_[82864]_ ,
    \new_[82868]_ , \new_[82869]_ , \new_[82872]_ , \new_[82875]_ ,
    \new_[82876]_ , \new_[82877]_ , \new_[82881]_ , \new_[82882]_ ,
    \new_[82885]_ , \new_[82888]_ , \new_[82889]_ , \new_[82890]_ ,
    \new_[82894]_ , \new_[82895]_ , \new_[82898]_ , \new_[82901]_ ,
    \new_[82902]_ , \new_[82903]_ , \new_[82907]_ , \new_[82908]_ ,
    \new_[82911]_ , \new_[82914]_ , \new_[82915]_ , \new_[82916]_ ,
    \new_[82920]_ , \new_[82921]_ , \new_[82924]_ , \new_[82927]_ ,
    \new_[82928]_ , \new_[82929]_ , \new_[82933]_ , \new_[82934]_ ,
    \new_[82937]_ , \new_[82940]_ , \new_[82941]_ , \new_[82942]_ ,
    \new_[82946]_ , \new_[82947]_ , \new_[82950]_ , \new_[82953]_ ,
    \new_[82954]_ , \new_[82955]_ , \new_[82959]_ , \new_[82960]_ ,
    \new_[82963]_ , \new_[82966]_ , \new_[82967]_ , \new_[82968]_ ,
    \new_[82972]_ , \new_[82973]_ , \new_[82976]_ , \new_[82979]_ ,
    \new_[82980]_ , \new_[82981]_ , \new_[82985]_ , \new_[82986]_ ,
    \new_[82989]_ , \new_[82992]_ , \new_[82993]_ , \new_[82994]_ ,
    \new_[82998]_ , \new_[82999]_ , \new_[83002]_ , \new_[83005]_ ,
    \new_[83006]_ , \new_[83007]_ , \new_[83011]_ , \new_[83012]_ ,
    \new_[83015]_ , \new_[83018]_ , \new_[83019]_ , \new_[83020]_ ,
    \new_[83024]_ , \new_[83025]_ , \new_[83028]_ , \new_[83031]_ ,
    \new_[83032]_ , \new_[83033]_ , \new_[83037]_ , \new_[83038]_ ,
    \new_[83041]_ , \new_[83044]_ , \new_[83045]_ , \new_[83046]_ ,
    \new_[83050]_ , \new_[83051]_ , \new_[83054]_ , \new_[83057]_ ,
    \new_[83058]_ , \new_[83059]_ , \new_[83063]_ , \new_[83064]_ ,
    \new_[83067]_ , \new_[83070]_ , \new_[83071]_ , \new_[83072]_ ,
    \new_[83076]_ , \new_[83077]_ , \new_[83080]_ , \new_[83083]_ ,
    \new_[83084]_ , \new_[83085]_ , \new_[83089]_ , \new_[83090]_ ,
    \new_[83093]_ , \new_[83096]_ , \new_[83097]_ , \new_[83098]_ ,
    \new_[83102]_ , \new_[83103]_ , \new_[83106]_ , \new_[83109]_ ,
    \new_[83110]_ , \new_[83111]_ , \new_[83115]_ , \new_[83116]_ ,
    \new_[83119]_ , \new_[83122]_ , \new_[83123]_ , \new_[83124]_ ,
    \new_[83128]_ , \new_[83129]_ , \new_[83132]_ , \new_[83135]_ ,
    \new_[83136]_ , \new_[83137]_ , \new_[83141]_ , \new_[83142]_ ,
    \new_[83145]_ , \new_[83148]_ , \new_[83149]_ , \new_[83150]_ ,
    \new_[83154]_ , \new_[83155]_ , \new_[83158]_ , \new_[83161]_ ,
    \new_[83162]_ , \new_[83163]_ , \new_[83167]_ , \new_[83168]_ ,
    \new_[83171]_ , \new_[83174]_ , \new_[83175]_ , \new_[83176]_ ,
    \new_[83180]_ , \new_[83181]_ , \new_[83184]_ , \new_[83187]_ ,
    \new_[83188]_ , \new_[83189]_ , \new_[83193]_ , \new_[83194]_ ,
    \new_[83197]_ , \new_[83200]_ , \new_[83201]_ , \new_[83202]_ ,
    \new_[83206]_ , \new_[83207]_ , \new_[83210]_ , \new_[83213]_ ,
    \new_[83214]_ , \new_[83215]_ , \new_[83219]_ , \new_[83220]_ ,
    \new_[83223]_ , \new_[83226]_ , \new_[83227]_ , \new_[83228]_ ,
    \new_[83232]_ , \new_[83233]_ , \new_[83236]_ , \new_[83239]_ ,
    \new_[83240]_ , \new_[83241]_ , \new_[83245]_ , \new_[83246]_ ,
    \new_[83249]_ , \new_[83252]_ , \new_[83253]_ , \new_[83254]_ ,
    \new_[83258]_ , \new_[83259]_ , \new_[83262]_ , \new_[83265]_ ,
    \new_[83266]_ , \new_[83267]_ , \new_[83271]_ , \new_[83272]_ ,
    \new_[83275]_ , \new_[83278]_ , \new_[83279]_ , \new_[83280]_ ,
    \new_[83284]_ , \new_[83285]_ , \new_[83288]_ , \new_[83291]_ ,
    \new_[83292]_ , \new_[83293]_ , \new_[83297]_ , \new_[83298]_ ,
    \new_[83301]_ , \new_[83304]_ , \new_[83305]_ , \new_[83306]_ ,
    \new_[83310]_ , \new_[83311]_ , \new_[83314]_ , \new_[83317]_ ,
    \new_[83318]_ , \new_[83319]_ , \new_[83323]_ , \new_[83324]_ ,
    \new_[83327]_ , \new_[83330]_ , \new_[83331]_ , \new_[83332]_ ,
    \new_[83336]_ , \new_[83337]_ , \new_[83340]_ , \new_[83343]_ ,
    \new_[83344]_ , \new_[83345]_ , \new_[83349]_ , \new_[83350]_ ,
    \new_[83353]_ , \new_[83356]_ , \new_[83357]_ , \new_[83358]_ ,
    \new_[83362]_ , \new_[83363]_ , \new_[83366]_ , \new_[83369]_ ,
    \new_[83370]_ , \new_[83371]_ , \new_[83375]_ , \new_[83376]_ ,
    \new_[83379]_ , \new_[83382]_ , \new_[83383]_ , \new_[83384]_ ,
    \new_[83388]_ , \new_[83389]_ , \new_[83392]_ , \new_[83395]_ ,
    \new_[83396]_ , \new_[83397]_ , \new_[83401]_ , \new_[83402]_ ,
    \new_[83405]_ , \new_[83408]_ , \new_[83409]_ , \new_[83410]_ ,
    \new_[83414]_ , \new_[83415]_ , \new_[83418]_ , \new_[83421]_ ,
    \new_[83422]_ , \new_[83423]_ , \new_[83427]_ , \new_[83428]_ ,
    \new_[83431]_ , \new_[83434]_ , \new_[83435]_ , \new_[83436]_ ,
    \new_[83440]_ , \new_[83441]_ , \new_[83444]_ , \new_[83447]_ ,
    \new_[83448]_ , \new_[83449]_ , \new_[83453]_ , \new_[83454]_ ,
    \new_[83457]_ , \new_[83460]_ , \new_[83461]_ , \new_[83462]_ ,
    \new_[83466]_ , \new_[83467]_ , \new_[83470]_ , \new_[83473]_ ,
    \new_[83474]_ , \new_[83475]_ , \new_[83479]_ , \new_[83480]_ ,
    \new_[83483]_ , \new_[83486]_ , \new_[83487]_ , \new_[83488]_ ,
    \new_[83492]_ , \new_[83493]_ , \new_[83496]_ , \new_[83499]_ ,
    \new_[83500]_ , \new_[83501]_ , \new_[83505]_ , \new_[83506]_ ,
    \new_[83509]_ , \new_[83512]_ , \new_[83513]_ , \new_[83514]_ ,
    \new_[83518]_ , \new_[83519]_ , \new_[83522]_ , \new_[83525]_ ,
    \new_[83526]_ , \new_[83527]_ , \new_[83531]_ , \new_[83532]_ ,
    \new_[83535]_ , \new_[83538]_ , \new_[83539]_ , \new_[83540]_ ,
    \new_[83544]_ , \new_[83545]_ , \new_[83548]_ , \new_[83551]_ ,
    \new_[83552]_ , \new_[83553]_ , \new_[83557]_ , \new_[83558]_ ,
    \new_[83561]_ , \new_[83564]_ , \new_[83565]_ , \new_[83566]_ ,
    \new_[83570]_ , \new_[83571]_ , \new_[83574]_ , \new_[83577]_ ,
    \new_[83578]_ , \new_[83579]_ , \new_[83583]_ , \new_[83584]_ ,
    \new_[83587]_ , \new_[83590]_ , \new_[83591]_ , \new_[83592]_ ,
    \new_[83596]_ , \new_[83597]_ , \new_[83600]_ , \new_[83603]_ ,
    \new_[83604]_ , \new_[83605]_ , \new_[83609]_ , \new_[83610]_ ,
    \new_[83613]_ , \new_[83616]_ , \new_[83617]_ , \new_[83618]_ ,
    \new_[83622]_ , \new_[83623]_ , \new_[83626]_ , \new_[83629]_ ,
    \new_[83630]_ , \new_[83631]_ , \new_[83635]_ , \new_[83636]_ ,
    \new_[83639]_ , \new_[83642]_ , \new_[83643]_ , \new_[83644]_ ,
    \new_[83648]_ , \new_[83649]_ , \new_[83652]_ , \new_[83655]_ ,
    \new_[83656]_ , \new_[83657]_ , \new_[83661]_ , \new_[83662]_ ,
    \new_[83665]_ , \new_[83668]_ , \new_[83669]_ , \new_[83670]_ ,
    \new_[83674]_ , \new_[83675]_ , \new_[83678]_ , \new_[83681]_ ,
    \new_[83682]_ , \new_[83683]_ , \new_[83687]_ , \new_[83688]_ ,
    \new_[83691]_ , \new_[83694]_ , \new_[83695]_ , \new_[83696]_ ,
    \new_[83700]_ , \new_[83701]_ , \new_[83704]_ , \new_[83707]_ ,
    \new_[83708]_ , \new_[83709]_ , \new_[83713]_ , \new_[83714]_ ,
    \new_[83717]_ , \new_[83720]_ , \new_[83721]_ , \new_[83722]_ ,
    \new_[83726]_ , \new_[83727]_ , \new_[83730]_ , \new_[83733]_ ,
    \new_[83734]_ , \new_[83735]_ , \new_[83739]_ , \new_[83740]_ ,
    \new_[83743]_ , \new_[83746]_ , \new_[83747]_ , \new_[83748]_ ,
    \new_[83752]_ , \new_[83753]_ , \new_[83756]_ , \new_[83759]_ ,
    \new_[83760]_ , \new_[83761]_ , \new_[83765]_ , \new_[83766]_ ,
    \new_[83769]_ , \new_[83772]_ , \new_[83773]_ , \new_[83774]_ ,
    \new_[83778]_ , \new_[83779]_ , \new_[83782]_ , \new_[83785]_ ,
    \new_[83786]_ , \new_[83787]_ , \new_[83791]_ , \new_[83792]_ ,
    \new_[83795]_ , \new_[83798]_ , \new_[83799]_ , \new_[83800]_ ,
    \new_[83804]_ , \new_[83805]_ , \new_[83808]_ , \new_[83811]_ ,
    \new_[83812]_ , \new_[83813]_ , \new_[83817]_ , \new_[83818]_ ,
    \new_[83821]_ , \new_[83824]_ , \new_[83825]_ , \new_[83826]_ ,
    \new_[83830]_ , \new_[83831]_ , \new_[83834]_ , \new_[83837]_ ,
    \new_[83838]_ , \new_[83839]_ , \new_[83843]_ , \new_[83844]_ ,
    \new_[83847]_ , \new_[83850]_ , \new_[83851]_ , \new_[83852]_ ,
    \new_[83856]_ , \new_[83857]_ , \new_[83860]_ , \new_[83863]_ ,
    \new_[83864]_ , \new_[83865]_ , \new_[83869]_ , \new_[83870]_ ,
    \new_[83873]_ , \new_[83876]_ , \new_[83877]_ , \new_[83878]_ ,
    \new_[83882]_ , \new_[83883]_ , \new_[83886]_ , \new_[83889]_ ,
    \new_[83890]_ , \new_[83891]_ , \new_[83895]_ , \new_[83896]_ ,
    \new_[83899]_ , \new_[83902]_ , \new_[83903]_ , \new_[83904]_ ,
    \new_[83908]_ , \new_[83909]_ , \new_[83912]_ , \new_[83915]_ ,
    \new_[83916]_ , \new_[83917]_ , \new_[83921]_ , \new_[83922]_ ,
    \new_[83925]_ , \new_[83928]_ , \new_[83929]_ , \new_[83930]_ ,
    \new_[83934]_ , \new_[83935]_ , \new_[83938]_ , \new_[83941]_ ,
    \new_[83942]_ , \new_[83943]_ , \new_[83947]_ , \new_[83948]_ ,
    \new_[83951]_ , \new_[83954]_ , \new_[83955]_ , \new_[83956]_ ,
    \new_[83960]_ , \new_[83961]_ , \new_[83964]_ , \new_[83967]_ ,
    \new_[83968]_ , \new_[83969]_ , \new_[83973]_ , \new_[83974]_ ,
    \new_[83977]_ , \new_[83980]_ , \new_[83981]_ , \new_[83982]_ ,
    \new_[83986]_ , \new_[83987]_ , \new_[83990]_ , \new_[83993]_ ,
    \new_[83994]_ , \new_[83995]_ , \new_[83999]_ , \new_[84000]_ ,
    \new_[84003]_ , \new_[84006]_ , \new_[84007]_ , \new_[84008]_ ,
    \new_[84012]_ , \new_[84013]_ , \new_[84016]_ , \new_[84019]_ ,
    \new_[84020]_ , \new_[84021]_ , \new_[84025]_ , \new_[84026]_ ,
    \new_[84029]_ , \new_[84032]_ , \new_[84033]_ , \new_[84034]_ ,
    \new_[84038]_ , \new_[84039]_ , \new_[84042]_ , \new_[84045]_ ,
    \new_[84046]_ , \new_[84047]_ , \new_[84051]_ , \new_[84052]_ ,
    \new_[84055]_ , \new_[84058]_ , \new_[84059]_ , \new_[84060]_ ,
    \new_[84064]_ , \new_[84065]_ , \new_[84068]_ , \new_[84071]_ ,
    \new_[84072]_ , \new_[84073]_ , \new_[84077]_ , \new_[84078]_ ,
    \new_[84081]_ , \new_[84084]_ , \new_[84085]_ , \new_[84086]_ ,
    \new_[84090]_ , \new_[84091]_ , \new_[84094]_ , \new_[84097]_ ,
    \new_[84098]_ , \new_[84099]_ , \new_[84103]_ , \new_[84104]_ ,
    \new_[84107]_ , \new_[84110]_ , \new_[84111]_ , \new_[84112]_ ,
    \new_[84116]_ , \new_[84117]_ , \new_[84120]_ , \new_[84123]_ ,
    \new_[84124]_ , \new_[84125]_ , \new_[84129]_ , \new_[84130]_ ,
    \new_[84133]_ , \new_[84136]_ , \new_[84137]_ , \new_[84138]_ ,
    \new_[84142]_ , \new_[84143]_ , \new_[84146]_ , \new_[84149]_ ,
    \new_[84150]_ , \new_[84151]_ , \new_[84155]_ , \new_[84156]_ ,
    \new_[84159]_ , \new_[84162]_ , \new_[84163]_ , \new_[84164]_ ,
    \new_[84168]_ , \new_[84169]_ , \new_[84172]_ , \new_[84175]_ ,
    \new_[84176]_ , \new_[84177]_ , \new_[84181]_ , \new_[84182]_ ,
    \new_[84185]_ , \new_[84188]_ , \new_[84189]_ , \new_[84190]_ ,
    \new_[84194]_ , \new_[84195]_ , \new_[84198]_ , \new_[84201]_ ,
    \new_[84202]_ , \new_[84203]_ , \new_[84207]_ , \new_[84208]_ ,
    \new_[84211]_ , \new_[84214]_ , \new_[84215]_ , \new_[84216]_ ,
    \new_[84220]_ , \new_[84221]_ , \new_[84224]_ , \new_[84227]_ ,
    \new_[84228]_ , \new_[84229]_ , \new_[84233]_ , \new_[84234]_ ,
    \new_[84237]_ , \new_[84240]_ , \new_[84241]_ , \new_[84242]_ ,
    \new_[84246]_ , \new_[84247]_ , \new_[84250]_ , \new_[84253]_ ,
    \new_[84254]_ , \new_[84255]_ , \new_[84259]_ , \new_[84260]_ ,
    \new_[84263]_ , \new_[84266]_ , \new_[84267]_ , \new_[84268]_ ,
    \new_[84272]_ , \new_[84273]_ , \new_[84276]_ , \new_[84279]_ ,
    \new_[84280]_ , \new_[84281]_ , \new_[84285]_ , \new_[84286]_ ,
    \new_[84289]_ , \new_[84292]_ , \new_[84293]_ , \new_[84294]_ ,
    \new_[84298]_ , \new_[84299]_ , \new_[84302]_ , \new_[84305]_ ,
    \new_[84306]_ , \new_[84307]_ , \new_[84311]_ , \new_[84312]_ ,
    \new_[84315]_ , \new_[84318]_ , \new_[84319]_ , \new_[84320]_ ,
    \new_[84324]_ , \new_[84325]_ , \new_[84328]_ , \new_[84331]_ ,
    \new_[84332]_ , \new_[84333]_ , \new_[84337]_ , \new_[84338]_ ,
    \new_[84341]_ , \new_[84344]_ , \new_[84345]_ , \new_[84346]_ ,
    \new_[84350]_ , \new_[84351]_ , \new_[84354]_ , \new_[84357]_ ,
    \new_[84358]_ , \new_[84359]_ , \new_[84363]_ , \new_[84364]_ ,
    \new_[84367]_ , \new_[84370]_ , \new_[84371]_ , \new_[84372]_ ,
    \new_[84376]_ , \new_[84377]_ , \new_[84380]_ , \new_[84383]_ ,
    \new_[84384]_ , \new_[84385]_ , \new_[84389]_ , \new_[84390]_ ,
    \new_[84393]_ , \new_[84396]_ , \new_[84397]_ , \new_[84398]_ ,
    \new_[84402]_ , \new_[84403]_ , \new_[84406]_ , \new_[84409]_ ,
    \new_[84410]_ , \new_[84411]_ , \new_[84415]_ , \new_[84416]_ ,
    \new_[84419]_ , \new_[84422]_ , \new_[84423]_ , \new_[84424]_ ,
    \new_[84428]_ , \new_[84429]_ , \new_[84432]_ , \new_[84435]_ ,
    \new_[84436]_ , \new_[84437]_ , \new_[84441]_ , \new_[84442]_ ,
    \new_[84445]_ , \new_[84448]_ , \new_[84449]_ , \new_[84450]_ ,
    \new_[84454]_ , \new_[84455]_ , \new_[84458]_ , \new_[84461]_ ,
    \new_[84462]_ , \new_[84463]_ , \new_[84467]_ , \new_[84468]_ ,
    \new_[84471]_ , \new_[84474]_ , \new_[84475]_ , \new_[84476]_ ,
    \new_[84480]_ , \new_[84481]_ , \new_[84484]_ , \new_[84487]_ ,
    \new_[84488]_ , \new_[84489]_ , \new_[84493]_ , \new_[84494]_ ,
    \new_[84497]_ , \new_[84500]_ , \new_[84501]_ , \new_[84502]_ ,
    \new_[84506]_ , \new_[84507]_ , \new_[84510]_ , \new_[84513]_ ,
    \new_[84514]_ , \new_[84515]_ , \new_[84519]_ , \new_[84520]_ ,
    \new_[84523]_ , \new_[84526]_ , \new_[84527]_ , \new_[84528]_ ,
    \new_[84532]_ , \new_[84533]_ , \new_[84536]_ , \new_[84539]_ ,
    \new_[84540]_ , \new_[84541]_ , \new_[84545]_ , \new_[84546]_ ,
    \new_[84549]_ , \new_[84552]_ , \new_[84553]_ , \new_[84554]_ ,
    \new_[84558]_ , \new_[84559]_ , \new_[84562]_ , \new_[84565]_ ,
    \new_[84566]_ , \new_[84567]_ , \new_[84571]_ , \new_[84572]_ ,
    \new_[84575]_ , \new_[84578]_ , \new_[84579]_ , \new_[84580]_ ,
    \new_[84584]_ , \new_[84585]_ , \new_[84588]_ , \new_[84591]_ ,
    \new_[84592]_ , \new_[84593]_ , \new_[84597]_ , \new_[84598]_ ,
    \new_[84601]_ , \new_[84604]_ , \new_[84605]_ , \new_[84606]_ ,
    \new_[84610]_ , \new_[84611]_ , \new_[84614]_ , \new_[84617]_ ,
    \new_[84618]_ , \new_[84619]_ , \new_[84623]_ , \new_[84624]_ ,
    \new_[84627]_ , \new_[84630]_ , \new_[84631]_ , \new_[84632]_ ,
    \new_[84636]_ , \new_[84637]_ , \new_[84640]_ , \new_[84643]_ ,
    \new_[84644]_ , \new_[84645]_ , \new_[84649]_ , \new_[84650]_ ,
    \new_[84653]_ , \new_[84656]_ , \new_[84657]_ , \new_[84658]_ ,
    \new_[84662]_ , \new_[84663]_ , \new_[84666]_ , \new_[84669]_ ,
    \new_[84670]_ , \new_[84671]_ , \new_[84675]_ , \new_[84676]_ ,
    \new_[84679]_ , \new_[84682]_ , \new_[84683]_ , \new_[84684]_ ,
    \new_[84688]_ , \new_[84689]_ , \new_[84692]_ , \new_[84695]_ ,
    \new_[84696]_ , \new_[84697]_ , \new_[84701]_ , \new_[84702]_ ,
    \new_[84705]_ , \new_[84708]_ , \new_[84709]_ , \new_[84710]_ ,
    \new_[84714]_ , \new_[84715]_ , \new_[84718]_ , \new_[84721]_ ,
    \new_[84722]_ , \new_[84723]_ , \new_[84727]_ , \new_[84728]_ ,
    \new_[84731]_ , \new_[84734]_ , \new_[84735]_ , \new_[84736]_ ,
    \new_[84740]_ , \new_[84741]_ , \new_[84744]_ , \new_[84747]_ ,
    \new_[84748]_ , \new_[84749]_ , \new_[84753]_ , \new_[84754]_ ,
    \new_[84757]_ , \new_[84760]_ , \new_[84761]_ , \new_[84762]_ ,
    \new_[84766]_ , \new_[84767]_ , \new_[84770]_ , \new_[84773]_ ,
    \new_[84774]_ , \new_[84775]_ , \new_[84779]_ , \new_[84780]_ ,
    \new_[84783]_ , \new_[84786]_ , \new_[84787]_ , \new_[84788]_ ,
    \new_[84792]_ , \new_[84793]_ , \new_[84796]_ , \new_[84799]_ ,
    \new_[84800]_ , \new_[84801]_ , \new_[84805]_ , \new_[84806]_ ,
    \new_[84809]_ , \new_[84812]_ , \new_[84813]_ , \new_[84814]_ ,
    \new_[84818]_ , \new_[84819]_ , \new_[84822]_ , \new_[84825]_ ,
    \new_[84826]_ , \new_[84827]_ , \new_[84831]_ , \new_[84832]_ ,
    \new_[84835]_ , \new_[84838]_ , \new_[84839]_ , \new_[84840]_ ,
    \new_[84844]_ , \new_[84845]_ , \new_[84848]_ , \new_[84851]_ ,
    \new_[84852]_ , \new_[84853]_ , \new_[84857]_ , \new_[84858]_ ,
    \new_[84861]_ , \new_[84864]_ , \new_[84865]_ , \new_[84866]_ ,
    \new_[84870]_ , \new_[84871]_ , \new_[84874]_ , \new_[84877]_ ,
    \new_[84878]_ , \new_[84879]_ , \new_[84883]_ , \new_[84884]_ ,
    \new_[84887]_ , \new_[84890]_ , \new_[84891]_ , \new_[84892]_ ,
    \new_[84896]_ , \new_[84897]_ , \new_[84900]_ , \new_[84903]_ ,
    \new_[84904]_ , \new_[84905]_ , \new_[84909]_ , \new_[84910]_ ,
    \new_[84913]_ , \new_[84916]_ , \new_[84917]_ , \new_[84918]_ ,
    \new_[84922]_ , \new_[84923]_ , \new_[84926]_ , \new_[84929]_ ,
    \new_[84930]_ , \new_[84931]_ , \new_[84935]_ , \new_[84936]_ ,
    \new_[84939]_ , \new_[84942]_ , \new_[84943]_ , \new_[84944]_ ,
    \new_[84948]_ , \new_[84949]_ , \new_[84952]_ , \new_[84955]_ ,
    \new_[84956]_ , \new_[84957]_ , \new_[84961]_ , \new_[84962]_ ,
    \new_[84965]_ , \new_[84968]_ , \new_[84969]_ , \new_[84970]_ ,
    \new_[84974]_ , \new_[84975]_ , \new_[84978]_ , \new_[84981]_ ,
    \new_[84982]_ , \new_[84983]_ , \new_[84987]_ , \new_[84988]_ ,
    \new_[84991]_ , \new_[84994]_ , \new_[84995]_ , \new_[84996]_ ,
    \new_[85000]_ , \new_[85001]_ , \new_[85004]_ , \new_[85007]_ ,
    \new_[85008]_ , \new_[85009]_ , \new_[85013]_ , \new_[85014]_ ,
    \new_[85017]_ , \new_[85020]_ , \new_[85021]_ , \new_[85022]_ ,
    \new_[85026]_ , \new_[85027]_ , \new_[85030]_ , \new_[85033]_ ,
    \new_[85034]_ , \new_[85035]_ , \new_[85039]_ , \new_[85040]_ ,
    \new_[85043]_ , \new_[85046]_ , \new_[85047]_ , \new_[85048]_ ,
    \new_[85052]_ , \new_[85053]_ , \new_[85056]_ , \new_[85059]_ ,
    \new_[85060]_ , \new_[85061]_ , \new_[85065]_ , \new_[85066]_ ,
    \new_[85069]_ , \new_[85072]_ , \new_[85073]_ , \new_[85074]_ ,
    \new_[85078]_ , \new_[85079]_ , \new_[85082]_ , \new_[85085]_ ,
    \new_[85086]_ , \new_[85087]_ , \new_[85091]_ , \new_[85092]_ ,
    \new_[85095]_ , \new_[85098]_ , \new_[85099]_ , \new_[85100]_ ,
    \new_[85104]_ , \new_[85105]_ , \new_[85108]_ , \new_[85111]_ ,
    \new_[85112]_ , \new_[85113]_ , \new_[85117]_ , \new_[85118]_ ,
    \new_[85121]_ , \new_[85124]_ , \new_[85125]_ , \new_[85126]_ ,
    \new_[85130]_ , \new_[85131]_ , \new_[85134]_ , \new_[85137]_ ,
    \new_[85138]_ , \new_[85139]_ , \new_[85143]_ , \new_[85144]_ ,
    \new_[85147]_ , \new_[85150]_ , \new_[85151]_ , \new_[85152]_ ,
    \new_[85156]_ , \new_[85157]_ , \new_[85160]_ , \new_[85163]_ ,
    \new_[85164]_ , \new_[85165]_ , \new_[85169]_ , \new_[85170]_ ,
    \new_[85173]_ , \new_[85176]_ , \new_[85177]_ , \new_[85178]_ ,
    \new_[85182]_ , \new_[85183]_ , \new_[85186]_ , \new_[85189]_ ,
    \new_[85190]_ , \new_[85191]_ , \new_[85195]_ , \new_[85196]_ ,
    \new_[85199]_ , \new_[85202]_ , \new_[85203]_ , \new_[85204]_ ,
    \new_[85208]_ , \new_[85209]_ , \new_[85212]_ , \new_[85215]_ ,
    \new_[85216]_ , \new_[85217]_ , \new_[85221]_ , \new_[85222]_ ,
    \new_[85225]_ , \new_[85228]_ , \new_[85229]_ , \new_[85230]_ ,
    \new_[85234]_ , \new_[85235]_ , \new_[85238]_ , \new_[85241]_ ,
    \new_[85242]_ , \new_[85243]_ , \new_[85247]_ , \new_[85248]_ ,
    \new_[85251]_ , \new_[85254]_ , \new_[85255]_ , \new_[85256]_ ,
    \new_[85260]_ , \new_[85261]_ , \new_[85264]_ , \new_[85267]_ ,
    \new_[85268]_ , \new_[85269]_ , \new_[85273]_ , \new_[85274]_ ,
    \new_[85277]_ , \new_[85280]_ , \new_[85281]_ , \new_[85282]_ ,
    \new_[85286]_ , \new_[85287]_ , \new_[85290]_ , \new_[85293]_ ,
    \new_[85294]_ , \new_[85295]_ , \new_[85299]_ , \new_[85300]_ ,
    \new_[85303]_ , \new_[85306]_ , \new_[85307]_ , \new_[85308]_ ,
    \new_[85312]_ , \new_[85313]_ , \new_[85316]_ , \new_[85319]_ ,
    \new_[85320]_ , \new_[85321]_ , \new_[85325]_ , \new_[85326]_ ,
    \new_[85329]_ , \new_[85332]_ , \new_[85333]_ , \new_[85334]_ ,
    \new_[85338]_ , \new_[85339]_ , \new_[85342]_ , \new_[85345]_ ,
    \new_[85346]_ , \new_[85347]_ , \new_[85351]_ , \new_[85352]_ ,
    \new_[85355]_ , \new_[85358]_ , \new_[85359]_ , \new_[85360]_ ,
    \new_[85364]_ , \new_[85365]_ , \new_[85368]_ , \new_[85371]_ ,
    \new_[85372]_ , \new_[85373]_ , \new_[85377]_ , \new_[85378]_ ,
    \new_[85381]_ , \new_[85384]_ , \new_[85385]_ , \new_[85386]_ ,
    \new_[85390]_ , \new_[85391]_ , \new_[85394]_ , \new_[85397]_ ,
    \new_[85398]_ , \new_[85399]_ , \new_[85403]_ , \new_[85404]_ ,
    \new_[85407]_ , \new_[85410]_ , \new_[85411]_ , \new_[85412]_ ,
    \new_[85416]_ , \new_[85417]_ , \new_[85420]_ , \new_[85423]_ ,
    \new_[85424]_ , \new_[85425]_ , \new_[85429]_ , \new_[85430]_ ,
    \new_[85433]_ , \new_[85436]_ , \new_[85437]_ , \new_[85438]_ ,
    \new_[85442]_ , \new_[85443]_ , \new_[85446]_ , \new_[85449]_ ,
    \new_[85450]_ , \new_[85451]_ , \new_[85455]_ , \new_[85456]_ ,
    \new_[85459]_ , \new_[85462]_ , \new_[85463]_ , \new_[85464]_ ,
    \new_[85468]_ , \new_[85469]_ , \new_[85472]_ , \new_[85475]_ ,
    \new_[85476]_ , \new_[85477]_ , \new_[85481]_ , \new_[85482]_ ,
    \new_[85485]_ , \new_[85488]_ , \new_[85489]_ , \new_[85490]_ ,
    \new_[85494]_ , \new_[85495]_ , \new_[85498]_ , \new_[85501]_ ,
    \new_[85502]_ , \new_[85503]_ , \new_[85507]_ , \new_[85508]_ ,
    \new_[85511]_ , \new_[85514]_ , \new_[85515]_ , \new_[85516]_ ,
    \new_[85520]_ , \new_[85521]_ , \new_[85524]_ , \new_[85527]_ ,
    \new_[85528]_ , \new_[85529]_ , \new_[85533]_ , \new_[85534]_ ,
    \new_[85537]_ , \new_[85540]_ , \new_[85541]_ , \new_[85542]_ ,
    \new_[85546]_ , \new_[85547]_ , \new_[85550]_ , \new_[85553]_ ,
    \new_[85554]_ , \new_[85555]_ , \new_[85559]_ , \new_[85560]_ ,
    \new_[85563]_ , \new_[85566]_ , \new_[85567]_ , \new_[85568]_ ,
    \new_[85572]_ , \new_[85573]_ , \new_[85576]_ , \new_[85579]_ ,
    \new_[85580]_ , \new_[85581]_ , \new_[85585]_ , \new_[85586]_ ,
    \new_[85589]_ , \new_[85592]_ , \new_[85593]_ , \new_[85594]_ ,
    \new_[85598]_ , \new_[85599]_ , \new_[85602]_ , \new_[85605]_ ,
    \new_[85606]_ , \new_[85607]_ , \new_[85611]_ , \new_[85612]_ ,
    \new_[85615]_ , \new_[85618]_ , \new_[85619]_ , \new_[85620]_ ,
    \new_[85624]_ , \new_[85625]_ , \new_[85628]_ , \new_[85631]_ ,
    \new_[85632]_ , \new_[85633]_ , \new_[85637]_ , \new_[85638]_ ,
    \new_[85641]_ , \new_[85644]_ , \new_[85645]_ , \new_[85646]_ ,
    \new_[85650]_ , \new_[85651]_ , \new_[85654]_ , \new_[85657]_ ,
    \new_[85658]_ , \new_[85659]_ , \new_[85663]_ , \new_[85664]_ ,
    \new_[85667]_ , \new_[85670]_ , \new_[85671]_ , \new_[85672]_ ,
    \new_[85676]_ , \new_[85677]_ , \new_[85680]_ , \new_[85683]_ ,
    \new_[85684]_ , \new_[85685]_ , \new_[85689]_ , \new_[85690]_ ,
    \new_[85693]_ , \new_[85696]_ , \new_[85697]_ , \new_[85698]_ ,
    \new_[85702]_ , \new_[85703]_ , \new_[85706]_ , \new_[85709]_ ,
    \new_[85710]_ , \new_[85711]_ , \new_[85715]_ , \new_[85716]_ ,
    \new_[85719]_ , \new_[85722]_ , \new_[85723]_ , \new_[85724]_ ,
    \new_[85728]_ , \new_[85729]_ , \new_[85732]_ , \new_[85735]_ ,
    \new_[85736]_ , \new_[85737]_ , \new_[85741]_ , \new_[85742]_ ,
    \new_[85745]_ , \new_[85748]_ , \new_[85749]_ , \new_[85750]_ ,
    \new_[85754]_ , \new_[85755]_ , \new_[85758]_ , \new_[85761]_ ,
    \new_[85762]_ , \new_[85763]_ , \new_[85767]_ , \new_[85768]_ ,
    \new_[85771]_ , \new_[85774]_ , \new_[85775]_ , \new_[85776]_ ,
    \new_[85780]_ , \new_[85781]_ , \new_[85784]_ , \new_[85787]_ ,
    \new_[85788]_ , \new_[85789]_ , \new_[85793]_ , \new_[85794]_ ,
    \new_[85797]_ , \new_[85800]_ , \new_[85801]_ , \new_[85802]_ ,
    \new_[85806]_ , \new_[85807]_ , \new_[85810]_ , \new_[85813]_ ,
    \new_[85814]_ , \new_[85815]_ , \new_[85819]_ , \new_[85820]_ ,
    \new_[85823]_ , \new_[85826]_ , \new_[85827]_ , \new_[85828]_ ,
    \new_[85832]_ , \new_[85833]_ , \new_[85836]_ , \new_[85839]_ ,
    \new_[85840]_ , \new_[85841]_ , \new_[85845]_ , \new_[85846]_ ,
    \new_[85849]_ , \new_[85852]_ , \new_[85853]_ , \new_[85854]_ ,
    \new_[85858]_ , \new_[85859]_ , \new_[85862]_ , \new_[85865]_ ,
    \new_[85866]_ , \new_[85867]_ , \new_[85871]_ , \new_[85872]_ ,
    \new_[85875]_ , \new_[85878]_ , \new_[85879]_ , \new_[85880]_ ,
    \new_[85884]_ , \new_[85885]_ , \new_[85888]_ , \new_[85891]_ ,
    \new_[85892]_ , \new_[85893]_ , \new_[85897]_ , \new_[85898]_ ,
    \new_[85901]_ , \new_[85904]_ , \new_[85905]_ , \new_[85906]_ ,
    \new_[85910]_ , \new_[85911]_ , \new_[85914]_ , \new_[85917]_ ,
    \new_[85918]_ , \new_[85919]_ , \new_[85923]_ , \new_[85924]_ ,
    \new_[85927]_ , \new_[85930]_ , \new_[85931]_ , \new_[85932]_ ,
    \new_[85936]_ , \new_[85937]_ , \new_[85940]_ , \new_[85943]_ ,
    \new_[85944]_ , \new_[85945]_ , \new_[85949]_ , \new_[85950]_ ,
    \new_[85953]_ , \new_[85956]_ , \new_[85957]_ , \new_[85958]_ ,
    \new_[85962]_ , \new_[85963]_ , \new_[85966]_ , \new_[85969]_ ,
    \new_[85970]_ , \new_[85971]_ , \new_[85975]_ , \new_[85976]_ ,
    \new_[85979]_ , \new_[85982]_ , \new_[85983]_ , \new_[85984]_ ,
    \new_[85988]_ , \new_[85989]_ , \new_[85992]_ , \new_[85995]_ ,
    \new_[85996]_ , \new_[85997]_ , \new_[86001]_ , \new_[86002]_ ,
    \new_[86005]_ , \new_[86008]_ , \new_[86009]_ , \new_[86010]_ ,
    \new_[86014]_ , \new_[86015]_ , \new_[86018]_ , \new_[86021]_ ,
    \new_[86022]_ , \new_[86023]_ , \new_[86027]_ , \new_[86028]_ ,
    \new_[86031]_ , \new_[86034]_ , \new_[86035]_ , \new_[86036]_ ,
    \new_[86040]_ , \new_[86041]_ , \new_[86044]_ , \new_[86047]_ ,
    \new_[86048]_ , \new_[86049]_ , \new_[86053]_ , \new_[86054]_ ,
    \new_[86057]_ , \new_[86060]_ , \new_[86061]_ , \new_[86062]_ ,
    \new_[86066]_ , \new_[86067]_ , \new_[86070]_ , \new_[86073]_ ,
    \new_[86074]_ , \new_[86075]_ , \new_[86079]_ , \new_[86080]_ ,
    \new_[86083]_ , \new_[86086]_ , \new_[86087]_ , \new_[86088]_ ,
    \new_[86092]_ , \new_[86093]_ , \new_[86096]_ , \new_[86099]_ ,
    \new_[86100]_ , \new_[86101]_ , \new_[86105]_ , \new_[86106]_ ,
    \new_[86109]_ , \new_[86112]_ , \new_[86113]_ , \new_[86114]_ ,
    \new_[86118]_ , \new_[86119]_ , \new_[86122]_ , \new_[86125]_ ,
    \new_[86126]_ , \new_[86127]_ , \new_[86131]_ , \new_[86132]_ ,
    \new_[86135]_ , \new_[86138]_ , \new_[86139]_ , \new_[86140]_ ,
    \new_[86144]_ , \new_[86145]_ , \new_[86148]_ , \new_[86151]_ ,
    \new_[86152]_ , \new_[86153]_ , \new_[86157]_ , \new_[86158]_ ,
    \new_[86161]_ , \new_[86164]_ , \new_[86165]_ , \new_[86166]_ ,
    \new_[86170]_ , \new_[86171]_ , \new_[86174]_ , \new_[86177]_ ,
    \new_[86178]_ , \new_[86179]_ , \new_[86183]_ , \new_[86184]_ ,
    \new_[86187]_ , \new_[86190]_ , \new_[86191]_ , \new_[86192]_ ,
    \new_[86196]_ , \new_[86197]_ , \new_[86200]_ , \new_[86203]_ ,
    \new_[86204]_ , \new_[86205]_ , \new_[86209]_ , \new_[86210]_ ,
    \new_[86213]_ , \new_[86216]_ , \new_[86217]_ , \new_[86218]_ ,
    \new_[86222]_ , \new_[86223]_ , \new_[86226]_ , \new_[86229]_ ,
    \new_[86230]_ , \new_[86231]_ , \new_[86235]_ , \new_[86236]_ ,
    \new_[86239]_ , \new_[86242]_ , \new_[86243]_ , \new_[86244]_ ,
    \new_[86248]_ , \new_[86249]_ , \new_[86252]_ , \new_[86255]_ ,
    \new_[86256]_ , \new_[86257]_ , \new_[86261]_ , \new_[86262]_ ,
    \new_[86265]_ , \new_[86268]_ , \new_[86269]_ , \new_[86270]_ ,
    \new_[86274]_ , \new_[86275]_ , \new_[86278]_ , \new_[86281]_ ,
    \new_[86282]_ , \new_[86283]_ , \new_[86287]_ , \new_[86288]_ ,
    \new_[86291]_ , \new_[86294]_ , \new_[86295]_ , \new_[86296]_ ,
    \new_[86300]_ , \new_[86301]_ , \new_[86304]_ , \new_[86307]_ ,
    \new_[86308]_ , \new_[86309]_ , \new_[86313]_ , \new_[86314]_ ,
    \new_[86317]_ , \new_[86320]_ , \new_[86321]_ , \new_[86322]_ ,
    \new_[86326]_ , \new_[86327]_ , \new_[86330]_ , \new_[86333]_ ,
    \new_[86334]_ , \new_[86335]_ , \new_[86339]_ , \new_[86340]_ ,
    \new_[86343]_ , \new_[86346]_ , \new_[86347]_ , \new_[86348]_ ,
    \new_[86352]_ , \new_[86353]_ , \new_[86356]_ , \new_[86359]_ ,
    \new_[86360]_ , \new_[86361]_ , \new_[86365]_ , \new_[86366]_ ,
    \new_[86369]_ , \new_[86372]_ , \new_[86373]_ , \new_[86374]_ ,
    \new_[86378]_ , \new_[86379]_ , \new_[86382]_ , \new_[86385]_ ,
    \new_[86386]_ , \new_[86387]_ , \new_[86391]_ , \new_[86392]_ ,
    \new_[86395]_ , \new_[86398]_ , \new_[86399]_ , \new_[86400]_ ,
    \new_[86404]_ , \new_[86405]_ , \new_[86408]_ , \new_[86411]_ ,
    \new_[86412]_ , \new_[86413]_ , \new_[86417]_ , \new_[86418]_ ,
    \new_[86421]_ , \new_[86424]_ , \new_[86425]_ , \new_[86426]_ ,
    \new_[86430]_ , \new_[86431]_ , \new_[86434]_ , \new_[86437]_ ,
    \new_[86438]_ , \new_[86439]_ , \new_[86443]_ , \new_[86444]_ ,
    \new_[86447]_ , \new_[86450]_ , \new_[86451]_ , \new_[86452]_ ,
    \new_[86456]_ , \new_[86457]_ , \new_[86460]_ , \new_[86463]_ ,
    \new_[86464]_ , \new_[86465]_ , \new_[86469]_ , \new_[86470]_ ,
    \new_[86473]_ , \new_[86476]_ , \new_[86477]_ , \new_[86478]_ ,
    \new_[86482]_ , \new_[86483]_ , \new_[86486]_ , \new_[86489]_ ,
    \new_[86490]_ , \new_[86491]_ , \new_[86495]_ , \new_[86496]_ ,
    \new_[86499]_ , \new_[86502]_ , \new_[86503]_ , \new_[86504]_ ,
    \new_[86508]_ , \new_[86509]_ , \new_[86512]_ , \new_[86515]_ ,
    \new_[86516]_ , \new_[86517]_ , \new_[86521]_ , \new_[86522]_ ,
    \new_[86525]_ , \new_[86528]_ , \new_[86529]_ , \new_[86530]_ ,
    \new_[86534]_ , \new_[86535]_ , \new_[86538]_ , \new_[86541]_ ,
    \new_[86542]_ , \new_[86543]_ , \new_[86547]_ , \new_[86548]_ ,
    \new_[86551]_ , \new_[86554]_ , \new_[86555]_ , \new_[86556]_ ,
    \new_[86560]_ , \new_[86561]_ , \new_[86564]_ , \new_[86567]_ ,
    \new_[86568]_ , \new_[86569]_ , \new_[86573]_ , \new_[86574]_ ,
    \new_[86577]_ , \new_[86580]_ , \new_[86581]_ , \new_[86582]_ ,
    \new_[86586]_ , \new_[86587]_ , \new_[86590]_ , \new_[86593]_ ,
    \new_[86594]_ , \new_[86595]_ , \new_[86599]_ , \new_[86600]_ ,
    \new_[86603]_ , \new_[86606]_ , \new_[86607]_ , \new_[86608]_ ,
    \new_[86612]_ , \new_[86613]_ , \new_[86616]_ , \new_[86619]_ ,
    \new_[86620]_ , \new_[86621]_ , \new_[86625]_ , \new_[86626]_ ,
    \new_[86629]_ , \new_[86632]_ , \new_[86633]_ , \new_[86634]_ ,
    \new_[86638]_ , \new_[86639]_ , \new_[86642]_ , \new_[86645]_ ,
    \new_[86646]_ , \new_[86647]_ , \new_[86651]_ , \new_[86652]_ ,
    \new_[86655]_ , \new_[86658]_ , \new_[86659]_ , \new_[86660]_ ,
    \new_[86664]_ , \new_[86665]_ , \new_[86668]_ , \new_[86671]_ ,
    \new_[86672]_ , \new_[86673]_ , \new_[86677]_ , \new_[86678]_ ,
    \new_[86681]_ , \new_[86684]_ , \new_[86685]_ , \new_[86686]_ ,
    \new_[86690]_ , \new_[86691]_ , \new_[86694]_ , \new_[86697]_ ,
    \new_[86698]_ , \new_[86699]_ , \new_[86703]_ , \new_[86704]_ ,
    \new_[86707]_ , \new_[86710]_ , \new_[86711]_ , \new_[86712]_ ,
    \new_[86716]_ , \new_[86717]_ , \new_[86720]_ , \new_[86723]_ ,
    \new_[86724]_ , \new_[86725]_ , \new_[86729]_ , \new_[86730]_ ,
    \new_[86733]_ , \new_[86736]_ , \new_[86737]_ , \new_[86738]_ ,
    \new_[86742]_ , \new_[86743]_ , \new_[86746]_ , \new_[86749]_ ,
    \new_[86750]_ , \new_[86751]_ , \new_[86755]_ , \new_[86756]_ ,
    \new_[86759]_ , \new_[86762]_ , \new_[86763]_ , \new_[86764]_ ,
    \new_[86768]_ , \new_[86769]_ , \new_[86772]_ , \new_[86775]_ ,
    \new_[86776]_ , \new_[86777]_ , \new_[86781]_ , \new_[86782]_ ,
    \new_[86785]_ , \new_[86788]_ , \new_[86789]_ , \new_[86790]_ ,
    \new_[86794]_ , \new_[86795]_ , \new_[86798]_ , \new_[86801]_ ,
    \new_[86802]_ , \new_[86803]_ , \new_[86806]_ , \new_[86809]_ ,
    \new_[86810]_ , \new_[86813]_ , \new_[86816]_ , \new_[86817]_ ,
    \new_[86818]_ , \new_[86822]_ , \new_[86823]_ , \new_[86826]_ ,
    \new_[86829]_ , \new_[86830]_ , \new_[86831]_ , \new_[86834]_ ,
    \new_[86837]_ , \new_[86838]_ , \new_[86841]_ , \new_[86844]_ ,
    \new_[86845]_ , \new_[86846]_ , \new_[86850]_ , \new_[86851]_ ,
    \new_[86854]_ , \new_[86857]_ , \new_[86858]_ , \new_[86859]_ ,
    \new_[86862]_ , \new_[86865]_ , \new_[86866]_ , \new_[86869]_ ,
    \new_[86872]_ , \new_[86873]_ , \new_[86874]_ , \new_[86878]_ ,
    \new_[86879]_ , \new_[86882]_ , \new_[86885]_ , \new_[86886]_ ,
    \new_[86887]_ , \new_[86890]_ , \new_[86893]_ , \new_[86894]_ ,
    \new_[86897]_ , \new_[86900]_ , \new_[86901]_ , \new_[86902]_ ,
    \new_[86906]_ , \new_[86907]_ , \new_[86910]_ , \new_[86913]_ ,
    \new_[86914]_ , \new_[86915]_ , \new_[86918]_ , \new_[86921]_ ,
    \new_[86922]_ , \new_[86925]_ , \new_[86928]_ , \new_[86929]_ ,
    \new_[86930]_ , \new_[86934]_ , \new_[86935]_ , \new_[86938]_ ,
    \new_[86941]_ , \new_[86942]_ , \new_[86943]_ , \new_[86946]_ ,
    \new_[86949]_ , \new_[86950]_ , \new_[86953]_ , \new_[86956]_ ,
    \new_[86957]_ , \new_[86958]_ , \new_[86962]_ , \new_[86963]_ ,
    \new_[86966]_ , \new_[86969]_ , \new_[86970]_ , \new_[86971]_ ,
    \new_[86974]_ , \new_[86977]_ , \new_[86978]_ , \new_[86981]_ ,
    \new_[86984]_ , \new_[86985]_ , \new_[86986]_ , \new_[86990]_ ,
    \new_[86991]_ , \new_[86994]_ , \new_[86997]_ , \new_[86998]_ ,
    \new_[86999]_ , \new_[87002]_ , \new_[87005]_ , \new_[87006]_ ,
    \new_[87009]_ , \new_[87012]_ , \new_[87013]_ , \new_[87014]_ ,
    \new_[87018]_ , \new_[87019]_ , \new_[87022]_ , \new_[87025]_ ,
    \new_[87026]_ , \new_[87027]_ , \new_[87030]_ , \new_[87033]_ ,
    \new_[87034]_ , \new_[87037]_ , \new_[87040]_ , \new_[87041]_ ,
    \new_[87042]_ , \new_[87046]_ , \new_[87047]_ , \new_[87050]_ ,
    \new_[87053]_ , \new_[87054]_ , \new_[87055]_ , \new_[87058]_ ,
    \new_[87061]_ , \new_[87062]_ , \new_[87065]_ , \new_[87068]_ ,
    \new_[87069]_ , \new_[87070]_ , \new_[87074]_ , \new_[87075]_ ,
    \new_[87078]_ , \new_[87081]_ , \new_[87082]_ , \new_[87083]_ ,
    \new_[87086]_ , \new_[87089]_ , \new_[87090]_ , \new_[87093]_ ,
    \new_[87096]_ , \new_[87097]_ , \new_[87098]_ , \new_[87102]_ ,
    \new_[87103]_ , \new_[87106]_ , \new_[87109]_ , \new_[87110]_ ,
    \new_[87111]_ , \new_[87114]_ , \new_[87117]_ , \new_[87118]_ ,
    \new_[87121]_ , \new_[87124]_ , \new_[87125]_ , \new_[87126]_ ,
    \new_[87130]_ , \new_[87131]_ , \new_[87134]_ , \new_[87137]_ ,
    \new_[87138]_ , \new_[87139]_ , \new_[87142]_ , \new_[87145]_ ,
    \new_[87146]_ , \new_[87149]_ , \new_[87152]_ , \new_[87153]_ ,
    \new_[87154]_ , \new_[87158]_ , \new_[87159]_ , \new_[87162]_ ,
    \new_[87165]_ , \new_[87166]_ , \new_[87167]_ , \new_[87170]_ ,
    \new_[87173]_ , \new_[87174]_ , \new_[87177]_ , \new_[87180]_ ,
    \new_[87181]_ , \new_[87182]_ , \new_[87186]_ , \new_[87187]_ ,
    \new_[87190]_ , \new_[87193]_ , \new_[87194]_ , \new_[87195]_ ,
    \new_[87198]_ , \new_[87201]_ , \new_[87202]_ , \new_[87205]_ ,
    \new_[87208]_ , \new_[87209]_ , \new_[87210]_ , \new_[87214]_ ,
    \new_[87215]_ , \new_[87218]_ , \new_[87221]_ , \new_[87222]_ ,
    \new_[87223]_ , \new_[87226]_ , \new_[87229]_ , \new_[87230]_ ,
    \new_[87233]_ , \new_[87236]_ , \new_[87237]_ , \new_[87238]_ ,
    \new_[87242]_ , \new_[87243]_ , \new_[87246]_ , \new_[87249]_ ,
    \new_[87250]_ , \new_[87251]_ , \new_[87254]_ , \new_[87257]_ ,
    \new_[87258]_ , \new_[87261]_ , \new_[87264]_ , \new_[87265]_ ,
    \new_[87266]_ , \new_[87270]_ , \new_[87271]_ , \new_[87274]_ ,
    \new_[87277]_ , \new_[87278]_ , \new_[87279]_ , \new_[87282]_ ,
    \new_[87285]_ , \new_[87286]_ , \new_[87289]_ , \new_[87292]_ ,
    \new_[87293]_ , \new_[87294]_ , \new_[87298]_ , \new_[87299]_ ,
    \new_[87302]_ , \new_[87305]_ , \new_[87306]_ , \new_[87307]_ ,
    \new_[87310]_ , \new_[87313]_ , \new_[87314]_ , \new_[87317]_ ,
    \new_[87320]_ , \new_[87321]_ , \new_[87322]_ , \new_[87326]_ ,
    \new_[87327]_ , \new_[87330]_ , \new_[87333]_ , \new_[87334]_ ,
    \new_[87335]_ , \new_[87338]_ , \new_[87341]_ , \new_[87342]_ ,
    \new_[87345]_ , \new_[87348]_ , \new_[87349]_ , \new_[87350]_ ,
    \new_[87354]_ , \new_[87355]_ , \new_[87358]_ , \new_[87361]_ ,
    \new_[87362]_ , \new_[87363]_ , \new_[87366]_ , \new_[87369]_ ,
    \new_[87370]_ , \new_[87373]_ , \new_[87376]_ , \new_[87377]_ ,
    \new_[87378]_ , \new_[87382]_ , \new_[87383]_ , \new_[87386]_ ,
    \new_[87389]_ , \new_[87390]_ , \new_[87391]_ , \new_[87394]_ ,
    \new_[87397]_ , \new_[87398]_ , \new_[87401]_ , \new_[87404]_ ,
    \new_[87405]_ , \new_[87406]_ , \new_[87410]_ , \new_[87411]_ ,
    \new_[87414]_ , \new_[87417]_ , \new_[87418]_ , \new_[87419]_ ,
    \new_[87422]_ , \new_[87425]_ , \new_[87426]_ , \new_[87429]_ ,
    \new_[87432]_ , \new_[87433]_ , \new_[87434]_ , \new_[87438]_ ,
    \new_[87439]_ , \new_[87442]_ , \new_[87445]_ , \new_[87446]_ ,
    \new_[87447]_ , \new_[87450]_ , \new_[87453]_ , \new_[87454]_ ,
    \new_[87457]_ , \new_[87460]_ , \new_[87461]_ , \new_[87462]_ ,
    \new_[87466]_ , \new_[87467]_ , \new_[87470]_ , \new_[87473]_ ,
    \new_[87474]_ , \new_[87475]_ , \new_[87478]_ , \new_[87481]_ ,
    \new_[87482]_ , \new_[87485]_ , \new_[87488]_ , \new_[87489]_ ,
    \new_[87490]_ , \new_[87494]_ , \new_[87495]_ , \new_[87498]_ ,
    \new_[87501]_ , \new_[87502]_ , \new_[87503]_ , \new_[87506]_ ,
    \new_[87509]_ , \new_[87510]_ , \new_[87513]_ , \new_[87516]_ ,
    \new_[87517]_ , \new_[87518]_ , \new_[87522]_ , \new_[87523]_ ,
    \new_[87526]_ , \new_[87529]_ , \new_[87530]_ , \new_[87531]_ ,
    \new_[87534]_ , \new_[87537]_ , \new_[87538]_ , \new_[87541]_ ,
    \new_[87544]_ , \new_[87545]_ , \new_[87546]_ , \new_[87550]_ ,
    \new_[87551]_ , \new_[87554]_ , \new_[87557]_ , \new_[87558]_ ,
    \new_[87559]_ , \new_[87562]_ , \new_[87565]_ , \new_[87566]_ ,
    \new_[87569]_ , \new_[87572]_ , \new_[87573]_ , \new_[87574]_ ,
    \new_[87578]_ , \new_[87579]_ , \new_[87582]_ , \new_[87585]_ ,
    \new_[87586]_ , \new_[87587]_ , \new_[87590]_ , \new_[87593]_ ,
    \new_[87594]_ , \new_[87597]_ , \new_[87600]_ , \new_[87601]_ ,
    \new_[87602]_ , \new_[87606]_ , \new_[87607]_ , \new_[87610]_ ,
    \new_[87613]_ , \new_[87614]_ , \new_[87615]_ , \new_[87618]_ ,
    \new_[87621]_ , \new_[87622]_ , \new_[87625]_ , \new_[87628]_ ,
    \new_[87629]_ , \new_[87630]_ , \new_[87634]_ , \new_[87635]_ ,
    \new_[87638]_ , \new_[87641]_ , \new_[87642]_ , \new_[87643]_ ,
    \new_[87646]_ , \new_[87649]_ , \new_[87650]_ , \new_[87653]_ ,
    \new_[87656]_ , \new_[87657]_ , \new_[87658]_ , \new_[87662]_ ,
    \new_[87663]_ , \new_[87666]_ , \new_[87669]_ , \new_[87670]_ ,
    \new_[87671]_ , \new_[87674]_ , \new_[87677]_ , \new_[87678]_ ,
    \new_[87681]_ , \new_[87684]_ , \new_[87685]_ , \new_[87686]_ ,
    \new_[87690]_ , \new_[87691]_ , \new_[87694]_ , \new_[87697]_ ,
    \new_[87698]_ , \new_[87699]_ , \new_[87702]_ , \new_[87705]_ ,
    \new_[87706]_ , \new_[87709]_ , \new_[87712]_ , \new_[87713]_ ,
    \new_[87714]_ , \new_[87718]_ , \new_[87719]_ , \new_[87722]_ ,
    \new_[87725]_ , \new_[87726]_ , \new_[87727]_ , \new_[87730]_ ,
    \new_[87733]_ , \new_[87734]_ , \new_[87737]_ , \new_[87740]_ ,
    \new_[87741]_ , \new_[87742]_ , \new_[87746]_ , \new_[87747]_ ,
    \new_[87750]_ , \new_[87753]_ , \new_[87754]_ , \new_[87755]_ ,
    \new_[87758]_ , \new_[87761]_ , \new_[87762]_ , \new_[87765]_ ,
    \new_[87768]_ , \new_[87769]_ , \new_[87770]_ , \new_[87774]_ ,
    \new_[87775]_ , \new_[87778]_ , \new_[87781]_ , \new_[87782]_ ,
    \new_[87783]_ , \new_[87786]_ , \new_[87789]_ , \new_[87790]_ ,
    \new_[87793]_ , \new_[87796]_ , \new_[87797]_ , \new_[87798]_ ,
    \new_[87802]_ , \new_[87803]_ , \new_[87806]_ , \new_[87809]_ ,
    \new_[87810]_ , \new_[87811]_ , \new_[87814]_ , \new_[87817]_ ,
    \new_[87818]_ , \new_[87821]_ , \new_[87824]_ , \new_[87825]_ ,
    \new_[87826]_ , \new_[87830]_ , \new_[87831]_ , \new_[87834]_ ,
    \new_[87837]_ , \new_[87838]_ , \new_[87839]_ , \new_[87842]_ ,
    \new_[87845]_ , \new_[87846]_ , \new_[87849]_ , \new_[87852]_ ,
    \new_[87853]_ , \new_[87854]_ , \new_[87858]_ , \new_[87859]_ ,
    \new_[87862]_ , \new_[87865]_ , \new_[87866]_ , \new_[87867]_ ,
    \new_[87870]_ , \new_[87873]_ , \new_[87874]_ , \new_[87877]_ ,
    \new_[87880]_ , \new_[87881]_ , \new_[87882]_ , \new_[87886]_ ,
    \new_[87887]_ , \new_[87890]_ , \new_[87893]_ , \new_[87894]_ ,
    \new_[87895]_ , \new_[87898]_ , \new_[87901]_ , \new_[87902]_ ,
    \new_[87905]_ , \new_[87908]_ , \new_[87909]_ , \new_[87910]_ ,
    \new_[87914]_ , \new_[87915]_ , \new_[87918]_ , \new_[87921]_ ,
    \new_[87922]_ , \new_[87923]_ , \new_[87926]_ , \new_[87929]_ ,
    \new_[87930]_ , \new_[87933]_ , \new_[87936]_ , \new_[87937]_ ,
    \new_[87938]_ , \new_[87942]_ , \new_[87943]_ , \new_[87946]_ ,
    \new_[87949]_ , \new_[87950]_ , \new_[87951]_ , \new_[87954]_ ,
    \new_[87957]_ , \new_[87958]_ , \new_[87961]_ , \new_[87964]_ ,
    \new_[87965]_ , \new_[87966]_ , \new_[87970]_ , \new_[87971]_ ,
    \new_[87974]_ , \new_[87977]_ , \new_[87978]_ , \new_[87979]_ ,
    \new_[87982]_ , \new_[87985]_ , \new_[87986]_ , \new_[87989]_ ,
    \new_[87992]_ , \new_[87993]_ , \new_[87994]_ , \new_[87998]_ ,
    \new_[87999]_ , \new_[88002]_ , \new_[88005]_ , \new_[88006]_ ,
    \new_[88007]_ , \new_[88010]_ , \new_[88013]_ , \new_[88014]_ ,
    \new_[88017]_ , \new_[88020]_ , \new_[88021]_ , \new_[88022]_ ,
    \new_[88026]_ , \new_[88027]_ , \new_[88030]_ , \new_[88033]_ ,
    \new_[88034]_ , \new_[88035]_ , \new_[88038]_ , \new_[88041]_ ,
    \new_[88042]_ , \new_[88045]_ , \new_[88048]_ , \new_[88049]_ ,
    \new_[88050]_ , \new_[88054]_ , \new_[88055]_ , \new_[88058]_ ,
    \new_[88061]_ , \new_[88062]_ , \new_[88063]_ , \new_[88066]_ ,
    \new_[88069]_ , \new_[88070]_ , \new_[88073]_ , \new_[88076]_ ,
    \new_[88077]_ , \new_[88078]_ , \new_[88082]_ , \new_[88083]_ ,
    \new_[88086]_ , \new_[88089]_ , \new_[88090]_ , \new_[88091]_ ,
    \new_[88094]_ , \new_[88097]_ , \new_[88098]_ , \new_[88101]_ ,
    \new_[88104]_ , \new_[88105]_ , \new_[88106]_ , \new_[88110]_ ,
    \new_[88111]_ , \new_[88114]_ , \new_[88117]_ , \new_[88118]_ ,
    \new_[88119]_ , \new_[88122]_ , \new_[88125]_ , \new_[88126]_ ,
    \new_[88129]_ , \new_[88132]_ , \new_[88133]_ , \new_[88134]_ ,
    \new_[88138]_ , \new_[88139]_ , \new_[88142]_ , \new_[88145]_ ,
    \new_[88146]_ , \new_[88147]_ , \new_[88150]_ , \new_[88153]_ ,
    \new_[88154]_ , \new_[88157]_ , \new_[88160]_ , \new_[88161]_ ,
    \new_[88162]_ , \new_[88166]_ , \new_[88167]_ , \new_[88170]_ ,
    \new_[88173]_ , \new_[88174]_ , \new_[88175]_ , \new_[88178]_ ,
    \new_[88181]_ , \new_[88182]_ , \new_[88185]_ , \new_[88188]_ ,
    \new_[88189]_ , \new_[88190]_ , \new_[88194]_ , \new_[88195]_ ,
    \new_[88198]_ , \new_[88201]_ , \new_[88202]_ , \new_[88203]_ ,
    \new_[88206]_ , \new_[88209]_ , \new_[88210]_ , \new_[88213]_ ,
    \new_[88216]_ , \new_[88217]_ , \new_[88218]_ , \new_[88222]_ ,
    \new_[88223]_ , \new_[88226]_ , \new_[88229]_ , \new_[88230]_ ,
    \new_[88231]_ , \new_[88234]_ , \new_[88237]_ , \new_[88238]_ ,
    \new_[88241]_ , \new_[88244]_ , \new_[88245]_ , \new_[88246]_ ,
    \new_[88250]_ , \new_[88251]_ , \new_[88254]_ , \new_[88257]_ ,
    \new_[88258]_ , \new_[88259]_ , \new_[88262]_ , \new_[88265]_ ,
    \new_[88266]_ , \new_[88269]_ , \new_[88272]_ , \new_[88273]_ ,
    \new_[88274]_ , \new_[88278]_ , \new_[88279]_ , \new_[88282]_ ,
    \new_[88285]_ , \new_[88286]_ , \new_[88287]_ , \new_[88290]_ ,
    \new_[88293]_ , \new_[88294]_ , \new_[88297]_ , \new_[88300]_ ,
    \new_[88301]_ , \new_[88302]_ , \new_[88306]_ , \new_[88307]_ ,
    \new_[88310]_ , \new_[88313]_ , \new_[88314]_ , \new_[88315]_ ,
    \new_[88318]_ , \new_[88321]_ , \new_[88322]_ , \new_[88325]_ ,
    \new_[88328]_ , \new_[88329]_ , \new_[88330]_ , \new_[88334]_ ,
    \new_[88335]_ , \new_[88338]_ , \new_[88341]_ , \new_[88342]_ ,
    \new_[88343]_ , \new_[88346]_ , \new_[88349]_ , \new_[88350]_ ,
    \new_[88353]_ , \new_[88356]_ , \new_[88357]_ , \new_[88358]_ ,
    \new_[88362]_ , \new_[88363]_ , \new_[88366]_ , \new_[88369]_ ,
    \new_[88370]_ , \new_[88371]_ , \new_[88374]_ , \new_[88377]_ ,
    \new_[88378]_ , \new_[88381]_ , \new_[88384]_ , \new_[88385]_ ,
    \new_[88386]_ , \new_[88390]_ , \new_[88391]_ , \new_[88394]_ ,
    \new_[88397]_ , \new_[88398]_ , \new_[88399]_ , \new_[88402]_ ,
    \new_[88405]_ , \new_[88406]_ , \new_[88409]_ , \new_[88412]_ ,
    \new_[88413]_ , \new_[88414]_ , \new_[88418]_ , \new_[88419]_ ,
    \new_[88422]_ , \new_[88425]_ , \new_[88426]_ , \new_[88427]_ ,
    \new_[88430]_ , \new_[88433]_ , \new_[88434]_ , \new_[88437]_ ,
    \new_[88440]_ , \new_[88441]_ , \new_[88442]_ , \new_[88446]_ ,
    \new_[88447]_ , \new_[88450]_ , \new_[88453]_ , \new_[88454]_ ,
    \new_[88455]_ , \new_[88458]_ , \new_[88461]_ , \new_[88462]_ ,
    \new_[88465]_ , \new_[88468]_ , \new_[88469]_ , \new_[88470]_ ,
    \new_[88474]_ , \new_[88475]_ , \new_[88478]_ , \new_[88481]_ ,
    \new_[88482]_ , \new_[88483]_ , \new_[88486]_ , \new_[88489]_ ,
    \new_[88490]_ , \new_[88493]_ , \new_[88496]_ , \new_[88497]_ ,
    \new_[88498]_ , \new_[88502]_ , \new_[88503]_ , \new_[88506]_ ,
    \new_[88509]_ , \new_[88510]_ , \new_[88511]_ , \new_[88514]_ ,
    \new_[88517]_ , \new_[88518]_ , \new_[88521]_ , \new_[88524]_ ,
    \new_[88525]_ , \new_[88526]_ , \new_[88530]_ , \new_[88531]_ ,
    \new_[88534]_ , \new_[88537]_ , \new_[88538]_ , \new_[88539]_ ,
    \new_[88542]_ , \new_[88545]_ , \new_[88546]_ , \new_[88549]_ ,
    \new_[88552]_ , \new_[88553]_ , \new_[88554]_ , \new_[88558]_ ,
    \new_[88559]_ , \new_[88562]_ , \new_[88565]_ , \new_[88566]_ ,
    \new_[88567]_ , \new_[88570]_ , \new_[88573]_ , \new_[88574]_ ,
    \new_[88577]_ , \new_[88580]_ , \new_[88581]_ , \new_[88582]_ ,
    \new_[88586]_ , \new_[88587]_ , \new_[88590]_ , \new_[88593]_ ,
    \new_[88594]_ , \new_[88595]_ , \new_[88598]_ , \new_[88601]_ ,
    \new_[88602]_ , \new_[88605]_ , \new_[88608]_ , \new_[88609]_ ,
    \new_[88610]_ , \new_[88614]_ , \new_[88615]_ , \new_[88618]_ ,
    \new_[88621]_ , \new_[88622]_ , \new_[88623]_ , \new_[88626]_ ,
    \new_[88629]_ , \new_[88630]_ , \new_[88633]_ , \new_[88636]_ ,
    \new_[88637]_ , \new_[88638]_ , \new_[88642]_ , \new_[88643]_ ,
    \new_[88646]_ , \new_[88649]_ , \new_[88650]_ , \new_[88651]_ ,
    \new_[88654]_ , \new_[88657]_ , \new_[88658]_ , \new_[88661]_ ,
    \new_[88664]_ , \new_[88665]_ , \new_[88666]_ , \new_[88670]_ ,
    \new_[88671]_ , \new_[88674]_ , \new_[88677]_ , \new_[88678]_ ,
    \new_[88679]_ , \new_[88682]_ , \new_[88685]_ , \new_[88686]_ ,
    \new_[88689]_ , \new_[88692]_ , \new_[88693]_ , \new_[88694]_ ,
    \new_[88698]_ , \new_[88699]_ , \new_[88702]_ , \new_[88705]_ ,
    \new_[88706]_ , \new_[88707]_ , \new_[88710]_ , \new_[88713]_ ,
    \new_[88714]_ , \new_[88717]_ , \new_[88720]_ , \new_[88721]_ ,
    \new_[88722]_ , \new_[88726]_ , \new_[88727]_ , \new_[88730]_ ,
    \new_[88733]_ , \new_[88734]_ , \new_[88735]_ , \new_[88738]_ ,
    \new_[88741]_ , \new_[88742]_ , \new_[88745]_ , \new_[88748]_ ,
    \new_[88749]_ , \new_[88750]_ , \new_[88754]_ , \new_[88755]_ ,
    \new_[88758]_ , \new_[88761]_ , \new_[88762]_ , \new_[88763]_ ,
    \new_[88766]_ , \new_[88769]_ , \new_[88770]_ , \new_[88773]_ ,
    \new_[88776]_ , \new_[88777]_ , \new_[88778]_ , \new_[88782]_ ,
    \new_[88783]_ , \new_[88786]_ , \new_[88789]_ , \new_[88790]_ ,
    \new_[88791]_ , \new_[88794]_ , \new_[88797]_ , \new_[88798]_ ,
    \new_[88801]_ , \new_[88804]_ , \new_[88805]_ , \new_[88806]_ ,
    \new_[88810]_ , \new_[88811]_ , \new_[88814]_ , \new_[88817]_ ,
    \new_[88818]_ , \new_[88819]_ , \new_[88822]_ , \new_[88825]_ ,
    \new_[88826]_ , \new_[88829]_ , \new_[88832]_ , \new_[88833]_ ,
    \new_[88834]_ , \new_[88838]_ , \new_[88839]_ , \new_[88842]_ ,
    \new_[88845]_ , \new_[88846]_ , \new_[88847]_ , \new_[88850]_ ,
    \new_[88853]_ , \new_[88854]_ , \new_[88857]_ , \new_[88860]_ ,
    \new_[88861]_ , \new_[88862]_ , \new_[88866]_ , \new_[88867]_ ,
    \new_[88870]_ , \new_[88873]_ , \new_[88874]_ , \new_[88875]_ ,
    \new_[88878]_ , \new_[88881]_ , \new_[88882]_ , \new_[88885]_ ,
    \new_[88888]_ , \new_[88889]_ , \new_[88890]_ , \new_[88894]_ ,
    \new_[88895]_ , \new_[88898]_ , \new_[88901]_ , \new_[88902]_ ,
    \new_[88903]_ , \new_[88906]_ , \new_[88909]_ , \new_[88910]_ ,
    \new_[88913]_ , \new_[88916]_ , \new_[88917]_ , \new_[88918]_ ,
    \new_[88922]_ , \new_[88923]_ , \new_[88926]_ , \new_[88929]_ ,
    \new_[88930]_ , \new_[88931]_ , \new_[88934]_ , \new_[88937]_ ,
    \new_[88938]_ , \new_[88941]_ , \new_[88944]_ , \new_[88945]_ ,
    \new_[88946]_ , \new_[88950]_ , \new_[88951]_ , \new_[88954]_ ,
    \new_[88957]_ , \new_[88958]_ , \new_[88959]_ , \new_[88962]_ ,
    \new_[88965]_ , \new_[88966]_ , \new_[88969]_ , \new_[88972]_ ,
    \new_[88973]_ , \new_[88974]_ , \new_[88978]_ , \new_[88979]_ ,
    \new_[88982]_ , \new_[88985]_ , \new_[88986]_ , \new_[88987]_ ,
    \new_[88990]_ , \new_[88993]_ , \new_[88994]_ , \new_[88997]_ ,
    \new_[89000]_ , \new_[89001]_ , \new_[89002]_ , \new_[89006]_ ,
    \new_[89007]_ , \new_[89010]_ , \new_[89013]_ , \new_[89014]_ ,
    \new_[89015]_ , \new_[89018]_ , \new_[89021]_ , \new_[89022]_ ,
    \new_[89025]_ , \new_[89028]_ , \new_[89029]_ , \new_[89030]_ ,
    \new_[89034]_ , \new_[89035]_ , \new_[89038]_ , \new_[89041]_ ,
    \new_[89042]_ , \new_[89043]_ , \new_[89046]_ , \new_[89049]_ ,
    \new_[89050]_ , \new_[89053]_ , \new_[89056]_ , \new_[89057]_ ,
    \new_[89058]_ , \new_[89062]_ , \new_[89063]_ , \new_[89066]_ ,
    \new_[89069]_ , \new_[89070]_ , \new_[89071]_ , \new_[89074]_ ,
    \new_[89077]_ , \new_[89078]_ , \new_[89081]_ , \new_[89084]_ ,
    \new_[89085]_ , \new_[89086]_ , \new_[89090]_ , \new_[89091]_ ,
    \new_[89094]_ , \new_[89097]_ , \new_[89098]_ , \new_[89099]_ ,
    \new_[89102]_ , \new_[89105]_ , \new_[89106]_ , \new_[89109]_ ,
    \new_[89112]_ , \new_[89113]_ , \new_[89114]_ , \new_[89118]_ ,
    \new_[89119]_ , \new_[89122]_ , \new_[89125]_ , \new_[89126]_ ,
    \new_[89127]_ , \new_[89130]_ , \new_[89133]_ , \new_[89134]_ ,
    \new_[89137]_ , \new_[89140]_ , \new_[89141]_ , \new_[89142]_ ,
    \new_[89146]_ , \new_[89147]_ , \new_[89150]_ , \new_[89153]_ ,
    \new_[89154]_ , \new_[89155]_ , \new_[89158]_ , \new_[89161]_ ,
    \new_[89162]_ , \new_[89165]_ , \new_[89168]_ , \new_[89169]_ ,
    \new_[89170]_ , \new_[89174]_ , \new_[89175]_ , \new_[89178]_ ,
    \new_[89181]_ , \new_[89182]_ , \new_[89183]_ , \new_[89186]_ ,
    \new_[89189]_ , \new_[89190]_ , \new_[89193]_ , \new_[89196]_ ,
    \new_[89197]_ , \new_[89198]_ , \new_[89202]_ , \new_[89203]_ ,
    \new_[89206]_ , \new_[89209]_ , \new_[89210]_ , \new_[89211]_ ,
    \new_[89214]_ , \new_[89217]_ , \new_[89218]_ , \new_[89221]_ ,
    \new_[89224]_ , \new_[89225]_ , \new_[89226]_ , \new_[89230]_ ,
    \new_[89231]_ , \new_[89234]_ , \new_[89237]_ , \new_[89238]_ ,
    \new_[89239]_ , \new_[89242]_ , \new_[89245]_ , \new_[89246]_ ,
    \new_[89249]_ , \new_[89252]_ , \new_[89253]_ , \new_[89254]_ ,
    \new_[89258]_ , \new_[89259]_ , \new_[89262]_ , \new_[89265]_ ,
    \new_[89266]_ , \new_[89267]_ , \new_[89270]_ , \new_[89273]_ ,
    \new_[89274]_ , \new_[89277]_ , \new_[89280]_ , \new_[89281]_ ,
    \new_[89282]_ , \new_[89286]_ , \new_[89287]_ , \new_[89290]_ ,
    \new_[89293]_ , \new_[89294]_ , \new_[89295]_ , \new_[89298]_ ,
    \new_[89301]_ , \new_[89302]_ , \new_[89305]_ , \new_[89308]_ ,
    \new_[89309]_ , \new_[89310]_ , \new_[89314]_ , \new_[89315]_ ,
    \new_[89318]_ , \new_[89321]_ , \new_[89322]_ , \new_[89323]_ ,
    \new_[89326]_ , \new_[89329]_ , \new_[89330]_ , \new_[89333]_ ,
    \new_[89336]_ , \new_[89337]_ , \new_[89338]_ , \new_[89342]_ ,
    \new_[89343]_ , \new_[89346]_ , \new_[89349]_ , \new_[89350]_ ,
    \new_[89351]_ , \new_[89354]_ , \new_[89357]_ , \new_[89358]_ ,
    \new_[89361]_ , \new_[89364]_ , \new_[89365]_ , \new_[89366]_ ,
    \new_[89370]_ , \new_[89371]_ , \new_[89374]_ , \new_[89377]_ ,
    \new_[89378]_ , \new_[89379]_ , \new_[89382]_ , \new_[89385]_ ,
    \new_[89386]_ , \new_[89389]_ , \new_[89392]_ , \new_[89393]_ ,
    \new_[89394]_ , \new_[89398]_ , \new_[89399]_ , \new_[89402]_ ,
    \new_[89405]_ , \new_[89406]_ , \new_[89407]_ , \new_[89410]_ ,
    \new_[89413]_ , \new_[89414]_ , \new_[89417]_ , \new_[89420]_ ,
    \new_[89421]_ , \new_[89422]_ , \new_[89426]_ , \new_[89427]_ ,
    \new_[89430]_ , \new_[89433]_ , \new_[89434]_ , \new_[89435]_ ,
    \new_[89438]_ , \new_[89441]_ , \new_[89442]_ , \new_[89445]_ ,
    \new_[89448]_ , \new_[89449]_ , \new_[89450]_ , \new_[89454]_ ,
    \new_[89455]_ , \new_[89458]_ , \new_[89461]_ , \new_[89462]_ ,
    \new_[89463]_ , \new_[89466]_ , \new_[89469]_ , \new_[89470]_ ,
    \new_[89473]_ , \new_[89476]_ , \new_[89477]_ , \new_[89478]_ ,
    \new_[89482]_ , \new_[89483]_ , \new_[89486]_ , \new_[89489]_ ,
    \new_[89490]_ , \new_[89491]_ , \new_[89494]_ , \new_[89497]_ ,
    \new_[89498]_ , \new_[89501]_ , \new_[89504]_ , \new_[89505]_ ,
    \new_[89506]_ , \new_[89510]_ , \new_[89511]_ , \new_[89514]_ ,
    \new_[89517]_ , \new_[89518]_ , \new_[89519]_ , \new_[89522]_ ,
    \new_[89525]_ , \new_[89526]_ , \new_[89529]_ , \new_[89532]_ ,
    \new_[89533]_ , \new_[89534]_ , \new_[89538]_ , \new_[89539]_ ,
    \new_[89542]_ , \new_[89545]_ , \new_[89546]_ , \new_[89547]_ ,
    \new_[89550]_ , \new_[89553]_ , \new_[89554]_ , \new_[89557]_ ,
    \new_[89560]_ , \new_[89561]_ , \new_[89562]_ , \new_[89566]_ ,
    \new_[89567]_ , \new_[89570]_ , \new_[89573]_ , \new_[89574]_ ,
    \new_[89575]_ , \new_[89578]_ , \new_[89581]_ , \new_[89582]_ ,
    \new_[89585]_ , \new_[89588]_ , \new_[89589]_ , \new_[89590]_ ,
    \new_[89594]_ , \new_[89595]_ , \new_[89598]_ , \new_[89601]_ ,
    \new_[89602]_ , \new_[89603]_ , \new_[89606]_ , \new_[89609]_ ,
    \new_[89610]_ , \new_[89613]_ , \new_[89616]_ , \new_[89617]_ ,
    \new_[89618]_ , \new_[89622]_ , \new_[89623]_ , \new_[89626]_ ,
    \new_[89629]_ , \new_[89630]_ , \new_[89631]_ , \new_[89634]_ ,
    \new_[89637]_ , \new_[89638]_ , \new_[89641]_ , \new_[89644]_ ,
    \new_[89645]_ , \new_[89646]_ , \new_[89650]_ , \new_[89651]_ ,
    \new_[89654]_ , \new_[89657]_ , \new_[89658]_ , \new_[89659]_ ,
    \new_[89662]_ , \new_[89665]_ , \new_[89666]_ , \new_[89669]_ ,
    \new_[89672]_ , \new_[89673]_ , \new_[89674]_ , \new_[89678]_ ,
    \new_[89679]_ , \new_[89682]_ , \new_[89685]_ , \new_[89686]_ ,
    \new_[89687]_ , \new_[89690]_ , \new_[89693]_ , \new_[89694]_ ,
    \new_[89697]_ , \new_[89700]_ , \new_[89701]_ , \new_[89702]_ ,
    \new_[89706]_ , \new_[89707]_ , \new_[89710]_ , \new_[89713]_ ,
    \new_[89714]_ , \new_[89715]_ , \new_[89718]_ , \new_[89721]_ ,
    \new_[89722]_ , \new_[89725]_ , \new_[89728]_ , \new_[89729]_ ,
    \new_[89730]_ , \new_[89734]_ , \new_[89735]_ , \new_[89738]_ ,
    \new_[89741]_ , \new_[89742]_ , \new_[89743]_ , \new_[89746]_ ,
    \new_[89749]_ , \new_[89750]_ , \new_[89753]_ , \new_[89756]_ ,
    \new_[89757]_ , \new_[89758]_ , \new_[89762]_ , \new_[89763]_ ,
    \new_[89766]_ , \new_[89769]_ , \new_[89770]_ , \new_[89771]_ ,
    \new_[89774]_ , \new_[89777]_ , \new_[89778]_ , \new_[89781]_ ,
    \new_[89784]_ , \new_[89785]_ , \new_[89786]_ , \new_[89790]_ ,
    \new_[89791]_ , \new_[89794]_ , \new_[89797]_ , \new_[89798]_ ,
    \new_[89799]_ , \new_[89802]_ , \new_[89805]_ , \new_[89806]_ ,
    \new_[89809]_ , \new_[89812]_ , \new_[89813]_ , \new_[89814]_ ,
    \new_[89818]_ , \new_[89819]_ , \new_[89822]_ , \new_[89825]_ ,
    \new_[89826]_ , \new_[89827]_ , \new_[89830]_ , \new_[89833]_ ,
    \new_[89834]_ , \new_[89837]_ , \new_[89840]_ , \new_[89841]_ ,
    \new_[89842]_ , \new_[89846]_ , \new_[89847]_ , \new_[89850]_ ,
    \new_[89853]_ , \new_[89854]_ , \new_[89855]_ , \new_[89858]_ ,
    \new_[89861]_ , \new_[89862]_ , \new_[89865]_ , \new_[89868]_ ,
    \new_[89869]_ , \new_[89870]_ , \new_[89874]_ , \new_[89875]_ ,
    \new_[89878]_ , \new_[89881]_ , \new_[89882]_ , \new_[89883]_ ,
    \new_[89886]_ , \new_[89889]_ , \new_[89890]_ , \new_[89893]_ ,
    \new_[89896]_ , \new_[89897]_ , \new_[89898]_ , \new_[89902]_ ,
    \new_[89903]_ , \new_[89906]_ , \new_[89909]_ , \new_[89910]_ ,
    \new_[89911]_ , \new_[89914]_ , \new_[89917]_ , \new_[89918]_ ,
    \new_[89921]_ , \new_[89924]_ , \new_[89925]_ , \new_[89926]_ ,
    \new_[89930]_ , \new_[89931]_ , \new_[89934]_ , \new_[89937]_ ,
    \new_[89938]_ , \new_[89939]_ , \new_[89942]_ , \new_[89945]_ ,
    \new_[89946]_ , \new_[89949]_ , \new_[89952]_ , \new_[89953]_ ,
    \new_[89954]_ , \new_[89958]_ , \new_[89959]_ , \new_[89962]_ ,
    \new_[89965]_ , \new_[89966]_ , \new_[89967]_ , \new_[89970]_ ,
    \new_[89973]_ , \new_[89974]_ , \new_[89977]_ , \new_[89980]_ ,
    \new_[89981]_ , \new_[89982]_ , \new_[89986]_ , \new_[89987]_ ,
    \new_[89990]_ , \new_[89993]_ , \new_[89994]_ , \new_[89995]_ ,
    \new_[89998]_ , \new_[90001]_ , \new_[90002]_ , \new_[90005]_ ,
    \new_[90008]_ , \new_[90009]_ , \new_[90010]_ , \new_[90014]_ ,
    \new_[90015]_ , \new_[90018]_ , \new_[90021]_ , \new_[90022]_ ,
    \new_[90023]_ , \new_[90026]_ , \new_[90029]_ , \new_[90030]_ ,
    \new_[90033]_ , \new_[90036]_ , \new_[90037]_ , \new_[90038]_ ,
    \new_[90042]_ , \new_[90043]_ , \new_[90046]_ , \new_[90049]_ ,
    \new_[90050]_ , \new_[90051]_ , \new_[90054]_ , \new_[90057]_ ,
    \new_[90058]_ , \new_[90061]_ , \new_[90064]_ , \new_[90065]_ ,
    \new_[90066]_ , \new_[90070]_ , \new_[90071]_ , \new_[90074]_ ,
    \new_[90077]_ , \new_[90078]_ , \new_[90079]_ , \new_[90082]_ ,
    \new_[90085]_ , \new_[90086]_ , \new_[90089]_ , \new_[90092]_ ,
    \new_[90093]_ , \new_[90094]_ , \new_[90098]_ , \new_[90099]_ ,
    \new_[90102]_ , \new_[90105]_ , \new_[90106]_ , \new_[90107]_ ,
    \new_[90110]_ , \new_[90113]_ , \new_[90114]_ , \new_[90117]_ ,
    \new_[90120]_ , \new_[90121]_ , \new_[90122]_ , \new_[90126]_ ,
    \new_[90127]_ , \new_[90130]_ , \new_[90133]_ , \new_[90134]_ ,
    \new_[90135]_ , \new_[90138]_ , \new_[90141]_ , \new_[90142]_ ,
    \new_[90145]_ , \new_[90148]_ , \new_[90149]_ , \new_[90150]_ ,
    \new_[90154]_ , \new_[90155]_ , \new_[90158]_ , \new_[90161]_ ,
    \new_[90162]_ , \new_[90163]_ , \new_[90166]_ , \new_[90169]_ ,
    \new_[90170]_ , \new_[90173]_ , \new_[90176]_ , \new_[90177]_ ,
    \new_[90178]_ , \new_[90182]_ , \new_[90183]_ , \new_[90186]_ ,
    \new_[90189]_ , \new_[90190]_ , \new_[90191]_ , \new_[90194]_ ,
    \new_[90197]_ , \new_[90198]_ , \new_[90201]_ , \new_[90204]_ ,
    \new_[90205]_ , \new_[90206]_ , \new_[90210]_ , \new_[90211]_ ,
    \new_[90214]_ , \new_[90217]_ , \new_[90218]_ , \new_[90219]_ ,
    \new_[90222]_ , \new_[90225]_ , \new_[90226]_ , \new_[90229]_ ,
    \new_[90232]_ , \new_[90233]_ , \new_[90234]_ , \new_[90238]_ ,
    \new_[90239]_ , \new_[90242]_ , \new_[90245]_ , \new_[90246]_ ,
    \new_[90247]_ , \new_[90250]_ , \new_[90253]_ , \new_[90254]_ ,
    \new_[90257]_ , \new_[90260]_ , \new_[90261]_ , \new_[90262]_ ,
    \new_[90266]_ , \new_[90267]_ , \new_[90270]_ , \new_[90273]_ ,
    \new_[90274]_ , \new_[90275]_ , \new_[90278]_ , \new_[90281]_ ,
    \new_[90282]_ , \new_[90285]_ , \new_[90288]_ , \new_[90289]_ ,
    \new_[90290]_ , \new_[90294]_ , \new_[90295]_ , \new_[90298]_ ,
    \new_[90301]_ , \new_[90302]_ , \new_[90303]_ , \new_[90306]_ ,
    \new_[90309]_ , \new_[90310]_ , \new_[90313]_ , \new_[90316]_ ,
    \new_[90317]_ , \new_[90318]_ , \new_[90322]_ , \new_[90323]_ ,
    \new_[90326]_ , \new_[90329]_ , \new_[90330]_ , \new_[90331]_ ,
    \new_[90334]_ , \new_[90337]_ , \new_[90338]_ , \new_[90341]_ ,
    \new_[90344]_ , \new_[90345]_ , \new_[90346]_ , \new_[90350]_ ,
    \new_[90351]_ , \new_[90354]_ , \new_[90357]_ , \new_[90358]_ ,
    \new_[90359]_ , \new_[90362]_ , \new_[90365]_ , \new_[90366]_ ,
    \new_[90369]_ , \new_[90372]_ , \new_[90373]_ , \new_[90374]_ ,
    \new_[90378]_ , \new_[90379]_ , \new_[90382]_ , \new_[90385]_ ,
    \new_[90386]_ , \new_[90387]_ , \new_[90390]_ , \new_[90393]_ ,
    \new_[90394]_ , \new_[90397]_ , \new_[90400]_ , \new_[90401]_ ,
    \new_[90402]_ , \new_[90406]_ , \new_[90407]_ , \new_[90410]_ ,
    \new_[90413]_ , \new_[90414]_ , \new_[90415]_ , \new_[90418]_ ,
    \new_[90421]_ , \new_[90422]_ , \new_[90425]_ , \new_[90428]_ ,
    \new_[90429]_ , \new_[90430]_ , \new_[90434]_ , \new_[90435]_ ,
    \new_[90438]_ , \new_[90441]_ , \new_[90442]_ , \new_[90443]_ ,
    \new_[90446]_ , \new_[90449]_ , \new_[90450]_ , \new_[90453]_ ,
    \new_[90456]_ , \new_[90457]_ , \new_[90458]_ , \new_[90462]_ ,
    \new_[90463]_ , \new_[90466]_ , \new_[90469]_ , \new_[90470]_ ,
    \new_[90471]_ , \new_[90474]_ , \new_[90477]_ , \new_[90478]_ ,
    \new_[90481]_ , \new_[90484]_ , \new_[90485]_ , \new_[90486]_ ,
    \new_[90490]_ , \new_[90491]_ , \new_[90494]_ , \new_[90497]_ ,
    \new_[90498]_ , \new_[90499]_ , \new_[90502]_ , \new_[90505]_ ,
    \new_[90506]_ , \new_[90509]_ , \new_[90512]_ , \new_[90513]_ ,
    \new_[90514]_ , \new_[90518]_ , \new_[90519]_ , \new_[90522]_ ,
    \new_[90525]_ , \new_[90526]_ , \new_[90527]_ , \new_[90530]_ ,
    \new_[90533]_ , \new_[90534]_ , \new_[90537]_ , \new_[90540]_ ,
    \new_[90541]_ , \new_[90542]_ , \new_[90546]_ , \new_[90547]_ ,
    \new_[90550]_ , \new_[90553]_ , \new_[90554]_ , \new_[90555]_ ,
    \new_[90558]_ , \new_[90561]_ , \new_[90562]_ , \new_[90565]_ ,
    \new_[90568]_ , \new_[90569]_ , \new_[90570]_ , \new_[90574]_ ,
    \new_[90575]_ , \new_[90578]_ , \new_[90581]_ , \new_[90582]_ ,
    \new_[90583]_ , \new_[90586]_ , \new_[90589]_ , \new_[90590]_ ,
    \new_[90593]_ , \new_[90596]_ , \new_[90597]_ , \new_[90598]_ ,
    \new_[90602]_ , \new_[90603]_ , \new_[90606]_ , \new_[90609]_ ,
    \new_[90610]_ , \new_[90611]_ , \new_[90614]_ , \new_[90617]_ ,
    \new_[90618]_ , \new_[90621]_ , \new_[90624]_ , \new_[90625]_ ,
    \new_[90626]_ , \new_[90630]_ , \new_[90631]_ , \new_[90634]_ ,
    \new_[90637]_ , \new_[90638]_ , \new_[90639]_ , \new_[90642]_ ,
    \new_[90645]_ , \new_[90646]_ , \new_[90649]_ , \new_[90652]_ ,
    \new_[90653]_ , \new_[90654]_ , \new_[90658]_ , \new_[90659]_ ,
    \new_[90662]_ , \new_[90665]_ , \new_[90666]_ , \new_[90667]_ ,
    \new_[90670]_ , \new_[90673]_ , \new_[90674]_ , \new_[90677]_ ,
    \new_[90680]_ , \new_[90681]_ , \new_[90682]_ , \new_[90686]_ ,
    \new_[90687]_ , \new_[90690]_ , \new_[90693]_ , \new_[90694]_ ,
    \new_[90695]_ , \new_[90698]_ , \new_[90701]_ , \new_[90702]_ ,
    \new_[90705]_ , \new_[90708]_ , \new_[90709]_ , \new_[90710]_ ,
    \new_[90714]_ , \new_[90715]_ , \new_[90718]_ , \new_[90721]_ ,
    \new_[90722]_ , \new_[90723]_ , \new_[90726]_ , \new_[90729]_ ,
    \new_[90730]_ , \new_[90733]_ , \new_[90736]_ , \new_[90737]_ ,
    \new_[90738]_ , \new_[90742]_ , \new_[90743]_ , \new_[90746]_ ,
    \new_[90749]_ , \new_[90750]_ , \new_[90751]_ , \new_[90754]_ ,
    \new_[90757]_ , \new_[90758]_ , \new_[90761]_ , \new_[90764]_ ,
    \new_[90765]_ , \new_[90766]_ , \new_[90770]_ , \new_[90771]_ ,
    \new_[90774]_ , \new_[90777]_ , \new_[90778]_ , \new_[90779]_ ,
    \new_[90782]_ , \new_[90785]_ , \new_[90786]_ , \new_[90789]_ ,
    \new_[90792]_ , \new_[90793]_ , \new_[90794]_ , \new_[90798]_ ,
    \new_[90799]_ , \new_[90802]_ , \new_[90805]_ , \new_[90806]_ ,
    \new_[90807]_ , \new_[90810]_ , \new_[90813]_ , \new_[90814]_ ,
    \new_[90817]_ , \new_[90820]_ , \new_[90821]_ , \new_[90822]_ ,
    \new_[90826]_ , \new_[90827]_ , \new_[90830]_ , \new_[90833]_ ,
    \new_[90834]_ , \new_[90835]_ , \new_[90838]_ , \new_[90841]_ ,
    \new_[90842]_ , \new_[90845]_ , \new_[90848]_ , \new_[90849]_ ,
    \new_[90850]_ , \new_[90854]_ , \new_[90855]_ , \new_[90858]_ ,
    \new_[90861]_ , \new_[90862]_ , \new_[90863]_ , \new_[90866]_ ,
    \new_[90869]_ , \new_[90870]_ , \new_[90873]_ , \new_[90876]_ ,
    \new_[90877]_ , \new_[90878]_ , \new_[90882]_ , \new_[90883]_ ,
    \new_[90886]_ , \new_[90889]_ , \new_[90890]_ , \new_[90891]_ ,
    \new_[90894]_ , \new_[90897]_ , \new_[90898]_ , \new_[90901]_ ,
    \new_[90904]_ , \new_[90905]_ , \new_[90906]_ , \new_[90910]_ ,
    \new_[90911]_ , \new_[90914]_ , \new_[90917]_ , \new_[90918]_ ,
    \new_[90919]_ , \new_[90922]_ , \new_[90925]_ , \new_[90926]_ ,
    \new_[90929]_ , \new_[90932]_ , \new_[90933]_ , \new_[90934]_ ,
    \new_[90938]_ , \new_[90939]_ , \new_[90942]_ , \new_[90945]_ ,
    \new_[90946]_ , \new_[90947]_ , \new_[90950]_ , \new_[90953]_ ,
    \new_[90954]_ , \new_[90957]_ , \new_[90960]_ , \new_[90961]_ ,
    \new_[90962]_ , \new_[90966]_ , \new_[90967]_ , \new_[90970]_ ,
    \new_[90973]_ , \new_[90974]_ , \new_[90975]_ , \new_[90978]_ ,
    \new_[90981]_ , \new_[90982]_ , \new_[90985]_ , \new_[90988]_ ,
    \new_[90989]_ , \new_[90990]_ , \new_[90994]_ , \new_[90995]_ ,
    \new_[90998]_ , \new_[91001]_ , \new_[91002]_ , \new_[91003]_ ,
    \new_[91006]_ , \new_[91009]_ , \new_[91010]_ , \new_[91013]_ ,
    \new_[91016]_ , \new_[91017]_ , \new_[91018]_ , \new_[91022]_ ,
    \new_[91023]_ , \new_[91026]_ , \new_[91029]_ , \new_[91030]_ ,
    \new_[91031]_ , \new_[91034]_ , \new_[91037]_ , \new_[91038]_ ,
    \new_[91041]_ , \new_[91044]_ , \new_[91045]_ , \new_[91046]_ ,
    \new_[91050]_ , \new_[91051]_ , \new_[91054]_ , \new_[91057]_ ,
    \new_[91058]_ , \new_[91059]_ , \new_[91062]_ , \new_[91065]_ ,
    \new_[91066]_ , \new_[91069]_ , \new_[91072]_ , \new_[91073]_ ,
    \new_[91074]_ , \new_[91078]_ , \new_[91079]_ , \new_[91082]_ ,
    \new_[91085]_ , \new_[91086]_ , \new_[91087]_ , \new_[91090]_ ,
    \new_[91093]_ , \new_[91094]_ , \new_[91097]_ , \new_[91100]_ ,
    \new_[91101]_ , \new_[91102]_ , \new_[91106]_ , \new_[91107]_ ,
    \new_[91110]_ , \new_[91113]_ , \new_[91114]_ , \new_[91115]_ ,
    \new_[91118]_ , \new_[91121]_ , \new_[91122]_ , \new_[91125]_ ,
    \new_[91128]_ , \new_[91129]_ , \new_[91130]_ , \new_[91134]_ ,
    \new_[91135]_ , \new_[91138]_ , \new_[91141]_ , \new_[91142]_ ,
    \new_[91143]_ , \new_[91146]_ , \new_[91149]_ , \new_[91150]_ ,
    \new_[91153]_ , \new_[91156]_ , \new_[91157]_ , \new_[91158]_ ,
    \new_[91162]_ , \new_[91163]_ , \new_[91166]_ , \new_[91169]_ ,
    \new_[91170]_ , \new_[91171]_ , \new_[91174]_ , \new_[91177]_ ,
    \new_[91178]_ , \new_[91181]_ , \new_[91184]_ , \new_[91185]_ ,
    \new_[91186]_ , \new_[91190]_ , \new_[91191]_ , \new_[91194]_ ,
    \new_[91197]_ , \new_[91198]_ , \new_[91199]_ , \new_[91202]_ ,
    \new_[91205]_ , \new_[91206]_ , \new_[91209]_ , \new_[91212]_ ,
    \new_[91213]_ , \new_[91214]_ , \new_[91218]_ , \new_[91219]_ ,
    \new_[91222]_ , \new_[91225]_ , \new_[91226]_ , \new_[91227]_ ,
    \new_[91230]_ , \new_[91233]_ , \new_[91234]_ , \new_[91237]_ ,
    \new_[91240]_ , \new_[91241]_ , \new_[91242]_ , \new_[91246]_ ,
    \new_[91247]_ , \new_[91250]_ , \new_[91253]_ , \new_[91254]_ ,
    \new_[91255]_ , \new_[91258]_ , \new_[91261]_ , \new_[91262]_ ,
    \new_[91265]_ , \new_[91268]_ , \new_[91269]_ , \new_[91270]_ ,
    \new_[91274]_ , \new_[91275]_ , \new_[91278]_ , \new_[91281]_ ,
    \new_[91282]_ , \new_[91283]_ , \new_[91286]_ , \new_[91289]_ ,
    \new_[91290]_ , \new_[91293]_ , \new_[91296]_ , \new_[91297]_ ,
    \new_[91298]_ , \new_[91302]_ , \new_[91303]_ , \new_[91306]_ ,
    \new_[91309]_ , \new_[91310]_ , \new_[91311]_ , \new_[91314]_ ,
    \new_[91317]_ , \new_[91318]_ , \new_[91321]_ , \new_[91324]_ ,
    \new_[91325]_ , \new_[91326]_ , \new_[91330]_ , \new_[91331]_ ,
    \new_[91334]_ , \new_[91337]_ , \new_[91338]_ , \new_[91339]_ ,
    \new_[91342]_ , \new_[91345]_ , \new_[91346]_ , \new_[91349]_ ,
    \new_[91352]_ , \new_[91353]_ , \new_[91354]_ , \new_[91358]_ ,
    \new_[91359]_ , \new_[91362]_ , \new_[91365]_ , \new_[91366]_ ,
    \new_[91367]_ , \new_[91370]_ , \new_[91373]_ , \new_[91374]_ ,
    \new_[91377]_ , \new_[91380]_ , \new_[91381]_ , \new_[91382]_ ,
    \new_[91386]_ , \new_[91387]_ , \new_[91390]_ , \new_[91393]_ ,
    \new_[91394]_ , \new_[91395]_ , \new_[91398]_ , \new_[91401]_ ,
    \new_[91402]_ , \new_[91405]_ , \new_[91408]_ , \new_[91409]_ ,
    \new_[91410]_ , \new_[91414]_ , \new_[91415]_ , \new_[91418]_ ,
    \new_[91421]_ , \new_[91422]_ , \new_[91423]_ , \new_[91426]_ ,
    \new_[91429]_ , \new_[91430]_ , \new_[91433]_ , \new_[91436]_ ,
    \new_[91437]_ , \new_[91438]_ , \new_[91442]_ , \new_[91443]_ ,
    \new_[91446]_ , \new_[91449]_ , \new_[91450]_ , \new_[91451]_ ,
    \new_[91454]_ , \new_[91457]_ , \new_[91458]_ , \new_[91461]_ ,
    \new_[91464]_ , \new_[91465]_ , \new_[91466]_ , \new_[91470]_ ,
    \new_[91471]_ , \new_[91474]_ , \new_[91477]_ , \new_[91478]_ ,
    \new_[91479]_ , \new_[91482]_ , \new_[91485]_ , \new_[91486]_ ,
    \new_[91489]_ , \new_[91492]_ , \new_[91493]_ , \new_[91494]_ ,
    \new_[91498]_ , \new_[91499]_ , \new_[91502]_ , \new_[91505]_ ,
    \new_[91506]_ , \new_[91507]_ , \new_[91510]_ , \new_[91513]_ ,
    \new_[91514]_ , \new_[91517]_ , \new_[91520]_ , \new_[91521]_ ,
    \new_[91522]_ , \new_[91526]_ , \new_[91527]_ , \new_[91530]_ ,
    \new_[91533]_ , \new_[91534]_ , \new_[91535]_ , \new_[91538]_ ,
    \new_[91541]_ , \new_[91542]_ , \new_[91545]_ , \new_[91548]_ ,
    \new_[91549]_ , \new_[91550]_ , \new_[91554]_ , \new_[91555]_ ,
    \new_[91558]_ , \new_[91561]_ , \new_[91562]_ , \new_[91563]_ ,
    \new_[91566]_ , \new_[91569]_ , \new_[91570]_ , \new_[91573]_ ,
    \new_[91576]_ , \new_[91577]_ , \new_[91578]_ , \new_[91582]_ ,
    \new_[91583]_ , \new_[91586]_ , \new_[91589]_ , \new_[91590]_ ,
    \new_[91591]_ , \new_[91594]_ , \new_[91597]_ , \new_[91598]_ ,
    \new_[91601]_ , \new_[91604]_ , \new_[91605]_ , \new_[91606]_ ,
    \new_[91610]_ , \new_[91611]_ , \new_[91614]_ , \new_[91617]_ ,
    \new_[91618]_ , \new_[91619]_ , \new_[91622]_ , \new_[91625]_ ,
    \new_[91626]_ , \new_[91629]_ , \new_[91632]_ , \new_[91633]_ ,
    \new_[91634]_ , \new_[91638]_ , \new_[91639]_ , \new_[91642]_ ,
    \new_[91645]_ , \new_[91646]_ , \new_[91647]_ , \new_[91650]_ ,
    \new_[91653]_ , \new_[91654]_ , \new_[91657]_ , \new_[91660]_ ,
    \new_[91661]_ , \new_[91662]_ , \new_[91666]_ , \new_[91667]_ ,
    \new_[91670]_ , \new_[91673]_ , \new_[91674]_ , \new_[91675]_ ,
    \new_[91678]_ , \new_[91681]_ , \new_[91682]_ , \new_[91685]_ ,
    \new_[91688]_ , \new_[91689]_ , \new_[91690]_ , \new_[91694]_ ,
    \new_[91695]_ , \new_[91698]_ , \new_[91701]_ , \new_[91702]_ ,
    \new_[91703]_ , \new_[91706]_ , \new_[91709]_ , \new_[91710]_ ,
    \new_[91713]_ , \new_[91716]_ , \new_[91717]_ , \new_[91718]_ ,
    \new_[91722]_ , \new_[91723]_ , \new_[91726]_ , \new_[91729]_ ,
    \new_[91730]_ , \new_[91731]_ , \new_[91734]_ , \new_[91737]_ ,
    \new_[91738]_ , \new_[91741]_ , \new_[91744]_ , \new_[91745]_ ,
    \new_[91746]_ , \new_[91750]_ , \new_[91751]_ , \new_[91754]_ ,
    \new_[91757]_ , \new_[91758]_ , \new_[91759]_ , \new_[91762]_ ,
    \new_[91765]_ , \new_[91766]_ , \new_[91769]_ , \new_[91772]_ ,
    \new_[91773]_ , \new_[91774]_ , \new_[91778]_ , \new_[91779]_ ,
    \new_[91782]_ , \new_[91785]_ , \new_[91786]_ , \new_[91787]_ ,
    \new_[91790]_ , \new_[91793]_ , \new_[91794]_ , \new_[91797]_ ,
    \new_[91800]_ , \new_[91801]_ , \new_[91802]_ , \new_[91806]_ ,
    \new_[91807]_ , \new_[91810]_ , \new_[91813]_ , \new_[91814]_ ,
    \new_[91815]_ , \new_[91818]_ , \new_[91821]_ , \new_[91822]_ ,
    \new_[91825]_ , \new_[91828]_ , \new_[91829]_ , \new_[91830]_ ,
    \new_[91834]_ , \new_[91835]_ , \new_[91838]_ , \new_[91841]_ ,
    \new_[91842]_ , \new_[91843]_ , \new_[91846]_ , \new_[91849]_ ,
    \new_[91850]_ , \new_[91853]_ , \new_[91856]_ , \new_[91857]_ ,
    \new_[91858]_ , \new_[91862]_ , \new_[91863]_ , \new_[91866]_ ,
    \new_[91869]_ , \new_[91870]_ , \new_[91871]_ , \new_[91874]_ ,
    \new_[91877]_ , \new_[91878]_ , \new_[91881]_ , \new_[91884]_ ,
    \new_[91885]_ , \new_[91886]_ , \new_[91890]_ , \new_[91891]_ ,
    \new_[91894]_ , \new_[91897]_ , \new_[91898]_ , \new_[91899]_ ,
    \new_[91902]_ , \new_[91905]_ , \new_[91906]_ , \new_[91909]_ ,
    \new_[91912]_ , \new_[91913]_ , \new_[91914]_ , \new_[91918]_ ,
    \new_[91919]_ , \new_[91922]_ , \new_[91925]_ , \new_[91926]_ ,
    \new_[91927]_ , \new_[91930]_ , \new_[91933]_ , \new_[91934]_ ,
    \new_[91937]_ , \new_[91940]_ , \new_[91941]_ , \new_[91942]_ ,
    \new_[91946]_ , \new_[91947]_ , \new_[91950]_ , \new_[91953]_ ,
    \new_[91954]_ , \new_[91955]_ , \new_[91958]_ , \new_[91961]_ ,
    \new_[91962]_ , \new_[91965]_ , \new_[91968]_ , \new_[91969]_ ,
    \new_[91970]_ , \new_[91974]_ , \new_[91975]_ , \new_[91978]_ ,
    \new_[91981]_ , \new_[91982]_ , \new_[91983]_ , \new_[91986]_ ,
    \new_[91989]_ , \new_[91990]_ , \new_[91993]_ , \new_[91996]_ ,
    \new_[91997]_ , \new_[91998]_ , \new_[92002]_ , \new_[92003]_ ,
    \new_[92006]_ , \new_[92009]_ , \new_[92010]_ , \new_[92011]_ ,
    \new_[92014]_ , \new_[92017]_ , \new_[92018]_ , \new_[92021]_ ,
    \new_[92024]_ , \new_[92025]_ , \new_[92026]_ , \new_[92030]_ ,
    \new_[92031]_ , \new_[92034]_ , \new_[92037]_ , \new_[92038]_ ,
    \new_[92039]_ , \new_[92042]_ , \new_[92045]_ , \new_[92046]_ ,
    \new_[92049]_ , \new_[92052]_ , \new_[92053]_ , \new_[92054]_ ,
    \new_[92058]_ , \new_[92059]_ , \new_[92062]_ , \new_[92065]_ ,
    \new_[92066]_ , \new_[92067]_ , \new_[92070]_ , \new_[92073]_ ,
    \new_[92074]_ , \new_[92077]_ , \new_[92080]_ , \new_[92081]_ ,
    \new_[92082]_ , \new_[92086]_ , \new_[92087]_ , \new_[92090]_ ,
    \new_[92093]_ , \new_[92094]_ , \new_[92095]_ , \new_[92098]_ ,
    \new_[92101]_ , \new_[92102]_ , \new_[92105]_ , \new_[92108]_ ,
    \new_[92109]_ , \new_[92110]_ , \new_[92114]_ , \new_[92115]_ ,
    \new_[92118]_ , \new_[92121]_ , \new_[92122]_ , \new_[92123]_ ,
    \new_[92126]_ , \new_[92129]_ , \new_[92130]_ , \new_[92133]_ ,
    \new_[92136]_ , \new_[92137]_ , \new_[92138]_ , \new_[92142]_ ,
    \new_[92143]_ , \new_[92146]_ , \new_[92149]_ , \new_[92150]_ ,
    \new_[92151]_ , \new_[92154]_ , \new_[92157]_ , \new_[92158]_ ,
    \new_[92161]_ , \new_[92164]_ , \new_[92165]_ , \new_[92166]_ ,
    \new_[92170]_ , \new_[92171]_ , \new_[92174]_ , \new_[92177]_ ,
    \new_[92178]_ , \new_[92179]_ , \new_[92182]_ , \new_[92185]_ ,
    \new_[92186]_ , \new_[92189]_ , \new_[92192]_ , \new_[92193]_ ,
    \new_[92194]_ , \new_[92198]_ , \new_[92199]_ , \new_[92202]_ ,
    \new_[92205]_ , \new_[92206]_ , \new_[92207]_ , \new_[92210]_ ,
    \new_[92213]_ , \new_[92214]_ , \new_[92217]_ , \new_[92220]_ ,
    \new_[92221]_ , \new_[92222]_ , \new_[92226]_ , \new_[92227]_ ,
    \new_[92230]_ , \new_[92233]_ , \new_[92234]_ , \new_[92235]_ ,
    \new_[92238]_ , \new_[92241]_ , \new_[92242]_ , \new_[92245]_ ,
    \new_[92248]_ , \new_[92249]_ , \new_[92250]_ , \new_[92254]_ ,
    \new_[92255]_ , \new_[92258]_ , \new_[92261]_ , \new_[92262]_ ,
    \new_[92263]_ , \new_[92266]_ , \new_[92269]_ , \new_[92270]_ ,
    \new_[92273]_ , \new_[92276]_ , \new_[92277]_ , \new_[92278]_ ,
    \new_[92282]_ , \new_[92283]_ , \new_[92286]_ , \new_[92289]_ ,
    \new_[92290]_ , \new_[92291]_ , \new_[92294]_ , \new_[92297]_ ,
    \new_[92298]_ , \new_[92301]_ , \new_[92304]_ , \new_[92305]_ ,
    \new_[92306]_ , \new_[92310]_ , \new_[92311]_ , \new_[92314]_ ,
    \new_[92317]_ , \new_[92318]_ , \new_[92319]_ , \new_[92322]_ ,
    \new_[92325]_ , \new_[92326]_ , \new_[92329]_ , \new_[92332]_ ,
    \new_[92333]_ , \new_[92334]_ , \new_[92338]_ , \new_[92339]_ ,
    \new_[92342]_ , \new_[92345]_ , \new_[92346]_ , \new_[92347]_ ,
    \new_[92350]_ , \new_[92353]_ , \new_[92354]_ , \new_[92357]_ ,
    \new_[92360]_ , \new_[92361]_ , \new_[92362]_ , \new_[92366]_ ,
    \new_[92367]_ , \new_[92370]_ , \new_[92373]_ , \new_[92374]_ ,
    \new_[92375]_ , \new_[92378]_ , \new_[92381]_ , \new_[92382]_ ,
    \new_[92385]_ , \new_[92388]_ , \new_[92389]_ , \new_[92390]_ ,
    \new_[92394]_ , \new_[92395]_ , \new_[92398]_ , \new_[92401]_ ,
    \new_[92402]_ , \new_[92403]_ , \new_[92406]_ , \new_[92409]_ ,
    \new_[92410]_ , \new_[92413]_ , \new_[92416]_ , \new_[92417]_ ,
    \new_[92418]_ , \new_[92422]_ , \new_[92423]_ , \new_[92426]_ ,
    \new_[92429]_ , \new_[92430]_ , \new_[92431]_ , \new_[92434]_ ,
    \new_[92437]_ , \new_[92438]_ , \new_[92441]_ , \new_[92444]_ ,
    \new_[92445]_ , \new_[92446]_ , \new_[92450]_ , \new_[92451]_ ,
    \new_[92454]_ , \new_[92457]_ , \new_[92458]_ , \new_[92459]_ ,
    \new_[92462]_ , \new_[92465]_ , \new_[92466]_ , \new_[92469]_ ,
    \new_[92472]_ , \new_[92473]_ , \new_[92474]_ , \new_[92478]_ ,
    \new_[92479]_ , \new_[92482]_ , \new_[92485]_ , \new_[92486]_ ,
    \new_[92487]_ , \new_[92490]_ , \new_[92493]_ , \new_[92494]_ ,
    \new_[92497]_ , \new_[92500]_ , \new_[92501]_ , \new_[92502]_ ,
    \new_[92506]_ , \new_[92507]_ , \new_[92510]_ , \new_[92513]_ ,
    \new_[92514]_ , \new_[92515]_ , \new_[92518]_ , \new_[92521]_ ,
    \new_[92522]_ , \new_[92525]_ , \new_[92528]_ , \new_[92529]_ ,
    \new_[92530]_ , \new_[92534]_ , \new_[92535]_ , \new_[92538]_ ,
    \new_[92541]_ , \new_[92542]_ , \new_[92543]_ , \new_[92546]_ ,
    \new_[92549]_ , \new_[92550]_ , \new_[92553]_ , \new_[92556]_ ,
    \new_[92557]_ , \new_[92558]_ , \new_[92562]_ , \new_[92563]_ ,
    \new_[92566]_ , \new_[92569]_ , \new_[92570]_ , \new_[92571]_ ,
    \new_[92574]_ , \new_[92577]_ , \new_[92578]_ , \new_[92581]_ ,
    \new_[92584]_ , \new_[92585]_ , \new_[92586]_ , \new_[92590]_ ,
    \new_[92591]_ , \new_[92594]_ , \new_[92597]_ , \new_[92598]_ ,
    \new_[92599]_ , \new_[92602]_ , \new_[92605]_ , \new_[92606]_ ,
    \new_[92609]_ , \new_[92612]_ , \new_[92613]_ , \new_[92614]_ ,
    \new_[92618]_ , \new_[92619]_ , \new_[92622]_ , \new_[92625]_ ,
    \new_[92626]_ , \new_[92627]_ , \new_[92630]_ , \new_[92633]_ ,
    \new_[92634]_ , \new_[92637]_ , \new_[92640]_ , \new_[92641]_ ,
    \new_[92642]_ , \new_[92646]_ , \new_[92647]_ , \new_[92650]_ ,
    \new_[92653]_ , \new_[92654]_ , \new_[92655]_ , \new_[92658]_ ,
    \new_[92661]_ , \new_[92662]_ , \new_[92665]_ , \new_[92668]_ ,
    \new_[92669]_ , \new_[92670]_ , \new_[92674]_ , \new_[92675]_ ,
    \new_[92678]_ , \new_[92681]_ , \new_[92682]_ , \new_[92683]_ ,
    \new_[92686]_ , \new_[92689]_ , \new_[92690]_ , \new_[92693]_ ,
    \new_[92696]_ , \new_[92697]_ , \new_[92698]_ , \new_[92702]_ ,
    \new_[92703]_ , \new_[92706]_ , \new_[92709]_ , \new_[92710]_ ,
    \new_[92711]_ , \new_[92714]_ , \new_[92717]_ , \new_[92718]_ ,
    \new_[92721]_ , \new_[92724]_ , \new_[92725]_ , \new_[92726]_ ,
    \new_[92730]_ , \new_[92731]_ , \new_[92734]_ , \new_[92737]_ ,
    \new_[92738]_ , \new_[92739]_ , \new_[92742]_ , \new_[92745]_ ,
    \new_[92746]_ , \new_[92749]_ , \new_[92752]_ , \new_[92753]_ ,
    \new_[92754]_ , \new_[92758]_ , \new_[92759]_ , \new_[92762]_ ,
    \new_[92765]_ , \new_[92766]_ , \new_[92767]_ , \new_[92770]_ ,
    \new_[92773]_ , \new_[92774]_ , \new_[92777]_ , \new_[92780]_ ,
    \new_[92781]_ , \new_[92782]_ , \new_[92786]_ , \new_[92787]_ ,
    \new_[92790]_ , \new_[92793]_ , \new_[92794]_ , \new_[92795]_ ,
    \new_[92798]_ , \new_[92801]_ , \new_[92802]_ , \new_[92805]_ ,
    \new_[92808]_ , \new_[92809]_ , \new_[92810]_ , \new_[92814]_ ,
    \new_[92815]_ , \new_[92818]_ , \new_[92821]_ , \new_[92822]_ ,
    \new_[92823]_ , \new_[92826]_ , \new_[92829]_ , \new_[92830]_ ,
    \new_[92833]_ , \new_[92836]_ , \new_[92837]_ , \new_[92838]_ ,
    \new_[92842]_ , \new_[92843]_ , \new_[92846]_ , \new_[92849]_ ,
    \new_[92850]_ , \new_[92851]_ , \new_[92854]_ , \new_[92857]_ ,
    \new_[92858]_ , \new_[92861]_ , \new_[92864]_ , \new_[92865]_ ,
    \new_[92866]_ , \new_[92870]_ , \new_[92871]_ , \new_[92874]_ ,
    \new_[92877]_ , \new_[92878]_ , \new_[92879]_ , \new_[92882]_ ,
    \new_[92885]_ , \new_[92886]_ , \new_[92889]_ , \new_[92892]_ ,
    \new_[92893]_ , \new_[92894]_ , \new_[92898]_ , \new_[92899]_ ,
    \new_[92902]_ , \new_[92905]_ , \new_[92906]_ , \new_[92907]_ ,
    \new_[92910]_ , \new_[92913]_ , \new_[92914]_ , \new_[92917]_ ,
    \new_[92920]_ , \new_[92921]_ , \new_[92922]_ , \new_[92926]_ ,
    \new_[92927]_ , \new_[92930]_ , \new_[92933]_ , \new_[92934]_ ,
    \new_[92935]_ , \new_[92938]_ , \new_[92941]_ , \new_[92942]_ ,
    \new_[92945]_ , \new_[92948]_ , \new_[92949]_ , \new_[92950]_ ,
    \new_[92954]_ , \new_[92955]_ , \new_[92958]_ , \new_[92961]_ ,
    \new_[92962]_ , \new_[92963]_ , \new_[92966]_ , \new_[92969]_ ,
    \new_[92970]_ , \new_[92973]_ , \new_[92976]_ , \new_[92977]_ ,
    \new_[92978]_ , \new_[92982]_ , \new_[92983]_ , \new_[92986]_ ,
    \new_[92989]_ , \new_[92990]_ , \new_[92991]_ , \new_[92994]_ ,
    \new_[92997]_ , \new_[92998]_ , \new_[93001]_ , \new_[93004]_ ,
    \new_[93005]_ , \new_[93006]_ , \new_[93010]_ , \new_[93011]_ ,
    \new_[93014]_ , \new_[93017]_ , \new_[93018]_ , \new_[93019]_ ,
    \new_[93022]_ , \new_[93025]_ , \new_[93026]_ , \new_[93029]_ ,
    \new_[93032]_ , \new_[93033]_ , \new_[93034]_ , \new_[93038]_ ,
    \new_[93039]_ , \new_[93042]_ , \new_[93045]_ , \new_[93046]_ ,
    \new_[93047]_ , \new_[93050]_ , \new_[93053]_ , \new_[93054]_ ,
    \new_[93057]_ , \new_[93060]_ , \new_[93061]_ , \new_[93062]_ ,
    \new_[93066]_ , \new_[93067]_ , \new_[93070]_ , \new_[93073]_ ,
    \new_[93074]_ , \new_[93075]_ , \new_[93078]_ , \new_[93081]_ ,
    \new_[93082]_ , \new_[93085]_ , \new_[93088]_ , \new_[93089]_ ,
    \new_[93090]_ , \new_[93094]_ , \new_[93095]_ , \new_[93098]_ ,
    \new_[93101]_ , \new_[93102]_ , \new_[93103]_ , \new_[93106]_ ,
    \new_[93109]_ , \new_[93110]_ , \new_[93113]_ , \new_[93116]_ ,
    \new_[93117]_ , \new_[93118]_ , \new_[93122]_ , \new_[93123]_ ,
    \new_[93126]_ , \new_[93129]_ , \new_[93130]_ , \new_[93131]_ ,
    \new_[93134]_ , \new_[93137]_ , \new_[93138]_ , \new_[93141]_ ,
    \new_[93144]_ , \new_[93145]_ , \new_[93146]_ , \new_[93150]_ ,
    \new_[93151]_ , \new_[93154]_ , \new_[93157]_ , \new_[93158]_ ,
    \new_[93159]_ , \new_[93162]_ , \new_[93165]_ , \new_[93166]_ ,
    \new_[93169]_ , \new_[93172]_ , \new_[93173]_ , \new_[93174]_ ,
    \new_[93178]_ , \new_[93179]_ , \new_[93182]_ , \new_[93185]_ ,
    \new_[93186]_ , \new_[93187]_ , \new_[93190]_ , \new_[93193]_ ,
    \new_[93194]_ , \new_[93197]_ , \new_[93200]_ , \new_[93201]_ ,
    \new_[93202]_ , \new_[93206]_ , \new_[93207]_ , \new_[93210]_ ,
    \new_[93213]_ , \new_[93214]_ , \new_[93215]_ , \new_[93218]_ ,
    \new_[93221]_ , \new_[93222]_ , \new_[93225]_ , \new_[93228]_ ,
    \new_[93229]_ , \new_[93230]_ , \new_[93234]_ , \new_[93235]_ ,
    \new_[93238]_ , \new_[93241]_ , \new_[93242]_ , \new_[93243]_ ,
    \new_[93246]_ , \new_[93249]_ , \new_[93250]_ , \new_[93253]_ ,
    \new_[93256]_ , \new_[93257]_ , \new_[93258]_ , \new_[93262]_ ,
    \new_[93263]_ , \new_[93266]_ , \new_[93269]_ , \new_[93270]_ ,
    \new_[93271]_ , \new_[93274]_ , \new_[93277]_ , \new_[93278]_ ,
    \new_[93281]_ , \new_[93284]_ , \new_[93285]_ , \new_[93286]_ ,
    \new_[93290]_ , \new_[93291]_ , \new_[93294]_ , \new_[93297]_ ,
    \new_[93298]_ , \new_[93299]_ , \new_[93302]_ , \new_[93305]_ ,
    \new_[93306]_ , \new_[93309]_ , \new_[93312]_ , \new_[93313]_ ,
    \new_[93314]_ , \new_[93318]_ , \new_[93319]_ , \new_[93322]_ ,
    \new_[93325]_ , \new_[93326]_ , \new_[93327]_ , \new_[93330]_ ,
    \new_[93333]_ , \new_[93334]_ , \new_[93337]_ , \new_[93340]_ ,
    \new_[93341]_ , \new_[93342]_ , \new_[93346]_ , \new_[93347]_ ,
    \new_[93350]_ , \new_[93353]_ , \new_[93354]_ , \new_[93355]_ ,
    \new_[93358]_ , \new_[93361]_ , \new_[93362]_ , \new_[93365]_ ,
    \new_[93368]_ , \new_[93369]_ , \new_[93370]_ , \new_[93374]_ ,
    \new_[93375]_ , \new_[93378]_ , \new_[93381]_ , \new_[93382]_ ,
    \new_[93383]_ , \new_[93386]_ , \new_[93389]_ , \new_[93390]_ ,
    \new_[93393]_ , \new_[93396]_ , \new_[93397]_ , \new_[93398]_ ,
    \new_[93402]_ , \new_[93403]_ , \new_[93406]_ , \new_[93409]_ ,
    \new_[93410]_ , \new_[93411]_ , \new_[93414]_ , \new_[93417]_ ,
    \new_[93418]_ , \new_[93421]_ , \new_[93424]_ , \new_[93425]_ ,
    \new_[93426]_ , \new_[93430]_ , \new_[93431]_ , \new_[93434]_ ,
    \new_[93437]_ , \new_[93438]_ , \new_[93439]_ , \new_[93442]_ ,
    \new_[93445]_ , \new_[93446]_ , \new_[93449]_ , \new_[93452]_ ,
    \new_[93453]_ , \new_[93454]_ , \new_[93458]_ , \new_[93459]_ ,
    \new_[93462]_ , \new_[93465]_ , \new_[93466]_ , \new_[93467]_ ,
    \new_[93470]_ , \new_[93473]_ , \new_[93474]_ , \new_[93477]_ ,
    \new_[93480]_ , \new_[93481]_ , \new_[93482]_ , \new_[93486]_ ,
    \new_[93487]_ , \new_[93490]_ , \new_[93493]_ , \new_[93494]_ ,
    \new_[93495]_ , \new_[93498]_ , \new_[93501]_ , \new_[93502]_ ,
    \new_[93505]_ , \new_[93508]_ , \new_[93509]_ , \new_[93510]_ ,
    \new_[93514]_ , \new_[93515]_ , \new_[93518]_ , \new_[93521]_ ,
    \new_[93522]_ , \new_[93523]_ , \new_[93526]_ , \new_[93529]_ ,
    \new_[93530]_ , \new_[93533]_ , \new_[93536]_ , \new_[93537]_ ,
    \new_[93538]_ , \new_[93542]_ , \new_[93543]_ , \new_[93546]_ ,
    \new_[93549]_ , \new_[93550]_ , \new_[93551]_ , \new_[93554]_ ,
    \new_[93557]_ , \new_[93558]_ , \new_[93561]_ , \new_[93564]_ ,
    \new_[93565]_ , \new_[93566]_ , \new_[93570]_ , \new_[93571]_ ,
    \new_[93574]_ , \new_[93577]_ , \new_[93578]_ , \new_[93579]_ ,
    \new_[93582]_ , \new_[93585]_ , \new_[93586]_ , \new_[93589]_ ,
    \new_[93592]_ , \new_[93593]_ , \new_[93594]_ , \new_[93598]_ ,
    \new_[93599]_ , \new_[93602]_ , \new_[93605]_ , \new_[93606]_ ,
    \new_[93607]_ , \new_[93610]_ , \new_[93613]_ , \new_[93614]_ ,
    \new_[93617]_ , \new_[93620]_ , \new_[93621]_ , \new_[93622]_ ,
    \new_[93626]_ , \new_[93627]_ , \new_[93630]_ , \new_[93633]_ ,
    \new_[93634]_ , \new_[93635]_ , \new_[93638]_ , \new_[93641]_ ,
    \new_[93642]_ , \new_[93645]_ , \new_[93648]_ , \new_[93649]_ ,
    \new_[93650]_ , \new_[93654]_ , \new_[93655]_ , \new_[93658]_ ,
    \new_[93661]_ , \new_[93662]_ , \new_[93663]_ , \new_[93666]_ ,
    \new_[93669]_ , \new_[93670]_ , \new_[93673]_ , \new_[93676]_ ,
    \new_[93677]_ , \new_[93678]_ , \new_[93682]_ , \new_[93683]_ ,
    \new_[93686]_ , \new_[93689]_ , \new_[93690]_ , \new_[93691]_ ,
    \new_[93694]_ , \new_[93697]_ , \new_[93698]_ , \new_[93701]_ ,
    \new_[93704]_ , \new_[93705]_ , \new_[93706]_ , \new_[93710]_ ,
    \new_[93711]_ , \new_[93714]_ , \new_[93717]_ , \new_[93718]_ ,
    \new_[93719]_ , \new_[93722]_ , \new_[93725]_ , \new_[93726]_ ,
    \new_[93729]_ , \new_[93732]_ , \new_[93733]_ , \new_[93734]_ ,
    \new_[93738]_ , \new_[93739]_ , \new_[93742]_ , \new_[93745]_ ,
    \new_[93746]_ , \new_[93747]_ , \new_[93750]_ , \new_[93753]_ ,
    \new_[93754]_ , \new_[93757]_ , \new_[93760]_ , \new_[93761]_ ,
    \new_[93762]_ , \new_[93766]_ , \new_[93767]_ , \new_[93770]_ ,
    \new_[93773]_ , \new_[93774]_ , \new_[93775]_ , \new_[93778]_ ,
    \new_[93781]_ , \new_[93782]_ , \new_[93785]_ , \new_[93788]_ ,
    \new_[93789]_ , \new_[93790]_ , \new_[93794]_ , \new_[93795]_ ,
    \new_[93798]_ , \new_[93801]_ , \new_[93802]_ , \new_[93803]_ ,
    \new_[93806]_ , \new_[93809]_ , \new_[93810]_ , \new_[93813]_ ,
    \new_[93816]_ , \new_[93817]_ , \new_[93818]_ , \new_[93822]_ ,
    \new_[93823]_ , \new_[93826]_ , \new_[93829]_ , \new_[93830]_ ,
    \new_[93831]_ , \new_[93834]_ , \new_[93837]_ , \new_[93838]_ ,
    \new_[93841]_ , \new_[93844]_ , \new_[93845]_ , \new_[93846]_ ,
    \new_[93850]_ , \new_[93851]_ , \new_[93854]_ , \new_[93857]_ ,
    \new_[93858]_ , \new_[93859]_ , \new_[93862]_ , \new_[93865]_ ,
    \new_[93866]_ , \new_[93869]_ , \new_[93872]_ , \new_[93873]_ ,
    \new_[93874]_ , \new_[93878]_ , \new_[93879]_ , \new_[93882]_ ,
    \new_[93885]_ , \new_[93886]_ , \new_[93887]_ , \new_[93890]_ ,
    \new_[93893]_ , \new_[93894]_ , \new_[93897]_ , \new_[93900]_ ,
    \new_[93901]_ , \new_[93902]_ , \new_[93906]_ , \new_[93907]_ ,
    \new_[93910]_ , \new_[93913]_ , \new_[93914]_ , \new_[93915]_ ,
    \new_[93918]_ , \new_[93921]_ , \new_[93922]_ , \new_[93925]_ ,
    \new_[93928]_ , \new_[93929]_ , \new_[93930]_ , \new_[93934]_ ,
    \new_[93935]_ , \new_[93938]_ , \new_[93941]_ , \new_[93942]_ ,
    \new_[93943]_ , \new_[93946]_ , \new_[93949]_ , \new_[93950]_ ,
    \new_[93953]_ , \new_[93956]_ , \new_[93957]_ , \new_[93958]_ ,
    \new_[93962]_ , \new_[93963]_ , \new_[93966]_ , \new_[93969]_ ,
    \new_[93970]_ , \new_[93971]_ , \new_[93974]_ , \new_[93977]_ ,
    \new_[93978]_ , \new_[93981]_ , \new_[93984]_ , \new_[93985]_ ,
    \new_[93986]_ , \new_[93990]_ , \new_[93991]_ , \new_[93994]_ ,
    \new_[93997]_ , \new_[93998]_ , \new_[93999]_ , \new_[94002]_ ,
    \new_[94005]_ , \new_[94006]_ , \new_[94009]_ , \new_[94012]_ ,
    \new_[94013]_ , \new_[94014]_ , \new_[94018]_ , \new_[94019]_ ,
    \new_[94022]_ , \new_[94025]_ , \new_[94026]_ , \new_[94027]_ ,
    \new_[94030]_ , \new_[94033]_ , \new_[94034]_ , \new_[94037]_ ,
    \new_[94040]_ , \new_[94041]_ , \new_[94042]_ , \new_[94046]_ ,
    \new_[94047]_ , \new_[94050]_ , \new_[94053]_ , \new_[94054]_ ,
    \new_[94055]_ , \new_[94058]_ , \new_[94061]_ , \new_[94062]_ ,
    \new_[94065]_ , \new_[94068]_ , \new_[94069]_ , \new_[94070]_ ,
    \new_[94074]_ , \new_[94075]_ , \new_[94078]_ , \new_[94081]_ ,
    \new_[94082]_ , \new_[94083]_ , \new_[94086]_ , \new_[94089]_ ,
    \new_[94090]_ , \new_[94093]_ , \new_[94096]_ , \new_[94097]_ ,
    \new_[94098]_ , \new_[94102]_ , \new_[94103]_ , \new_[94106]_ ,
    \new_[94109]_ , \new_[94110]_ , \new_[94111]_ , \new_[94114]_ ,
    \new_[94117]_ , \new_[94118]_ , \new_[94121]_ , \new_[94124]_ ,
    \new_[94125]_ , \new_[94126]_ , \new_[94130]_ , \new_[94131]_ ,
    \new_[94134]_ , \new_[94137]_ , \new_[94138]_ , \new_[94139]_ ,
    \new_[94142]_ , \new_[94145]_ , \new_[94146]_ , \new_[94149]_ ,
    \new_[94152]_ , \new_[94153]_ , \new_[94154]_ , \new_[94158]_ ,
    \new_[94159]_ , \new_[94162]_ , \new_[94165]_ , \new_[94166]_ ,
    \new_[94167]_ , \new_[94170]_ , \new_[94173]_ , \new_[94174]_ ,
    \new_[94177]_ , \new_[94180]_ , \new_[94181]_ , \new_[94182]_ ,
    \new_[94186]_ , \new_[94187]_ , \new_[94190]_ , \new_[94193]_ ,
    \new_[94194]_ , \new_[94195]_ , \new_[94198]_ , \new_[94201]_ ,
    \new_[94202]_ , \new_[94205]_ , \new_[94208]_ , \new_[94209]_ ,
    \new_[94210]_ , \new_[94214]_ , \new_[94215]_ , \new_[94218]_ ,
    \new_[94221]_ , \new_[94222]_ , \new_[94223]_ , \new_[94226]_ ,
    \new_[94229]_ , \new_[94230]_ , \new_[94233]_ , \new_[94236]_ ,
    \new_[94237]_ , \new_[94238]_ , \new_[94242]_ , \new_[94243]_ ,
    \new_[94246]_ , \new_[94249]_ , \new_[94250]_ , \new_[94251]_ ,
    \new_[94254]_ , \new_[94257]_ , \new_[94258]_ , \new_[94261]_ ,
    \new_[94264]_ , \new_[94265]_ , \new_[94266]_ , \new_[94270]_ ,
    \new_[94271]_ , \new_[94274]_ , \new_[94277]_ , \new_[94278]_ ,
    \new_[94279]_ , \new_[94282]_ , \new_[94285]_ , \new_[94286]_ ,
    \new_[94289]_ , \new_[94292]_ , \new_[94293]_ , \new_[94294]_ ,
    \new_[94298]_ , \new_[94299]_ , \new_[94302]_ , \new_[94305]_ ,
    \new_[94306]_ , \new_[94307]_ , \new_[94310]_ , \new_[94313]_ ,
    \new_[94314]_ , \new_[94317]_ , \new_[94320]_ , \new_[94321]_ ,
    \new_[94322]_ , \new_[94326]_ , \new_[94327]_ , \new_[94330]_ ,
    \new_[94333]_ , \new_[94334]_ , \new_[94335]_ , \new_[94338]_ ,
    \new_[94341]_ , \new_[94342]_ , \new_[94345]_ , \new_[94348]_ ,
    \new_[94349]_ , \new_[94350]_ , \new_[94354]_ , \new_[94355]_ ,
    \new_[94358]_ , \new_[94361]_ , \new_[94362]_ , \new_[94363]_ ,
    \new_[94366]_ , \new_[94369]_ , \new_[94370]_ , \new_[94373]_ ,
    \new_[94376]_ , \new_[94377]_ , \new_[94378]_ , \new_[94382]_ ,
    \new_[94383]_ , \new_[94386]_ , \new_[94389]_ , \new_[94390]_ ,
    \new_[94391]_ , \new_[94394]_ , \new_[94397]_ , \new_[94398]_ ,
    \new_[94401]_ , \new_[94404]_ , \new_[94405]_ , \new_[94406]_ ,
    \new_[94410]_ , \new_[94411]_ , \new_[94414]_ , \new_[94417]_ ,
    \new_[94418]_ , \new_[94419]_ , \new_[94422]_ , \new_[94425]_ ,
    \new_[94426]_ , \new_[94429]_ , \new_[94432]_ , \new_[94433]_ ,
    \new_[94434]_ , \new_[94438]_ , \new_[94439]_ , \new_[94442]_ ,
    \new_[94445]_ , \new_[94446]_ , \new_[94447]_ , \new_[94450]_ ,
    \new_[94453]_ , \new_[94454]_ , \new_[94457]_ , \new_[94460]_ ,
    \new_[94461]_ , \new_[94462]_ , \new_[94466]_ , \new_[94467]_ ,
    \new_[94470]_ , \new_[94473]_ , \new_[94474]_ , \new_[94475]_ ,
    \new_[94478]_ , \new_[94481]_ , \new_[94482]_ , \new_[94485]_ ,
    \new_[94488]_ , \new_[94489]_ , \new_[94490]_ , \new_[94494]_ ,
    \new_[94495]_ , \new_[94498]_ , \new_[94501]_ , \new_[94502]_ ,
    \new_[94503]_ , \new_[94506]_ , \new_[94509]_ , \new_[94510]_ ,
    \new_[94513]_ , \new_[94516]_ , \new_[94517]_ , \new_[94518]_ ,
    \new_[94522]_ , \new_[94523]_ , \new_[94526]_ , \new_[94529]_ ,
    \new_[94530]_ , \new_[94531]_ , \new_[94534]_ , \new_[94537]_ ,
    \new_[94538]_ , \new_[94541]_ , \new_[94544]_ , \new_[94545]_ ,
    \new_[94546]_ , \new_[94550]_ , \new_[94551]_ , \new_[94554]_ ,
    \new_[94557]_ , \new_[94558]_ , \new_[94559]_ , \new_[94562]_ ,
    \new_[94565]_ , \new_[94566]_ , \new_[94569]_ , \new_[94572]_ ,
    \new_[94573]_ , \new_[94574]_ , \new_[94578]_ , \new_[94579]_ ,
    \new_[94582]_ , \new_[94585]_ , \new_[94586]_ , \new_[94587]_ ,
    \new_[94590]_ , \new_[94593]_ , \new_[94594]_ , \new_[94597]_ ,
    \new_[94600]_ , \new_[94601]_ , \new_[94602]_ , \new_[94606]_ ,
    \new_[94607]_ , \new_[94610]_ , \new_[94613]_ , \new_[94614]_ ,
    \new_[94615]_ , \new_[94618]_ , \new_[94621]_ , \new_[94622]_ ,
    \new_[94625]_ , \new_[94628]_ , \new_[94629]_ , \new_[94630]_ ,
    \new_[94634]_ , \new_[94635]_ , \new_[94638]_ , \new_[94641]_ ,
    \new_[94642]_ , \new_[94643]_ , \new_[94646]_ , \new_[94649]_ ,
    \new_[94650]_ , \new_[94653]_ , \new_[94656]_ , \new_[94657]_ ,
    \new_[94658]_ , \new_[94662]_ , \new_[94663]_ , \new_[94666]_ ,
    \new_[94669]_ , \new_[94670]_ , \new_[94671]_ , \new_[94674]_ ,
    \new_[94677]_ , \new_[94678]_ , \new_[94681]_ , \new_[94684]_ ,
    \new_[94685]_ , \new_[94686]_ , \new_[94690]_ , \new_[94691]_ ,
    \new_[94694]_ , \new_[94697]_ , \new_[94698]_ , \new_[94699]_ ,
    \new_[94702]_ , \new_[94705]_ , \new_[94706]_ , \new_[94709]_ ,
    \new_[94712]_ , \new_[94713]_ , \new_[94714]_ , \new_[94718]_ ,
    \new_[94719]_ , \new_[94722]_ , \new_[94725]_ , \new_[94726]_ ,
    \new_[94727]_ , \new_[94730]_ , \new_[94733]_ , \new_[94734]_ ,
    \new_[94737]_ , \new_[94740]_ , \new_[94741]_ , \new_[94742]_ ,
    \new_[94746]_ , \new_[94747]_ , \new_[94750]_ , \new_[94753]_ ,
    \new_[94754]_ , \new_[94755]_ , \new_[94758]_ , \new_[94761]_ ,
    \new_[94762]_ , \new_[94765]_ , \new_[94768]_ , \new_[94769]_ ,
    \new_[94770]_ , \new_[94774]_ , \new_[94775]_ , \new_[94778]_ ,
    \new_[94781]_ , \new_[94782]_ , \new_[94783]_ , \new_[94786]_ ,
    \new_[94789]_ , \new_[94790]_ , \new_[94793]_ , \new_[94796]_ ,
    \new_[94797]_ , \new_[94798]_ , \new_[94802]_ , \new_[94803]_ ,
    \new_[94806]_ , \new_[94809]_ , \new_[94810]_ , \new_[94811]_ ,
    \new_[94814]_ , \new_[94817]_ , \new_[94818]_ , \new_[94821]_ ,
    \new_[94824]_ , \new_[94825]_ , \new_[94826]_ , \new_[94830]_ ,
    \new_[94831]_ , \new_[94834]_ , \new_[94837]_ , \new_[94838]_ ,
    \new_[94839]_ , \new_[94842]_ , \new_[94845]_ , \new_[94846]_ ,
    \new_[94849]_ , \new_[94852]_ , \new_[94853]_ , \new_[94854]_ ,
    \new_[94858]_ , \new_[94859]_ , \new_[94862]_ , \new_[94865]_ ,
    \new_[94866]_ , \new_[94867]_ , \new_[94870]_ , \new_[94873]_ ,
    \new_[94874]_ , \new_[94877]_ , \new_[94880]_ , \new_[94881]_ ,
    \new_[94882]_ , \new_[94886]_ , \new_[94887]_ , \new_[94890]_ ,
    \new_[94893]_ , \new_[94894]_ , \new_[94895]_ , \new_[94898]_ ,
    \new_[94901]_ , \new_[94902]_ , \new_[94905]_ , \new_[94908]_ ,
    \new_[94909]_ , \new_[94910]_ , \new_[94914]_ , \new_[94915]_ ,
    \new_[94918]_ , \new_[94921]_ , \new_[94922]_ , \new_[94923]_ ,
    \new_[94926]_ , \new_[94929]_ , \new_[94930]_ , \new_[94933]_ ,
    \new_[94936]_ , \new_[94937]_ , \new_[94938]_ , \new_[94942]_ ,
    \new_[94943]_ , \new_[94946]_ , \new_[94949]_ , \new_[94950]_ ,
    \new_[94951]_ , \new_[94954]_ , \new_[94957]_ , \new_[94958]_ ,
    \new_[94961]_ , \new_[94964]_ , \new_[94965]_ , \new_[94966]_ ,
    \new_[94970]_ , \new_[94971]_ , \new_[94974]_ , \new_[94977]_ ,
    \new_[94978]_ , \new_[94979]_ , \new_[94982]_ , \new_[94985]_ ,
    \new_[94986]_ , \new_[94989]_ , \new_[94992]_ , \new_[94993]_ ,
    \new_[94994]_ , \new_[94998]_ , \new_[94999]_ , \new_[95002]_ ,
    \new_[95005]_ , \new_[95006]_ , \new_[95007]_ , \new_[95010]_ ,
    \new_[95013]_ , \new_[95014]_ , \new_[95017]_ , \new_[95020]_ ,
    \new_[95021]_ , \new_[95022]_ , \new_[95026]_ , \new_[95027]_ ,
    \new_[95030]_ , \new_[95033]_ , \new_[95034]_ , \new_[95035]_ ,
    \new_[95038]_ , \new_[95041]_ , \new_[95042]_ , \new_[95045]_ ,
    \new_[95048]_ , \new_[95049]_ , \new_[95050]_ , \new_[95054]_ ,
    \new_[95055]_ , \new_[95058]_ , \new_[95061]_ , \new_[95062]_ ,
    \new_[95063]_ , \new_[95066]_ , \new_[95069]_ , \new_[95070]_ ,
    \new_[95073]_ , \new_[95076]_ , \new_[95077]_ , \new_[95078]_ ,
    \new_[95082]_ , \new_[95083]_ , \new_[95086]_ , \new_[95089]_ ,
    \new_[95090]_ , \new_[95091]_ , \new_[95094]_ , \new_[95097]_ ,
    \new_[95098]_ , \new_[95101]_ , \new_[95104]_ , \new_[95105]_ ,
    \new_[95106]_ , \new_[95110]_ , \new_[95111]_ , \new_[95114]_ ,
    \new_[95117]_ , \new_[95118]_ , \new_[95119]_ , \new_[95122]_ ,
    \new_[95125]_ , \new_[95126]_ , \new_[95129]_ , \new_[95132]_ ,
    \new_[95133]_ , \new_[95134]_ , \new_[95138]_ , \new_[95139]_ ,
    \new_[95142]_ , \new_[95145]_ , \new_[95146]_ , \new_[95147]_ ,
    \new_[95150]_ , \new_[95153]_ , \new_[95154]_ , \new_[95157]_ ,
    \new_[95160]_ , \new_[95161]_ , \new_[95162]_ , \new_[95166]_ ,
    \new_[95167]_ , \new_[95170]_ , \new_[95173]_ , \new_[95174]_ ,
    \new_[95175]_ , \new_[95178]_ , \new_[95181]_ , \new_[95182]_ ,
    \new_[95185]_ , \new_[95188]_ , \new_[95189]_ , \new_[95190]_ ,
    \new_[95194]_ , \new_[95195]_ , \new_[95198]_ , \new_[95201]_ ,
    \new_[95202]_ , \new_[95203]_ , \new_[95206]_ , \new_[95209]_ ,
    \new_[95210]_ , \new_[95213]_ , \new_[95216]_ , \new_[95217]_ ,
    \new_[95218]_ , \new_[95222]_ , \new_[95223]_ , \new_[95226]_ ,
    \new_[95229]_ , \new_[95230]_ , \new_[95231]_ , \new_[95234]_ ,
    \new_[95237]_ , \new_[95238]_ , \new_[95241]_ , \new_[95244]_ ,
    \new_[95245]_ , \new_[95246]_ , \new_[95250]_ , \new_[95251]_ ,
    \new_[95254]_ , \new_[95257]_ , \new_[95258]_ , \new_[95259]_ ,
    \new_[95262]_ , \new_[95265]_ , \new_[95266]_ , \new_[95269]_ ,
    \new_[95272]_ , \new_[95273]_ , \new_[95274]_ , \new_[95278]_ ,
    \new_[95279]_ , \new_[95282]_ , \new_[95285]_ , \new_[95286]_ ,
    \new_[95287]_ , \new_[95290]_ , \new_[95293]_ , \new_[95294]_ ,
    \new_[95297]_ , \new_[95300]_ , \new_[95301]_ , \new_[95302]_ ,
    \new_[95306]_ , \new_[95307]_ , \new_[95310]_ , \new_[95313]_ ,
    \new_[95314]_ , \new_[95315]_ , \new_[95318]_ , \new_[95321]_ ,
    \new_[95322]_ , \new_[95325]_ , \new_[95328]_ , \new_[95329]_ ,
    \new_[95330]_ , \new_[95334]_ , \new_[95335]_ , \new_[95338]_ ,
    \new_[95341]_ , \new_[95342]_ , \new_[95343]_ , \new_[95346]_ ,
    \new_[95349]_ , \new_[95350]_ , \new_[95353]_ , \new_[95356]_ ,
    \new_[95357]_ , \new_[95358]_ , \new_[95362]_ , \new_[95363]_ ,
    \new_[95366]_ , \new_[95369]_ , \new_[95370]_ , \new_[95371]_ ,
    \new_[95374]_ , \new_[95377]_ , \new_[95378]_ , \new_[95381]_ ,
    \new_[95384]_ , \new_[95385]_ , \new_[95386]_ , \new_[95390]_ ,
    \new_[95391]_ , \new_[95394]_ , \new_[95397]_ , \new_[95398]_ ,
    \new_[95399]_ , \new_[95402]_ , \new_[95405]_ , \new_[95406]_ ,
    \new_[95409]_ , \new_[95412]_ , \new_[95413]_ , \new_[95414]_ ,
    \new_[95418]_ , \new_[95419]_ , \new_[95422]_ , \new_[95425]_ ,
    \new_[95426]_ , \new_[95427]_ , \new_[95430]_ , \new_[95433]_ ,
    \new_[95434]_ , \new_[95437]_ , \new_[95440]_ , \new_[95441]_ ,
    \new_[95442]_ , \new_[95446]_ , \new_[95447]_ , \new_[95450]_ ,
    \new_[95453]_ , \new_[95454]_ , \new_[95455]_ , \new_[95458]_ ,
    \new_[95461]_ , \new_[95462]_ , \new_[95465]_ , \new_[95468]_ ,
    \new_[95469]_ , \new_[95470]_ , \new_[95474]_ , \new_[95475]_ ,
    \new_[95478]_ , \new_[95481]_ , \new_[95482]_ , \new_[95483]_ ,
    \new_[95486]_ , \new_[95489]_ , \new_[95490]_ , \new_[95493]_ ,
    \new_[95496]_ , \new_[95497]_ , \new_[95498]_ , \new_[95502]_ ,
    \new_[95503]_ , \new_[95506]_ , \new_[95509]_ , \new_[95510]_ ,
    \new_[95511]_ , \new_[95514]_ , \new_[95517]_ , \new_[95518]_ ,
    \new_[95521]_ , \new_[95524]_ , \new_[95525]_ , \new_[95526]_ ,
    \new_[95530]_ , \new_[95531]_ , \new_[95534]_ , \new_[95537]_ ,
    \new_[95538]_ , \new_[95539]_ , \new_[95542]_ , \new_[95545]_ ,
    \new_[95546]_ , \new_[95549]_ , \new_[95552]_ , \new_[95553]_ ,
    \new_[95554]_ , \new_[95558]_ , \new_[95559]_ , \new_[95562]_ ,
    \new_[95565]_ , \new_[95566]_ , \new_[95567]_ , \new_[95570]_ ,
    \new_[95573]_ , \new_[95574]_ , \new_[95577]_ , \new_[95580]_ ,
    \new_[95581]_ , \new_[95582]_ , \new_[95586]_ , \new_[95587]_ ,
    \new_[95590]_ , \new_[95593]_ , \new_[95594]_ , \new_[95595]_ ,
    \new_[95598]_ , \new_[95601]_ , \new_[95602]_ , \new_[95605]_ ,
    \new_[95608]_ , \new_[95609]_ , \new_[95610]_ , \new_[95614]_ ,
    \new_[95615]_ , \new_[95618]_ , \new_[95621]_ , \new_[95622]_ ,
    \new_[95623]_ , \new_[95626]_ , \new_[95629]_ , \new_[95630]_ ,
    \new_[95633]_ , \new_[95636]_ , \new_[95637]_ , \new_[95638]_ ,
    \new_[95642]_ , \new_[95643]_ , \new_[95646]_ , \new_[95649]_ ,
    \new_[95650]_ , \new_[95651]_ , \new_[95654]_ , \new_[95657]_ ,
    \new_[95658]_ , \new_[95661]_ , \new_[95664]_ , \new_[95665]_ ,
    \new_[95666]_ , \new_[95670]_ , \new_[95671]_ , \new_[95674]_ ,
    \new_[95677]_ , \new_[95678]_ , \new_[95679]_ , \new_[95682]_ ,
    \new_[95685]_ , \new_[95686]_ , \new_[95689]_ , \new_[95692]_ ,
    \new_[95693]_ , \new_[95694]_ , \new_[95698]_ , \new_[95699]_ ,
    \new_[95702]_ , \new_[95705]_ , \new_[95706]_ , \new_[95707]_ ,
    \new_[95710]_ , \new_[95713]_ , \new_[95714]_ , \new_[95717]_ ,
    \new_[95720]_ , \new_[95721]_ , \new_[95722]_ , \new_[95726]_ ,
    \new_[95727]_ , \new_[95730]_ , \new_[95733]_ , \new_[95734]_ ,
    \new_[95735]_ , \new_[95738]_ , \new_[95741]_ , \new_[95742]_ ,
    \new_[95745]_ , \new_[95748]_ , \new_[95749]_ , \new_[95750]_ ,
    \new_[95754]_ , \new_[95755]_ , \new_[95758]_ , \new_[95761]_ ,
    \new_[95762]_ , \new_[95763]_ , \new_[95766]_ , \new_[95769]_ ,
    \new_[95770]_ , \new_[95773]_ , \new_[95776]_ , \new_[95777]_ ,
    \new_[95778]_ , \new_[95782]_ , \new_[95783]_ , \new_[95786]_ ,
    \new_[95789]_ , \new_[95790]_ , \new_[95791]_ , \new_[95794]_ ,
    \new_[95797]_ , \new_[95798]_ , \new_[95801]_ , \new_[95804]_ ,
    \new_[95805]_ , \new_[95806]_ , \new_[95810]_ , \new_[95811]_ ,
    \new_[95814]_ , \new_[95817]_ , \new_[95818]_ , \new_[95819]_ ,
    \new_[95822]_ , \new_[95825]_ , \new_[95826]_ , \new_[95829]_ ,
    \new_[95832]_ , \new_[95833]_ , \new_[95834]_ , \new_[95838]_ ,
    \new_[95839]_ , \new_[95842]_ , \new_[95845]_ , \new_[95846]_ ,
    \new_[95847]_ , \new_[95850]_ , \new_[95853]_ , \new_[95854]_ ,
    \new_[95857]_ , \new_[95860]_ , \new_[95861]_ , \new_[95862]_ ,
    \new_[95866]_ , \new_[95867]_ , \new_[95870]_ , \new_[95873]_ ,
    \new_[95874]_ , \new_[95875]_ , \new_[95878]_ , \new_[95881]_ ,
    \new_[95882]_ , \new_[95885]_ , \new_[95888]_ , \new_[95889]_ ,
    \new_[95890]_ , \new_[95894]_ , \new_[95895]_ , \new_[95898]_ ,
    \new_[95901]_ , \new_[95902]_ , \new_[95903]_ , \new_[95906]_ ,
    \new_[95909]_ , \new_[95910]_ , \new_[95913]_ , \new_[95916]_ ,
    \new_[95917]_ , \new_[95918]_ , \new_[95922]_ , \new_[95923]_ ,
    \new_[95926]_ , \new_[95929]_ , \new_[95930]_ , \new_[95931]_ ,
    \new_[95934]_ , \new_[95937]_ , \new_[95938]_ , \new_[95941]_ ,
    \new_[95944]_ , \new_[95945]_ , \new_[95946]_ , \new_[95950]_ ,
    \new_[95951]_ , \new_[95954]_ , \new_[95957]_ , \new_[95958]_ ,
    \new_[95959]_ , \new_[95962]_ , \new_[95965]_ , \new_[95966]_ ,
    \new_[95969]_ , \new_[95972]_ , \new_[95973]_ , \new_[95974]_ ,
    \new_[95978]_ , \new_[95979]_ , \new_[95982]_ , \new_[95985]_ ,
    \new_[95986]_ , \new_[95987]_ , \new_[95990]_ , \new_[95993]_ ,
    \new_[95994]_ , \new_[95997]_ , \new_[96000]_ , \new_[96001]_ ,
    \new_[96002]_ , \new_[96006]_ , \new_[96007]_ , \new_[96010]_ ,
    \new_[96013]_ , \new_[96014]_ , \new_[96015]_ , \new_[96018]_ ,
    \new_[96021]_ , \new_[96022]_ , \new_[96025]_ , \new_[96028]_ ,
    \new_[96029]_ , \new_[96030]_ , \new_[96034]_ , \new_[96035]_ ,
    \new_[96038]_ , \new_[96041]_ , \new_[96042]_ , \new_[96043]_ ,
    \new_[96046]_ , \new_[96049]_ , \new_[96050]_ , \new_[96053]_ ,
    \new_[96056]_ , \new_[96057]_ , \new_[96058]_ , \new_[96062]_ ,
    \new_[96063]_ , \new_[96066]_ , \new_[96069]_ , \new_[96070]_ ,
    \new_[96071]_ , \new_[96074]_ , \new_[96077]_ , \new_[96078]_ ,
    \new_[96081]_ , \new_[96084]_ , \new_[96085]_ , \new_[96086]_ ,
    \new_[96090]_ , \new_[96091]_ , \new_[96094]_ , \new_[96097]_ ,
    \new_[96098]_ , \new_[96099]_ , \new_[96102]_ , \new_[96105]_ ,
    \new_[96106]_ , \new_[96109]_ , \new_[96112]_ , \new_[96113]_ ,
    \new_[96114]_ , \new_[96118]_ , \new_[96119]_ , \new_[96122]_ ,
    \new_[96125]_ , \new_[96126]_ , \new_[96127]_ , \new_[96130]_ ,
    \new_[96133]_ , \new_[96134]_ , \new_[96137]_ , \new_[96140]_ ,
    \new_[96141]_ , \new_[96142]_ , \new_[96146]_ , \new_[96147]_ ,
    \new_[96150]_ , \new_[96153]_ , \new_[96154]_ , \new_[96155]_ ,
    \new_[96158]_ , \new_[96161]_ , \new_[96162]_ , \new_[96165]_ ,
    \new_[96168]_ , \new_[96169]_ , \new_[96170]_ , \new_[96174]_ ,
    \new_[96175]_ , \new_[96178]_ , \new_[96181]_ , \new_[96182]_ ,
    \new_[96183]_ , \new_[96186]_ , \new_[96189]_ , \new_[96190]_ ,
    \new_[96193]_ , \new_[96196]_ , \new_[96197]_ , \new_[96198]_ ,
    \new_[96202]_ , \new_[96203]_ , \new_[96206]_ , \new_[96209]_ ,
    \new_[96210]_ , \new_[96211]_ , \new_[96214]_ , \new_[96217]_ ,
    \new_[96218]_ , \new_[96221]_ , \new_[96224]_ , \new_[96225]_ ,
    \new_[96226]_ , \new_[96230]_ , \new_[96231]_ , \new_[96234]_ ,
    \new_[96237]_ , \new_[96238]_ , \new_[96239]_ , \new_[96242]_ ,
    \new_[96245]_ , \new_[96246]_ , \new_[96249]_ , \new_[96252]_ ,
    \new_[96253]_ , \new_[96254]_ , \new_[96258]_ , \new_[96259]_ ,
    \new_[96262]_ , \new_[96265]_ , \new_[96266]_ , \new_[96267]_ ,
    \new_[96270]_ , \new_[96273]_ , \new_[96274]_ , \new_[96277]_ ,
    \new_[96280]_ , \new_[96281]_ , \new_[96282]_ , \new_[96286]_ ,
    \new_[96287]_ , \new_[96290]_ , \new_[96293]_ , \new_[96294]_ ,
    \new_[96295]_ , \new_[96298]_ , \new_[96301]_ , \new_[96302]_ ,
    \new_[96305]_ , \new_[96308]_ , \new_[96309]_ , \new_[96310]_ ,
    \new_[96314]_ , \new_[96315]_ , \new_[96318]_ , \new_[96321]_ ,
    \new_[96322]_ , \new_[96323]_ , \new_[96326]_ , \new_[96329]_ ,
    \new_[96330]_ , \new_[96333]_ , \new_[96336]_ , \new_[96337]_ ,
    \new_[96338]_ , \new_[96342]_ , \new_[96343]_ , \new_[96346]_ ,
    \new_[96349]_ , \new_[96350]_ , \new_[96351]_ , \new_[96354]_ ,
    \new_[96357]_ , \new_[96358]_ , \new_[96361]_ , \new_[96364]_ ,
    \new_[96365]_ , \new_[96366]_ , \new_[96370]_ , \new_[96371]_ ,
    \new_[96374]_ , \new_[96377]_ , \new_[96378]_ , \new_[96379]_ ,
    \new_[96382]_ , \new_[96385]_ , \new_[96386]_ , \new_[96389]_ ,
    \new_[96392]_ , \new_[96393]_ , \new_[96394]_ , \new_[96398]_ ,
    \new_[96399]_ , \new_[96402]_ , \new_[96405]_ , \new_[96406]_ ,
    \new_[96407]_ , \new_[96410]_ , \new_[96413]_ , \new_[96414]_ ,
    \new_[96417]_ , \new_[96420]_ , \new_[96421]_ , \new_[96422]_ ,
    \new_[96426]_ , \new_[96427]_ , \new_[96430]_ , \new_[96433]_ ,
    \new_[96434]_ , \new_[96435]_ , \new_[96438]_ , \new_[96441]_ ,
    \new_[96442]_ , \new_[96445]_ , \new_[96448]_ , \new_[96449]_ ,
    \new_[96450]_ , \new_[96454]_ , \new_[96455]_ , \new_[96458]_ ,
    \new_[96461]_ , \new_[96462]_ , \new_[96463]_ , \new_[96466]_ ,
    \new_[96469]_ , \new_[96470]_ , \new_[96473]_ , \new_[96476]_ ,
    \new_[96477]_ , \new_[96478]_ , \new_[96482]_ , \new_[96483]_ ,
    \new_[96486]_ , \new_[96489]_ , \new_[96490]_ , \new_[96491]_ ,
    \new_[96494]_ , \new_[96497]_ , \new_[96498]_ , \new_[96501]_ ,
    \new_[96504]_ , \new_[96505]_ , \new_[96506]_ , \new_[96510]_ ,
    \new_[96511]_ , \new_[96514]_ , \new_[96517]_ , \new_[96518]_ ,
    \new_[96519]_ , \new_[96522]_ , \new_[96525]_ , \new_[96526]_ ,
    \new_[96529]_ , \new_[96532]_ , \new_[96533]_ , \new_[96534]_ ,
    \new_[96538]_ , \new_[96539]_ , \new_[96542]_ , \new_[96545]_ ,
    \new_[96546]_ , \new_[96547]_ , \new_[96550]_ , \new_[96553]_ ,
    \new_[96554]_ , \new_[96557]_ , \new_[96560]_ , \new_[96561]_ ,
    \new_[96562]_ , \new_[96566]_ , \new_[96567]_ , \new_[96570]_ ,
    \new_[96573]_ , \new_[96574]_ , \new_[96575]_ , \new_[96578]_ ,
    \new_[96581]_ , \new_[96582]_ , \new_[96585]_ , \new_[96588]_ ,
    \new_[96589]_ , \new_[96590]_ , \new_[96594]_ , \new_[96595]_ ,
    \new_[96598]_ , \new_[96601]_ , \new_[96602]_ , \new_[96603]_ ,
    \new_[96606]_ , \new_[96609]_ , \new_[96610]_ , \new_[96613]_ ,
    \new_[96616]_ , \new_[96617]_ , \new_[96618]_ , \new_[96622]_ ,
    \new_[96623]_ , \new_[96626]_ , \new_[96629]_ , \new_[96630]_ ,
    \new_[96631]_ , \new_[96634]_ , \new_[96637]_ , \new_[96638]_ ,
    \new_[96641]_ , \new_[96644]_ , \new_[96645]_ , \new_[96646]_ ,
    \new_[96650]_ , \new_[96651]_ , \new_[96654]_ , \new_[96657]_ ,
    \new_[96658]_ , \new_[96659]_ , \new_[96662]_ , \new_[96665]_ ,
    \new_[96666]_ , \new_[96669]_ , \new_[96672]_ , \new_[96673]_ ,
    \new_[96674]_ , \new_[96678]_ , \new_[96679]_ , \new_[96682]_ ,
    \new_[96685]_ , \new_[96686]_ , \new_[96687]_ , \new_[96690]_ ,
    \new_[96693]_ , \new_[96694]_ , \new_[96697]_ , \new_[96700]_ ,
    \new_[96701]_ , \new_[96702]_ , \new_[96706]_ , \new_[96707]_ ,
    \new_[96710]_ , \new_[96713]_ , \new_[96714]_ , \new_[96715]_ ,
    \new_[96718]_ , \new_[96721]_ , \new_[96722]_ , \new_[96725]_ ,
    \new_[96728]_ , \new_[96729]_ , \new_[96730]_ , \new_[96734]_ ,
    \new_[96735]_ , \new_[96738]_ , \new_[96741]_ , \new_[96742]_ ,
    \new_[96743]_ , \new_[96746]_ , \new_[96749]_ , \new_[96750]_ ,
    \new_[96753]_ , \new_[96756]_ , \new_[96757]_ , \new_[96758]_ ,
    \new_[96762]_ , \new_[96763]_ , \new_[96766]_ , \new_[96769]_ ,
    \new_[96770]_ , \new_[96771]_ , \new_[96774]_ , \new_[96777]_ ,
    \new_[96778]_ , \new_[96781]_ , \new_[96784]_ , \new_[96785]_ ,
    \new_[96786]_ , \new_[96790]_ , \new_[96791]_ , \new_[96794]_ ,
    \new_[96797]_ , \new_[96798]_ , \new_[96799]_ , \new_[96802]_ ,
    \new_[96805]_ , \new_[96806]_ , \new_[96809]_ , \new_[96812]_ ,
    \new_[96813]_ , \new_[96814]_ , \new_[96818]_ , \new_[96819]_ ,
    \new_[96822]_ , \new_[96825]_ , \new_[96826]_ , \new_[96827]_ ,
    \new_[96830]_ , \new_[96833]_ , \new_[96834]_ , \new_[96837]_ ,
    \new_[96840]_ , \new_[96841]_ , \new_[96842]_ , \new_[96846]_ ,
    \new_[96847]_ , \new_[96850]_ , \new_[96853]_ , \new_[96854]_ ,
    \new_[96855]_ , \new_[96858]_ , \new_[96861]_ , \new_[96862]_ ,
    \new_[96865]_ , \new_[96868]_ , \new_[96869]_ , \new_[96870]_ ,
    \new_[96874]_ , \new_[96875]_ , \new_[96878]_ , \new_[96881]_ ,
    \new_[96882]_ , \new_[96883]_ , \new_[96886]_ , \new_[96889]_ ,
    \new_[96890]_ , \new_[96893]_ , \new_[96896]_ , \new_[96897]_ ,
    \new_[96898]_ , \new_[96902]_ , \new_[96903]_ , \new_[96906]_ ,
    \new_[96909]_ , \new_[96910]_ , \new_[96911]_ , \new_[96914]_ ,
    \new_[96917]_ , \new_[96918]_ , \new_[96921]_ , \new_[96924]_ ,
    \new_[96925]_ , \new_[96926]_ , \new_[96930]_ , \new_[96931]_ ,
    \new_[96934]_ , \new_[96937]_ , \new_[96938]_ , \new_[96939]_ ,
    \new_[96942]_ , \new_[96945]_ , \new_[96946]_ , \new_[96949]_ ,
    \new_[96952]_ , \new_[96953]_ , \new_[96954]_ , \new_[96958]_ ,
    \new_[96959]_ , \new_[96962]_ , \new_[96965]_ , \new_[96966]_ ,
    \new_[96967]_ , \new_[96970]_ , \new_[96973]_ , \new_[96974]_ ,
    \new_[96977]_ , \new_[96980]_ , \new_[96981]_ , \new_[96982]_ ,
    \new_[96986]_ , \new_[96987]_ , \new_[96990]_ , \new_[96993]_ ,
    \new_[96994]_ , \new_[96995]_ , \new_[96998]_ , \new_[97001]_ ,
    \new_[97002]_ , \new_[97005]_ , \new_[97008]_ , \new_[97009]_ ,
    \new_[97010]_ , \new_[97014]_ , \new_[97015]_ , \new_[97018]_ ,
    \new_[97021]_ , \new_[97022]_ , \new_[97023]_ , \new_[97026]_ ,
    \new_[97029]_ , \new_[97030]_ , \new_[97033]_ , \new_[97036]_ ,
    \new_[97037]_ , \new_[97038]_ , \new_[97042]_ , \new_[97043]_ ,
    \new_[97046]_ , \new_[97049]_ , \new_[97050]_ , \new_[97051]_ ,
    \new_[97054]_ , \new_[97057]_ , \new_[97058]_ , \new_[97061]_ ,
    \new_[97064]_ , \new_[97065]_ , \new_[97066]_ , \new_[97070]_ ,
    \new_[97071]_ , \new_[97074]_ , \new_[97077]_ , \new_[97078]_ ,
    \new_[97079]_ , \new_[97082]_ , \new_[97085]_ , \new_[97086]_ ,
    \new_[97089]_ , \new_[97092]_ , \new_[97093]_ , \new_[97094]_ ,
    \new_[97098]_ , \new_[97099]_ , \new_[97102]_ , \new_[97105]_ ,
    \new_[97106]_ , \new_[97107]_ , \new_[97110]_ , \new_[97113]_ ,
    \new_[97114]_ , \new_[97117]_ , \new_[97120]_ , \new_[97121]_ ,
    \new_[97122]_ , \new_[97126]_ , \new_[97127]_ , \new_[97130]_ ,
    \new_[97133]_ , \new_[97134]_ , \new_[97135]_ , \new_[97138]_ ,
    \new_[97141]_ , \new_[97142]_ , \new_[97145]_ , \new_[97148]_ ,
    \new_[97149]_ , \new_[97150]_ , \new_[97154]_ , \new_[97155]_ ,
    \new_[97158]_ , \new_[97161]_ , \new_[97162]_ , \new_[97163]_ ,
    \new_[97166]_ , \new_[97169]_ , \new_[97170]_ , \new_[97173]_ ,
    \new_[97176]_ , \new_[97177]_ , \new_[97178]_ , \new_[97182]_ ,
    \new_[97183]_ , \new_[97186]_ , \new_[97189]_ , \new_[97190]_ ,
    \new_[97191]_ , \new_[97194]_ , \new_[97197]_ , \new_[97198]_ ,
    \new_[97201]_ , \new_[97204]_ , \new_[97205]_ , \new_[97206]_ ,
    \new_[97210]_ , \new_[97211]_ , \new_[97214]_ , \new_[97217]_ ,
    \new_[97218]_ , \new_[97219]_ , \new_[97222]_ , \new_[97225]_ ,
    \new_[97226]_ , \new_[97229]_ , \new_[97232]_ , \new_[97233]_ ,
    \new_[97234]_ , \new_[97238]_ , \new_[97239]_ , \new_[97242]_ ,
    \new_[97245]_ , \new_[97246]_ , \new_[97247]_ , \new_[97250]_ ,
    \new_[97253]_ , \new_[97254]_ , \new_[97257]_ , \new_[97260]_ ,
    \new_[97261]_ , \new_[97262]_ , \new_[97266]_ , \new_[97267]_ ,
    \new_[97270]_ , \new_[97273]_ , \new_[97274]_ , \new_[97275]_ ,
    \new_[97278]_ , \new_[97281]_ , \new_[97282]_ , \new_[97285]_ ,
    \new_[97288]_ , \new_[97289]_ , \new_[97290]_ , \new_[97294]_ ,
    \new_[97295]_ , \new_[97298]_ , \new_[97301]_ , \new_[97302]_ ,
    \new_[97303]_ , \new_[97306]_ , \new_[97309]_ , \new_[97310]_ ,
    \new_[97313]_ , \new_[97316]_ , \new_[97317]_ , \new_[97318]_ ,
    \new_[97322]_ , \new_[97323]_ , \new_[97326]_ , \new_[97329]_ ,
    \new_[97330]_ , \new_[97331]_ , \new_[97334]_ , \new_[97337]_ ,
    \new_[97338]_ , \new_[97341]_ , \new_[97344]_ , \new_[97345]_ ,
    \new_[97346]_ , \new_[97350]_ , \new_[97351]_ , \new_[97354]_ ,
    \new_[97357]_ , \new_[97358]_ , \new_[97359]_ , \new_[97362]_ ,
    \new_[97365]_ , \new_[97366]_ , \new_[97369]_ , \new_[97372]_ ,
    \new_[97373]_ , \new_[97374]_ , \new_[97378]_ , \new_[97379]_ ,
    \new_[97382]_ , \new_[97385]_ , \new_[97386]_ , \new_[97387]_ ,
    \new_[97390]_ , \new_[97393]_ , \new_[97394]_ , \new_[97397]_ ,
    \new_[97400]_ , \new_[97401]_ , \new_[97402]_ , \new_[97406]_ ,
    \new_[97407]_ , \new_[97410]_ , \new_[97413]_ , \new_[97414]_ ,
    \new_[97415]_ , \new_[97418]_ , \new_[97421]_ , \new_[97422]_ ,
    \new_[97425]_ , \new_[97428]_ , \new_[97429]_ , \new_[97430]_ ,
    \new_[97434]_ , \new_[97435]_ , \new_[97438]_ , \new_[97441]_ ,
    \new_[97442]_ , \new_[97443]_ , \new_[97446]_ , \new_[97449]_ ,
    \new_[97450]_ , \new_[97453]_ , \new_[97456]_ , \new_[97457]_ ,
    \new_[97458]_ , \new_[97462]_ , \new_[97463]_ , \new_[97466]_ ,
    \new_[97469]_ , \new_[97470]_ , \new_[97471]_ , \new_[97474]_ ,
    \new_[97477]_ , \new_[97478]_ , \new_[97481]_ , \new_[97484]_ ,
    \new_[97485]_ , \new_[97486]_ , \new_[97490]_ , \new_[97491]_ ,
    \new_[97494]_ , \new_[97497]_ , \new_[97498]_ , \new_[97499]_ ,
    \new_[97502]_ , \new_[97505]_ , \new_[97506]_ , \new_[97509]_ ,
    \new_[97512]_ , \new_[97513]_ , \new_[97514]_ , \new_[97518]_ ,
    \new_[97519]_ , \new_[97522]_ , \new_[97525]_ , \new_[97526]_ ,
    \new_[97527]_ , \new_[97530]_ , \new_[97533]_ , \new_[97534]_ ,
    \new_[97537]_ , \new_[97540]_ , \new_[97541]_ , \new_[97542]_ ,
    \new_[97545]_ , \new_[97548]_ , \new_[97549]_ , \new_[97552]_ ,
    \new_[97555]_ , \new_[97556]_ , \new_[97557]_ , \new_[97560]_ ,
    \new_[97563]_ , \new_[97564]_ , \new_[97567]_ , \new_[97570]_ ,
    \new_[97571]_ , \new_[97572]_ , \new_[97575]_ , \new_[97578]_ ,
    \new_[97579]_ , \new_[97582]_ , \new_[97585]_ , \new_[97586]_ ,
    \new_[97587]_ , \new_[97590]_ , \new_[97593]_ , \new_[97594]_ ,
    \new_[97597]_ , \new_[97600]_ , \new_[97601]_ , \new_[97602]_ ,
    \new_[97605]_ , \new_[97608]_ , \new_[97609]_ , \new_[97612]_ ,
    \new_[97615]_ , \new_[97616]_ , \new_[97617]_ , \new_[97620]_ ,
    \new_[97623]_ , \new_[97624]_ , \new_[97627]_ , \new_[97630]_ ,
    \new_[97631]_ , \new_[97632]_ , \new_[97635]_ , \new_[97638]_ ,
    \new_[97639]_ , \new_[97642]_ , \new_[97645]_ , \new_[97646]_ ,
    \new_[97647]_ , \new_[97650]_ , \new_[97653]_ , \new_[97654]_ ,
    \new_[97657]_ , \new_[97660]_ , \new_[97661]_ , \new_[97662]_ ,
    \new_[97665]_ , \new_[97668]_ , \new_[97669]_ , \new_[97672]_ ,
    \new_[97675]_ , \new_[97676]_ , \new_[97677]_ , \new_[97680]_ ,
    \new_[97683]_ , \new_[97684]_ , \new_[97687]_ , \new_[97690]_ ,
    \new_[97691]_ , \new_[97692]_ , \new_[97695]_ , \new_[97698]_ ,
    \new_[97699]_ , \new_[97702]_ , \new_[97705]_ , \new_[97706]_ ,
    \new_[97707]_ , \new_[97710]_ , \new_[97713]_ , \new_[97714]_ ,
    \new_[97717]_ , \new_[97720]_ , \new_[97721]_ , \new_[97722]_ ,
    \new_[97725]_ , \new_[97728]_ , \new_[97729]_ , \new_[97732]_ ,
    \new_[97735]_ , \new_[97736]_ , \new_[97737]_ , \new_[97740]_ ,
    \new_[97743]_ , \new_[97744]_ , \new_[97747]_ , \new_[97750]_ ,
    \new_[97751]_ , \new_[97752]_ , \new_[97755]_ , \new_[97758]_ ,
    \new_[97759]_ , \new_[97762]_ , \new_[97765]_ , \new_[97766]_ ,
    \new_[97767]_ , \new_[97770]_ , \new_[97773]_ , \new_[97774]_ ,
    \new_[97777]_ , \new_[97780]_ , \new_[97781]_ , \new_[97782]_ ,
    \new_[97785]_ , \new_[97788]_ , \new_[97789]_ , \new_[97792]_ ,
    \new_[97795]_ , \new_[97796]_ , \new_[97797]_ , \new_[97800]_ ,
    \new_[97803]_ , \new_[97804]_ , \new_[97807]_ , \new_[97810]_ ,
    \new_[97811]_ , \new_[97812]_ , \new_[97815]_ , \new_[97818]_ ,
    \new_[97819]_ , \new_[97822]_ , \new_[97825]_ , \new_[97826]_ ,
    \new_[97827]_ , \new_[97830]_ , \new_[97833]_ , \new_[97834]_ ,
    \new_[97837]_ , \new_[97840]_ , \new_[97841]_ , \new_[97842]_ ,
    \new_[97845]_ , \new_[97848]_ , \new_[97849]_ , \new_[97852]_ ,
    \new_[97855]_ , \new_[97856]_ , \new_[97857]_ , \new_[97860]_ ,
    \new_[97863]_ , \new_[97864]_ , \new_[97867]_ , \new_[97870]_ ,
    \new_[97871]_ , \new_[97872]_ , \new_[97875]_ , \new_[97878]_ ,
    \new_[97879]_ , \new_[97882]_ , \new_[97885]_ , \new_[97886]_ ,
    \new_[97887]_ , \new_[97890]_ , \new_[97893]_ , \new_[97894]_ ,
    \new_[97897]_ , \new_[97900]_ , \new_[97901]_ , \new_[97902]_ ,
    \new_[97905]_ , \new_[97908]_ , \new_[97909]_ , \new_[97912]_ ,
    \new_[97915]_ , \new_[97916]_ , \new_[97917]_ , \new_[97920]_ ,
    \new_[97923]_ , \new_[97924]_ , \new_[97927]_ , \new_[97930]_ ,
    \new_[97931]_ , \new_[97932]_ , \new_[97935]_ , \new_[97938]_ ,
    \new_[97939]_ , \new_[97942]_ , \new_[97945]_ , \new_[97946]_ ,
    \new_[97947]_ , \new_[97950]_ , \new_[97953]_ , \new_[97954]_ ,
    \new_[97957]_ , \new_[97960]_ , \new_[97961]_ , \new_[97962]_ ,
    \new_[97965]_ , \new_[97968]_ , \new_[97969]_ , \new_[97972]_ ,
    \new_[97975]_ , \new_[97976]_ , \new_[97977]_ , \new_[97980]_ ,
    \new_[97983]_ , \new_[97984]_ , \new_[97987]_ , \new_[97990]_ ,
    \new_[97991]_ , \new_[97992]_ , \new_[97995]_ , \new_[97998]_ ,
    \new_[97999]_ , \new_[98002]_ , \new_[98005]_ , \new_[98006]_ ,
    \new_[98007]_ , \new_[98010]_ , \new_[98013]_ , \new_[98014]_ ,
    \new_[98017]_ , \new_[98020]_ , \new_[98021]_ , \new_[98022]_ ,
    \new_[98025]_ , \new_[98028]_ , \new_[98029]_ , \new_[98032]_ ,
    \new_[98035]_ , \new_[98036]_ , \new_[98037]_ , \new_[98040]_ ,
    \new_[98043]_ , \new_[98044]_ , \new_[98047]_ , \new_[98050]_ ,
    \new_[98051]_ , \new_[98052]_ , \new_[98055]_ , \new_[98058]_ ,
    \new_[98059]_ , \new_[98062]_ , \new_[98065]_ , \new_[98066]_ ,
    \new_[98067]_ , \new_[98070]_ , \new_[98073]_ , \new_[98074]_ ,
    \new_[98077]_ , \new_[98080]_ , \new_[98081]_ , \new_[98082]_ ,
    \new_[98085]_ , \new_[98088]_ , \new_[98089]_ , \new_[98092]_ ,
    \new_[98095]_ , \new_[98096]_ , \new_[98097]_ , \new_[98100]_ ,
    \new_[98103]_ , \new_[98104]_ , \new_[98107]_ , \new_[98110]_ ,
    \new_[98111]_ , \new_[98112]_ , \new_[98115]_ , \new_[98118]_ ,
    \new_[98119]_ , \new_[98122]_ , \new_[98125]_ , \new_[98126]_ ,
    \new_[98127]_ , \new_[98130]_ , \new_[98133]_ , \new_[98134]_ ,
    \new_[98137]_ , \new_[98140]_ , \new_[98141]_ , \new_[98142]_ ,
    \new_[98145]_ , \new_[98148]_ , \new_[98149]_ , \new_[98152]_ ,
    \new_[98155]_ , \new_[98156]_ , \new_[98157]_ , \new_[98160]_ ,
    \new_[98163]_ , \new_[98164]_ , \new_[98167]_ , \new_[98170]_ ,
    \new_[98171]_ , \new_[98172]_ , \new_[98175]_ , \new_[98178]_ ,
    \new_[98179]_ , \new_[98182]_ , \new_[98185]_ , \new_[98186]_ ,
    \new_[98187]_ , \new_[98190]_ , \new_[98193]_ , \new_[98194]_ ,
    \new_[98197]_ , \new_[98200]_ , \new_[98201]_ , \new_[98202]_ ,
    \new_[98205]_ , \new_[98208]_ , \new_[98209]_ , \new_[98212]_ ,
    \new_[98215]_ , \new_[98216]_ , \new_[98217]_ , \new_[98220]_ ,
    \new_[98223]_ , \new_[98224]_ , \new_[98227]_ , \new_[98230]_ ,
    \new_[98231]_ , \new_[98232]_ , \new_[98235]_ , \new_[98238]_ ,
    \new_[98239]_ , \new_[98242]_ , \new_[98245]_ , \new_[98246]_ ,
    \new_[98247]_ , \new_[98250]_ , \new_[98253]_ , \new_[98254]_ ,
    \new_[98257]_ , \new_[98260]_ , \new_[98261]_ , \new_[98262]_ ,
    \new_[98265]_ , \new_[98268]_ , \new_[98269]_ , \new_[98272]_ ,
    \new_[98275]_ , \new_[98276]_ , \new_[98277]_ , \new_[98280]_ ,
    \new_[98283]_ , \new_[98284]_ , \new_[98287]_ , \new_[98290]_ ,
    \new_[98291]_ , \new_[98292]_ , \new_[98295]_ , \new_[98298]_ ,
    \new_[98299]_ , \new_[98302]_ , \new_[98305]_ , \new_[98306]_ ,
    \new_[98307]_ , \new_[98310]_ , \new_[98313]_ , \new_[98314]_ ,
    \new_[98317]_ , \new_[98320]_ , \new_[98321]_ , \new_[98322]_ ,
    \new_[98325]_ , \new_[98328]_ , \new_[98329]_ , \new_[98332]_ ,
    \new_[98335]_ , \new_[98336]_ , \new_[98337]_ , \new_[98340]_ ,
    \new_[98343]_ , \new_[98344]_ , \new_[98347]_ , \new_[98350]_ ,
    \new_[98351]_ , \new_[98352]_ , \new_[98355]_ , \new_[98358]_ ,
    \new_[98359]_ , \new_[98362]_ , \new_[98365]_ , \new_[98366]_ ,
    \new_[98367]_ , \new_[98370]_ , \new_[98373]_ , \new_[98374]_ ,
    \new_[98377]_ , \new_[98380]_ , \new_[98381]_ , \new_[98382]_ ,
    \new_[98385]_ , \new_[98388]_ , \new_[98389]_ , \new_[98392]_ ,
    \new_[98395]_ , \new_[98396]_ , \new_[98397]_ , \new_[98400]_ ,
    \new_[98403]_ , \new_[98404]_ , \new_[98407]_ , \new_[98410]_ ,
    \new_[98411]_ , \new_[98412]_ , \new_[98415]_ , \new_[98418]_ ,
    \new_[98419]_ , \new_[98422]_ , \new_[98425]_ , \new_[98426]_ ,
    \new_[98427]_ , \new_[98430]_ , \new_[98433]_ , \new_[98434]_ ,
    \new_[98437]_ , \new_[98440]_ , \new_[98441]_ , \new_[98442]_ ,
    \new_[98445]_ , \new_[98448]_ , \new_[98449]_ , \new_[98452]_ ,
    \new_[98455]_ , \new_[98456]_ , \new_[98457]_ , \new_[98460]_ ,
    \new_[98463]_ , \new_[98464]_ , \new_[98467]_ , \new_[98470]_ ,
    \new_[98471]_ , \new_[98472]_ , \new_[98475]_ , \new_[98478]_ ,
    \new_[98479]_ , \new_[98482]_ , \new_[98485]_ , \new_[98486]_ ,
    \new_[98487]_ , \new_[98490]_ , \new_[98493]_ , \new_[98494]_ ,
    \new_[98497]_ , \new_[98500]_ , \new_[98501]_ , \new_[98502]_ ,
    \new_[98505]_ , \new_[98508]_ , \new_[98509]_ , \new_[98512]_ ,
    \new_[98515]_ , \new_[98516]_ , \new_[98517]_ , \new_[98520]_ ,
    \new_[98523]_ , \new_[98524]_ , \new_[98527]_ , \new_[98530]_ ,
    \new_[98531]_ , \new_[98532]_ , \new_[98535]_ , \new_[98538]_ ,
    \new_[98539]_ , \new_[98542]_ , \new_[98545]_ , \new_[98546]_ ,
    \new_[98547]_ , \new_[98550]_ , \new_[98553]_ , \new_[98554]_ ,
    \new_[98557]_ , \new_[98560]_ , \new_[98561]_ , \new_[98562]_ ,
    \new_[98565]_ , \new_[98568]_ , \new_[98569]_ , \new_[98572]_ ,
    \new_[98575]_ , \new_[98576]_ , \new_[98577]_ , \new_[98580]_ ,
    \new_[98583]_ , \new_[98584]_ , \new_[98587]_ , \new_[98590]_ ,
    \new_[98591]_ , \new_[98592]_ , \new_[98595]_ , \new_[98598]_ ,
    \new_[98599]_ , \new_[98602]_ , \new_[98605]_ , \new_[98606]_ ,
    \new_[98607]_ , \new_[98610]_ , \new_[98613]_ , \new_[98614]_ ,
    \new_[98617]_ , \new_[98620]_ , \new_[98621]_ , \new_[98622]_ ,
    \new_[98625]_ , \new_[98628]_ , \new_[98629]_ , \new_[98632]_ ,
    \new_[98635]_ , \new_[98636]_ , \new_[98637]_ , \new_[98640]_ ,
    \new_[98643]_ , \new_[98644]_ , \new_[98647]_ , \new_[98650]_ ,
    \new_[98651]_ , \new_[98652]_ , \new_[98655]_ , \new_[98658]_ ,
    \new_[98659]_ , \new_[98662]_ , \new_[98665]_ , \new_[98666]_ ,
    \new_[98667]_ , \new_[98670]_ , \new_[98673]_ , \new_[98674]_ ,
    \new_[98677]_ , \new_[98680]_ , \new_[98681]_ , \new_[98682]_ ,
    \new_[98685]_ , \new_[98688]_ , \new_[98689]_ , \new_[98692]_ ,
    \new_[98695]_ , \new_[98696]_ , \new_[98697]_ , \new_[98700]_ ,
    \new_[98703]_ , \new_[98704]_ , \new_[98707]_ , \new_[98710]_ ,
    \new_[98711]_ , \new_[98712]_ , \new_[98715]_ , \new_[98718]_ ,
    \new_[98719]_ , \new_[98722]_ , \new_[98725]_ , \new_[98726]_ ,
    \new_[98727]_ , \new_[98730]_ , \new_[98733]_ , \new_[98734]_ ,
    \new_[98737]_ , \new_[98740]_ , \new_[98741]_ , \new_[98742]_ ,
    \new_[98745]_ , \new_[98748]_ , \new_[98749]_ , \new_[98752]_ ,
    \new_[98755]_ , \new_[98756]_ , \new_[98757]_ , \new_[98760]_ ,
    \new_[98763]_ , \new_[98764]_ , \new_[98767]_ , \new_[98770]_ ,
    \new_[98771]_ , \new_[98772]_ , \new_[98775]_ , \new_[98778]_ ,
    \new_[98779]_ , \new_[98782]_ , \new_[98785]_ , \new_[98786]_ ,
    \new_[98787]_ , \new_[98790]_ , \new_[98793]_ , \new_[98794]_ ,
    \new_[98797]_ , \new_[98800]_ , \new_[98801]_ , \new_[98802]_ ,
    \new_[98805]_ , \new_[98808]_ , \new_[98809]_ , \new_[98812]_ ,
    \new_[98815]_ , \new_[98816]_ , \new_[98817]_ , \new_[98820]_ ,
    \new_[98823]_ , \new_[98824]_ , \new_[98827]_ , \new_[98830]_ ,
    \new_[98831]_ , \new_[98832]_ , \new_[98835]_ , \new_[98838]_ ,
    \new_[98839]_ , \new_[98842]_ , \new_[98845]_ , \new_[98846]_ ,
    \new_[98847]_ , \new_[98850]_ , \new_[98853]_ , \new_[98854]_ ,
    \new_[98857]_ , \new_[98860]_ , \new_[98861]_ , \new_[98862]_ ,
    \new_[98865]_ , \new_[98868]_ , \new_[98869]_ , \new_[98872]_ ,
    \new_[98875]_ , \new_[98876]_ , \new_[98877]_ , \new_[98880]_ ,
    \new_[98883]_ , \new_[98884]_ , \new_[98887]_ , \new_[98890]_ ,
    \new_[98891]_ , \new_[98892]_ , \new_[98895]_ , \new_[98898]_ ,
    \new_[98899]_ , \new_[98902]_ , \new_[98905]_ , \new_[98906]_ ,
    \new_[98907]_ , \new_[98910]_ , \new_[98913]_ , \new_[98914]_ ,
    \new_[98917]_ , \new_[98920]_ , \new_[98921]_ , \new_[98922]_ ,
    \new_[98925]_ , \new_[98928]_ , \new_[98929]_ , \new_[98932]_ ,
    \new_[98935]_ , \new_[98936]_ , \new_[98937]_ , \new_[98940]_ ,
    \new_[98943]_ , \new_[98944]_ , \new_[98947]_ , \new_[98950]_ ,
    \new_[98951]_ , \new_[98952]_ , \new_[98955]_ , \new_[98958]_ ,
    \new_[98959]_ , \new_[98962]_ , \new_[98965]_ , \new_[98966]_ ,
    \new_[98967]_ , \new_[98970]_ , \new_[98973]_ , \new_[98974]_ ,
    \new_[98977]_ , \new_[98980]_ , \new_[98981]_ , \new_[98982]_ ,
    \new_[98985]_ , \new_[98988]_ , \new_[98989]_ , \new_[98992]_ ,
    \new_[98995]_ , \new_[98996]_ , \new_[98997]_ , \new_[99000]_ ,
    \new_[99003]_ , \new_[99004]_ , \new_[99007]_ , \new_[99010]_ ,
    \new_[99011]_ , \new_[99012]_ , \new_[99015]_ , \new_[99018]_ ,
    \new_[99019]_ , \new_[99022]_ , \new_[99025]_ , \new_[99026]_ ,
    \new_[99027]_ , \new_[99030]_ , \new_[99033]_ , \new_[99034]_ ,
    \new_[99037]_ , \new_[99040]_ , \new_[99041]_ , \new_[99042]_ ,
    \new_[99045]_ , \new_[99048]_ , \new_[99049]_ , \new_[99052]_ ,
    \new_[99055]_ , \new_[99056]_ , \new_[99057]_ , \new_[99060]_ ,
    \new_[99063]_ , \new_[99064]_ , \new_[99067]_ , \new_[99070]_ ,
    \new_[99071]_ , \new_[99072]_ , \new_[99075]_ , \new_[99078]_ ,
    \new_[99079]_ , \new_[99082]_ , \new_[99085]_ , \new_[99086]_ ,
    \new_[99087]_ , \new_[99090]_ , \new_[99093]_ , \new_[99094]_ ,
    \new_[99097]_ , \new_[99100]_ , \new_[99101]_ , \new_[99102]_ ,
    \new_[99105]_ , \new_[99108]_ , \new_[99109]_ , \new_[99112]_ ,
    \new_[99115]_ , \new_[99116]_ , \new_[99117]_ , \new_[99120]_ ,
    \new_[99123]_ , \new_[99124]_ , \new_[99127]_ , \new_[99130]_ ,
    \new_[99131]_ , \new_[99132]_ , \new_[99135]_ , \new_[99138]_ ,
    \new_[99139]_ , \new_[99142]_ , \new_[99145]_ , \new_[99146]_ ,
    \new_[99147]_ , \new_[99150]_ , \new_[99153]_ , \new_[99154]_ ,
    \new_[99157]_ , \new_[99160]_ , \new_[99161]_ , \new_[99162]_ ,
    \new_[99165]_ , \new_[99168]_ , \new_[99169]_ , \new_[99172]_ ,
    \new_[99175]_ , \new_[99176]_ , \new_[99177]_ , \new_[99180]_ ,
    \new_[99183]_ , \new_[99184]_ , \new_[99187]_ , \new_[99190]_ ,
    \new_[99191]_ , \new_[99192]_ , \new_[99195]_ , \new_[99198]_ ,
    \new_[99199]_ , \new_[99202]_ , \new_[99205]_ , \new_[99206]_ ,
    \new_[99207]_ , \new_[99210]_ , \new_[99213]_ , \new_[99214]_ ,
    \new_[99217]_ , \new_[99220]_ , \new_[99221]_ , \new_[99222]_ ,
    \new_[99225]_ , \new_[99228]_ , \new_[99229]_ , \new_[99232]_ ,
    \new_[99235]_ , \new_[99236]_ , \new_[99237]_ , \new_[99240]_ ,
    \new_[99243]_ , \new_[99244]_ , \new_[99247]_ , \new_[99250]_ ,
    \new_[99251]_ , \new_[99252]_ , \new_[99255]_ , \new_[99258]_ ,
    \new_[99259]_ , \new_[99262]_ , \new_[99265]_ , \new_[99266]_ ,
    \new_[99267]_ , \new_[99270]_ , \new_[99273]_ , \new_[99274]_ ,
    \new_[99277]_ , \new_[99280]_ , \new_[99281]_ , \new_[99282]_ ,
    \new_[99285]_ , \new_[99288]_ , \new_[99289]_ , \new_[99292]_ ,
    \new_[99295]_ , \new_[99296]_ , \new_[99297]_ , \new_[99300]_ ,
    \new_[99303]_ , \new_[99304]_ , \new_[99307]_ , \new_[99310]_ ,
    \new_[99311]_ , \new_[99312]_ , \new_[99315]_ , \new_[99318]_ ,
    \new_[99319]_ , \new_[99322]_ , \new_[99325]_ , \new_[99326]_ ,
    \new_[99327]_ , \new_[99330]_ , \new_[99333]_ , \new_[99334]_ ,
    \new_[99337]_ , \new_[99340]_ , \new_[99341]_ , \new_[99342]_ ,
    \new_[99345]_ , \new_[99348]_ , \new_[99349]_ , \new_[99352]_ ,
    \new_[99355]_ , \new_[99356]_ , \new_[99357]_ , \new_[99360]_ ,
    \new_[99363]_ , \new_[99364]_ , \new_[99367]_ , \new_[99370]_ ,
    \new_[99371]_ , \new_[99372]_ , \new_[99375]_ , \new_[99378]_ ,
    \new_[99379]_ , \new_[99382]_ , \new_[99385]_ , \new_[99386]_ ,
    \new_[99387]_ , \new_[99390]_ , \new_[99393]_ , \new_[99394]_ ,
    \new_[99397]_ , \new_[99400]_ , \new_[99401]_ , \new_[99402]_ ,
    \new_[99405]_ , \new_[99408]_ , \new_[99409]_ , \new_[99412]_ ,
    \new_[99415]_ , \new_[99416]_ , \new_[99417]_ , \new_[99420]_ ,
    \new_[99423]_ , \new_[99424]_ , \new_[99427]_ , \new_[99430]_ ,
    \new_[99431]_ , \new_[99432]_ , \new_[99435]_ , \new_[99438]_ ,
    \new_[99439]_ , \new_[99442]_ , \new_[99445]_ , \new_[99446]_ ,
    \new_[99447]_ , \new_[99450]_ , \new_[99453]_ , \new_[99454]_ ,
    \new_[99457]_ , \new_[99460]_ , \new_[99461]_ , \new_[99462]_ ,
    \new_[99465]_ , \new_[99468]_ , \new_[99469]_ , \new_[99472]_ ,
    \new_[99475]_ , \new_[99476]_ , \new_[99477]_ , \new_[99480]_ ,
    \new_[99483]_ , \new_[99484]_ , \new_[99487]_ , \new_[99490]_ ,
    \new_[99491]_ , \new_[99492]_ , \new_[99495]_ , \new_[99498]_ ,
    \new_[99499]_ , \new_[99502]_ , \new_[99505]_ , \new_[99506]_ ,
    \new_[99507]_ , \new_[99510]_ , \new_[99513]_ , \new_[99514]_ ,
    \new_[99517]_ , \new_[99520]_ , \new_[99521]_ , \new_[99522]_ ,
    \new_[99525]_ , \new_[99528]_ , \new_[99529]_ , \new_[99532]_ ,
    \new_[99535]_ , \new_[99536]_ , \new_[99537]_ , \new_[99540]_ ,
    \new_[99543]_ , \new_[99544]_ , \new_[99547]_ , \new_[99550]_ ,
    \new_[99551]_ , \new_[99552]_ , \new_[99555]_ , \new_[99558]_ ,
    \new_[99559]_ , \new_[99562]_ , \new_[99565]_ , \new_[99566]_ ,
    \new_[99567]_ , \new_[99570]_ , \new_[99573]_ , \new_[99574]_ ,
    \new_[99577]_ , \new_[99580]_ , \new_[99581]_ , \new_[99582]_ ,
    \new_[99585]_ , \new_[99588]_ , \new_[99589]_ , \new_[99592]_ ,
    \new_[99595]_ , \new_[99596]_ , \new_[99597]_ , \new_[99600]_ ,
    \new_[99603]_ , \new_[99604]_ , \new_[99607]_ , \new_[99610]_ ,
    \new_[99611]_ , \new_[99612]_ , \new_[99615]_ , \new_[99618]_ ,
    \new_[99619]_ , \new_[99622]_ , \new_[99625]_ , \new_[99626]_ ,
    \new_[99627]_ , \new_[99630]_ , \new_[99633]_ , \new_[99634]_ ,
    \new_[99637]_ , \new_[99640]_ , \new_[99641]_ , \new_[99642]_ ,
    \new_[99645]_ , \new_[99648]_ , \new_[99649]_ , \new_[99652]_ ,
    \new_[99655]_ , \new_[99656]_ , \new_[99657]_ , \new_[99660]_ ,
    \new_[99663]_ , \new_[99664]_ , \new_[99667]_ , \new_[99670]_ ,
    \new_[99671]_ , \new_[99672]_ , \new_[99675]_ , \new_[99678]_ ,
    \new_[99679]_ , \new_[99682]_ , \new_[99685]_ , \new_[99686]_ ,
    \new_[99687]_ , \new_[99690]_ , \new_[99693]_ , \new_[99694]_ ,
    \new_[99697]_ , \new_[99700]_ , \new_[99701]_ , \new_[99702]_ ,
    \new_[99705]_ , \new_[99708]_ , \new_[99709]_ , \new_[99712]_ ,
    \new_[99715]_ , \new_[99716]_ , \new_[99717]_ , \new_[99720]_ ,
    \new_[99723]_ , \new_[99724]_ , \new_[99727]_ , \new_[99730]_ ,
    \new_[99731]_ , \new_[99732]_ , \new_[99735]_ , \new_[99738]_ ,
    \new_[99739]_ , \new_[99742]_ , \new_[99745]_ , \new_[99746]_ ,
    \new_[99747]_ , \new_[99750]_ , \new_[99753]_ , \new_[99754]_ ,
    \new_[99757]_ , \new_[99760]_ , \new_[99761]_ , \new_[99762]_ ,
    \new_[99765]_ , \new_[99768]_ , \new_[99769]_ , \new_[99772]_ ,
    \new_[99775]_ , \new_[99776]_ , \new_[99777]_ , \new_[99780]_ ,
    \new_[99783]_ , \new_[99784]_ , \new_[99787]_ , \new_[99790]_ ,
    \new_[99791]_ , \new_[99792]_ , \new_[99795]_ , \new_[99798]_ ,
    \new_[99799]_ , \new_[99802]_ , \new_[99805]_ , \new_[99806]_ ,
    \new_[99807]_ , \new_[99810]_ , \new_[99813]_ , \new_[99814]_ ,
    \new_[99817]_ , \new_[99820]_ , \new_[99821]_ , \new_[99822]_ ,
    \new_[99825]_ , \new_[99828]_ , \new_[99829]_ , \new_[99832]_ ,
    \new_[99835]_ , \new_[99836]_ , \new_[99837]_ , \new_[99840]_ ,
    \new_[99843]_ , \new_[99844]_ , \new_[99847]_ , \new_[99850]_ ,
    \new_[99851]_ , \new_[99852]_ , \new_[99855]_ , \new_[99858]_ ,
    \new_[99859]_ , \new_[99862]_ , \new_[99865]_ , \new_[99866]_ ,
    \new_[99867]_ , \new_[99870]_ , \new_[99873]_ , \new_[99874]_ ,
    \new_[99877]_ , \new_[99880]_ , \new_[99881]_ , \new_[99882]_ ,
    \new_[99885]_ , \new_[99888]_ , \new_[99889]_ , \new_[99892]_ ,
    \new_[99895]_ , \new_[99896]_ , \new_[99897]_ , \new_[99900]_ ,
    \new_[99903]_ , \new_[99904]_ , \new_[99907]_ , \new_[99910]_ ,
    \new_[99911]_ , \new_[99912]_ , \new_[99915]_ , \new_[99918]_ ,
    \new_[99919]_ , \new_[99922]_ , \new_[99925]_ , \new_[99926]_ ,
    \new_[99927]_ , \new_[99930]_ , \new_[99933]_ , \new_[99934]_ ,
    \new_[99937]_ , \new_[99940]_ , \new_[99941]_ , \new_[99942]_ ,
    \new_[99945]_ , \new_[99948]_ , \new_[99949]_ , \new_[99952]_ ,
    \new_[99955]_ , \new_[99956]_ , \new_[99957]_ , \new_[99960]_ ,
    \new_[99963]_ , \new_[99964]_ , \new_[99967]_ , \new_[99970]_ ,
    \new_[99971]_ , \new_[99972]_ , \new_[99975]_ , \new_[99978]_ ,
    \new_[99979]_ , \new_[99982]_ , \new_[99985]_ , \new_[99986]_ ,
    \new_[99987]_ , \new_[99990]_ , \new_[99993]_ , \new_[99994]_ ,
    \new_[99997]_ , \new_[100000]_ , \new_[100001]_ , \new_[100002]_ ,
    \new_[100005]_ , \new_[100008]_ , \new_[100009]_ , \new_[100012]_ ,
    \new_[100015]_ , \new_[100016]_ , \new_[100017]_ , \new_[100020]_ ,
    \new_[100023]_ , \new_[100024]_ , \new_[100027]_ , \new_[100030]_ ,
    \new_[100031]_ , \new_[100032]_ , \new_[100035]_ , \new_[100038]_ ,
    \new_[100039]_ , \new_[100042]_ , \new_[100045]_ , \new_[100046]_ ,
    \new_[100047]_ , \new_[100050]_ , \new_[100053]_ , \new_[100054]_ ,
    \new_[100057]_ , \new_[100060]_ , \new_[100061]_ , \new_[100062]_ ,
    \new_[100065]_ , \new_[100068]_ , \new_[100069]_ , \new_[100072]_ ,
    \new_[100075]_ , \new_[100076]_ , \new_[100077]_ , \new_[100080]_ ,
    \new_[100083]_ , \new_[100084]_ , \new_[100087]_ , \new_[100090]_ ,
    \new_[100091]_ , \new_[100092]_ , \new_[100095]_ , \new_[100098]_ ,
    \new_[100099]_ , \new_[100102]_ , \new_[100105]_ , \new_[100106]_ ,
    \new_[100107]_ , \new_[100110]_ , \new_[100113]_ , \new_[100114]_ ,
    \new_[100117]_ , \new_[100120]_ , \new_[100121]_ , \new_[100122]_ ,
    \new_[100125]_ , \new_[100128]_ , \new_[100129]_ , \new_[100132]_ ,
    \new_[100135]_ , \new_[100136]_ , \new_[100137]_ , \new_[100140]_ ,
    \new_[100143]_ , \new_[100144]_ , \new_[100147]_ , \new_[100150]_ ,
    \new_[100151]_ , \new_[100152]_ , \new_[100155]_ , \new_[100158]_ ,
    \new_[100159]_ , \new_[100162]_ , \new_[100165]_ , \new_[100166]_ ,
    \new_[100167]_ , \new_[100170]_ , \new_[100173]_ , \new_[100174]_ ,
    \new_[100177]_ , \new_[100180]_ , \new_[100181]_ , \new_[100182]_ ,
    \new_[100185]_ , \new_[100188]_ , \new_[100189]_ , \new_[100192]_ ,
    \new_[100195]_ , \new_[100196]_ , \new_[100197]_ , \new_[100200]_ ,
    \new_[100203]_ , \new_[100204]_ , \new_[100207]_ , \new_[100210]_ ,
    \new_[100211]_ , \new_[100212]_ , \new_[100215]_ , \new_[100218]_ ,
    \new_[100219]_ , \new_[100222]_ , \new_[100225]_ , \new_[100226]_ ,
    \new_[100227]_ , \new_[100230]_ , \new_[100233]_ , \new_[100234]_ ,
    \new_[100237]_ , \new_[100240]_ , \new_[100241]_ , \new_[100242]_ ,
    \new_[100245]_ , \new_[100248]_ , \new_[100249]_ , \new_[100252]_ ,
    \new_[100255]_ , \new_[100256]_ , \new_[100257]_ , \new_[100260]_ ,
    \new_[100263]_ , \new_[100264]_ , \new_[100267]_ , \new_[100270]_ ,
    \new_[100271]_ , \new_[100272]_ , \new_[100275]_ , \new_[100278]_ ,
    \new_[100279]_ , \new_[100282]_ , \new_[100285]_ , \new_[100286]_ ,
    \new_[100287]_ , \new_[100290]_ , \new_[100293]_ , \new_[100294]_ ,
    \new_[100297]_ , \new_[100300]_ , \new_[100301]_ , \new_[100302]_ ,
    \new_[100305]_ , \new_[100308]_ , \new_[100309]_ , \new_[100312]_ ,
    \new_[100315]_ , \new_[100316]_ , \new_[100317]_ , \new_[100320]_ ,
    \new_[100323]_ , \new_[100324]_ , \new_[100327]_ , \new_[100330]_ ,
    \new_[100331]_ , \new_[100332]_ , \new_[100335]_ , \new_[100338]_ ,
    \new_[100339]_ , \new_[100342]_ , \new_[100345]_ , \new_[100346]_ ,
    \new_[100347]_ , \new_[100350]_ , \new_[100353]_ , \new_[100354]_ ,
    \new_[100357]_ , \new_[100360]_ , \new_[100361]_ , \new_[100362]_ ,
    \new_[100365]_ , \new_[100368]_ , \new_[100369]_ , \new_[100372]_ ,
    \new_[100375]_ , \new_[100376]_ , \new_[100377]_ , \new_[100380]_ ,
    \new_[100383]_ , \new_[100384]_ , \new_[100387]_ , \new_[100390]_ ,
    \new_[100391]_ , \new_[100392]_ , \new_[100395]_ , \new_[100398]_ ,
    \new_[100399]_ , \new_[100402]_ , \new_[100405]_ , \new_[100406]_ ,
    \new_[100407]_ , \new_[100410]_ , \new_[100413]_ , \new_[100414]_ ,
    \new_[100417]_ , \new_[100420]_ , \new_[100421]_ , \new_[100422]_ ,
    \new_[100425]_ , \new_[100428]_ , \new_[100429]_ , \new_[100432]_ ,
    \new_[100435]_ , \new_[100436]_ , \new_[100437]_ , \new_[100440]_ ,
    \new_[100443]_ , \new_[100444]_ , \new_[100447]_ , \new_[100450]_ ,
    \new_[100451]_ , \new_[100452]_ , \new_[100455]_ , \new_[100458]_ ,
    \new_[100459]_ , \new_[100462]_ , \new_[100465]_ , \new_[100466]_ ,
    \new_[100467]_ , \new_[100470]_ , \new_[100473]_ , \new_[100474]_ ,
    \new_[100477]_ , \new_[100480]_ , \new_[100481]_ , \new_[100482]_ ,
    \new_[100485]_ , \new_[100488]_ , \new_[100489]_ , \new_[100492]_ ,
    \new_[100495]_ , \new_[100496]_ , \new_[100497]_ , \new_[100500]_ ,
    \new_[100503]_ , \new_[100504]_ , \new_[100507]_ , \new_[100510]_ ,
    \new_[100511]_ , \new_[100512]_ , \new_[100515]_ , \new_[100518]_ ,
    \new_[100519]_ , \new_[100522]_ , \new_[100525]_ , \new_[100526]_ ,
    \new_[100527]_ , \new_[100530]_ , \new_[100533]_ , \new_[100534]_ ,
    \new_[100537]_ , \new_[100540]_ , \new_[100541]_ , \new_[100542]_ ,
    \new_[100545]_ , \new_[100548]_ , \new_[100549]_ , \new_[100552]_ ,
    \new_[100555]_ , \new_[100556]_ , \new_[100557]_ , \new_[100560]_ ,
    \new_[100563]_ , \new_[100564]_ , \new_[100567]_ , \new_[100570]_ ,
    \new_[100571]_ , \new_[100572]_ , \new_[100575]_ , \new_[100578]_ ,
    \new_[100579]_ , \new_[100582]_ , \new_[100585]_ , \new_[100586]_ ,
    \new_[100587]_ , \new_[100590]_ , \new_[100593]_ , \new_[100594]_ ,
    \new_[100597]_ , \new_[100600]_ , \new_[100601]_ , \new_[100602]_ ,
    \new_[100605]_ , \new_[100608]_ , \new_[100609]_ , \new_[100612]_ ,
    \new_[100615]_ , \new_[100616]_ , \new_[100617]_ , \new_[100620]_ ,
    \new_[100623]_ , \new_[100624]_ , \new_[100627]_ , \new_[100630]_ ,
    \new_[100631]_ , \new_[100632]_ , \new_[100635]_ , \new_[100638]_ ,
    \new_[100639]_ , \new_[100642]_ , \new_[100645]_ , \new_[100646]_ ,
    \new_[100647]_ , \new_[100650]_ , \new_[100653]_ , \new_[100654]_ ,
    \new_[100657]_ , \new_[100660]_ , \new_[100661]_ , \new_[100662]_ ,
    \new_[100665]_ , \new_[100668]_ , \new_[100669]_ , \new_[100672]_ ,
    \new_[100675]_ , \new_[100676]_ , \new_[100677]_ , \new_[100680]_ ,
    \new_[100683]_ , \new_[100684]_ , \new_[100687]_ , \new_[100690]_ ,
    \new_[100691]_ , \new_[100692]_ , \new_[100695]_ , \new_[100698]_ ,
    \new_[100699]_ , \new_[100702]_ , \new_[100705]_ , \new_[100706]_ ,
    \new_[100707]_ , \new_[100710]_ , \new_[100713]_ , \new_[100714]_ ,
    \new_[100717]_ , \new_[100720]_ , \new_[100721]_ , \new_[100722]_ ,
    \new_[100725]_ , \new_[100728]_ , \new_[100729]_ , \new_[100732]_ ,
    \new_[100735]_ , \new_[100736]_ , \new_[100737]_ , \new_[100740]_ ,
    \new_[100743]_ , \new_[100744]_ , \new_[100747]_ , \new_[100750]_ ,
    \new_[100751]_ , \new_[100752]_ , \new_[100755]_ , \new_[100758]_ ,
    \new_[100759]_ , \new_[100762]_ , \new_[100765]_ , \new_[100766]_ ,
    \new_[100767]_ , \new_[100770]_ , \new_[100773]_ , \new_[100774]_ ,
    \new_[100777]_ , \new_[100780]_ , \new_[100781]_ , \new_[100782]_ ,
    \new_[100785]_ , \new_[100788]_ , \new_[100789]_ , \new_[100792]_ ,
    \new_[100795]_ , \new_[100796]_ , \new_[100797]_ , \new_[100800]_ ,
    \new_[100803]_ , \new_[100804]_ , \new_[100807]_ , \new_[100810]_ ,
    \new_[100811]_ , \new_[100812]_ , \new_[100815]_ , \new_[100818]_ ,
    \new_[100819]_ , \new_[100822]_ , \new_[100825]_ , \new_[100826]_ ,
    \new_[100827]_ , \new_[100830]_ , \new_[100833]_ , \new_[100834]_ ,
    \new_[100837]_ , \new_[100840]_ , \new_[100841]_ , \new_[100842]_ ,
    \new_[100845]_ , \new_[100848]_ , \new_[100849]_ , \new_[100852]_ ,
    \new_[100855]_ , \new_[100856]_ , \new_[100857]_ , \new_[100860]_ ,
    \new_[100863]_ , \new_[100864]_ , \new_[100867]_ , \new_[100870]_ ,
    \new_[100871]_ , \new_[100872]_ , \new_[100875]_ , \new_[100878]_ ,
    \new_[100879]_ , \new_[100882]_ , \new_[100885]_ , \new_[100886]_ ,
    \new_[100887]_ , \new_[100890]_ , \new_[100893]_ , \new_[100894]_ ,
    \new_[100897]_ , \new_[100900]_ , \new_[100901]_ , \new_[100902]_ ,
    \new_[100905]_ , \new_[100908]_ , \new_[100909]_ , \new_[100912]_ ,
    \new_[100915]_ , \new_[100916]_ , \new_[100917]_ , \new_[100920]_ ,
    \new_[100923]_ , \new_[100924]_ , \new_[100927]_ , \new_[100930]_ ,
    \new_[100931]_ , \new_[100932]_ , \new_[100935]_ , \new_[100938]_ ,
    \new_[100939]_ , \new_[100942]_ , \new_[100945]_ , \new_[100946]_ ,
    \new_[100947]_ , \new_[100950]_ , \new_[100953]_ , \new_[100954]_ ,
    \new_[100957]_ , \new_[100960]_ , \new_[100961]_ , \new_[100962]_ ,
    \new_[100965]_ , \new_[100968]_ , \new_[100969]_ , \new_[100972]_ ,
    \new_[100975]_ , \new_[100976]_ , \new_[100977]_ , \new_[100980]_ ,
    \new_[100983]_ , \new_[100984]_ , \new_[100987]_ , \new_[100991]_ ,
    \new_[100992]_ , \new_[100993]_ , \new_[100994]_ , \new_[100997]_ ,
    \new_[101000]_ , \new_[101001]_ , \new_[101004]_ , \new_[101007]_ ,
    \new_[101008]_ , \new_[101009]_ , \new_[101012]_ , \new_[101015]_ ,
    \new_[101016]_ , \new_[101019]_ , \new_[101023]_ , \new_[101024]_ ,
    \new_[101025]_ , \new_[101026]_ , \new_[101029]_ , \new_[101032]_ ,
    \new_[101033]_ , \new_[101036]_ , \new_[101039]_ , \new_[101040]_ ,
    \new_[101041]_ , \new_[101044]_ , \new_[101047]_ , \new_[101048]_ ,
    \new_[101051]_ , \new_[101055]_ , \new_[101056]_ , \new_[101057]_ ,
    \new_[101058]_ , \new_[101061]_ , \new_[101064]_ , \new_[101065]_ ,
    \new_[101068]_ , \new_[101071]_ , \new_[101072]_ , \new_[101073]_ ,
    \new_[101076]_ , \new_[101079]_ , \new_[101080]_ , \new_[101083]_ ,
    \new_[101087]_ , \new_[101088]_ , \new_[101089]_ , \new_[101090]_ ,
    \new_[101093]_ , \new_[101096]_ , \new_[101097]_ , \new_[101100]_ ,
    \new_[101103]_ , \new_[101104]_ , \new_[101105]_ , \new_[101108]_ ,
    \new_[101111]_ , \new_[101112]_ , \new_[101115]_ , \new_[101119]_ ,
    \new_[101120]_ , \new_[101121]_ , \new_[101122]_ , \new_[101125]_ ,
    \new_[101128]_ , \new_[101129]_ , \new_[101132]_ , \new_[101135]_ ,
    \new_[101136]_ , \new_[101137]_ , \new_[101140]_ , \new_[101143]_ ,
    \new_[101144]_ , \new_[101147]_ , \new_[101151]_ , \new_[101152]_ ,
    \new_[101153]_ , \new_[101154]_ ;
  assign A109 = \new_[11314]_  | \new_[7543]_ ;
  assign \new_[1]_  = \new_[101154]_  & \new_[101137]_ ;
  assign \new_[2]_  = \new_[101122]_  & \new_[101105]_ ;
  assign \new_[3]_  = \new_[101090]_  & \new_[101073]_ ;
  assign \new_[4]_  = \new_[101058]_  & \new_[101041]_ ;
  assign \new_[5]_  = \new_[101026]_  & \new_[101009]_ ;
  assign \new_[6]_  = \new_[100994]_  & \new_[100977]_ ;
  assign \new_[7]_  = \new_[100962]_  & \new_[100947]_ ;
  assign \new_[8]_  = \new_[100932]_  & \new_[100917]_ ;
  assign \new_[9]_  = \new_[100902]_  & \new_[100887]_ ;
  assign \new_[10]_  = \new_[100872]_  & \new_[100857]_ ;
  assign \new_[11]_  = \new_[100842]_  & \new_[100827]_ ;
  assign \new_[12]_  = \new_[100812]_  & \new_[100797]_ ;
  assign \new_[13]_  = \new_[100782]_  & \new_[100767]_ ;
  assign \new_[14]_  = \new_[100752]_  & \new_[100737]_ ;
  assign \new_[15]_  = \new_[100722]_  & \new_[100707]_ ;
  assign \new_[16]_  = \new_[100692]_  & \new_[100677]_ ;
  assign \new_[17]_  = \new_[100662]_  & \new_[100647]_ ;
  assign \new_[18]_  = \new_[100632]_  & \new_[100617]_ ;
  assign \new_[19]_  = \new_[100602]_  & \new_[100587]_ ;
  assign \new_[20]_  = \new_[100572]_  & \new_[100557]_ ;
  assign \new_[21]_  = \new_[100542]_  & \new_[100527]_ ;
  assign \new_[22]_  = \new_[100512]_  & \new_[100497]_ ;
  assign \new_[23]_  = \new_[100482]_  & \new_[100467]_ ;
  assign \new_[24]_  = \new_[100452]_  & \new_[100437]_ ;
  assign \new_[25]_  = \new_[100422]_  & \new_[100407]_ ;
  assign \new_[26]_  = \new_[100392]_  & \new_[100377]_ ;
  assign \new_[27]_  = \new_[100362]_  & \new_[100347]_ ;
  assign \new_[28]_  = \new_[100332]_  & \new_[100317]_ ;
  assign \new_[29]_  = \new_[100302]_  & \new_[100287]_ ;
  assign \new_[30]_  = \new_[100272]_  & \new_[100257]_ ;
  assign \new_[31]_  = \new_[100242]_  & \new_[100227]_ ;
  assign \new_[32]_  = \new_[100212]_  & \new_[100197]_ ;
  assign \new_[33]_  = \new_[100182]_  & \new_[100167]_ ;
  assign \new_[34]_  = \new_[100152]_  & \new_[100137]_ ;
  assign \new_[35]_  = \new_[100122]_  & \new_[100107]_ ;
  assign \new_[36]_  = \new_[100092]_  & \new_[100077]_ ;
  assign \new_[37]_  = \new_[100062]_  & \new_[100047]_ ;
  assign \new_[38]_  = \new_[100032]_  & \new_[100017]_ ;
  assign \new_[39]_  = \new_[100002]_  & \new_[99987]_ ;
  assign \new_[40]_  = \new_[99972]_  & \new_[99957]_ ;
  assign \new_[41]_  = \new_[99942]_  & \new_[99927]_ ;
  assign \new_[42]_  = \new_[99912]_  & \new_[99897]_ ;
  assign \new_[43]_  = \new_[99882]_  & \new_[99867]_ ;
  assign \new_[44]_  = \new_[99852]_  & \new_[99837]_ ;
  assign \new_[45]_  = \new_[99822]_  & \new_[99807]_ ;
  assign \new_[46]_  = \new_[99792]_  & \new_[99777]_ ;
  assign \new_[47]_  = \new_[99762]_  & \new_[99747]_ ;
  assign \new_[48]_  = \new_[99732]_  & \new_[99717]_ ;
  assign \new_[49]_  = \new_[99702]_  & \new_[99687]_ ;
  assign \new_[50]_  = \new_[99672]_  & \new_[99657]_ ;
  assign \new_[51]_  = \new_[99642]_  & \new_[99627]_ ;
  assign \new_[52]_  = \new_[99612]_  & \new_[99597]_ ;
  assign \new_[53]_  = \new_[99582]_  & \new_[99567]_ ;
  assign \new_[54]_  = \new_[99552]_  & \new_[99537]_ ;
  assign \new_[55]_  = \new_[99522]_  & \new_[99507]_ ;
  assign \new_[56]_  = \new_[99492]_  & \new_[99477]_ ;
  assign \new_[57]_  = \new_[99462]_  & \new_[99447]_ ;
  assign \new_[58]_  = \new_[99432]_  & \new_[99417]_ ;
  assign \new_[59]_  = \new_[99402]_  & \new_[99387]_ ;
  assign \new_[60]_  = \new_[99372]_  & \new_[99357]_ ;
  assign \new_[61]_  = \new_[99342]_  & \new_[99327]_ ;
  assign \new_[62]_  = \new_[99312]_  & \new_[99297]_ ;
  assign \new_[63]_  = \new_[99282]_  & \new_[99267]_ ;
  assign \new_[64]_  = \new_[99252]_  & \new_[99237]_ ;
  assign \new_[65]_  = \new_[99222]_  & \new_[99207]_ ;
  assign \new_[66]_  = \new_[99192]_  & \new_[99177]_ ;
  assign \new_[67]_  = \new_[99162]_  & \new_[99147]_ ;
  assign \new_[68]_  = \new_[99132]_  & \new_[99117]_ ;
  assign \new_[69]_  = \new_[99102]_  & \new_[99087]_ ;
  assign \new_[70]_  = \new_[99072]_  & \new_[99057]_ ;
  assign \new_[71]_  = \new_[99042]_  & \new_[99027]_ ;
  assign \new_[72]_  = \new_[99012]_  & \new_[98997]_ ;
  assign \new_[73]_  = \new_[98982]_  & \new_[98967]_ ;
  assign \new_[74]_  = \new_[98952]_  & \new_[98937]_ ;
  assign \new_[75]_  = \new_[98922]_  & \new_[98907]_ ;
  assign \new_[76]_  = \new_[98892]_  & \new_[98877]_ ;
  assign \new_[77]_  = \new_[98862]_  & \new_[98847]_ ;
  assign \new_[78]_  = \new_[98832]_  & \new_[98817]_ ;
  assign \new_[79]_  = \new_[98802]_  & \new_[98787]_ ;
  assign \new_[80]_  = \new_[98772]_  & \new_[98757]_ ;
  assign \new_[81]_  = \new_[98742]_  & \new_[98727]_ ;
  assign \new_[82]_  = \new_[98712]_  & \new_[98697]_ ;
  assign \new_[83]_  = \new_[98682]_  & \new_[98667]_ ;
  assign \new_[84]_  = \new_[98652]_  & \new_[98637]_ ;
  assign \new_[85]_  = \new_[98622]_  & \new_[98607]_ ;
  assign \new_[86]_  = \new_[98592]_  & \new_[98577]_ ;
  assign \new_[87]_  = \new_[98562]_  & \new_[98547]_ ;
  assign \new_[88]_  = \new_[98532]_  & \new_[98517]_ ;
  assign \new_[89]_  = \new_[98502]_  & \new_[98487]_ ;
  assign \new_[90]_  = \new_[98472]_  & \new_[98457]_ ;
  assign \new_[91]_  = \new_[98442]_  & \new_[98427]_ ;
  assign \new_[92]_  = \new_[98412]_  & \new_[98397]_ ;
  assign \new_[93]_  = \new_[98382]_  & \new_[98367]_ ;
  assign \new_[94]_  = \new_[98352]_  & \new_[98337]_ ;
  assign \new_[95]_  = \new_[98322]_  & \new_[98307]_ ;
  assign \new_[96]_  = \new_[98292]_  & \new_[98277]_ ;
  assign \new_[97]_  = \new_[98262]_  & \new_[98247]_ ;
  assign \new_[98]_  = \new_[98232]_  & \new_[98217]_ ;
  assign \new_[99]_  = \new_[98202]_  & \new_[98187]_ ;
  assign \new_[100]_  = \new_[98172]_  & \new_[98157]_ ;
  assign \new_[101]_  = \new_[98142]_  & \new_[98127]_ ;
  assign \new_[102]_  = \new_[98112]_  & \new_[98097]_ ;
  assign \new_[103]_  = \new_[98082]_  & \new_[98067]_ ;
  assign \new_[104]_  = \new_[98052]_  & \new_[98037]_ ;
  assign \new_[105]_  = \new_[98022]_  & \new_[98007]_ ;
  assign \new_[106]_  = \new_[97992]_  & \new_[97977]_ ;
  assign \new_[107]_  = \new_[97962]_  & \new_[97947]_ ;
  assign \new_[108]_  = \new_[97932]_  & \new_[97917]_ ;
  assign \new_[109]_  = \new_[97902]_  & \new_[97887]_ ;
  assign \new_[110]_  = \new_[97872]_  & \new_[97857]_ ;
  assign \new_[111]_  = \new_[97842]_  & \new_[97827]_ ;
  assign \new_[112]_  = \new_[97812]_  & \new_[97797]_ ;
  assign \new_[113]_  = \new_[97782]_  & \new_[97767]_ ;
  assign \new_[114]_  = \new_[97752]_  & \new_[97737]_ ;
  assign \new_[115]_  = \new_[97722]_  & \new_[97707]_ ;
  assign \new_[116]_  = \new_[97692]_  & \new_[97677]_ ;
  assign \new_[117]_  = \new_[97662]_  & \new_[97647]_ ;
  assign \new_[118]_  = \new_[97632]_  & \new_[97617]_ ;
  assign \new_[119]_  = \new_[97602]_  & \new_[97587]_ ;
  assign \new_[120]_  = \new_[97572]_  & \new_[97557]_ ;
  assign \new_[121]_  = \new_[97542]_  & \new_[97527]_ ;
  assign \new_[122]_  = \new_[97514]_  & \new_[97499]_ ;
  assign \new_[123]_  = \new_[97486]_  & \new_[97471]_ ;
  assign \new_[124]_  = \new_[97458]_  & \new_[97443]_ ;
  assign \new_[125]_  = \new_[97430]_  & \new_[97415]_ ;
  assign \new_[126]_  = \new_[97402]_  & \new_[97387]_ ;
  assign \new_[127]_  = \new_[97374]_  & \new_[97359]_ ;
  assign \new_[128]_  = \new_[97346]_  & \new_[97331]_ ;
  assign \new_[129]_  = \new_[97318]_  & \new_[97303]_ ;
  assign \new_[130]_  = \new_[97290]_  & \new_[97275]_ ;
  assign \new_[131]_  = \new_[97262]_  & \new_[97247]_ ;
  assign \new_[132]_  = \new_[97234]_  & \new_[97219]_ ;
  assign \new_[133]_  = \new_[97206]_  & \new_[97191]_ ;
  assign \new_[134]_  = \new_[97178]_  & \new_[97163]_ ;
  assign \new_[135]_  = \new_[97150]_  & \new_[97135]_ ;
  assign \new_[136]_  = \new_[97122]_  & \new_[97107]_ ;
  assign \new_[137]_  = \new_[97094]_  & \new_[97079]_ ;
  assign \new_[138]_  = \new_[97066]_  & \new_[97051]_ ;
  assign \new_[139]_  = \new_[97038]_  & \new_[97023]_ ;
  assign \new_[140]_  = \new_[97010]_  & \new_[96995]_ ;
  assign \new_[141]_  = \new_[96982]_  & \new_[96967]_ ;
  assign \new_[142]_  = \new_[96954]_  & \new_[96939]_ ;
  assign \new_[143]_  = \new_[96926]_  & \new_[96911]_ ;
  assign \new_[144]_  = \new_[96898]_  & \new_[96883]_ ;
  assign \new_[145]_  = \new_[96870]_  & \new_[96855]_ ;
  assign \new_[146]_  = \new_[96842]_  & \new_[96827]_ ;
  assign \new_[147]_  = \new_[96814]_  & \new_[96799]_ ;
  assign \new_[148]_  = \new_[96786]_  & \new_[96771]_ ;
  assign \new_[149]_  = \new_[96758]_  & \new_[96743]_ ;
  assign \new_[150]_  = \new_[96730]_  & \new_[96715]_ ;
  assign \new_[151]_  = \new_[96702]_  & \new_[96687]_ ;
  assign \new_[152]_  = \new_[96674]_  & \new_[96659]_ ;
  assign \new_[153]_  = \new_[96646]_  & \new_[96631]_ ;
  assign \new_[154]_  = \new_[96618]_  & \new_[96603]_ ;
  assign \new_[155]_  = \new_[96590]_  & \new_[96575]_ ;
  assign \new_[156]_  = \new_[96562]_  & \new_[96547]_ ;
  assign \new_[157]_  = \new_[96534]_  & \new_[96519]_ ;
  assign \new_[158]_  = \new_[96506]_  & \new_[96491]_ ;
  assign \new_[159]_  = \new_[96478]_  & \new_[96463]_ ;
  assign \new_[160]_  = \new_[96450]_  & \new_[96435]_ ;
  assign \new_[161]_  = \new_[96422]_  & \new_[96407]_ ;
  assign \new_[162]_  = \new_[96394]_  & \new_[96379]_ ;
  assign \new_[163]_  = \new_[96366]_  & \new_[96351]_ ;
  assign \new_[164]_  = \new_[96338]_  & \new_[96323]_ ;
  assign \new_[165]_  = \new_[96310]_  & \new_[96295]_ ;
  assign \new_[166]_  = \new_[96282]_  & \new_[96267]_ ;
  assign \new_[167]_  = \new_[96254]_  & \new_[96239]_ ;
  assign \new_[168]_  = \new_[96226]_  & \new_[96211]_ ;
  assign \new_[169]_  = \new_[96198]_  & \new_[96183]_ ;
  assign \new_[170]_  = \new_[96170]_  & \new_[96155]_ ;
  assign \new_[171]_  = \new_[96142]_  & \new_[96127]_ ;
  assign \new_[172]_  = \new_[96114]_  & \new_[96099]_ ;
  assign \new_[173]_  = \new_[96086]_  & \new_[96071]_ ;
  assign \new_[174]_  = \new_[96058]_  & \new_[96043]_ ;
  assign \new_[175]_  = \new_[96030]_  & \new_[96015]_ ;
  assign \new_[176]_  = \new_[96002]_  & \new_[95987]_ ;
  assign \new_[177]_  = \new_[95974]_  & \new_[95959]_ ;
  assign \new_[178]_  = \new_[95946]_  & \new_[95931]_ ;
  assign \new_[179]_  = \new_[95918]_  & \new_[95903]_ ;
  assign \new_[180]_  = \new_[95890]_  & \new_[95875]_ ;
  assign \new_[181]_  = \new_[95862]_  & \new_[95847]_ ;
  assign \new_[182]_  = \new_[95834]_  & \new_[95819]_ ;
  assign \new_[183]_  = \new_[95806]_  & \new_[95791]_ ;
  assign \new_[184]_  = \new_[95778]_  & \new_[95763]_ ;
  assign \new_[185]_  = \new_[95750]_  & \new_[95735]_ ;
  assign \new_[186]_  = \new_[95722]_  & \new_[95707]_ ;
  assign \new_[187]_  = \new_[95694]_  & \new_[95679]_ ;
  assign \new_[188]_  = \new_[95666]_  & \new_[95651]_ ;
  assign \new_[189]_  = \new_[95638]_  & \new_[95623]_ ;
  assign \new_[190]_  = \new_[95610]_  & \new_[95595]_ ;
  assign \new_[191]_  = \new_[95582]_  & \new_[95567]_ ;
  assign \new_[192]_  = \new_[95554]_  & \new_[95539]_ ;
  assign \new_[193]_  = \new_[95526]_  & \new_[95511]_ ;
  assign \new_[194]_  = \new_[95498]_  & \new_[95483]_ ;
  assign \new_[195]_  = \new_[95470]_  & \new_[95455]_ ;
  assign \new_[196]_  = \new_[95442]_  & \new_[95427]_ ;
  assign \new_[197]_  = \new_[95414]_  & \new_[95399]_ ;
  assign \new_[198]_  = \new_[95386]_  & \new_[95371]_ ;
  assign \new_[199]_  = \new_[95358]_  & \new_[95343]_ ;
  assign \new_[200]_  = \new_[95330]_  & \new_[95315]_ ;
  assign \new_[201]_  = \new_[95302]_  & \new_[95287]_ ;
  assign \new_[202]_  = \new_[95274]_  & \new_[95259]_ ;
  assign \new_[203]_  = \new_[95246]_  & \new_[95231]_ ;
  assign \new_[204]_  = \new_[95218]_  & \new_[95203]_ ;
  assign \new_[205]_  = \new_[95190]_  & \new_[95175]_ ;
  assign \new_[206]_  = \new_[95162]_  & \new_[95147]_ ;
  assign \new_[207]_  = \new_[95134]_  & \new_[95119]_ ;
  assign \new_[208]_  = \new_[95106]_  & \new_[95091]_ ;
  assign \new_[209]_  = \new_[95078]_  & \new_[95063]_ ;
  assign \new_[210]_  = \new_[95050]_  & \new_[95035]_ ;
  assign \new_[211]_  = \new_[95022]_  & \new_[95007]_ ;
  assign \new_[212]_  = \new_[94994]_  & \new_[94979]_ ;
  assign \new_[213]_  = \new_[94966]_  & \new_[94951]_ ;
  assign \new_[214]_  = \new_[94938]_  & \new_[94923]_ ;
  assign \new_[215]_  = \new_[94910]_  & \new_[94895]_ ;
  assign \new_[216]_  = \new_[94882]_  & \new_[94867]_ ;
  assign \new_[217]_  = \new_[94854]_  & \new_[94839]_ ;
  assign \new_[218]_  = \new_[94826]_  & \new_[94811]_ ;
  assign \new_[219]_  = \new_[94798]_  & \new_[94783]_ ;
  assign \new_[220]_  = \new_[94770]_  & \new_[94755]_ ;
  assign \new_[221]_  = \new_[94742]_  & \new_[94727]_ ;
  assign \new_[222]_  = \new_[94714]_  & \new_[94699]_ ;
  assign \new_[223]_  = \new_[94686]_  & \new_[94671]_ ;
  assign \new_[224]_  = \new_[94658]_  & \new_[94643]_ ;
  assign \new_[225]_  = \new_[94630]_  & \new_[94615]_ ;
  assign \new_[226]_  = \new_[94602]_  & \new_[94587]_ ;
  assign \new_[227]_  = \new_[94574]_  & \new_[94559]_ ;
  assign \new_[228]_  = \new_[94546]_  & \new_[94531]_ ;
  assign \new_[229]_  = \new_[94518]_  & \new_[94503]_ ;
  assign \new_[230]_  = \new_[94490]_  & \new_[94475]_ ;
  assign \new_[231]_  = \new_[94462]_  & \new_[94447]_ ;
  assign \new_[232]_  = \new_[94434]_  & \new_[94419]_ ;
  assign \new_[233]_  = \new_[94406]_  & \new_[94391]_ ;
  assign \new_[234]_  = \new_[94378]_  & \new_[94363]_ ;
  assign \new_[235]_  = \new_[94350]_  & \new_[94335]_ ;
  assign \new_[236]_  = \new_[94322]_  & \new_[94307]_ ;
  assign \new_[237]_  = \new_[94294]_  & \new_[94279]_ ;
  assign \new_[238]_  = \new_[94266]_  & \new_[94251]_ ;
  assign \new_[239]_  = \new_[94238]_  & \new_[94223]_ ;
  assign \new_[240]_  = \new_[94210]_  & \new_[94195]_ ;
  assign \new_[241]_  = \new_[94182]_  & \new_[94167]_ ;
  assign \new_[242]_  = \new_[94154]_  & \new_[94139]_ ;
  assign \new_[243]_  = \new_[94126]_  & \new_[94111]_ ;
  assign \new_[244]_  = \new_[94098]_  & \new_[94083]_ ;
  assign \new_[245]_  = \new_[94070]_  & \new_[94055]_ ;
  assign \new_[246]_  = \new_[94042]_  & \new_[94027]_ ;
  assign \new_[247]_  = \new_[94014]_  & \new_[93999]_ ;
  assign \new_[248]_  = \new_[93986]_  & \new_[93971]_ ;
  assign \new_[249]_  = \new_[93958]_  & \new_[93943]_ ;
  assign \new_[250]_  = \new_[93930]_  & \new_[93915]_ ;
  assign \new_[251]_  = \new_[93902]_  & \new_[93887]_ ;
  assign \new_[252]_  = \new_[93874]_  & \new_[93859]_ ;
  assign \new_[253]_  = \new_[93846]_  & \new_[93831]_ ;
  assign \new_[254]_  = \new_[93818]_  & \new_[93803]_ ;
  assign \new_[255]_  = \new_[93790]_  & \new_[93775]_ ;
  assign \new_[256]_  = \new_[93762]_  & \new_[93747]_ ;
  assign \new_[257]_  = \new_[93734]_  & \new_[93719]_ ;
  assign \new_[258]_  = \new_[93706]_  & \new_[93691]_ ;
  assign \new_[259]_  = \new_[93678]_  & \new_[93663]_ ;
  assign \new_[260]_  = \new_[93650]_  & \new_[93635]_ ;
  assign \new_[261]_  = \new_[93622]_  & \new_[93607]_ ;
  assign \new_[262]_  = \new_[93594]_  & \new_[93579]_ ;
  assign \new_[263]_  = \new_[93566]_  & \new_[93551]_ ;
  assign \new_[264]_  = \new_[93538]_  & \new_[93523]_ ;
  assign \new_[265]_  = \new_[93510]_  & \new_[93495]_ ;
  assign \new_[266]_  = \new_[93482]_  & \new_[93467]_ ;
  assign \new_[267]_  = \new_[93454]_  & \new_[93439]_ ;
  assign \new_[268]_  = \new_[93426]_  & \new_[93411]_ ;
  assign \new_[269]_  = \new_[93398]_  & \new_[93383]_ ;
  assign \new_[270]_  = \new_[93370]_  & \new_[93355]_ ;
  assign \new_[271]_  = \new_[93342]_  & \new_[93327]_ ;
  assign \new_[272]_  = \new_[93314]_  & \new_[93299]_ ;
  assign \new_[273]_  = \new_[93286]_  & \new_[93271]_ ;
  assign \new_[274]_  = \new_[93258]_  & \new_[93243]_ ;
  assign \new_[275]_  = \new_[93230]_  & \new_[93215]_ ;
  assign \new_[276]_  = \new_[93202]_  & \new_[93187]_ ;
  assign \new_[277]_  = \new_[93174]_  & \new_[93159]_ ;
  assign \new_[278]_  = \new_[93146]_  & \new_[93131]_ ;
  assign \new_[279]_  = \new_[93118]_  & \new_[93103]_ ;
  assign \new_[280]_  = \new_[93090]_  & \new_[93075]_ ;
  assign \new_[281]_  = \new_[93062]_  & \new_[93047]_ ;
  assign \new_[282]_  = \new_[93034]_  & \new_[93019]_ ;
  assign \new_[283]_  = \new_[93006]_  & \new_[92991]_ ;
  assign \new_[284]_  = \new_[92978]_  & \new_[92963]_ ;
  assign \new_[285]_  = \new_[92950]_  & \new_[92935]_ ;
  assign \new_[286]_  = \new_[92922]_  & \new_[92907]_ ;
  assign \new_[287]_  = \new_[92894]_  & \new_[92879]_ ;
  assign \new_[288]_  = \new_[92866]_  & \new_[92851]_ ;
  assign \new_[289]_  = \new_[92838]_  & \new_[92823]_ ;
  assign \new_[290]_  = \new_[92810]_  & \new_[92795]_ ;
  assign \new_[291]_  = \new_[92782]_  & \new_[92767]_ ;
  assign \new_[292]_  = \new_[92754]_  & \new_[92739]_ ;
  assign \new_[293]_  = \new_[92726]_  & \new_[92711]_ ;
  assign \new_[294]_  = \new_[92698]_  & \new_[92683]_ ;
  assign \new_[295]_  = \new_[92670]_  & \new_[92655]_ ;
  assign \new_[296]_  = \new_[92642]_  & \new_[92627]_ ;
  assign \new_[297]_  = \new_[92614]_  & \new_[92599]_ ;
  assign \new_[298]_  = \new_[92586]_  & \new_[92571]_ ;
  assign \new_[299]_  = \new_[92558]_  & \new_[92543]_ ;
  assign \new_[300]_  = \new_[92530]_  & \new_[92515]_ ;
  assign \new_[301]_  = \new_[92502]_  & \new_[92487]_ ;
  assign \new_[302]_  = \new_[92474]_  & \new_[92459]_ ;
  assign \new_[303]_  = \new_[92446]_  & \new_[92431]_ ;
  assign \new_[304]_  = \new_[92418]_  & \new_[92403]_ ;
  assign \new_[305]_  = \new_[92390]_  & \new_[92375]_ ;
  assign \new_[306]_  = \new_[92362]_  & \new_[92347]_ ;
  assign \new_[307]_  = \new_[92334]_  & \new_[92319]_ ;
  assign \new_[308]_  = \new_[92306]_  & \new_[92291]_ ;
  assign \new_[309]_  = \new_[92278]_  & \new_[92263]_ ;
  assign \new_[310]_  = \new_[92250]_  & \new_[92235]_ ;
  assign \new_[311]_  = \new_[92222]_  & \new_[92207]_ ;
  assign \new_[312]_  = \new_[92194]_  & \new_[92179]_ ;
  assign \new_[313]_  = \new_[92166]_  & \new_[92151]_ ;
  assign \new_[314]_  = \new_[92138]_  & \new_[92123]_ ;
  assign \new_[315]_  = \new_[92110]_  & \new_[92095]_ ;
  assign \new_[316]_  = \new_[92082]_  & \new_[92067]_ ;
  assign \new_[317]_  = \new_[92054]_  & \new_[92039]_ ;
  assign \new_[318]_  = \new_[92026]_  & \new_[92011]_ ;
  assign \new_[319]_  = \new_[91998]_  & \new_[91983]_ ;
  assign \new_[320]_  = \new_[91970]_  & \new_[91955]_ ;
  assign \new_[321]_  = \new_[91942]_  & \new_[91927]_ ;
  assign \new_[322]_  = \new_[91914]_  & \new_[91899]_ ;
  assign \new_[323]_  = \new_[91886]_  & \new_[91871]_ ;
  assign \new_[324]_  = \new_[91858]_  & \new_[91843]_ ;
  assign \new_[325]_  = \new_[91830]_  & \new_[91815]_ ;
  assign \new_[326]_  = \new_[91802]_  & \new_[91787]_ ;
  assign \new_[327]_  = \new_[91774]_  & \new_[91759]_ ;
  assign \new_[328]_  = \new_[91746]_  & \new_[91731]_ ;
  assign \new_[329]_  = \new_[91718]_  & \new_[91703]_ ;
  assign \new_[330]_  = \new_[91690]_  & \new_[91675]_ ;
  assign \new_[331]_  = \new_[91662]_  & \new_[91647]_ ;
  assign \new_[332]_  = \new_[91634]_  & \new_[91619]_ ;
  assign \new_[333]_  = \new_[91606]_  & \new_[91591]_ ;
  assign \new_[334]_  = \new_[91578]_  & \new_[91563]_ ;
  assign \new_[335]_  = \new_[91550]_  & \new_[91535]_ ;
  assign \new_[336]_  = \new_[91522]_  & \new_[91507]_ ;
  assign \new_[337]_  = \new_[91494]_  & \new_[91479]_ ;
  assign \new_[338]_  = \new_[91466]_  & \new_[91451]_ ;
  assign \new_[339]_  = \new_[91438]_  & \new_[91423]_ ;
  assign \new_[340]_  = \new_[91410]_  & \new_[91395]_ ;
  assign \new_[341]_  = \new_[91382]_  & \new_[91367]_ ;
  assign \new_[342]_  = \new_[91354]_  & \new_[91339]_ ;
  assign \new_[343]_  = \new_[91326]_  & \new_[91311]_ ;
  assign \new_[344]_  = \new_[91298]_  & \new_[91283]_ ;
  assign \new_[345]_  = \new_[91270]_  & \new_[91255]_ ;
  assign \new_[346]_  = \new_[91242]_  & \new_[91227]_ ;
  assign \new_[347]_  = \new_[91214]_  & \new_[91199]_ ;
  assign \new_[348]_  = \new_[91186]_  & \new_[91171]_ ;
  assign \new_[349]_  = \new_[91158]_  & \new_[91143]_ ;
  assign \new_[350]_  = \new_[91130]_  & \new_[91115]_ ;
  assign \new_[351]_  = \new_[91102]_  & \new_[91087]_ ;
  assign \new_[352]_  = \new_[91074]_  & \new_[91059]_ ;
  assign \new_[353]_  = \new_[91046]_  & \new_[91031]_ ;
  assign \new_[354]_  = \new_[91018]_  & \new_[91003]_ ;
  assign \new_[355]_  = \new_[90990]_  & \new_[90975]_ ;
  assign \new_[356]_  = \new_[90962]_  & \new_[90947]_ ;
  assign \new_[357]_  = \new_[90934]_  & \new_[90919]_ ;
  assign \new_[358]_  = \new_[90906]_  & \new_[90891]_ ;
  assign \new_[359]_  = \new_[90878]_  & \new_[90863]_ ;
  assign \new_[360]_  = \new_[90850]_  & \new_[90835]_ ;
  assign \new_[361]_  = \new_[90822]_  & \new_[90807]_ ;
  assign \new_[362]_  = \new_[90794]_  & \new_[90779]_ ;
  assign \new_[363]_  = \new_[90766]_  & \new_[90751]_ ;
  assign \new_[364]_  = \new_[90738]_  & \new_[90723]_ ;
  assign \new_[365]_  = \new_[90710]_  & \new_[90695]_ ;
  assign \new_[366]_  = \new_[90682]_  & \new_[90667]_ ;
  assign \new_[367]_  = \new_[90654]_  & \new_[90639]_ ;
  assign \new_[368]_  = \new_[90626]_  & \new_[90611]_ ;
  assign \new_[369]_  = \new_[90598]_  & \new_[90583]_ ;
  assign \new_[370]_  = \new_[90570]_  & \new_[90555]_ ;
  assign \new_[371]_  = \new_[90542]_  & \new_[90527]_ ;
  assign \new_[372]_  = \new_[90514]_  & \new_[90499]_ ;
  assign \new_[373]_  = \new_[90486]_  & \new_[90471]_ ;
  assign \new_[374]_  = \new_[90458]_  & \new_[90443]_ ;
  assign \new_[375]_  = \new_[90430]_  & \new_[90415]_ ;
  assign \new_[376]_  = \new_[90402]_  & \new_[90387]_ ;
  assign \new_[377]_  = \new_[90374]_  & \new_[90359]_ ;
  assign \new_[378]_  = \new_[90346]_  & \new_[90331]_ ;
  assign \new_[379]_  = \new_[90318]_  & \new_[90303]_ ;
  assign \new_[380]_  = \new_[90290]_  & \new_[90275]_ ;
  assign \new_[381]_  = \new_[90262]_  & \new_[90247]_ ;
  assign \new_[382]_  = \new_[90234]_  & \new_[90219]_ ;
  assign \new_[383]_  = \new_[90206]_  & \new_[90191]_ ;
  assign \new_[384]_  = \new_[90178]_  & \new_[90163]_ ;
  assign \new_[385]_  = \new_[90150]_  & \new_[90135]_ ;
  assign \new_[386]_  = \new_[90122]_  & \new_[90107]_ ;
  assign \new_[387]_  = \new_[90094]_  & \new_[90079]_ ;
  assign \new_[388]_  = \new_[90066]_  & \new_[90051]_ ;
  assign \new_[389]_  = \new_[90038]_  & \new_[90023]_ ;
  assign \new_[390]_  = \new_[90010]_  & \new_[89995]_ ;
  assign \new_[391]_  = \new_[89982]_  & \new_[89967]_ ;
  assign \new_[392]_  = \new_[89954]_  & \new_[89939]_ ;
  assign \new_[393]_  = \new_[89926]_  & \new_[89911]_ ;
  assign \new_[394]_  = \new_[89898]_  & \new_[89883]_ ;
  assign \new_[395]_  = \new_[89870]_  & \new_[89855]_ ;
  assign \new_[396]_  = \new_[89842]_  & \new_[89827]_ ;
  assign \new_[397]_  = \new_[89814]_  & \new_[89799]_ ;
  assign \new_[398]_  = \new_[89786]_  & \new_[89771]_ ;
  assign \new_[399]_  = \new_[89758]_  & \new_[89743]_ ;
  assign \new_[400]_  = \new_[89730]_  & \new_[89715]_ ;
  assign \new_[401]_  = \new_[89702]_  & \new_[89687]_ ;
  assign \new_[402]_  = \new_[89674]_  & \new_[89659]_ ;
  assign \new_[403]_  = \new_[89646]_  & \new_[89631]_ ;
  assign \new_[404]_  = \new_[89618]_  & \new_[89603]_ ;
  assign \new_[405]_  = \new_[89590]_  & \new_[89575]_ ;
  assign \new_[406]_  = \new_[89562]_  & \new_[89547]_ ;
  assign \new_[407]_  = \new_[89534]_  & \new_[89519]_ ;
  assign \new_[408]_  = \new_[89506]_  & \new_[89491]_ ;
  assign \new_[409]_  = \new_[89478]_  & \new_[89463]_ ;
  assign \new_[410]_  = \new_[89450]_  & \new_[89435]_ ;
  assign \new_[411]_  = \new_[89422]_  & \new_[89407]_ ;
  assign \new_[412]_  = \new_[89394]_  & \new_[89379]_ ;
  assign \new_[413]_  = \new_[89366]_  & \new_[89351]_ ;
  assign \new_[414]_  = \new_[89338]_  & \new_[89323]_ ;
  assign \new_[415]_  = \new_[89310]_  & \new_[89295]_ ;
  assign \new_[416]_  = \new_[89282]_  & \new_[89267]_ ;
  assign \new_[417]_  = \new_[89254]_  & \new_[89239]_ ;
  assign \new_[418]_  = \new_[89226]_  & \new_[89211]_ ;
  assign \new_[419]_  = \new_[89198]_  & \new_[89183]_ ;
  assign \new_[420]_  = \new_[89170]_  & \new_[89155]_ ;
  assign \new_[421]_  = \new_[89142]_  & \new_[89127]_ ;
  assign \new_[422]_  = \new_[89114]_  & \new_[89099]_ ;
  assign \new_[423]_  = \new_[89086]_  & \new_[89071]_ ;
  assign \new_[424]_  = \new_[89058]_  & \new_[89043]_ ;
  assign \new_[425]_  = \new_[89030]_  & \new_[89015]_ ;
  assign \new_[426]_  = \new_[89002]_  & \new_[88987]_ ;
  assign \new_[427]_  = \new_[88974]_  & \new_[88959]_ ;
  assign \new_[428]_  = \new_[88946]_  & \new_[88931]_ ;
  assign \new_[429]_  = \new_[88918]_  & \new_[88903]_ ;
  assign \new_[430]_  = \new_[88890]_  & \new_[88875]_ ;
  assign \new_[431]_  = \new_[88862]_  & \new_[88847]_ ;
  assign \new_[432]_  = \new_[88834]_  & \new_[88819]_ ;
  assign \new_[433]_  = \new_[88806]_  & \new_[88791]_ ;
  assign \new_[434]_  = \new_[88778]_  & \new_[88763]_ ;
  assign \new_[435]_  = \new_[88750]_  & \new_[88735]_ ;
  assign \new_[436]_  = \new_[88722]_  & \new_[88707]_ ;
  assign \new_[437]_  = \new_[88694]_  & \new_[88679]_ ;
  assign \new_[438]_  = \new_[88666]_  & \new_[88651]_ ;
  assign \new_[439]_  = \new_[88638]_  & \new_[88623]_ ;
  assign \new_[440]_  = \new_[88610]_  & \new_[88595]_ ;
  assign \new_[441]_  = \new_[88582]_  & \new_[88567]_ ;
  assign \new_[442]_  = \new_[88554]_  & \new_[88539]_ ;
  assign \new_[443]_  = \new_[88526]_  & \new_[88511]_ ;
  assign \new_[444]_  = \new_[88498]_  & \new_[88483]_ ;
  assign \new_[445]_  = \new_[88470]_  & \new_[88455]_ ;
  assign \new_[446]_  = \new_[88442]_  & \new_[88427]_ ;
  assign \new_[447]_  = \new_[88414]_  & \new_[88399]_ ;
  assign \new_[448]_  = \new_[88386]_  & \new_[88371]_ ;
  assign \new_[449]_  = \new_[88358]_  & \new_[88343]_ ;
  assign \new_[450]_  = \new_[88330]_  & \new_[88315]_ ;
  assign \new_[451]_  = \new_[88302]_  & \new_[88287]_ ;
  assign \new_[452]_  = \new_[88274]_  & \new_[88259]_ ;
  assign \new_[453]_  = \new_[88246]_  & \new_[88231]_ ;
  assign \new_[454]_  = \new_[88218]_  & \new_[88203]_ ;
  assign \new_[455]_  = \new_[88190]_  & \new_[88175]_ ;
  assign \new_[456]_  = \new_[88162]_  & \new_[88147]_ ;
  assign \new_[457]_  = \new_[88134]_  & \new_[88119]_ ;
  assign \new_[458]_  = \new_[88106]_  & \new_[88091]_ ;
  assign \new_[459]_  = \new_[88078]_  & \new_[88063]_ ;
  assign \new_[460]_  = \new_[88050]_  & \new_[88035]_ ;
  assign \new_[461]_  = \new_[88022]_  & \new_[88007]_ ;
  assign \new_[462]_  = \new_[87994]_  & \new_[87979]_ ;
  assign \new_[463]_  = \new_[87966]_  & \new_[87951]_ ;
  assign \new_[464]_  = \new_[87938]_  & \new_[87923]_ ;
  assign \new_[465]_  = \new_[87910]_  & \new_[87895]_ ;
  assign \new_[466]_  = \new_[87882]_  & \new_[87867]_ ;
  assign \new_[467]_  = \new_[87854]_  & \new_[87839]_ ;
  assign \new_[468]_  = \new_[87826]_  & \new_[87811]_ ;
  assign \new_[469]_  = \new_[87798]_  & \new_[87783]_ ;
  assign \new_[470]_  = \new_[87770]_  & \new_[87755]_ ;
  assign \new_[471]_  = \new_[87742]_  & \new_[87727]_ ;
  assign \new_[472]_  = \new_[87714]_  & \new_[87699]_ ;
  assign \new_[473]_  = \new_[87686]_  & \new_[87671]_ ;
  assign \new_[474]_  = \new_[87658]_  & \new_[87643]_ ;
  assign \new_[475]_  = \new_[87630]_  & \new_[87615]_ ;
  assign \new_[476]_  = \new_[87602]_  & \new_[87587]_ ;
  assign \new_[477]_  = \new_[87574]_  & \new_[87559]_ ;
  assign \new_[478]_  = \new_[87546]_  & \new_[87531]_ ;
  assign \new_[479]_  = \new_[87518]_  & \new_[87503]_ ;
  assign \new_[480]_  = \new_[87490]_  & \new_[87475]_ ;
  assign \new_[481]_  = \new_[87462]_  & \new_[87447]_ ;
  assign \new_[482]_  = \new_[87434]_  & \new_[87419]_ ;
  assign \new_[483]_  = \new_[87406]_  & \new_[87391]_ ;
  assign \new_[484]_  = \new_[87378]_  & \new_[87363]_ ;
  assign \new_[485]_  = \new_[87350]_  & \new_[87335]_ ;
  assign \new_[486]_  = \new_[87322]_  & \new_[87307]_ ;
  assign \new_[487]_  = \new_[87294]_  & \new_[87279]_ ;
  assign \new_[488]_  = \new_[87266]_  & \new_[87251]_ ;
  assign \new_[489]_  = \new_[87238]_  & \new_[87223]_ ;
  assign \new_[490]_  = \new_[87210]_  & \new_[87195]_ ;
  assign \new_[491]_  = \new_[87182]_  & \new_[87167]_ ;
  assign \new_[492]_  = \new_[87154]_  & \new_[87139]_ ;
  assign \new_[493]_  = \new_[87126]_  & \new_[87111]_ ;
  assign \new_[494]_  = \new_[87098]_  & \new_[87083]_ ;
  assign \new_[495]_  = \new_[87070]_  & \new_[87055]_ ;
  assign \new_[496]_  = \new_[87042]_  & \new_[87027]_ ;
  assign \new_[497]_  = \new_[87014]_  & \new_[86999]_ ;
  assign \new_[498]_  = \new_[86986]_  & \new_[86971]_ ;
  assign \new_[499]_  = \new_[86958]_  & \new_[86943]_ ;
  assign \new_[500]_  = \new_[86930]_  & \new_[86915]_ ;
  assign \new_[501]_  = \new_[86902]_  & \new_[86887]_ ;
  assign \new_[502]_  = \new_[86874]_  & \new_[86859]_ ;
  assign \new_[503]_  = \new_[86846]_  & \new_[86831]_ ;
  assign \new_[504]_  = \new_[86818]_  & \new_[86803]_ ;
  assign \new_[505]_  = \new_[86790]_  & \new_[86777]_ ;
  assign \new_[506]_  = \new_[86764]_  & \new_[86751]_ ;
  assign \new_[507]_  = \new_[86738]_  & \new_[86725]_ ;
  assign \new_[508]_  = \new_[86712]_  & \new_[86699]_ ;
  assign \new_[509]_  = \new_[86686]_  & \new_[86673]_ ;
  assign \new_[510]_  = \new_[86660]_  & \new_[86647]_ ;
  assign \new_[511]_  = \new_[86634]_  & \new_[86621]_ ;
  assign \new_[512]_  = \new_[86608]_  & \new_[86595]_ ;
  assign \new_[513]_  = \new_[86582]_  & \new_[86569]_ ;
  assign \new_[514]_  = \new_[86556]_  & \new_[86543]_ ;
  assign \new_[515]_  = \new_[86530]_  & \new_[86517]_ ;
  assign \new_[516]_  = \new_[86504]_  & \new_[86491]_ ;
  assign \new_[517]_  = \new_[86478]_  & \new_[86465]_ ;
  assign \new_[518]_  = \new_[86452]_  & \new_[86439]_ ;
  assign \new_[519]_  = \new_[86426]_  & \new_[86413]_ ;
  assign \new_[520]_  = \new_[86400]_  & \new_[86387]_ ;
  assign \new_[521]_  = \new_[86374]_  & \new_[86361]_ ;
  assign \new_[522]_  = \new_[86348]_  & \new_[86335]_ ;
  assign \new_[523]_  = \new_[86322]_  & \new_[86309]_ ;
  assign \new_[524]_  = \new_[86296]_  & \new_[86283]_ ;
  assign \new_[525]_  = \new_[86270]_  & \new_[86257]_ ;
  assign \new_[526]_  = \new_[86244]_  & \new_[86231]_ ;
  assign \new_[527]_  = \new_[86218]_  & \new_[86205]_ ;
  assign \new_[528]_  = \new_[86192]_  & \new_[86179]_ ;
  assign \new_[529]_  = \new_[86166]_  & \new_[86153]_ ;
  assign \new_[530]_  = \new_[86140]_  & \new_[86127]_ ;
  assign \new_[531]_  = \new_[86114]_  & \new_[86101]_ ;
  assign \new_[532]_  = \new_[86088]_  & \new_[86075]_ ;
  assign \new_[533]_  = \new_[86062]_  & \new_[86049]_ ;
  assign \new_[534]_  = \new_[86036]_  & \new_[86023]_ ;
  assign \new_[535]_  = \new_[86010]_  & \new_[85997]_ ;
  assign \new_[536]_  = \new_[85984]_  & \new_[85971]_ ;
  assign \new_[537]_  = \new_[85958]_  & \new_[85945]_ ;
  assign \new_[538]_  = \new_[85932]_  & \new_[85919]_ ;
  assign \new_[539]_  = \new_[85906]_  & \new_[85893]_ ;
  assign \new_[540]_  = \new_[85880]_  & \new_[85867]_ ;
  assign \new_[541]_  = \new_[85854]_  & \new_[85841]_ ;
  assign \new_[542]_  = \new_[85828]_  & \new_[85815]_ ;
  assign \new_[543]_  = \new_[85802]_  & \new_[85789]_ ;
  assign \new_[544]_  = \new_[85776]_  & \new_[85763]_ ;
  assign \new_[545]_  = \new_[85750]_  & \new_[85737]_ ;
  assign \new_[546]_  = \new_[85724]_  & \new_[85711]_ ;
  assign \new_[547]_  = \new_[85698]_  & \new_[85685]_ ;
  assign \new_[548]_  = \new_[85672]_  & \new_[85659]_ ;
  assign \new_[549]_  = \new_[85646]_  & \new_[85633]_ ;
  assign \new_[550]_  = \new_[85620]_  & \new_[85607]_ ;
  assign \new_[551]_  = \new_[85594]_  & \new_[85581]_ ;
  assign \new_[552]_  = \new_[85568]_  & \new_[85555]_ ;
  assign \new_[553]_  = \new_[85542]_  & \new_[85529]_ ;
  assign \new_[554]_  = \new_[85516]_  & \new_[85503]_ ;
  assign \new_[555]_  = \new_[85490]_  & \new_[85477]_ ;
  assign \new_[556]_  = \new_[85464]_  & \new_[85451]_ ;
  assign \new_[557]_  = \new_[85438]_  & \new_[85425]_ ;
  assign \new_[558]_  = \new_[85412]_  & \new_[85399]_ ;
  assign \new_[559]_  = \new_[85386]_  & \new_[85373]_ ;
  assign \new_[560]_  = \new_[85360]_  & \new_[85347]_ ;
  assign \new_[561]_  = \new_[85334]_  & \new_[85321]_ ;
  assign \new_[562]_  = \new_[85308]_  & \new_[85295]_ ;
  assign \new_[563]_  = \new_[85282]_  & \new_[85269]_ ;
  assign \new_[564]_  = \new_[85256]_  & \new_[85243]_ ;
  assign \new_[565]_  = \new_[85230]_  & \new_[85217]_ ;
  assign \new_[566]_  = \new_[85204]_  & \new_[85191]_ ;
  assign \new_[567]_  = \new_[85178]_  & \new_[85165]_ ;
  assign \new_[568]_  = \new_[85152]_  & \new_[85139]_ ;
  assign \new_[569]_  = \new_[85126]_  & \new_[85113]_ ;
  assign \new_[570]_  = \new_[85100]_  & \new_[85087]_ ;
  assign \new_[571]_  = \new_[85074]_  & \new_[85061]_ ;
  assign \new_[572]_  = \new_[85048]_  & \new_[85035]_ ;
  assign \new_[573]_  = \new_[85022]_  & \new_[85009]_ ;
  assign \new_[574]_  = \new_[84996]_  & \new_[84983]_ ;
  assign \new_[575]_  = \new_[84970]_  & \new_[84957]_ ;
  assign \new_[576]_  = \new_[84944]_  & \new_[84931]_ ;
  assign \new_[577]_  = \new_[84918]_  & \new_[84905]_ ;
  assign \new_[578]_  = \new_[84892]_  & \new_[84879]_ ;
  assign \new_[579]_  = \new_[84866]_  & \new_[84853]_ ;
  assign \new_[580]_  = \new_[84840]_  & \new_[84827]_ ;
  assign \new_[581]_  = \new_[84814]_  & \new_[84801]_ ;
  assign \new_[582]_  = \new_[84788]_  & \new_[84775]_ ;
  assign \new_[583]_  = \new_[84762]_  & \new_[84749]_ ;
  assign \new_[584]_  = \new_[84736]_  & \new_[84723]_ ;
  assign \new_[585]_  = \new_[84710]_  & \new_[84697]_ ;
  assign \new_[586]_  = \new_[84684]_  & \new_[84671]_ ;
  assign \new_[587]_  = \new_[84658]_  & \new_[84645]_ ;
  assign \new_[588]_  = \new_[84632]_  & \new_[84619]_ ;
  assign \new_[589]_  = \new_[84606]_  & \new_[84593]_ ;
  assign \new_[590]_  = \new_[84580]_  & \new_[84567]_ ;
  assign \new_[591]_  = \new_[84554]_  & \new_[84541]_ ;
  assign \new_[592]_  = \new_[84528]_  & \new_[84515]_ ;
  assign \new_[593]_  = \new_[84502]_  & \new_[84489]_ ;
  assign \new_[594]_  = \new_[84476]_  & \new_[84463]_ ;
  assign \new_[595]_  = \new_[84450]_  & \new_[84437]_ ;
  assign \new_[596]_  = \new_[84424]_  & \new_[84411]_ ;
  assign \new_[597]_  = \new_[84398]_  & \new_[84385]_ ;
  assign \new_[598]_  = \new_[84372]_  & \new_[84359]_ ;
  assign \new_[599]_  = \new_[84346]_  & \new_[84333]_ ;
  assign \new_[600]_  = \new_[84320]_  & \new_[84307]_ ;
  assign \new_[601]_  = \new_[84294]_  & \new_[84281]_ ;
  assign \new_[602]_  = \new_[84268]_  & \new_[84255]_ ;
  assign \new_[603]_  = \new_[84242]_  & \new_[84229]_ ;
  assign \new_[604]_  = \new_[84216]_  & \new_[84203]_ ;
  assign \new_[605]_  = \new_[84190]_  & \new_[84177]_ ;
  assign \new_[606]_  = \new_[84164]_  & \new_[84151]_ ;
  assign \new_[607]_  = \new_[84138]_  & \new_[84125]_ ;
  assign \new_[608]_  = \new_[84112]_  & \new_[84099]_ ;
  assign \new_[609]_  = \new_[84086]_  & \new_[84073]_ ;
  assign \new_[610]_  = \new_[84060]_  & \new_[84047]_ ;
  assign \new_[611]_  = \new_[84034]_  & \new_[84021]_ ;
  assign \new_[612]_  = \new_[84008]_  & \new_[83995]_ ;
  assign \new_[613]_  = \new_[83982]_  & \new_[83969]_ ;
  assign \new_[614]_  = \new_[83956]_  & \new_[83943]_ ;
  assign \new_[615]_  = \new_[83930]_  & \new_[83917]_ ;
  assign \new_[616]_  = \new_[83904]_  & \new_[83891]_ ;
  assign \new_[617]_  = \new_[83878]_  & \new_[83865]_ ;
  assign \new_[618]_  = \new_[83852]_  & \new_[83839]_ ;
  assign \new_[619]_  = \new_[83826]_  & \new_[83813]_ ;
  assign \new_[620]_  = \new_[83800]_  & \new_[83787]_ ;
  assign \new_[621]_  = \new_[83774]_  & \new_[83761]_ ;
  assign \new_[622]_  = \new_[83748]_  & \new_[83735]_ ;
  assign \new_[623]_  = \new_[83722]_  & \new_[83709]_ ;
  assign \new_[624]_  = \new_[83696]_  & \new_[83683]_ ;
  assign \new_[625]_  = \new_[83670]_  & \new_[83657]_ ;
  assign \new_[626]_  = \new_[83644]_  & \new_[83631]_ ;
  assign \new_[627]_  = \new_[83618]_  & \new_[83605]_ ;
  assign \new_[628]_  = \new_[83592]_  & \new_[83579]_ ;
  assign \new_[629]_  = \new_[83566]_  & \new_[83553]_ ;
  assign \new_[630]_  = \new_[83540]_  & \new_[83527]_ ;
  assign \new_[631]_  = \new_[83514]_  & \new_[83501]_ ;
  assign \new_[632]_  = \new_[83488]_  & \new_[83475]_ ;
  assign \new_[633]_  = \new_[83462]_  & \new_[83449]_ ;
  assign \new_[634]_  = \new_[83436]_  & \new_[83423]_ ;
  assign \new_[635]_  = \new_[83410]_  & \new_[83397]_ ;
  assign \new_[636]_  = \new_[83384]_  & \new_[83371]_ ;
  assign \new_[637]_  = \new_[83358]_  & \new_[83345]_ ;
  assign \new_[638]_  = \new_[83332]_  & \new_[83319]_ ;
  assign \new_[639]_  = \new_[83306]_  & \new_[83293]_ ;
  assign \new_[640]_  = \new_[83280]_  & \new_[83267]_ ;
  assign \new_[641]_  = \new_[83254]_  & \new_[83241]_ ;
  assign \new_[642]_  = \new_[83228]_  & \new_[83215]_ ;
  assign \new_[643]_  = \new_[83202]_  & \new_[83189]_ ;
  assign \new_[644]_  = \new_[83176]_  & \new_[83163]_ ;
  assign \new_[645]_  = \new_[83150]_  & \new_[83137]_ ;
  assign \new_[646]_  = \new_[83124]_  & \new_[83111]_ ;
  assign \new_[647]_  = \new_[83098]_  & \new_[83085]_ ;
  assign \new_[648]_  = \new_[83072]_  & \new_[83059]_ ;
  assign \new_[649]_  = \new_[83046]_  & \new_[83033]_ ;
  assign \new_[650]_  = \new_[83020]_  & \new_[83007]_ ;
  assign \new_[651]_  = \new_[82994]_  & \new_[82981]_ ;
  assign \new_[652]_  = \new_[82968]_  & \new_[82955]_ ;
  assign \new_[653]_  = \new_[82942]_  & \new_[82929]_ ;
  assign \new_[654]_  = \new_[82916]_  & \new_[82903]_ ;
  assign \new_[655]_  = \new_[82890]_  & \new_[82877]_ ;
  assign \new_[656]_  = \new_[82864]_  & \new_[82851]_ ;
  assign \new_[657]_  = \new_[82838]_  & \new_[82825]_ ;
  assign \new_[658]_  = \new_[82812]_  & \new_[82799]_ ;
  assign \new_[659]_  = \new_[82786]_  & \new_[82773]_ ;
  assign \new_[660]_  = \new_[82760]_  & \new_[82747]_ ;
  assign \new_[661]_  = \new_[82734]_  & \new_[82721]_ ;
  assign \new_[662]_  = \new_[82708]_  & \new_[82695]_ ;
  assign \new_[663]_  = \new_[82682]_  & \new_[82669]_ ;
  assign \new_[664]_  = \new_[82656]_  & \new_[82643]_ ;
  assign \new_[665]_  = \new_[82630]_  & \new_[82617]_ ;
  assign \new_[666]_  = \new_[82604]_  & \new_[82591]_ ;
  assign \new_[667]_  = \new_[82578]_  & \new_[82565]_ ;
  assign \new_[668]_  = \new_[82552]_  & \new_[82539]_ ;
  assign \new_[669]_  = \new_[82526]_  & \new_[82513]_ ;
  assign \new_[670]_  = \new_[82500]_  & \new_[82487]_ ;
  assign \new_[671]_  = \new_[82474]_  & \new_[82461]_ ;
  assign \new_[672]_  = \new_[82448]_  & \new_[82435]_ ;
  assign \new_[673]_  = \new_[82422]_  & \new_[82409]_ ;
  assign \new_[674]_  = \new_[82396]_  & \new_[82383]_ ;
  assign \new_[675]_  = \new_[82370]_  & \new_[82357]_ ;
  assign \new_[676]_  = \new_[82344]_  & \new_[82331]_ ;
  assign \new_[677]_  = \new_[82318]_  & \new_[82305]_ ;
  assign \new_[678]_  = \new_[82292]_  & \new_[82279]_ ;
  assign \new_[679]_  = \new_[82266]_  & \new_[82253]_ ;
  assign \new_[680]_  = \new_[82240]_  & \new_[82227]_ ;
  assign \new_[681]_  = \new_[82214]_  & \new_[82201]_ ;
  assign \new_[682]_  = \new_[82188]_  & \new_[82175]_ ;
  assign \new_[683]_  = \new_[82162]_  & \new_[82149]_ ;
  assign \new_[684]_  = \new_[82136]_  & \new_[82123]_ ;
  assign \new_[685]_  = \new_[82110]_  & \new_[82097]_ ;
  assign \new_[686]_  = \new_[82084]_  & \new_[82071]_ ;
  assign \new_[687]_  = \new_[82058]_  & \new_[82045]_ ;
  assign \new_[688]_  = \new_[82032]_  & \new_[82019]_ ;
  assign \new_[689]_  = \new_[82006]_  & \new_[81993]_ ;
  assign \new_[690]_  = \new_[81980]_  & \new_[81967]_ ;
  assign \new_[691]_  = \new_[81954]_  & \new_[81941]_ ;
  assign \new_[692]_  = \new_[81928]_  & \new_[81915]_ ;
  assign \new_[693]_  = \new_[81902]_  & \new_[81889]_ ;
  assign \new_[694]_  = \new_[81876]_  & \new_[81863]_ ;
  assign \new_[695]_  = \new_[81850]_  & \new_[81837]_ ;
  assign \new_[696]_  = \new_[81824]_  & \new_[81811]_ ;
  assign \new_[697]_  = \new_[81798]_  & \new_[81785]_ ;
  assign \new_[698]_  = \new_[81772]_  & \new_[81759]_ ;
  assign \new_[699]_  = \new_[81746]_  & \new_[81733]_ ;
  assign \new_[700]_  = \new_[81720]_  & \new_[81707]_ ;
  assign \new_[701]_  = \new_[81694]_  & \new_[81681]_ ;
  assign \new_[702]_  = \new_[81668]_  & \new_[81655]_ ;
  assign \new_[703]_  = \new_[81642]_  & \new_[81629]_ ;
  assign \new_[704]_  = \new_[81616]_  & \new_[81603]_ ;
  assign \new_[705]_  = \new_[81590]_  & \new_[81577]_ ;
  assign \new_[706]_  = \new_[81564]_  & \new_[81551]_ ;
  assign \new_[707]_  = \new_[81538]_  & \new_[81525]_ ;
  assign \new_[708]_  = \new_[81512]_  & \new_[81499]_ ;
  assign \new_[709]_  = \new_[81486]_  & \new_[81473]_ ;
  assign \new_[710]_  = \new_[81460]_  & \new_[81447]_ ;
  assign \new_[711]_  = \new_[81434]_  & \new_[81421]_ ;
  assign \new_[712]_  = \new_[81408]_  & \new_[81395]_ ;
  assign \new_[713]_  = \new_[81382]_  & \new_[81369]_ ;
  assign \new_[714]_  = \new_[81356]_  & \new_[81343]_ ;
  assign \new_[715]_  = \new_[81330]_  & \new_[81317]_ ;
  assign \new_[716]_  = \new_[81304]_  & \new_[81291]_ ;
  assign \new_[717]_  = \new_[81278]_  & \new_[81265]_ ;
  assign \new_[718]_  = \new_[81252]_  & \new_[81239]_ ;
  assign \new_[719]_  = \new_[81226]_  & \new_[81213]_ ;
  assign \new_[720]_  = \new_[81200]_  & \new_[81187]_ ;
  assign \new_[721]_  = \new_[81174]_  & \new_[81161]_ ;
  assign \new_[722]_  = \new_[81148]_  & \new_[81135]_ ;
  assign \new_[723]_  = \new_[81122]_  & \new_[81109]_ ;
  assign \new_[724]_  = \new_[81096]_  & \new_[81083]_ ;
  assign \new_[725]_  = \new_[81070]_  & \new_[81057]_ ;
  assign \new_[726]_  = \new_[81044]_  & \new_[81031]_ ;
  assign \new_[727]_  = \new_[81018]_  & \new_[81005]_ ;
  assign \new_[728]_  = \new_[80992]_  & \new_[80979]_ ;
  assign \new_[729]_  = \new_[80966]_  & \new_[80953]_ ;
  assign \new_[730]_  = \new_[80940]_  & \new_[80927]_ ;
  assign \new_[731]_  = \new_[80914]_  & \new_[80901]_ ;
  assign \new_[732]_  = \new_[80888]_  & \new_[80875]_ ;
  assign \new_[733]_  = \new_[80862]_  & \new_[80849]_ ;
  assign \new_[734]_  = \new_[80836]_  & \new_[80823]_ ;
  assign \new_[735]_  = \new_[80810]_  & \new_[80797]_ ;
  assign \new_[736]_  = \new_[80784]_  & \new_[80771]_ ;
  assign \new_[737]_  = \new_[80758]_  & \new_[80745]_ ;
  assign \new_[738]_  = \new_[80732]_  & \new_[80719]_ ;
  assign \new_[739]_  = \new_[80706]_  & \new_[80693]_ ;
  assign \new_[740]_  = \new_[80680]_  & \new_[80667]_ ;
  assign \new_[741]_  = \new_[80654]_  & \new_[80641]_ ;
  assign \new_[742]_  = \new_[80628]_  & \new_[80615]_ ;
  assign \new_[743]_  = \new_[80602]_  & \new_[80589]_ ;
  assign \new_[744]_  = \new_[80576]_  & \new_[80563]_ ;
  assign \new_[745]_  = \new_[80550]_  & \new_[80537]_ ;
  assign \new_[746]_  = \new_[80524]_  & \new_[80511]_ ;
  assign \new_[747]_  = \new_[80498]_  & \new_[80485]_ ;
  assign \new_[748]_  = \new_[80472]_  & \new_[80459]_ ;
  assign \new_[749]_  = \new_[80446]_  & \new_[80433]_ ;
  assign \new_[750]_  = \new_[80420]_  & \new_[80407]_ ;
  assign \new_[751]_  = \new_[80394]_  & \new_[80381]_ ;
  assign \new_[752]_  = \new_[80368]_  & \new_[80355]_ ;
  assign \new_[753]_  = \new_[80342]_  & \new_[80329]_ ;
  assign \new_[754]_  = \new_[80316]_  & \new_[80303]_ ;
  assign \new_[755]_  = \new_[80290]_  & \new_[80277]_ ;
  assign \new_[756]_  = \new_[80264]_  & \new_[80251]_ ;
  assign \new_[757]_  = \new_[80238]_  & \new_[80225]_ ;
  assign \new_[758]_  = \new_[80212]_  & \new_[80199]_ ;
  assign \new_[759]_  = \new_[80186]_  & \new_[80173]_ ;
  assign \new_[760]_  = \new_[80160]_  & \new_[80147]_ ;
  assign \new_[761]_  = \new_[80134]_  & \new_[80121]_ ;
  assign \new_[762]_  = \new_[80108]_  & \new_[80095]_ ;
  assign \new_[763]_  = \new_[80082]_  & \new_[80069]_ ;
  assign \new_[764]_  = \new_[80056]_  & \new_[80043]_ ;
  assign \new_[765]_  = \new_[80030]_  & \new_[80017]_ ;
  assign \new_[766]_  = \new_[80004]_  & \new_[79991]_ ;
  assign \new_[767]_  = \new_[79978]_  & \new_[79965]_ ;
  assign \new_[768]_  = \new_[79952]_  & \new_[79939]_ ;
  assign \new_[769]_  = \new_[79926]_  & \new_[79913]_ ;
  assign \new_[770]_  = \new_[79900]_  & \new_[79887]_ ;
  assign \new_[771]_  = \new_[79874]_  & \new_[79861]_ ;
  assign \new_[772]_  = \new_[79848]_  & \new_[79835]_ ;
  assign \new_[773]_  = \new_[79822]_  & \new_[79809]_ ;
  assign \new_[774]_  = \new_[79796]_  & \new_[79783]_ ;
  assign \new_[775]_  = \new_[79770]_  & \new_[79757]_ ;
  assign \new_[776]_  = \new_[79744]_  & \new_[79731]_ ;
  assign \new_[777]_  = \new_[79718]_  & \new_[79705]_ ;
  assign \new_[778]_  = \new_[79692]_  & \new_[79679]_ ;
  assign \new_[779]_  = \new_[79666]_  & \new_[79653]_ ;
  assign \new_[780]_  = \new_[79640]_  & \new_[79627]_ ;
  assign \new_[781]_  = \new_[79614]_  & \new_[79601]_ ;
  assign \new_[782]_  = \new_[79588]_  & \new_[79575]_ ;
  assign \new_[783]_  = \new_[79562]_  & \new_[79549]_ ;
  assign \new_[784]_  = \new_[79536]_  & \new_[79523]_ ;
  assign \new_[785]_  = \new_[79510]_  & \new_[79497]_ ;
  assign \new_[786]_  = \new_[79484]_  & \new_[79471]_ ;
  assign \new_[787]_  = \new_[79458]_  & \new_[79445]_ ;
  assign \new_[788]_  = \new_[79432]_  & \new_[79419]_ ;
  assign \new_[789]_  = \new_[79406]_  & \new_[79393]_ ;
  assign \new_[790]_  = \new_[79380]_  & \new_[79367]_ ;
  assign \new_[791]_  = \new_[79354]_  & \new_[79341]_ ;
  assign \new_[792]_  = \new_[79328]_  & \new_[79315]_ ;
  assign \new_[793]_  = \new_[79302]_  & \new_[79289]_ ;
  assign \new_[794]_  = \new_[79276]_  & \new_[79263]_ ;
  assign \new_[795]_  = \new_[79250]_  & \new_[79237]_ ;
  assign \new_[796]_  = \new_[79224]_  & \new_[79211]_ ;
  assign \new_[797]_  = \new_[79198]_  & \new_[79185]_ ;
  assign \new_[798]_  = \new_[79172]_  & \new_[79159]_ ;
  assign \new_[799]_  = \new_[79146]_  & \new_[79133]_ ;
  assign \new_[800]_  = \new_[79120]_  & \new_[79107]_ ;
  assign \new_[801]_  = \new_[79094]_  & \new_[79081]_ ;
  assign \new_[802]_  = \new_[79068]_  & \new_[79055]_ ;
  assign \new_[803]_  = \new_[79042]_  & \new_[79029]_ ;
  assign \new_[804]_  = \new_[79016]_  & \new_[79003]_ ;
  assign \new_[805]_  = \new_[78990]_  & \new_[78977]_ ;
  assign \new_[806]_  = \new_[78964]_  & \new_[78951]_ ;
  assign \new_[807]_  = \new_[78938]_  & \new_[78925]_ ;
  assign \new_[808]_  = \new_[78912]_  & \new_[78899]_ ;
  assign \new_[809]_  = \new_[78886]_  & \new_[78873]_ ;
  assign \new_[810]_  = \new_[78860]_  & \new_[78847]_ ;
  assign \new_[811]_  = \new_[78834]_  & \new_[78821]_ ;
  assign \new_[812]_  = \new_[78808]_  & \new_[78795]_ ;
  assign \new_[813]_  = \new_[78782]_  & \new_[78769]_ ;
  assign \new_[814]_  = \new_[78756]_  & \new_[78743]_ ;
  assign \new_[815]_  = \new_[78730]_  & \new_[78717]_ ;
  assign \new_[816]_  = \new_[78704]_  & \new_[78691]_ ;
  assign \new_[817]_  = \new_[78678]_  & \new_[78665]_ ;
  assign \new_[818]_  = \new_[78652]_  & \new_[78639]_ ;
  assign \new_[819]_  = \new_[78626]_  & \new_[78613]_ ;
  assign \new_[820]_  = \new_[78600]_  & \new_[78587]_ ;
  assign \new_[821]_  = \new_[78574]_  & \new_[78561]_ ;
  assign \new_[822]_  = \new_[78548]_  & \new_[78535]_ ;
  assign \new_[823]_  = \new_[78522]_  & \new_[78509]_ ;
  assign \new_[824]_  = \new_[78496]_  & \new_[78483]_ ;
  assign \new_[825]_  = \new_[78470]_  & \new_[78457]_ ;
  assign \new_[826]_  = \new_[78444]_  & \new_[78431]_ ;
  assign \new_[827]_  = \new_[78418]_  & \new_[78405]_ ;
  assign \new_[828]_  = \new_[78392]_  & \new_[78379]_ ;
  assign \new_[829]_  = \new_[78366]_  & \new_[78353]_ ;
  assign \new_[830]_  = \new_[78340]_  & \new_[78327]_ ;
  assign \new_[831]_  = \new_[78314]_  & \new_[78301]_ ;
  assign \new_[832]_  = \new_[78288]_  & \new_[78275]_ ;
  assign \new_[833]_  = \new_[78262]_  & \new_[78249]_ ;
  assign \new_[834]_  = \new_[78236]_  & \new_[78223]_ ;
  assign \new_[835]_  = \new_[78210]_  & \new_[78197]_ ;
  assign \new_[836]_  = \new_[78184]_  & \new_[78171]_ ;
  assign \new_[837]_  = \new_[78158]_  & \new_[78145]_ ;
  assign \new_[838]_  = \new_[78132]_  & \new_[78119]_ ;
  assign \new_[839]_  = \new_[78106]_  & \new_[78093]_ ;
  assign \new_[840]_  = \new_[78080]_  & \new_[78067]_ ;
  assign \new_[841]_  = \new_[78054]_  & \new_[78041]_ ;
  assign \new_[842]_  = \new_[78028]_  & \new_[78015]_ ;
  assign \new_[843]_  = \new_[78002]_  & \new_[77989]_ ;
  assign \new_[844]_  = \new_[77976]_  & \new_[77963]_ ;
  assign \new_[845]_  = \new_[77950]_  & \new_[77937]_ ;
  assign \new_[846]_  = \new_[77924]_  & \new_[77911]_ ;
  assign \new_[847]_  = \new_[77898]_  & \new_[77885]_ ;
  assign \new_[848]_  = \new_[77872]_  & \new_[77859]_ ;
  assign \new_[849]_  = \new_[77846]_  & \new_[77833]_ ;
  assign \new_[850]_  = \new_[77820]_  & \new_[77807]_ ;
  assign \new_[851]_  = \new_[77794]_  & \new_[77781]_ ;
  assign \new_[852]_  = \new_[77768]_  & \new_[77755]_ ;
  assign \new_[853]_  = \new_[77742]_  & \new_[77729]_ ;
  assign \new_[854]_  = \new_[77716]_  & \new_[77703]_ ;
  assign \new_[855]_  = \new_[77690]_  & \new_[77677]_ ;
  assign \new_[856]_  = \new_[77664]_  & \new_[77651]_ ;
  assign \new_[857]_  = \new_[77638]_  & \new_[77625]_ ;
  assign \new_[858]_  = \new_[77612]_  & \new_[77599]_ ;
  assign \new_[859]_  = \new_[77586]_  & \new_[77573]_ ;
  assign \new_[860]_  = \new_[77560]_  & \new_[77547]_ ;
  assign \new_[861]_  = \new_[77534]_  & \new_[77521]_ ;
  assign \new_[862]_  = \new_[77508]_  & \new_[77495]_ ;
  assign \new_[863]_  = \new_[77482]_  & \new_[77469]_ ;
  assign \new_[864]_  = \new_[77456]_  & \new_[77443]_ ;
  assign \new_[865]_  = \new_[77430]_  & \new_[77417]_ ;
  assign \new_[866]_  = \new_[77404]_  & \new_[77391]_ ;
  assign \new_[867]_  = \new_[77378]_  & \new_[77365]_ ;
  assign \new_[868]_  = \new_[77352]_  & \new_[77339]_ ;
  assign \new_[869]_  = \new_[77326]_  & \new_[77313]_ ;
  assign \new_[870]_  = \new_[77300]_  & \new_[77287]_ ;
  assign \new_[871]_  = \new_[77274]_  & \new_[77261]_ ;
  assign \new_[872]_  = \new_[77248]_  & \new_[77235]_ ;
  assign \new_[873]_  = \new_[77222]_  & \new_[77209]_ ;
  assign \new_[874]_  = \new_[77196]_  & \new_[77183]_ ;
  assign \new_[875]_  = \new_[77170]_  & \new_[77157]_ ;
  assign \new_[876]_  = \new_[77144]_  & \new_[77131]_ ;
  assign \new_[877]_  = \new_[77118]_  & \new_[77105]_ ;
  assign \new_[878]_  = \new_[77092]_  & \new_[77079]_ ;
  assign \new_[879]_  = \new_[77066]_  & \new_[77053]_ ;
  assign \new_[880]_  = \new_[77040]_  & \new_[77027]_ ;
  assign \new_[881]_  = \new_[77014]_  & \new_[77001]_ ;
  assign \new_[882]_  = \new_[76988]_  & \new_[76975]_ ;
  assign \new_[883]_  = \new_[76962]_  & \new_[76949]_ ;
  assign \new_[884]_  = \new_[76936]_  & \new_[76923]_ ;
  assign \new_[885]_  = \new_[76910]_  & \new_[76897]_ ;
  assign \new_[886]_  = \new_[76884]_  & \new_[76871]_ ;
  assign \new_[887]_  = \new_[76858]_  & \new_[76845]_ ;
  assign \new_[888]_  = \new_[76832]_  & \new_[76819]_ ;
  assign \new_[889]_  = \new_[76806]_  & \new_[76793]_ ;
  assign \new_[890]_  = \new_[76780]_  & \new_[76767]_ ;
  assign \new_[891]_  = \new_[76754]_  & \new_[76741]_ ;
  assign \new_[892]_  = \new_[76728]_  & \new_[76715]_ ;
  assign \new_[893]_  = \new_[76702]_  & \new_[76689]_ ;
  assign \new_[894]_  = \new_[76676]_  & \new_[76663]_ ;
  assign \new_[895]_  = \new_[76650]_  & \new_[76637]_ ;
  assign \new_[896]_  = \new_[76624]_  & \new_[76611]_ ;
  assign \new_[897]_  = \new_[76598]_  & \new_[76585]_ ;
  assign \new_[898]_  = \new_[76572]_  & \new_[76559]_ ;
  assign \new_[899]_  = \new_[76546]_  & \new_[76533]_ ;
  assign \new_[900]_  = \new_[76520]_  & \new_[76507]_ ;
  assign \new_[901]_  = \new_[76494]_  & \new_[76481]_ ;
  assign \new_[902]_  = \new_[76468]_  & \new_[76455]_ ;
  assign \new_[903]_  = \new_[76442]_  & \new_[76429]_ ;
  assign \new_[904]_  = \new_[76416]_  & \new_[76403]_ ;
  assign \new_[905]_  = \new_[76390]_  & \new_[76377]_ ;
  assign \new_[906]_  = \new_[76364]_  & \new_[76351]_ ;
  assign \new_[907]_  = \new_[76338]_  & \new_[76325]_ ;
  assign \new_[908]_  = \new_[76312]_  & \new_[76299]_ ;
  assign \new_[909]_  = \new_[76286]_  & \new_[76273]_ ;
  assign \new_[910]_  = \new_[76260]_  & \new_[76247]_ ;
  assign \new_[911]_  = \new_[76234]_  & \new_[76221]_ ;
  assign \new_[912]_  = \new_[76208]_  & \new_[76195]_ ;
  assign \new_[913]_  = \new_[76182]_  & \new_[76169]_ ;
  assign \new_[914]_  = \new_[76156]_  & \new_[76143]_ ;
  assign \new_[915]_  = \new_[76130]_  & \new_[76117]_ ;
  assign \new_[916]_  = \new_[76104]_  & \new_[76091]_ ;
  assign \new_[917]_  = \new_[76078]_  & \new_[76065]_ ;
  assign \new_[918]_  = \new_[76052]_  & \new_[76039]_ ;
  assign \new_[919]_  = \new_[76026]_  & \new_[76013]_ ;
  assign \new_[920]_  = \new_[76000]_  & \new_[75987]_ ;
  assign \new_[921]_  = \new_[75974]_  & \new_[75961]_ ;
  assign \new_[922]_  = \new_[75948]_  & \new_[75935]_ ;
  assign \new_[923]_  = \new_[75922]_  & \new_[75909]_ ;
  assign \new_[924]_  = \new_[75896]_  & \new_[75883]_ ;
  assign \new_[925]_  = \new_[75870]_  & \new_[75857]_ ;
  assign \new_[926]_  = \new_[75844]_  & \new_[75831]_ ;
  assign \new_[927]_  = \new_[75818]_  & \new_[75805]_ ;
  assign \new_[928]_  = \new_[75792]_  & \new_[75779]_ ;
  assign \new_[929]_  = \new_[75766]_  & \new_[75753]_ ;
  assign \new_[930]_  = \new_[75740]_  & \new_[75727]_ ;
  assign \new_[931]_  = \new_[75714]_  & \new_[75701]_ ;
  assign \new_[932]_  = \new_[75688]_  & \new_[75675]_ ;
  assign \new_[933]_  = \new_[75662]_  & \new_[75649]_ ;
  assign \new_[934]_  = \new_[75636]_  & \new_[75623]_ ;
  assign \new_[935]_  = \new_[75610]_  & \new_[75597]_ ;
  assign \new_[936]_  = \new_[75584]_  & \new_[75571]_ ;
  assign \new_[937]_  = \new_[75558]_  & \new_[75545]_ ;
  assign \new_[938]_  = \new_[75532]_  & \new_[75519]_ ;
  assign \new_[939]_  = \new_[75506]_  & \new_[75493]_ ;
  assign \new_[940]_  = \new_[75480]_  & \new_[75467]_ ;
  assign \new_[941]_  = \new_[75454]_  & \new_[75441]_ ;
  assign \new_[942]_  = \new_[75428]_  & \new_[75415]_ ;
  assign \new_[943]_  = \new_[75402]_  & \new_[75389]_ ;
  assign \new_[944]_  = \new_[75376]_  & \new_[75363]_ ;
  assign \new_[945]_  = \new_[75350]_  & \new_[75337]_ ;
  assign \new_[946]_  = \new_[75324]_  & \new_[75311]_ ;
  assign \new_[947]_  = \new_[75298]_  & \new_[75285]_ ;
  assign \new_[948]_  = \new_[75272]_  & \new_[75259]_ ;
  assign \new_[949]_  = \new_[75246]_  & \new_[75233]_ ;
  assign \new_[950]_  = \new_[75220]_  & \new_[75207]_ ;
  assign \new_[951]_  = \new_[75194]_  & \new_[75181]_ ;
  assign \new_[952]_  = \new_[75168]_  & \new_[75155]_ ;
  assign \new_[953]_  = \new_[75142]_  & \new_[75129]_ ;
  assign \new_[954]_  = \new_[75116]_  & \new_[75103]_ ;
  assign \new_[955]_  = \new_[75090]_  & \new_[75077]_ ;
  assign \new_[956]_  = \new_[75064]_  & \new_[75051]_ ;
  assign \new_[957]_  = \new_[75038]_  & \new_[75025]_ ;
  assign \new_[958]_  = \new_[75012]_  & \new_[74999]_ ;
  assign \new_[959]_  = \new_[74986]_  & \new_[74973]_ ;
  assign \new_[960]_  = \new_[74960]_  & \new_[74947]_ ;
  assign \new_[961]_  = \new_[74934]_  & \new_[74921]_ ;
  assign \new_[962]_  = \new_[74908]_  & \new_[74895]_ ;
  assign \new_[963]_  = \new_[74882]_  & \new_[74869]_ ;
  assign \new_[964]_  = \new_[74856]_  & \new_[74843]_ ;
  assign \new_[965]_  = \new_[74830]_  & \new_[74817]_ ;
  assign \new_[966]_  = \new_[74804]_  & \new_[74791]_ ;
  assign \new_[967]_  = \new_[74778]_  & \new_[74765]_ ;
  assign \new_[968]_  = \new_[74752]_  & \new_[74739]_ ;
  assign \new_[969]_  = \new_[74726]_  & \new_[74713]_ ;
  assign \new_[970]_  = \new_[74700]_  & \new_[74687]_ ;
  assign \new_[971]_  = \new_[74674]_  & \new_[74661]_ ;
  assign \new_[972]_  = \new_[74648]_  & \new_[74635]_ ;
  assign \new_[973]_  = \new_[74622]_  & \new_[74609]_ ;
  assign \new_[974]_  = \new_[74596]_  & \new_[74583]_ ;
  assign \new_[975]_  = \new_[74570]_  & \new_[74557]_ ;
  assign \new_[976]_  = \new_[74544]_  & \new_[74531]_ ;
  assign \new_[977]_  = \new_[74518]_  & \new_[74505]_ ;
  assign \new_[978]_  = \new_[74492]_  & \new_[74479]_ ;
  assign \new_[979]_  = \new_[74466]_  & \new_[74453]_ ;
  assign \new_[980]_  = \new_[74440]_  & \new_[74427]_ ;
  assign \new_[981]_  = \new_[74414]_  & \new_[74401]_ ;
  assign \new_[982]_  = \new_[74388]_  & \new_[74375]_ ;
  assign \new_[983]_  = \new_[74362]_  & \new_[74349]_ ;
  assign \new_[984]_  = \new_[74336]_  & \new_[74323]_ ;
  assign \new_[985]_  = \new_[74310]_  & \new_[74297]_ ;
  assign \new_[986]_  = \new_[74284]_  & \new_[74271]_ ;
  assign \new_[987]_  = \new_[74258]_  & \new_[74245]_ ;
  assign \new_[988]_  = \new_[74232]_  & \new_[74219]_ ;
  assign \new_[989]_  = \new_[74206]_  & \new_[74193]_ ;
  assign \new_[990]_  = \new_[74180]_  & \new_[74167]_ ;
  assign \new_[991]_  = \new_[74154]_  & \new_[74141]_ ;
  assign \new_[992]_  = \new_[74128]_  & \new_[74115]_ ;
  assign \new_[993]_  = \new_[74102]_  & \new_[74089]_ ;
  assign \new_[994]_  = \new_[74076]_  & \new_[74063]_ ;
  assign \new_[995]_  = \new_[74050]_  & \new_[74037]_ ;
  assign \new_[996]_  = \new_[74024]_  & \new_[74011]_ ;
  assign \new_[997]_  = \new_[73998]_  & \new_[73985]_ ;
  assign \new_[998]_  = \new_[73972]_  & \new_[73959]_ ;
  assign \new_[999]_  = \new_[73946]_  & \new_[73933]_ ;
  assign \new_[1000]_  = \new_[73920]_  & \new_[73907]_ ;
  assign \new_[1001]_  = \new_[73894]_  & \new_[73881]_ ;
  assign \new_[1002]_  = \new_[73868]_  & \new_[73855]_ ;
  assign \new_[1003]_  = \new_[73842]_  & \new_[73829]_ ;
  assign \new_[1004]_  = \new_[73816]_  & \new_[73803]_ ;
  assign \new_[1005]_  = \new_[73790]_  & \new_[73777]_ ;
  assign \new_[1006]_  = \new_[73764]_  & \new_[73751]_ ;
  assign \new_[1007]_  = \new_[73738]_  & \new_[73725]_ ;
  assign \new_[1008]_  = \new_[73712]_  & \new_[73699]_ ;
  assign \new_[1009]_  = \new_[73686]_  & \new_[73673]_ ;
  assign \new_[1010]_  = \new_[73660]_  & \new_[73647]_ ;
  assign \new_[1011]_  = \new_[73634]_  & \new_[73621]_ ;
  assign \new_[1012]_  = \new_[73608]_  & \new_[73595]_ ;
  assign \new_[1013]_  = \new_[73582]_  & \new_[73569]_ ;
  assign \new_[1014]_  = \new_[73556]_  & \new_[73543]_ ;
  assign \new_[1015]_  = \new_[73530]_  & \new_[73517]_ ;
  assign \new_[1016]_  = \new_[73504]_  & \new_[73491]_ ;
  assign \new_[1017]_  = \new_[73478]_  & \new_[73465]_ ;
  assign \new_[1018]_  = \new_[73452]_  & \new_[73439]_ ;
  assign \new_[1019]_  = \new_[73426]_  & \new_[73413]_ ;
  assign \new_[1020]_  = \new_[73400]_  & \new_[73387]_ ;
  assign \new_[1021]_  = \new_[73374]_  & \new_[73361]_ ;
  assign \new_[1022]_  = \new_[73348]_  & \new_[73335]_ ;
  assign \new_[1023]_  = \new_[73322]_  & \new_[73309]_ ;
  assign \new_[1024]_  = \new_[73296]_  & \new_[73283]_ ;
  assign \new_[1025]_  = \new_[73270]_  & \new_[73257]_ ;
  assign \new_[1026]_  = \new_[73244]_  & \new_[73231]_ ;
  assign \new_[1027]_  = \new_[73218]_  & \new_[73205]_ ;
  assign \new_[1028]_  = \new_[73192]_  & \new_[73179]_ ;
  assign \new_[1029]_  = \new_[73166]_  & \new_[73153]_ ;
  assign \new_[1030]_  = \new_[73140]_  & \new_[73127]_ ;
  assign \new_[1031]_  = \new_[73114]_  & \new_[73101]_ ;
  assign \new_[1032]_  = \new_[73088]_  & \new_[73075]_ ;
  assign \new_[1033]_  = \new_[73062]_  & \new_[73049]_ ;
  assign \new_[1034]_  = \new_[73036]_  & \new_[73023]_ ;
  assign \new_[1035]_  = \new_[73010]_  & \new_[72997]_ ;
  assign \new_[1036]_  = \new_[72984]_  & \new_[72971]_ ;
  assign \new_[1037]_  = \new_[72958]_  & \new_[72945]_ ;
  assign \new_[1038]_  = \new_[72932]_  & \new_[72919]_ ;
  assign \new_[1039]_  = \new_[72906]_  & \new_[72893]_ ;
  assign \new_[1040]_  = \new_[72880]_  & \new_[72867]_ ;
  assign \new_[1041]_  = \new_[72854]_  & \new_[72841]_ ;
  assign \new_[1042]_  = \new_[72828]_  & \new_[72815]_ ;
  assign \new_[1043]_  = \new_[72802]_  & \new_[72789]_ ;
  assign \new_[1044]_  = \new_[72776]_  & \new_[72763]_ ;
  assign \new_[1045]_  = \new_[72750]_  & \new_[72737]_ ;
  assign \new_[1046]_  = \new_[72724]_  & \new_[72711]_ ;
  assign \new_[1047]_  = \new_[72698]_  & \new_[72685]_ ;
  assign \new_[1048]_  = \new_[72672]_  & \new_[72659]_ ;
  assign \new_[1049]_  = \new_[72646]_  & \new_[72633]_ ;
  assign \new_[1050]_  = \new_[72620]_  & \new_[72607]_ ;
  assign \new_[1051]_  = \new_[72594]_  & \new_[72581]_ ;
  assign \new_[1052]_  = \new_[72568]_  & \new_[72555]_ ;
  assign \new_[1053]_  = \new_[72542]_  & \new_[72529]_ ;
  assign \new_[1054]_  = \new_[72516]_  & \new_[72503]_ ;
  assign \new_[1055]_  = \new_[72490]_  & \new_[72477]_ ;
  assign \new_[1056]_  = \new_[72464]_  & \new_[72451]_ ;
  assign \new_[1057]_  = \new_[72438]_  & \new_[72425]_ ;
  assign \new_[1058]_  = \new_[72412]_  & \new_[72399]_ ;
  assign \new_[1059]_  = \new_[72386]_  & \new_[72373]_ ;
  assign \new_[1060]_  = \new_[72360]_  & \new_[72347]_ ;
  assign \new_[1061]_  = \new_[72334]_  & \new_[72321]_ ;
  assign \new_[1062]_  = \new_[72308]_  & \new_[72295]_ ;
  assign \new_[1063]_  = \new_[72282]_  & \new_[72269]_ ;
  assign \new_[1064]_  = \new_[72256]_  & \new_[72243]_ ;
  assign \new_[1065]_  = \new_[72230]_  & \new_[72217]_ ;
  assign \new_[1066]_  = \new_[72204]_  & \new_[72191]_ ;
  assign \new_[1067]_  = \new_[72178]_  & \new_[72165]_ ;
  assign \new_[1068]_  = \new_[72152]_  & \new_[72139]_ ;
  assign \new_[1069]_  = \new_[72126]_  & \new_[72113]_ ;
  assign \new_[1070]_  = \new_[72100]_  & \new_[72087]_ ;
  assign \new_[1071]_  = \new_[72074]_  & \new_[72061]_ ;
  assign \new_[1072]_  = \new_[72048]_  & \new_[72035]_ ;
  assign \new_[1073]_  = \new_[72022]_  & \new_[72009]_ ;
  assign \new_[1074]_  = \new_[71996]_  & \new_[71983]_ ;
  assign \new_[1075]_  = \new_[71970]_  & \new_[71957]_ ;
  assign \new_[1076]_  = \new_[71944]_  & \new_[71931]_ ;
  assign \new_[1077]_  = \new_[71918]_  & \new_[71905]_ ;
  assign \new_[1078]_  = \new_[71892]_  & \new_[71879]_ ;
  assign \new_[1079]_  = \new_[71866]_  & \new_[71853]_ ;
  assign \new_[1080]_  = \new_[71840]_  & \new_[71827]_ ;
  assign \new_[1081]_  = \new_[71814]_  & \new_[71801]_ ;
  assign \new_[1082]_  = \new_[71788]_  & \new_[71775]_ ;
  assign \new_[1083]_  = \new_[71762]_  & \new_[71749]_ ;
  assign \new_[1084]_  = \new_[71736]_  & \new_[71723]_ ;
  assign \new_[1085]_  = \new_[71710]_  & \new_[71697]_ ;
  assign \new_[1086]_  = \new_[71684]_  & \new_[71671]_ ;
  assign \new_[1087]_  = \new_[71658]_  & \new_[71645]_ ;
  assign \new_[1088]_  = \new_[71632]_  & \new_[71619]_ ;
  assign \new_[1089]_  = \new_[71606]_  & \new_[71593]_ ;
  assign \new_[1090]_  = \new_[71580]_  & \new_[71567]_ ;
  assign \new_[1091]_  = \new_[71554]_  & \new_[71541]_ ;
  assign \new_[1092]_  = \new_[71528]_  & \new_[71515]_ ;
  assign \new_[1093]_  = \new_[71502]_  & \new_[71489]_ ;
  assign \new_[1094]_  = \new_[71476]_  & \new_[71463]_ ;
  assign \new_[1095]_  = \new_[71450]_  & \new_[71437]_ ;
  assign \new_[1096]_  = \new_[71424]_  & \new_[71411]_ ;
  assign \new_[1097]_  = \new_[71398]_  & \new_[71385]_ ;
  assign \new_[1098]_  = \new_[71372]_  & \new_[71359]_ ;
  assign \new_[1099]_  = \new_[71346]_  & \new_[71333]_ ;
  assign \new_[1100]_  = \new_[71320]_  & \new_[71307]_ ;
  assign \new_[1101]_  = \new_[71294]_  & \new_[71281]_ ;
  assign \new_[1102]_  = \new_[71268]_  & \new_[71255]_ ;
  assign \new_[1103]_  = \new_[71242]_  & \new_[71229]_ ;
  assign \new_[1104]_  = \new_[71216]_  & \new_[71203]_ ;
  assign \new_[1105]_  = \new_[71190]_  & \new_[71177]_ ;
  assign \new_[1106]_  = \new_[71164]_  & \new_[71151]_ ;
  assign \new_[1107]_  = \new_[71138]_  & \new_[71125]_ ;
  assign \new_[1108]_  = \new_[71112]_  & \new_[71099]_ ;
  assign \new_[1109]_  = \new_[71086]_  & \new_[71073]_ ;
  assign \new_[1110]_  = \new_[71060]_  & \new_[71047]_ ;
  assign \new_[1111]_  = \new_[71034]_  & \new_[71021]_ ;
  assign \new_[1112]_  = \new_[71008]_  & \new_[70995]_ ;
  assign \new_[1113]_  = \new_[70982]_  & \new_[70969]_ ;
  assign \new_[1114]_  = \new_[70956]_  & \new_[70943]_ ;
  assign \new_[1115]_  = \new_[70930]_  & \new_[70917]_ ;
  assign \new_[1116]_  = \new_[70904]_  & \new_[70891]_ ;
  assign \new_[1117]_  = \new_[70878]_  & \new_[70865]_ ;
  assign \new_[1118]_  = \new_[70852]_  & \new_[70839]_ ;
  assign \new_[1119]_  = \new_[70826]_  & \new_[70813]_ ;
  assign \new_[1120]_  = \new_[70800]_  & \new_[70787]_ ;
  assign \new_[1121]_  = \new_[70774]_  & \new_[70761]_ ;
  assign \new_[1122]_  = \new_[70748]_  & \new_[70735]_ ;
  assign \new_[1123]_  = \new_[70722]_  & \new_[70709]_ ;
  assign \new_[1124]_  = \new_[70696]_  & \new_[70683]_ ;
  assign \new_[1125]_  = \new_[70670]_  & \new_[70657]_ ;
  assign \new_[1126]_  = \new_[70644]_  & \new_[70631]_ ;
  assign \new_[1127]_  = \new_[70618]_  & \new_[70605]_ ;
  assign \new_[1128]_  = \new_[70592]_  & \new_[70579]_ ;
  assign \new_[1129]_  = \new_[70566]_  & \new_[70553]_ ;
  assign \new_[1130]_  = \new_[70540]_  & \new_[70527]_ ;
  assign \new_[1131]_  = \new_[70514]_  & \new_[70501]_ ;
  assign \new_[1132]_  = \new_[70488]_  & \new_[70475]_ ;
  assign \new_[1133]_  = \new_[70462]_  & \new_[70449]_ ;
  assign \new_[1134]_  = \new_[70436]_  & \new_[70423]_ ;
  assign \new_[1135]_  = \new_[70410]_  & \new_[70397]_ ;
  assign \new_[1136]_  = \new_[70384]_  & \new_[70371]_ ;
  assign \new_[1137]_  = \new_[70358]_  & \new_[70345]_ ;
  assign \new_[1138]_  = \new_[70332]_  & \new_[70319]_ ;
  assign \new_[1139]_  = \new_[70306]_  & \new_[70293]_ ;
  assign \new_[1140]_  = \new_[70280]_  & \new_[70267]_ ;
  assign \new_[1141]_  = \new_[70254]_  & \new_[70241]_ ;
  assign \new_[1142]_  = \new_[70228]_  & \new_[70215]_ ;
  assign \new_[1143]_  = \new_[70202]_  & \new_[70189]_ ;
  assign \new_[1144]_  = \new_[70176]_  & \new_[70163]_ ;
  assign \new_[1145]_  = \new_[70150]_  & \new_[70137]_ ;
  assign \new_[1146]_  = \new_[70124]_  & \new_[70111]_ ;
  assign \new_[1147]_  = \new_[70098]_  & \new_[70085]_ ;
  assign \new_[1148]_  = \new_[70072]_  & \new_[70059]_ ;
  assign \new_[1149]_  = \new_[70046]_  & \new_[70033]_ ;
  assign \new_[1150]_  = \new_[70020]_  & \new_[70007]_ ;
  assign \new_[1151]_  = \new_[69994]_  & \new_[69981]_ ;
  assign \new_[1152]_  = \new_[69968]_  & \new_[69955]_ ;
  assign \new_[1153]_  = \new_[69942]_  & \new_[69929]_ ;
  assign \new_[1154]_  = \new_[69916]_  & \new_[69903]_ ;
  assign \new_[1155]_  = \new_[69890]_  & \new_[69877]_ ;
  assign \new_[1156]_  = \new_[69864]_  & \new_[69851]_ ;
  assign \new_[1157]_  = \new_[69838]_  & \new_[69825]_ ;
  assign \new_[1158]_  = \new_[69812]_  & \new_[69799]_ ;
  assign \new_[1159]_  = \new_[69786]_  & \new_[69773]_ ;
  assign \new_[1160]_  = \new_[69760]_  & \new_[69747]_ ;
  assign \new_[1161]_  = \new_[69734]_  & \new_[69721]_ ;
  assign \new_[1162]_  = \new_[69708]_  & \new_[69695]_ ;
  assign \new_[1163]_  = \new_[69682]_  & \new_[69669]_ ;
  assign \new_[1164]_  = \new_[69656]_  & \new_[69643]_ ;
  assign \new_[1165]_  = \new_[69630]_  & \new_[69617]_ ;
  assign \new_[1166]_  = \new_[69604]_  & \new_[69591]_ ;
  assign \new_[1167]_  = \new_[69578]_  & \new_[69565]_ ;
  assign \new_[1168]_  = \new_[69552]_  & \new_[69539]_ ;
  assign \new_[1169]_  = \new_[69526]_  & \new_[69513]_ ;
  assign \new_[1170]_  = \new_[69500]_  & \new_[69487]_ ;
  assign \new_[1171]_  = \new_[69474]_  & \new_[69461]_ ;
  assign \new_[1172]_  = \new_[69448]_  & \new_[69435]_ ;
  assign \new_[1173]_  = \new_[69422]_  & \new_[69409]_ ;
  assign \new_[1174]_  = \new_[69396]_  & \new_[69383]_ ;
  assign \new_[1175]_  = \new_[69370]_  & \new_[69357]_ ;
  assign \new_[1176]_  = \new_[69344]_  & \new_[69331]_ ;
  assign \new_[1177]_  = \new_[69318]_  & \new_[69305]_ ;
  assign \new_[1178]_  = \new_[69292]_  & \new_[69279]_ ;
  assign \new_[1179]_  = \new_[69266]_  & \new_[69253]_ ;
  assign \new_[1180]_  = \new_[69240]_  & \new_[69227]_ ;
  assign \new_[1181]_  = \new_[69214]_  & \new_[69201]_ ;
  assign \new_[1182]_  = \new_[69188]_  & \new_[69175]_ ;
  assign \new_[1183]_  = \new_[69162]_  & \new_[69149]_ ;
  assign \new_[1184]_  = \new_[69136]_  & \new_[69123]_ ;
  assign \new_[1185]_  = \new_[69110]_  & \new_[69097]_ ;
  assign \new_[1186]_  = \new_[69084]_  & \new_[69071]_ ;
  assign \new_[1187]_  = \new_[69058]_  & \new_[69045]_ ;
  assign \new_[1188]_  = \new_[69032]_  & \new_[69019]_ ;
  assign \new_[1189]_  = \new_[69006]_  & \new_[68993]_ ;
  assign \new_[1190]_  = \new_[68980]_  & \new_[68967]_ ;
  assign \new_[1191]_  = \new_[68954]_  & \new_[68941]_ ;
  assign \new_[1192]_  = \new_[68928]_  & \new_[68915]_ ;
  assign \new_[1193]_  = \new_[68902]_  & \new_[68889]_ ;
  assign \new_[1194]_  = \new_[68876]_  & \new_[68863]_ ;
  assign \new_[1195]_  = \new_[68850]_  & \new_[68837]_ ;
  assign \new_[1196]_  = \new_[68824]_  & \new_[68811]_ ;
  assign \new_[1197]_  = \new_[68798]_  & \new_[68785]_ ;
  assign \new_[1198]_  = \new_[68772]_  & \new_[68759]_ ;
  assign \new_[1199]_  = \new_[68746]_  & \new_[68733]_ ;
  assign \new_[1200]_  = \new_[68720]_  & \new_[68707]_ ;
  assign \new_[1201]_  = \new_[68694]_  & \new_[68681]_ ;
  assign \new_[1202]_  = \new_[68668]_  & \new_[68655]_ ;
  assign \new_[1203]_  = \new_[68642]_  & \new_[68629]_ ;
  assign \new_[1204]_  = \new_[68616]_  & \new_[68603]_ ;
  assign \new_[1205]_  = \new_[68590]_  & \new_[68577]_ ;
  assign \new_[1206]_  = \new_[68564]_  & \new_[68551]_ ;
  assign \new_[1207]_  = \new_[68538]_  & \new_[68525]_ ;
  assign \new_[1208]_  = \new_[68512]_  & \new_[68499]_ ;
  assign \new_[1209]_  = \new_[68486]_  & \new_[68473]_ ;
  assign \new_[1210]_  = \new_[68460]_  & \new_[68447]_ ;
  assign \new_[1211]_  = \new_[68434]_  & \new_[68421]_ ;
  assign \new_[1212]_  = \new_[68408]_  & \new_[68395]_ ;
  assign \new_[1213]_  = \new_[68382]_  & \new_[68369]_ ;
  assign \new_[1214]_  = \new_[68356]_  & \new_[68343]_ ;
  assign \new_[1215]_  = \new_[68330]_  & \new_[68317]_ ;
  assign \new_[1216]_  = \new_[68304]_  & \new_[68291]_ ;
  assign \new_[1217]_  = \new_[68278]_  & \new_[68265]_ ;
  assign \new_[1218]_  = \new_[68252]_  & \new_[68239]_ ;
  assign \new_[1219]_  = \new_[68226]_  & \new_[68213]_ ;
  assign \new_[1220]_  = \new_[68200]_  & \new_[68187]_ ;
  assign \new_[1221]_  = \new_[68174]_  & \new_[68161]_ ;
  assign \new_[1222]_  = \new_[68148]_  & \new_[68135]_ ;
  assign \new_[1223]_  = \new_[68122]_  & \new_[68109]_ ;
  assign \new_[1224]_  = \new_[68096]_  & \new_[68083]_ ;
  assign \new_[1225]_  = \new_[68070]_  & \new_[68057]_ ;
  assign \new_[1226]_  = \new_[68044]_  & \new_[68031]_ ;
  assign \new_[1227]_  = \new_[68018]_  & \new_[68005]_ ;
  assign \new_[1228]_  = \new_[67992]_  & \new_[67979]_ ;
  assign \new_[1229]_  = \new_[67966]_  & \new_[67953]_ ;
  assign \new_[1230]_  = \new_[67940]_  & \new_[67927]_ ;
  assign \new_[1231]_  = \new_[67914]_  & \new_[67901]_ ;
  assign \new_[1232]_  = \new_[67888]_  & \new_[67875]_ ;
  assign \new_[1233]_  = \new_[67862]_  & \new_[67849]_ ;
  assign \new_[1234]_  = \new_[67836]_  & \new_[67823]_ ;
  assign \new_[1235]_  = \new_[67810]_  & \new_[67797]_ ;
  assign \new_[1236]_  = \new_[67784]_  & \new_[67771]_ ;
  assign \new_[1237]_  = \new_[67758]_  & \new_[67745]_ ;
  assign \new_[1238]_  = \new_[67732]_  & \new_[67719]_ ;
  assign \new_[1239]_  = \new_[67706]_  & \new_[67693]_ ;
  assign \new_[1240]_  = \new_[67680]_  & \new_[67667]_ ;
  assign \new_[1241]_  = \new_[67654]_  & \new_[67641]_ ;
  assign \new_[1242]_  = \new_[67628]_  & \new_[67615]_ ;
  assign \new_[1243]_  = \new_[67602]_  & \new_[67589]_ ;
  assign \new_[1244]_  = \new_[67576]_  & \new_[67563]_ ;
  assign \new_[1245]_  = \new_[67550]_  & \new_[67537]_ ;
  assign \new_[1246]_  = \new_[67524]_  & \new_[67511]_ ;
  assign \new_[1247]_  = \new_[67498]_  & \new_[67485]_ ;
  assign \new_[1248]_  = \new_[67472]_  & \new_[67459]_ ;
  assign \new_[1249]_  = \new_[67446]_  & \new_[67433]_ ;
  assign \new_[1250]_  = \new_[67420]_  & \new_[67407]_ ;
  assign \new_[1251]_  = \new_[67394]_  & \new_[67381]_ ;
  assign \new_[1252]_  = \new_[67368]_  & \new_[67355]_ ;
  assign \new_[1253]_  = \new_[67342]_  & \new_[67329]_ ;
  assign \new_[1254]_  = \new_[67316]_  & \new_[67303]_ ;
  assign \new_[1255]_  = \new_[67290]_  & \new_[67277]_ ;
  assign \new_[1256]_  = \new_[67264]_  & \new_[67251]_ ;
  assign \new_[1257]_  = \new_[67238]_  & \new_[67225]_ ;
  assign \new_[1258]_  = \new_[67212]_  & \new_[67199]_ ;
  assign \new_[1259]_  = \new_[67186]_  & \new_[67173]_ ;
  assign \new_[1260]_  = \new_[67160]_  & \new_[67147]_ ;
  assign \new_[1261]_  = \new_[67134]_  & \new_[67121]_ ;
  assign \new_[1262]_  = \new_[67108]_  & \new_[67095]_ ;
  assign \new_[1263]_  = \new_[67082]_  & \new_[67069]_ ;
  assign \new_[1264]_  = \new_[67056]_  & \new_[67043]_ ;
  assign \new_[1265]_  = \new_[67030]_  & \new_[67017]_ ;
  assign \new_[1266]_  = \new_[67004]_  & \new_[66991]_ ;
  assign \new_[1267]_  = \new_[66978]_  & \new_[66965]_ ;
  assign \new_[1268]_  = \new_[66952]_  & \new_[66939]_ ;
  assign \new_[1269]_  = \new_[66926]_  & \new_[66913]_ ;
  assign \new_[1270]_  = \new_[66900]_  & \new_[66887]_ ;
  assign \new_[1271]_  = \new_[66874]_  & \new_[66861]_ ;
  assign \new_[1272]_  = \new_[66848]_  & \new_[66835]_ ;
  assign \new_[1273]_  = \new_[66822]_  & \new_[66809]_ ;
  assign \new_[1274]_  = \new_[66796]_  & \new_[66783]_ ;
  assign \new_[1275]_  = \new_[66770]_  & \new_[66757]_ ;
  assign \new_[1276]_  = \new_[66744]_  & \new_[66731]_ ;
  assign \new_[1277]_  = \new_[66718]_  & \new_[66705]_ ;
  assign \new_[1278]_  = \new_[66692]_  & \new_[66679]_ ;
  assign \new_[1279]_  = \new_[66666]_  & \new_[66653]_ ;
  assign \new_[1280]_  = \new_[66640]_  & \new_[66627]_ ;
  assign \new_[1281]_  = \new_[66614]_  & \new_[66601]_ ;
  assign \new_[1282]_  = \new_[66588]_  & \new_[66575]_ ;
  assign \new_[1283]_  = \new_[66562]_  & \new_[66549]_ ;
  assign \new_[1284]_  = \new_[66536]_  & \new_[66523]_ ;
  assign \new_[1285]_  = \new_[66510]_  & \new_[66497]_ ;
  assign \new_[1286]_  = \new_[66484]_  & \new_[66471]_ ;
  assign \new_[1287]_  = \new_[66458]_  & \new_[66445]_ ;
  assign \new_[1288]_  = \new_[66432]_  & \new_[66419]_ ;
  assign \new_[1289]_  = \new_[66406]_  & \new_[66393]_ ;
  assign \new_[1290]_  = \new_[66380]_  & \new_[66367]_ ;
  assign \new_[1291]_  = \new_[66354]_  & \new_[66341]_ ;
  assign \new_[1292]_  = \new_[66328]_  & \new_[66315]_ ;
  assign \new_[1293]_  = \new_[66302]_  & \new_[66289]_ ;
  assign \new_[1294]_  = \new_[66276]_  & \new_[66263]_ ;
  assign \new_[1295]_  = \new_[66250]_  & \new_[66237]_ ;
  assign \new_[1296]_  = \new_[66224]_  & \new_[66211]_ ;
  assign \new_[1297]_  = \new_[66198]_  & \new_[66185]_ ;
  assign \new_[1298]_  = \new_[66172]_  & \new_[66159]_ ;
  assign \new_[1299]_  = \new_[66146]_  & \new_[66133]_ ;
  assign \new_[1300]_  = \new_[66120]_  & \new_[66107]_ ;
  assign \new_[1301]_  = \new_[66094]_  & \new_[66081]_ ;
  assign \new_[1302]_  = \new_[66068]_  & \new_[66055]_ ;
  assign \new_[1303]_  = \new_[66042]_  & \new_[66029]_ ;
  assign \new_[1304]_  = \new_[66016]_  & \new_[66003]_ ;
  assign \new_[1305]_  = \new_[65990]_  & \new_[65977]_ ;
  assign \new_[1306]_  = \new_[65964]_  & \new_[65951]_ ;
  assign \new_[1307]_  = \new_[65938]_  & \new_[65925]_ ;
  assign \new_[1308]_  = \new_[65912]_  & \new_[65899]_ ;
  assign \new_[1309]_  = \new_[65886]_  & \new_[65873]_ ;
  assign \new_[1310]_  = \new_[65860]_  & \new_[65847]_ ;
  assign \new_[1311]_  = \new_[65834]_  & \new_[65821]_ ;
  assign \new_[1312]_  = \new_[65808]_  & \new_[65795]_ ;
  assign \new_[1313]_  = \new_[65782]_  & \new_[65769]_ ;
  assign \new_[1314]_  = \new_[65756]_  & \new_[65743]_ ;
  assign \new_[1315]_  = \new_[65730]_  & \new_[65717]_ ;
  assign \new_[1316]_  = \new_[65704]_  & \new_[65691]_ ;
  assign \new_[1317]_  = \new_[65678]_  & \new_[65665]_ ;
  assign \new_[1318]_  = \new_[65652]_  & \new_[65639]_ ;
  assign \new_[1319]_  = \new_[65626]_  & \new_[65613]_ ;
  assign \new_[1320]_  = \new_[65600]_  & \new_[65587]_ ;
  assign \new_[1321]_  = \new_[65574]_  & \new_[65561]_ ;
  assign \new_[1322]_  = \new_[65548]_  & \new_[65535]_ ;
  assign \new_[1323]_  = \new_[65522]_  & \new_[65509]_ ;
  assign \new_[1324]_  = \new_[65496]_  & \new_[65483]_ ;
  assign \new_[1325]_  = \new_[65470]_  & \new_[65457]_ ;
  assign \new_[1326]_  = \new_[65444]_  & \new_[65431]_ ;
  assign \new_[1327]_  = \new_[65418]_  & \new_[65405]_ ;
  assign \new_[1328]_  = \new_[65392]_  & \new_[65379]_ ;
  assign \new_[1329]_  = \new_[65366]_  & \new_[65353]_ ;
  assign \new_[1330]_  = \new_[65340]_  & \new_[65327]_ ;
  assign \new_[1331]_  = \new_[65314]_  & \new_[65301]_ ;
  assign \new_[1332]_  = \new_[65288]_  & \new_[65275]_ ;
  assign \new_[1333]_  = \new_[65262]_  & \new_[65249]_ ;
  assign \new_[1334]_  = \new_[65236]_  & \new_[65223]_ ;
  assign \new_[1335]_  = \new_[65210]_  & \new_[65197]_ ;
  assign \new_[1336]_  = \new_[65184]_  & \new_[65171]_ ;
  assign \new_[1337]_  = \new_[65158]_  & \new_[65145]_ ;
  assign \new_[1338]_  = \new_[65132]_  & \new_[65119]_ ;
  assign \new_[1339]_  = \new_[65106]_  & \new_[65093]_ ;
  assign \new_[1340]_  = \new_[65080]_  & \new_[65067]_ ;
  assign \new_[1341]_  = \new_[65054]_  & \new_[65041]_ ;
  assign \new_[1342]_  = \new_[65028]_  & \new_[65015]_ ;
  assign \new_[1343]_  = \new_[65002]_  & \new_[64989]_ ;
  assign \new_[1344]_  = \new_[64976]_  & \new_[64963]_ ;
  assign \new_[1345]_  = \new_[64950]_  & \new_[64937]_ ;
  assign \new_[1346]_  = \new_[64924]_  & \new_[64911]_ ;
  assign \new_[1347]_  = \new_[64898]_  & \new_[64885]_ ;
  assign \new_[1348]_  = \new_[64872]_  & \new_[64859]_ ;
  assign \new_[1349]_  = \new_[64846]_  & \new_[64833]_ ;
  assign \new_[1350]_  = \new_[64820]_  & \new_[64807]_ ;
  assign \new_[1351]_  = \new_[64794]_  & \new_[64781]_ ;
  assign \new_[1352]_  = \new_[64768]_  & \new_[64755]_ ;
  assign \new_[1353]_  = \new_[64742]_  & \new_[64729]_ ;
  assign \new_[1354]_  = \new_[64716]_  & \new_[64703]_ ;
  assign \new_[1355]_  = \new_[64690]_  & \new_[64677]_ ;
  assign \new_[1356]_  = \new_[64664]_  & \new_[64651]_ ;
  assign \new_[1357]_  = \new_[64638]_  & \new_[64625]_ ;
  assign \new_[1358]_  = \new_[64614]_  & \new_[64601]_ ;
  assign \new_[1359]_  = \new_[64590]_  & \new_[64577]_ ;
  assign \new_[1360]_  = \new_[64566]_  & \new_[64553]_ ;
  assign \new_[1361]_  = \new_[64542]_  & \new_[64529]_ ;
  assign \new_[1362]_  = \new_[64518]_  & \new_[64505]_ ;
  assign \new_[1363]_  = \new_[64494]_  & \new_[64481]_ ;
  assign \new_[1364]_  = \new_[64470]_  & \new_[64457]_ ;
  assign \new_[1365]_  = \new_[64446]_  & \new_[64433]_ ;
  assign \new_[1366]_  = \new_[64422]_  & \new_[64409]_ ;
  assign \new_[1367]_  = \new_[64398]_  & \new_[64385]_ ;
  assign \new_[1368]_  = \new_[64374]_  & \new_[64361]_ ;
  assign \new_[1369]_  = \new_[64350]_  & \new_[64337]_ ;
  assign \new_[1370]_  = \new_[64326]_  & \new_[64313]_ ;
  assign \new_[1371]_  = \new_[64302]_  & \new_[64289]_ ;
  assign \new_[1372]_  = \new_[64278]_  & \new_[64265]_ ;
  assign \new_[1373]_  = \new_[64254]_  & \new_[64241]_ ;
  assign \new_[1374]_  = \new_[64230]_  & \new_[64217]_ ;
  assign \new_[1375]_  = \new_[64206]_  & \new_[64193]_ ;
  assign \new_[1376]_  = \new_[64182]_  & \new_[64169]_ ;
  assign \new_[1377]_  = \new_[64158]_  & \new_[64145]_ ;
  assign \new_[1378]_  = \new_[64134]_  & \new_[64121]_ ;
  assign \new_[1379]_  = \new_[64110]_  & \new_[64097]_ ;
  assign \new_[1380]_  = \new_[64086]_  & \new_[64073]_ ;
  assign \new_[1381]_  = \new_[64062]_  & \new_[64049]_ ;
  assign \new_[1382]_  = \new_[64038]_  & \new_[64025]_ ;
  assign \new_[1383]_  = \new_[64014]_  & \new_[64001]_ ;
  assign \new_[1384]_  = \new_[63990]_  & \new_[63977]_ ;
  assign \new_[1385]_  = \new_[63966]_  & \new_[63953]_ ;
  assign \new_[1386]_  = \new_[63942]_  & \new_[63929]_ ;
  assign \new_[1387]_  = \new_[63918]_  & \new_[63905]_ ;
  assign \new_[1388]_  = \new_[63894]_  & \new_[63881]_ ;
  assign \new_[1389]_  = \new_[63870]_  & \new_[63857]_ ;
  assign \new_[1390]_  = \new_[63846]_  & \new_[63833]_ ;
  assign \new_[1391]_  = \new_[63822]_  & \new_[63809]_ ;
  assign \new_[1392]_  = \new_[63798]_  & \new_[63785]_ ;
  assign \new_[1393]_  = \new_[63774]_  & \new_[63761]_ ;
  assign \new_[1394]_  = \new_[63750]_  & \new_[63737]_ ;
  assign \new_[1395]_  = \new_[63726]_  & \new_[63713]_ ;
  assign \new_[1396]_  = \new_[63702]_  & \new_[63689]_ ;
  assign \new_[1397]_  = \new_[63678]_  & \new_[63665]_ ;
  assign \new_[1398]_  = \new_[63654]_  & \new_[63641]_ ;
  assign \new_[1399]_  = \new_[63630]_  & \new_[63617]_ ;
  assign \new_[1400]_  = \new_[63606]_  & \new_[63593]_ ;
  assign \new_[1401]_  = \new_[63582]_  & \new_[63569]_ ;
  assign \new_[1402]_  = \new_[63558]_  & \new_[63545]_ ;
  assign \new_[1403]_  = \new_[63534]_  & \new_[63521]_ ;
  assign \new_[1404]_  = \new_[63510]_  & \new_[63497]_ ;
  assign \new_[1405]_  = \new_[63486]_  & \new_[63473]_ ;
  assign \new_[1406]_  = \new_[63462]_  & \new_[63449]_ ;
  assign \new_[1407]_  = \new_[63438]_  & \new_[63425]_ ;
  assign \new_[1408]_  = \new_[63414]_  & \new_[63401]_ ;
  assign \new_[1409]_  = \new_[63390]_  & \new_[63377]_ ;
  assign \new_[1410]_  = \new_[63366]_  & \new_[63353]_ ;
  assign \new_[1411]_  = \new_[63342]_  & \new_[63329]_ ;
  assign \new_[1412]_  = \new_[63318]_  & \new_[63305]_ ;
  assign \new_[1413]_  = \new_[63294]_  & \new_[63281]_ ;
  assign \new_[1414]_  = \new_[63270]_  & \new_[63257]_ ;
  assign \new_[1415]_  = \new_[63246]_  & \new_[63233]_ ;
  assign \new_[1416]_  = \new_[63222]_  & \new_[63209]_ ;
  assign \new_[1417]_  = \new_[63198]_  & \new_[63185]_ ;
  assign \new_[1418]_  = \new_[63174]_  & \new_[63161]_ ;
  assign \new_[1419]_  = \new_[63150]_  & \new_[63137]_ ;
  assign \new_[1420]_  = \new_[63126]_  & \new_[63113]_ ;
  assign \new_[1421]_  = \new_[63102]_  & \new_[63089]_ ;
  assign \new_[1422]_  = \new_[63078]_  & \new_[63065]_ ;
  assign \new_[1423]_  = \new_[63054]_  & \new_[63041]_ ;
  assign \new_[1424]_  = \new_[63030]_  & \new_[63017]_ ;
  assign \new_[1425]_  = \new_[63006]_  & \new_[62993]_ ;
  assign \new_[1426]_  = \new_[62982]_  & \new_[62969]_ ;
  assign \new_[1427]_  = \new_[62958]_  & \new_[62945]_ ;
  assign \new_[1428]_  = \new_[62934]_  & \new_[62921]_ ;
  assign \new_[1429]_  = \new_[62910]_  & \new_[62897]_ ;
  assign \new_[1430]_  = \new_[62886]_  & \new_[62873]_ ;
  assign \new_[1431]_  = \new_[62862]_  & \new_[62849]_ ;
  assign \new_[1432]_  = \new_[62838]_  & \new_[62825]_ ;
  assign \new_[1433]_  = \new_[62814]_  & \new_[62801]_ ;
  assign \new_[1434]_  = \new_[62790]_  & \new_[62777]_ ;
  assign \new_[1435]_  = \new_[62766]_  & \new_[62753]_ ;
  assign \new_[1436]_  = \new_[62742]_  & \new_[62729]_ ;
  assign \new_[1437]_  = \new_[62718]_  & \new_[62705]_ ;
  assign \new_[1438]_  = \new_[62694]_  & \new_[62681]_ ;
  assign \new_[1439]_  = \new_[62670]_  & \new_[62657]_ ;
  assign \new_[1440]_  = \new_[62646]_  & \new_[62633]_ ;
  assign \new_[1441]_  = \new_[62622]_  & \new_[62609]_ ;
  assign \new_[1442]_  = \new_[62598]_  & \new_[62585]_ ;
  assign \new_[1443]_  = \new_[62574]_  & \new_[62561]_ ;
  assign \new_[1444]_  = \new_[62550]_  & \new_[62537]_ ;
  assign \new_[1445]_  = \new_[62526]_  & \new_[62513]_ ;
  assign \new_[1446]_  = \new_[62502]_  & \new_[62489]_ ;
  assign \new_[1447]_  = \new_[62478]_  & \new_[62465]_ ;
  assign \new_[1448]_  = \new_[62454]_  & \new_[62441]_ ;
  assign \new_[1449]_  = \new_[62430]_  & \new_[62417]_ ;
  assign \new_[1450]_  = \new_[62406]_  & \new_[62393]_ ;
  assign \new_[1451]_  = \new_[62382]_  & \new_[62369]_ ;
  assign \new_[1452]_  = \new_[62358]_  & \new_[62345]_ ;
  assign \new_[1453]_  = \new_[62334]_  & \new_[62321]_ ;
  assign \new_[1454]_  = \new_[62310]_  & \new_[62297]_ ;
  assign \new_[1455]_  = \new_[62286]_  & \new_[62273]_ ;
  assign \new_[1456]_  = \new_[62262]_  & \new_[62249]_ ;
  assign \new_[1457]_  = \new_[62238]_  & \new_[62225]_ ;
  assign \new_[1458]_  = \new_[62214]_  & \new_[62201]_ ;
  assign \new_[1459]_  = \new_[62190]_  & \new_[62177]_ ;
  assign \new_[1460]_  = \new_[62166]_  & \new_[62153]_ ;
  assign \new_[1461]_  = \new_[62142]_  & \new_[62129]_ ;
  assign \new_[1462]_  = \new_[62118]_  & \new_[62105]_ ;
  assign \new_[1463]_  = \new_[62094]_  & \new_[62081]_ ;
  assign \new_[1464]_  = \new_[62070]_  & \new_[62057]_ ;
  assign \new_[1465]_  = \new_[62046]_  & \new_[62033]_ ;
  assign \new_[1466]_  = \new_[62022]_  & \new_[62009]_ ;
  assign \new_[1467]_  = \new_[61998]_  & \new_[61985]_ ;
  assign \new_[1468]_  = \new_[61974]_  & \new_[61961]_ ;
  assign \new_[1469]_  = \new_[61950]_  & \new_[61937]_ ;
  assign \new_[1470]_  = \new_[61926]_  & \new_[61913]_ ;
  assign \new_[1471]_  = \new_[61902]_  & \new_[61889]_ ;
  assign \new_[1472]_  = \new_[61878]_  & \new_[61865]_ ;
  assign \new_[1473]_  = \new_[61854]_  & \new_[61841]_ ;
  assign \new_[1474]_  = \new_[61830]_  & \new_[61817]_ ;
  assign \new_[1475]_  = \new_[61806]_  & \new_[61793]_ ;
  assign \new_[1476]_  = \new_[61782]_  & \new_[61769]_ ;
  assign \new_[1477]_  = \new_[61758]_  & \new_[61745]_ ;
  assign \new_[1478]_  = \new_[61734]_  & \new_[61721]_ ;
  assign \new_[1479]_  = \new_[61710]_  & \new_[61697]_ ;
  assign \new_[1480]_  = \new_[61686]_  & \new_[61673]_ ;
  assign \new_[1481]_  = \new_[61662]_  & \new_[61649]_ ;
  assign \new_[1482]_  = \new_[61638]_  & \new_[61625]_ ;
  assign \new_[1483]_  = \new_[61614]_  & \new_[61601]_ ;
  assign \new_[1484]_  = \new_[61590]_  & \new_[61577]_ ;
  assign \new_[1485]_  = \new_[61566]_  & \new_[61553]_ ;
  assign \new_[1486]_  = \new_[61542]_  & \new_[61529]_ ;
  assign \new_[1487]_  = \new_[61518]_  & \new_[61505]_ ;
  assign \new_[1488]_  = \new_[61494]_  & \new_[61481]_ ;
  assign \new_[1489]_  = \new_[61470]_  & \new_[61457]_ ;
  assign \new_[1490]_  = \new_[61446]_  & \new_[61433]_ ;
  assign \new_[1491]_  = \new_[61422]_  & \new_[61409]_ ;
  assign \new_[1492]_  = \new_[61398]_  & \new_[61385]_ ;
  assign \new_[1493]_  = \new_[61374]_  & \new_[61361]_ ;
  assign \new_[1494]_  = \new_[61350]_  & \new_[61337]_ ;
  assign \new_[1495]_  = \new_[61326]_  & \new_[61313]_ ;
  assign \new_[1496]_  = \new_[61302]_  & \new_[61289]_ ;
  assign \new_[1497]_  = \new_[61278]_  & \new_[61265]_ ;
  assign \new_[1498]_  = \new_[61254]_  & \new_[61241]_ ;
  assign \new_[1499]_  = \new_[61230]_  & \new_[61217]_ ;
  assign \new_[1500]_  = \new_[61206]_  & \new_[61193]_ ;
  assign \new_[1501]_  = \new_[61182]_  & \new_[61169]_ ;
  assign \new_[1502]_  = \new_[61158]_  & \new_[61145]_ ;
  assign \new_[1503]_  = \new_[61134]_  & \new_[61121]_ ;
  assign \new_[1504]_  = \new_[61110]_  & \new_[61097]_ ;
  assign \new_[1505]_  = \new_[61086]_  & \new_[61073]_ ;
  assign \new_[1506]_  = \new_[61062]_  & \new_[61049]_ ;
  assign \new_[1507]_  = \new_[61038]_  & \new_[61025]_ ;
  assign \new_[1508]_  = \new_[61014]_  & \new_[61001]_ ;
  assign \new_[1509]_  = \new_[60990]_  & \new_[60977]_ ;
  assign \new_[1510]_  = \new_[60966]_  & \new_[60953]_ ;
  assign \new_[1511]_  = \new_[60942]_  & \new_[60929]_ ;
  assign \new_[1512]_  = \new_[60918]_  & \new_[60905]_ ;
  assign \new_[1513]_  = \new_[60894]_  & \new_[60881]_ ;
  assign \new_[1514]_  = \new_[60870]_  & \new_[60857]_ ;
  assign \new_[1515]_  = \new_[60846]_  & \new_[60833]_ ;
  assign \new_[1516]_  = \new_[60822]_  & \new_[60809]_ ;
  assign \new_[1517]_  = \new_[60798]_  & \new_[60785]_ ;
  assign \new_[1518]_  = \new_[60774]_  & \new_[60761]_ ;
  assign \new_[1519]_  = \new_[60750]_  & \new_[60737]_ ;
  assign \new_[1520]_  = \new_[60726]_  & \new_[60713]_ ;
  assign \new_[1521]_  = \new_[60702]_  & \new_[60689]_ ;
  assign \new_[1522]_  = \new_[60678]_  & \new_[60665]_ ;
  assign \new_[1523]_  = \new_[60654]_  & \new_[60641]_ ;
  assign \new_[1524]_  = \new_[60630]_  & \new_[60617]_ ;
  assign \new_[1525]_  = \new_[60606]_  & \new_[60593]_ ;
  assign \new_[1526]_  = \new_[60582]_  & \new_[60569]_ ;
  assign \new_[1527]_  = \new_[60558]_  & \new_[60545]_ ;
  assign \new_[1528]_  = \new_[60534]_  & \new_[60521]_ ;
  assign \new_[1529]_  = \new_[60510]_  & \new_[60497]_ ;
  assign \new_[1530]_  = \new_[60486]_  & \new_[60473]_ ;
  assign \new_[1531]_  = \new_[60462]_  & \new_[60449]_ ;
  assign \new_[1532]_  = \new_[60438]_  & \new_[60425]_ ;
  assign \new_[1533]_  = \new_[60414]_  & \new_[60401]_ ;
  assign \new_[1534]_  = \new_[60390]_  & \new_[60377]_ ;
  assign \new_[1535]_  = \new_[60366]_  & \new_[60353]_ ;
  assign \new_[1536]_  = \new_[60342]_  & \new_[60329]_ ;
  assign \new_[1537]_  = \new_[60318]_  & \new_[60305]_ ;
  assign \new_[1538]_  = \new_[60294]_  & \new_[60281]_ ;
  assign \new_[1539]_  = \new_[60270]_  & \new_[60257]_ ;
  assign \new_[1540]_  = \new_[60246]_  & \new_[60233]_ ;
  assign \new_[1541]_  = \new_[60222]_  & \new_[60209]_ ;
  assign \new_[1542]_  = \new_[60198]_  & \new_[60185]_ ;
  assign \new_[1543]_  = \new_[60174]_  & \new_[60161]_ ;
  assign \new_[1544]_  = \new_[60150]_  & \new_[60137]_ ;
  assign \new_[1545]_  = \new_[60126]_  & \new_[60113]_ ;
  assign \new_[1546]_  = \new_[60102]_  & \new_[60089]_ ;
  assign \new_[1547]_  = \new_[60078]_  & \new_[60065]_ ;
  assign \new_[1548]_  = \new_[60054]_  & \new_[60041]_ ;
  assign \new_[1549]_  = \new_[60030]_  & \new_[60017]_ ;
  assign \new_[1550]_  = \new_[60006]_  & \new_[59993]_ ;
  assign \new_[1551]_  = \new_[59982]_  & \new_[59969]_ ;
  assign \new_[1552]_  = \new_[59958]_  & \new_[59945]_ ;
  assign \new_[1553]_  = \new_[59934]_  & \new_[59921]_ ;
  assign \new_[1554]_  = \new_[59910]_  & \new_[59897]_ ;
  assign \new_[1555]_  = \new_[59886]_  & \new_[59873]_ ;
  assign \new_[1556]_  = \new_[59862]_  & \new_[59849]_ ;
  assign \new_[1557]_  = \new_[59838]_  & \new_[59825]_ ;
  assign \new_[1558]_  = \new_[59814]_  & \new_[59801]_ ;
  assign \new_[1559]_  = \new_[59790]_  & \new_[59777]_ ;
  assign \new_[1560]_  = \new_[59766]_  & \new_[59753]_ ;
  assign \new_[1561]_  = \new_[59742]_  & \new_[59729]_ ;
  assign \new_[1562]_  = \new_[59718]_  & \new_[59705]_ ;
  assign \new_[1563]_  = \new_[59694]_  & \new_[59681]_ ;
  assign \new_[1564]_  = \new_[59670]_  & \new_[59657]_ ;
  assign \new_[1565]_  = \new_[59646]_  & \new_[59633]_ ;
  assign \new_[1566]_  = \new_[59622]_  & \new_[59609]_ ;
  assign \new_[1567]_  = \new_[59598]_  & \new_[59585]_ ;
  assign \new_[1568]_  = \new_[59574]_  & \new_[59561]_ ;
  assign \new_[1569]_  = \new_[59550]_  & \new_[59537]_ ;
  assign \new_[1570]_  = \new_[59526]_  & \new_[59513]_ ;
  assign \new_[1571]_  = \new_[59502]_  & \new_[59489]_ ;
  assign \new_[1572]_  = \new_[59478]_  & \new_[59465]_ ;
  assign \new_[1573]_  = \new_[59454]_  & \new_[59441]_ ;
  assign \new_[1574]_  = \new_[59430]_  & \new_[59417]_ ;
  assign \new_[1575]_  = \new_[59406]_  & \new_[59393]_ ;
  assign \new_[1576]_  = \new_[59382]_  & \new_[59369]_ ;
  assign \new_[1577]_  = \new_[59358]_  & \new_[59345]_ ;
  assign \new_[1578]_  = \new_[59334]_  & \new_[59321]_ ;
  assign \new_[1579]_  = \new_[59310]_  & \new_[59297]_ ;
  assign \new_[1580]_  = \new_[59286]_  & \new_[59273]_ ;
  assign \new_[1581]_  = \new_[59262]_  & \new_[59249]_ ;
  assign \new_[1582]_  = \new_[59238]_  & \new_[59225]_ ;
  assign \new_[1583]_  = \new_[59214]_  & \new_[59201]_ ;
  assign \new_[1584]_  = \new_[59190]_  & \new_[59177]_ ;
  assign \new_[1585]_  = \new_[59166]_  & \new_[59153]_ ;
  assign \new_[1586]_  = \new_[59142]_  & \new_[59129]_ ;
  assign \new_[1587]_  = \new_[59118]_  & \new_[59105]_ ;
  assign \new_[1588]_  = \new_[59094]_  & \new_[59081]_ ;
  assign \new_[1589]_  = \new_[59070]_  & \new_[59057]_ ;
  assign \new_[1590]_  = \new_[59046]_  & \new_[59033]_ ;
  assign \new_[1591]_  = \new_[59022]_  & \new_[59009]_ ;
  assign \new_[1592]_  = \new_[58998]_  & \new_[58985]_ ;
  assign \new_[1593]_  = \new_[58974]_  & \new_[58961]_ ;
  assign \new_[1594]_  = \new_[58950]_  & \new_[58937]_ ;
  assign \new_[1595]_  = \new_[58926]_  & \new_[58913]_ ;
  assign \new_[1596]_  = \new_[58902]_  & \new_[58889]_ ;
  assign \new_[1597]_  = \new_[58878]_  & \new_[58865]_ ;
  assign \new_[1598]_  = \new_[58854]_  & \new_[58841]_ ;
  assign \new_[1599]_  = \new_[58830]_  & \new_[58817]_ ;
  assign \new_[1600]_  = \new_[58806]_  & \new_[58793]_ ;
  assign \new_[1601]_  = \new_[58782]_  & \new_[58769]_ ;
  assign \new_[1602]_  = \new_[58758]_  & \new_[58745]_ ;
  assign \new_[1603]_  = \new_[58734]_  & \new_[58721]_ ;
  assign \new_[1604]_  = \new_[58710]_  & \new_[58697]_ ;
  assign \new_[1605]_  = \new_[58686]_  & \new_[58673]_ ;
  assign \new_[1606]_  = \new_[58662]_  & \new_[58649]_ ;
  assign \new_[1607]_  = \new_[58638]_  & \new_[58625]_ ;
  assign \new_[1608]_  = \new_[58614]_  & \new_[58601]_ ;
  assign \new_[1609]_  = \new_[58590]_  & \new_[58577]_ ;
  assign \new_[1610]_  = \new_[58566]_  & \new_[58553]_ ;
  assign \new_[1611]_  = \new_[58542]_  & \new_[58529]_ ;
  assign \new_[1612]_  = \new_[58518]_  & \new_[58505]_ ;
  assign \new_[1613]_  = \new_[58494]_  & \new_[58481]_ ;
  assign \new_[1614]_  = \new_[58470]_  & \new_[58457]_ ;
  assign \new_[1615]_  = \new_[58446]_  & \new_[58433]_ ;
  assign \new_[1616]_  = \new_[58422]_  & \new_[58409]_ ;
  assign \new_[1617]_  = \new_[58398]_  & \new_[58385]_ ;
  assign \new_[1618]_  = \new_[58374]_  & \new_[58361]_ ;
  assign \new_[1619]_  = \new_[58350]_  & \new_[58337]_ ;
  assign \new_[1620]_  = \new_[58326]_  & \new_[58313]_ ;
  assign \new_[1621]_  = \new_[58302]_  & \new_[58289]_ ;
  assign \new_[1622]_  = \new_[58278]_  & \new_[58265]_ ;
  assign \new_[1623]_  = \new_[58254]_  & \new_[58241]_ ;
  assign \new_[1624]_  = \new_[58230]_  & \new_[58217]_ ;
  assign \new_[1625]_  = \new_[58206]_  & \new_[58193]_ ;
  assign \new_[1626]_  = \new_[58182]_  & \new_[58169]_ ;
  assign \new_[1627]_  = \new_[58158]_  & \new_[58145]_ ;
  assign \new_[1628]_  = \new_[58134]_  & \new_[58121]_ ;
  assign \new_[1629]_  = \new_[58110]_  & \new_[58097]_ ;
  assign \new_[1630]_  = \new_[58086]_  & \new_[58073]_ ;
  assign \new_[1631]_  = \new_[58062]_  & \new_[58049]_ ;
  assign \new_[1632]_  = \new_[58038]_  & \new_[58025]_ ;
  assign \new_[1633]_  = \new_[58014]_  & \new_[58001]_ ;
  assign \new_[1634]_  = \new_[57990]_  & \new_[57977]_ ;
  assign \new_[1635]_  = \new_[57966]_  & \new_[57953]_ ;
  assign \new_[1636]_  = \new_[57942]_  & \new_[57929]_ ;
  assign \new_[1637]_  = \new_[57918]_  & \new_[57905]_ ;
  assign \new_[1638]_  = \new_[57894]_  & \new_[57881]_ ;
  assign \new_[1639]_  = \new_[57870]_  & \new_[57857]_ ;
  assign \new_[1640]_  = \new_[57846]_  & \new_[57833]_ ;
  assign \new_[1641]_  = \new_[57822]_  & \new_[57809]_ ;
  assign \new_[1642]_  = \new_[57798]_  & \new_[57785]_ ;
  assign \new_[1643]_  = \new_[57774]_  & \new_[57761]_ ;
  assign \new_[1644]_  = \new_[57750]_  & \new_[57737]_ ;
  assign \new_[1645]_  = \new_[57726]_  & \new_[57713]_ ;
  assign \new_[1646]_  = \new_[57702]_  & \new_[57689]_ ;
  assign \new_[1647]_  = \new_[57678]_  & \new_[57665]_ ;
  assign \new_[1648]_  = \new_[57654]_  & \new_[57641]_ ;
  assign \new_[1649]_  = \new_[57630]_  & \new_[57617]_ ;
  assign \new_[1650]_  = \new_[57606]_  & \new_[57593]_ ;
  assign \new_[1651]_  = \new_[57582]_  & \new_[57569]_ ;
  assign \new_[1652]_  = \new_[57558]_  & \new_[57545]_ ;
  assign \new_[1653]_  = \new_[57534]_  & \new_[57521]_ ;
  assign \new_[1654]_  = \new_[57510]_  & \new_[57497]_ ;
  assign \new_[1655]_  = \new_[57486]_  & \new_[57473]_ ;
  assign \new_[1656]_  = \new_[57462]_  & \new_[57449]_ ;
  assign \new_[1657]_  = \new_[57438]_  & \new_[57425]_ ;
  assign \new_[1658]_  = \new_[57414]_  & \new_[57401]_ ;
  assign \new_[1659]_  = \new_[57390]_  & \new_[57377]_ ;
  assign \new_[1660]_  = \new_[57366]_  & \new_[57353]_ ;
  assign \new_[1661]_  = \new_[57342]_  & \new_[57329]_ ;
  assign \new_[1662]_  = \new_[57318]_  & \new_[57305]_ ;
  assign \new_[1663]_  = \new_[57294]_  & \new_[57281]_ ;
  assign \new_[1664]_  = \new_[57270]_  & \new_[57257]_ ;
  assign \new_[1665]_  = \new_[57246]_  & \new_[57233]_ ;
  assign \new_[1666]_  = \new_[57222]_  & \new_[57209]_ ;
  assign \new_[1667]_  = \new_[57198]_  & \new_[57185]_ ;
  assign \new_[1668]_  = \new_[57174]_  & \new_[57161]_ ;
  assign \new_[1669]_  = \new_[57150]_  & \new_[57137]_ ;
  assign \new_[1670]_  = \new_[57126]_  & \new_[57113]_ ;
  assign \new_[1671]_  = \new_[57102]_  & \new_[57089]_ ;
  assign \new_[1672]_  = \new_[57078]_  & \new_[57065]_ ;
  assign \new_[1673]_  = \new_[57054]_  & \new_[57041]_ ;
  assign \new_[1674]_  = \new_[57030]_  & \new_[57017]_ ;
  assign \new_[1675]_  = \new_[57006]_  & \new_[56993]_ ;
  assign \new_[1676]_  = \new_[56982]_  & \new_[56969]_ ;
  assign \new_[1677]_  = \new_[56958]_  & \new_[56945]_ ;
  assign \new_[1678]_  = \new_[56934]_  & \new_[56921]_ ;
  assign \new_[1679]_  = \new_[56910]_  & \new_[56897]_ ;
  assign \new_[1680]_  = \new_[56886]_  & \new_[56873]_ ;
  assign \new_[1681]_  = \new_[56862]_  & \new_[56849]_ ;
  assign \new_[1682]_  = \new_[56838]_  & \new_[56825]_ ;
  assign \new_[1683]_  = \new_[56814]_  & \new_[56801]_ ;
  assign \new_[1684]_  = \new_[56790]_  & \new_[56777]_ ;
  assign \new_[1685]_  = \new_[56766]_  & \new_[56753]_ ;
  assign \new_[1686]_  = \new_[56742]_  & \new_[56729]_ ;
  assign \new_[1687]_  = \new_[56718]_  & \new_[56705]_ ;
  assign \new_[1688]_  = \new_[56694]_  & \new_[56681]_ ;
  assign \new_[1689]_  = \new_[56670]_  & \new_[56657]_ ;
  assign \new_[1690]_  = \new_[56646]_  & \new_[56633]_ ;
  assign \new_[1691]_  = \new_[56622]_  & \new_[56609]_ ;
  assign \new_[1692]_  = \new_[56598]_  & \new_[56585]_ ;
  assign \new_[1693]_  = \new_[56574]_  & \new_[56561]_ ;
  assign \new_[1694]_  = \new_[56550]_  & \new_[56537]_ ;
  assign \new_[1695]_  = \new_[56526]_  & \new_[56513]_ ;
  assign \new_[1696]_  = \new_[56502]_  & \new_[56489]_ ;
  assign \new_[1697]_  = \new_[56478]_  & \new_[56465]_ ;
  assign \new_[1698]_  = \new_[56454]_  & \new_[56441]_ ;
  assign \new_[1699]_  = \new_[56430]_  & \new_[56417]_ ;
  assign \new_[1700]_  = \new_[56406]_  & \new_[56393]_ ;
  assign \new_[1701]_  = \new_[56382]_  & \new_[56369]_ ;
  assign \new_[1702]_  = \new_[56358]_  & \new_[56345]_ ;
  assign \new_[1703]_  = \new_[56334]_  & \new_[56321]_ ;
  assign \new_[1704]_  = \new_[56310]_  & \new_[56297]_ ;
  assign \new_[1705]_  = \new_[56286]_  & \new_[56273]_ ;
  assign \new_[1706]_  = \new_[56262]_  & \new_[56249]_ ;
  assign \new_[1707]_  = \new_[56238]_  & \new_[56225]_ ;
  assign \new_[1708]_  = \new_[56214]_  & \new_[56201]_ ;
  assign \new_[1709]_  = \new_[56190]_  & \new_[56177]_ ;
  assign \new_[1710]_  = \new_[56166]_  & \new_[56153]_ ;
  assign \new_[1711]_  = \new_[56142]_  & \new_[56129]_ ;
  assign \new_[1712]_  = \new_[56118]_  & \new_[56105]_ ;
  assign \new_[1713]_  = \new_[56094]_  & \new_[56081]_ ;
  assign \new_[1714]_  = \new_[56070]_  & \new_[56057]_ ;
  assign \new_[1715]_  = \new_[56046]_  & \new_[56033]_ ;
  assign \new_[1716]_  = \new_[56022]_  & \new_[56009]_ ;
  assign \new_[1717]_  = \new_[55998]_  & \new_[55985]_ ;
  assign \new_[1718]_  = \new_[55974]_  & \new_[55961]_ ;
  assign \new_[1719]_  = \new_[55950]_  & \new_[55937]_ ;
  assign \new_[1720]_  = \new_[55926]_  & \new_[55913]_ ;
  assign \new_[1721]_  = \new_[55902]_  & \new_[55889]_ ;
  assign \new_[1722]_  = \new_[55878]_  & \new_[55865]_ ;
  assign \new_[1723]_  = \new_[55854]_  & \new_[55841]_ ;
  assign \new_[1724]_  = \new_[55830]_  & \new_[55817]_ ;
  assign \new_[1725]_  = \new_[55806]_  & \new_[55793]_ ;
  assign \new_[1726]_  = \new_[55782]_  & \new_[55769]_ ;
  assign \new_[1727]_  = \new_[55758]_  & \new_[55745]_ ;
  assign \new_[1728]_  = \new_[55734]_  & \new_[55721]_ ;
  assign \new_[1729]_  = \new_[55710]_  & \new_[55697]_ ;
  assign \new_[1730]_  = \new_[55686]_  & \new_[55673]_ ;
  assign \new_[1731]_  = \new_[55662]_  & \new_[55649]_ ;
  assign \new_[1732]_  = \new_[55638]_  & \new_[55625]_ ;
  assign \new_[1733]_  = \new_[55614]_  & \new_[55601]_ ;
  assign \new_[1734]_  = \new_[55590]_  & \new_[55577]_ ;
  assign \new_[1735]_  = \new_[55566]_  & \new_[55553]_ ;
  assign \new_[1736]_  = \new_[55542]_  & \new_[55529]_ ;
  assign \new_[1737]_  = \new_[55518]_  & \new_[55505]_ ;
  assign \new_[1738]_  = \new_[55494]_  & \new_[55481]_ ;
  assign \new_[1739]_  = \new_[55470]_  & \new_[55457]_ ;
  assign \new_[1740]_  = \new_[55446]_  & \new_[55433]_ ;
  assign \new_[1741]_  = \new_[55422]_  & \new_[55409]_ ;
  assign \new_[1742]_  = \new_[55398]_  & \new_[55385]_ ;
  assign \new_[1743]_  = \new_[55374]_  & \new_[55361]_ ;
  assign \new_[1744]_  = \new_[55350]_  & \new_[55337]_ ;
  assign \new_[1745]_  = \new_[55326]_  & \new_[55313]_ ;
  assign \new_[1746]_  = \new_[55302]_  & \new_[55289]_ ;
  assign \new_[1747]_  = \new_[55278]_  & \new_[55265]_ ;
  assign \new_[1748]_  = \new_[55254]_  & \new_[55241]_ ;
  assign \new_[1749]_  = \new_[55230]_  & \new_[55217]_ ;
  assign \new_[1750]_  = \new_[55206]_  & \new_[55193]_ ;
  assign \new_[1751]_  = \new_[55182]_  & \new_[55169]_ ;
  assign \new_[1752]_  = \new_[55158]_  & \new_[55145]_ ;
  assign \new_[1753]_  = \new_[55134]_  & \new_[55121]_ ;
  assign \new_[1754]_  = \new_[55110]_  & \new_[55097]_ ;
  assign \new_[1755]_  = \new_[55086]_  & \new_[55073]_ ;
  assign \new_[1756]_  = \new_[55062]_  & \new_[55049]_ ;
  assign \new_[1757]_  = \new_[55038]_  & \new_[55025]_ ;
  assign \new_[1758]_  = \new_[55014]_  & \new_[55001]_ ;
  assign \new_[1759]_  = \new_[54990]_  & \new_[54977]_ ;
  assign \new_[1760]_  = \new_[54966]_  & \new_[54953]_ ;
  assign \new_[1761]_  = \new_[54942]_  & \new_[54929]_ ;
  assign \new_[1762]_  = \new_[54918]_  & \new_[54905]_ ;
  assign \new_[1763]_  = \new_[54894]_  & \new_[54881]_ ;
  assign \new_[1764]_  = \new_[54870]_  & \new_[54857]_ ;
  assign \new_[1765]_  = \new_[54846]_  & \new_[54833]_ ;
  assign \new_[1766]_  = \new_[54822]_  & \new_[54809]_ ;
  assign \new_[1767]_  = \new_[54798]_  & \new_[54785]_ ;
  assign \new_[1768]_  = \new_[54774]_  & \new_[54761]_ ;
  assign \new_[1769]_  = \new_[54750]_  & \new_[54737]_ ;
  assign \new_[1770]_  = \new_[54726]_  & \new_[54713]_ ;
  assign \new_[1771]_  = \new_[54702]_  & \new_[54689]_ ;
  assign \new_[1772]_  = \new_[54678]_  & \new_[54665]_ ;
  assign \new_[1773]_  = \new_[54654]_  & \new_[54641]_ ;
  assign \new_[1774]_  = \new_[54630]_  & \new_[54617]_ ;
  assign \new_[1775]_  = \new_[54606]_  & \new_[54593]_ ;
  assign \new_[1776]_  = \new_[54582]_  & \new_[54569]_ ;
  assign \new_[1777]_  = \new_[54558]_  & \new_[54545]_ ;
  assign \new_[1778]_  = \new_[54534]_  & \new_[54521]_ ;
  assign \new_[1779]_  = \new_[54510]_  & \new_[54497]_ ;
  assign \new_[1780]_  = \new_[54486]_  & \new_[54473]_ ;
  assign \new_[1781]_  = \new_[54462]_  & \new_[54449]_ ;
  assign \new_[1782]_  = \new_[54438]_  & \new_[54425]_ ;
  assign \new_[1783]_  = \new_[54414]_  & \new_[54401]_ ;
  assign \new_[1784]_  = \new_[54390]_  & \new_[54377]_ ;
  assign \new_[1785]_  = \new_[54366]_  & \new_[54353]_ ;
  assign \new_[1786]_  = \new_[54342]_  & \new_[54329]_ ;
  assign \new_[1787]_  = \new_[54318]_  & \new_[54305]_ ;
  assign \new_[1788]_  = \new_[54294]_  & \new_[54281]_ ;
  assign \new_[1789]_  = \new_[54270]_  & \new_[54257]_ ;
  assign \new_[1790]_  = \new_[54246]_  & \new_[54233]_ ;
  assign \new_[1791]_  = \new_[54222]_  & \new_[54209]_ ;
  assign \new_[1792]_  = \new_[54198]_  & \new_[54185]_ ;
  assign \new_[1793]_  = \new_[54174]_  & \new_[54161]_ ;
  assign \new_[1794]_  = \new_[54150]_  & \new_[54137]_ ;
  assign \new_[1795]_  = \new_[54126]_  & \new_[54113]_ ;
  assign \new_[1796]_  = \new_[54102]_  & \new_[54089]_ ;
  assign \new_[1797]_  = \new_[54078]_  & \new_[54065]_ ;
  assign \new_[1798]_  = \new_[54054]_  & \new_[54041]_ ;
  assign \new_[1799]_  = \new_[54030]_  & \new_[54017]_ ;
  assign \new_[1800]_  = \new_[54006]_  & \new_[53993]_ ;
  assign \new_[1801]_  = \new_[53982]_  & \new_[53969]_ ;
  assign \new_[1802]_  = \new_[53958]_  & \new_[53945]_ ;
  assign \new_[1803]_  = \new_[53934]_  & \new_[53921]_ ;
  assign \new_[1804]_  = \new_[53910]_  & \new_[53897]_ ;
  assign \new_[1805]_  = \new_[53886]_  & \new_[53873]_ ;
  assign \new_[1806]_  = \new_[53862]_  & \new_[53849]_ ;
  assign \new_[1807]_  = \new_[53838]_  & \new_[53825]_ ;
  assign \new_[1808]_  = \new_[53814]_  & \new_[53801]_ ;
  assign \new_[1809]_  = \new_[53790]_  & \new_[53777]_ ;
  assign \new_[1810]_  = \new_[53766]_  & \new_[53753]_ ;
  assign \new_[1811]_  = \new_[53742]_  & \new_[53729]_ ;
  assign \new_[1812]_  = \new_[53718]_  & \new_[53705]_ ;
  assign \new_[1813]_  = \new_[53694]_  & \new_[53681]_ ;
  assign \new_[1814]_  = \new_[53670]_  & \new_[53657]_ ;
  assign \new_[1815]_  = \new_[53646]_  & \new_[53633]_ ;
  assign \new_[1816]_  = \new_[53622]_  & \new_[53609]_ ;
  assign \new_[1817]_  = \new_[53598]_  & \new_[53585]_ ;
  assign \new_[1818]_  = \new_[53574]_  & \new_[53561]_ ;
  assign \new_[1819]_  = \new_[53550]_  & \new_[53537]_ ;
  assign \new_[1820]_  = \new_[53526]_  & \new_[53513]_ ;
  assign \new_[1821]_  = \new_[53502]_  & \new_[53489]_ ;
  assign \new_[1822]_  = \new_[53478]_  & \new_[53465]_ ;
  assign \new_[1823]_  = \new_[53454]_  & \new_[53441]_ ;
  assign \new_[1824]_  = \new_[53430]_  & \new_[53417]_ ;
  assign \new_[1825]_  = \new_[53406]_  & \new_[53393]_ ;
  assign \new_[1826]_  = \new_[53382]_  & \new_[53369]_ ;
  assign \new_[1827]_  = \new_[53358]_  & \new_[53345]_ ;
  assign \new_[1828]_  = \new_[53334]_  & \new_[53321]_ ;
  assign \new_[1829]_  = \new_[53310]_  & \new_[53297]_ ;
  assign \new_[1830]_  = \new_[53286]_  & \new_[53273]_ ;
  assign \new_[1831]_  = \new_[53262]_  & \new_[53249]_ ;
  assign \new_[1832]_  = \new_[53238]_  & \new_[53225]_ ;
  assign \new_[1833]_  = \new_[53214]_  & \new_[53201]_ ;
  assign \new_[1834]_  = \new_[53190]_  & \new_[53177]_ ;
  assign \new_[1835]_  = \new_[53166]_  & \new_[53153]_ ;
  assign \new_[1836]_  = \new_[53142]_  & \new_[53129]_ ;
  assign \new_[1837]_  = \new_[53118]_  & \new_[53105]_ ;
  assign \new_[1838]_  = \new_[53094]_  & \new_[53081]_ ;
  assign \new_[1839]_  = \new_[53070]_  & \new_[53057]_ ;
  assign \new_[1840]_  = \new_[53046]_  & \new_[53033]_ ;
  assign \new_[1841]_  = \new_[53022]_  & \new_[53009]_ ;
  assign \new_[1842]_  = \new_[52998]_  & \new_[52985]_ ;
  assign \new_[1843]_  = \new_[52974]_  & \new_[52961]_ ;
  assign \new_[1844]_  = \new_[52950]_  & \new_[52937]_ ;
  assign \new_[1845]_  = \new_[52926]_  & \new_[52913]_ ;
  assign \new_[1846]_  = \new_[52902]_  & \new_[52889]_ ;
  assign \new_[1847]_  = \new_[52878]_  & \new_[52865]_ ;
  assign \new_[1848]_  = \new_[52854]_  & \new_[52841]_ ;
  assign \new_[1849]_  = \new_[52830]_  & \new_[52817]_ ;
  assign \new_[1850]_  = \new_[52806]_  & \new_[52793]_ ;
  assign \new_[1851]_  = \new_[52782]_  & \new_[52769]_ ;
  assign \new_[1852]_  = \new_[52758]_  & \new_[52745]_ ;
  assign \new_[1853]_  = \new_[52734]_  & \new_[52721]_ ;
  assign \new_[1854]_  = \new_[52710]_  & \new_[52697]_ ;
  assign \new_[1855]_  = \new_[52686]_  & \new_[52673]_ ;
  assign \new_[1856]_  = \new_[52662]_  & \new_[52649]_ ;
  assign \new_[1857]_  = \new_[52638]_  & \new_[52625]_ ;
  assign \new_[1858]_  = \new_[52614]_  & \new_[52601]_ ;
  assign \new_[1859]_  = \new_[52590]_  & \new_[52577]_ ;
  assign \new_[1860]_  = \new_[52566]_  & \new_[52553]_ ;
  assign \new_[1861]_  = \new_[52542]_  & \new_[52529]_ ;
  assign \new_[1862]_  = \new_[52518]_  & \new_[52505]_ ;
  assign \new_[1863]_  = \new_[52494]_  & \new_[52481]_ ;
  assign \new_[1864]_  = \new_[52470]_  & \new_[52457]_ ;
  assign \new_[1865]_  = \new_[52446]_  & \new_[52433]_ ;
  assign \new_[1866]_  = \new_[52422]_  & \new_[52409]_ ;
  assign \new_[1867]_  = \new_[52398]_  & \new_[52385]_ ;
  assign \new_[1868]_  = \new_[52374]_  & \new_[52361]_ ;
  assign \new_[1869]_  = \new_[52350]_  & \new_[52337]_ ;
  assign \new_[1870]_  = \new_[52326]_  & \new_[52313]_ ;
  assign \new_[1871]_  = \new_[52302]_  & \new_[52289]_ ;
  assign \new_[1872]_  = \new_[52278]_  & \new_[52265]_ ;
  assign \new_[1873]_  = \new_[52254]_  & \new_[52241]_ ;
  assign \new_[1874]_  = \new_[52230]_  & \new_[52217]_ ;
  assign \new_[1875]_  = \new_[52206]_  & \new_[52193]_ ;
  assign \new_[1876]_  = \new_[52182]_  & \new_[52169]_ ;
  assign \new_[1877]_  = \new_[52158]_  & \new_[52145]_ ;
  assign \new_[1878]_  = \new_[52134]_  & \new_[52121]_ ;
  assign \new_[1879]_  = \new_[52110]_  & \new_[52097]_ ;
  assign \new_[1880]_  = \new_[52086]_  & \new_[52073]_ ;
  assign \new_[1881]_  = \new_[52062]_  & \new_[52049]_ ;
  assign \new_[1882]_  = \new_[52038]_  & \new_[52025]_ ;
  assign \new_[1883]_  = \new_[52014]_  & \new_[52001]_ ;
  assign \new_[1884]_  = \new_[51990]_  & \new_[51977]_ ;
  assign \new_[1885]_  = \new_[51966]_  & \new_[51953]_ ;
  assign \new_[1886]_  = \new_[51942]_  & \new_[51929]_ ;
  assign \new_[1887]_  = \new_[51918]_  & \new_[51905]_ ;
  assign \new_[1888]_  = \new_[51894]_  & \new_[51881]_ ;
  assign \new_[1889]_  = \new_[51870]_  & \new_[51857]_ ;
  assign \new_[1890]_  = \new_[51846]_  & \new_[51833]_ ;
  assign \new_[1891]_  = \new_[51822]_  & \new_[51809]_ ;
  assign \new_[1892]_  = \new_[51798]_  & \new_[51785]_ ;
  assign \new_[1893]_  = \new_[51774]_  & \new_[51761]_ ;
  assign \new_[1894]_  = \new_[51750]_  & \new_[51737]_ ;
  assign \new_[1895]_  = \new_[51726]_  & \new_[51713]_ ;
  assign \new_[1896]_  = \new_[51702]_  & \new_[51689]_ ;
  assign \new_[1897]_  = \new_[51678]_  & \new_[51665]_ ;
  assign \new_[1898]_  = \new_[51654]_  & \new_[51641]_ ;
  assign \new_[1899]_  = \new_[51630]_  & \new_[51617]_ ;
  assign \new_[1900]_  = \new_[51606]_  & \new_[51593]_ ;
  assign \new_[1901]_  = \new_[51582]_  & \new_[51569]_ ;
  assign \new_[1902]_  = \new_[51558]_  & \new_[51545]_ ;
  assign \new_[1903]_  = \new_[51534]_  & \new_[51521]_ ;
  assign \new_[1904]_  = \new_[51510]_  & \new_[51497]_ ;
  assign \new_[1905]_  = \new_[51486]_  & \new_[51473]_ ;
  assign \new_[1906]_  = \new_[51462]_  & \new_[51449]_ ;
  assign \new_[1907]_  = \new_[51438]_  & \new_[51425]_ ;
  assign \new_[1908]_  = \new_[51414]_  & \new_[51401]_ ;
  assign \new_[1909]_  = \new_[51390]_  & \new_[51377]_ ;
  assign \new_[1910]_  = \new_[51366]_  & \new_[51353]_ ;
  assign \new_[1911]_  = \new_[51342]_  & \new_[51329]_ ;
  assign \new_[1912]_  = \new_[51318]_  & \new_[51305]_ ;
  assign \new_[1913]_  = \new_[51294]_  & \new_[51281]_ ;
  assign \new_[1914]_  = \new_[51270]_  & \new_[51257]_ ;
  assign \new_[1915]_  = \new_[51246]_  & \new_[51233]_ ;
  assign \new_[1916]_  = \new_[51222]_  & \new_[51209]_ ;
  assign \new_[1917]_  = \new_[51198]_  & \new_[51185]_ ;
  assign \new_[1918]_  = \new_[51174]_  & \new_[51161]_ ;
  assign \new_[1919]_  = \new_[51150]_  & \new_[51137]_ ;
  assign \new_[1920]_  = \new_[51126]_  & \new_[51113]_ ;
  assign \new_[1921]_  = \new_[51102]_  & \new_[51089]_ ;
  assign \new_[1922]_  = \new_[51078]_  & \new_[51065]_ ;
  assign \new_[1923]_  = \new_[51054]_  & \new_[51041]_ ;
  assign \new_[1924]_  = \new_[51030]_  & \new_[51017]_ ;
  assign \new_[1925]_  = \new_[51006]_  & \new_[50993]_ ;
  assign \new_[1926]_  = \new_[50982]_  & \new_[50969]_ ;
  assign \new_[1927]_  = \new_[50958]_  & \new_[50945]_ ;
  assign \new_[1928]_  = \new_[50934]_  & \new_[50921]_ ;
  assign \new_[1929]_  = \new_[50910]_  & \new_[50897]_ ;
  assign \new_[1930]_  = \new_[50886]_  & \new_[50873]_ ;
  assign \new_[1931]_  = \new_[50862]_  & \new_[50849]_ ;
  assign \new_[1932]_  = \new_[50838]_  & \new_[50825]_ ;
  assign \new_[1933]_  = \new_[50814]_  & \new_[50801]_ ;
  assign \new_[1934]_  = \new_[50790]_  & \new_[50777]_ ;
  assign \new_[1935]_  = \new_[50766]_  & \new_[50753]_ ;
  assign \new_[1936]_  = \new_[50742]_  & \new_[50729]_ ;
  assign \new_[1937]_  = \new_[50718]_  & \new_[50705]_ ;
  assign \new_[1938]_  = \new_[50694]_  & \new_[50681]_ ;
  assign \new_[1939]_  = \new_[50670]_  & \new_[50657]_ ;
  assign \new_[1940]_  = \new_[50646]_  & \new_[50633]_ ;
  assign \new_[1941]_  = \new_[50622]_  & \new_[50609]_ ;
  assign \new_[1942]_  = \new_[50598]_  & \new_[50585]_ ;
  assign \new_[1943]_  = \new_[50574]_  & \new_[50561]_ ;
  assign \new_[1944]_  = \new_[50550]_  & \new_[50537]_ ;
  assign \new_[1945]_  = \new_[50526]_  & \new_[50513]_ ;
  assign \new_[1946]_  = \new_[50502]_  & \new_[50489]_ ;
  assign \new_[1947]_  = \new_[50478]_  & \new_[50465]_ ;
  assign \new_[1948]_  = \new_[50454]_  & \new_[50441]_ ;
  assign \new_[1949]_  = \new_[50430]_  & \new_[50417]_ ;
  assign \new_[1950]_  = \new_[50406]_  & \new_[50393]_ ;
  assign \new_[1951]_  = \new_[50382]_  & \new_[50369]_ ;
  assign \new_[1952]_  = \new_[50358]_  & \new_[50345]_ ;
  assign \new_[1953]_  = \new_[50334]_  & \new_[50321]_ ;
  assign \new_[1954]_  = \new_[50310]_  & \new_[50297]_ ;
  assign \new_[1955]_  = \new_[50286]_  & \new_[50273]_ ;
  assign \new_[1956]_  = \new_[50262]_  & \new_[50249]_ ;
  assign \new_[1957]_  = \new_[50238]_  & \new_[50225]_ ;
  assign \new_[1958]_  = \new_[50214]_  & \new_[50201]_ ;
  assign \new_[1959]_  = \new_[50190]_  & \new_[50177]_ ;
  assign \new_[1960]_  = \new_[50166]_  & \new_[50153]_ ;
  assign \new_[1961]_  = \new_[50142]_  & \new_[50129]_ ;
  assign \new_[1962]_  = \new_[50118]_  & \new_[50105]_ ;
  assign \new_[1963]_  = \new_[50094]_  & \new_[50081]_ ;
  assign \new_[1964]_  = \new_[50070]_  & \new_[50057]_ ;
  assign \new_[1965]_  = \new_[50046]_  & \new_[50033]_ ;
  assign \new_[1966]_  = \new_[50022]_  & \new_[50009]_ ;
  assign \new_[1967]_  = \new_[49998]_  & \new_[49985]_ ;
  assign \new_[1968]_  = \new_[49974]_  & \new_[49961]_ ;
  assign \new_[1969]_  = \new_[49950]_  & \new_[49937]_ ;
  assign \new_[1970]_  = \new_[49926]_  & \new_[49913]_ ;
  assign \new_[1971]_  = \new_[49902]_  & \new_[49889]_ ;
  assign \new_[1972]_  = \new_[49878]_  & \new_[49865]_ ;
  assign \new_[1973]_  = \new_[49854]_  & \new_[49841]_ ;
  assign \new_[1974]_  = \new_[49830]_  & \new_[49817]_ ;
  assign \new_[1975]_  = \new_[49806]_  & \new_[49793]_ ;
  assign \new_[1976]_  = \new_[49782]_  & \new_[49769]_ ;
  assign \new_[1977]_  = \new_[49758]_  & \new_[49745]_ ;
  assign \new_[1978]_  = \new_[49734]_  & \new_[49721]_ ;
  assign \new_[1979]_  = \new_[49710]_  & \new_[49697]_ ;
  assign \new_[1980]_  = \new_[49686]_  & \new_[49673]_ ;
  assign \new_[1981]_  = \new_[49662]_  & \new_[49649]_ ;
  assign \new_[1982]_  = \new_[49638]_  & \new_[49625]_ ;
  assign \new_[1983]_  = \new_[49614]_  & \new_[49601]_ ;
  assign \new_[1984]_  = \new_[49590]_  & \new_[49577]_ ;
  assign \new_[1985]_  = \new_[49566]_  & \new_[49553]_ ;
  assign \new_[1986]_  = \new_[49542]_  & \new_[49529]_ ;
  assign \new_[1987]_  = \new_[49518]_  & \new_[49505]_ ;
  assign \new_[1988]_  = \new_[49494]_  & \new_[49481]_ ;
  assign \new_[1989]_  = \new_[49470]_  & \new_[49457]_ ;
  assign \new_[1990]_  = \new_[49446]_  & \new_[49433]_ ;
  assign \new_[1991]_  = \new_[49422]_  & \new_[49409]_ ;
  assign \new_[1992]_  = \new_[49398]_  & \new_[49385]_ ;
  assign \new_[1993]_  = \new_[49374]_  & \new_[49361]_ ;
  assign \new_[1994]_  = \new_[49350]_  & \new_[49337]_ ;
  assign \new_[1995]_  = \new_[49326]_  & \new_[49313]_ ;
  assign \new_[1996]_  = \new_[49302]_  & \new_[49289]_ ;
  assign \new_[1997]_  = \new_[49278]_  & \new_[49265]_ ;
  assign \new_[1998]_  = \new_[49254]_  & \new_[49241]_ ;
  assign \new_[1999]_  = \new_[49230]_  & \new_[49217]_ ;
  assign \new_[2000]_  = \new_[49206]_  & \new_[49193]_ ;
  assign \new_[2001]_  = \new_[49182]_  & \new_[49169]_ ;
  assign \new_[2002]_  = \new_[49158]_  & \new_[49145]_ ;
  assign \new_[2003]_  = \new_[49134]_  & \new_[49121]_ ;
  assign \new_[2004]_  = \new_[49110]_  & \new_[49097]_ ;
  assign \new_[2005]_  = \new_[49086]_  & \new_[49073]_ ;
  assign \new_[2006]_  = \new_[49062]_  & \new_[49049]_ ;
  assign \new_[2007]_  = \new_[49038]_  & \new_[49025]_ ;
  assign \new_[2008]_  = \new_[49014]_  & \new_[49001]_ ;
  assign \new_[2009]_  = \new_[48990]_  & \new_[48977]_ ;
  assign \new_[2010]_  = \new_[48966]_  & \new_[48953]_ ;
  assign \new_[2011]_  = \new_[48942]_  & \new_[48929]_ ;
  assign \new_[2012]_  = \new_[48918]_  & \new_[48905]_ ;
  assign \new_[2013]_  = \new_[48894]_  & \new_[48881]_ ;
  assign \new_[2014]_  = \new_[48870]_  & \new_[48857]_ ;
  assign \new_[2015]_  = \new_[48846]_  & \new_[48833]_ ;
  assign \new_[2016]_  = \new_[48822]_  & \new_[48809]_ ;
  assign \new_[2017]_  = \new_[48798]_  & \new_[48785]_ ;
  assign \new_[2018]_  = \new_[48774]_  & \new_[48761]_ ;
  assign \new_[2019]_  = \new_[48750]_  & \new_[48737]_ ;
  assign \new_[2020]_  = \new_[48726]_  & \new_[48713]_ ;
  assign \new_[2021]_  = \new_[48702]_  & \new_[48689]_ ;
  assign \new_[2022]_  = \new_[48678]_  & \new_[48665]_ ;
  assign \new_[2023]_  = \new_[48654]_  & \new_[48641]_ ;
  assign \new_[2024]_  = \new_[48630]_  & \new_[48617]_ ;
  assign \new_[2025]_  = \new_[48606]_  & \new_[48593]_ ;
  assign \new_[2026]_  = \new_[48582]_  & \new_[48569]_ ;
  assign \new_[2027]_  = \new_[48558]_  & \new_[48545]_ ;
  assign \new_[2028]_  = \new_[48534]_  & \new_[48521]_ ;
  assign \new_[2029]_  = \new_[48510]_  & \new_[48497]_ ;
  assign \new_[2030]_  = \new_[48486]_  & \new_[48473]_ ;
  assign \new_[2031]_  = \new_[48462]_  & \new_[48449]_ ;
  assign \new_[2032]_  = \new_[48438]_  & \new_[48425]_ ;
  assign \new_[2033]_  = \new_[48414]_  & \new_[48401]_ ;
  assign \new_[2034]_  = \new_[48390]_  & \new_[48377]_ ;
  assign \new_[2035]_  = \new_[48366]_  & \new_[48353]_ ;
  assign \new_[2036]_  = \new_[48342]_  & \new_[48329]_ ;
  assign \new_[2037]_  = \new_[48318]_  & \new_[48305]_ ;
  assign \new_[2038]_  = \new_[48294]_  & \new_[48281]_ ;
  assign \new_[2039]_  = \new_[48270]_  & \new_[48257]_ ;
  assign \new_[2040]_  = \new_[48246]_  & \new_[48233]_ ;
  assign \new_[2041]_  = \new_[48222]_  & \new_[48209]_ ;
  assign \new_[2042]_  = \new_[48198]_  & \new_[48185]_ ;
  assign \new_[2043]_  = \new_[48174]_  & \new_[48161]_ ;
  assign \new_[2044]_  = \new_[48150]_  & \new_[48137]_ ;
  assign \new_[2045]_  = \new_[48126]_  & \new_[48113]_ ;
  assign \new_[2046]_  = \new_[48102]_  & \new_[48089]_ ;
  assign \new_[2047]_  = \new_[48078]_  & \new_[48065]_ ;
  assign \new_[2048]_  = \new_[48054]_  & \new_[48041]_ ;
  assign \new_[2049]_  = \new_[48030]_  & \new_[48017]_ ;
  assign \new_[2050]_  = \new_[48006]_  & \new_[47993]_ ;
  assign \new_[2051]_  = \new_[47982]_  & \new_[47969]_ ;
  assign \new_[2052]_  = \new_[47958]_  & \new_[47945]_ ;
  assign \new_[2053]_  = \new_[47934]_  & \new_[47921]_ ;
  assign \new_[2054]_  = \new_[47910]_  & \new_[47897]_ ;
  assign \new_[2055]_  = \new_[47886]_  & \new_[47873]_ ;
  assign \new_[2056]_  = \new_[47862]_  & \new_[47849]_ ;
  assign \new_[2057]_  = \new_[47838]_  & \new_[47825]_ ;
  assign \new_[2058]_  = \new_[47814]_  & \new_[47801]_ ;
  assign \new_[2059]_  = \new_[47790]_  & \new_[47777]_ ;
  assign \new_[2060]_  = \new_[47766]_  & \new_[47753]_ ;
  assign \new_[2061]_  = \new_[47742]_  & \new_[47729]_ ;
  assign \new_[2062]_  = \new_[47718]_  & \new_[47705]_ ;
  assign \new_[2063]_  = \new_[47694]_  & \new_[47681]_ ;
  assign \new_[2064]_  = \new_[47670]_  & \new_[47657]_ ;
  assign \new_[2065]_  = \new_[47646]_  & \new_[47633]_ ;
  assign \new_[2066]_  = \new_[47622]_  & \new_[47609]_ ;
  assign \new_[2067]_  = \new_[47598]_  & \new_[47585]_ ;
  assign \new_[2068]_  = \new_[47574]_  & \new_[47561]_ ;
  assign \new_[2069]_  = \new_[47550]_  & \new_[47537]_ ;
  assign \new_[2070]_  = \new_[47526]_  & \new_[47513]_ ;
  assign \new_[2071]_  = \new_[47502]_  & \new_[47489]_ ;
  assign \new_[2072]_  = \new_[47478]_  & \new_[47465]_ ;
  assign \new_[2073]_  = \new_[47454]_  & \new_[47441]_ ;
  assign \new_[2074]_  = \new_[47430]_  & \new_[47417]_ ;
  assign \new_[2075]_  = \new_[47406]_  & \new_[47393]_ ;
  assign \new_[2076]_  = \new_[47382]_  & \new_[47369]_ ;
  assign \new_[2077]_  = \new_[47358]_  & \new_[47345]_ ;
  assign \new_[2078]_  = \new_[47334]_  & \new_[47321]_ ;
  assign \new_[2079]_  = \new_[47310]_  & \new_[47297]_ ;
  assign \new_[2080]_  = \new_[47286]_  & \new_[47273]_ ;
  assign \new_[2081]_  = \new_[47262]_  & \new_[47249]_ ;
  assign \new_[2082]_  = \new_[47238]_  & \new_[47225]_ ;
  assign \new_[2083]_  = \new_[47214]_  & \new_[47201]_ ;
  assign \new_[2084]_  = \new_[47190]_  & \new_[47177]_ ;
  assign \new_[2085]_  = \new_[47166]_  & \new_[47153]_ ;
  assign \new_[2086]_  = \new_[47142]_  & \new_[47129]_ ;
  assign \new_[2087]_  = \new_[47118]_  & \new_[47105]_ ;
  assign \new_[2088]_  = \new_[47094]_  & \new_[47081]_ ;
  assign \new_[2089]_  = \new_[47070]_  & \new_[47057]_ ;
  assign \new_[2090]_  = \new_[47046]_  & \new_[47033]_ ;
  assign \new_[2091]_  = \new_[47022]_  & \new_[47009]_ ;
  assign \new_[2092]_  = \new_[46998]_  & \new_[46985]_ ;
  assign \new_[2093]_  = \new_[46974]_  & \new_[46961]_ ;
  assign \new_[2094]_  = \new_[46950]_  & \new_[46937]_ ;
  assign \new_[2095]_  = \new_[46926]_  & \new_[46913]_ ;
  assign \new_[2096]_  = \new_[46902]_  & \new_[46889]_ ;
  assign \new_[2097]_  = \new_[46878]_  & \new_[46865]_ ;
  assign \new_[2098]_  = \new_[46854]_  & \new_[46841]_ ;
  assign \new_[2099]_  = \new_[46830]_  & \new_[46817]_ ;
  assign \new_[2100]_  = \new_[46806]_  & \new_[46793]_ ;
  assign \new_[2101]_  = \new_[46782]_  & \new_[46769]_ ;
  assign \new_[2102]_  = \new_[46758]_  & \new_[46745]_ ;
  assign \new_[2103]_  = \new_[46734]_  & \new_[46721]_ ;
  assign \new_[2104]_  = \new_[46710]_  & \new_[46697]_ ;
  assign \new_[2105]_  = \new_[46686]_  & \new_[46673]_ ;
  assign \new_[2106]_  = \new_[46662]_  & \new_[46649]_ ;
  assign \new_[2107]_  = \new_[46638]_  & \new_[46625]_ ;
  assign \new_[2108]_  = \new_[46614]_  & \new_[46601]_ ;
  assign \new_[2109]_  = \new_[46590]_  & \new_[46577]_ ;
  assign \new_[2110]_  = \new_[46566]_  & \new_[46553]_ ;
  assign \new_[2111]_  = \new_[46542]_  & \new_[46529]_ ;
  assign \new_[2112]_  = \new_[46518]_  & \new_[46505]_ ;
  assign \new_[2113]_  = \new_[46494]_  & \new_[46481]_ ;
  assign \new_[2114]_  = \new_[46470]_  & \new_[46457]_ ;
  assign \new_[2115]_  = \new_[46446]_  & \new_[46433]_ ;
  assign \new_[2116]_  = \new_[46422]_  & \new_[46409]_ ;
  assign \new_[2117]_  = \new_[46398]_  & \new_[46385]_ ;
  assign \new_[2118]_  = \new_[46374]_  & \new_[46361]_ ;
  assign \new_[2119]_  = \new_[46350]_  & \new_[46337]_ ;
  assign \new_[2120]_  = \new_[46326]_  & \new_[46313]_ ;
  assign \new_[2121]_  = \new_[46302]_  & \new_[46289]_ ;
  assign \new_[2122]_  = \new_[46278]_  & \new_[46265]_ ;
  assign \new_[2123]_  = \new_[46254]_  & \new_[46241]_ ;
  assign \new_[2124]_  = \new_[46230]_  & \new_[46217]_ ;
  assign \new_[2125]_  = \new_[46206]_  & \new_[46193]_ ;
  assign \new_[2126]_  = \new_[46182]_  & \new_[46169]_ ;
  assign \new_[2127]_  = \new_[46158]_  & \new_[46145]_ ;
  assign \new_[2128]_  = \new_[46134]_  & \new_[46121]_ ;
  assign \new_[2129]_  = \new_[46110]_  & \new_[46097]_ ;
  assign \new_[2130]_  = \new_[46086]_  & \new_[46073]_ ;
  assign \new_[2131]_  = \new_[46062]_  & \new_[46049]_ ;
  assign \new_[2132]_  = \new_[46038]_  & \new_[46025]_ ;
  assign \new_[2133]_  = \new_[46014]_  & \new_[46001]_ ;
  assign \new_[2134]_  = \new_[45990]_  & \new_[45977]_ ;
  assign \new_[2135]_  = \new_[45966]_  & \new_[45953]_ ;
  assign \new_[2136]_  = \new_[45942]_  & \new_[45929]_ ;
  assign \new_[2137]_  = \new_[45918]_  & \new_[45905]_ ;
  assign \new_[2138]_  = \new_[45894]_  & \new_[45881]_ ;
  assign \new_[2139]_  = \new_[45870]_  & \new_[45857]_ ;
  assign \new_[2140]_  = \new_[45846]_  & \new_[45833]_ ;
  assign \new_[2141]_  = \new_[45822]_  & \new_[45809]_ ;
  assign \new_[2142]_  = \new_[45798]_  & \new_[45785]_ ;
  assign \new_[2143]_  = \new_[45774]_  & \new_[45761]_ ;
  assign \new_[2144]_  = \new_[45750]_  & \new_[45737]_ ;
  assign \new_[2145]_  = \new_[45726]_  & \new_[45713]_ ;
  assign \new_[2146]_  = \new_[45702]_  & \new_[45689]_ ;
  assign \new_[2147]_  = \new_[45678]_  & \new_[45665]_ ;
  assign \new_[2148]_  = \new_[45654]_  & \new_[45641]_ ;
  assign \new_[2149]_  = \new_[45630]_  & \new_[45617]_ ;
  assign \new_[2150]_  = \new_[45606]_  & \new_[45593]_ ;
  assign \new_[2151]_  = \new_[45582]_  & \new_[45569]_ ;
  assign \new_[2152]_  = \new_[45558]_  & \new_[45545]_ ;
  assign \new_[2153]_  = \new_[45534]_  & \new_[45521]_ ;
  assign \new_[2154]_  = \new_[45510]_  & \new_[45497]_ ;
  assign \new_[2155]_  = \new_[45486]_  & \new_[45473]_ ;
  assign \new_[2156]_  = \new_[45462]_  & \new_[45449]_ ;
  assign \new_[2157]_  = \new_[45438]_  & \new_[45425]_ ;
  assign \new_[2158]_  = \new_[45414]_  & \new_[45401]_ ;
  assign \new_[2159]_  = \new_[45390]_  & \new_[45377]_ ;
  assign \new_[2160]_  = \new_[45366]_  & \new_[45353]_ ;
  assign \new_[2161]_  = \new_[45342]_  & \new_[45329]_ ;
  assign \new_[2162]_  = \new_[45318]_  & \new_[45305]_ ;
  assign \new_[2163]_  = \new_[45294]_  & \new_[45281]_ ;
  assign \new_[2164]_  = \new_[45270]_  & \new_[45257]_ ;
  assign \new_[2165]_  = \new_[45246]_  & \new_[45233]_ ;
  assign \new_[2166]_  = \new_[45222]_  & \new_[45209]_ ;
  assign \new_[2167]_  = \new_[45198]_  & \new_[45185]_ ;
  assign \new_[2168]_  = \new_[45174]_  & \new_[45161]_ ;
  assign \new_[2169]_  = \new_[45150]_  & \new_[45137]_ ;
  assign \new_[2170]_  = \new_[45126]_  & \new_[45113]_ ;
  assign \new_[2171]_  = \new_[45102]_  & \new_[45089]_ ;
  assign \new_[2172]_  = \new_[45078]_  & \new_[45065]_ ;
  assign \new_[2173]_  = \new_[45054]_  & \new_[45041]_ ;
  assign \new_[2174]_  = \new_[45030]_  & \new_[45017]_ ;
  assign \new_[2175]_  = \new_[45006]_  & \new_[44993]_ ;
  assign \new_[2176]_  = \new_[44982]_  & \new_[44969]_ ;
  assign \new_[2177]_  = \new_[44958]_  & \new_[44945]_ ;
  assign \new_[2178]_  = \new_[44934]_  & \new_[44921]_ ;
  assign \new_[2179]_  = \new_[44910]_  & \new_[44897]_ ;
  assign \new_[2180]_  = \new_[44886]_  & \new_[44873]_ ;
  assign \new_[2181]_  = \new_[44862]_  & \new_[44849]_ ;
  assign \new_[2182]_  = \new_[44838]_  & \new_[44825]_ ;
  assign \new_[2183]_  = \new_[44814]_  & \new_[44801]_ ;
  assign \new_[2184]_  = \new_[44790]_  & \new_[44777]_ ;
  assign \new_[2185]_  = \new_[44766]_  & \new_[44753]_ ;
  assign \new_[2186]_  = \new_[44742]_  & \new_[44729]_ ;
  assign \new_[2187]_  = \new_[44718]_  & \new_[44705]_ ;
  assign \new_[2188]_  = \new_[44694]_  & \new_[44681]_ ;
  assign \new_[2189]_  = \new_[44670]_  & \new_[44657]_ ;
  assign \new_[2190]_  = \new_[44646]_  & \new_[44633]_ ;
  assign \new_[2191]_  = \new_[44622]_  & \new_[44609]_ ;
  assign \new_[2192]_  = \new_[44598]_  & \new_[44585]_ ;
  assign \new_[2193]_  = \new_[44574]_  & \new_[44561]_ ;
  assign \new_[2194]_  = \new_[44550]_  & \new_[44537]_ ;
  assign \new_[2195]_  = \new_[44526]_  & \new_[44513]_ ;
  assign \new_[2196]_  = \new_[44502]_  & \new_[44489]_ ;
  assign \new_[2197]_  = \new_[44478]_  & \new_[44465]_ ;
  assign \new_[2198]_  = \new_[44454]_  & \new_[44441]_ ;
  assign \new_[2199]_  = \new_[44430]_  & \new_[44417]_ ;
  assign \new_[2200]_  = \new_[44406]_  & \new_[44393]_ ;
  assign \new_[2201]_  = \new_[44382]_  & \new_[44369]_ ;
  assign \new_[2202]_  = \new_[44358]_  & \new_[44345]_ ;
  assign \new_[2203]_  = \new_[44334]_  & \new_[44321]_ ;
  assign \new_[2204]_  = \new_[44310]_  & \new_[44297]_ ;
  assign \new_[2205]_  = \new_[44286]_  & \new_[44273]_ ;
  assign \new_[2206]_  = \new_[44262]_  & \new_[44249]_ ;
  assign \new_[2207]_  = \new_[44238]_  & \new_[44225]_ ;
  assign \new_[2208]_  = \new_[44214]_  & \new_[44201]_ ;
  assign \new_[2209]_  = \new_[44190]_  & \new_[44177]_ ;
  assign \new_[2210]_  = \new_[44166]_  & \new_[44153]_ ;
  assign \new_[2211]_  = \new_[44142]_  & \new_[44129]_ ;
  assign \new_[2212]_  = \new_[44118]_  & \new_[44105]_ ;
  assign \new_[2213]_  = \new_[44094]_  & \new_[44081]_ ;
  assign \new_[2214]_  = \new_[44070]_  & \new_[44057]_ ;
  assign \new_[2215]_  = \new_[44046]_  & \new_[44033]_ ;
  assign \new_[2216]_  = \new_[44022]_  & \new_[44009]_ ;
  assign \new_[2217]_  = \new_[43998]_  & \new_[43985]_ ;
  assign \new_[2218]_  = \new_[43974]_  & \new_[43961]_ ;
  assign \new_[2219]_  = \new_[43950]_  & \new_[43937]_ ;
  assign \new_[2220]_  = \new_[43926]_  & \new_[43913]_ ;
  assign \new_[2221]_  = \new_[43902]_  & \new_[43889]_ ;
  assign \new_[2222]_  = \new_[43878]_  & \new_[43865]_ ;
  assign \new_[2223]_  = \new_[43854]_  & \new_[43841]_ ;
  assign \new_[2224]_  = \new_[43830]_  & \new_[43817]_ ;
  assign \new_[2225]_  = \new_[43806]_  & \new_[43793]_ ;
  assign \new_[2226]_  = \new_[43782]_  & \new_[43769]_ ;
  assign \new_[2227]_  = \new_[43758]_  & \new_[43745]_ ;
  assign \new_[2228]_  = \new_[43734]_  & \new_[43721]_ ;
  assign \new_[2229]_  = \new_[43710]_  & \new_[43697]_ ;
  assign \new_[2230]_  = \new_[43686]_  & \new_[43673]_ ;
  assign \new_[2231]_  = \new_[43662]_  & \new_[43649]_ ;
  assign \new_[2232]_  = \new_[43638]_  & \new_[43625]_ ;
  assign \new_[2233]_  = \new_[43614]_  & \new_[43601]_ ;
  assign \new_[2234]_  = \new_[43590]_  & \new_[43577]_ ;
  assign \new_[2235]_  = \new_[43566]_  & \new_[43553]_ ;
  assign \new_[2236]_  = \new_[43542]_  & \new_[43529]_ ;
  assign \new_[2237]_  = \new_[43518]_  & \new_[43505]_ ;
  assign \new_[2238]_  = \new_[43494]_  & \new_[43481]_ ;
  assign \new_[2239]_  = \new_[43470]_  & \new_[43457]_ ;
  assign \new_[2240]_  = \new_[43446]_  & \new_[43433]_ ;
  assign \new_[2241]_  = \new_[43422]_  & \new_[43409]_ ;
  assign \new_[2242]_  = \new_[43398]_  & \new_[43385]_ ;
  assign \new_[2243]_  = \new_[43374]_  & \new_[43361]_ ;
  assign \new_[2244]_  = \new_[43350]_  & \new_[43337]_ ;
  assign \new_[2245]_  = \new_[43326]_  & \new_[43313]_ ;
  assign \new_[2246]_  = \new_[43302]_  & \new_[43289]_ ;
  assign \new_[2247]_  = \new_[43278]_  & \new_[43265]_ ;
  assign \new_[2248]_  = \new_[43254]_  & \new_[43241]_ ;
  assign \new_[2249]_  = \new_[43230]_  & \new_[43217]_ ;
  assign \new_[2250]_  = \new_[43206]_  & \new_[43193]_ ;
  assign \new_[2251]_  = \new_[43182]_  & \new_[43169]_ ;
  assign \new_[2252]_  = \new_[43158]_  & \new_[43145]_ ;
  assign \new_[2253]_  = \new_[43134]_  & \new_[43121]_ ;
  assign \new_[2254]_  = \new_[43110]_  & \new_[43097]_ ;
  assign \new_[2255]_  = \new_[43086]_  & \new_[43073]_ ;
  assign \new_[2256]_  = \new_[43062]_  & \new_[43049]_ ;
  assign \new_[2257]_  = \new_[43038]_  & \new_[43025]_ ;
  assign \new_[2258]_  = \new_[43014]_  & \new_[43001]_ ;
  assign \new_[2259]_  = \new_[42990]_  & \new_[42977]_ ;
  assign \new_[2260]_  = \new_[42966]_  & \new_[42953]_ ;
  assign \new_[2261]_  = \new_[42942]_  & \new_[42929]_ ;
  assign \new_[2262]_  = \new_[42918]_  & \new_[42905]_ ;
  assign \new_[2263]_  = \new_[42894]_  & \new_[42881]_ ;
  assign \new_[2264]_  = \new_[42870]_  & \new_[42857]_ ;
  assign \new_[2265]_  = \new_[42846]_  & \new_[42833]_ ;
  assign \new_[2266]_  = \new_[42822]_  & \new_[42809]_ ;
  assign \new_[2267]_  = \new_[42798]_  & \new_[42785]_ ;
  assign \new_[2268]_  = \new_[42774]_  & \new_[42761]_ ;
  assign \new_[2269]_  = \new_[42750]_  & \new_[42737]_ ;
  assign \new_[2270]_  = \new_[42726]_  & \new_[42713]_ ;
  assign \new_[2271]_  = \new_[42702]_  & \new_[42689]_ ;
  assign \new_[2272]_  = \new_[42678]_  & \new_[42665]_ ;
  assign \new_[2273]_  = \new_[42654]_  & \new_[42641]_ ;
  assign \new_[2274]_  = \new_[42630]_  & \new_[42617]_ ;
  assign \new_[2275]_  = \new_[42606]_  & \new_[42593]_ ;
  assign \new_[2276]_  = \new_[42582]_  & \new_[42569]_ ;
  assign \new_[2277]_  = \new_[42558]_  & \new_[42545]_ ;
  assign \new_[2278]_  = \new_[42534]_  & \new_[42521]_ ;
  assign \new_[2279]_  = \new_[42510]_  & \new_[42497]_ ;
  assign \new_[2280]_  = \new_[42486]_  & \new_[42473]_ ;
  assign \new_[2281]_  = \new_[42462]_  & \new_[42449]_ ;
  assign \new_[2282]_  = \new_[42438]_  & \new_[42425]_ ;
  assign \new_[2283]_  = \new_[42414]_  & \new_[42401]_ ;
  assign \new_[2284]_  = \new_[42390]_  & \new_[42377]_ ;
  assign \new_[2285]_  = \new_[42366]_  & \new_[42353]_ ;
  assign \new_[2286]_  = \new_[42342]_  & \new_[42329]_ ;
  assign \new_[2287]_  = \new_[42318]_  & \new_[42305]_ ;
  assign \new_[2288]_  = \new_[42294]_  & \new_[42281]_ ;
  assign \new_[2289]_  = \new_[42270]_  & \new_[42257]_ ;
  assign \new_[2290]_  = \new_[42246]_  & \new_[42233]_ ;
  assign \new_[2291]_  = \new_[42222]_  & \new_[42209]_ ;
  assign \new_[2292]_  = \new_[42198]_  & \new_[42185]_ ;
  assign \new_[2293]_  = \new_[42174]_  & \new_[42161]_ ;
  assign \new_[2294]_  = \new_[42150]_  & \new_[42137]_ ;
  assign \new_[2295]_  = \new_[42126]_  & \new_[42113]_ ;
  assign \new_[2296]_  = \new_[42102]_  & \new_[42089]_ ;
  assign \new_[2297]_  = \new_[42078]_  & \new_[42065]_ ;
  assign \new_[2298]_  = \new_[42054]_  & \new_[42041]_ ;
  assign \new_[2299]_  = \new_[42030]_  & \new_[42017]_ ;
  assign \new_[2300]_  = \new_[42006]_  & \new_[41993]_ ;
  assign \new_[2301]_  = \new_[41982]_  & \new_[41969]_ ;
  assign \new_[2302]_  = \new_[41958]_  & \new_[41945]_ ;
  assign \new_[2303]_  = \new_[41934]_  & \new_[41921]_ ;
  assign \new_[2304]_  = \new_[41910]_  & \new_[41897]_ ;
  assign \new_[2305]_  = \new_[41886]_  & \new_[41873]_ ;
  assign \new_[2306]_  = \new_[41862]_  & \new_[41849]_ ;
  assign \new_[2307]_  = \new_[41838]_  & \new_[41825]_ ;
  assign \new_[2308]_  = \new_[41814]_  & \new_[41801]_ ;
  assign \new_[2309]_  = \new_[41790]_  & \new_[41777]_ ;
  assign \new_[2310]_  = \new_[41766]_  & \new_[41753]_ ;
  assign \new_[2311]_  = \new_[41742]_  & \new_[41729]_ ;
  assign \new_[2312]_  = \new_[41718]_  & \new_[41705]_ ;
  assign \new_[2313]_  = \new_[41694]_  & \new_[41681]_ ;
  assign \new_[2314]_  = \new_[41670]_  & \new_[41657]_ ;
  assign \new_[2315]_  = \new_[41646]_  & \new_[41633]_ ;
  assign \new_[2316]_  = \new_[41622]_  & \new_[41609]_ ;
  assign \new_[2317]_  = \new_[41598]_  & \new_[41585]_ ;
  assign \new_[2318]_  = \new_[41574]_  & \new_[41561]_ ;
  assign \new_[2319]_  = \new_[41550]_  & \new_[41537]_ ;
  assign \new_[2320]_  = \new_[41526]_  & \new_[41513]_ ;
  assign \new_[2321]_  = \new_[41502]_  & \new_[41489]_ ;
  assign \new_[2322]_  = \new_[41478]_  & \new_[41465]_ ;
  assign \new_[2323]_  = \new_[41454]_  & \new_[41441]_ ;
  assign \new_[2324]_  = \new_[41430]_  & \new_[41417]_ ;
  assign \new_[2325]_  = \new_[41406]_  & \new_[41393]_ ;
  assign \new_[2326]_  = \new_[41382]_  & \new_[41369]_ ;
  assign \new_[2327]_  = \new_[41358]_  & \new_[41345]_ ;
  assign \new_[2328]_  = \new_[41334]_  & \new_[41321]_ ;
  assign \new_[2329]_  = \new_[41310]_  & \new_[41299]_ ;
  assign \new_[2330]_  = \new_[41288]_  & \new_[41277]_ ;
  assign \new_[2331]_  = \new_[41266]_  & \new_[41255]_ ;
  assign \new_[2332]_  = \new_[41244]_  & \new_[41233]_ ;
  assign \new_[2333]_  = \new_[41222]_  & \new_[41211]_ ;
  assign \new_[2334]_  = \new_[41200]_  & \new_[41189]_ ;
  assign \new_[2335]_  = \new_[41178]_  & \new_[41167]_ ;
  assign \new_[2336]_  = \new_[41156]_  & \new_[41145]_ ;
  assign \new_[2337]_  = \new_[41134]_  & \new_[41123]_ ;
  assign \new_[2338]_  = \new_[41112]_  & \new_[41101]_ ;
  assign \new_[2339]_  = \new_[41090]_  & \new_[41079]_ ;
  assign \new_[2340]_  = \new_[41068]_  & \new_[41057]_ ;
  assign \new_[2341]_  = \new_[41046]_  & \new_[41035]_ ;
  assign \new_[2342]_  = \new_[41024]_  & \new_[41013]_ ;
  assign \new_[2343]_  = \new_[41002]_  & \new_[40991]_ ;
  assign \new_[2344]_  = \new_[40980]_  & \new_[40969]_ ;
  assign \new_[2345]_  = \new_[40958]_  & \new_[40947]_ ;
  assign \new_[2346]_  = \new_[40936]_  & \new_[40925]_ ;
  assign \new_[2347]_  = \new_[40914]_  & \new_[40903]_ ;
  assign \new_[2348]_  = \new_[40892]_  & \new_[40881]_ ;
  assign \new_[2349]_  = \new_[40870]_  & \new_[40859]_ ;
  assign \new_[2350]_  = \new_[40848]_  & \new_[40837]_ ;
  assign \new_[2351]_  = \new_[40826]_  & \new_[40815]_ ;
  assign \new_[2352]_  = \new_[40804]_  & \new_[40793]_ ;
  assign \new_[2353]_  = \new_[40782]_  & \new_[40771]_ ;
  assign \new_[2354]_  = \new_[40760]_  & \new_[40749]_ ;
  assign \new_[2355]_  = \new_[40738]_  & \new_[40727]_ ;
  assign \new_[2356]_  = \new_[40716]_  & \new_[40705]_ ;
  assign \new_[2357]_  = \new_[40694]_  & \new_[40683]_ ;
  assign \new_[2358]_  = \new_[40672]_  & \new_[40661]_ ;
  assign \new_[2359]_  = \new_[40650]_  & \new_[40639]_ ;
  assign \new_[2360]_  = \new_[40628]_  & \new_[40617]_ ;
  assign \new_[2361]_  = \new_[40606]_  & \new_[40595]_ ;
  assign \new_[2362]_  = \new_[40584]_  & \new_[40573]_ ;
  assign \new_[2363]_  = \new_[40562]_  & \new_[40551]_ ;
  assign \new_[2364]_  = \new_[40540]_  & \new_[40529]_ ;
  assign \new_[2365]_  = \new_[40518]_  & \new_[40507]_ ;
  assign \new_[2366]_  = \new_[40496]_  & \new_[40485]_ ;
  assign \new_[2367]_  = \new_[40474]_  & \new_[40463]_ ;
  assign \new_[2368]_  = \new_[40452]_  & \new_[40441]_ ;
  assign \new_[2369]_  = \new_[40430]_  & \new_[40419]_ ;
  assign \new_[2370]_  = \new_[40408]_  & \new_[40397]_ ;
  assign \new_[2371]_  = \new_[40386]_  & \new_[40375]_ ;
  assign \new_[2372]_  = \new_[40364]_  & \new_[40353]_ ;
  assign \new_[2373]_  = \new_[40342]_  & \new_[40331]_ ;
  assign \new_[2374]_  = \new_[40320]_  & \new_[40309]_ ;
  assign \new_[2375]_  = \new_[40298]_  & \new_[40287]_ ;
  assign \new_[2376]_  = \new_[40276]_  & \new_[40265]_ ;
  assign \new_[2377]_  = \new_[40254]_  & \new_[40243]_ ;
  assign \new_[2378]_  = \new_[40232]_  & \new_[40221]_ ;
  assign \new_[2379]_  = \new_[40210]_  & \new_[40199]_ ;
  assign \new_[2380]_  = \new_[40188]_  & \new_[40177]_ ;
  assign \new_[2381]_  = \new_[40166]_  & \new_[40155]_ ;
  assign \new_[2382]_  = \new_[40144]_  & \new_[40133]_ ;
  assign \new_[2383]_  = \new_[40122]_  & \new_[40111]_ ;
  assign \new_[2384]_  = \new_[40100]_  & \new_[40089]_ ;
  assign \new_[2385]_  = \new_[40078]_  & \new_[40067]_ ;
  assign \new_[2386]_  = \new_[40056]_  & \new_[40045]_ ;
  assign \new_[2387]_  = \new_[40034]_  & \new_[40023]_ ;
  assign \new_[2388]_  = \new_[40012]_  & \new_[40001]_ ;
  assign \new_[2389]_  = \new_[39990]_  & \new_[39979]_ ;
  assign \new_[2390]_  = \new_[39968]_  & \new_[39957]_ ;
  assign \new_[2391]_  = \new_[39946]_  & \new_[39935]_ ;
  assign \new_[2392]_  = \new_[39924]_  & \new_[39913]_ ;
  assign \new_[2393]_  = \new_[39902]_  & \new_[39891]_ ;
  assign \new_[2394]_  = \new_[39880]_  & \new_[39869]_ ;
  assign \new_[2395]_  = \new_[39858]_  & \new_[39847]_ ;
  assign \new_[2396]_  = \new_[39836]_  & \new_[39825]_ ;
  assign \new_[2397]_  = \new_[39814]_  & \new_[39803]_ ;
  assign \new_[2398]_  = \new_[39792]_  & \new_[39781]_ ;
  assign \new_[2399]_  = \new_[39770]_  & \new_[39759]_ ;
  assign \new_[2400]_  = \new_[39748]_  & \new_[39737]_ ;
  assign \new_[2401]_  = \new_[39726]_  & \new_[39715]_ ;
  assign \new_[2402]_  = \new_[39704]_  & \new_[39693]_ ;
  assign \new_[2403]_  = \new_[39682]_  & \new_[39671]_ ;
  assign \new_[2404]_  = \new_[39660]_  & \new_[39649]_ ;
  assign \new_[2405]_  = \new_[39638]_  & \new_[39627]_ ;
  assign \new_[2406]_  = \new_[39616]_  & \new_[39605]_ ;
  assign \new_[2407]_  = \new_[39594]_  & \new_[39583]_ ;
  assign \new_[2408]_  = \new_[39572]_  & \new_[39561]_ ;
  assign \new_[2409]_  = \new_[39550]_  & \new_[39539]_ ;
  assign \new_[2410]_  = \new_[39528]_  & \new_[39517]_ ;
  assign \new_[2411]_  = \new_[39506]_  & \new_[39495]_ ;
  assign \new_[2412]_  = \new_[39484]_  & \new_[39473]_ ;
  assign \new_[2413]_  = \new_[39462]_  & \new_[39451]_ ;
  assign \new_[2414]_  = \new_[39440]_  & \new_[39429]_ ;
  assign \new_[2415]_  = \new_[39418]_  & \new_[39407]_ ;
  assign \new_[2416]_  = \new_[39396]_  & \new_[39385]_ ;
  assign \new_[2417]_  = \new_[39374]_  & \new_[39363]_ ;
  assign \new_[2418]_  = \new_[39352]_  & \new_[39341]_ ;
  assign \new_[2419]_  = \new_[39330]_  & \new_[39319]_ ;
  assign \new_[2420]_  = \new_[39308]_  & \new_[39297]_ ;
  assign \new_[2421]_  = \new_[39286]_  & \new_[39275]_ ;
  assign \new_[2422]_  = \new_[39264]_  & \new_[39253]_ ;
  assign \new_[2423]_  = \new_[39242]_  & \new_[39231]_ ;
  assign \new_[2424]_  = \new_[39220]_  & \new_[39209]_ ;
  assign \new_[2425]_  = \new_[39198]_  & \new_[39187]_ ;
  assign \new_[2426]_  = \new_[39176]_  & \new_[39165]_ ;
  assign \new_[2427]_  = \new_[39154]_  & \new_[39143]_ ;
  assign \new_[2428]_  = \new_[39132]_  & \new_[39121]_ ;
  assign \new_[2429]_  = \new_[39110]_  & \new_[39099]_ ;
  assign \new_[2430]_  = \new_[39088]_  & \new_[39077]_ ;
  assign \new_[2431]_  = \new_[39066]_  & \new_[39055]_ ;
  assign \new_[2432]_  = \new_[39044]_  & \new_[39033]_ ;
  assign \new_[2433]_  = \new_[39022]_  & \new_[39011]_ ;
  assign \new_[2434]_  = \new_[39000]_  & \new_[38989]_ ;
  assign \new_[2435]_  = \new_[38978]_  & \new_[38967]_ ;
  assign \new_[2436]_  = \new_[38956]_  & \new_[38945]_ ;
  assign \new_[2437]_  = \new_[38934]_  & \new_[38923]_ ;
  assign \new_[2438]_  = \new_[38912]_  & \new_[38901]_ ;
  assign \new_[2439]_  = \new_[38890]_  & \new_[38879]_ ;
  assign \new_[2440]_  = \new_[38868]_  & \new_[38857]_ ;
  assign \new_[2441]_  = \new_[38846]_  & \new_[38835]_ ;
  assign \new_[2442]_  = \new_[38824]_  & \new_[38813]_ ;
  assign \new_[2443]_  = \new_[38802]_  & \new_[38791]_ ;
  assign \new_[2444]_  = \new_[38780]_  & \new_[38769]_ ;
  assign \new_[2445]_  = \new_[38758]_  & \new_[38747]_ ;
  assign \new_[2446]_  = \new_[38736]_  & \new_[38725]_ ;
  assign \new_[2447]_  = \new_[38714]_  & \new_[38703]_ ;
  assign \new_[2448]_  = \new_[38692]_  & \new_[38681]_ ;
  assign \new_[2449]_  = \new_[38670]_  & \new_[38659]_ ;
  assign \new_[2450]_  = \new_[38648]_  & \new_[38637]_ ;
  assign \new_[2451]_  = \new_[38626]_  & \new_[38615]_ ;
  assign \new_[2452]_  = \new_[38604]_  & \new_[38593]_ ;
  assign \new_[2453]_  = \new_[38582]_  & \new_[38571]_ ;
  assign \new_[2454]_  = \new_[38560]_  & \new_[38549]_ ;
  assign \new_[2455]_  = \new_[38538]_  & \new_[38527]_ ;
  assign \new_[2456]_  = \new_[38516]_  & \new_[38505]_ ;
  assign \new_[2457]_  = \new_[38494]_  & \new_[38483]_ ;
  assign \new_[2458]_  = \new_[38472]_  & \new_[38461]_ ;
  assign \new_[2459]_  = \new_[38450]_  & \new_[38439]_ ;
  assign \new_[2460]_  = \new_[38428]_  & \new_[38417]_ ;
  assign \new_[2461]_  = \new_[38406]_  & \new_[38395]_ ;
  assign \new_[2462]_  = \new_[38384]_  & \new_[38373]_ ;
  assign \new_[2463]_  = \new_[38362]_  & \new_[38351]_ ;
  assign \new_[2464]_  = \new_[38340]_  & \new_[38329]_ ;
  assign \new_[2465]_  = \new_[38318]_  & \new_[38307]_ ;
  assign \new_[2466]_  = \new_[38296]_  & \new_[38285]_ ;
  assign \new_[2467]_  = \new_[38274]_  & \new_[38263]_ ;
  assign \new_[2468]_  = \new_[38252]_  & \new_[38241]_ ;
  assign \new_[2469]_  = \new_[38230]_  & \new_[38219]_ ;
  assign \new_[2470]_  = \new_[38208]_  & \new_[38197]_ ;
  assign \new_[2471]_  = \new_[38186]_  & \new_[38175]_ ;
  assign \new_[2472]_  = \new_[38164]_  & \new_[38153]_ ;
  assign \new_[2473]_  = \new_[38142]_  & \new_[38131]_ ;
  assign \new_[2474]_  = \new_[38120]_  & \new_[38109]_ ;
  assign \new_[2475]_  = \new_[38098]_  & \new_[38087]_ ;
  assign \new_[2476]_  = \new_[38076]_  & \new_[38065]_ ;
  assign \new_[2477]_  = \new_[38054]_  & \new_[38043]_ ;
  assign \new_[2478]_  = \new_[38032]_  & \new_[38021]_ ;
  assign \new_[2479]_  = \new_[38010]_  & \new_[37999]_ ;
  assign \new_[2480]_  = \new_[37988]_  & \new_[37977]_ ;
  assign \new_[2481]_  = \new_[37966]_  & \new_[37955]_ ;
  assign \new_[2482]_  = \new_[37944]_  & \new_[37933]_ ;
  assign \new_[2483]_  = \new_[37922]_  & \new_[37911]_ ;
  assign \new_[2484]_  = \new_[37900]_  & \new_[37889]_ ;
  assign \new_[2485]_  = \new_[37878]_  & \new_[37867]_ ;
  assign \new_[2486]_  = \new_[37856]_  & \new_[37845]_ ;
  assign \new_[2487]_  = \new_[37834]_  & \new_[37823]_ ;
  assign \new_[2488]_  = \new_[37812]_  & \new_[37801]_ ;
  assign \new_[2489]_  = \new_[37790]_  & \new_[37779]_ ;
  assign \new_[2490]_  = \new_[37768]_  & \new_[37757]_ ;
  assign \new_[2491]_  = \new_[37746]_  & \new_[37735]_ ;
  assign \new_[2492]_  = \new_[37724]_  & \new_[37713]_ ;
  assign \new_[2493]_  = \new_[37702]_  & \new_[37691]_ ;
  assign \new_[2494]_  = \new_[37680]_  & \new_[37669]_ ;
  assign \new_[2495]_  = \new_[37658]_  & \new_[37647]_ ;
  assign \new_[2496]_  = \new_[37636]_  & \new_[37625]_ ;
  assign \new_[2497]_  = \new_[37614]_  & \new_[37603]_ ;
  assign \new_[2498]_  = \new_[37592]_  & \new_[37581]_ ;
  assign \new_[2499]_  = \new_[37570]_  & \new_[37559]_ ;
  assign \new_[2500]_  = \new_[37548]_  & \new_[37537]_ ;
  assign \new_[2501]_  = \new_[37526]_  & \new_[37515]_ ;
  assign \new_[2502]_  = \new_[37504]_  & \new_[37493]_ ;
  assign \new_[2503]_  = \new_[37482]_  & \new_[37471]_ ;
  assign \new_[2504]_  = \new_[37460]_  & \new_[37449]_ ;
  assign \new_[2505]_  = \new_[37438]_  & \new_[37427]_ ;
  assign \new_[2506]_  = \new_[37416]_  & \new_[37405]_ ;
  assign \new_[2507]_  = \new_[37394]_  & \new_[37383]_ ;
  assign \new_[2508]_  = \new_[37372]_  & \new_[37361]_ ;
  assign \new_[2509]_  = \new_[37350]_  & \new_[37339]_ ;
  assign \new_[2510]_  = \new_[37328]_  & \new_[37317]_ ;
  assign \new_[2511]_  = \new_[37306]_  & \new_[37295]_ ;
  assign \new_[2512]_  = \new_[37284]_  & \new_[37273]_ ;
  assign \new_[2513]_  = \new_[37262]_  & \new_[37251]_ ;
  assign \new_[2514]_  = \new_[37240]_  & \new_[37229]_ ;
  assign \new_[2515]_  = \new_[37218]_  & \new_[37207]_ ;
  assign \new_[2516]_  = \new_[37196]_  & \new_[37185]_ ;
  assign \new_[2517]_  = \new_[37174]_  & \new_[37163]_ ;
  assign \new_[2518]_  = \new_[37152]_  & \new_[37141]_ ;
  assign \new_[2519]_  = \new_[37130]_  & \new_[37119]_ ;
  assign \new_[2520]_  = \new_[37108]_  & \new_[37097]_ ;
  assign \new_[2521]_  = \new_[37086]_  & \new_[37075]_ ;
  assign \new_[2522]_  = \new_[37064]_  & \new_[37053]_ ;
  assign \new_[2523]_  = \new_[37042]_  & \new_[37031]_ ;
  assign \new_[2524]_  = \new_[37020]_  & \new_[37009]_ ;
  assign \new_[2525]_  = \new_[36998]_  & \new_[36987]_ ;
  assign \new_[2526]_  = \new_[36976]_  & \new_[36965]_ ;
  assign \new_[2527]_  = \new_[36954]_  & \new_[36943]_ ;
  assign \new_[2528]_  = \new_[36932]_  & \new_[36921]_ ;
  assign \new_[2529]_  = \new_[36910]_  & \new_[36899]_ ;
  assign \new_[2530]_  = \new_[36888]_  & \new_[36877]_ ;
  assign \new_[2531]_  = \new_[36866]_  & \new_[36855]_ ;
  assign \new_[2532]_  = \new_[36844]_  & \new_[36833]_ ;
  assign \new_[2533]_  = \new_[36822]_  & \new_[36811]_ ;
  assign \new_[2534]_  = \new_[36800]_  & \new_[36789]_ ;
  assign \new_[2535]_  = \new_[36778]_  & \new_[36767]_ ;
  assign \new_[2536]_  = \new_[36756]_  & \new_[36745]_ ;
  assign \new_[2537]_  = \new_[36734]_  & \new_[36723]_ ;
  assign \new_[2538]_  = \new_[36712]_  & \new_[36701]_ ;
  assign \new_[2539]_  = \new_[36690]_  & \new_[36679]_ ;
  assign \new_[2540]_  = \new_[36668]_  & \new_[36657]_ ;
  assign \new_[2541]_  = \new_[36646]_  & \new_[36635]_ ;
  assign \new_[2542]_  = \new_[36624]_  & \new_[36613]_ ;
  assign \new_[2543]_  = \new_[36602]_  & \new_[36591]_ ;
  assign \new_[2544]_  = \new_[36580]_  & \new_[36569]_ ;
  assign \new_[2545]_  = \new_[36558]_  & \new_[36547]_ ;
  assign \new_[2546]_  = \new_[36536]_  & \new_[36525]_ ;
  assign \new_[2547]_  = \new_[36514]_  & \new_[36503]_ ;
  assign \new_[2548]_  = \new_[36492]_  & \new_[36481]_ ;
  assign \new_[2549]_  = \new_[36470]_  & \new_[36459]_ ;
  assign \new_[2550]_  = \new_[36448]_  & \new_[36437]_ ;
  assign \new_[2551]_  = \new_[36426]_  & \new_[36415]_ ;
  assign \new_[2552]_  = \new_[36404]_  & \new_[36393]_ ;
  assign \new_[2553]_  = \new_[36382]_  & \new_[36371]_ ;
  assign \new_[2554]_  = \new_[36360]_  & \new_[36349]_ ;
  assign \new_[2555]_  = \new_[36338]_  & \new_[36327]_ ;
  assign \new_[2556]_  = \new_[36316]_  & \new_[36305]_ ;
  assign \new_[2557]_  = \new_[36294]_  & \new_[36283]_ ;
  assign \new_[2558]_  = \new_[36272]_  & \new_[36261]_ ;
  assign \new_[2559]_  = \new_[36250]_  & \new_[36239]_ ;
  assign \new_[2560]_  = \new_[36228]_  & \new_[36217]_ ;
  assign \new_[2561]_  = \new_[36206]_  & \new_[36195]_ ;
  assign \new_[2562]_  = \new_[36184]_  & \new_[36173]_ ;
  assign \new_[2563]_  = \new_[36162]_  & \new_[36151]_ ;
  assign \new_[2564]_  = \new_[36140]_  & \new_[36129]_ ;
  assign \new_[2565]_  = \new_[36118]_  & \new_[36107]_ ;
  assign \new_[2566]_  = \new_[36096]_  & \new_[36085]_ ;
  assign \new_[2567]_  = \new_[36074]_  & \new_[36063]_ ;
  assign \new_[2568]_  = \new_[36052]_  & \new_[36041]_ ;
  assign \new_[2569]_  = \new_[36030]_  & \new_[36019]_ ;
  assign \new_[2570]_  = \new_[36008]_  & \new_[35997]_ ;
  assign \new_[2571]_  = \new_[35986]_  & \new_[35975]_ ;
  assign \new_[2572]_  = \new_[35964]_  & \new_[35953]_ ;
  assign \new_[2573]_  = \new_[35942]_  & \new_[35931]_ ;
  assign \new_[2574]_  = \new_[35920]_  & \new_[35909]_ ;
  assign \new_[2575]_  = \new_[35898]_  & \new_[35887]_ ;
  assign \new_[2576]_  = \new_[35876]_  & \new_[35865]_ ;
  assign \new_[2577]_  = \new_[35854]_  & \new_[35843]_ ;
  assign \new_[2578]_  = \new_[35832]_  & \new_[35821]_ ;
  assign \new_[2579]_  = \new_[35810]_  & \new_[35799]_ ;
  assign \new_[2580]_  = \new_[35788]_  & \new_[35777]_ ;
  assign \new_[2581]_  = \new_[35766]_  & \new_[35755]_ ;
  assign \new_[2582]_  = \new_[35744]_  & \new_[35733]_ ;
  assign \new_[2583]_  = \new_[35722]_  & \new_[35711]_ ;
  assign \new_[2584]_  = \new_[35700]_  & \new_[35689]_ ;
  assign \new_[2585]_  = \new_[35678]_  & \new_[35667]_ ;
  assign \new_[2586]_  = \new_[35656]_  & \new_[35645]_ ;
  assign \new_[2587]_  = \new_[35634]_  & \new_[35623]_ ;
  assign \new_[2588]_  = \new_[35612]_  & \new_[35601]_ ;
  assign \new_[2589]_  = \new_[35590]_  & \new_[35579]_ ;
  assign \new_[2590]_  = \new_[35568]_  & \new_[35557]_ ;
  assign \new_[2591]_  = \new_[35546]_  & \new_[35535]_ ;
  assign \new_[2592]_  = \new_[35524]_  & \new_[35513]_ ;
  assign \new_[2593]_  = \new_[35502]_  & \new_[35491]_ ;
  assign \new_[2594]_  = \new_[35480]_  & \new_[35469]_ ;
  assign \new_[2595]_  = \new_[35458]_  & \new_[35447]_ ;
  assign \new_[2596]_  = \new_[35436]_  & \new_[35425]_ ;
  assign \new_[2597]_  = \new_[35414]_  & \new_[35403]_ ;
  assign \new_[2598]_  = \new_[35392]_  & \new_[35381]_ ;
  assign \new_[2599]_  = \new_[35370]_  & \new_[35359]_ ;
  assign \new_[2600]_  = \new_[35348]_  & \new_[35337]_ ;
  assign \new_[2601]_  = \new_[35326]_  & \new_[35315]_ ;
  assign \new_[2602]_  = \new_[35304]_  & \new_[35293]_ ;
  assign \new_[2603]_  = \new_[35282]_  & \new_[35271]_ ;
  assign \new_[2604]_  = \new_[35260]_  & \new_[35249]_ ;
  assign \new_[2605]_  = \new_[35238]_  & \new_[35227]_ ;
  assign \new_[2606]_  = \new_[35216]_  & \new_[35205]_ ;
  assign \new_[2607]_  = \new_[35194]_  & \new_[35183]_ ;
  assign \new_[2608]_  = \new_[35172]_  & \new_[35161]_ ;
  assign \new_[2609]_  = \new_[35150]_  & \new_[35139]_ ;
  assign \new_[2610]_  = \new_[35128]_  & \new_[35117]_ ;
  assign \new_[2611]_  = \new_[35106]_  & \new_[35095]_ ;
  assign \new_[2612]_  = \new_[35084]_  & \new_[35073]_ ;
  assign \new_[2613]_  = \new_[35062]_  & \new_[35051]_ ;
  assign \new_[2614]_  = \new_[35040]_  & \new_[35029]_ ;
  assign \new_[2615]_  = \new_[35018]_  & \new_[35007]_ ;
  assign \new_[2616]_  = \new_[34996]_  & \new_[34985]_ ;
  assign \new_[2617]_  = \new_[34974]_  & \new_[34963]_ ;
  assign \new_[2618]_  = \new_[34952]_  & \new_[34941]_ ;
  assign \new_[2619]_  = \new_[34930]_  & \new_[34919]_ ;
  assign \new_[2620]_  = \new_[34908]_  & \new_[34897]_ ;
  assign \new_[2621]_  = \new_[34886]_  & \new_[34875]_ ;
  assign \new_[2622]_  = \new_[34864]_  & \new_[34853]_ ;
  assign \new_[2623]_  = \new_[34842]_  & \new_[34831]_ ;
  assign \new_[2624]_  = \new_[34820]_  & \new_[34809]_ ;
  assign \new_[2625]_  = \new_[34798]_  & \new_[34787]_ ;
  assign \new_[2626]_  = \new_[34776]_  & \new_[34765]_ ;
  assign \new_[2627]_  = \new_[34754]_  & \new_[34743]_ ;
  assign \new_[2628]_  = \new_[34732]_  & \new_[34721]_ ;
  assign \new_[2629]_  = \new_[34710]_  & \new_[34699]_ ;
  assign \new_[2630]_  = \new_[34688]_  & \new_[34677]_ ;
  assign \new_[2631]_  = \new_[34666]_  & \new_[34655]_ ;
  assign \new_[2632]_  = \new_[34644]_  & \new_[34633]_ ;
  assign \new_[2633]_  = \new_[34622]_  & \new_[34611]_ ;
  assign \new_[2634]_  = \new_[34600]_  & \new_[34589]_ ;
  assign \new_[2635]_  = \new_[34578]_  & \new_[34567]_ ;
  assign \new_[2636]_  = \new_[34556]_  & \new_[34545]_ ;
  assign \new_[2637]_  = \new_[34534]_  & \new_[34523]_ ;
  assign \new_[2638]_  = \new_[34512]_  & \new_[34501]_ ;
  assign \new_[2639]_  = \new_[34490]_  & \new_[34479]_ ;
  assign \new_[2640]_  = \new_[34468]_  & \new_[34457]_ ;
  assign \new_[2641]_  = \new_[34446]_  & \new_[34435]_ ;
  assign \new_[2642]_  = \new_[34424]_  & \new_[34413]_ ;
  assign \new_[2643]_  = \new_[34402]_  & \new_[34391]_ ;
  assign \new_[2644]_  = \new_[34380]_  & \new_[34369]_ ;
  assign \new_[2645]_  = \new_[34358]_  & \new_[34347]_ ;
  assign \new_[2646]_  = \new_[34336]_  & \new_[34325]_ ;
  assign \new_[2647]_  = \new_[34314]_  & \new_[34303]_ ;
  assign \new_[2648]_  = \new_[34292]_  & \new_[34281]_ ;
  assign \new_[2649]_  = \new_[34270]_  & \new_[34259]_ ;
  assign \new_[2650]_  = \new_[34248]_  & \new_[34237]_ ;
  assign \new_[2651]_  = \new_[34226]_  & \new_[34215]_ ;
  assign \new_[2652]_  = \new_[34204]_  & \new_[34193]_ ;
  assign \new_[2653]_  = \new_[34182]_  & \new_[34171]_ ;
  assign \new_[2654]_  = \new_[34160]_  & \new_[34149]_ ;
  assign \new_[2655]_  = \new_[34138]_  & \new_[34127]_ ;
  assign \new_[2656]_  = \new_[34116]_  & \new_[34105]_ ;
  assign \new_[2657]_  = \new_[34094]_  & \new_[34083]_ ;
  assign \new_[2658]_  = \new_[34072]_  & \new_[34061]_ ;
  assign \new_[2659]_  = \new_[34050]_  & \new_[34039]_ ;
  assign \new_[2660]_  = \new_[34028]_  & \new_[34017]_ ;
  assign \new_[2661]_  = \new_[34006]_  & \new_[33995]_ ;
  assign \new_[2662]_  = \new_[33984]_  & \new_[33973]_ ;
  assign \new_[2663]_  = \new_[33962]_  & \new_[33951]_ ;
  assign \new_[2664]_  = \new_[33940]_  & \new_[33929]_ ;
  assign \new_[2665]_  = \new_[33918]_  & \new_[33907]_ ;
  assign \new_[2666]_  = \new_[33896]_  & \new_[33885]_ ;
  assign \new_[2667]_  = \new_[33874]_  & \new_[33863]_ ;
  assign \new_[2668]_  = \new_[33852]_  & \new_[33841]_ ;
  assign \new_[2669]_  = \new_[33830]_  & \new_[33819]_ ;
  assign \new_[2670]_  = \new_[33808]_  & \new_[33797]_ ;
  assign \new_[2671]_  = \new_[33786]_  & \new_[33775]_ ;
  assign \new_[2672]_  = \new_[33764]_  & \new_[33753]_ ;
  assign \new_[2673]_  = \new_[33742]_  & \new_[33731]_ ;
  assign \new_[2674]_  = \new_[33720]_  & \new_[33709]_ ;
  assign \new_[2675]_  = \new_[33698]_  & \new_[33687]_ ;
  assign \new_[2676]_  = \new_[33676]_  & \new_[33665]_ ;
  assign \new_[2677]_  = \new_[33654]_  & \new_[33643]_ ;
  assign \new_[2678]_  = \new_[33632]_  & \new_[33621]_ ;
  assign \new_[2679]_  = \new_[33610]_  & \new_[33599]_ ;
  assign \new_[2680]_  = \new_[33588]_  & \new_[33577]_ ;
  assign \new_[2681]_  = \new_[33566]_  & \new_[33555]_ ;
  assign \new_[2682]_  = \new_[33544]_  & \new_[33533]_ ;
  assign \new_[2683]_  = \new_[33522]_  & \new_[33511]_ ;
  assign \new_[2684]_  = \new_[33500]_  & \new_[33489]_ ;
  assign \new_[2685]_  = \new_[33478]_  & \new_[33467]_ ;
  assign \new_[2686]_  = \new_[33456]_  & \new_[33445]_ ;
  assign \new_[2687]_  = \new_[33434]_  & \new_[33423]_ ;
  assign \new_[2688]_  = \new_[33412]_  & \new_[33401]_ ;
  assign \new_[2689]_  = \new_[33390]_  & \new_[33379]_ ;
  assign \new_[2690]_  = \new_[33368]_  & \new_[33357]_ ;
  assign \new_[2691]_  = \new_[33346]_  & \new_[33335]_ ;
  assign \new_[2692]_  = \new_[33324]_  & \new_[33313]_ ;
  assign \new_[2693]_  = \new_[33302]_  & \new_[33291]_ ;
  assign \new_[2694]_  = \new_[33280]_  & \new_[33269]_ ;
  assign \new_[2695]_  = \new_[33258]_  & \new_[33247]_ ;
  assign \new_[2696]_  = \new_[33236]_  & \new_[33225]_ ;
  assign \new_[2697]_  = \new_[33214]_  & \new_[33203]_ ;
  assign \new_[2698]_  = \new_[33192]_  & \new_[33181]_ ;
  assign \new_[2699]_  = \new_[33170]_  & \new_[33159]_ ;
  assign \new_[2700]_  = \new_[33148]_  & \new_[33137]_ ;
  assign \new_[2701]_  = \new_[33126]_  & \new_[33115]_ ;
  assign \new_[2702]_  = \new_[33104]_  & \new_[33093]_ ;
  assign \new_[2703]_  = \new_[33082]_  & \new_[33071]_ ;
  assign \new_[2704]_  = \new_[33060]_  & \new_[33049]_ ;
  assign \new_[2705]_  = \new_[33038]_  & \new_[33027]_ ;
  assign \new_[2706]_  = \new_[33016]_  & \new_[33005]_ ;
  assign \new_[2707]_  = \new_[32994]_  & \new_[32983]_ ;
  assign \new_[2708]_  = \new_[32972]_  & \new_[32961]_ ;
  assign \new_[2709]_  = \new_[32950]_  & \new_[32939]_ ;
  assign \new_[2710]_  = \new_[32928]_  & \new_[32917]_ ;
  assign \new_[2711]_  = \new_[32906]_  & \new_[32895]_ ;
  assign \new_[2712]_  = \new_[32884]_  & \new_[32873]_ ;
  assign \new_[2713]_  = \new_[32862]_  & \new_[32851]_ ;
  assign \new_[2714]_  = \new_[32840]_  & \new_[32829]_ ;
  assign \new_[2715]_  = \new_[32818]_  & \new_[32807]_ ;
  assign \new_[2716]_  = \new_[32796]_  & \new_[32785]_ ;
  assign \new_[2717]_  = \new_[32774]_  & \new_[32763]_ ;
  assign \new_[2718]_  = \new_[32752]_  & \new_[32741]_ ;
  assign \new_[2719]_  = \new_[32730]_  & \new_[32719]_ ;
  assign \new_[2720]_  = \new_[32708]_  & \new_[32697]_ ;
  assign \new_[2721]_  = \new_[32686]_  & \new_[32675]_ ;
  assign \new_[2722]_  = \new_[32664]_  & \new_[32653]_ ;
  assign \new_[2723]_  = \new_[32642]_  & \new_[32631]_ ;
  assign \new_[2724]_  = \new_[32620]_  & \new_[32609]_ ;
  assign \new_[2725]_  = \new_[32598]_  & \new_[32587]_ ;
  assign \new_[2726]_  = \new_[32576]_  & \new_[32565]_ ;
  assign \new_[2727]_  = \new_[32554]_  & \new_[32543]_ ;
  assign \new_[2728]_  = \new_[32532]_  & \new_[32521]_ ;
  assign \new_[2729]_  = \new_[32510]_  & \new_[32499]_ ;
  assign \new_[2730]_  = \new_[32488]_  & \new_[32477]_ ;
  assign \new_[2731]_  = \new_[32466]_  & \new_[32455]_ ;
  assign \new_[2732]_  = \new_[32444]_  & \new_[32433]_ ;
  assign \new_[2733]_  = \new_[32422]_  & \new_[32411]_ ;
  assign \new_[2734]_  = \new_[32400]_  & \new_[32389]_ ;
  assign \new_[2735]_  = \new_[32378]_  & \new_[32367]_ ;
  assign \new_[2736]_  = \new_[32356]_  & \new_[32345]_ ;
  assign \new_[2737]_  = \new_[32334]_  & \new_[32323]_ ;
  assign \new_[2738]_  = \new_[32312]_  & \new_[32301]_ ;
  assign \new_[2739]_  = \new_[32290]_  & \new_[32279]_ ;
  assign \new_[2740]_  = \new_[32268]_  & \new_[32257]_ ;
  assign \new_[2741]_  = \new_[32246]_  & \new_[32235]_ ;
  assign \new_[2742]_  = \new_[32224]_  & \new_[32213]_ ;
  assign \new_[2743]_  = \new_[32202]_  & \new_[32191]_ ;
  assign \new_[2744]_  = \new_[32180]_  & \new_[32169]_ ;
  assign \new_[2745]_  = \new_[32158]_  & \new_[32147]_ ;
  assign \new_[2746]_  = \new_[32136]_  & \new_[32125]_ ;
  assign \new_[2747]_  = \new_[32114]_  & \new_[32103]_ ;
  assign \new_[2748]_  = \new_[32092]_  & \new_[32081]_ ;
  assign \new_[2749]_  = \new_[32070]_  & \new_[32059]_ ;
  assign \new_[2750]_  = \new_[32048]_  & \new_[32037]_ ;
  assign \new_[2751]_  = \new_[32026]_  & \new_[32015]_ ;
  assign \new_[2752]_  = \new_[32004]_  & \new_[31993]_ ;
  assign \new_[2753]_  = \new_[31982]_  & \new_[31971]_ ;
  assign \new_[2754]_  = \new_[31960]_  & \new_[31949]_ ;
  assign \new_[2755]_  = \new_[31938]_  & \new_[31927]_ ;
  assign \new_[2756]_  = \new_[31916]_  & \new_[31905]_ ;
  assign \new_[2757]_  = \new_[31894]_  & \new_[31883]_ ;
  assign \new_[2758]_  = \new_[31872]_  & \new_[31861]_ ;
  assign \new_[2759]_  = \new_[31850]_  & \new_[31839]_ ;
  assign \new_[2760]_  = \new_[31828]_  & \new_[31817]_ ;
  assign \new_[2761]_  = \new_[31806]_  & \new_[31795]_ ;
  assign \new_[2762]_  = \new_[31784]_  & \new_[31773]_ ;
  assign \new_[2763]_  = \new_[31762]_  & \new_[31751]_ ;
  assign \new_[2764]_  = \new_[31740]_  & \new_[31729]_ ;
  assign \new_[2765]_  = \new_[31718]_  & \new_[31707]_ ;
  assign \new_[2766]_  = \new_[31696]_  & \new_[31685]_ ;
  assign \new_[2767]_  = \new_[31674]_  & \new_[31663]_ ;
  assign \new_[2768]_  = \new_[31652]_  & \new_[31641]_ ;
  assign \new_[2769]_  = \new_[31630]_  & \new_[31619]_ ;
  assign \new_[2770]_  = \new_[31608]_  & \new_[31597]_ ;
  assign \new_[2771]_  = \new_[31586]_  & \new_[31575]_ ;
  assign \new_[2772]_  = \new_[31564]_  & \new_[31553]_ ;
  assign \new_[2773]_  = \new_[31542]_  & \new_[31531]_ ;
  assign \new_[2774]_  = \new_[31520]_  & \new_[31509]_ ;
  assign \new_[2775]_  = \new_[31498]_  & \new_[31487]_ ;
  assign \new_[2776]_  = \new_[31476]_  & \new_[31465]_ ;
  assign \new_[2777]_  = \new_[31454]_  & \new_[31443]_ ;
  assign \new_[2778]_  = \new_[31432]_  & \new_[31421]_ ;
  assign \new_[2779]_  = \new_[31410]_  & \new_[31399]_ ;
  assign \new_[2780]_  = \new_[31388]_  & \new_[31377]_ ;
  assign \new_[2781]_  = \new_[31366]_  & \new_[31355]_ ;
  assign \new_[2782]_  = \new_[31344]_  & \new_[31333]_ ;
  assign \new_[2783]_  = \new_[31322]_  & \new_[31311]_ ;
  assign \new_[2784]_  = \new_[31300]_  & \new_[31289]_ ;
  assign \new_[2785]_  = \new_[31278]_  & \new_[31267]_ ;
  assign \new_[2786]_  = \new_[31256]_  & \new_[31245]_ ;
  assign \new_[2787]_  = \new_[31234]_  & \new_[31223]_ ;
  assign \new_[2788]_  = \new_[31212]_  & \new_[31201]_ ;
  assign \new_[2789]_  = \new_[31190]_  & \new_[31179]_ ;
  assign \new_[2790]_  = \new_[31168]_  & \new_[31157]_ ;
  assign \new_[2791]_  = \new_[31146]_  & \new_[31135]_ ;
  assign \new_[2792]_  = \new_[31124]_  & \new_[31113]_ ;
  assign \new_[2793]_  = \new_[31102]_  & \new_[31091]_ ;
  assign \new_[2794]_  = \new_[31080]_  & \new_[31069]_ ;
  assign \new_[2795]_  = \new_[31058]_  & \new_[31047]_ ;
  assign \new_[2796]_  = \new_[31036]_  & \new_[31025]_ ;
  assign \new_[2797]_  = \new_[31014]_  & \new_[31003]_ ;
  assign \new_[2798]_  = \new_[30992]_  & \new_[30981]_ ;
  assign \new_[2799]_  = \new_[30970]_  & \new_[30959]_ ;
  assign \new_[2800]_  = \new_[30948]_  & \new_[30937]_ ;
  assign \new_[2801]_  = \new_[30926]_  & \new_[30915]_ ;
  assign \new_[2802]_  = \new_[30904]_  & \new_[30893]_ ;
  assign \new_[2803]_  = \new_[30882]_  & \new_[30871]_ ;
  assign \new_[2804]_  = \new_[30860]_  & \new_[30849]_ ;
  assign \new_[2805]_  = \new_[30838]_  & \new_[30827]_ ;
  assign \new_[2806]_  = \new_[30816]_  & \new_[30805]_ ;
  assign \new_[2807]_  = \new_[30794]_  & \new_[30783]_ ;
  assign \new_[2808]_  = \new_[30772]_  & \new_[30761]_ ;
  assign \new_[2809]_  = \new_[30750]_  & \new_[30739]_ ;
  assign \new_[2810]_  = \new_[30728]_  & \new_[30717]_ ;
  assign \new_[2811]_  = \new_[30706]_  & \new_[30695]_ ;
  assign \new_[2812]_  = \new_[30684]_  & \new_[30673]_ ;
  assign \new_[2813]_  = \new_[30662]_  & \new_[30651]_ ;
  assign \new_[2814]_  = \new_[30640]_  & \new_[30629]_ ;
  assign \new_[2815]_  = \new_[30618]_  & \new_[30607]_ ;
  assign \new_[2816]_  = \new_[30596]_  & \new_[30585]_ ;
  assign \new_[2817]_  = \new_[30574]_  & \new_[30563]_ ;
  assign \new_[2818]_  = \new_[30552]_  & \new_[30541]_ ;
  assign \new_[2819]_  = \new_[30530]_  & \new_[30519]_ ;
  assign \new_[2820]_  = \new_[30508]_  & \new_[30497]_ ;
  assign \new_[2821]_  = \new_[30486]_  & \new_[30475]_ ;
  assign \new_[2822]_  = \new_[30464]_  & \new_[30453]_ ;
  assign \new_[2823]_  = \new_[30442]_  & \new_[30431]_ ;
  assign \new_[2824]_  = \new_[30420]_  & \new_[30409]_ ;
  assign \new_[2825]_  = \new_[30398]_  & \new_[30387]_ ;
  assign \new_[2826]_  = \new_[30376]_  & \new_[30365]_ ;
  assign \new_[2827]_  = \new_[30354]_  & \new_[30343]_ ;
  assign \new_[2828]_  = \new_[30332]_  & \new_[30321]_ ;
  assign \new_[2829]_  = \new_[30310]_  & \new_[30299]_ ;
  assign \new_[2830]_  = \new_[30288]_  & \new_[30277]_ ;
  assign \new_[2831]_  = \new_[30266]_  & \new_[30255]_ ;
  assign \new_[2832]_  = \new_[30244]_  & \new_[30233]_ ;
  assign \new_[2833]_  = \new_[30222]_  & \new_[30211]_ ;
  assign \new_[2834]_  = \new_[30200]_  & \new_[30189]_ ;
  assign \new_[2835]_  = \new_[30178]_  & \new_[30167]_ ;
  assign \new_[2836]_  = \new_[30156]_  & \new_[30145]_ ;
  assign \new_[2837]_  = \new_[30134]_  & \new_[30123]_ ;
  assign \new_[2838]_  = \new_[30112]_  & \new_[30101]_ ;
  assign \new_[2839]_  = \new_[30090]_  & \new_[30079]_ ;
  assign \new_[2840]_  = \new_[30068]_  & \new_[30057]_ ;
  assign \new_[2841]_  = \new_[30046]_  & \new_[30035]_ ;
  assign \new_[2842]_  = \new_[30024]_  & \new_[30013]_ ;
  assign \new_[2843]_  = \new_[30002]_  & \new_[29991]_ ;
  assign \new_[2844]_  = \new_[29980]_  & \new_[29969]_ ;
  assign \new_[2845]_  = \new_[29958]_  & \new_[29947]_ ;
  assign \new_[2846]_  = \new_[29936]_  & \new_[29925]_ ;
  assign \new_[2847]_  = \new_[29914]_  & \new_[29903]_ ;
  assign \new_[2848]_  = \new_[29892]_  & \new_[29881]_ ;
  assign \new_[2849]_  = \new_[29870]_  & \new_[29859]_ ;
  assign \new_[2850]_  = \new_[29848]_  & \new_[29837]_ ;
  assign \new_[2851]_  = \new_[29826]_  & \new_[29815]_ ;
  assign \new_[2852]_  = \new_[29804]_  & \new_[29793]_ ;
  assign \new_[2853]_  = \new_[29782]_  & \new_[29771]_ ;
  assign \new_[2854]_  = \new_[29760]_  & \new_[29749]_ ;
  assign \new_[2855]_  = \new_[29738]_  & \new_[29727]_ ;
  assign \new_[2856]_  = \new_[29716]_  & \new_[29705]_ ;
  assign \new_[2857]_  = \new_[29694]_  & \new_[29683]_ ;
  assign \new_[2858]_  = \new_[29672]_  & \new_[29661]_ ;
  assign \new_[2859]_  = \new_[29650]_  & \new_[29639]_ ;
  assign \new_[2860]_  = \new_[29628]_  & \new_[29617]_ ;
  assign \new_[2861]_  = \new_[29606]_  & \new_[29595]_ ;
  assign \new_[2862]_  = \new_[29584]_  & \new_[29573]_ ;
  assign \new_[2863]_  = \new_[29562]_  & \new_[29551]_ ;
  assign \new_[2864]_  = \new_[29540]_  & \new_[29529]_ ;
  assign \new_[2865]_  = \new_[29518]_  & \new_[29507]_ ;
  assign \new_[2866]_  = \new_[29496]_  & \new_[29485]_ ;
  assign \new_[2867]_  = \new_[29474]_  & \new_[29463]_ ;
  assign \new_[2868]_  = \new_[29452]_  & \new_[29441]_ ;
  assign \new_[2869]_  = \new_[29430]_  & \new_[29419]_ ;
  assign \new_[2870]_  = \new_[29408]_  & \new_[29397]_ ;
  assign \new_[2871]_  = \new_[29386]_  & \new_[29375]_ ;
  assign \new_[2872]_  = \new_[29364]_  & \new_[29353]_ ;
  assign \new_[2873]_  = \new_[29342]_  & \new_[29331]_ ;
  assign \new_[2874]_  = \new_[29320]_  & \new_[29309]_ ;
  assign \new_[2875]_  = \new_[29298]_  & \new_[29287]_ ;
  assign \new_[2876]_  = \new_[29276]_  & \new_[29265]_ ;
  assign \new_[2877]_  = \new_[29254]_  & \new_[29243]_ ;
  assign \new_[2878]_  = \new_[29232]_  & \new_[29221]_ ;
  assign \new_[2879]_  = \new_[29210]_  & \new_[29199]_ ;
  assign \new_[2880]_  = \new_[29188]_  & \new_[29177]_ ;
  assign \new_[2881]_  = \new_[29166]_  & \new_[29155]_ ;
  assign \new_[2882]_  = \new_[29144]_  & \new_[29133]_ ;
  assign \new_[2883]_  = \new_[29122]_  & \new_[29111]_ ;
  assign \new_[2884]_  = \new_[29100]_  & \new_[29089]_ ;
  assign \new_[2885]_  = \new_[29078]_  & \new_[29067]_ ;
  assign \new_[2886]_  = \new_[29056]_  & \new_[29045]_ ;
  assign \new_[2887]_  = \new_[29034]_  & \new_[29023]_ ;
  assign \new_[2888]_  = \new_[29012]_  & \new_[29001]_ ;
  assign \new_[2889]_  = \new_[28990]_  & \new_[28979]_ ;
  assign \new_[2890]_  = \new_[28968]_  & \new_[28957]_ ;
  assign \new_[2891]_  = \new_[28946]_  & \new_[28935]_ ;
  assign \new_[2892]_  = \new_[28924]_  & \new_[28913]_ ;
  assign \new_[2893]_  = \new_[28902]_  & \new_[28891]_ ;
  assign \new_[2894]_  = \new_[28880]_  & \new_[28869]_ ;
  assign \new_[2895]_  = \new_[28858]_  & \new_[28847]_ ;
  assign \new_[2896]_  = \new_[28836]_  & \new_[28825]_ ;
  assign \new_[2897]_  = \new_[28814]_  & \new_[28803]_ ;
  assign \new_[2898]_  = \new_[28792]_  & \new_[28781]_ ;
  assign \new_[2899]_  = \new_[28770]_  & \new_[28759]_ ;
  assign \new_[2900]_  = \new_[28748]_  & \new_[28737]_ ;
  assign \new_[2901]_  = \new_[28726]_  & \new_[28715]_ ;
  assign \new_[2902]_  = \new_[28704]_  & \new_[28693]_ ;
  assign \new_[2903]_  = \new_[28682]_  & \new_[28671]_ ;
  assign \new_[2904]_  = \new_[28660]_  & \new_[28649]_ ;
  assign \new_[2905]_  = \new_[28638]_  & \new_[28627]_ ;
  assign \new_[2906]_  = \new_[28616]_  & \new_[28605]_ ;
  assign \new_[2907]_  = \new_[28594]_  & \new_[28583]_ ;
  assign \new_[2908]_  = \new_[28572]_  & \new_[28561]_ ;
  assign \new_[2909]_  = \new_[28550]_  & \new_[28539]_ ;
  assign \new_[2910]_  = \new_[28528]_  & \new_[28517]_ ;
  assign \new_[2911]_  = \new_[28506]_  & \new_[28495]_ ;
  assign \new_[2912]_  = \new_[28484]_  & \new_[28473]_ ;
  assign \new_[2913]_  = \new_[28462]_  & \new_[28451]_ ;
  assign \new_[2914]_  = \new_[28440]_  & \new_[28429]_ ;
  assign \new_[2915]_  = \new_[28418]_  & \new_[28407]_ ;
  assign \new_[2916]_  = \new_[28396]_  & \new_[28385]_ ;
  assign \new_[2917]_  = \new_[28374]_  & \new_[28363]_ ;
  assign \new_[2918]_  = \new_[28352]_  & \new_[28341]_ ;
  assign \new_[2919]_  = \new_[28330]_  & \new_[28319]_ ;
  assign \new_[2920]_  = \new_[28308]_  & \new_[28297]_ ;
  assign \new_[2921]_  = \new_[28286]_  & \new_[28275]_ ;
  assign \new_[2922]_  = \new_[28264]_  & \new_[28253]_ ;
  assign \new_[2923]_  = \new_[28242]_  & \new_[28231]_ ;
  assign \new_[2924]_  = \new_[28220]_  & \new_[28209]_ ;
  assign \new_[2925]_  = \new_[28198]_  & \new_[28187]_ ;
  assign \new_[2926]_  = \new_[28176]_  & \new_[28165]_ ;
  assign \new_[2927]_  = \new_[28154]_  & \new_[28143]_ ;
  assign \new_[2928]_  = \new_[28132]_  & \new_[28121]_ ;
  assign \new_[2929]_  = \new_[28110]_  & \new_[28099]_ ;
  assign \new_[2930]_  = \new_[28088]_  & \new_[28077]_ ;
  assign \new_[2931]_  = \new_[28066]_  & \new_[28055]_ ;
  assign \new_[2932]_  = \new_[28044]_  & \new_[28033]_ ;
  assign \new_[2933]_  = \new_[28022]_  & \new_[28011]_ ;
  assign \new_[2934]_  = \new_[28000]_  & \new_[27989]_ ;
  assign \new_[2935]_  = \new_[27978]_  & \new_[27967]_ ;
  assign \new_[2936]_  = \new_[27956]_  & \new_[27945]_ ;
  assign \new_[2937]_  = \new_[27934]_  & \new_[27923]_ ;
  assign \new_[2938]_  = \new_[27912]_  & \new_[27901]_ ;
  assign \new_[2939]_  = \new_[27890]_  & \new_[27879]_ ;
  assign \new_[2940]_  = \new_[27868]_  & \new_[27857]_ ;
  assign \new_[2941]_  = \new_[27846]_  & \new_[27835]_ ;
  assign \new_[2942]_  = \new_[27824]_  & \new_[27813]_ ;
  assign \new_[2943]_  = \new_[27802]_  & \new_[27791]_ ;
  assign \new_[2944]_  = \new_[27780]_  & \new_[27769]_ ;
  assign \new_[2945]_  = \new_[27758]_  & \new_[27747]_ ;
  assign \new_[2946]_  = \new_[27736]_  & \new_[27725]_ ;
  assign \new_[2947]_  = \new_[27714]_  & \new_[27703]_ ;
  assign \new_[2948]_  = \new_[27692]_  & \new_[27681]_ ;
  assign \new_[2949]_  = \new_[27670]_  & \new_[27659]_ ;
  assign \new_[2950]_  = \new_[27648]_  & \new_[27637]_ ;
  assign \new_[2951]_  = \new_[27626]_  & \new_[27615]_ ;
  assign \new_[2952]_  = \new_[27604]_  & \new_[27593]_ ;
  assign \new_[2953]_  = \new_[27582]_  & \new_[27571]_ ;
  assign \new_[2954]_  = \new_[27560]_  & \new_[27549]_ ;
  assign \new_[2955]_  = \new_[27538]_  & \new_[27527]_ ;
  assign \new_[2956]_  = \new_[27516]_  & \new_[27505]_ ;
  assign \new_[2957]_  = \new_[27494]_  & \new_[27483]_ ;
  assign \new_[2958]_  = \new_[27472]_  & \new_[27461]_ ;
  assign \new_[2959]_  = \new_[27450]_  & \new_[27439]_ ;
  assign \new_[2960]_  = \new_[27428]_  & \new_[27417]_ ;
  assign \new_[2961]_  = \new_[27406]_  & \new_[27395]_ ;
  assign \new_[2962]_  = \new_[27384]_  & \new_[27373]_ ;
  assign \new_[2963]_  = \new_[27362]_  & \new_[27351]_ ;
  assign \new_[2964]_  = \new_[27340]_  & \new_[27329]_ ;
  assign \new_[2965]_  = \new_[27318]_  & \new_[27307]_ ;
  assign \new_[2966]_  = \new_[27296]_  & \new_[27285]_ ;
  assign \new_[2967]_  = \new_[27274]_  & \new_[27263]_ ;
  assign \new_[2968]_  = \new_[27252]_  & \new_[27241]_ ;
  assign \new_[2969]_  = \new_[27230]_  & \new_[27219]_ ;
  assign \new_[2970]_  = \new_[27208]_  & \new_[27197]_ ;
  assign \new_[2971]_  = \new_[27186]_  & \new_[27175]_ ;
  assign \new_[2972]_  = \new_[27164]_  & \new_[27153]_ ;
  assign \new_[2973]_  = \new_[27142]_  & \new_[27131]_ ;
  assign \new_[2974]_  = \new_[27120]_  & \new_[27109]_ ;
  assign \new_[2975]_  = \new_[27098]_  & \new_[27087]_ ;
  assign \new_[2976]_  = \new_[27076]_  & \new_[27065]_ ;
  assign \new_[2977]_  = \new_[27054]_  & \new_[27043]_ ;
  assign \new_[2978]_  = \new_[27032]_  & \new_[27021]_ ;
  assign \new_[2979]_  = \new_[27010]_  & \new_[26999]_ ;
  assign \new_[2980]_  = \new_[26988]_  & \new_[26977]_ ;
  assign \new_[2981]_  = \new_[26966]_  & \new_[26955]_ ;
  assign \new_[2982]_  = \new_[26944]_  & \new_[26933]_ ;
  assign \new_[2983]_  = \new_[26922]_  & \new_[26911]_ ;
  assign \new_[2984]_  = \new_[26900]_  & \new_[26889]_ ;
  assign \new_[2985]_  = \new_[26878]_  & \new_[26867]_ ;
  assign \new_[2986]_  = \new_[26856]_  & \new_[26845]_ ;
  assign \new_[2987]_  = \new_[26834]_  & \new_[26823]_ ;
  assign \new_[2988]_  = \new_[26812]_  & \new_[26801]_ ;
  assign \new_[2989]_  = \new_[26790]_  & \new_[26779]_ ;
  assign \new_[2990]_  = \new_[26768]_  & \new_[26757]_ ;
  assign \new_[2991]_  = \new_[26746]_  & \new_[26735]_ ;
  assign \new_[2992]_  = \new_[26724]_  & \new_[26713]_ ;
  assign \new_[2993]_  = \new_[26702]_  & \new_[26691]_ ;
  assign \new_[2994]_  = \new_[26680]_  & \new_[26669]_ ;
  assign \new_[2995]_  = \new_[26658]_  & \new_[26647]_ ;
  assign \new_[2996]_  = \new_[26636]_  & \new_[26625]_ ;
  assign \new_[2997]_  = \new_[26614]_  & \new_[26603]_ ;
  assign \new_[2998]_  = \new_[26592]_  & \new_[26581]_ ;
  assign \new_[2999]_  = \new_[26570]_  & \new_[26559]_ ;
  assign \new_[3000]_  = \new_[26548]_  & \new_[26537]_ ;
  assign \new_[3001]_  = \new_[26526]_  & \new_[26515]_ ;
  assign \new_[3002]_  = \new_[26504]_  & \new_[26493]_ ;
  assign \new_[3003]_  = \new_[26482]_  & \new_[26471]_ ;
  assign \new_[3004]_  = \new_[26460]_  & \new_[26449]_ ;
  assign \new_[3005]_  = \new_[26438]_  & \new_[26427]_ ;
  assign \new_[3006]_  = \new_[26416]_  & \new_[26405]_ ;
  assign \new_[3007]_  = \new_[26394]_  & \new_[26383]_ ;
  assign \new_[3008]_  = \new_[26372]_  & \new_[26361]_ ;
  assign \new_[3009]_  = \new_[26350]_  & \new_[26339]_ ;
  assign \new_[3010]_  = \new_[26328]_  & \new_[26317]_ ;
  assign \new_[3011]_  = \new_[26306]_  & \new_[26295]_ ;
  assign \new_[3012]_  = \new_[26284]_  & \new_[26273]_ ;
  assign \new_[3013]_  = \new_[26262]_  & \new_[26251]_ ;
  assign \new_[3014]_  = \new_[26240]_  & \new_[26229]_ ;
  assign \new_[3015]_  = \new_[26218]_  & \new_[26207]_ ;
  assign \new_[3016]_  = \new_[26196]_  & \new_[26185]_ ;
  assign \new_[3017]_  = \new_[26174]_  & \new_[26163]_ ;
  assign \new_[3018]_  = \new_[26152]_  & \new_[26141]_ ;
  assign \new_[3019]_  = \new_[26130]_  & \new_[26119]_ ;
  assign \new_[3020]_  = \new_[26108]_  & \new_[26097]_ ;
  assign \new_[3021]_  = \new_[26086]_  & \new_[26075]_ ;
  assign \new_[3022]_  = \new_[26064]_  & \new_[26053]_ ;
  assign \new_[3023]_  = \new_[26042]_  & \new_[26031]_ ;
  assign \new_[3024]_  = \new_[26020]_  & \new_[26009]_ ;
  assign \new_[3025]_  = \new_[25998]_  & \new_[25987]_ ;
  assign \new_[3026]_  = \new_[25976]_  & \new_[25965]_ ;
  assign \new_[3027]_  = \new_[25954]_  & \new_[25943]_ ;
  assign \new_[3028]_  = \new_[25932]_  & \new_[25921]_ ;
  assign \new_[3029]_  = \new_[25910]_  & \new_[25899]_ ;
  assign \new_[3030]_  = \new_[25888]_  & \new_[25877]_ ;
  assign \new_[3031]_  = \new_[25866]_  & \new_[25855]_ ;
  assign \new_[3032]_  = \new_[25844]_  & \new_[25833]_ ;
  assign \new_[3033]_  = \new_[25822]_  & \new_[25811]_ ;
  assign \new_[3034]_  = \new_[25800]_  & \new_[25789]_ ;
  assign \new_[3035]_  = \new_[25778]_  & \new_[25767]_ ;
  assign \new_[3036]_  = \new_[25756]_  & \new_[25745]_ ;
  assign \new_[3037]_  = \new_[25734]_  & \new_[25723]_ ;
  assign \new_[3038]_  = \new_[25712]_  & \new_[25701]_ ;
  assign \new_[3039]_  = \new_[25690]_  & \new_[25679]_ ;
  assign \new_[3040]_  = \new_[25668]_  & \new_[25657]_ ;
  assign \new_[3041]_  = \new_[25646]_  & \new_[25635]_ ;
  assign \new_[3042]_  = \new_[25624]_  & \new_[25613]_ ;
  assign \new_[3043]_  = \new_[25602]_  & \new_[25591]_ ;
  assign \new_[3044]_  = \new_[25580]_  & \new_[25569]_ ;
  assign \new_[3045]_  = \new_[25558]_  & \new_[25547]_ ;
  assign \new_[3046]_  = \new_[25536]_  & \new_[25525]_ ;
  assign \new_[3047]_  = \new_[25514]_  & \new_[25503]_ ;
  assign \new_[3048]_  = \new_[25492]_  & \new_[25481]_ ;
  assign \new_[3049]_  = \new_[25470]_  & \new_[25459]_ ;
  assign \new_[3050]_  = \new_[25448]_  & \new_[25437]_ ;
  assign \new_[3051]_  = \new_[25426]_  & \new_[25415]_ ;
  assign \new_[3052]_  = \new_[25404]_  & \new_[25393]_ ;
  assign \new_[3053]_  = \new_[25382]_  & \new_[25371]_ ;
  assign \new_[3054]_  = \new_[25360]_  & \new_[25349]_ ;
  assign \new_[3055]_  = \new_[25338]_  & \new_[25327]_ ;
  assign \new_[3056]_  = \new_[25316]_  & \new_[25305]_ ;
  assign \new_[3057]_  = \new_[25294]_  & \new_[25283]_ ;
  assign \new_[3058]_  = \new_[25272]_  & \new_[25261]_ ;
  assign \new_[3059]_  = \new_[25250]_  & \new_[25239]_ ;
  assign \new_[3060]_  = \new_[25228]_  & \new_[25217]_ ;
  assign \new_[3061]_  = \new_[25206]_  & \new_[25195]_ ;
  assign \new_[3062]_  = \new_[25184]_  & \new_[25173]_ ;
  assign \new_[3063]_  = \new_[25162]_  & \new_[25151]_ ;
  assign \new_[3064]_  = \new_[25140]_  & \new_[25129]_ ;
  assign \new_[3065]_  = \new_[25118]_  & \new_[25107]_ ;
  assign \new_[3066]_  = \new_[25096]_  & \new_[25085]_ ;
  assign \new_[3067]_  = \new_[25074]_  & \new_[25063]_ ;
  assign \new_[3068]_  = \new_[25052]_  & \new_[25041]_ ;
  assign \new_[3069]_  = \new_[25030]_  & \new_[25019]_ ;
  assign \new_[3070]_  = \new_[25008]_  & \new_[24997]_ ;
  assign \new_[3071]_  = \new_[24986]_  & \new_[24975]_ ;
  assign \new_[3072]_  = \new_[24964]_  & \new_[24953]_ ;
  assign \new_[3073]_  = \new_[24942]_  & \new_[24931]_ ;
  assign \new_[3074]_  = \new_[24920]_  & \new_[24909]_ ;
  assign \new_[3075]_  = \new_[24898]_  & \new_[24887]_ ;
  assign \new_[3076]_  = \new_[24876]_  & \new_[24865]_ ;
  assign \new_[3077]_  = \new_[24854]_  & \new_[24843]_ ;
  assign \new_[3078]_  = \new_[24832]_  & \new_[24821]_ ;
  assign \new_[3079]_  = \new_[24810]_  & \new_[24799]_ ;
  assign \new_[3080]_  = \new_[24788]_  & \new_[24777]_ ;
  assign \new_[3081]_  = \new_[24766]_  & \new_[24755]_ ;
  assign \new_[3082]_  = \new_[24744]_  & \new_[24733]_ ;
  assign \new_[3083]_  = \new_[24722]_  & \new_[24711]_ ;
  assign \new_[3084]_  = \new_[24700]_  & \new_[24689]_ ;
  assign \new_[3085]_  = \new_[24678]_  & \new_[24667]_ ;
  assign \new_[3086]_  = \new_[24656]_  & \new_[24645]_ ;
  assign \new_[3087]_  = \new_[24634]_  & \new_[24623]_ ;
  assign \new_[3088]_  = \new_[24612]_  & \new_[24601]_ ;
  assign \new_[3089]_  = \new_[24590]_  & \new_[24579]_ ;
  assign \new_[3090]_  = \new_[24568]_  & \new_[24557]_ ;
  assign \new_[3091]_  = \new_[24546]_  & \new_[24535]_ ;
  assign \new_[3092]_  = \new_[24524]_  & \new_[24513]_ ;
  assign \new_[3093]_  = \new_[24502]_  & \new_[24491]_ ;
  assign \new_[3094]_  = \new_[24480]_  & \new_[24469]_ ;
  assign \new_[3095]_  = \new_[24458]_  & \new_[24447]_ ;
  assign \new_[3096]_  = \new_[24436]_  & \new_[24425]_ ;
  assign \new_[3097]_  = \new_[24414]_  & \new_[24403]_ ;
  assign \new_[3098]_  = \new_[24392]_  & \new_[24381]_ ;
  assign \new_[3099]_  = \new_[24370]_  & \new_[24359]_ ;
  assign \new_[3100]_  = \new_[24348]_  & \new_[24337]_ ;
  assign \new_[3101]_  = \new_[24326]_  & \new_[24315]_ ;
  assign \new_[3102]_  = \new_[24304]_  & \new_[24293]_ ;
  assign \new_[3103]_  = \new_[24282]_  & \new_[24271]_ ;
  assign \new_[3104]_  = \new_[24260]_  & \new_[24249]_ ;
  assign \new_[3105]_  = \new_[24238]_  & \new_[24227]_ ;
  assign \new_[3106]_  = \new_[24216]_  & \new_[24205]_ ;
  assign \new_[3107]_  = \new_[24194]_  & \new_[24183]_ ;
  assign \new_[3108]_  = \new_[24172]_  & \new_[24161]_ ;
  assign \new_[3109]_  = \new_[24150]_  & \new_[24139]_ ;
  assign \new_[3110]_  = \new_[24128]_  & \new_[24117]_ ;
  assign \new_[3111]_  = \new_[24106]_  & \new_[24095]_ ;
  assign \new_[3112]_  = \new_[24084]_  & \new_[24073]_ ;
  assign \new_[3113]_  = \new_[24062]_  & \new_[24051]_ ;
  assign \new_[3114]_  = \new_[24040]_  & \new_[24029]_ ;
  assign \new_[3115]_  = \new_[24018]_  & \new_[24007]_ ;
  assign \new_[3116]_  = \new_[23996]_  & \new_[23985]_ ;
  assign \new_[3117]_  = \new_[23974]_  & \new_[23963]_ ;
  assign \new_[3118]_  = \new_[23952]_  & \new_[23941]_ ;
  assign \new_[3119]_  = \new_[23930]_  & \new_[23919]_ ;
  assign \new_[3120]_  = \new_[23908]_  & \new_[23897]_ ;
  assign \new_[3121]_  = \new_[23886]_  & \new_[23875]_ ;
  assign \new_[3122]_  = \new_[23864]_  & \new_[23853]_ ;
  assign \new_[3123]_  = \new_[23842]_  & \new_[23831]_ ;
  assign \new_[3124]_  = \new_[23820]_  & \new_[23809]_ ;
  assign \new_[3125]_  = \new_[23798]_  & \new_[23787]_ ;
  assign \new_[3126]_  = \new_[23776]_  & \new_[23765]_ ;
  assign \new_[3127]_  = \new_[23754]_  & \new_[23743]_ ;
  assign \new_[3128]_  = \new_[23732]_  & \new_[23721]_ ;
  assign \new_[3129]_  = \new_[23710]_  & \new_[23699]_ ;
  assign \new_[3130]_  = \new_[23688]_  & \new_[23677]_ ;
  assign \new_[3131]_  = \new_[23666]_  & \new_[23655]_ ;
  assign \new_[3132]_  = \new_[23644]_  & \new_[23633]_ ;
  assign \new_[3133]_  = \new_[23622]_  & \new_[23611]_ ;
  assign \new_[3134]_  = \new_[23600]_  & \new_[23589]_ ;
  assign \new_[3135]_  = \new_[23578]_  & \new_[23567]_ ;
  assign \new_[3136]_  = \new_[23556]_  & \new_[23545]_ ;
  assign \new_[3137]_  = \new_[23534]_  & \new_[23523]_ ;
  assign \new_[3138]_  = \new_[23512]_  & \new_[23501]_ ;
  assign \new_[3139]_  = \new_[23490]_  & \new_[23479]_ ;
  assign \new_[3140]_  = \new_[23468]_  & \new_[23457]_ ;
  assign \new_[3141]_  = \new_[23446]_  & \new_[23435]_ ;
  assign \new_[3142]_  = \new_[23424]_  & \new_[23413]_ ;
  assign \new_[3143]_  = \new_[23402]_  & \new_[23391]_ ;
  assign \new_[3144]_  = \new_[23380]_  & \new_[23369]_ ;
  assign \new_[3145]_  = \new_[23358]_  & \new_[23347]_ ;
  assign \new_[3146]_  = \new_[23336]_  & \new_[23325]_ ;
  assign \new_[3147]_  = \new_[23314]_  & \new_[23303]_ ;
  assign \new_[3148]_  = \new_[23292]_  & \new_[23281]_ ;
  assign \new_[3149]_  = \new_[23270]_  & \new_[23259]_ ;
  assign \new_[3150]_  = \new_[23248]_  & \new_[23237]_ ;
  assign \new_[3151]_  = \new_[23226]_  & \new_[23215]_ ;
  assign \new_[3152]_  = \new_[23204]_  & \new_[23193]_ ;
  assign \new_[3153]_  = \new_[23182]_  & \new_[23171]_ ;
  assign \new_[3154]_  = \new_[23160]_  & \new_[23149]_ ;
  assign \new_[3155]_  = \new_[23138]_  & \new_[23127]_ ;
  assign \new_[3156]_  = \new_[23116]_  & \new_[23105]_ ;
  assign \new_[3157]_  = \new_[23094]_  & \new_[23083]_ ;
  assign \new_[3158]_  = \new_[23072]_  & \new_[23061]_ ;
  assign \new_[3159]_  = \new_[23050]_  & \new_[23039]_ ;
  assign \new_[3160]_  = \new_[23028]_  & \new_[23017]_ ;
  assign \new_[3161]_  = \new_[23006]_  & \new_[22995]_ ;
  assign \new_[3162]_  = \new_[22984]_  & \new_[22973]_ ;
  assign \new_[3163]_  = \new_[22962]_  & \new_[22951]_ ;
  assign \new_[3164]_  = \new_[22940]_  & \new_[22929]_ ;
  assign \new_[3165]_  = \new_[22918]_  & \new_[22907]_ ;
  assign \new_[3166]_  = \new_[22896]_  & \new_[22885]_ ;
  assign \new_[3167]_  = \new_[22874]_  & \new_[22863]_ ;
  assign \new_[3168]_  = \new_[22852]_  & \new_[22841]_ ;
  assign \new_[3169]_  = \new_[22830]_  & \new_[22819]_ ;
  assign \new_[3170]_  = \new_[22808]_  & \new_[22797]_ ;
  assign \new_[3171]_  = \new_[22786]_  & \new_[22775]_ ;
  assign \new_[3172]_  = \new_[22764]_  & \new_[22753]_ ;
  assign \new_[3173]_  = \new_[22742]_  & \new_[22731]_ ;
  assign \new_[3174]_  = \new_[22720]_  & \new_[22709]_ ;
  assign \new_[3175]_  = \new_[22698]_  & \new_[22687]_ ;
  assign \new_[3176]_  = \new_[22676]_  & \new_[22665]_ ;
  assign \new_[3177]_  = \new_[22654]_  & \new_[22643]_ ;
  assign \new_[3178]_  = \new_[22632]_  & \new_[22621]_ ;
  assign \new_[3179]_  = \new_[22610]_  & \new_[22599]_ ;
  assign \new_[3180]_  = \new_[22588]_  & \new_[22577]_ ;
  assign \new_[3181]_  = \new_[22566]_  & \new_[22555]_ ;
  assign \new_[3182]_  = \new_[22544]_  & \new_[22533]_ ;
  assign \new_[3183]_  = \new_[22522]_  & \new_[22511]_ ;
  assign \new_[3184]_  = \new_[22500]_  & \new_[22489]_ ;
  assign \new_[3185]_  = \new_[22478]_  & \new_[22467]_ ;
  assign \new_[3186]_  = \new_[22458]_  & \new_[22447]_ ;
  assign \new_[3187]_  = \new_[22438]_  & \new_[22427]_ ;
  assign \new_[3188]_  = \new_[22418]_  & \new_[22407]_ ;
  assign \new_[3189]_  = \new_[22398]_  & \new_[22387]_ ;
  assign \new_[3190]_  = \new_[22378]_  & \new_[22367]_ ;
  assign \new_[3191]_  = \new_[22358]_  & \new_[22347]_ ;
  assign \new_[3192]_  = \new_[22338]_  & \new_[22327]_ ;
  assign \new_[3193]_  = \new_[22318]_  & \new_[22307]_ ;
  assign \new_[3194]_  = \new_[22298]_  & \new_[22287]_ ;
  assign \new_[3195]_  = \new_[22278]_  & \new_[22267]_ ;
  assign \new_[3196]_  = \new_[22258]_  & \new_[22247]_ ;
  assign \new_[3197]_  = \new_[22238]_  & \new_[22227]_ ;
  assign \new_[3198]_  = \new_[22218]_  & \new_[22207]_ ;
  assign \new_[3199]_  = \new_[22198]_  & \new_[22187]_ ;
  assign \new_[3200]_  = \new_[22178]_  & \new_[22167]_ ;
  assign \new_[3201]_  = \new_[22158]_  & \new_[22147]_ ;
  assign \new_[3202]_  = \new_[22138]_  & \new_[22127]_ ;
  assign \new_[3203]_  = \new_[22118]_  & \new_[22107]_ ;
  assign \new_[3204]_  = \new_[22098]_  & \new_[22087]_ ;
  assign \new_[3205]_  = \new_[22078]_  & \new_[22067]_ ;
  assign \new_[3206]_  = \new_[22058]_  & \new_[22047]_ ;
  assign \new_[3207]_  = \new_[22038]_  & \new_[22027]_ ;
  assign \new_[3208]_  = \new_[22018]_  & \new_[22007]_ ;
  assign \new_[3209]_  = \new_[21998]_  & \new_[21987]_ ;
  assign \new_[3210]_  = \new_[21978]_  & \new_[21967]_ ;
  assign \new_[3211]_  = \new_[21958]_  & \new_[21947]_ ;
  assign \new_[3212]_  = \new_[21938]_  & \new_[21927]_ ;
  assign \new_[3213]_  = \new_[21918]_  & \new_[21907]_ ;
  assign \new_[3214]_  = \new_[21898]_  & \new_[21887]_ ;
  assign \new_[3215]_  = \new_[21878]_  & \new_[21867]_ ;
  assign \new_[3216]_  = \new_[21858]_  & \new_[21847]_ ;
  assign \new_[3217]_  = \new_[21838]_  & \new_[21827]_ ;
  assign \new_[3218]_  = \new_[21818]_  & \new_[21807]_ ;
  assign \new_[3219]_  = \new_[21798]_  & \new_[21787]_ ;
  assign \new_[3220]_  = \new_[21778]_  & \new_[21767]_ ;
  assign \new_[3221]_  = \new_[21758]_  & \new_[21747]_ ;
  assign \new_[3222]_  = \new_[21738]_  & \new_[21727]_ ;
  assign \new_[3223]_  = \new_[21718]_  & \new_[21707]_ ;
  assign \new_[3224]_  = \new_[21698]_  & \new_[21687]_ ;
  assign \new_[3225]_  = \new_[21678]_  & \new_[21667]_ ;
  assign \new_[3226]_  = \new_[21658]_  & \new_[21647]_ ;
  assign \new_[3227]_  = \new_[21638]_  & \new_[21627]_ ;
  assign \new_[3228]_  = \new_[21618]_  & \new_[21607]_ ;
  assign \new_[3229]_  = \new_[21598]_  & \new_[21587]_ ;
  assign \new_[3230]_  = \new_[21578]_  & \new_[21567]_ ;
  assign \new_[3231]_  = \new_[21558]_  & \new_[21547]_ ;
  assign \new_[3232]_  = \new_[21538]_  & \new_[21527]_ ;
  assign \new_[3233]_  = \new_[21518]_  & \new_[21507]_ ;
  assign \new_[3234]_  = \new_[21498]_  & \new_[21487]_ ;
  assign \new_[3235]_  = \new_[21478]_  & \new_[21467]_ ;
  assign \new_[3236]_  = \new_[21458]_  & \new_[21447]_ ;
  assign \new_[3237]_  = \new_[21438]_  & \new_[21427]_ ;
  assign \new_[3238]_  = \new_[21418]_  & \new_[21407]_ ;
  assign \new_[3239]_  = \new_[21398]_  & \new_[21387]_ ;
  assign \new_[3240]_  = \new_[21378]_  & \new_[21367]_ ;
  assign \new_[3241]_  = \new_[21358]_  & \new_[21347]_ ;
  assign \new_[3242]_  = \new_[21338]_  & \new_[21327]_ ;
  assign \new_[3243]_  = \new_[21318]_  & \new_[21307]_ ;
  assign \new_[3244]_  = \new_[21298]_  & \new_[21287]_ ;
  assign \new_[3245]_  = \new_[21278]_  & \new_[21267]_ ;
  assign \new_[3246]_  = \new_[21258]_  & \new_[21247]_ ;
  assign \new_[3247]_  = \new_[21238]_  & \new_[21227]_ ;
  assign \new_[3248]_  = \new_[21218]_  & \new_[21207]_ ;
  assign \new_[3249]_  = \new_[21198]_  & \new_[21187]_ ;
  assign \new_[3250]_  = \new_[21178]_  & \new_[21167]_ ;
  assign \new_[3251]_  = \new_[21158]_  & \new_[21147]_ ;
  assign \new_[3252]_  = \new_[21138]_  & \new_[21127]_ ;
  assign \new_[3253]_  = \new_[21118]_  & \new_[21107]_ ;
  assign \new_[3254]_  = \new_[21098]_  & \new_[21087]_ ;
  assign \new_[3255]_  = \new_[21078]_  & \new_[21067]_ ;
  assign \new_[3256]_  = \new_[21058]_  & \new_[21047]_ ;
  assign \new_[3257]_  = \new_[21038]_  & \new_[21027]_ ;
  assign \new_[3258]_  = \new_[21018]_  & \new_[21007]_ ;
  assign \new_[3259]_  = \new_[20998]_  & \new_[20987]_ ;
  assign \new_[3260]_  = \new_[20978]_  & \new_[20967]_ ;
  assign \new_[3261]_  = \new_[20958]_  & \new_[20947]_ ;
  assign \new_[3262]_  = \new_[20938]_  & \new_[20927]_ ;
  assign \new_[3263]_  = \new_[20918]_  & \new_[20907]_ ;
  assign \new_[3264]_  = \new_[20898]_  & \new_[20887]_ ;
  assign \new_[3265]_  = \new_[20878]_  & \new_[20867]_ ;
  assign \new_[3266]_  = \new_[20858]_  & \new_[20847]_ ;
  assign \new_[3267]_  = \new_[20838]_  & \new_[20827]_ ;
  assign \new_[3268]_  = \new_[20818]_  & \new_[20807]_ ;
  assign \new_[3269]_  = \new_[20798]_  & \new_[20787]_ ;
  assign \new_[3270]_  = \new_[20778]_  & \new_[20767]_ ;
  assign \new_[3271]_  = \new_[20758]_  & \new_[20747]_ ;
  assign \new_[3272]_  = \new_[20738]_  & \new_[20727]_ ;
  assign \new_[3273]_  = \new_[20718]_  & \new_[20707]_ ;
  assign \new_[3274]_  = \new_[20698]_  & \new_[20687]_ ;
  assign \new_[3275]_  = \new_[20678]_  & \new_[20667]_ ;
  assign \new_[3276]_  = \new_[20658]_  & \new_[20647]_ ;
  assign \new_[3277]_  = \new_[20638]_  & \new_[20627]_ ;
  assign \new_[3278]_  = \new_[20618]_  & \new_[20607]_ ;
  assign \new_[3279]_  = \new_[20598]_  & \new_[20587]_ ;
  assign \new_[3280]_  = \new_[20578]_  & \new_[20567]_ ;
  assign \new_[3281]_  = \new_[20558]_  & \new_[20547]_ ;
  assign \new_[3282]_  = \new_[20538]_  & \new_[20527]_ ;
  assign \new_[3283]_  = \new_[20518]_  & \new_[20507]_ ;
  assign \new_[3284]_  = \new_[20498]_  & \new_[20487]_ ;
  assign \new_[3285]_  = \new_[20478]_  & \new_[20467]_ ;
  assign \new_[3286]_  = \new_[20458]_  & \new_[20447]_ ;
  assign \new_[3287]_  = \new_[20438]_  & \new_[20427]_ ;
  assign \new_[3288]_  = \new_[20418]_  & \new_[20407]_ ;
  assign \new_[3289]_  = \new_[20398]_  & \new_[20387]_ ;
  assign \new_[3290]_  = \new_[20378]_  & \new_[20367]_ ;
  assign \new_[3291]_  = \new_[20358]_  & \new_[20347]_ ;
  assign \new_[3292]_  = \new_[20338]_  & \new_[20327]_ ;
  assign \new_[3293]_  = \new_[20318]_  & \new_[20307]_ ;
  assign \new_[3294]_  = \new_[20298]_  & \new_[20287]_ ;
  assign \new_[3295]_  = \new_[20278]_  & \new_[20267]_ ;
  assign \new_[3296]_  = \new_[20258]_  & \new_[20247]_ ;
  assign \new_[3297]_  = \new_[20238]_  & \new_[20227]_ ;
  assign \new_[3298]_  = \new_[20218]_  & \new_[20207]_ ;
  assign \new_[3299]_  = \new_[20198]_  & \new_[20187]_ ;
  assign \new_[3300]_  = \new_[20178]_  & \new_[20167]_ ;
  assign \new_[3301]_  = \new_[20158]_  & \new_[20147]_ ;
  assign \new_[3302]_  = \new_[20138]_  & \new_[20127]_ ;
  assign \new_[3303]_  = \new_[20118]_  & \new_[20107]_ ;
  assign \new_[3304]_  = \new_[20098]_  & \new_[20087]_ ;
  assign \new_[3305]_  = \new_[20078]_  & \new_[20067]_ ;
  assign \new_[3306]_  = \new_[20058]_  & \new_[20047]_ ;
  assign \new_[3307]_  = \new_[20038]_  & \new_[20027]_ ;
  assign \new_[3308]_  = \new_[20018]_  & \new_[20007]_ ;
  assign \new_[3309]_  = \new_[19998]_  & \new_[19987]_ ;
  assign \new_[3310]_  = \new_[19978]_  & \new_[19967]_ ;
  assign \new_[3311]_  = \new_[19958]_  & \new_[19947]_ ;
  assign \new_[3312]_  = \new_[19938]_  & \new_[19927]_ ;
  assign \new_[3313]_  = \new_[19918]_  & \new_[19907]_ ;
  assign \new_[3314]_  = \new_[19898]_  & \new_[19887]_ ;
  assign \new_[3315]_  = \new_[19878]_  & \new_[19867]_ ;
  assign \new_[3316]_  = \new_[19858]_  & \new_[19847]_ ;
  assign \new_[3317]_  = \new_[19838]_  & \new_[19827]_ ;
  assign \new_[3318]_  = \new_[19818]_  & \new_[19807]_ ;
  assign \new_[3319]_  = \new_[19798]_  & \new_[19787]_ ;
  assign \new_[3320]_  = \new_[19778]_  & \new_[19767]_ ;
  assign \new_[3321]_  = \new_[19758]_  & \new_[19747]_ ;
  assign \new_[3322]_  = \new_[19738]_  & \new_[19727]_ ;
  assign \new_[3323]_  = \new_[19718]_  & \new_[19707]_ ;
  assign \new_[3324]_  = \new_[19698]_  & \new_[19687]_ ;
  assign \new_[3325]_  = \new_[19678]_  & \new_[19667]_ ;
  assign \new_[3326]_  = \new_[19658]_  & \new_[19647]_ ;
  assign \new_[3327]_  = \new_[19638]_  & \new_[19627]_ ;
  assign \new_[3328]_  = \new_[19618]_  & \new_[19607]_ ;
  assign \new_[3329]_  = \new_[19598]_  & \new_[19587]_ ;
  assign \new_[3330]_  = \new_[19578]_  & \new_[19567]_ ;
  assign \new_[3331]_  = \new_[19558]_  & \new_[19547]_ ;
  assign \new_[3332]_  = \new_[19538]_  & \new_[19527]_ ;
  assign \new_[3333]_  = \new_[19518]_  & \new_[19507]_ ;
  assign \new_[3334]_  = \new_[19498]_  & \new_[19487]_ ;
  assign \new_[3335]_  = \new_[19478]_  & \new_[19467]_ ;
  assign \new_[3336]_  = \new_[19458]_  & \new_[19447]_ ;
  assign \new_[3337]_  = \new_[19438]_  & \new_[19427]_ ;
  assign \new_[3338]_  = \new_[19418]_  & \new_[19407]_ ;
  assign \new_[3339]_  = \new_[19398]_  & \new_[19387]_ ;
  assign \new_[3340]_  = \new_[19378]_  & \new_[19367]_ ;
  assign \new_[3341]_  = \new_[19358]_  & \new_[19347]_ ;
  assign \new_[3342]_  = \new_[19338]_  & \new_[19327]_ ;
  assign \new_[3343]_  = \new_[19318]_  & \new_[19307]_ ;
  assign \new_[3344]_  = \new_[19298]_  & \new_[19287]_ ;
  assign \new_[3345]_  = \new_[19278]_  & \new_[19267]_ ;
  assign \new_[3346]_  = \new_[19258]_  & \new_[19247]_ ;
  assign \new_[3347]_  = \new_[19238]_  & \new_[19227]_ ;
  assign \new_[3348]_  = \new_[19218]_  & \new_[19207]_ ;
  assign \new_[3349]_  = \new_[19198]_  & \new_[19187]_ ;
  assign \new_[3350]_  = \new_[19178]_  & \new_[19167]_ ;
  assign \new_[3351]_  = \new_[19158]_  & \new_[19147]_ ;
  assign \new_[3352]_  = \new_[19138]_  & \new_[19127]_ ;
  assign \new_[3353]_  = \new_[19118]_  & \new_[19107]_ ;
  assign \new_[3354]_  = \new_[19098]_  & \new_[19087]_ ;
  assign \new_[3355]_  = \new_[19078]_  & \new_[19067]_ ;
  assign \new_[3356]_  = \new_[19058]_  & \new_[19047]_ ;
  assign \new_[3357]_  = \new_[19038]_  & \new_[19027]_ ;
  assign \new_[3358]_  = \new_[19018]_  & \new_[19007]_ ;
  assign \new_[3359]_  = \new_[18998]_  & \new_[18987]_ ;
  assign \new_[3360]_  = \new_[18978]_  & \new_[18967]_ ;
  assign \new_[3361]_  = \new_[18958]_  & \new_[18947]_ ;
  assign \new_[3362]_  = \new_[18938]_  & \new_[18927]_ ;
  assign \new_[3363]_  = \new_[18918]_  & \new_[18907]_ ;
  assign \new_[3364]_  = \new_[18898]_  & \new_[18887]_ ;
  assign \new_[3365]_  = \new_[18878]_  & \new_[18867]_ ;
  assign \new_[3366]_  = \new_[18858]_  & \new_[18847]_ ;
  assign \new_[3367]_  = \new_[18838]_  & \new_[18827]_ ;
  assign \new_[3368]_  = \new_[18818]_  & \new_[18807]_ ;
  assign \new_[3369]_  = \new_[18798]_  & \new_[18787]_ ;
  assign \new_[3370]_  = \new_[18778]_  & \new_[18767]_ ;
  assign \new_[3371]_  = \new_[18758]_  & \new_[18747]_ ;
  assign \new_[3372]_  = \new_[18738]_  & \new_[18727]_ ;
  assign \new_[3373]_  = \new_[18718]_  & \new_[18707]_ ;
  assign \new_[3374]_  = \new_[18698]_  & \new_[18687]_ ;
  assign \new_[3375]_  = \new_[18678]_  & \new_[18667]_ ;
  assign \new_[3376]_  = \new_[18658]_  & \new_[18647]_ ;
  assign \new_[3377]_  = \new_[18638]_  & \new_[18627]_ ;
  assign \new_[3378]_  = \new_[18618]_  & \new_[18607]_ ;
  assign \new_[3379]_  = \new_[18598]_  & \new_[18587]_ ;
  assign \new_[3380]_  = \new_[18578]_  & \new_[18567]_ ;
  assign \new_[3381]_  = \new_[18558]_  & \new_[18547]_ ;
  assign \new_[3382]_  = \new_[18538]_  & \new_[18527]_ ;
  assign \new_[3383]_  = \new_[18518]_  & \new_[18507]_ ;
  assign \new_[3384]_  = \new_[18498]_  & \new_[18487]_ ;
  assign \new_[3385]_  = \new_[18478]_  & \new_[18467]_ ;
  assign \new_[3386]_  = \new_[18458]_  & \new_[18447]_ ;
  assign \new_[3387]_  = \new_[18438]_  & \new_[18427]_ ;
  assign \new_[3388]_  = \new_[18418]_  & \new_[18407]_ ;
  assign \new_[3389]_  = \new_[18398]_  & \new_[18387]_ ;
  assign \new_[3390]_  = \new_[18378]_  & \new_[18367]_ ;
  assign \new_[3391]_  = \new_[18358]_  & \new_[18347]_ ;
  assign \new_[3392]_  = \new_[18338]_  & \new_[18327]_ ;
  assign \new_[3393]_  = \new_[18318]_  & \new_[18307]_ ;
  assign \new_[3394]_  = \new_[18298]_  & \new_[18287]_ ;
  assign \new_[3395]_  = \new_[18278]_  & \new_[18267]_ ;
  assign \new_[3396]_  = \new_[18258]_  & \new_[18247]_ ;
  assign \new_[3397]_  = \new_[18238]_  & \new_[18227]_ ;
  assign \new_[3398]_  = \new_[18218]_  & \new_[18207]_ ;
  assign \new_[3399]_  = \new_[18198]_  & \new_[18187]_ ;
  assign \new_[3400]_  = \new_[18178]_  & \new_[18167]_ ;
  assign \new_[3401]_  = \new_[18158]_  & \new_[18147]_ ;
  assign \new_[3402]_  = \new_[18138]_  & \new_[18127]_ ;
  assign \new_[3403]_  = \new_[18118]_  & \new_[18107]_ ;
  assign \new_[3404]_  = \new_[18098]_  & \new_[18087]_ ;
  assign \new_[3405]_  = \new_[18078]_  & \new_[18067]_ ;
  assign \new_[3406]_  = \new_[18058]_  & \new_[18047]_ ;
  assign \new_[3407]_  = \new_[18038]_  & \new_[18027]_ ;
  assign \new_[3408]_  = \new_[18018]_  & \new_[18007]_ ;
  assign \new_[3409]_  = \new_[17998]_  & \new_[17987]_ ;
  assign \new_[3410]_  = \new_[17978]_  & \new_[17967]_ ;
  assign \new_[3411]_  = \new_[17958]_  & \new_[17947]_ ;
  assign \new_[3412]_  = \new_[17938]_  & \new_[17927]_ ;
  assign \new_[3413]_  = \new_[17918]_  & \new_[17907]_ ;
  assign \new_[3414]_  = \new_[17898]_  & \new_[17887]_ ;
  assign \new_[3415]_  = \new_[17878]_  & \new_[17867]_ ;
  assign \new_[3416]_  = \new_[17858]_  & \new_[17847]_ ;
  assign \new_[3417]_  = \new_[17838]_  & \new_[17827]_ ;
  assign \new_[3418]_  = \new_[17818]_  & \new_[17807]_ ;
  assign \new_[3419]_  = \new_[17798]_  & \new_[17787]_ ;
  assign \new_[3420]_  = \new_[17778]_  & \new_[17767]_ ;
  assign \new_[3421]_  = \new_[17758]_  & \new_[17747]_ ;
  assign \new_[3422]_  = \new_[17738]_  & \new_[17727]_ ;
  assign \new_[3423]_  = \new_[17718]_  & \new_[17707]_ ;
  assign \new_[3424]_  = \new_[17698]_  & \new_[17687]_ ;
  assign \new_[3425]_  = \new_[17678]_  & \new_[17667]_ ;
  assign \new_[3426]_  = \new_[17658]_  & \new_[17647]_ ;
  assign \new_[3427]_  = \new_[17638]_  & \new_[17627]_ ;
  assign \new_[3428]_  = \new_[17618]_  & \new_[17607]_ ;
  assign \new_[3429]_  = \new_[17598]_  & \new_[17587]_ ;
  assign \new_[3430]_  = \new_[17578]_  & \new_[17567]_ ;
  assign \new_[3431]_  = \new_[17558]_  & \new_[17547]_ ;
  assign \new_[3432]_  = \new_[17538]_  & \new_[17527]_ ;
  assign \new_[3433]_  = \new_[17518]_  & \new_[17507]_ ;
  assign \new_[3434]_  = \new_[17498]_  & \new_[17487]_ ;
  assign \new_[3435]_  = \new_[17478]_  & \new_[17467]_ ;
  assign \new_[3436]_  = \new_[17458]_  & \new_[17447]_ ;
  assign \new_[3437]_  = \new_[17438]_  & \new_[17427]_ ;
  assign \new_[3438]_  = \new_[17418]_  & \new_[17407]_ ;
  assign \new_[3439]_  = \new_[17398]_  & \new_[17387]_ ;
  assign \new_[3440]_  = \new_[17378]_  & \new_[17367]_ ;
  assign \new_[3441]_  = \new_[17358]_  & \new_[17347]_ ;
  assign \new_[3442]_  = \new_[17338]_  & \new_[17327]_ ;
  assign \new_[3443]_  = \new_[17318]_  & \new_[17307]_ ;
  assign \new_[3444]_  = \new_[17298]_  & \new_[17287]_ ;
  assign \new_[3445]_  = \new_[17278]_  & \new_[17267]_ ;
  assign \new_[3446]_  = \new_[17258]_  & \new_[17247]_ ;
  assign \new_[3447]_  = \new_[17238]_  & \new_[17227]_ ;
  assign \new_[3448]_  = \new_[17218]_  & \new_[17207]_ ;
  assign \new_[3449]_  = \new_[17198]_  & \new_[17187]_ ;
  assign \new_[3450]_  = \new_[17178]_  & \new_[17167]_ ;
  assign \new_[3451]_  = \new_[17158]_  & \new_[17147]_ ;
  assign \new_[3452]_  = \new_[17138]_  & \new_[17127]_ ;
  assign \new_[3453]_  = \new_[17118]_  & \new_[17107]_ ;
  assign \new_[3454]_  = \new_[17098]_  & \new_[17087]_ ;
  assign \new_[3455]_  = \new_[17078]_  & \new_[17067]_ ;
  assign \new_[3456]_  = \new_[17058]_  & \new_[17047]_ ;
  assign \new_[3457]_  = \new_[17038]_  & \new_[17027]_ ;
  assign \new_[3458]_  = \new_[17018]_  & \new_[17007]_ ;
  assign \new_[3459]_  = \new_[16998]_  & \new_[16987]_ ;
  assign \new_[3460]_  = \new_[16978]_  & \new_[16967]_ ;
  assign \new_[3461]_  = \new_[16958]_  & \new_[16947]_ ;
  assign \new_[3462]_  = \new_[16938]_  & \new_[16927]_ ;
  assign \new_[3463]_  = \new_[16918]_  & \new_[16907]_ ;
  assign \new_[3464]_  = \new_[16898]_  & \new_[16887]_ ;
  assign \new_[3465]_  = \new_[16878]_  & \new_[16867]_ ;
  assign \new_[3466]_  = \new_[16858]_  & \new_[16847]_ ;
  assign \new_[3467]_  = \new_[16838]_  & \new_[16827]_ ;
  assign \new_[3468]_  = \new_[16818]_  & \new_[16807]_ ;
  assign \new_[3469]_  = \new_[16798]_  & \new_[16787]_ ;
  assign \new_[3470]_  = \new_[16778]_  & \new_[16767]_ ;
  assign \new_[3471]_  = \new_[16758]_  & \new_[16747]_ ;
  assign \new_[3472]_  = \new_[16738]_  & \new_[16727]_ ;
  assign \new_[3473]_  = \new_[16718]_  & \new_[16707]_ ;
  assign \new_[3474]_  = \new_[16698]_  & \new_[16687]_ ;
  assign \new_[3475]_  = \new_[16678]_  & \new_[16667]_ ;
  assign \new_[3476]_  = \new_[16658]_  & \new_[16647]_ ;
  assign \new_[3477]_  = \new_[16638]_  & \new_[16627]_ ;
  assign \new_[3478]_  = \new_[16618]_  & \new_[16607]_ ;
  assign \new_[3479]_  = \new_[16598]_  & \new_[16587]_ ;
  assign \new_[3480]_  = \new_[16578]_  & \new_[16567]_ ;
  assign \new_[3481]_  = \new_[16558]_  & \new_[16547]_ ;
  assign \new_[3482]_  = \new_[16538]_  & \new_[16527]_ ;
  assign \new_[3483]_  = \new_[16518]_  & \new_[16507]_ ;
  assign \new_[3484]_  = \new_[16498]_  & \new_[16487]_ ;
  assign \new_[3485]_  = \new_[16478]_  & \new_[16467]_ ;
  assign \new_[3486]_  = \new_[16458]_  & \new_[16447]_ ;
  assign \new_[3487]_  = \new_[16438]_  & \new_[16427]_ ;
  assign \new_[3488]_  = \new_[16418]_  & \new_[16407]_ ;
  assign \new_[3489]_  = \new_[16398]_  & \new_[16387]_ ;
  assign \new_[3490]_  = \new_[16378]_  & \new_[16367]_ ;
  assign \new_[3491]_  = \new_[16358]_  & \new_[16347]_ ;
  assign \new_[3492]_  = \new_[16338]_  & \new_[16327]_ ;
  assign \new_[3493]_  = \new_[16318]_  & \new_[16307]_ ;
  assign \new_[3494]_  = \new_[16298]_  & \new_[16287]_ ;
  assign \new_[3495]_  = \new_[16278]_  & \new_[16267]_ ;
  assign \new_[3496]_  = \new_[16258]_  & \new_[16247]_ ;
  assign \new_[3497]_  = \new_[16238]_  & \new_[16227]_ ;
  assign \new_[3498]_  = \new_[16218]_  & \new_[16207]_ ;
  assign \new_[3499]_  = \new_[16198]_  & \new_[16187]_ ;
  assign \new_[3500]_  = \new_[16178]_  & \new_[16167]_ ;
  assign \new_[3501]_  = \new_[16158]_  & \new_[16147]_ ;
  assign \new_[3502]_  = \new_[16138]_  & \new_[16127]_ ;
  assign \new_[3503]_  = \new_[16118]_  & \new_[16107]_ ;
  assign \new_[3504]_  = \new_[16098]_  & \new_[16087]_ ;
  assign \new_[3505]_  = \new_[16078]_  & \new_[16067]_ ;
  assign \new_[3506]_  = \new_[16058]_  & \new_[16047]_ ;
  assign \new_[3507]_  = \new_[16038]_  & \new_[16029]_ ;
  assign \new_[3508]_  = \new_[16020]_  & \new_[16011]_ ;
  assign \new_[3509]_  = \new_[16002]_  & \new_[15993]_ ;
  assign \new_[3510]_  = \new_[15984]_  & \new_[15975]_ ;
  assign \new_[3511]_  = \new_[15966]_  & \new_[15957]_ ;
  assign \new_[3512]_  = \new_[15948]_  & \new_[15939]_ ;
  assign \new_[3513]_  = \new_[15930]_  & \new_[15921]_ ;
  assign \new_[3514]_  = \new_[15912]_  & \new_[15903]_ ;
  assign \new_[3515]_  = \new_[15894]_  & \new_[15885]_ ;
  assign \new_[3516]_  = \new_[15876]_  & \new_[15867]_ ;
  assign \new_[3517]_  = \new_[15858]_  & \new_[15849]_ ;
  assign \new_[3518]_  = \new_[15840]_  & \new_[15831]_ ;
  assign \new_[3519]_  = \new_[15822]_  & \new_[15813]_ ;
  assign \new_[3520]_  = \new_[15804]_  & \new_[15795]_ ;
  assign \new_[3521]_  = \new_[15786]_  & \new_[15777]_ ;
  assign \new_[3522]_  = \new_[15768]_  & \new_[15759]_ ;
  assign \new_[3523]_  = \new_[15750]_  & \new_[15741]_ ;
  assign \new_[3524]_  = \new_[15732]_  & \new_[15723]_ ;
  assign \new_[3525]_  = \new_[15714]_  & \new_[15705]_ ;
  assign \new_[3526]_  = \new_[15696]_  & \new_[15687]_ ;
  assign \new_[3527]_  = \new_[15678]_  & \new_[15669]_ ;
  assign \new_[3528]_  = \new_[15660]_  & \new_[15651]_ ;
  assign \new_[3529]_  = \new_[15642]_  & \new_[15633]_ ;
  assign \new_[3530]_  = \new_[15624]_  & \new_[15615]_ ;
  assign \new_[3531]_  = \new_[15606]_  & \new_[15597]_ ;
  assign \new_[3532]_  = \new_[15588]_  & \new_[15579]_ ;
  assign \new_[3533]_  = \new_[15570]_  & \new_[15561]_ ;
  assign \new_[3534]_  = \new_[15552]_  & \new_[15543]_ ;
  assign \new_[3535]_  = \new_[15534]_  & \new_[15525]_ ;
  assign \new_[3536]_  = \new_[15516]_  & \new_[15507]_ ;
  assign \new_[3537]_  = \new_[15498]_  & \new_[15489]_ ;
  assign \new_[3538]_  = \new_[15480]_  & \new_[15471]_ ;
  assign \new_[3539]_  = \new_[15462]_  & \new_[15453]_ ;
  assign \new_[3540]_  = \new_[15444]_  & \new_[15435]_ ;
  assign \new_[3541]_  = \new_[15426]_  & \new_[15417]_ ;
  assign \new_[3542]_  = \new_[15408]_  & \new_[15399]_ ;
  assign \new_[3543]_  = \new_[15390]_  & \new_[15381]_ ;
  assign \new_[3544]_  = \new_[15372]_  & \new_[15363]_ ;
  assign \new_[3545]_  = \new_[15354]_  & \new_[15345]_ ;
  assign \new_[3546]_  = \new_[15336]_  & \new_[15327]_ ;
  assign \new_[3547]_  = \new_[15318]_  & \new_[15309]_ ;
  assign \new_[3548]_  = \new_[15300]_  & \new_[15291]_ ;
  assign \new_[3549]_  = \new_[15282]_  & \new_[15273]_ ;
  assign \new_[3550]_  = \new_[15264]_  & \new_[15255]_ ;
  assign \new_[3551]_  = \new_[15246]_  & \new_[15237]_ ;
  assign \new_[3552]_  = \new_[15228]_  & \new_[15219]_ ;
  assign \new_[3553]_  = \new_[15210]_  & \new_[15201]_ ;
  assign \new_[3554]_  = \new_[15192]_  & \new_[15183]_ ;
  assign \new_[3555]_  = \new_[15174]_  & \new_[15165]_ ;
  assign \new_[3556]_  = \new_[15156]_  & \new_[15147]_ ;
  assign \new_[3557]_  = \new_[15138]_  & \new_[15129]_ ;
  assign \new_[3558]_  = \new_[15120]_  & \new_[15111]_ ;
  assign \new_[3559]_  = \new_[15102]_  & \new_[15093]_ ;
  assign \new_[3560]_  = \new_[15084]_  & \new_[15075]_ ;
  assign \new_[3561]_  = \new_[15066]_  & \new_[15057]_ ;
  assign \new_[3562]_  = \new_[15048]_  & \new_[15039]_ ;
  assign \new_[3563]_  = \new_[15030]_  & \new_[15021]_ ;
  assign \new_[3564]_  = \new_[15012]_  & \new_[15003]_ ;
  assign \new_[3565]_  = \new_[14994]_  & \new_[14985]_ ;
  assign \new_[3566]_  = \new_[14976]_  & \new_[14967]_ ;
  assign \new_[3567]_  = \new_[14958]_  & \new_[14949]_ ;
  assign \new_[3568]_  = \new_[14940]_  & \new_[14931]_ ;
  assign \new_[3569]_  = \new_[14922]_  & \new_[14913]_ ;
  assign \new_[3570]_  = \new_[14904]_  & \new_[14895]_ ;
  assign \new_[3571]_  = \new_[14886]_  & \new_[14877]_ ;
  assign \new_[3572]_  = \new_[14868]_  & \new_[14859]_ ;
  assign \new_[3573]_  = \new_[14850]_  & \new_[14841]_ ;
  assign \new_[3574]_  = \new_[14832]_  & \new_[14823]_ ;
  assign \new_[3575]_  = \new_[14814]_  & \new_[14805]_ ;
  assign \new_[3576]_  = \new_[14796]_  & \new_[14787]_ ;
  assign \new_[3577]_  = \new_[14778]_  & \new_[14769]_ ;
  assign \new_[3578]_  = \new_[14760]_  & \new_[14751]_ ;
  assign \new_[3579]_  = \new_[14742]_  & \new_[14733]_ ;
  assign \new_[3580]_  = \new_[14724]_  & \new_[14715]_ ;
  assign \new_[3581]_  = \new_[14706]_  & \new_[14697]_ ;
  assign \new_[3582]_  = \new_[14688]_  & \new_[14679]_ ;
  assign \new_[3583]_  = \new_[14670]_  & \new_[14661]_ ;
  assign \new_[3584]_  = \new_[14652]_  & \new_[14643]_ ;
  assign \new_[3585]_  = \new_[14634]_  & \new_[14625]_ ;
  assign \new_[3586]_  = \new_[14616]_  & \new_[14607]_ ;
  assign \new_[3587]_  = \new_[14598]_  & \new_[14589]_ ;
  assign \new_[3588]_  = \new_[14580]_  & \new_[14571]_ ;
  assign \new_[3589]_  = \new_[14562]_  & \new_[14553]_ ;
  assign \new_[3590]_  = \new_[14544]_  & \new_[14535]_ ;
  assign \new_[3591]_  = \new_[14526]_  & \new_[14517]_ ;
  assign \new_[3592]_  = \new_[14508]_  & \new_[14499]_ ;
  assign \new_[3593]_  = \new_[14490]_  & \new_[14481]_ ;
  assign \new_[3594]_  = \new_[14472]_  & \new_[14463]_ ;
  assign \new_[3595]_  = \new_[14454]_  & \new_[14445]_ ;
  assign \new_[3596]_  = \new_[14436]_  & \new_[14427]_ ;
  assign \new_[3597]_  = \new_[14418]_  & \new_[14409]_ ;
  assign \new_[3598]_  = \new_[14400]_  & \new_[14391]_ ;
  assign \new_[3599]_  = \new_[14382]_  & \new_[14373]_ ;
  assign \new_[3600]_  = \new_[14364]_  & \new_[14355]_ ;
  assign \new_[3601]_  = \new_[14346]_  & \new_[14337]_ ;
  assign \new_[3602]_  = \new_[14328]_  & \new_[14319]_ ;
  assign \new_[3603]_  = \new_[14310]_  & \new_[14301]_ ;
  assign \new_[3604]_  = \new_[14292]_  & \new_[14283]_ ;
  assign \new_[3605]_  = \new_[14274]_  & \new_[14265]_ ;
  assign \new_[3606]_  = \new_[14256]_  & \new_[14247]_ ;
  assign \new_[3607]_  = \new_[14238]_  & \new_[14229]_ ;
  assign \new_[3608]_  = \new_[14220]_  & \new_[14211]_ ;
  assign \new_[3609]_  = \new_[14202]_  & \new_[14193]_ ;
  assign \new_[3610]_  = \new_[14184]_  & \new_[14175]_ ;
  assign \new_[3611]_  = \new_[14166]_  & \new_[14157]_ ;
  assign \new_[3612]_  = \new_[14148]_  & \new_[14139]_ ;
  assign \new_[3613]_  = \new_[14130]_  & \new_[14121]_ ;
  assign \new_[3614]_  = \new_[14112]_  & \new_[14103]_ ;
  assign \new_[3615]_  = \new_[14094]_  & \new_[14085]_ ;
  assign \new_[3616]_  = \new_[14076]_  & \new_[14067]_ ;
  assign \new_[3617]_  = \new_[14058]_  & \new_[14049]_ ;
  assign \new_[3618]_  = \new_[14040]_  & \new_[14031]_ ;
  assign \new_[3619]_  = \new_[14022]_  & \new_[14013]_ ;
  assign \new_[3620]_  = \new_[14004]_  & \new_[13995]_ ;
  assign \new_[3621]_  = \new_[13986]_  & \new_[13977]_ ;
  assign \new_[3622]_  = \new_[13968]_  & \new_[13959]_ ;
  assign \new_[3623]_  = \new_[13950]_  & \new_[13941]_ ;
  assign \new_[3624]_  = \new_[13932]_  & \new_[13923]_ ;
  assign \new_[3625]_  = \new_[13914]_  & \new_[13905]_ ;
  assign \new_[3626]_  = \new_[13896]_  & \new_[13887]_ ;
  assign \new_[3627]_  = \new_[13878]_  & \new_[13869]_ ;
  assign \new_[3628]_  = \new_[13860]_  & \new_[13851]_ ;
  assign \new_[3629]_  = \new_[13842]_  & \new_[13833]_ ;
  assign \new_[3630]_  = \new_[13824]_  & \new_[13815]_ ;
  assign \new_[3631]_  = \new_[13806]_  & \new_[13797]_ ;
  assign \new_[3632]_  = \new_[13788]_  & \new_[13779]_ ;
  assign \new_[3633]_  = \new_[13770]_  & \new_[13761]_ ;
  assign \new_[3634]_  = \new_[13752]_  & \new_[13743]_ ;
  assign \new_[3635]_  = \new_[13734]_  & \new_[13725]_ ;
  assign \new_[3636]_  = \new_[13716]_  & \new_[13707]_ ;
  assign \new_[3637]_  = \new_[13698]_  & \new_[13689]_ ;
  assign \new_[3638]_  = \new_[13680]_  & \new_[13671]_ ;
  assign \new_[3639]_  = \new_[13662]_  & \new_[13653]_ ;
  assign \new_[3640]_  = \new_[13644]_  & \new_[13635]_ ;
  assign \new_[3641]_  = \new_[13626]_  & \new_[13617]_ ;
  assign \new_[3642]_  = \new_[13608]_  & \new_[13599]_ ;
  assign \new_[3643]_  = \new_[13590]_  & \new_[13581]_ ;
  assign \new_[3644]_  = \new_[13572]_  & \new_[13563]_ ;
  assign \new_[3645]_  = \new_[13554]_  & \new_[13545]_ ;
  assign \new_[3646]_  = \new_[13536]_  & \new_[13527]_ ;
  assign \new_[3647]_  = \new_[13518]_  & \new_[13509]_ ;
  assign \new_[3648]_  = \new_[13500]_  & \new_[13491]_ ;
  assign \new_[3649]_  = \new_[13482]_  & \new_[13473]_ ;
  assign \new_[3650]_  = \new_[13464]_  & \new_[13455]_ ;
  assign \new_[3651]_  = \new_[13446]_  & \new_[13437]_ ;
  assign \new_[3652]_  = \new_[13428]_  & \new_[13419]_ ;
  assign \new_[3653]_  = \new_[13410]_  & \new_[13401]_ ;
  assign \new_[3654]_  = \new_[13392]_  & \new_[13383]_ ;
  assign \new_[3655]_  = \new_[13374]_  & \new_[13365]_ ;
  assign \new_[3656]_  = \new_[13356]_  & \new_[13347]_ ;
  assign \new_[3657]_  = \new_[13338]_  & \new_[13329]_ ;
  assign \new_[3658]_  = \new_[13320]_  & \new_[13311]_ ;
  assign \new_[3659]_  = \new_[13302]_  & \new_[13293]_ ;
  assign \new_[3660]_  = \new_[13284]_  & \new_[13275]_ ;
  assign \new_[3661]_  = \new_[13266]_  & \new_[13257]_ ;
  assign \new_[3662]_  = \new_[13248]_  & \new_[13239]_ ;
  assign \new_[3663]_  = \new_[13230]_  & \new_[13221]_ ;
  assign \new_[3664]_  = \new_[13212]_  & \new_[13203]_ ;
  assign \new_[3665]_  = \new_[13194]_  & \new_[13185]_ ;
  assign \new_[3666]_  = \new_[13176]_  & \new_[13167]_ ;
  assign \new_[3667]_  = \new_[13158]_  & \new_[13149]_ ;
  assign \new_[3668]_  = \new_[13140]_  & \new_[13131]_ ;
  assign \new_[3669]_  = \new_[13122]_  & \new_[13113]_ ;
  assign \new_[3670]_  = \new_[13104]_  & \new_[13095]_ ;
  assign \new_[3671]_  = \new_[13086]_  & \new_[13077]_ ;
  assign \new_[3672]_  = \new_[13068]_  & \new_[13059]_ ;
  assign \new_[3673]_  = \new_[13050]_  & \new_[13041]_ ;
  assign \new_[3674]_  = \new_[13032]_  & \new_[13023]_ ;
  assign \new_[3675]_  = \new_[13014]_  & \new_[13005]_ ;
  assign \new_[3676]_  = \new_[12996]_  & \new_[12987]_ ;
  assign \new_[3677]_  = \new_[12978]_  & \new_[12969]_ ;
  assign \new_[3678]_  = \new_[12960]_  & \new_[12951]_ ;
  assign \new_[3679]_  = \new_[12942]_  & \new_[12933]_ ;
  assign \new_[3680]_  = \new_[12924]_  & \new_[12915]_ ;
  assign \new_[3681]_  = \new_[12906]_  & \new_[12897]_ ;
  assign \new_[3682]_  = \new_[12888]_  & \new_[12879]_ ;
  assign \new_[3683]_  = \new_[12870]_  & \new_[12861]_ ;
  assign \new_[3684]_  = \new_[12852]_  & \new_[12843]_ ;
  assign \new_[3685]_  = \new_[12834]_  & \new_[12825]_ ;
  assign \new_[3686]_  = \new_[12816]_  & \new_[12807]_ ;
  assign \new_[3687]_  = \new_[12798]_  & \new_[12789]_ ;
  assign \new_[3688]_  = \new_[12780]_  & \new_[12771]_ ;
  assign \new_[3689]_  = \new_[12762]_  & \new_[12753]_ ;
  assign \new_[3690]_  = \new_[12744]_  & \new_[12735]_ ;
  assign \new_[3691]_  = \new_[12726]_  & \new_[12717]_ ;
  assign \new_[3692]_  = \new_[12708]_  & \new_[12699]_ ;
  assign \new_[3693]_  = \new_[12690]_  & \new_[12681]_ ;
  assign \new_[3694]_  = \new_[12672]_  & \new_[12663]_ ;
  assign \new_[3695]_  = \new_[12654]_  & \new_[12645]_ ;
  assign \new_[3696]_  = \new_[12636]_  & \new_[12627]_ ;
  assign \new_[3697]_  = \new_[12618]_  & \new_[12609]_ ;
  assign \new_[3698]_  = \new_[12600]_  & \new_[12591]_ ;
  assign \new_[3699]_  = \new_[12582]_  & \new_[12573]_ ;
  assign \new_[3700]_  = \new_[12564]_  & \new_[12555]_ ;
  assign \new_[3701]_  = \new_[12546]_  & \new_[12537]_ ;
  assign \new_[3702]_  = \new_[12528]_  & \new_[12519]_ ;
  assign \new_[3703]_  = \new_[12510]_  & \new_[12501]_ ;
  assign \new_[3704]_  = \new_[12492]_  & \new_[12483]_ ;
  assign \new_[3705]_  = \new_[12474]_  & \new_[12465]_ ;
  assign \new_[3706]_  = \new_[12456]_  & \new_[12447]_ ;
  assign \new_[3707]_  = \new_[12438]_  & \new_[12429]_ ;
  assign \new_[3708]_  = \new_[12420]_  & \new_[12411]_ ;
  assign \new_[3709]_  = \new_[12402]_  & \new_[12393]_ ;
  assign \new_[3710]_  = \new_[12384]_  & \new_[12375]_ ;
  assign \new_[3711]_  = \new_[12366]_  & \new_[12357]_ ;
  assign \new_[3712]_  = \new_[12348]_  & \new_[12339]_ ;
  assign \new_[3713]_  = \new_[12330]_  & \new_[12321]_ ;
  assign \new_[3714]_  = \new_[12312]_  & \new_[12303]_ ;
  assign \new_[3715]_  = \new_[12294]_  & \new_[12285]_ ;
  assign \new_[3716]_  = \new_[12276]_  & \new_[12267]_ ;
  assign \new_[3717]_  = \new_[12258]_  & \new_[12249]_ ;
  assign \new_[3718]_  = \new_[12240]_  & \new_[12231]_ ;
  assign \new_[3719]_  = \new_[12222]_  & \new_[12213]_ ;
  assign \new_[3720]_  = \new_[12204]_  & \new_[12195]_ ;
  assign \new_[3721]_  = \new_[12186]_  & \new_[12177]_ ;
  assign \new_[3722]_  = \new_[12168]_  & \new_[12159]_ ;
  assign \new_[3723]_  = \new_[12150]_  & \new_[12141]_ ;
  assign \new_[3724]_  = \new_[12132]_  & \new_[12123]_ ;
  assign \new_[3725]_  = \new_[12114]_  & \new_[12105]_ ;
  assign \new_[3726]_  = \new_[12096]_  & \new_[12087]_ ;
  assign \new_[3727]_  = \new_[12078]_  & \new_[12069]_ ;
  assign \new_[3728]_  = \new_[12060]_  & \new_[12051]_ ;
  assign \new_[3729]_  = \new_[12042]_  & \new_[12033]_ ;
  assign \new_[3730]_  = \new_[12024]_  & \new_[12015]_ ;
  assign \new_[3731]_  = \new_[12006]_  & \new_[11997]_ ;
  assign \new_[3732]_  = \new_[11988]_  & \new_[11979]_ ;
  assign \new_[3733]_  = \new_[11970]_  & \new_[11961]_ ;
  assign \new_[3734]_  = \new_[11952]_  & \new_[11943]_ ;
  assign \new_[3735]_  = \new_[11934]_  & \new_[11925]_ ;
  assign \new_[3736]_  = \new_[11916]_  & \new_[11907]_ ;
  assign \new_[3737]_  = \new_[11898]_  & \new_[11889]_ ;
  assign \new_[3738]_  = \new_[11880]_  & \new_[11871]_ ;
  assign \new_[3739]_  = \new_[11862]_  & \new_[11853]_ ;
  assign \new_[3740]_  = \new_[11844]_  & \new_[11835]_ ;
  assign \new_[3741]_  = \new_[11826]_  & \new_[11817]_ ;
  assign \new_[3742]_  = \new_[11808]_  & \new_[11799]_ ;
  assign \new_[3743]_  = \new_[11790]_  & \new_[11781]_ ;
  assign \new_[3744]_  = \new_[11772]_  & \new_[11763]_ ;
  assign \new_[3745]_  = \new_[11754]_  & \new_[11745]_ ;
  assign \new_[3746]_  = \new_[11736]_  & \new_[11727]_ ;
  assign \new_[3747]_  = \new_[11718]_  & \new_[11709]_ ;
  assign \new_[3748]_  = \new_[11700]_  & \new_[11691]_ ;
  assign \new_[3749]_  = \new_[11682]_  & \new_[11673]_ ;
  assign \new_[3750]_  = \new_[11664]_  & \new_[11655]_ ;
  assign \new_[3751]_  = \new_[11646]_  & \new_[11637]_ ;
  assign \new_[3752]_  = \new_[11628]_  & \new_[11619]_ ;
  assign \new_[3753]_  = \new_[11610]_  & \new_[11601]_ ;
  assign \new_[3754]_  = \new_[11594]_  & \new_[11585]_ ;
  assign \new_[3755]_  = \new_[11578]_  & \new_[11569]_ ;
  assign \new_[3756]_  = \new_[11562]_  & \new_[11553]_ ;
  assign \new_[3757]_  = \new_[11546]_  & \new_[11537]_ ;
  assign \new_[3758]_  = \new_[11530]_  & \new_[11521]_ ;
  assign \new_[3759]_  = \new_[11514]_  & \new_[11505]_ ;
  assign \new_[3760]_  = \new_[11498]_  & \new_[11489]_ ;
  assign \new_[3761]_  = \new_[11482]_  & \new_[11475]_ ;
  assign \new_[3762]_  = \new_[11468]_  & \new_[11461]_ ;
  assign \new_[3763]_  = \new_[11454]_  & \new_[11447]_ ;
  assign \new_[3764]_  = \new_[11440]_  & \new_[11433]_ ;
  assign \new_[3765]_  = \new_[11426]_  & \new_[11419]_ ;
  assign \new_[3766]_  = \new_[11412]_  & \new_[11405]_ ;
  assign \new_[3767]_  = \new_[11398]_  & \new_[11391]_ ;
  assign \new_[3768]_  = \new_[11384]_  & \new_[11377]_ ;
  assign \new_[3769]_  = \new_[11370]_  & \new_[11363]_ ;
  assign \new_[3770]_  = \new_[11356]_  & \new_[11349]_ ;
  assign \new_[3771]_  = \new_[11342]_  & \new_[11335]_ ;
  assign \new_[3772]_  = \new_[11328]_  & \new_[11321]_ ;
  assign \new_[3776]_  = \new_[3770]_  | \new_[3771]_ ;
  assign \new_[3777]_  = \new_[3772]_  | \new_[3776]_ ;
  assign \new_[3780]_  = \new_[3768]_  | \new_[3769]_ ;
  assign \new_[3783]_  = \new_[3766]_  | \new_[3767]_ ;
  assign \new_[3784]_  = \new_[3783]_  | \new_[3780]_ ;
  assign \new_[3785]_  = \new_[3784]_  | \new_[3777]_ ;
  assign \new_[3789]_  = \new_[3763]_  | \new_[3764]_ ;
  assign \new_[3790]_  = \new_[3765]_  | \new_[3789]_ ;
  assign \new_[3793]_  = \new_[3761]_  | \new_[3762]_ ;
  assign \new_[3796]_  = \new_[3759]_  | \new_[3760]_ ;
  assign \new_[3797]_  = \new_[3796]_  | \new_[3793]_ ;
  assign \new_[3798]_  = \new_[3797]_  | \new_[3790]_ ;
  assign \new_[3799]_  = \new_[3798]_  | \new_[3785]_ ;
  assign \new_[3803]_  = \new_[3756]_  | \new_[3757]_ ;
  assign \new_[3804]_  = \new_[3758]_  | \new_[3803]_ ;
  assign \new_[3807]_  = \new_[3754]_  | \new_[3755]_ ;
  assign \new_[3810]_  = \new_[3752]_  | \new_[3753]_ ;
  assign \new_[3811]_  = \new_[3810]_  | \new_[3807]_ ;
  assign \new_[3812]_  = \new_[3811]_  | \new_[3804]_ ;
  assign \new_[3815]_  = \new_[3750]_  | \new_[3751]_ ;
  assign \new_[3818]_  = \new_[3748]_  | \new_[3749]_ ;
  assign \new_[3819]_  = \new_[3818]_  | \new_[3815]_ ;
  assign \new_[3822]_  = \new_[3746]_  | \new_[3747]_ ;
  assign \new_[3825]_  = \new_[3744]_  | \new_[3745]_ ;
  assign \new_[3826]_  = \new_[3825]_  | \new_[3822]_ ;
  assign \new_[3827]_  = \new_[3826]_  | \new_[3819]_ ;
  assign \new_[3828]_  = \new_[3827]_  | \new_[3812]_ ;
  assign \new_[3829]_  = \new_[3828]_  | \new_[3799]_ ;
  assign \new_[3833]_  = \new_[3741]_  | \new_[3742]_ ;
  assign \new_[3834]_  = \new_[3743]_  | \new_[3833]_ ;
  assign \new_[3837]_  = \new_[3739]_  | \new_[3740]_ ;
  assign \new_[3840]_  = \new_[3737]_  | \new_[3738]_ ;
  assign \new_[3841]_  = \new_[3840]_  | \new_[3837]_ ;
  assign \new_[3842]_  = \new_[3841]_  | \new_[3834]_ ;
  assign \new_[3846]_  = \new_[3734]_  | \new_[3735]_ ;
  assign \new_[3847]_  = \new_[3736]_  | \new_[3846]_ ;
  assign \new_[3850]_  = \new_[3732]_  | \new_[3733]_ ;
  assign \new_[3853]_  = \new_[3730]_  | \new_[3731]_ ;
  assign \new_[3854]_  = \new_[3853]_  | \new_[3850]_ ;
  assign \new_[3855]_  = \new_[3854]_  | \new_[3847]_ ;
  assign \new_[3856]_  = \new_[3855]_  | \new_[3842]_ ;
  assign \new_[3860]_  = \new_[3727]_  | \new_[3728]_ ;
  assign \new_[3861]_  = \new_[3729]_  | \new_[3860]_ ;
  assign \new_[3864]_  = \new_[3725]_  | \new_[3726]_ ;
  assign \new_[3867]_  = \new_[3723]_  | \new_[3724]_ ;
  assign \new_[3868]_  = \new_[3867]_  | \new_[3864]_ ;
  assign \new_[3869]_  = \new_[3868]_  | \new_[3861]_ ;
  assign \new_[3872]_  = \new_[3721]_  | \new_[3722]_ ;
  assign \new_[3875]_  = \new_[3719]_  | \new_[3720]_ ;
  assign \new_[3876]_  = \new_[3875]_  | \new_[3872]_ ;
  assign \new_[3879]_  = \new_[3717]_  | \new_[3718]_ ;
  assign \new_[3882]_  = \new_[3715]_  | \new_[3716]_ ;
  assign \new_[3883]_  = \new_[3882]_  | \new_[3879]_ ;
  assign \new_[3884]_  = \new_[3883]_  | \new_[3876]_ ;
  assign \new_[3885]_  = \new_[3884]_  | \new_[3869]_ ;
  assign \new_[3886]_  = \new_[3885]_  | \new_[3856]_ ;
  assign \new_[3887]_  = \new_[3886]_  | \new_[3829]_ ;
  assign \new_[3891]_  = \new_[3712]_  | \new_[3713]_ ;
  assign \new_[3892]_  = \new_[3714]_  | \new_[3891]_ ;
  assign \new_[3895]_  = \new_[3710]_  | \new_[3711]_ ;
  assign \new_[3898]_  = \new_[3708]_  | \new_[3709]_ ;
  assign \new_[3899]_  = \new_[3898]_  | \new_[3895]_ ;
  assign \new_[3900]_  = \new_[3899]_  | \new_[3892]_ ;
  assign \new_[3904]_  = \new_[3705]_  | \new_[3706]_ ;
  assign \new_[3905]_  = \new_[3707]_  | \new_[3904]_ ;
  assign \new_[3908]_  = \new_[3703]_  | \new_[3704]_ ;
  assign \new_[3911]_  = \new_[3701]_  | \new_[3702]_ ;
  assign \new_[3912]_  = \new_[3911]_  | \new_[3908]_ ;
  assign \new_[3913]_  = \new_[3912]_  | \new_[3905]_ ;
  assign \new_[3914]_  = \new_[3913]_  | \new_[3900]_ ;
  assign \new_[3918]_  = \new_[3698]_  | \new_[3699]_ ;
  assign \new_[3919]_  = \new_[3700]_  | \new_[3918]_ ;
  assign \new_[3922]_  = \new_[3696]_  | \new_[3697]_ ;
  assign \new_[3925]_  = \new_[3694]_  | \new_[3695]_ ;
  assign \new_[3926]_  = \new_[3925]_  | \new_[3922]_ ;
  assign \new_[3927]_  = \new_[3926]_  | \new_[3919]_ ;
  assign \new_[3930]_  = \new_[3692]_  | \new_[3693]_ ;
  assign \new_[3933]_  = \new_[3690]_  | \new_[3691]_ ;
  assign \new_[3934]_  = \new_[3933]_  | \new_[3930]_ ;
  assign \new_[3937]_  = \new_[3688]_  | \new_[3689]_ ;
  assign \new_[3940]_  = \new_[3686]_  | \new_[3687]_ ;
  assign \new_[3941]_  = \new_[3940]_  | \new_[3937]_ ;
  assign \new_[3942]_  = \new_[3941]_  | \new_[3934]_ ;
  assign \new_[3943]_  = \new_[3942]_  | \new_[3927]_ ;
  assign \new_[3944]_  = \new_[3943]_  | \new_[3914]_ ;
  assign \new_[3948]_  = \new_[3683]_  | \new_[3684]_ ;
  assign \new_[3949]_  = \new_[3685]_  | \new_[3948]_ ;
  assign \new_[3952]_  = \new_[3681]_  | \new_[3682]_ ;
  assign \new_[3955]_  = \new_[3679]_  | \new_[3680]_ ;
  assign \new_[3956]_  = \new_[3955]_  | \new_[3952]_ ;
  assign \new_[3957]_  = \new_[3956]_  | \new_[3949]_ ;
  assign \new_[3960]_  = \new_[3677]_  | \new_[3678]_ ;
  assign \new_[3963]_  = \new_[3675]_  | \new_[3676]_ ;
  assign \new_[3964]_  = \new_[3963]_  | \new_[3960]_ ;
  assign \new_[3967]_  = \new_[3673]_  | \new_[3674]_ ;
  assign \new_[3970]_  = \new_[3671]_  | \new_[3672]_ ;
  assign \new_[3971]_  = \new_[3970]_  | \new_[3967]_ ;
  assign \new_[3972]_  = \new_[3971]_  | \new_[3964]_ ;
  assign \new_[3973]_  = \new_[3972]_  | \new_[3957]_ ;
  assign \new_[3977]_  = \new_[3668]_  | \new_[3669]_ ;
  assign \new_[3978]_  = \new_[3670]_  | \new_[3977]_ ;
  assign \new_[3981]_  = \new_[3666]_  | \new_[3667]_ ;
  assign \new_[3984]_  = \new_[3664]_  | \new_[3665]_ ;
  assign \new_[3985]_  = \new_[3984]_  | \new_[3981]_ ;
  assign \new_[3986]_  = \new_[3985]_  | \new_[3978]_ ;
  assign \new_[3989]_  = \new_[3662]_  | \new_[3663]_ ;
  assign \new_[3992]_  = \new_[3660]_  | \new_[3661]_ ;
  assign \new_[3993]_  = \new_[3992]_  | \new_[3989]_ ;
  assign \new_[3996]_  = \new_[3658]_  | \new_[3659]_ ;
  assign \new_[3999]_  = \new_[3656]_  | \new_[3657]_ ;
  assign \new_[4000]_  = \new_[3999]_  | \new_[3996]_ ;
  assign \new_[4001]_  = \new_[4000]_  | \new_[3993]_ ;
  assign \new_[4002]_  = \new_[4001]_  | \new_[3986]_ ;
  assign \new_[4003]_  = \new_[4002]_  | \new_[3973]_ ;
  assign \new_[4004]_  = \new_[4003]_  | \new_[3944]_ ;
  assign \new_[4005]_  = \new_[4004]_  | \new_[3887]_ ;
  assign \new_[4009]_  = \new_[3653]_  | \new_[3654]_ ;
  assign \new_[4010]_  = \new_[3655]_  | \new_[4009]_ ;
  assign \new_[4013]_  = \new_[3651]_  | \new_[3652]_ ;
  assign \new_[4016]_  = \new_[3649]_  | \new_[3650]_ ;
  assign \new_[4017]_  = \new_[4016]_  | \new_[4013]_ ;
  assign \new_[4018]_  = \new_[4017]_  | \new_[4010]_ ;
  assign \new_[4022]_  = \new_[3646]_  | \new_[3647]_ ;
  assign \new_[4023]_  = \new_[3648]_  | \new_[4022]_ ;
  assign \new_[4026]_  = \new_[3644]_  | \new_[3645]_ ;
  assign \new_[4029]_  = \new_[3642]_  | \new_[3643]_ ;
  assign \new_[4030]_  = \new_[4029]_  | \new_[4026]_ ;
  assign \new_[4031]_  = \new_[4030]_  | \new_[4023]_ ;
  assign \new_[4032]_  = \new_[4031]_  | \new_[4018]_ ;
  assign \new_[4036]_  = \new_[3639]_  | \new_[3640]_ ;
  assign \new_[4037]_  = \new_[3641]_  | \new_[4036]_ ;
  assign \new_[4040]_  = \new_[3637]_  | \new_[3638]_ ;
  assign \new_[4043]_  = \new_[3635]_  | \new_[3636]_ ;
  assign \new_[4044]_  = \new_[4043]_  | \new_[4040]_ ;
  assign \new_[4045]_  = \new_[4044]_  | \new_[4037]_ ;
  assign \new_[4048]_  = \new_[3633]_  | \new_[3634]_ ;
  assign \new_[4051]_  = \new_[3631]_  | \new_[3632]_ ;
  assign \new_[4052]_  = \new_[4051]_  | \new_[4048]_ ;
  assign \new_[4055]_  = \new_[3629]_  | \new_[3630]_ ;
  assign \new_[4058]_  = \new_[3627]_  | \new_[3628]_ ;
  assign \new_[4059]_  = \new_[4058]_  | \new_[4055]_ ;
  assign \new_[4060]_  = \new_[4059]_  | \new_[4052]_ ;
  assign \new_[4061]_  = \new_[4060]_  | \new_[4045]_ ;
  assign \new_[4062]_  = \new_[4061]_  | \new_[4032]_ ;
  assign \new_[4066]_  = \new_[3624]_  | \new_[3625]_ ;
  assign \new_[4067]_  = \new_[3626]_  | \new_[4066]_ ;
  assign \new_[4070]_  = \new_[3622]_  | \new_[3623]_ ;
  assign \new_[4073]_  = \new_[3620]_  | \new_[3621]_ ;
  assign \new_[4074]_  = \new_[4073]_  | \new_[4070]_ ;
  assign \new_[4075]_  = \new_[4074]_  | \new_[4067]_ ;
  assign \new_[4078]_  = \new_[3618]_  | \new_[3619]_ ;
  assign \new_[4081]_  = \new_[3616]_  | \new_[3617]_ ;
  assign \new_[4082]_  = \new_[4081]_  | \new_[4078]_ ;
  assign \new_[4085]_  = \new_[3614]_  | \new_[3615]_ ;
  assign \new_[4088]_  = \new_[3612]_  | \new_[3613]_ ;
  assign \new_[4089]_  = \new_[4088]_  | \new_[4085]_ ;
  assign \new_[4090]_  = \new_[4089]_  | \new_[4082]_ ;
  assign \new_[4091]_  = \new_[4090]_  | \new_[4075]_ ;
  assign \new_[4095]_  = \new_[3609]_  | \new_[3610]_ ;
  assign \new_[4096]_  = \new_[3611]_  | \new_[4095]_ ;
  assign \new_[4099]_  = \new_[3607]_  | \new_[3608]_ ;
  assign \new_[4102]_  = \new_[3605]_  | \new_[3606]_ ;
  assign \new_[4103]_  = \new_[4102]_  | \new_[4099]_ ;
  assign \new_[4104]_  = \new_[4103]_  | \new_[4096]_ ;
  assign \new_[4107]_  = \new_[3603]_  | \new_[3604]_ ;
  assign \new_[4110]_  = \new_[3601]_  | \new_[3602]_ ;
  assign \new_[4111]_  = \new_[4110]_  | \new_[4107]_ ;
  assign \new_[4114]_  = \new_[3599]_  | \new_[3600]_ ;
  assign \new_[4117]_  = \new_[3597]_  | \new_[3598]_ ;
  assign \new_[4118]_  = \new_[4117]_  | \new_[4114]_ ;
  assign \new_[4119]_  = \new_[4118]_  | \new_[4111]_ ;
  assign \new_[4120]_  = \new_[4119]_  | \new_[4104]_ ;
  assign \new_[4121]_  = \new_[4120]_  | \new_[4091]_ ;
  assign \new_[4122]_  = \new_[4121]_  | \new_[4062]_ ;
  assign \new_[4126]_  = \new_[3594]_  | \new_[3595]_ ;
  assign \new_[4127]_  = \new_[3596]_  | \new_[4126]_ ;
  assign \new_[4130]_  = \new_[3592]_  | \new_[3593]_ ;
  assign \new_[4133]_  = \new_[3590]_  | \new_[3591]_ ;
  assign \new_[4134]_  = \new_[4133]_  | \new_[4130]_ ;
  assign \new_[4135]_  = \new_[4134]_  | \new_[4127]_ ;
  assign \new_[4139]_  = \new_[3587]_  | \new_[3588]_ ;
  assign \new_[4140]_  = \new_[3589]_  | \new_[4139]_ ;
  assign \new_[4143]_  = \new_[3585]_  | \new_[3586]_ ;
  assign \new_[4146]_  = \new_[3583]_  | \new_[3584]_ ;
  assign \new_[4147]_  = \new_[4146]_  | \new_[4143]_ ;
  assign \new_[4148]_  = \new_[4147]_  | \new_[4140]_ ;
  assign \new_[4149]_  = \new_[4148]_  | \new_[4135]_ ;
  assign \new_[4153]_  = \new_[3580]_  | \new_[3581]_ ;
  assign \new_[4154]_  = \new_[3582]_  | \new_[4153]_ ;
  assign \new_[4157]_  = \new_[3578]_  | \new_[3579]_ ;
  assign \new_[4160]_  = \new_[3576]_  | \new_[3577]_ ;
  assign \new_[4161]_  = \new_[4160]_  | \new_[4157]_ ;
  assign \new_[4162]_  = \new_[4161]_  | \new_[4154]_ ;
  assign \new_[4165]_  = \new_[3574]_  | \new_[3575]_ ;
  assign \new_[4168]_  = \new_[3572]_  | \new_[3573]_ ;
  assign \new_[4169]_  = \new_[4168]_  | \new_[4165]_ ;
  assign \new_[4172]_  = \new_[3570]_  | \new_[3571]_ ;
  assign \new_[4175]_  = \new_[3568]_  | \new_[3569]_ ;
  assign \new_[4176]_  = \new_[4175]_  | \new_[4172]_ ;
  assign \new_[4177]_  = \new_[4176]_  | \new_[4169]_ ;
  assign \new_[4178]_  = \new_[4177]_  | \new_[4162]_ ;
  assign \new_[4179]_  = \new_[4178]_  | \new_[4149]_ ;
  assign \new_[4183]_  = \new_[3565]_  | \new_[3566]_ ;
  assign \new_[4184]_  = \new_[3567]_  | \new_[4183]_ ;
  assign \new_[4187]_  = \new_[3563]_  | \new_[3564]_ ;
  assign \new_[4190]_  = \new_[3561]_  | \new_[3562]_ ;
  assign \new_[4191]_  = \new_[4190]_  | \new_[4187]_ ;
  assign \new_[4192]_  = \new_[4191]_  | \new_[4184]_ ;
  assign \new_[4195]_  = \new_[3559]_  | \new_[3560]_ ;
  assign \new_[4198]_  = \new_[3557]_  | \new_[3558]_ ;
  assign \new_[4199]_  = \new_[4198]_  | \new_[4195]_ ;
  assign \new_[4202]_  = \new_[3555]_  | \new_[3556]_ ;
  assign \new_[4205]_  = \new_[3553]_  | \new_[3554]_ ;
  assign \new_[4206]_  = \new_[4205]_  | \new_[4202]_ ;
  assign \new_[4207]_  = \new_[4206]_  | \new_[4199]_ ;
  assign \new_[4208]_  = \new_[4207]_  | \new_[4192]_ ;
  assign \new_[4212]_  = \new_[3550]_  | \new_[3551]_ ;
  assign \new_[4213]_  = \new_[3552]_  | \new_[4212]_ ;
  assign \new_[4216]_  = \new_[3548]_  | \new_[3549]_ ;
  assign \new_[4219]_  = \new_[3546]_  | \new_[3547]_ ;
  assign \new_[4220]_  = \new_[4219]_  | \new_[4216]_ ;
  assign \new_[4221]_  = \new_[4220]_  | \new_[4213]_ ;
  assign \new_[4224]_  = \new_[3544]_  | \new_[3545]_ ;
  assign \new_[4227]_  = \new_[3542]_  | \new_[3543]_ ;
  assign \new_[4228]_  = \new_[4227]_  | \new_[4224]_ ;
  assign \new_[4231]_  = \new_[3540]_  | \new_[3541]_ ;
  assign \new_[4234]_  = \new_[3538]_  | \new_[3539]_ ;
  assign \new_[4235]_  = \new_[4234]_  | \new_[4231]_ ;
  assign \new_[4236]_  = \new_[4235]_  | \new_[4228]_ ;
  assign \new_[4237]_  = \new_[4236]_  | \new_[4221]_ ;
  assign \new_[4238]_  = \new_[4237]_  | \new_[4208]_ ;
  assign \new_[4239]_  = \new_[4238]_  | \new_[4179]_ ;
  assign \new_[4240]_  = \new_[4239]_  | \new_[4122]_ ;
  assign \new_[4241]_  = \new_[4240]_  | \new_[4005]_ ;
  assign \new_[4245]_  = \new_[3535]_  | \new_[3536]_ ;
  assign \new_[4246]_  = \new_[3537]_  | \new_[4245]_ ;
  assign \new_[4249]_  = \new_[3533]_  | \new_[3534]_ ;
  assign \new_[4252]_  = \new_[3531]_  | \new_[3532]_ ;
  assign \new_[4253]_  = \new_[4252]_  | \new_[4249]_ ;
  assign \new_[4254]_  = \new_[4253]_  | \new_[4246]_ ;
  assign \new_[4258]_  = \new_[3528]_  | \new_[3529]_ ;
  assign \new_[4259]_  = \new_[3530]_  | \new_[4258]_ ;
  assign \new_[4262]_  = \new_[3526]_  | \new_[3527]_ ;
  assign \new_[4265]_  = \new_[3524]_  | \new_[3525]_ ;
  assign \new_[4266]_  = \new_[4265]_  | \new_[4262]_ ;
  assign \new_[4267]_  = \new_[4266]_  | \new_[4259]_ ;
  assign \new_[4268]_  = \new_[4267]_  | \new_[4254]_ ;
  assign \new_[4272]_  = \new_[3521]_  | \new_[3522]_ ;
  assign \new_[4273]_  = \new_[3523]_  | \new_[4272]_ ;
  assign \new_[4276]_  = \new_[3519]_  | \new_[3520]_ ;
  assign \new_[4279]_  = \new_[3517]_  | \new_[3518]_ ;
  assign \new_[4280]_  = \new_[4279]_  | \new_[4276]_ ;
  assign \new_[4281]_  = \new_[4280]_  | \new_[4273]_ ;
  assign \new_[4284]_  = \new_[3515]_  | \new_[3516]_ ;
  assign \new_[4287]_  = \new_[3513]_  | \new_[3514]_ ;
  assign \new_[4288]_  = \new_[4287]_  | \new_[4284]_ ;
  assign \new_[4291]_  = \new_[3511]_  | \new_[3512]_ ;
  assign \new_[4294]_  = \new_[3509]_  | \new_[3510]_ ;
  assign \new_[4295]_  = \new_[4294]_  | \new_[4291]_ ;
  assign \new_[4296]_  = \new_[4295]_  | \new_[4288]_ ;
  assign \new_[4297]_  = \new_[4296]_  | \new_[4281]_ ;
  assign \new_[4298]_  = \new_[4297]_  | \new_[4268]_ ;
  assign \new_[4302]_  = \new_[3506]_  | \new_[3507]_ ;
  assign \new_[4303]_  = \new_[3508]_  | \new_[4302]_ ;
  assign \new_[4306]_  = \new_[3504]_  | \new_[3505]_ ;
  assign \new_[4309]_  = \new_[3502]_  | \new_[3503]_ ;
  assign \new_[4310]_  = \new_[4309]_  | \new_[4306]_ ;
  assign \new_[4311]_  = \new_[4310]_  | \new_[4303]_ ;
  assign \new_[4314]_  = \new_[3500]_  | \new_[3501]_ ;
  assign \new_[4317]_  = \new_[3498]_  | \new_[3499]_ ;
  assign \new_[4318]_  = \new_[4317]_  | \new_[4314]_ ;
  assign \new_[4321]_  = \new_[3496]_  | \new_[3497]_ ;
  assign \new_[4324]_  = \new_[3494]_  | \new_[3495]_ ;
  assign \new_[4325]_  = \new_[4324]_  | \new_[4321]_ ;
  assign \new_[4326]_  = \new_[4325]_  | \new_[4318]_ ;
  assign \new_[4327]_  = \new_[4326]_  | \new_[4311]_ ;
  assign \new_[4331]_  = \new_[3491]_  | \new_[3492]_ ;
  assign \new_[4332]_  = \new_[3493]_  | \new_[4331]_ ;
  assign \new_[4335]_  = \new_[3489]_  | \new_[3490]_ ;
  assign \new_[4338]_  = \new_[3487]_  | \new_[3488]_ ;
  assign \new_[4339]_  = \new_[4338]_  | \new_[4335]_ ;
  assign \new_[4340]_  = \new_[4339]_  | \new_[4332]_ ;
  assign \new_[4343]_  = \new_[3485]_  | \new_[3486]_ ;
  assign \new_[4346]_  = \new_[3483]_  | \new_[3484]_ ;
  assign \new_[4347]_  = \new_[4346]_  | \new_[4343]_ ;
  assign \new_[4350]_  = \new_[3481]_  | \new_[3482]_ ;
  assign \new_[4353]_  = \new_[3479]_  | \new_[3480]_ ;
  assign \new_[4354]_  = \new_[4353]_  | \new_[4350]_ ;
  assign \new_[4355]_  = \new_[4354]_  | \new_[4347]_ ;
  assign \new_[4356]_  = \new_[4355]_  | \new_[4340]_ ;
  assign \new_[4357]_  = \new_[4356]_  | \new_[4327]_ ;
  assign \new_[4358]_  = \new_[4357]_  | \new_[4298]_ ;
  assign \new_[4362]_  = \new_[3476]_  | \new_[3477]_ ;
  assign \new_[4363]_  = \new_[3478]_  | \new_[4362]_ ;
  assign \new_[4366]_  = \new_[3474]_  | \new_[3475]_ ;
  assign \new_[4369]_  = \new_[3472]_  | \new_[3473]_ ;
  assign \new_[4370]_  = \new_[4369]_  | \new_[4366]_ ;
  assign \new_[4371]_  = \new_[4370]_  | \new_[4363]_ ;
  assign \new_[4375]_  = \new_[3469]_  | \new_[3470]_ ;
  assign \new_[4376]_  = \new_[3471]_  | \new_[4375]_ ;
  assign \new_[4379]_  = \new_[3467]_  | \new_[3468]_ ;
  assign \new_[4382]_  = \new_[3465]_  | \new_[3466]_ ;
  assign \new_[4383]_  = \new_[4382]_  | \new_[4379]_ ;
  assign \new_[4384]_  = \new_[4383]_  | \new_[4376]_ ;
  assign \new_[4385]_  = \new_[4384]_  | \new_[4371]_ ;
  assign \new_[4389]_  = \new_[3462]_  | \new_[3463]_ ;
  assign \new_[4390]_  = \new_[3464]_  | \new_[4389]_ ;
  assign \new_[4393]_  = \new_[3460]_  | \new_[3461]_ ;
  assign \new_[4396]_  = \new_[3458]_  | \new_[3459]_ ;
  assign \new_[4397]_  = \new_[4396]_  | \new_[4393]_ ;
  assign \new_[4398]_  = \new_[4397]_  | \new_[4390]_ ;
  assign \new_[4401]_  = \new_[3456]_  | \new_[3457]_ ;
  assign \new_[4404]_  = \new_[3454]_  | \new_[3455]_ ;
  assign \new_[4405]_  = \new_[4404]_  | \new_[4401]_ ;
  assign \new_[4408]_  = \new_[3452]_  | \new_[3453]_ ;
  assign \new_[4411]_  = \new_[3450]_  | \new_[3451]_ ;
  assign \new_[4412]_  = \new_[4411]_  | \new_[4408]_ ;
  assign \new_[4413]_  = \new_[4412]_  | \new_[4405]_ ;
  assign \new_[4414]_  = \new_[4413]_  | \new_[4398]_ ;
  assign \new_[4415]_  = \new_[4414]_  | \new_[4385]_ ;
  assign \new_[4419]_  = \new_[3447]_  | \new_[3448]_ ;
  assign \new_[4420]_  = \new_[3449]_  | \new_[4419]_ ;
  assign \new_[4423]_  = \new_[3445]_  | \new_[3446]_ ;
  assign \new_[4426]_  = \new_[3443]_  | \new_[3444]_ ;
  assign \new_[4427]_  = \new_[4426]_  | \new_[4423]_ ;
  assign \new_[4428]_  = \new_[4427]_  | \new_[4420]_ ;
  assign \new_[4431]_  = \new_[3441]_  | \new_[3442]_ ;
  assign \new_[4434]_  = \new_[3439]_  | \new_[3440]_ ;
  assign \new_[4435]_  = \new_[4434]_  | \new_[4431]_ ;
  assign \new_[4438]_  = \new_[3437]_  | \new_[3438]_ ;
  assign \new_[4441]_  = \new_[3435]_  | \new_[3436]_ ;
  assign \new_[4442]_  = \new_[4441]_  | \new_[4438]_ ;
  assign \new_[4443]_  = \new_[4442]_  | \new_[4435]_ ;
  assign \new_[4444]_  = \new_[4443]_  | \new_[4428]_ ;
  assign \new_[4448]_  = \new_[3432]_  | \new_[3433]_ ;
  assign \new_[4449]_  = \new_[3434]_  | \new_[4448]_ ;
  assign \new_[4452]_  = \new_[3430]_  | \new_[3431]_ ;
  assign \new_[4455]_  = \new_[3428]_  | \new_[3429]_ ;
  assign \new_[4456]_  = \new_[4455]_  | \new_[4452]_ ;
  assign \new_[4457]_  = \new_[4456]_  | \new_[4449]_ ;
  assign \new_[4460]_  = \new_[3426]_  | \new_[3427]_ ;
  assign \new_[4463]_  = \new_[3424]_  | \new_[3425]_ ;
  assign \new_[4464]_  = \new_[4463]_  | \new_[4460]_ ;
  assign \new_[4467]_  = \new_[3422]_  | \new_[3423]_ ;
  assign \new_[4470]_  = \new_[3420]_  | \new_[3421]_ ;
  assign \new_[4471]_  = \new_[4470]_  | \new_[4467]_ ;
  assign \new_[4472]_  = \new_[4471]_  | \new_[4464]_ ;
  assign \new_[4473]_  = \new_[4472]_  | \new_[4457]_ ;
  assign \new_[4474]_  = \new_[4473]_  | \new_[4444]_ ;
  assign \new_[4475]_  = \new_[4474]_  | \new_[4415]_ ;
  assign \new_[4476]_  = \new_[4475]_  | \new_[4358]_ ;
  assign \new_[4480]_  = \new_[3417]_  | \new_[3418]_ ;
  assign \new_[4481]_  = \new_[3419]_  | \new_[4480]_ ;
  assign \new_[4484]_  = \new_[3415]_  | \new_[3416]_ ;
  assign \new_[4487]_  = \new_[3413]_  | \new_[3414]_ ;
  assign \new_[4488]_  = \new_[4487]_  | \new_[4484]_ ;
  assign \new_[4489]_  = \new_[4488]_  | \new_[4481]_ ;
  assign \new_[4493]_  = \new_[3410]_  | \new_[3411]_ ;
  assign \new_[4494]_  = \new_[3412]_  | \new_[4493]_ ;
  assign \new_[4497]_  = \new_[3408]_  | \new_[3409]_ ;
  assign \new_[4500]_  = \new_[3406]_  | \new_[3407]_ ;
  assign \new_[4501]_  = \new_[4500]_  | \new_[4497]_ ;
  assign \new_[4502]_  = \new_[4501]_  | \new_[4494]_ ;
  assign \new_[4503]_  = \new_[4502]_  | \new_[4489]_ ;
  assign \new_[4507]_  = \new_[3403]_  | \new_[3404]_ ;
  assign \new_[4508]_  = \new_[3405]_  | \new_[4507]_ ;
  assign \new_[4511]_  = \new_[3401]_  | \new_[3402]_ ;
  assign \new_[4514]_  = \new_[3399]_  | \new_[3400]_ ;
  assign \new_[4515]_  = \new_[4514]_  | \new_[4511]_ ;
  assign \new_[4516]_  = \new_[4515]_  | \new_[4508]_ ;
  assign \new_[4519]_  = \new_[3397]_  | \new_[3398]_ ;
  assign \new_[4522]_  = \new_[3395]_  | \new_[3396]_ ;
  assign \new_[4523]_  = \new_[4522]_  | \new_[4519]_ ;
  assign \new_[4526]_  = \new_[3393]_  | \new_[3394]_ ;
  assign \new_[4529]_  = \new_[3391]_  | \new_[3392]_ ;
  assign \new_[4530]_  = \new_[4529]_  | \new_[4526]_ ;
  assign \new_[4531]_  = \new_[4530]_  | \new_[4523]_ ;
  assign \new_[4532]_  = \new_[4531]_  | \new_[4516]_ ;
  assign \new_[4533]_  = \new_[4532]_  | \new_[4503]_ ;
  assign \new_[4537]_  = \new_[3388]_  | \new_[3389]_ ;
  assign \new_[4538]_  = \new_[3390]_  | \new_[4537]_ ;
  assign \new_[4541]_  = \new_[3386]_  | \new_[3387]_ ;
  assign \new_[4544]_  = \new_[3384]_  | \new_[3385]_ ;
  assign \new_[4545]_  = \new_[4544]_  | \new_[4541]_ ;
  assign \new_[4546]_  = \new_[4545]_  | \new_[4538]_ ;
  assign \new_[4549]_  = \new_[3382]_  | \new_[3383]_ ;
  assign \new_[4552]_  = \new_[3380]_  | \new_[3381]_ ;
  assign \new_[4553]_  = \new_[4552]_  | \new_[4549]_ ;
  assign \new_[4556]_  = \new_[3378]_  | \new_[3379]_ ;
  assign \new_[4559]_  = \new_[3376]_  | \new_[3377]_ ;
  assign \new_[4560]_  = \new_[4559]_  | \new_[4556]_ ;
  assign \new_[4561]_  = \new_[4560]_  | \new_[4553]_ ;
  assign \new_[4562]_  = \new_[4561]_  | \new_[4546]_ ;
  assign \new_[4566]_  = \new_[3373]_  | \new_[3374]_ ;
  assign \new_[4567]_  = \new_[3375]_  | \new_[4566]_ ;
  assign \new_[4570]_  = \new_[3371]_  | \new_[3372]_ ;
  assign \new_[4573]_  = \new_[3369]_  | \new_[3370]_ ;
  assign \new_[4574]_  = \new_[4573]_  | \new_[4570]_ ;
  assign \new_[4575]_  = \new_[4574]_  | \new_[4567]_ ;
  assign \new_[4578]_  = \new_[3367]_  | \new_[3368]_ ;
  assign \new_[4581]_  = \new_[3365]_  | \new_[3366]_ ;
  assign \new_[4582]_  = \new_[4581]_  | \new_[4578]_ ;
  assign \new_[4585]_  = \new_[3363]_  | \new_[3364]_ ;
  assign \new_[4588]_  = \new_[3361]_  | \new_[3362]_ ;
  assign \new_[4589]_  = \new_[4588]_  | \new_[4585]_ ;
  assign \new_[4590]_  = \new_[4589]_  | \new_[4582]_ ;
  assign \new_[4591]_  = \new_[4590]_  | \new_[4575]_ ;
  assign \new_[4592]_  = \new_[4591]_  | \new_[4562]_ ;
  assign \new_[4593]_  = \new_[4592]_  | \new_[4533]_ ;
  assign \new_[4597]_  = \new_[3358]_  | \new_[3359]_ ;
  assign \new_[4598]_  = \new_[3360]_  | \new_[4597]_ ;
  assign \new_[4601]_  = \new_[3356]_  | \new_[3357]_ ;
  assign \new_[4604]_  = \new_[3354]_  | \new_[3355]_ ;
  assign \new_[4605]_  = \new_[4604]_  | \new_[4601]_ ;
  assign \new_[4606]_  = \new_[4605]_  | \new_[4598]_ ;
  assign \new_[4610]_  = \new_[3351]_  | \new_[3352]_ ;
  assign \new_[4611]_  = \new_[3353]_  | \new_[4610]_ ;
  assign \new_[4614]_  = \new_[3349]_  | \new_[3350]_ ;
  assign \new_[4617]_  = \new_[3347]_  | \new_[3348]_ ;
  assign \new_[4618]_  = \new_[4617]_  | \new_[4614]_ ;
  assign \new_[4619]_  = \new_[4618]_  | \new_[4611]_ ;
  assign \new_[4620]_  = \new_[4619]_  | \new_[4606]_ ;
  assign \new_[4624]_  = \new_[3344]_  | \new_[3345]_ ;
  assign \new_[4625]_  = \new_[3346]_  | \new_[4624]_ ;
  assign \new_[4628]_  = \new_[3342]_  | \new_[3343]_ ;
  assign \new_[4631]_  = \new_[3340]_  | \new_[3341]_ ;
  assign \new_[4632]_  = \new_[4631]_  | \new_[4628]_ ;
  assign \new_[4633]_  = \new_[4632]_  | \new_[4625]_ ;
  assign \new_[4636]_  = \new_[3338]_  | \new_[3339]_ ;
  assign \new_[4639]_  = \new_[3336]_  | \new_[3337]_ ;
  assign \new_[4640]_  = \new_[4639]_  | \new_[4636]_ ;
  assign \new_[4643]_  = \new_[3334]_  | \new_[3335]_ ;
  assign \new_[4646]_  = \new_[3332]_  | \new_[3333]_ ;
  assign \new_[4647]_  = \new_[4646]_  | \new_[4643]_ ;
  assign \new_[4648]_  = \new_[4647]_  | \new_[4640]_ ;
  assign \new_[4649]_  = \new_[4648]_  | \new_[4633]_ ;
  assign \new_[4650]_  = \new_[4649]_  | \new_[4620]_ ;
  assign \new_[4654]_  = \new_[3329]_  | \new_[3330]_ ;
  assign \new_[4655]_  = \new_[3331]_  | \new_[4654]_ ;
  assign \new_[4658]_  = \new_[3327]_  | \new_[3328]_ ;
  assign \new_[4661]_  = \new_[3325]_  | \new_[3326]_ ;
  assign \new_[4662]_  = \new_[4661]_  | \new_[4658]_ ;
  assign \new_[4663]_  = \new_[4662]_  | \new_[4655]_ ;
  assign \new_[4666]_  = \new_[3323]_  | \new_[3324]_ ;
  assign \new_[4669]_  = \new_[3321]_  | \new_[3322]_ ;
  assign \new_[4670]_  = \new_[4669]_  | \new_[4666]_ ;
  assign \new_[4673]_  = \new_[3319]_  | \new_[3320]_ ;
  assign \new_[4676]_  = \new_[3317]_  | \new_[3318]_ ;
  assign \new_[4677]_  = \new_[4676]_  | \new_[4673]_ ;
  assign \new_[4678]_  = \new_[4677]_  | \new_[4670]_ ;
  assign \new_[4679]_  = \new_[4678]_  | \new_[4663]_ ;
  assign \new_[4683]_  = \new_[3314]_  | \new_[3315]_ ;
  assign \new_[4684]_  = \new_[3316]_  | \new_[4683]_ ;
  assign \new_[4687]_  = \new_[3312]_  | \new_[3313]_ ;
  assign \new_[4690]_  = \new_[3310]_  | \new_[3311]_ ;
  assign \new_[4691]_  = \new_[4690]_  | \new_[4687]_ ;
  assign \new_[4692]_  = \new_[4691]_  | \new_[4684]_ ;
  assign \new_[4695]_  = \new_[3308]_  | \new_[3309]_ ;
  assign \new_[4698]_  = \new_[3306]_  | \new_[3307]_ ;
  assign \new_[4699]_  = \new_[4698]_  | \new_[4695]_ ;
  assign \new_[4702]_  = \new_[3304]_  | \new_[3305]_ ;
  assign \new_[4705]_  = \new_[3302]_  | \new_[3303]_ ;
  assign \new_[4706]_  = \new_[4705]_  | \new_[4702]_ ;
  assign \new_[4707]_  = \new_[4706]_  | \new_[4699]_ ;
  assign \new_[4708]_  = \new_[4707]_  | \new_[4692]_ ;
  assign \new_[4709]_  = \new_[4708]_  | \new_[4679]_ ;
  assign \new_[4710]_  = \new_[4709]_  | \new_[4650]_ ;
  assign \new_[4711]_  = \new_[4710]_  | \new_[4593]_ ;
  assign \new_[4712]_  = \new_[4711]_  | \new_[4476]_ ;
  assign \new_[4713]_  = \new_[4712]_  | \new_[4241]_ ;
  assign \new_[4717]_  = \new_[3299]_  | \new_[3300]_ ;
  assign \new_[4718]_  = \new_[3301]_  | \new_[4717]_ ;
  assign \new_[4721]_  = \new_[3297]_  | \new_[3298]_ ;
  assign \new_[4724]_  = \new_[3295]_  | \new_[3296]_ ;
  assign \new_[4725]_  = \new_[4724]_  | \new_[4721]_ ;
  assign \new_[4726]_  = \new_[4725]_  | \new_[4718]_ ;
  assign \new_[4730]_  = \new_[3292]_  | \new_[3293]_ ;
  assign \new_[4731]_  = \new_[3294]_  | \new_[4730]_ ;
  assign \new_[4734]_  = \new_[3290]_  | \new_[3291]_ ;
  assign \new_[4737]_  = \new_[3288]_  | \new_[3289]_ ;
  assign \new_[4738]_  = \new_[4737]_  | \new_[4734]_ ;
  assign \new_[4739]_  = \new_[4738]_  | \new_[4731]_ ;
  assign \new_[4740]_  = \new_[4739]_  | \new_[4726]_ ;
  assign \new_[4744]_  = \new_[3285]_  | \new_[3286]_ ;
  assign \new_[4745]_  = \new_[3287]_  | \new_[4744]_ ;
  assign \new_[4748]_  = \new_[3283]_  | \new_[3284]_ ;
  assign \new_[4751]_  = \new_[3281]_  | \new_[3282]_ ;
  assign \new_[4752]_  = \new_[4751]_  | \new_[4748]_ ;
  assign \new_[4753]_  = \new_[4752]_  | \new_[4745]_ ;
  assign \new_[4756]_  = \new_[3279]_  | \new_[3280]_ ;
  assign \new_[4759]_  = \new_[3277]_  | \new_[3278]_ ;
  assign \new_[4760]_  = \new_[4759]_  | \new_[4756]_ ;
  assign \new_[4763]_  = \new_[3275]_  | \new_[3276]_ ;
  assign \new_[4766]_  = \new_[3273]_  | \new_[3274]_ ;
  assign \new_[4767]_  = \new_[4766]_  | \new_[4763]_ ;
  assign \new_[4768]_  = \new_[4767]_  | \new_[4760]_ ;
  assign \new_[4769]_  = \new_[4768]_  | \new_[4753]_ ;
  assign \new_[4770]_  = \new_[4769]_  | \new_[4740]_ ;
  assign \new_[4774]_  = \new_[3270]_  | \new_[3271]_ ;
  assign \new_[4775]_  = \new_[3272]_  | \new_[4774]_ ;
  assign \new_[4778]_  = \new_[3268]_  | \new_[3269]_ ;
  assign \new_[4781]_  = \new_[3266]_  | \new_[3267]_ ;
  assign \new_[4782]_  = \new_[4781]_  | \new_[4778]_ ;
  assign \new_[4783]_  = \new_[4782]_  | \new_[4775]_ ;
  assign \new_[4786]_  = \new_[3264]_  | \new_[3265]_ ;
  assign \new_[4789]_  = \new_[3262]_  | \new_[3263]_ ;
  assign \new_[4790]_  = \new_[4789]_  | \new_[4786]_ ;
  assign \new_[4793]_  = \new_[3260]_  | \new_[3261]_ ;
  assign \new_[4796]_  = \new_[3258]_  | \new_[3259]_ ;
  assign \new_[4797]_  = \new_[4796]_  | \new_[4793]_ ;
  assign \new_[4798]_  = \new_[4797]_  | \new_[4790]_ ;
  assign \new_[4799]_  = \new_[4798]_  | \new_[4783]_ ;
  assign \new_[4803]_  = \new_[3255]_  | \new_[3256]_ ;
  assign \new_[4804]_  = \new_[3257]_  | \new_[4803]_ ;
  assign \new_[4807]_  = \new_[3253]_  | \new_[3254]_ ;
  assign \new_[4810]_  = \new_[3251]_  | \new_[3252]_ ;
  assign \new_[4811]_  = \new_[4810]_  | \new_[4807]_ ;
  assign \new_[4812]_  = \new_[4811]_  | \new_[4804]_ ;
  assign \new_[4815]_  = \new_[3249]_  | \new_[3250]_ ;
  assign \new_[4818]_  = \new_[3247]_  | \new_[3248]_ ;
  assign \new_[4819]_  = \new_[4818]_  | \new_[4815]_ ;
  assign \new_[4822]_  = \new_[3245]_  | \new_[3246]_ ;
  assign \new_[4825]_  = \new_[3243]_  | \new_[3244]_ ;
  assign \new_[4826]_  = \new_[4825]_  | \new_[4822]_ ;
  assign \new_[4827]_  = \new_[4826]_  | \new_[4819]_ ;
  assign \new_[4828]_  = \new_[4827]_  | \new_[4812]_ ;
  assign \new_[4829]_  = \new_[4828]_  | \new_[4799]_ ;
  assign \new_[4830]_  = \new_[4829]_  | \new_[4770]_ ;
  assign \new_[4834]_  = \new_[3240]_  | \new_[3241]_ ;
  assign \new_[4835]_  = \new_[3242]_  | \new_[4834]_ ;
  assign \new_[4838]_  = \new_[3238]_  | \new_[3239]_ ;
  assign \new_[4841]_  = \new_[3236]_  | \new_[3237]_ ;
  assign \new_[4842]_  = \new_[4841]_  | \new_[4838]_ ;
  assign \new_[4843]_  = \new_[4842]_  | \new_[4835]_ ;
  assign \new_[4847]_  = \new_[3233]_  | \new_[3234]_ ;
  assign \new_[4848]_  = \new_[3235]_  | \new_[4847]_ ;
  assign \new_[4851]_  = \new_[3231]_  | \new_[3232]_ ;
  assign \new_[4854]_  = \new_[3229]_  | \new_[3230]_ ;
  assign \new_[4855]_  = \new_[4854]_  | \new_[4851]_ ;
  assign \new_[4856]_  = \new_[4855]_  | \new_[4848]_ ;
  assign \new_[4857]_  = \new_[4856]_  | \new_[4843]_ ;
  assign \new_[4861]_  = \new_[3226]_  | \new_[3227]_ ;
  assign \new_[4862]_  = \new_[3228]_  | \new_[4861]_ ;
  assign \new_[4865]_  = \new_[3224]_  | \new_[3225]_ ;
  assign \new_[4868]_  = \new_[3222]_  | \new_[3223]_ ;
  assign \new_[4869]_  = \new_[4868]_  | \new_[4865]_ ;
  assign \new_[4870]_  = \new_[4869]_  | \new_[4862]_ ;
  assign \new_[4873]_  = \new_[3220]_  | \new_[3221]_ ;
  assign \new_[4876]_  = \new_[3218]_  | \new_[3219]_ ;
  assign \new_[4877]_  = \new_[4876]_  | \new_[4873]_ ;
  assign \new_[4880]_  = \new_[3216]_  | \new_[3217]_ ;
  assign \new_[4883]_  = \new_[3214]_  | \new_[3215]_ ;
  assign \new_[4884]_  = \new_[4883]_  | \new_[4880]_ ;
  assign \new_[4885]_  = \new_[4884]_  | \new_[4877]_ ;
  assign \new_[4886]_  = \new_[4885]_  | \new_[4870]_ ;
  assign \new_[4887]_  = \new_[4886]_  | \new_[4857]_ ;
  assign \new_[4891]_  = \new_[3211]_  | \new_[3212]_ ;
  assign \new_[4892]_  = \new_[3213]_  | \new_[4891]_ ;
  assign \new_[4895]_  = \new_[3209]_  | \new_[3210]_ ;
  assign \new_[4898]_  = \new_[3207]_  | \new_[3208]_ ;
  assign \new_[4899]_  = \new_[4898]_  | \new_[4895]_ ;
  assign \new_[4900]_  = \new_[4899]_  | \new_[4892]_ ;
  assign \new_[4903]_  = \new_[3205]_  | \new_[3206]_ ;
  assign \new_[4906]_  = \new_[3203]_  | \new_[3204]_ ;
  assign \new_[4907]_  = \new_[4906]_  | \new_[4903]_ ;
  assign \new_[4910]_  = \new_[3201]_  | \new_[3202]_ ;
  assign \new_[4913]_  = \new_[3199]_  | \new_[3200]_ ;
  assign \new_[4914]_  = \new_[4913]_  | \new_[4910]_ ;
  assign \new_[4915]_  = \new_[4914]_  | \new_[4907]_ ;
  assign \new_[4916]_  = \new_[4915]_  | \new_[4900]_ ;
  assign \new_[4920]_  = \new_[3196]_  | \new_[3197]_ ;
  assign \new_[4921]_  = \new_[3198]_  | \new_[4920]_ ;
  assign \new_[4924]_  = \new_[3194]_  | \new_[3195]_ ;
  assign \new_[4927]_  = \new_[3192]_  | \new_[3193]_ ;
  assign \new_[4928]_  = \new_[4927]_  | \new_[4924]_ ;
  assign \new_[4929]_  = \new_[4928]_  | \new_[4921]_ ;
  assign \new_[4932]_  = \new_[3190]_  | \new_[3191]_ ;
  assign \new_[4935]_  = \new_[3188]_  | \new_[3189]_ ;
  assign \new_[4936]_  = \new_[4935]_  | \new_[4932]_ ;
  assign \new_[4939]_  = \new_[3186]_  | \new_[3187]_ ;
  assign \new_[4942]_  = \new_[3184]_  | \new_[3185]_ ;
  assign \new_[4943]_  = \new_[4942]_  | \new_[4939]_ ;
  assign \new_[4944]_  = \new_[4943]_  | \new_[4936]_ ;
  assign \new_[4945]_  = \new_[4944]_  | \new_[4929]_ ;
  assign \new_[4946]_  = \new_[4945]_  | \new_[4916]_ ;
  assign \new_[4947]_  = \new_[4946]_  | \new_[4887]_ ;
  assign \new_[4948]_  = \new_[4947]_  | \new_[4830]_ ;
  assign \new_[4952]_  = \new_[3181]_  | \new_[3182]_ ;
  assign \new_[4953]_  = \new_[3183]_  | \new_[4952]_ ;
  assign \new_[4956]_  = \new_[3179]_  | \new_[3180]_ ;
  assign \new_[4959]_  = \new_[3177]_  | \new_[3178]_ ;
  assign \new_[4960]_  = \new_[4959]_  | \new_[4956]_ ;
  assign \new_[4961]_  = \new_[4960]_  | \new_[4953]_ ;
  assign \new_[4965]_  = \new_[3174]_  | \new_[3175]_ ;
  assign \new_[4966]_  = \new_[3176]_  | \new_[4965]_ ;
  assign \new_[4969]_  = \new_[3172]_  | \new_[3173]_ ;
  assign \new_[4972]_  = \new_[3170]_  | \new_[3171]_ ;
  assign \new_[4973]_  = \new_[4972]_  | \new_[4969]_ ;
  assign \new_[4974]_  = \new_[4973]_  | \new_[4966]_ ;
  assign \new_[4975]_  = \new_[4974]_  | \new_[4961]_ ;
  assign \new_[4979]_  = \new_[3167]_  | \new_[3168]_ ;
  assign \new_[4980]_  = \new_[3169]_  | \new_[4979]_ ;
  assign \new_[4983]_  = \new_[3165]_  | \new_[3166]_ ;
  assign \new_[4986]_  = \new_[3163]_  | \new_[3164]_ ;
  assign \new_[4987]_  = \new_[4986]_  | \new_[4983]_ ;
  assign \new_[4988]_  = \new_[4987]_  | \new_[4980]_ ;
  assign \new_[4991]_  = \new_[3161]_  | \new_[3162]_ ;
  assign \new_[4994]_  = \new_[3159]_  | \new_[3160]_ ;
  assign \new_[4995]_  = \new_[4994]_  | \new_[4991]_ ;
  assign \new_[4998]_  = \new_[3157]_  | \new_[3158]_ ;
  assign \new_[5001]_  = \new_[3155]_  | \new_[3156]_ ;
  assign \new_[5002]_  = \new_[5001]_  | \new_[4998]_ ;
  assign \new_[5003]_  = \new_[5002]_  | \new_[4995]_ ;
  assign \new_[5004]_  = \new_[5003]_  | \new_[4988]_ ;
  assign \new_[5005]_  = \new_[5004]_  | \new_[4975]_ ;
  assign \new_[5009]_  = \new_[3152]_  | \new_[3153]_ ;
  assign \new_[5010]_  = \new_[3154]_  | \new_[5009]_ ;
  assign \new_[5013]_  = \new_[3150]_  | \new_[3151]_ ;
  assign \new_[5016]_  = \new_[3148]_  | \new_[3149]_ ;
  assign \new_[5017]_  = \new_[5016]_  | \new_[5013]_ ;
  assign \new_[5018]_  = \new_[5017]_  | \new_[5010]_ ;
  assign \new_[5021]_  = \new_[3146]_  | \new_[3147]_ ;
  assign \new_[5024]_  = \new_[3144]_  | \new_[3145]_ ;
  assign \new_[5025]_  = \new_[5024]_  | \new_[5021]_ ;
  assign \new_[5028]_  = \new_[3142]_  | \new_[3143]_ ;
  assign \new_[5031]_  = \new_[3140]_  | \new_[3141]_ ;
  assign \new_[5032]_  = \new_[5031]_  | \new_[5028]_ ;
  assign \new_[5033]_  = \new_[5032]_  | \new_[5025]_ ;
  assign \new_[5034]_  = \new_[5033]_  | \new_[5018]_ ;
  assign \new_[5038]_  = \new_[3137]_  | \new_[3138]_ ;
  assign \new_[5039]_  = \new_[3139]_  | \new_[5038]_ ;
  assign \new_[5042]_  = \new_[3135]_  | \new_[3136]_ ;
  assign \new_[5045]_  = \new_[3133]_  | \new_[3134]_ ;
  assign \new_[5046]_  = \new_[5045]_  | \new_[5042]_ ;
  assign \new_[5047]_  = \new_[5046]_  | \new_[5039]_ ;
  assign \new_[5050]_  = \new_[3131]_  | \new_[3132]_ ;
  assign \new_[5053]_  = \new_[3129]_  | \new_[3130]_ ;
  assign \new_[5054]_  = \new_[5053]_  | \new_[5050]_ ;
  assign \new_[5057]_  = \new_[3127]_  | \new_[3128]_ ;
  assign \new_[5060]_  = \new_[3125]_  | \new_[3126]_ ;
  assign \new_[5061]_  = \new_[5060]_  | \new_[5057]_ ;
  assign \new_[5062]_  = \new_[5061]_  | \new_[5054]_ ;
  assign \new_[5063]_  = \new_[5062]_  | \new_[5047]_ ;
  assign \new_[5064]_  = \new_[5063]_  | \new_[5034]_ ;
  assign \new_[5065]_  = \new_[5064]_  | \new_[5005]_ ;
  assign \new_[5069]_  = \new_[3122]_  | \new_[3123]_ ;
  assign \new_[5070]_  = \new_[3124]_  | \new_[5069]_ ;
  assign \new_[5073]_  = \new_[3120]_  | \new_[3121]_ ;
  assign \new_[5076]_  = \new_[3118]_  | \new_[3119]_ ;
  assign \new_[5077]_  = \new_[5076]_  | \new_[5073]_ ;
  assign \new_[5078]_  = \new_[5077]_  | \new_[5070]_ ;
  assign \new_[5082]_  = \new_[3115]_  | \new_[3116]_ ;
  assign \new_[5083]_  = \new_[3117]_  | \new_[5082]_ ;
  assign \new_[5086]_  = \new_[3113]_  | \new_[3114]_ ;
  assign \new_[5089]_  = \new_[3111]_  | \new_[3112]_ ;
  assign \new_[5090]_  = \new_[5089]_  | \new_[5086]_ ;
  assign \new_[5091]_  = \new_[5090]_  | \new_[5083]_ ;
  assign \new_[5092]_  = \new_[5091]_  | \new_[5078]_ ;
  assign \new_[5096]_  = \new_[3108]_  | \new_[3109]_ ;
  assign \new_[5097]_  = \new_[3110]_  | \new_[5096]_ ;
  assign \new_[5100]_  = \new_[3106]_  | \new_[3107]_ ;
  assign \new_[5103]_  = \new_[3104]_  | \new_[3105]_ ;
  assign \new_[5104]_  = \new_[5103]_  | \new_[5100]_ ;
  assign \new_[5105]_  = \new_[5104]_  | \new_[5097]_ ;
  assign \new_[5108]_  = \new_[3102]_  | \new_[3103]_ ;
  assign \new_[5111]_  = \new_[3100]_  | \new_[3101]_ ;
  assign \new_[5112]_  = \new_[5111]_  | \new_[5108]_ ;
  assign \new_[5115]_  = \new_[3098]_  | \new_[3099]_ ;
  assign \new_[5118]_  = \new_[3096]_  | \new_[3097]_ ;
  assign \new_[5119]_  = \new_[5118]_  | \new_[5115]_ ;
  assign \new_[5120]_  = \new_[5119]_  | \new_[5112]_ ;
  assign \new_[5121]_  = \new_[5120]_  | \new_[5105]_ ;
  assign \new_[5122]_  = \new_[5121]_  | \new_[5092]_ ;
  assign \new_[5126]_  = \new_[3093]_  | \new_[3094]_ ;
  assign \new_[5127]_  = \new_[3095]_  | \new_[5126]_ ;
  assign \new_[5130]_  = \new_[3091]_  | \new_[3092]_ ;
  assign \new_[5133]_  = \new_[3089]_  | \new_[3090]_ ;
  assign \new_[5134]_  = \new_[5133]_  | \new_[5130]_ ;
  assign \new_[5135]_  = \new_[5134]_  | \new_[5127]_ ;
  assign \new_[5138]_  = \new_[3087]_  | \new_[3088]_ ;
  assign \new_[5141]_  = \new_[3085]_  | \new_[3086]_ ;
  assign \new_[5142]_  = \new_[5141]_  | \new_[5138]_ ;
  assign \new_[5145]_  = \new_[3083]_  | \new_[3084]_ ;
  assign \new_[5148]_  = \new_[3081]_  | \new_[3082]_ ;
  assign \new_[5149]_  = \new_[5148]_  | \new_[5145]_ ;
  assign \new_[5150]_  = \new_[5149]_  | \new_[5142]_ ;
  assign \new_[5151]_  = \new_[5150]_  | \new_[5135]_ ;
  assign \new_[5155]_  = \new_[3078]_  | \new_[3079]_ ;
  assign \new_[5156]_  = \new_[3080]_  | \new_[5155]_ ;
  assign \new_[5159]_  = \new_[3076]_  | \new_[3077]_ ;
  assign \new_[5162]_  = \new_[3074]_  | \new_[3075]_ ;
  assign \new_[5163]_  = \new_[5162]_  | \new_[5159]_ ;
  assign \new_[5164]_  = \new_[5163]_  | \new_[5156]_ ;
  assign \new_[5167]_  = \new_[3072]_  | \new_[3073]_ ;
  assign \new_[5170]_  = \new_[3070]_  | \new_[3071]_ ;
  assign \new_[5171]_  = \new_[5170]_  | \new_[5167]_ ;
  assign \new_[5174]_  = \new_[3068]_  | \new_[3069]_ ;
  assign \new_[5177]_  = \new_[3066]_  | \new_[3067]_ ;
  assign \new_[5178]_  = \new_[5177]_  | \new_[5174]_ ;
  assign \new_[5179]_  = \new_[5178]_  | \new_[5171]_ ;
  assign \new_[5180]_  = \new_[5179]_  | \new_[5164]_ ;
  assign \new_[5181]_  = \new_[5180]_  | \new_[5151]_ ;
  assign \new_[5182]_  = \new_[5181]_  | \new_[5122]_ ;
  assign \new_[5183]_  = \new_[5182]_  | \new_[5065]_ ;
  assign \new_[5184]_  = \new_[5183]_  | \new_[4948]_ ;
  assign \new_[5188]_  = \new_[3063]_  | \new_[3064]_ ;
  assign \new_[5189]_  = \new_[3065]_  | \new_[5188]_ ;
  assign \new_[5192]_  = \new_[3061]_  | \new_[3062]_ ;
  assign \new_[5195]_  = \new_[3059]_  | \new_[3060]_ ;
  assign \new_[5196]_  = \new_[5195]_  | \new_[5192]_ ;
  assign \new_[5197]_  = \new_[5196]_  | \new_[5189]_ ;
  assign \new_[5201]_  = \new_[3056]_  | \new_[3057]_ ;
  assign \new_[5202]_  = \new_[3058]_  | \new_[5201]_ ;
  assign \new_[5205]_  = \new_[3054]_  | \new_[3055]_ ;
  assign \new_[5208]_  = \new_[3052]_  | \new_[3053]_ ;
  assign \new_[5209]_  = \new_[5208]_  | \new_[5205]_ ;
  assign \new_[5210]_  = \new_[5209]_  | \new_[5202]_ ;
  assign \new_[5211]_  = \new_[5210]_  | \new_[5197]_ ;
  assign \new_[5215]_  = \new_[3049]_  | \new_[3050]_ ;
  assign \new_[5216]_  = \new_[3051]_  | \new_[5215]_ ;
  assign \new_[5219]_  = \new_[3047]_  | \new_[3048]_ ;
  assign \new_[5222]_  = \new_[3045]_  | \new_[3046]_ ;
  assign \new_[5223]_  = \new_[5222]_  | \new_[5219]_ ;
  assign \new_[5224]_  = \new_[5223]_  | \new_[5216]_ ;
  assign \new_[5227]_  = \new_[3043]_  | \new_[3044]_ ;
  assign \new_[5230]_  = \new_[3041]_  | \new_[3042]_ ;
  assign \new_[5231]_  = \new_[5230]_  | \new_[5227]_ ;
  assign \new_[5234]_  = \new_[3039]_  | \new_[3040]_ ;
  assign \new_[5237]_  = \new_[3037]_  | \new_[3038]_ ;
  assign \new_[5238]_  = \new_[5237]_  | \new_[5234]_ ;
  assign \new_[5239]_  = \new_[5238]_  | \new_[5231]_ ;
  assign \new_[5240]_  = \new_[5239]_  | \new_[5224]_ ;
  assign \new_[5241]_  = \new_[5240]_  | \new_[5211]_ ;
  assign \new_[5245]_  = \new_[3034]_  | \new_[3035]_ ;
  assign \new_[5246]_  = \new_[3036]_  | \new_[5245]_ ;
  assign \new_[5249]_  = \new_[3032]_  | \new_[3033]_ ;
  assign \new_[5252]_  = \new_[3030]_  | \new_[3031]_ ;
  assign \new_[5253]_  = \new_[5252]_  | \new_[5249]_ ;
  assign \new_[5254]_  = \new_[5253]_  | \new_[5246]_ ;
  assign \new_[5257]_  = \new_[3028]_  | \new_[3029]_ ;
  assign \new_[5260]_  = \new_[3026]_  | \new_[3027]_ ;
  assign \new_[5261]_  = \new_[5260]_  | \new_[5257]_ ;
  assign \new_[5264]_  = \new_[3024]_  | \new_[3025]_ ;
  assign \new_[5267]_  = \new_[3022]_  | \new_[3023]_ ;
  assign \new_[5268]_  = \new_[5267]_  | \new_[5264]_ ;
  assign \new_[5269]_  = \new_[5268]_  | \new_[5261]_ ;
  assign \new_[5270]_  = \new_[5269]_  | \new_[5254]_ ;
  assign \new_[5274]_  = \new_[3019]_  | \new_[3020]_ ;
  assign \new_[5275]_  = \new_[3021]_  | \new_[5274]_ ;
  assign \new_[5278]_  = \new_[3017]_  | \new_[3018]_ ;
  assign \new_[5281]_  = \new_[3015]_  | \new_[3016]_ ;
  assign \new_[5282]_  = \new_[5281]_  | \new_[5278]_ ;
  assign \new_[5283]_  = \new_[5282]_  | \new_[5275]_ ;
  assign \new_[5286]_  = \new_[3013]_  | \new_[3014]_ ;
  assign \new_[5289]_  = \new_[3011]_  | \new_[3012]_ ;
  assign \new_[5290]_  = \new_[5289]_  | \new_[5286]_ ;
  assign \new_[5293]_  = \new_[3009]_  | \new_[3010]_ ;
  assign \new_[5296]_  = \new_[3007]_  | \new_[3008]_ ;
  assign \new_[5297]_  = \new_[5296]_  | \new_[5293]_ ;
  assign \new_[5298]_  = \new_[5297]_  | \new_[5290]_ ;
  assign \new_[5299]_  = \new_[5298]_  | \new_[5283]_ ;
  assign \new_[5300]_  = \new_[5299]_  | \new_[5270]_ ;
  assign \new_[5301]_  = \new_[5300]_  | \new_[5241]_ ;
  assign \new_[5305]_  = \new_[3004]_  | \new_[3005]_ ;
  assign \new_[5306]_  = \new_[3006]_  | \new_[5305]_ ;
  assign \new_[5309]_  = \new_[3002]_  | \new_[3003]_ ;
  assign \new_[5312]_  = \new_[3000]_  | \new_[3001]_ ;
  assign \new_[5313]_  = \new_[5312]_  | \new_[5309]_ ;
  assign \new_[5314]_  = \new_[5313]_  | \new_[5306]_ ;
  assign \new_[5318]_  = \new_[2997]_  | \new_[2998]_ ;
  assign \new_[5319]_  = \new_[2999]_  | \new_[5318]_ ;
  assign \new_[5322]_  = \new_[2995]_  | \new_[2996]_ ;
  assign \new_[5325]_  = \new_[2993]_  | \new_[2994]_ ;
  assign \new_[5326]_  = \new_[5325]_  | \new_[5322]_ ;
  assign \new_[5327]_  = \new_[5326]_  | \new_[5319]_ ;
  assign \new_[5328]_  = \new_[5327]_  | \new_[5314]_ ;
  assign \new_[5332]_  = \new_[2990]_  | \new_[2991]_ ;
  assign \new_[5333]_  = \new_[2992]_  | \new_[5332]_ ;
  assign \new_[5336]_  = \new_[2988]_  | \new_[2989]_ ;
  assign \new_[5339]_  = \new_[2986]_  | \new_[2987]_ ;
  assign \new_[5340]_  = \new_[5339]_  | \new_[5336]_ ;
  assign \new_[5341]_  = \new_[5340]_  | \new_[5333]_ ;
  assign \new_[5344]_  = \new_[2984]_  | \new_[2985]_ ;
  assign \new_[5347]_  = \new_[2982]_  | \new_[2983]_ ;
  assign \new_[5348]_  = \new_[5347]_  | \new_[5344]_ ;
  assign \new_[5351]_  = \new_[2980]_  | \new_[2981]_ ;
  assign \new_[5354]_  = \new_[2978]_  | \new_[2979]_ ;
  assign \new_[5355]_  = \new_[5354]_  | \new_[5351]_ ;
  assign \new_[5356]_  = \new_[5355]_  | \new_[5348]_ ;
  assign \new_[5357]_  = \new_[5356]_  | \new_[5341]_ ;
  assign \new_[5358]_  = \new_[5357]_  | \new_[5328]_ ;
  assign \new_[5362]_  = \new_[2975]_  | \new_[2976]_ ;
  assign \new_[5363]_  = \new_[2977]_  | \new_[5362]_ ;
  assign \new_[5366]_  = \new_[2973]_  | \new_[2974]_ ;
  assign \new_[5369]_  = \new_[2971]_  | \new_[2972]_ ;
  assign \new_[5370]_  = \new_[5369]_  | \new_[5366]_ ;
  assign \new_[5371]_  = \new_[5370]_  | \new_[5363]_ ;
  assign \new_[5374]_  = \new_[2969]_  | \new_[2970]_ ;
  assign \new_[5377]_  = \new_[2967]_  | \new_[2968]_ ;
  assign \new_[5378]_  = \new_[5377]_  | \new_[5374]_ ;
  assign \new_[5381]_  = \new_[2965]_  | \new_[2966]_ ;
  assign \new_[5384]_  = \new_[2963]_  | \new_[2964]_ ;
  assign \new_[5385]_  = \new_[5384]_  | \new_[5381]_ ;
  assign \new_[5386]_  = \new_[5385]_  | \new_[5378]_ ;
  assign \new_[5387]_  = \new_[5386]_  | \new_[5371]_ ;
  assign \new_[5391]_  = \new_[2960]_  | \new_[2961]_ ;
  assign \new_[5392]_  = \new_[2962]_  | \new_[5391]_ ;
  assign \new_[5395]_  = \new_[2958]_  | \new_[2959]_ ;
  assign \new_[5398]_  = \new_[2956]_  | \new_[2957]_ ;
  assign \new_[5399]_  = \new_[5398]_  | \new_[5395]_ ;
  assign \new_[5400]_  = \new_[5399]_  | \new_[5392]_ ;
  assign \new_[5403]_  = \new_[2954]_  | \new_[2955]_ ;
  assign \new_[5406]_  = \new_[2952]_  | \new_[2953]_ ;
  assign \new_[5407]_  = \new_[5406]_  | \new_[5403]_ ;
  assign \new_[5410]_  = \new_[2950]_  | \new_[2951]_ ;
  assign \new_[5413]_  = \new_[2948]_  | \new_[2949]_ ;
  assign \new_[5414]_  = \new_[5413]_  | \new_[5410]_ ;
  assign \new_[5415]_  = \new_[5414]_  | \new_[5407]_ ;
  assign \new_[5416]_  = \new_[5415]_  | \new_[5400]_ ;
  assign \new_[5417]_  = \new_[5416]_  | \new_[5387]_ ;
  assign \new_[5418]_  = \new_[5417]_  | \new_[5358]_ ;
  assign \new_[5419]_  = \new_[5418]_  | \new_[5301]_ ;
  assign \new_[5423]_  = \new_[2945]_  | \new_[2946]_ ;
  assign \new_[5424]_  = \new_[2947]_  | \new_[5423]_ ;
  assign \new_[5427]_  = \new_[2943]_  | \new_[2944]_ ;
  assign \new_[5430]_  = \new_[2941]_  | \new_[2942]_ ;
  assign \new_[5431]_  = \new_[5430]_  | \new_[5427]_ ;
  assign \new_[5432]_  = \new_[5431]_  | \new_[5424]_ ;
  assign \new_[5436]_  = \new_[2938]_  | \new_[2939]_ ;
  assign \new_[5437]_  = \new_[2940]_  | \new_[5436]_ ;
  assign \new_[5440]_  = \new_[2936]_  | \new_[2937]_ ;
  assign \new_[5443]_  = \new_[2934]_  | \new_[2935]_ ;
  assign \new_[5444]_  = \new_[5443]_  | \new_[5440]_ ;
  assign \new_[5445]_  = \new_[5444]_  | \new_[5437]_ ;
  assign \new_[5446]_  = \new_[5445]_  | \new_[5432]_ ;
  assign \new_[5450]_  = \new_[2931]_  | \new_[2932]_ ;
  assign \new_[5451]_  = \new_[2933]_  | \new_[5450]_ ;
  assign \new_[5454]_  = \new_[2929]_  | \new_[2930]_ ;
  assign \new_[5457]_  = \new_[2927]_  | \new_[2928]_ ;
  assign \new_[5458]_  = \new_[5457]_  | \new_[5454]_ ;
  assign \new_[5459]_  = \new_[5458]_  | \new_[5451]_ ;
  assign \new_[5462]_  = \new_[2925]_  | \new_[2926]_ ;
  assign \new_[5465]_  = \new_[2923]_  | \new_[2924]_ ;
  assign \new_[5466]_  = \new_[5465]_  | \new_[5462]_ ;
  assign \new_[5469]_  = \new_[2921]_  | \new_[2922]_ ;
  assign \new_[5472]_  = \new_[2919]_  | \new_[2920]_ ;
  assign \new_[5473]_  = \new_[5472]_  | \new_[5469]_ ;
  assign \new_[5474]_  = \new_[5473]_  | \new_[5466]_ ;
  assign \new_[5475]_  = \new_[5474]_  | \new_[5459]_ ;
  assign \new_[5476]_  = \new_[5475]_  | \new_[5446]_ ;
  assign \new_[5480]_  = \new_[2916]_  | \new_[2917]_ ;
  assign \new_[5481]_  = \new_[2918]_  | \new_[5480]_ ;
  assign \new_[5484]_  = \new_[2914]_  | \new_[2915]_ ;
  assign \new_[5487]_  = \new_[2912]_  | \new_[2913]_ ;
  assign \new_[5488]_  = \new_[5487]_  | \new_[5484]_ ;
  assign \new_[5489]_  = \new_[5488]_  | \new_[5481]_ ;
  assign \new_[5492]_  = \new_[2910]_  | \new_[2911]_ ;
  assign \new_[5495]_  = \new_[2908]_  | \new_[2909]_ ;
  assign \new_[5496]_  = \new_[5495]_  | \new_[5492]_ ;
  assign \new_[5499]_  = \new_[2906]_  | \new_[2907]_ ;
  assign \new_[5502]_  = \new_[2904]_  | \new_[2905]_ ;
  assign \new_[5503]_  = \new_[5502]_  | \new_[5499]_ ;
  assign \new_[5504]_  = \new_[5503]_  | \new_[5496]_ ;
  assign \new_[5505]_  = \new_[5504]_  | \new_[5489]_ ;
  assign \new_[5509]_  = \new_[2901]_  | \new_[2902]_ ;
  assign \new_[5510]_  = \new_[2903]_  | \new_[5509]_ ;
  assign \new_[5513]_  = \new_[2899]_  | \new_[2900]_ ;
  assign \new_[5516]_  = \new_[2897]_  | \new_[2898]_ ;
  assign \new_[5517]_  = \new_[5516]_  | \new_[5513]_ ;
  assign \new_[5518]_  = \new_[5517]_  | \new_[5510]_ ;
  assign \new_[5521]_  = \new_[2895]_  | \new_[2896]_ ;
  assign \new_[5524]_  = \new_[2893]_  | \new_[2894]_ ;
  assign \new_[5525]_  = \new_[5524]_  | \new_[5521]_ ;
  assign \new_[5528]_  = \new_[2891]_  | \new_[2892]_ ;
  assign \new_[5531]_  = \new_[2889]_  | \new_[2890]_ ;
  assign \new_[5532]_  = \new_[5531]_  | \new_[5528]_ ;
  assign \new_[5533]_  = \new_[5532]_  | \new_[5525]_ ;
  assign \new_[5534]_  = \new_[5533]_  | \new_[5518]_ ;
  assign \new_[5535]_  = \new_[5534]_  | \new_[5505]_ ;
  assign \new_[5536]_  = \new_[5535]_  | \new_[5476]_ ;
  assign \new_[5540]_  = \new_[2886]_  | \new_[2887]_ ;
  assign \new_[5541]_  = \new_[2888]_  | \new_[5540]_ ;
  assign \new_[5544]_  = \new_[2884]_  | \new_[2885]_ ;
  assign \new_[5547]_  = \new_[2882]_  | \new_[2883]_ ;
  assign \new_[5548]_  = \new_[5547]_  | \new_[5544]_ ;
  assign \new_[5549]_  = \new_[5548]_  | \new_[5541]_ ;
  assign \new_[5553]_  = \new_[2879]_  | \new_[2880]_ ;
  assign \new_[5554]_  = \new_[2881]_  | \new_[5553]_ ;
  assign \new_[5557]_  = \new_[2877]_  | \new_[2878]_ ;
  assign \new_[5560]_  = \new_[2875]_  | \new_[2876]_ ;
  assign \new_[5561]_  = \new_[5560]_  | \new_[5557]_ ;
  assign \new_[5562]_  = \new_[5561]_  | \new_[5554]_ ;
  assign \new_[5563]_  = \new_[5562]_  | \new_[5549]_ ;
  assign \new_[5567]_  = \new_[2872]_  | \new_[2873]_ ;
  assign \new_[5568]_  = \new_[2874]_  | \new_[5567]_ ;
  assign \new_[5571]_  = \new_[2870]_  | \new_[2871]_ ;
  assign \new_[5574]_  = \new_[2868]_  | \new_[2869]_ ;
  assign \new_[5575]_  = \new_[5574]_  | \new_[5571]_ ;
  assign \new_[5576]_  = \new_[5575]_  | \new_[5568]_ ;
  assign \new_[5579]_  = \new_[2866]_  | \new_[2867]_ ;
  assign \new_[5582]_  = \new_[2864]_  | \new_[2865]_ ;
  assign \new_[5583]_  = \new_[5582]_  | \new_[5579]_ ;
  assign \new_[5586]_  = \new_[2862]_  | \new_[2863]_ ;
  assign \new_[5589]_  = \new_[2860]_  | \new_[2861]_ ;
  assign \new_[5590]_  = \new_[5589]_  | \new_[5586]_ ;
  assign \new_[5591]_  = \new_[5590]_  | \new_[5583]_ ;
  assign \new_[5592]_  = \new_[5591]_  | \new_[5576]_ ;
  assign \new_[5593]_  = \new_[5592]_  | \new_[5563]_ ;
  assign \new_[5597]_  = \new_[2857]_  | \new_[2858]_ ;
  assign \new_[5598]_  = \new_[2859]_  | \new_[5597]_ ;
  assign \new_[5601]_  = \new_[2855]_  | \new_[2856]_ ;
  assign \new_[5604]_  = \new_[2853]_  | \new_[2854]_ ;
  assign \new_[5605]_  = \new_[5604]_  | \new_[5601]_ ;
  assign \new_[5606]_  = \new_[5605]_  | \new_[5598]_ ;
  assign \new_[5609]_  = \new_[2851]_  | \new_[2852]_ ;
  assign \new_[5612]_  = \new_[2849]_  | \new_[2850]_ ;
  assign \new_[5613]_  = \new_[5612]_  | \new_[5609]_ ;
  assign \new_[5616]_  = \new_[2847]_  | \new_[2848]_ ;
  assign \new_[5619]_  = \new_[2845]_  | \new_[2846]_ ;
  assign \new_[5620]_  = \new_[5619]_  | \new_[5616]_ ;
  assign \new_[5621]_  = \new_[5620]_  | \new_[5613]_ ;
  assign \new_[5622]_  = \new_[5621]_  | \new_[5606]_ ;
  assign \new_[5626]_  = \new_[2842]_  | \new_[2843]_ ;
  assign \new_[5627]_  = \new_[2844]_  | \new_[5626]_ ;
  assign \new_[5630]_  = \new_[2840]_  | \new_[2841]_ ;
  assign \new_[5633]_  = \new_[2838]_  | \new_[2839]_ ;
  assign \new_[5634]_  = \new_[5633]_  | \new_[5630]_ ;
  assign \new_[5635]_  = \new_[5634]_  | \new_[5627]_ ;
  assign \new_[5638]_  = \new_[2836]_  | \new_[2837]_ ;
  assign \new_[5641]_  = \new_[2834]_  | \new_[2835]_ ;
  assign \new_[5642]_  = \new_[5641]_  | \new_[5638]_ ;
  assign \new_[5645]_  = \new_[2832]_  | \new_[2833]_ ;
  assign \new_[5648]_  = \new_[2830]_  | \new_[2831]_ ;
  assign \new_[5649]_  = \new_[5648]_  | \new_[5645]_ ;
  assign \new_[5650]_  = \new_[5649]_  | \new_[5642]_ ;
  assign \new_[5651]_  = \new_[5650]_  | \new_[5635]_ ;
  assign \new_[5652]_  = \new_[5651]_  | \new_[5622]_ ;
  assign \new_[5653]_  = \new_[5652]_  | \new_[5593]_ ;
  assign \new_[5654]_  = \new_[5653]_  | \new_[5536]_ ;
  assign \new_[5655]_  = \new_[5654]_  | \new_[5419]_ ;
  assign \new_[5656]_  = \new_[5655]_  | \new_[5184]_ ;
  assign \new_[5657]_  = \new_[5656]_  | \new_[4713]_ ;
  assign \new_[5661]_  = \new_[2827]_  | \new_[2828]_ ;
  assign \new_[5662]_  = \new_[2829]_  | \new_[5661]_ ;
  assign \new_[5665]_  = \new_[2825]_  | \new_[2826]_ ;
  assign \new_[5668]_  = \new_[2823]_  | \new_[2824]_ ;
  assign \new_[5669]_  = \new_[5668]_  | \new_[5665]_ ;
  assign \new_[5670]_  = \new_[5669]_  | \new_[5662]_ ;
  assign \new_[5674]_  = \new_[2820]_  | \new_[2821]_ ;
  assign \new_[5675]_  = \new_[2822]_  | \new_[5674]_ ;
  assign \new_[5678]_  = \new_[2818]_  | \new_[2819]_ ;
  assign \new_[5681]_  = \new_[2816]_  | \new_[2817]_ ;
  assign \new_[5682]_  = \new_[5681]_  | \new_[5678]_ ;
  assign \new_[5683]_  = \new_[5682]_  | \new_[5675]_ ;
  assign \new_[5684]_  = \new_[5683]_  | \new_[5670]_ ;
  assign \new_[5688]_  = \new_[2813]_  | \new_[2814]_ ;
  assign \new_[5689]_  = \new_[2815]_  | \new_[5688]_ ;
  assign \new_[5692]_  = \new_[2811]_  | \new_[2812]_ ;
  assign \new_[5695]_  = \new_[2809]_  | \new_[2810]_ ;
  assign \new_[5696]_  = \new_[5695]_  | \new_[5692]_ ;
  assign \new_[5697]_  = \new_[5696]_  | \new_[5689]_ ;
  assign \new_[5700]_  = \new_[2807]_  | \new_[2808]_ ;
  assign \new_[5703]_  = \new_[2805]_  | \new_[2806]_ ;
  assign \new_[5704]_  = \new_[5703]_  | \new_[5700]_ ;
  assign \new_[5707]_  = \new_[2803]_  | \new_[2804]_ ;
  assign \new_[5710]_  = \new_[2801]_  | \new_[2802]_ ;
  assign \new_[5711]_  = \new_[5710]_  | \new_[5707]_ ;
  assign \new_[5712]_  = \new_[5711]_  | \new_[5704]_ ;
  assign \new_[5713]_  = \new_[5712]_  | \new_[5697]_ ;
  assign \new_[5714]_  = \new_[5713]_  | \new_[5684]_ ;
  assign \new_[5718]_  = \new_[2798]_  | \new_[2799]_ ;
  assign \new_[5719]_  = \new_[2800]_  | \new_[5718]_ ;
  assign \new_[5722]_  = \new_[2796]_  | \new_[2797]_ ;
  assign \new_[5725]_  = \new_[2794]_  | \new_[2795]_ ;
  assign \new_[5726]_  = \new_[5725]_  | \new_[5722]_ ;
  assign \new_[5727]_  = \new_[5726]_  | \new_[5719]_ ;
  assign \new_[5731]_  = \new_[2791]_  | \new_[2792]_ ;
  assign \new_[5732]_  = \new_[2793]_  | \new_[5731]_ ;
  assign \new_[5735]_  = \new_[2789]_  | \new_[2790]_ ;
  assign \new_[5738]_  = \new_[2787]_  | \new_[2788]_ ;
  assign \new_[5739]_  = \new_[5738]_  | \new_[5735]_ ;
  assign \new_[5740]_  = \new_[5739]_  | \new_[5732]_ ;
  assign \new_[5741]_  = \new_[5740]_  | \new_[5727]_ ;
  assign \new_[5745]_  = \new_[2784]_  | \new_[2785]_ ;
  assign \new_[5746]_  = \new_[2786]_  | \new_[5745]_ ;
  assign \new_[5749]_  = \new_[2782]_  | \new_[2783]_ ;
  assign \new_[5752]_  = \new_[2780]_  | \new_[2781]_ ;
  assign \new_[5753]_  = \new_[5752]_  | \new_[5749]_ ;
  assign \new_[5754]_  = \new_[5753]_  | \new_[5746]_ ;
  assign \new_[5757]_  = \new_[2778]_  | \new_[2779]_ ;
  assign \new_[5760]_  = \new_[2776]_  | \new_[2777]_ ;
  assign \new_[5761]_  = \new_[5760]_  | \new_[5757]_ ;
  assign \new_[5764]_  = \new_[2774]_  | \new_[2775]_ ;
  assign \new_[5767]_  = \new_[2772]_  | \new_[2773]_ ;
  assign \new_[5768]_  = \new_[5767]_  | \new_[5764]_ ;
  assign \new_[5769]_  = \new_[5768]_  | \new_[5761]_ ;
  assign \new_[5770]_  = \new_[5769]_  | \new_[5754]_ ;
  assign \new_[5771]_  = \new_[5770]_  | \new_[5741]_ ;
  assign \new_[5772]_  = \new_[5771]_  | \new_[5714]_ ;
  assign \new_[5776]_  = \new_[2769]_  | \new_[2770]_ ;
  assign \new_[5777]_  = \new_[2771]_  | \new_[5776]_ ;
  assign \new_[5780]_  = \new_[2767]_  | \new_[2768]_ ;
  assign \new_[5783]_  = \new_[2765]_  | \new_[2766]_ ;
  assign \new_[5784]_  = \new_[5783]_  | \new_[5780]_ ;
  assign \new_[5785]_  = \new_[5784]_  | \new_[5777]_ ;
  assign \new_[5789]_  = \new_[2762]_  | \new_[2763]_ ;
  assign \new_[5790]_  = \new_[2764]_  | \new_[5789]_ ;
  assign \new_[5793]_  = \new_[2760]_  | \new_[2761]_ ;
  assign \new_[5796]_  = \new_[2758]_  | \new_[2759]_ ;
  assign \new_[5797]_  = \new_[5796]_  | \new_[5793]_ ;
  assign \new_[5798]_  = \new_[5797]_  | \new_[5790]_ ;
  assign \new_[5799]_  = \new_[5798]_  | \new_[5785]_ ;
  assign \new_[5803]_  = \new_[2755]_  | \new_[2756]_ ;
  assign \new_[5804]_  = \new_[2757]_  | \new_[5803]_ ;
  assign \new_[5807]_  = \new_[2753]_  | \new_[2754]_ ;
  assign \new_[5810]_  = \new_[2751]_  | \new_[2752]_ ;
  assign \new_[5811]_  = \new_[5810]_  | \new_[5807]_ ;
  assign \new_[5812]_  = \new_[5811]_  | \new_[5804]_ ;
  assign \new_[5815]_  = \new_[2749]_  | \new_[2750]_ ;
  assign \new_[5818]_  = \new_[2747]_  | \new_[2748]_ ;
  assign \new_[5819]_  = \new_[5818]_  | \new_[5815]_ ;
  assign \new_[5822]_  = \new_[2745]_  | \new_[2746]_ ;
  assign \new_[5825]_  = \new_[2743]_  | \new_[2744]_ ;
  assign \new_[5826]_  = \new_[5825]_  | \new_[5822]_ ;
  assign \new_[5827]_  = \new_[5826]_  | \new_[5819]_ ;
  assign \new_[5828]_  = \new_[5827]_  | \new_[5812]_ ;
  assign \new_[5829]_  = \new_[5828]_  | \new_[5799]_ ;
  assign \new_[5833]_  = \new_[2740]_  | \new_[2741]_ ;
  assign \new_[5834]_  = \new_[2742]_  | \new_[5833]_ ;
  assign \new_[5837]_  = \new_[2738]_  | \new_[2739]_ ;
  assign \new_[5840]_  = \new_[2736]_  | \new_[2737]_ ;
  assign \new_[5841]_  = \new_[5840]_  | \new_[5837]_ ;
  assign \new_[5842]_  = \new_[5841]_  | \new_[5834]_ ;
  assign \new_[5845]_  = \new_[2734]_  | \new_[2735]_ ;
  assign \new_[5848]_  = \new_[2732]_  | \new_[2733]_ ;
  assign \new_[5849]_  = \new_[5848]_  | \new_[5845]_ ;
  assign \new_[5852]_  = \new_[2730]_  | \new_[2731]_ ;
  assign \new_[5855]_  = \new_[2728]_  | \new_[2729]_ ;
  assign \new_[5856]_  = \new_[5855]_  | \new_[5852]_ ;
  assign \new_[5857]_  = \new_[5856]_  | \new_[5849]_ ;
  assign \new_[5858]_  = \new_[5857]_  | \new_[5842]_ ;
  assign \new_[5862]_  = \new_[2725]_  | \new_[2726]_ ;
  assign \new_[5863]_  = \new_[2727]_  | \new_[5862]_ ;
  assign \new_[5866]_  = \new_[2723]_  | \new_[2724]_ ;
  assign \new_[5869]_  = \new_[2721]_  | \new_[2722]_ ;
  assign \new_[5870]_  = \new_[5869]_  | \new_[5866]_ ;
  assign \new_[5871]_  = \new_[5870]_  | \new_[5863]_ ;
  assign \new_[5874]_  = \new_[2719]_  | \new_[2720]_ ;
  assign \new_[5877]_  = \new_[2717]_  | \new_[2718]_ ;
  assign \new_[5878]_  = \new_[5877]_  | \new_[5874]_ ;
  assign \new_[5881]_  = \new_[2715]_  | \new_[2716]_ ;
  assign \new_[5884]_  = \new_[2713]_  | \new_[2714]_ ;
  assign \new_[5885]_  = \new_[5884]_  | \new_[5881]_ ;
  assign \new_[5886]_  = \new_[5885]_  | \new_[5878]_ ;
  assign \new_[5887]_  = \new_[5886]_  | \new_[5871]_ ;
  assign \new_[5888]_  = \new_[5887]_  | \new_[5858]_ ;
  assign \new_[5889]_  = \new_[5888]_  | \new_[5829]_ ;
  assign \new_[5890]_  = \new_[5889]_  | \new_[5772]_ ;
  assign \new_[5894]_  = \new_[2710]_  | \new_[2711]_ ;
  assign \new_[5895]_  = \new_[2712]_  | \new_[5894]_ ;
  assign \new_[5898]_  = \new_[2708]_  | \new_[2709]_ ;
  assign \new_[5901]_  = \new_[2706]_  | \new_[2707]_ ;
  assign \new_[5902]_  = \new_[5901]_  | \new_[5898]_ ;
  assign \new_[5903]_  = \new_[5902]_  | \new_[5895]_ ;
  assign \new_[5907]_  = \new_[2703]_  | \new_[2704]_ ;
  assign \new_[5908]_  = \new_[2705]_  | \new_[5907]_ ;
  assign \new_[5911]_  = \new_[2701]_  | \new_[2702]_ ;
  assign \new_[5914]_  = \new_[2699]_  | \new_[2700]_ ;
  assign \new_[5915]_  = \new_[5914]_  | \new_[5911]_ ;
  assign \new_[5916]_  = \new_[5915]_  | \new_[5908]_ ;
  assign \new_[5917]_  = \new_[5916]_  | \new_[5903]_ ;
  assign \new_[5921]_  = \new_[2696]_  | \new_[2697]_ ;
  assign \new_[5922]_  = \new_[2698]_  | \new_[5921]_ ;
  assign \new_[5925]_  = \new_[2694]_  | \new_[2695]_ ;
  assign \new_[5928]_  = \new_[2692]_  | \new_[2693]_ ;
  assign \new_[5929]_  = \new_[5928]_  | \new_[5925]_ ;
  assign \new_[5930]_  = \new_[5929]_  | \new_[5922]_ ;
  assign \new_[5933]_  = \new_[2690]_  | \new_[2691]_ ;
  assign \new_[5936]_  = \new_[2688]_  | \new_[2689]_ ;
  assign \new_[5937]_  = \new_[5936]_  | \new_[5933]_ ;
  assign \new_[5940]_  = \new_[2686]_  | \new_[2687]_ ;
  assign \new_[5943]_  = \new_[2684]_  | \new_[2685]_ ;
  assign \new_[5944]_  = \new_[5943]_  | \new_[5940]_ ;
  assign \new_[5945]_  = \new_[5944]_  | \new_[5937]_ ;
  assign \new_[5946]_  = \new_[5945]_  | \new_[5930]_ ;
  assign \new_[5947]_  = \new_[5946]_  | \new_[5917]_ ;
  assign \new_[5951]_  = \new_[2681]_  | \new_[2682]_ ;
  assign \new_[5952]_  = \new_[2683]_  | \new_[5951]_ ;
  assign \new_[5955]_  = \new_[2679]_  | \new_[2680]_ ;
  assign \new_[5958]_  = \new_[2677]_  | \new_[2678]_ ;
  assign \new_[5959]_  = \new_[5958]_  | \new_[5955]_ ;
  assign \new_[5960]_  = \new_[5959]_  | \new_[5952]_ ;
  assign \new_[5963]_  = \new_[2675]_  | \new_[2676]_ ;
  assign \new_[5966]_  = \new_[2673]_  | \new_[2674]_ ;
  assign \new_[5967]_  = \new_[5966]_  | \new_[5963]_ ;
  assign \new_[5970]_  = \new_[2671]_  | \new_[2672]_ ;
  assign \new_[5973]_  = \new_[2669]_  | \new_[2670]_ ;
  assign \new_[5974]_  = \new_[5973]_  | \new_[5970]_ ;
  assign \new_[5975]_  = \new_[5974]_  | \new_[5967]_ ;
  assign \new_[5976]_  = \new_[5975]_  | \new_[5960]_ ;
  assign \new_[5980]_  = \new_[2666]_  | \new_[2667]_ ;
  assign \new_[5981]_  = \new_[2668]_  | \new_[5980]_ ;
  assign \new_[5984]_  = \new_[2664]_  | \new_[2665]_ ;
  assign \new_[5987]_  = \new_[2662]_  | \new_[2663]_ ;
  assign \new_[5988]_  = \new_[5987]_  | \new_[5984]_ ;
  assign \new_[5989]_  = \new_[5988]_  | \new_[5981]_ ;
  assign \new_[5992]_  = \new_[2660]_  | \new_[2661]_ ;
  assign \new_[5995]_  = \new_[2658]_  | \new_[2659]_ ;
  assign \new_[5996]_  = \new_[5995]_  | \new_[5992]_ ;
  assign \new_[5999]_  = \new_[2656]_  | \new_[2657]_ ;
  assign \new_[6002]_  = \new_[2654]_  | \new_[2655]_ ;
  assign \new_[6003]_  = \new_[6002]_  | \new_[5999]_ ;
  assign \new_[6004]_  = \new_[6003]_  | \new_[5996]_ ;
  assign \new_[6005]_  = \new_[6004]_  | \new_[5989]_ ;
  assign \new_[6006]_  = \new_[6005]_  | \new_[5976]_ ;
  assign \new_[6007]_  = \new_[6006]_  | \new_[5947]_ ;
  assign \new_[6011]_  = \new_[2651]_  | \new_[2652]_ ;
  assign \new_[6012]_  = \new_[2653]_  | \new_[6011]_ ;
  assign \new_[6015]_  = \new_[2649]_  | \new_[2650]_ ;
  assign \new_[6018]_  = \new_[2647]_  | \new_[2648]_ ;
  assign \new_[6019]_  = \new_[6018]_  | \new_[6015]_ ;
  assign \new_[6020]_  = \new_[6019]_  | \new_[6012]_ ;
  assign \new_[6024]_  = \new_[2644]_  | \new_[2645]_ ;
  assign \new_[6025]_  = \new_[2646]_  | \new_[6024]_ ;
  assign \new_[6028]_  = \new_[2642]_  | \new_[2643]_ ;
  assign \new_[6031]_  = \new_[2640]_  | \new_[2641]_ ;
  assign \new_[6032]_  = \new_[6031]_  | \new_[6028]_ ;
  assign \new_[6033]_  = \new_[6032]_  | \new_[6025]_ ;
  assign \new_[6034]_  = \new_[6033]_  | \new_[6020]_ ;
  assign \new_[6038]_  = \new_[2637]_  | \new_[2638]_ ;
  assign \new_[6039]_  = \new_[2639]_  | \new_[6038]_ ;
  assign \new_[6042]_  = \new_[2635]_  | \new_[2636]_ ;
  assign \new_[6045]_  = \new_[2633]_  | \new_[2634]_ ;
  assign \new_[6046]_  = \new_[6045]_  | \new_[6042]_ ;
  assign \new_[6047]_  = \new_[6046]_  | \new_[6039]_ ;
  assign \new_[6050]_  = \new_[2631]_  | \new_[2632]_ ;
  assign \new_[6053]_  = \new_[2629]_  | \new_[2630]_ ;
  assign \new_[6054]_  = \new_[6053]_  | \new_[6050]_ ;
  assign \new_[6057]_  = \new_[2627]_  | \new_[2628]_ ;
  assign \new_[6060]_  = \new_[2625]_  | \new_[2626]_ ;
  assign \new_[6061]_  = \new_[6060]_  | \new_[6057]_ ;
  assign \new_[6062]_  = \new_[6061]_  | \new_[6054]_ ;
  assign \new_[6063]_  = \new_[6062]_  | \new_[6047]_ ;
  assign \new_[6064]_  = \new_[6063]_  | \new_[6034]_ ;
  assign \new_[6068]_  = \new_[2622]_  | \new_[2623]_ ;
  assign \new_[6069]_  = \new_[2624]_  | \new_[6068]_ ;
  assign \new_[6072]_  = \new_[2620]_  | \new_[2621]_ ;
  assign \new_[6075]_  = \new_[2618]_  | \new_[2619]_ ;
  assign \new_[6076]_  = \new_[6075]_  | \new_[6072]_ ;
  assign \new_[6077]_  = \new_[6076]_  | \new_[6069]_ ;
  assign \new_[6080]_  = \new_[2616]_  | \new_[2617]_ ;
  assign \new_[6083]_  = \new_[2614]_  | \new_[2615]_ ;
  assign \new_[6084]_  = \new_[6083]_  | \new_[6080]_ ;
  assign \new_[6087]_  = \new_[2612]_  | \new_[2613]_ ;
  assign \new_[6090]_  = \new_[2610]_  | \new_[2611]_ ;
  assign \new_[6091]_  = \new_[6090]_  | \new_[6087]_ ;
  assign \new_[6092]_  = \new_[6091]_  | \new_[6084]_ ;
  assign \new_[6093]_  = \new_[6092]_  | \new_[6077]_ ;
  assign \new_[6097]_  = \new_[2607]_  | \new_[2608]_ ;
  assign \new_[6098]_  = \new_[2609]_  | \new_[6097]_ ;
  assign \new_[6101]_  = \new_[2605]_  | \new_[2606]_ ;
  assign \new_[6104]_  = \new_[2603]_  | \new_[2604]_ ;
  assign \new_[6105]_  = \new_[6104]_  | \new_[6101]_ ;
  assign \new_[6106]_  = \new_[6105]_  | \new_[6098]_ ;
  assign \new_[6109]_  = \new_[2601]_  | \new_[2602]_ ;
  assign \new_[6112]_  = \new_[2599]_  | \new_[2600]_ ;
  assign \new_[6113]_  = \new_[6112]_  | \new_[6109]_ ;
  assign \new_[6116]_  = \new_[2597]_  | \new_[2598]_ ;
  assign \new_[6119]_  = \new_[2595]_  | \new_[2596]_ ;
  assign \new_[6120]_  = \new_[6119]_  | \new_[6116]_ ;
  assign \new_[6121]_  = \new_[6120]_  | \new_[6113]_ ;
  assign \new_[6122]_  = \new_[6121]_  | \new_[6106]_ ;
  assign \new_[6123]_  = \new_[6122]_  | \new_[6093]_ ;
  assign \new_[6124]_  = \new_[6123]_  | \new_[6064]_ ;
  assign \new_[6125]_  = \new_[6124]_  | \new_[6007]_ ;
  assign \new_[6126]_  = \new_[6125]_  | \new_[5890]_ ;
  assign \new_[6130]_  = \new_[2592]_  | \new_[2593]_ ;
  assign \new_[6131]_  = \new_[2594]_  | \new_[6130]_ ;
  assign \new_[6134]_  = \new_[2590]_  | \new_[2591]_ ;
  assign \new_[6137]_  = \new_[2588]_  | \new_[2589]_ ;
  assign \new_[6138]_  = \new_[6137]_  | \new_[6134]_ ;
  assign \new_[6139]_  = \new_[6138]_  | \new_[6131]_ ;
  assign \new_[6143]_  = \new_[2585]_  | \new_[2586]_ ;
  assign \new_[6144]_  = \new_[2587]_  | \new_[6143]_ ;
  assign \new_[6147]_  = \new_[2583]_  | \new_[2584]_ ;
  assign \new_[6150]_  = \new_[2581]_  | \new_[2582]_ ;
  assign \new_[6151]_  = \new_[6150]_  | \new_[6147]_ ;
  assign \new_[6152]_  = \new_[6151]_  | \new_[6144]_ ;
  assign \new_[6153]_  = \new_[6152]_  | \new_[6139]_ ;
  assign \new_[6157]_  = \new_[2578]_  | \new_[2579]_ ;
  assign \new_[6158]_  = \new_[2580]_  | \new_[6157]_ ;
  assign \new_[6161]_  = \new_[2576]_  | \new_[2577]_ ;
  assign \new_[6164]_  = \new_[2574]_  | \new_[2575]_ ;
  assign \new_[6165]_  = \new_[6164]_  | \new_[6161]_ ;
  assign \new_[6166]_  = \new_[6165]_  | \new_[6158]_ ;
  assign \new_[6169]_  = \new_[2572]_  | \new_[2573]_ ;
  assign \new_[6172]_  = \new_[2570]_  | \new_[2571]_ ;
  assign \new_[6173]_  = \new_[6172]_  | \new_[6169]_ ;
  assign \new_[6176]_  = \new_[2568]_  | \new_[2569]_ ;
  assign \new_[6179]_  = \new_[2566]_  | \new_[2567]_ ;
  assign \new_[6180]_  = \new_[6179]_  | \new_[6176]_ ;
  assign \new_[6181]_  = \new_[6180]_  | \new_[6173]_ ;
  assign \new_[6182]_  = \new_[6181]_  | \new_[6166]_ ;
  assign \new_[6183]_  = \new_[6182]_  | \new_[6153]_ ;
  assign \new_[6187]_  = \new_[2563]_  | \new_[2564]_ ;
  assign \new_[6188]_  = \new_[2565]_  | \new_[6187]_ ;
  assign \new_[6191]_  = \new_[2561]_  | \new_[2562]_ ;
  assign \new_[6194]_  = \new_[2559]_  | \new_[2560]_ ;
  assign \new_[6195]_  = \new_[6194]_  | \new_[6191]_ ;
  assign \new_[6196]_  = \new_[6195]_  | \new_[6188]_ ;
  assign \new_[6199]_  = \new_[2557]_  | \new_[2558]_ ;
  assign \new_[6202]_  = \new_[2555]_  | \new_[2556]_ ;
  assign \new_[6203]_  = \new_[6202]_  | \new_[6199]_ ;
  assign \new_[6206]_  = \new_[2553]_  | \new_[2554]_ ;
  assign \new_[6209]_  = \new_[2551]_  | \new_[2552]_ ;
  assign \new_[6210]_  = \new_[6209]_  | \new_[6206]_ ;
  assign \new_[6211]_  = \new_[6210]_  | \new_[6203]_ ;
  assign \new_[6212]_  = \new_[6211]_  | \new_[6196]_ ;
  assign \new_[6216]_  = \new_[2548]_  | \new_[2549]_ ;
  assign \new_[6217]_  = \new_[2550]_  | \new_[6216]_ ;
  assign \new_[6220]_  = \new_[2546]_  | \new_[2547]_ ;
  assign \new_[6223]_  = \new_[2544]_  | \new_[2545]_ ;
  assign \new_[6224]_  = \new_[6223]_  | \new_[6220]_ ;
  assign \new_[6225]_  = \new_[6224]_  | \new_[6217]_ ;
  assign \new_[6228]_  = \new_[2542]_  | \new_[2543]_ ;
  assign \new_[6231]_  = \new_[2540]_  | \new_[2541]_ ;
  assign \new_[6232]_  = \new_[6231]_  | \new_[6228]_ ;
  assign \new_[6235]_  = \new_[2538]_  | \new_[2539]_ ;
  assign \new_[6238]_  = \new_[2536]_  | \new_[2537]_ ;
  assign \new_[6239]_  = \new_[6238]_  | \new_[6235]_ ;
  assign \new_[6240]_  = \new_[6239]_  | \new_[6232]_ ;
  assign \new_[6241]_  = \new_[6240]_  | \new_[6225]_ ;
  assign \new_[6242]_  = \new_[6241]_  | \new_[6212]_ ;
  assign \new_[6243]_  = \new_[6242]_  | \new_[6183]_ ;
  assign \new_[6247]_  = \new_[2533]_  | \new_[2534]_ ;
  assign \new_[6248]_  = \new_[2535]_  | \new_[6247]_ ;
  assign \new_[6251]_  = \new_[2531]_  | \new_[2532]_ ;
  assign \new_[6254]_  = \new_[2529]_  | \new_[2530]_ ;
  assign \new_[6255]_  = \new_[6254]_  | \new_[6251]_ ;
  assign \new_[6256]_  = \new_[6255]_  | \new_[6248]_ ;
  assign \new_[6260]_  = \new_[2526]_  | \new_[2527]_ ;
  assign \new_[6261]_  = \new_[2528]_  | \new_[6260]_ ;
  assign \new_[6264]_  = \new_[2524]_  | \new_[2525]_ ;
  assign \new_[6267]_  = \new_[2522]_  | \new_[2523]_ ;
  assign \new_[6268]_  = \new_[6267]_  | \new_[6264]_ ;
  assign \new_[6269]_  = \new_[6268]_  | \new_[6261]_ ;
  assign \new_[6270]_  = \new_[6269]_  | \new_[6256]_ ;
  assign \new_[6274]_  = \new_[2519]_  | \new_[2520]_ ;
  assign \new_[6275]_  = \new_[2521]_  | \new_[6274]_ ;
  assign \new_[6278]_  = \new_[2517]_  | \new_[2518]_ ;
  assign \new_[6281]_  = \new_[2515]_  | \new_[2516]_ ;
  assign \new_[6282]_  = \new_[6281]_  | \new_[6278]_ ;
  assign \new_[6283]_  = \new_[6282]_  | \new_[6275]_ ;
  assign \new_[6286]_  = \new_[2513]_  | \new_[2514]_ ;
  assign \new_[6289]_  = \new_[2511]_  | \new_[2512]_ ;
  assign \new_[6290]_  = \new_[6289]_  | \new_[6286]_ ;
  assign \new_[6293]_  = \new_[2509]_  | \new_[2510]_ ;
  assign \new_[6296]_  = \new_[2507]_  | \new_[2508]_ ;
  assign \new_[6297]_  = \new_[6296]_  | \new_[6293]_ ;
  assign \new_[6298]_  = \new_[6297]_  | \new_[6290]_ ;
  assign \new_[6299]_  = \new_[6298]_  | \new_[6283]_ ;
  assign \new_[6300]_  = \new_[6299]_  | \new_[6270]_ ;
  assign \new_[6304]_  = \new_[2504]_  | \new_[2505]_ ;
  assign \new_[6305]_  = \new_[2506]_  | \new_[6304]_ ;
  assign \new_[6308]_  = \new_[2502]_  | \new_[2503]_ ;
  assign \new_[6311]_  = \new_[2500]_  | \new_[2501]_ ;
  assign \new_[6312]_  = \new_[6311]_  | \new_[6308]_ ;
  assign \new_[6313]_  = \new_[6312]_  | \new_[6305]_ ;
  assign \new_[6316]_  = \new_[2498]_  | \new_[2499]_ ;
  assign \new_[6319]_  = \new_[2496]_  | \new_[2497]_ ;
  assign \new_[6320]_  = \new_[6319]_  | \new_[6316]_ ;
  assign \new_[6323]_  = \new_[2494]_  | \new_[2495]_ ;
  assign \new_[6326]_  = \new_[2492]_  | \new_[2493]_ ;
  assign \new_[6327]_  = \new_[6326]_  | \new_[6323]_ ;
  assign \new_[6328]_  = \new_[6327]_  | \new_[6320]_ ;
  assign \new_[6329]_  = \new_[6328]_  | \new_[6313]_ ;
  assign \new_[6333]_  = \new_[2489]_  | \new_[2490]_ ;
  assign \new_[6334]_  = \new_[2491]_  | \new_[6333]_ ;
  assign \new_[6337]_  = \new_[2487]_  | \new_[2488]_ ;
  assign \new_[6340]_  = \new_[2485]_  | \new_[2486]_ ;
  assign \new_[6341]_  = \new_[6340]_  | \new_[6337]_ ;
  assign \new_[6342]_  = \new_[6341]_  | \new_[6334]_ ;
  assign \new_[6345]_  = \new_[2483]_  | \new_[2484]_ ;
  assign \new_[6348]_  = \new_[2481]_  | \new_[2482]_ ;
  assign \new_[6349]_  = \new_[6348]_  | \new_[6345]_ ;
  assign \new_[6352]_  = \new_[2479]_  | \new_[2480]_ ;
  assign \new_[6355]_  = \new_[2477]_  | \new_[2478]_ ;
  assign \new_[6356]_  = \new_[6355]_  | \new_[6352]_ ;
  assign \new_[6357]_  = \new_[6356]_  | \new_[6349]_ ;
  assign \new_[6358]_  = \new_[6357]_  | \new_[6342]_ ;
  assign \new_[6359]_  = \new_[6358]_  | \new_[6329]_ ;
  assign \new_[6360]_  = \new_[6359]_  | \new_[6300]_ ;
  assign \new_[6361]_  = \new_[6360]_  | \new_[6243]_ ;
  assign \new_[6365]_  = \new_[2474]_  | \new_[2475]_ ;
  assign \new_[6366]_  = \new_[2476]_  | \new_[6365]_ ;
  assign \new_[6369]_  = \new_[2472]_  | \new_[2473]_ ;
  assign \new_[6372]_  = \new_[2470]_  | \new_[2471]_ ;
  assign \new_[6373]_  = \new_[6372]_  | \new_[6369]_ ;
  assign \new_[6374]_  = \new_[6373]_  | \new_[6366]_ ;
  assign \new_[6378]_  = \new_[2467]_  | \new_[2468]_ ;
  assign \new_[6379]_  = \new_[2469]_  | \new_[6378]_ ;
  assign \new_[6382]_  = \new_[2465]_  | \new_[2466]_ ;
  assign \new_[6385]_  = \new_[2463]_  | \new_[2464]_ ;
  assign \new_[6386]_  = \new_[6385]_  | \new_[6382]_ ;
  assign \new_[6387]_  = \new_[6386]_  | \new_[6379]_ ;
  assign \new_[6388]_  = \new_[6387]_  | \new_[6374]_ ;
  assign \new_[6392]_  = \new_[2460]_  | \new_[2461]_ ;
  assign \new_[6393]_  = \new_[2462]_  | \new_[6392]_ ;
  assign \new_[6396]_  = \new_[2458]_  | \new_[2459]_ ;
  assign \new_[6399]_  = \new_[2456]_  | \new_[2457]_ ;
  assign \new_[6400]_  = \new_[6399]_  | \new_[6396]_ ;
  assign \new_[6401]_  = \new_[6400]_  | \new_[6393]_ ;
  assign \new_[6404]_  = \new_[2454]_  | \new_[2455]_ ;
  assign \new_[6407]_  = \new_[2452]_  | \new_[2453]_ ;
  assign \new_[6408]_  = \new_[6407]_  | \new_[6404]_ ;
  assign \new_[6411]_  = \new_[2450]_  | \new_[2451]_ ;
  assign \new_[6414]_  = \new_[2448]_  | \new_[2449]_ ;
  assign \new_[6415]_  = \new_[6414]_  | \new_[6411]_ ;
  assign \new_[6416]_  = \new_[6415]_  | \new_[6408]_ ;
  assign \new_[6417]_  = \new_[6416]_  | \new_[6401]_ ;
  assign \new_[6418]_  = \new_[6417]_  | \new_[6388]_ ;
  assign \new_[6422]_  = \new_[2445]_  | \new_[2446]_ ;
  assign \new_[6423]_  = \new_[2447]_  | \new_[6422]_ ;
  assign \new_[6426]_  = \new_[2443]_  | \new_[2444]_ ;
  assign \new_[6429]_  = \new_[2441]_  | \new_[2442]_ ;
  assign \new_[6430]_  = \new_[6429]_  | \new_[6426]_ ;
  assign \new_[6431]_  = \new_[6430]_  | \new_[6423]_ ;
  assign \new_[6434]_  = \new_[2439]_  | \new_[2440]_ ;
  assign \new_[6437]_  = \new_[2437]_  | \new_[2438]_ ;
  assign \new_[6438]_  = \new_[6437]_  | \new_[6434]_ ;
  assign \new_[6441]_  = \new_[2435]_  | \new_[2436]_ ;
  assign \new_[6444]_  = \new_[2433]_  | \new_[2434]_ ;
  assign \new_[6445]_  = \new_[6444]_  | \new_[6441]_ ;
  assign \new_[6446]_  = \new_[6445]_  | \new_[6438]_ ;
  assign \new_[6447]_  = \new_[6446]_  | \new_[6431]_ ;
  assign \new_[6451]_  = \new_[2430]_  | \new_[2431]_ ;
  assign \new_[6452]_  = \new_[2432]_  | \new_[6451]_ ;
  assign \new_[6455]_  = \new_[2428]_  | \new_[2429]_ ;
  assign \new_[6458]_  = \new_[2426]_  | \new_[2427]_ ;
  assign \new_[6459]_  = \new_[6458]_  | \new_[6455]_ ;
  assign \new_[6460]_  = \new_[6459]_  | \new_[6452]_ ;
  assign \new_[6463]_  = \new_[2424]_  | \new_[2425]_ ;
  assign \new_[6466]_  = \new_[2422]_  | \new_[2423]_ ;
  assign \new_[6467]_  = \new_[6466]_  | \new_[6463]_ ;
  assign \new_[6470]_  = \new_[2420]_  | \new_[2421]_ ;
  assign \new_[6473]_  = \new_[2418]_  | \new_[2419]_ ;
  assign \new_[6474]_  = \new_[6473]_  | \new_[6470]_ ;
  assign \new_[6475]_  = \new_[6474]_  | \new_[6467]_ ;
  assign \new_[6476]_  = \new_[6475]_  | \new_[6460]_ ;
  assign \new_[6477]_  = \new_[6476]_  | \new_[6447]_ ;
  assign \new_[6478]_  = \new_[6477]_  | \new_[6418]_ ;
  assign \new_[6482]_  = \new_[2415]_  | \new_[2416]_ ;
  assign \new_[6483]_  = \new_[2417]_  | \new_[6482]_ ;
  assign \new_[6486]_  = \new_[2413]_  | \new_[2414]_ ;
  assign \new_[6489]_  = \new_[2411]_  | \new_[2412]_ ;
  assign \new_[6490]_  = \new_[6489]_  | \new_[6486]_ ;
  assign \new_[6491]_  = \new_[6490]_  | \new_[6483]_ ;
  assign \new_[6495]_  = \new_[2408]_  | \new_[2409]_ ;
  assign \new_[6496]_  = \new_[2410]_  | \new_[6495]_ ;
  assign \new_[6499]_  = \new_[2406]_  | \new_[2407]_ ;
  assign \new_[6502]_  = \new_[2404]_  | \new_[2405]_ ;
  assign \new_[6503]_  = \new_[6502]_  | \new_[6499]_ ;
  assign \new_[6504]_  = \new_[6503]_  | \new_[6496]_ ;
  assign \new_[6505]_  = \new_[6504]_  | \new_[6491]_ ;
  assign \new_[6509]_  = \new_[2401]_  | \new_[2402]_ ;
  assign \new_[6510]_  = \new_[2403]_  | \new_[6509]_ ;
  assign \new_[6513]_  = \new_[2399]_  | \new_[2400]_ ;
  assign \new_[6516]_  = \new_[2397]_  | \new_[2398]_ ;
  assign \new_[6517]_  = \new_[6516]_  | \new_[6513]_ ;
  assign \new_[6518]_  = \new_[6517]_  | \new_[6510]_ ;
  assign \new_[6521]_  = \new_[2395]_  | \new_[2396]_ ;
  assign \new_[6524]_  = \new_[2393]_  | \new_[2394]_ ;
  assign \new_[6525]_  = \new_[6524]_  | \new_[6521]_ ;
  assign \new_[6528]_  = \new_[2391]_  | \new_[2392]_ ;
  assign \new_[6531]_  = \new_[2389]_  | \new_[2390]_ ;
  assign \new_[6532]_  = \new_[6531]_  | \new_[6528]_ ;
  assign \new_[6533]_  = \new_[6532]_  | \new_[6525]_ ;
  assign \new_[6534]_  = \new_[6533]_  | \new_[6518]_ ;
  assign \new_[6535]_  = \new_[6534]_  | \new_[6505]_ ;
  assign \new_[6539]_  = \new_[2386]_  | \new_[2387]_ ;
  assign \new_[6540]_  = \new_[2388]_  | \new_[6539]_ ;
  assign \new_[6543]_  = \new_[2384]_  | \new_[2385]_ ;
  assign \new_[6546]_  = \new_[2382]_  | \new_[2383]_ ;
  assign \new_[6547]_  = \new_[6546]_  | \new_[6543]_ ;
  assign \new_[6548]_  = \new_[6547]_  | \new_[6540]_ ;
  assign \new_[6551]_  = \new_[2380]_  | \new_[2381]_ ;
  assign \new_[6554]_  = \new_[2378]_  | \new_[2379]_ ;
  assign \new_[6555]_  = \new_[6554]_  | \new_[6551]_ ;
  assign \new_[6558]_  = \new_[2376]_  | \new_[2377]_ ;
  assign \new_[6561]_  = \new_[2374]_  | \new_[2375]_ ;
  assign \new_[6562]_  = \new_[6561]_  | \new_[6558]_ ;
  assign \new_[6563]_  = \new_[6562]_  | \new_[6555]_ ;
  assign \new_[6564]_  = \new_[6563]_  | \new_[6548]_ ;
  assign \new_[6568]_  = \new_[2371]_  | \new_[2372]_ ;
  assign \new_[6569]_  = \new_[2373]_  | \new_[6568]_ ;
  assign \new_[6572]_  = \new_[2369]_  | \new_[2370]_ ;
  assign \new_[6575]_  = \new_[2367]_  | \new_[2368]_ ;
  assign \new_[6576]_  = \new_[6575]_  | \new_[6572]_ ;
  assign \new_[6577]_  = \new_[6576]_  | \new_[6569]_ ;
  assign \new_[6580]_  = \new_[2365]_  | \new_[2366]_ ;
  assign \new_[6583]_  = \new_[2363]_  | \new_[2364]_ ;
  assign \new_[6584]_  = \new_[6583]_  | \new_[6580]_ ;
  assign \new_[6587]_  = \new_[2361]_  | \new_[2362]_ ;
  assign \new_[6590]_  = \new_[2359]_  | \new_[2360]_ ;
  assign \new_[6591]_  = \new_[6590]_  | \new_[6587]_ ;
  assign \new_[6592]_  = \new_[6591]_  | \new_[6584]_ ;
  assign \new_[6593]_  = \new_[6592]_  | \new_[6577]_ ;
  assign \new_[6594]_  = \new_[6593]_  | \new_[6564]_ ;
  assign \new_[6595]_  = \new_[6594]_  | \new_[6535]_ ;
  assign \new_[6596]_  = \new_[6595]_  | \new_[6478]_ ;
  assign \new_[6597]_  = \new_[6596]_  | \new_[6361]_ ;
  assign \new_[6598]_  = \new_[6597]_  | \new_[6126]_ ;
  assign \new_[6602]_  = \new_[2356]_  | \new_[2357]_ ;
  assign \new_[6603]_  = \new_[2358]_  | \new_[6602]_ ;
  assign \new_[6606]_  = \new_[2354]_  | \new_[2355]_ ;
  assign \new_[6609]_  = \new_[2352]_  | \new_[2353]_ ;
  assign \new_[6610]_  = \new_[6609]_  | \new_[6606]_ ;
  assign \new_[6611]_  = \new_[6610]_  | \new_[6603]_ ;
  assign \new_[6615]_  = \new_[2349]_  | \new_[2350]_ ;
  assign \new_[6616]_  = \new_[2351]_  | \new_[6615]_ ;
  assign \new_[6619]_  = \new_[2347]_  | \new_[2348]_ ;
  assign \new_[6622]_  = \new_[2345]_  | \new_[2346]_ ;
  assign \new_[6623]_  = \new_[6622]_  | \new_[6619]_ ;
  assign \new_[6624]_  = \new_[6623]_  | \new_[6616]_ ;
  assign \new_[6625]_  = \new_[6624]_  | \new_[6611]_ ;
  assign \new_[6629]_  = \new_[2342]_  | \new_[2343]_ ;
  assign \new_[6630]_  = \new_[2344]_  | \new_[6629]_ ;
  assign \new_[6633]_  = \new_[2340]_  | \new_[2341]_ ;
  assign \new_[6636]_  = \new_[2338]_  | \new_[2339]_ ;
  assign \new_[6637]_  = \new_[6636]_  | \new_[6633]_ ;
  assign \new_[6638]_  = \new_[6637]_  | \new_[6630]_ ;
  assign \new_[6641]_  = \new_[2336]_  | \new_[2337]_ ;
  assign \new_[6644]_  = \new_[2334]_  | \new_[2335]_ ;
  assign \new_[6645]_  = \new_[6644]_  | \new_[6641]_ ;
  assign \new_[6648]_  = \new_[2332]_  | \new_[2333]_ ;
  assign \new_[6651]_  = \new_[2330]_  | \new_[2331]_ ;
  assign \new_[6652]_  = \new_[6651]_  | \new_[6648]_ ;
  assign \new_[6653]_  = \new_[6652]_  | \new_[6645]_ ;
  assign \new_[6654]_  = \new_[6653]_  | \new_[6638]_ ;
  assign \new_[6655]_  = \new_[6654]_  | \new_[6625]_ ;
  assign \new_[6659]_  = \new_[2327]_  | \new_[2328]_ ;
  assign \new_[6660]_  = \new_[2329]_  | \new_[6659]_ ;
  assign \new_[6663]_  = \new_[2325]_  | \new_[2326]_ ;
  assign \new_[6666]_  = \new_[2323]_  | \new_[2324]_ ;
  assign \new_[6667]_  = \new_[6666]_  | \new_[6663]_ ;
  assign \new_[6668]_  = \new_[6667]_  | \new_[6660]_ ;
  assign \new_[6671]_  = \new_[2321]_  | \new_[2322]_ ;
  assign \new_[6674]_  = \new_[2319]_  | \new_[2320]_ ;
  assign \new_[6675]_  = \new_[6674]_  | \new_[6671]_ ;
  assign \new_[6678]_  = \new_[2317]_  | \new_[2318]_ ;
  assign \new_[6681]_  = \new_[2315]_  | \new_[2316]_ ;
  assign \new_[6682]_  = \new_[6681]_  | \new_[6678]_ ;
  assign \new_[6683]_  = \new_[6682]_  | \new_[6675]_ ;
  assign \new_[6684]_  = \new_[6683]_  | \new_[6668]_ ;
  assign \new_[6688]_  = \new_[2312]_  | \new_[2313]_ ;
  assign \new_[6689]_  = \new_[2314]_  | \new_[6688]_ ;
  assign \new_[6692]_  = \new_[2310]_  | \new_[2311]_ ;
  assign \new_[6695]_  = \new_[2308]_  | \new_[2309]_ ;
  assign \new_[6696]_  = \new_[6695]_  | \new_[6692]_ ;
  assign \new_[6697]_  = \new_[6696]_  | \new_[6689]_ ;
  assign \new_[6700]_  = \new_[2306]_  | \new_[2307]_ ;
  assign \new_[6703]_  = \new_[2304]_  | \new_[2305]_ ;
  assign \new_[6704]_  = \new_[6703]_  | \new_[6700]_ ;
  assign \new_[6707]_  = \new_[2302]_  | \new_[2303]_ ;
  assign \new_[6710]_  = \new_[2300]_  | \new_[2301]_ ;
  assign \new_[6711]_  = \new_[6710]_  | \new_[6707]_ ;
  assign \new_[6712]_  = \new_[6711]_  | \new_[6704]_ ;
  assign \new_[6713]_  = \new_[6712]_  | \new_[6697]_ ;
  assign \new_[6714]_  = \new_[6713]_  | \new_[6684]_ ;
  assign \new_[6715]_  = \new_[6714]_  | \new_[6655]_ ;
  assign \new_[6719]_  = \new_[2297]_  | \new_[2298]_ ;
  assign \new_[6720]_  = \new_[2299]_  | \new_[6719]_ ;
  assign \new_[6723]_  = \new_[2295]_  | \new_[2296]_ ;
  assign \new_[6726]_  = \new_[2293]_  | \new_[2294]_ ;
  assign \new_[6727]_  = \new_[6726]_  | \new_[6723]_ ;
  assign \new_[6728]_  = \new_[6727]_  | \new_[6720]_ ;
  assign \new_[6732]_  = \new_[2290]_  | \new_[2291]_ ;
  assign \new_[6733]_  = \new_[2292]_  | \new_[6732]_ ;
  assign \new_[6736]_  = \new_[2288]_  | \new_[2289]_ ;
  assign \new_[6739]_  = \new_[2286]_  | \new_[2287]_ ;
  assign \new_[6740]_  = \new_[6739]_  | \new_[6736]_ ;
  assign \new_[6741]_  = \new_[6740]_  | \new_[6733]_ ;
  assign \new_[6742]_  = \new_[6741]_  | \new_[6728]_ ;
  assign \new_[6746]_  = \new_[2283]_  | \new_[2284]_ ;
  assign \new_[6747]_  = \new_[2285]_  | \new_[6746]_ ;
  assign \new_[6750]_  = \new_[2281]_  | \new_[2282]_ ;
  assign \new_[6753]_  = \new_[2279]_  | \new_[2280]_ ;
  assign \new_[6754]_  = \new_[6753]_  | \new_[6750]_ ;
  assign \new_[6755]_  = \new_[6754]_  | \new_[6747]_ ;
  assign \new_[6758]_  = \new_[2277]_  | \new_[2278]_ ;
  assign \new_[6761]_  = \new_[2275]_  | \new_[2276]_ ;
  assign \new_[6762]_  = \new_[6761]_  | \new_[6758]_ ;
  assign \new_[6765]_  = \new_[2273]_  | \new_[2274]_ ;
  assign \new_[6768]_  = \new_[2271]_  | \new_[2272]_ ;
  assign \new_[6769]_  = \new_[6768]_  | \new_[6765]_ ;
  assign \new_[6770]_  = \new_[6769]_  | \new_[6762]_ ;
  assign \new_[6771]_  = \new_[6770]_  | \new_[6755]_ ;
  assign \new_[6772]_  = \new_[6771]_  | \new_[6742]_ ;
  assign \new_[6776]_  = \new_[2268]_  | \new_[2269]_ ;
  assign \new_[6777]_  = \new_[2270]_  | \new_[6776]_ ;
  assign \new_[6780]_  = \new_[2266]_  | \new_[2267]_ ;
  assign \new_[6783]_  = \new_[2264]_  | \new_[2265]_ ;
  assign \new_[6784]_  = \new_[6783]_  | \new_[6780]_ ;
  assign \new_[6785]_  = \new_[6784]_  | \new_[6777]_ ;
  assign \new_[6788]_  = \new_[2262]_  | \new_[2263]_ ;
  assign \new_[6791]_  = \new_[2260]_  | \new_[2261]_ ;
  assign \new_[6792]_  = \new_[6791]_  | \new_[6788]_ ;
  assign \new_[6795]_  = \new_[2258]_  | \new_[2259]_ ;
  assign \new_[6798]_  = \new_[2256]_  | \new_[2257]_ ;
  assign \new_[6799]_  = \new_[6798]_  | \new_[6795]_ ;
  assign \new_[6800]_  = \new_[6799]_  | \new_[6792]_ ;
  assign \new_[6801]_  = \new_[6800]_  | \new_[6785]_ ;
  assign \new_[6805]_  = \new_[2253]_  | \new_[2254]_ ;
  assign \new_[6806]_  = \new_[2255]_  | \new_[6805]_ ;
  assign \new_[6809]_  = \new_[2251]_  | \new_[2252]_ ;
  assign \new_[6812]_  = \new_[2249]_  | \new_[2250]_ ;
  assign \new_[6813]_  = \new_[6812]_  | \new_[6809]_ ;
  assign \new_[6814]_  = \new_[6813]_  | \new_[6806]_ ;
  assign \new_[6817]_  = \new_[2247]_  | \new_[2248]_ ;
  assign \new_[6820]_  = \new_[2245]_  | \new_[2246]_ ;
  assign \new_[6821]_  = \new_[6820]_  | \new_[6817]_ ;
  assign \new_[6824]_  = \new_[2243]_  | \new_[2244]_ ;
  assign \new_[6827]_  = \new_[2241]_  | \new_[2242]_ ;
  assign \new_[6828]_  = \new_[6827]_  | \new_[6824]_ ;
  assign \new_[6829]_  = \new_[6828]_  | \new_[6821]_ ;
  assign \new_[6830]_  = \new_[6829]_  | \new_[6814]_ ;
  assign \new_[6831]_  = \new_[6830]_  | \new_[6801]_ ;
  assign \new_[6832]_  = \new_[6831]_  | \new_[6772]_ ;
  assign \new_[6833]_  = \new_[6832]_  | \new_[6715]_ ;
  assign \new_[6837]_  = \new_[2238]_  | \new_[2239]_ ;
  assign \new_[6838]_  = \new_[2240]_  | \new_[6837]_ ;
  assign \new_[6841]_  = \new_[2236]_  | \new_[2237]_ ;
  assign \new_[6844]_  = \new_[2234]_  | \new_[2235]_ ;
  assign \new_[6845]_  = \new_[6844]_  | \new_[6841]_ ;
  assign \new_[6846]_  = \new_[6845]_  | \new_[6838]_ ;
  assign \new_[6850]_  = \new_[2231]_  | \new_[2232]_ ;
  assign \new_[6851]_  = \new_[2233]_  | \new_[6850]_ ;
  assign \new_[6854]_  = \new_[2229]_  | \new_[2230]_ ;
  assign \new_[6857]_  = \new_[2227]_  | \new_[2228]_ ;
  assign \new_[6858]_  = \new_[6857]_  | \new_[6854]_ ;
  assign \new_[6859]_  = \new_[6858]_  | \new_[6851]_ ;
  assign \new_[6860]_  = \new_[6859]_  | \new_[6846]_ ;
  assign \new_[6864]_  = \new_[2224]_  | \new_[2225]_ ;
  assign \new_[6865]_  = \new_[2226]_  | \new_[6864]_ ;
  assign \new_[6868]_  = \new_[2222]_  | \new_[2223]_ ;
  assign \new_[6871]_  = \new_[2220]_  | \new_[2221]_ ;
  assign \new_[6872]_  = \new_[6871]_  | \new_[6868]_ ;
  assign \new_[6873]_  = \new_[6872]_  | \new_[6865]_ ;
  assign \new_[6876]_  = \new_[2218]_  | \new_[2219]_ ;
  assign \new_[6879]_  = \new_[2216]_  | \new_[2217]_ ;
  assign \new_[6880]_  = \new_[6879]_  | \new_[6876]_ ;
  assign \new_[6883]_  = \new_[2214]_  | \new_[2215]_ ;
  assign \new_[6886]_  = \new_[2212]_  | \new_[2213]_ ;
  assign \new_[6887]_  = \new_[6886]_  | \new_[6883]_ ;
  assign \new_[6888]_  = \new_[6887]_  | \new_[6880]_ ;
  assign \new_[6889]_  = \new_[6888]_  | \new_[6873]_ ;
  assign \new_[6890]_  = \new_[6889]_  | \new_[6860]_ ;
  assign \new_[6894]_  = \new_[2209]_  | \new_[2210]_ ;
  assign \new_[6895]_  = \new_[2211]_  | \new_[6894]_ ;
  assign \new_[6898]_  = \new_[2207]_  | \new_[2208]_ ;
  assign \new_[6901]_  = \new_[2205]_  | \new_[2206]_ ;
  assign \new_[6902]_  = \new_[6901]_  | \new_[6898]_ ;
  assign \new_[6903]_  = \new_[6902]_  | \new_[6895]_ ;
  assign \new_[6906]_  = \new_[2203]_  | \new_[2204]_ ;
  assign \new_[6909]_  = \new_[2201]_  | \new_[2202]_ ;
  assign \new_[6910]_  = \new_[6909]_  | \new_[6906]_ ;
  assign \new_[6913]_  = \new_[2199]_  | \new_[2200]_ ;
  assign \new_[6916]_  = \new_[2197]_  | \new_[2198]_ ;
  assign \new_[6917]_  = \new_[6916]_  | \new_[6913]_ ;
  assign \new_[6918]_  = \new_[6917]_  | \new_[6910]_ ;
  assign \new_[6919]_  = \new_[6918]_  | \new_[6903]_ ;
  assign \new_[6923]_  = \new_[2194]_  | \new_[2195]_ ;
  assign \new_[6924]_  = \new_[2196]_  | \new_[6923]_ ;
  assign \new_[6927]_  = \new_[2192]_  | \new_[2193]_ ;
  assign \new_[6930]_  = \new_[2190]_  | \new_[2191]_ ;
  assign \new_[6931]_  = \new_[6930]_  | \new_[6927]_ ;
  assign \new_[6932]_  = \new_[6931]_  | \new_[6924]_ ;
  assign \new_[6935]_  = \new_[2188]_  | \new_[2189]_ ;
  assign \new_[6938]_  = \new_[2186]_  | \new_[2187]_ ;
  assign \new_[6939]_  = \new_[6938]_  | \new_[6935]_ ;
  assign \new_[6942]_  = \new_[2184]_  | \new_[2185]_ ;
  assign \new_[6945]_  = \new_[2182]_  | \new_[2183]_ ;
  assign \new_[6946]_  = \new_[6945]_  | \new_[6942]_ ;
  assign \new_[6947]_  = \new_[6946]_  | \new_[6939]_ ;
  assign \new_[6948]_  = \new_[6947]_  | \new_[6932]_ ;
  assign \new_[6949]_  = \new_[6948]_  | \new_[6919]_ ;
  assign \new_[6950]_  = \new_[6949]_  | \new_[6890]_ ;
  assign \new_[6954]_  = \new_[2179]_  | \new_[2180]_ ;
  assign \new_[6955]_  = \new_[2181]_  | \new_[6954]_ ;
  assign \new_[6958]_  = \new_[2177]_  | \new_[2178]_ ;
  assign \new_[6961]_  = \new_[2175]_  | \new_[2176]_ ;
  assign \new_[6962]_  = \new_[6961]_  | \new_[6958]_ ;
  assign \new_[6963]_  = \new_[6962]_  | \new_[6955]_ ;
  assign \new_[6967]_  = \new_[2172]_  | \new_[2173]_ ;
  assign \new_[6968]_  = \new_[2174]_  | \new_[6967]_ ;
  assign \new_[6971]_  = \new_[2170]_  | \new_[2171]_ ;
  assign \new_[6974]_  = \new_[2168]_  | \new_[2169]_ ;
  assign \new_[6975]_  = \new_[6974]_  | \new_[6971]_ ;
  assign \new_[6976]_  = \new_[6975]_  | \new_[6968]_ ;
  assign \new_[6977]_  = \new_[6976]_  | \new_[6963]_ ;
  assign \new_[6981]_  = \new_[2165]_  | \new_[2166]_ ;
  assign \new_[6982]_  = \new_[2167]_  | \new_[6981]_ ;
  assign \new_[6985]_  = \new_[2163]_  | \new_[2164]_ ;
  assign \new_[6988]_  = \new_[2161]_  | \new_[2162]_ ;
  assign \new_[6989]_  = \new_[6988]_  | \new_[6985]_ ;
  assign \new_[6990]_  = \new_[6989]_  | \new_[6982]_ ;
  assign \new_[6993]_  = \new_[2159]_  | \new_[2160]_ ;
  assign \new_[6996]_  = \new_[2157]_  | \new_[2158]_ ;
  assign \new_[6997]_  = \new_[6996]_  | \new_[6993]_ ;
  assign \new_[7000]_  = \new_[2155]_  | \new_[2156]_ ;
  assign \new_[7003]_  = \new_[2153]_  | \new_[2154]_ ;
  assign \new_[7004]_  = \new_[7003]_  | \new_[7000]_ ;
  assign \new_[7005]_  = \new_[7004]_  | \new_[6997]_ ;
  assign \new_[7006]_  = \new_[7005]_  | \new_[6990]_ ;
  assign \new_[7007]_  = \new_[7006]_  | \new_[6977]_ ;
  assign \new_[7011]_  = \new_[2150]_  | \new_[2151]_ ;
  assign \new_[7012]_  = \new_[2152]_  | \new_[7011]_ ;
  assign \new_[7015]_  = \new_[2148]_  | \new_[2149]_ ;
  assign \new_[7018]_  = \new_[2146]_  | \new_[2147]_ ;
  assign \new_[7019]_  = \new_[7018]_  | \new_[7015]_ ;
  assign \new_[7020]_  = \new_[7019]_  | \new_[7012]_ ;
  assign \new_[7023]_  = \new_[2144]_  | \new_[2145]_ ;
  assign \new_[7026]_  = \new_[2142]_  | \new_[2143]_ ;
  assign \new_[7027]_  = \new_[7026]_  | \new_[7023]_ ;
  assign \new_[7030]_  = \new_[2140]_  | \new_[2141]_ ;
  assign \new_[7033]_  = \new_[2138]_  | \new_[2139]_ ;
  assign \new_[7034]_  = \new_[7033]_  | \new_[7030]_ ;
  assign \new_[7035]_  = \new_[7034]_  | \new_[7027]_ ;
  assign \new_[7036]_  = \new_[7035]_  | \new_[7020]_ ;
  assign \new_[7040]_  = \new_[2135]_  | \new_[2136]_ ;
  assign \new_[7041]_  = \new_[2137]_  | \new_[7040]_ ;
  assign \new_[7044]_  = \new_[2133]_  | \new_[2134]_ ;
  assign \new_[7047]_  = \new_[2131]_  | \new_[2132]_ ;
  assign \new_[7048]_  = \new_[7047]_  | \new_[7044]_ ;
  assign \new_[7049]_  = \new_[7048]_  | \new_[7041]_ ;
  assign \new_[7052]_  = \new_[2129]_  | \new_[2130]_ ;
  assign \new_[7055]_  = \new_[2127]_  | \new_[2128]_ ;
  assign \new_[7056]_  = \new_[7055]_  | \new_[7052]_ ;
  assign \new_[7059]_  = \new_[2125]_  | \new_[2126]_ ;
  assign \new_[7062]_  = \new_[2123]_  | \new_[2124]_ ;
  assign \new_[7063]_  = \new_[7062]_  | \new_[7059]_ ;
  assign \new_[7064]_  = \new_[7063]_  | \new_[7056]_ ;
  assign \new_[7065]_  = \new_[7064]_  | \new_[7049]_ ;
  assign \new_[7066]_  = \new_[7065]_  | \new_[7036]_ ;
  assign \new_[7067]_  = \new_[7066]_  | \new_[7007]_ ;
  assign \new_[7068]_  = \new_[7067]_  | \new_[6950]_ ;
  assign \new_[7069]_  = \new_[7068]_  | \new_[6833]_ ;
  assign \new_[7073]_  = \new_[2120]_  | \new_[2121]_ ;
  assign \new_[7074]_  = \new_[2122]_  | \new_[7073]_ ;
  assign \new_[7077]_  = \new_[2118]_  | \new_[2119]_ ;
  assign \new_[7080]_  = \new_[2116]_  | \new_[2117]_ ;
  assign \new_[7081]_  = \new_[7080]_  | \new_[7077]_ ;
  assign \new_[7082]_  = \new_[7081]_  | \new_[7074]_ ;
  assign \new_[7086]_  = \new_[2113]_  | \new_[2114]_ ;
  assign \new_[7087]_  = \new_[2115]_  | \new_[7086]_ ;
  assign \new_[7090]_  = \new_[2111]_  | \new_[2112]_ ;
  assign \new_[7093]_  = \new_[2109]_  | \new_[2110]_ ;
  assign \new_[7094]_  = \new_[7093]_  | \new_[7090]_ ;
  assign \new_[7095]_  = \new_[7094]_  | \new_[7087]_ ;
  assign \new_[7096]_  = \new_[7095]_  | \new_[7082]_ ;
  assign \new_[7100]_  = \new_[2106]_  | \new_[2107]_ ;
  assign \new_[7101]_  = \new_[2108]_  | \new_[7100]_ ;
  assign \new_[7104]_  = \new_[2104]_  | \new_[2105]_ ;
  assign \new_[7107]_  = \new_[2102]_  | \new_[2103]_ ;
  assign \new_[7108]_  = \new_[7107]_  | \new_[7104]_ ;
  assign \new_[7109]_  = \new_[7108]_  | \new_[7101]_ ;
  assign \new_[7112]_  = \new_[2100]_  | \new_[2101]_ ;
  assign \new_[7115]_  = \new_[2098]_  | \new_[2099]_ ;
  assign \new_[7116]_  = \new_[7115]_  | \new_[7112]_ ;
  assign \new_[7119]_  = \new_[2096]_  | \new_[2097]_ ;
  assign \new_[7122]_  = \new_[2094]_  | \new_[2095]_ ;
  assign \new_[7123]_  = \new_[7122]_  | \new_[7119]_ ;
  assign \new_[7124]_  = \new_[7123]_  | \new_[7116]_ ;
  assign \new_[7125]_  = \new_[7124]_  | \new_[7109]_ ;
  assign \new_[7126]_  = \new_[7125]_  | \new_[7096]_ ;
  assign \new_[7130]_  = \new_[2091]_  | \new_[2092]_ ;
  assign \new_[7131]_  = \new_[2093]_  | \new_[7130]_ ;
  assign \new_[7134]_  = \new_[2089]_  | \new_[2090]_ ;
  assign \new_[7137]_  = \new_[2087]_  | \new_[2088]_ ;
  assign \new_[7138]_  = \new_[7137]_  | \new_[7134]_ ;
  assign \new_[7139]_  = \new_[7138]_  | \new_[7131]_ ;
  assign \new_[7142]_  = \new_[2085]_  | \new_[2086]_ ;
  assign \new_[7145]_  = \new_[2083]_  | \new_[2084]_ ;
  assign \new_[7146]_  = \new_[7145]_  | \new_[7142]_ ;
  assign \new_[7149]_  = \new_[2081]_  | \new_[2082]_ ;
  assign \new_[7152]_  = \new_[2079]_  | \new_[2080]_ ;
  assign \new_[7153]_  = \new_[7152]_  | \new_[7149]_ ;
  assign \new_[7154]_  = \new_[7153]_  | \new_[7146]_ ;
  assign \new_[7155]_  = \new_[7154]_  | \new_[7139]_ ;
  assign \new_[7159]_  = \new_[2076]_  | \new_[2077]_ ;
  assign \new_[7160]_  = \new_[2078]_  | \new_[7159]_ ;
  assign \new_[7163]_  = \new_[2074]_  | \new_[2075]_ ;
  assign \new_[7166]_  = \new_[2072]_  | \new_[2073]_ ;
  assign \new_[7167]_  = \new_[7166]_  | \new_[7163]_ ;
  assign \new_[7168]_  = \new_[7167]_  | \new_[7160]_ ;
  assign \new_[7171]_  = \new_[2070]_  | \new_[2071]_ ;
  assign \new_[7174]_  = \new_[2068]_  | \new_[2069]_ ;
  assign \new_[7175]_  = \new_[7174]_  | \new_[7171]_ ;
  assign \new_[7178]_  = \new_[2066]_  | \new_[2067]_ ;
  assign \new_[7181]_  = \new_[2064]_  | \new_[2065]_ ;
  assign \new_[7182]_  = \new_[7181]_  | \new_[7178]_ ;
  assign \new_[7183]_  = \new_[7182]_  | \new_[7175]_ ;
  assign \new_[7184]_  = \new_[7183]_  | \new_[7168]_ ;
  assign \new_[7185]_  = \new_[7184]_  | \new_[7155]_ ;
  assign \new_[7186]_  = \new_[7185]_  | \new_[7126]_ ;
  assign \new_[7190]_  = \new_[2061]_  | \new_[2062]_ ;
  assign \new_[7191]_  = \new_[2063]_  | \new_[7190]_ ;
  assign \new_[7194]_  = \new_[2059]_  | \new_[2060]_ ;
  assign \new_[7197]_  = \new_[2057]_  | \new_[2058]_ ;
  assign \new_[7198]_  = \new_[7197]_  | \new_[7194]_ ;
  assign \new_[7199]_  = \new_[7198]_  | \new_[7191]_ ;
  assign \new_[7203]_  = \new_[2054]_  | \new_[2055]_ ;
  assign \new_[7204]_  = \new_[2056]_  | \new_[7203]_ ;
  assign \new_[7207]_  = \new_[2052]_  | \new_[2053]_ ;
  assign \new_[7210]_  = \new_[2050]_  | \new_[2051]_ ;
  assign \new_[7211]_  = \new_[7210]_  | \new_[7207]_ ;
  assign \new_[7212]_  = \new_[7211]_  | \new_[7204]_ ;
  assign \new_[7213]_  = \new_[7212]_  | \new_[7199]_ ;
  assign \new_[7217]_  = \new_[2047]_  | \new_[2048]_ ;
  assign \new_[7218]_  = \new_[2049]_  | \new_[7217]_ ;
  assign \new_[7221]_  = \new_[2045]_  | \new_[2046]_ ;
  assign \new_[7224]_  = \new_[2043]_  | \new_[2044]_ ;
  assign \new_[7225]_  = \new_[7224]_  | \new_[7221]_ ;
  assign \new_[7226]_  = \new_[7225]_  | \new_[7218]_ ;
  assign \new_[7229]_  = \new_[2041]_  | \new_[2042]_ ;
  assign \new_[7232]_  = \new_[2039]_  | \new_[2040]_ ;
  assign \new_[7233]_  = \new_[7232]_  | \new_[7229]_ ;
  assign \new_[7236]_  = \new_[2037]_  | \new_[2038]_ ;
  assign \new_[7239]_  = \new_[2035]_  | \new_[2036]_ ;
  assign \new_[7240]_  = \new_[7239]_  | \new_[7236]_ ;
  assign \new_[7241]_  = \new_[7240]_  | \new_[7233]_ ;
  assign \new_[7242]_  = \new_[7241]_  | \new_[7226]_ ;
  assign \new_[7243]_  = \new_[7242]_  | \new_[7213]_ ;
  assign \new_[7247]_  = \new_[2032]_  | \new_[2033]_ ;
  assign \new_[7248]_  = \new_[2034]_  | \new_[7247]_ ;
  assign \new_[7251]_  = \new_[2030]_  | \new_[2031]_ ;
  assign \new_[7254]_  = \new_[2028]_  | \new_[2029]_ ;
  assign \new_[7255]_  = \new_[7254]_  | \new_[7251]_ ;
  assign \new_[7256]_  = \new_[7255]_  | \new_[7248]_ ;
  assign \new_[7259]_  = \new_[2026]_  | \new_[2027]_ ;
  assign \new_[7262]_  = \new_[2024]_  | \new_[2025]_ ;
  assign \new_[7263]_  = \new_[7262]_  | \new_[7259]_ ;
  assign \new_[7266]_  = \new_[2022]_  | \new_[2023]_ ;
  assign \new_[7269]_  = \new_[2020]_  | \new_[2021]_ ;
  assign \new_[7270]_  = \new_[7269]_  | \new_[7266]_ ;
  assign \new_[7271]_  = \new_[7270]_  | \new_[7263]_ ;
  assign \new_[7272]_  = \new_[7271]_  | \new_[7256]_ ;
  assign \new_[7276]_  = \new_[2017]_  | \new_[2018]_ ;
  assign \new_[7277]_  = \new_[2019]_  | \new_[7276]_ ;
  assign \new_[7280]_  = \new_[2015]_  | \new_[2016]_ ;
  assign \new_[7283]_  = \new_[2013]_  | \new_[2014]_ ;
  assign \new_[7284]_  = \new_[7283]_  | \new_[7280]_ ;
  assign \new_[7285]_  = \new_[7284]_  | \new_[7277]_ ;
  assign \new_[7288]_  = \new_[2011]_  | \new_[2012]_ ;
  assign \new_[7291]_  = \new_[2009]_  | \new_[2010]_ ;
  assign \new_[7292]_  = \new_[7291]_  | \new_[7288]_ ;
  assign \new_[7295]_  = \new_[2007]_  | \new_[2008]_ ;
  assign \new_[7298]_  = \new_[2005]_  | \new_[2006]_ ;
  assign \new_[7299]_  = \new_[7298]_  | \new_[7295]_ ;
  assign \new_[7300]_  = \new_[7299]_  | \new_[7292]_ ;
  assign \new_[7301]_  = \new_[7300]_  | \new_[7285]_ ;
  assign \new_[7302]_  = \new_[7301]_  | \new_[7272]_ ;
  assign \new_[7303]_  = \new_[7302]_  | \new_[7243]_ ;
  assign \new_[7304]_  = \new_[7303]_  | \new_[7186]_ ;
  assign \new_[7308]_  = \new_[2002]_  | \new_[2003]_ ;
  assign \new_[7309]_  = \new_[2004]_  | \new_[7308]_ ;
  assign \new_[7312]_  = \new_[2000]_  | \new_[2001]_ ;
  assign \new_[7315]_  = \new_[1998]_  | \new_[1999]_ ;
  assign \new_[7316]_  = \new_[7315]_  | \new_[7312]_ ;
  assign \new_[7317]_  = \new_[7316]_  | \new_[7309]_ ;
  assign \new_[7321]_  = \new_[1995]_  | \new_[1996]_ ;
  assign \new_[7322]_  = \new_[1997]_  | \new_[7321]_ ;
  assign \new_[7325]_  = \new_[1993]_  | \new_[1994]_ ;
  assign \new_[7328]_  = \new_[1991]_  | \new_[1992]_ ;
  assign \new_[7329]_  = \new_[7328]_  | \new_[7325]_ ;
  assign \new_[7330]_  = \new_[7329]_  | \new_[7322]_ ;
  assign \new_[7331]_  = \new_[7330]_  | \new_[7317]_ ;
  assign \new_[7335]_  = \new_[1988]_  | \new_[1989]_ ;
  assign \new_[7336]_  = \new_[1990]_  | \new_[7335]_ ;
  assign \new_[7339]_  = \new_[1986]_  | \new_[1987]_ ;
  assign \new_[7342]_  = \new_[1984]_  | \new_[1985]_ ;
  assign \new_[7343]_  = \new_[7342]_  | \new_[7339]_ ;
  assign \new_[7344]_  = \new_[7343]_  | \new_[7336]_ ;
  assign \new_[7347]_  = \new_[1982]_  | \new_[1983]_ ;
  assign \new_[7350]_  = \new_[1980]_  | \new_[1981]_ ;
  assign \new_[7351]_  = \new_[7350]_  | \new_[7347]_ ;
  assign \new_[7354]_  = \new_[1978]_  | \new_[1979]_ ;
  assign \new_[7357]_  = \new_[1976]_  | \new_[1977]_ ;
  assign \new_[7358]_  = \new_[7357]_  | \new_[7354]_ ;
  assign \new_[7359]_  = \new_[7358]_  | \new_[7351]_ ;
  assign \new_[7360]_  = \new_[7359]_  | \new_[7344]_ ;
  assign \new_[7361]_  = \new_[7360]_  | \new_[7331]_ ;
  assign \new_[7365]_  = \new_[1973]_  | \new_[1974]_ ;
  assign \new_[7366]_  = \new_[1975]_  | \new_[7365]_ ;
  assign \new_[7369]_  = \new_[1971]_  | \new_[1972]_ ;
  assign \new_[7372]_  = \new_[1969]_  | \new_[1970]_ ;
  assign \new_[7373]_  = \new_[7372]_  | \new_[7369]_ ;
  assign \new_[7374]_  = \new_[7373]_  | \new_[7366]_ ;
  assign \new_[7377]_  = \new_[1967]_  | \new_[1968]_ ;
  assign \new_[7380]_  = \new_[1965]_  | \new_[1966]_ ;
  assign \new_[7381]_  = \new_[7380]_  | \new_[7377]_ ;
  assign \new_[7384]_  = \new_[1963]_  | \new_[1964]_ ;
  assign \new_[7387]_  = \new_[1961]_  | \new_[1962]_ ;
  assign \new_[7388]_  = \new_[7387]_  | \new_[7384]_ ;
  assign \new_[7389]_  = \new_[7388]_  | \new_[7381]_ ;
  assign \new_[7390]_  = \new_[7389]_  | \new_[7374]_ ;
  assign \new_[7394]_  = \new_[1958]_  | \new_[1959]_ ;
  assign \new_[7395]_  = \new_[1960]_  | \new_[7394]_ ;
  assign \new_[7398]_  = \new_[1956]_  | \new_[1957]_ ;
  assign \new_[7401]_  = \new_[1954]_  | \new_[1955]_ ;
  assign \new_[7402]_  = \new_[7401]_  | \new_[7398]_ ;
  assign \new_[7403]_  = \new_[7402]_  | \new_[7395]_ ;
  assign \new_[7406]_  = \new_[1952]_  | \new_[1953]_ ;
  assign \new_[7409]_  = \new_[1950]_  | \new_[1951]_ ;
  assign \new_[7410]_  = \new_[7409]_  | \new_[7406]_ ;
  assign \new_[7413]_  = \new_[1948]_  | \new_[1949]_ ;
  assign \new_[7416]_  = \new_[1946]_  | \new_[1947]_ ;
  assign \new_[7417]_  = \new_[7416]_  | \new_[7413]_ ;
  assign \new_[7418]_  = \new_[7417]_  | \new_[7410]_ ;
  assign \new_[7419]_  = \new_[7418]_  | \new_[7403]_ ;
  assign \new_[7420]_  = \new_[7419]_  | \new_[7390]_ ;
  assign \new_[7421]_  = \new_[7420]_  | \new_[7361]_ ;
  assign \new_[7425]_  = \new_[1943]_  | \new_[1944]_ ;
  assign \new_[7426]_  = \new_[1945]_  | \new_[7425]_ ;
  assign \new_[7429]_  = \new_[1941]_  | \new_[1942]_ ;
  assign \new_[7432]_  = \new_[1939]_  | \new_[1940]_ ;
  assign \new_[7433]_  = \new_[7432]_  | \new_[7429]_ ;
  assign \new_[7434]_  = \new_[7433]_  | \new_[7426]_ ;
  assign \new_[7438]_  = \new_[1936]_  | \new_[1937]_ ;
  assign \new_[7439]_  = \new_[1938]_  | \new_[7438]_ ;
  assign \new_[7442]_  = \new_[1934]_  | \new_[1935]_ ;
  assign \new_[7445]_  = \new_[1932]_  | \new_[1933]_ ;
  assign \new_[7446]_  = \new_[7445]_  | \new_[7442]_ ;
  assign \new_[7447]_  = \new_[7446]_  | \new_[7439]_ ;
  assign \new_[7448]_  = \new_[7447]_  | \new_[7434]_ ;
  assign \new_[7452]_  = \new_[1929]_  | \new_[1930]_ ;
  assign \new_[7453]_  = \new_[1931]_  | \new_[7452]_ ;
  assign \new_[7456]_  = \new_[1927]_  | \new_[1928]_ ;
  assign \new_[7459]_  = \new_[1925]_  | \new_[1926]_ ;
  assign \new_[7460]_  = \new_[7459]_  | \new_[7456]_ ;
  assign \new_[7461]_  = \new_[7460]_  | \new_[7453]_ ;
  assign \new_[7464]_  = \new_[1923]_  | \new_[1924]_ ;
  assign \new_[7467]_  = \new_[1921]_  | \new_[1922]_ ;
  assign \new_[7468]_  = \new_[7467]_  | \new_[7464]_ ;
  assign \new_[7471]_  = \new_[1919]_  | \new_[1920]_ ;
  assign \new_[7474]_  = \new_[1917]_  | \new_[1918]_ ;
  assign \new_[7475]_  = \new_[7474]_  | \new_[7471]_ ;
  assign \new_[7476]_  = \new_[7475]_  | \new_[7468]_ ;
  assign \new_[7477]_  = \new_[7476]_  | \new_[7461]_ ;
  assign \new_[7478]_  = \new_[7477]_  | \new_[7448]_ ;
  assign \new_[7482]_  = \new_[1914]_  | \new_[1915]_ ;
  assign \new_[7483]_  = \new_[1916]_  | \new_[7482]_ ;
  assign \new_[7486]_  = \new_[1912]_  | \new_[1913]_ ;
  assign \new_[7489]_  = \new_[1910]_  | \new_[1911]_ ;
  assign \new_[7490]_  = \new_[7489]_  | \new_[7486]_ ;
  assign \new_[7491]_  = \new_[7490]_  | \new_[7483]_ ;
  assign \new_[7494]_  = \new_[1908]_  | \new_[1909]_ ;
  assign \new_[7497]_  = \new_[1906]_  | \new_[1907]_ ;
  assign \new_[7498]_  = \new_[7497]_  | \new_[7494]_ ;
  assign \new_[7501]_  = \new_[1904]_  | \new_[1905]_ ;
  assign \new_[7504]_  = \new_[1902]_  | \new_[1903]_ ;
  assign \new_[7505]_  = \new_[7504]_  | \new_[7501]_ ;
  assign \new_[7506]_  = \new_[7505]_  | \new_[7498]_ ;
  assign \new_[7507]_  = \new_[7506]_  | \new_[7491]_ ;
  assign \new_[7511]_  = \new_[1899]_  | \new_[1900]_ ;
  assign \new_[7512]_  = \new_[1901]_  | \new_[7511]_ ;
  assign \new_[7515]_  = \new_[1897]_  | \new_[1898]_ ;
  assign \new_[7518]_  = \new_[1895]_  | \new_[1896]_ ;
  assign \new_[7519]_  = \new_[7518]_  | \new_[7515]_ ;
  assign \new_[7520]_  = \new_[7519]_  | \new_[7512]_ ;
  assign \new_[7523]_  = \new_[1893]_  | \new_[1894]_ ;
  assign \new_[7526]_  = \new_[1891]_  | \new_[1892]_ ;
  assign \new_[7527]_  = \new_[7526]_  | \new_[7523]_ ;
  assign \new_[7530]_  = \new_[1889]_  | \new_[1890]_ ;
  assign \new_[7533]_  = \new_[1887]_  | \new_[1888]_ ;
  assign \new_[7534]_  = \new_[7533]_  | \new_[7530]_ ;
  assign \new_[7535]_  = \new_[7534]_  | \new_[7527]_ ;
  assign \new_[7536]_  = \new_[7535]_  | \new_[7520]_ ;
  assign \new_[7537]_  = \new_[7536]_  | \new_[7507]_ ;
  assign \new_[7538]_  = \new_[7537]_  | \new_[7478]_ ;
  assign \new_[7539]_  = \new_[7538]_  | \new_[7421]_ ;
  assign \new_[7540]_  = \new_[7539]_  | \new_[7304]_ ;
  assign \new_[7541]_  = \new_[7540]_  | \new_[7069]_ ;
  assign \new_[7542]_  = \new_[7541]_  | \new_[6598]_ ;
  assign \new_[7543]_  = \new_[7542]_  | \new_[5657]_ ;
  assign \new_[7547]_  = \new_[1884]_  | \new_[1885]_ ;
  assign \new_[7548]_  = \new_[1886]_  | \new_[7547]_ ;
  assign \new_[7551]_  = \new_[1882]_  | \new_[1883]_ ;
  assign \new_[7554]_  = \new_[1880]_  | \new_[1881]_ ;
  assign \new_[7555]_  = \new_[7554]_  | \new_[7551]_ ;
  assign \new_[7556]_  = \new_[7555]_  | \new_[7548]_ ;
  assign \new_[7560]_  = \new_[1877]_  | \new_[1878]_ ;
  assign \new_[7561]_  = \new_[1879]_  | \new_[7560]_ ;
  assign \new_[7564]_  = \new_[1875]_  | \new_[1876]_ ;
  assign \new_[7567]_  = \new_[1873]_  | \new_[1874]_ ;
  assign \new_[7568]_  = \new_[7567]_  | \new_[7564]_ ;
  assign \new_[7569]_  = \new_[7568]_  | \new_[7561]_ ;
  assign \new_[7570]_  = \new_[7569]_  | \new_[7556]_ ;
  assign \new_[7574]_  = \new_[1870]_  | \new_[1871]_ ;
  assign \new_[7575]_  = \new_[1872]_  | \new_[7574]_ ;
  assign \new_[7578]_  = \new_[1868]_  | \new_[1869]_ ;
  assign \new_[7581]_  = \new_[1866]_  | \new_[1867]_ ;
  assign \new_[7582]_  = \new_[7581]_  | \new_[7578]_ ;
  assign \new_[7583]_  = \new_[7582]_  | \new_[7575]_ ;
  assign \new_[7586]_  = \new_[1864]_  | \new_[1865]_ ;
  assign \new_[7589]_  = \new_[1862]_  | \new_[1863]_ ;
  assign \new_[7590]_  = \new_[7589]_  | \new_[7586]_ ;
  assign \new_[7593]_  = \new_[1860]_  | \new_[1861]_ ;
  assign \new_[7596]_  = \new_[1858]_  | \new_[1859]_ ;
  assign \new_[7597]_  = \new_[7596]_  | \new_[7593]_ ;
  assign \new_[7598]_  = \new_[7597]_  | \new_[7590]_ ;
  assign \new_[7599]_  = \new_[7598]_  | \new_[7583]_ ;
  assign \new_[7600]_  = \new_[7599]_  | \new_[7570]_ ;
  assign \new_[7604]_  = \new_[1855]_  | \new_[1856]_ ;
  assign \new_[7605]_  = \new_[1857]_  | \new_[7604]_ ;
  assign \new_[7608]_  = \new_[1853]_  | \new_[1854]_ ;
  assign \new_[7611]_  = \new_[1851]_  | \new_[1852]_ ;
  assign \new_[7612]_  = \new_[7611]_  | \new_[7608]_ ;
  assign \new_[7613]_  = \new_[7612]_  | \new_[7605]_ ;
  assign \new_[7617]_  = \new_[1848]_  | \new_[1849]_ ;
  assign \new_[7618]_  = \new_[1850]_  | \new_[7617]_ ;
  assign \new_[7621]_  = \new_[1846]_  | \new_[1847]_ ;
  assign \new_[7624]_  = \new_[1844]_  | \new_[1845]_ ;
  assign \new_[7625]_  = \new_[7624]_  | \new_[7621]_ ;
  assign \new_[7626]_  = \new_[7625]_  | \new_[7618]_ ;
  assign \new_[7627]_  = \new_[7626]_  | \new_[7613]_ ;
  assign \new_[7631]_  = \new_[1841]_  | \new_[1842]_ ;
  assign \new_[7632]_  = \new_[1843]_  | \new_[7631]_ ;
  assign \new_[7635]_  = \new_[1839]_  | \new_[1840]_ ;
  assign \new_[7638]_  = \new_[1837]_  | \new_[1838]_ ;
  assign \new_[7639]_  = \new_[7638]_  | \new_[7635]_ ;
  assign \new_[7640]_  = \new_[7639]_  | \new_[7632]_ ;
  assign \new_[7643]_  = \new_[1835]_  | \new_[1836]_ ;
  assign \new_[7646]_  = \new_[1833]_  | \new_[1834]_ ;
  assign \new_[7647]_  = \new_[7646]_  | \new_[7643]_ ;
  assign \new_[7650]_  = \new_[1831]_  | \new_[1832]_ ;
  assign \new_[7653]_  = \new_[1829]_  | \new_[1830]_ ;
  assign \new_[7654]_  = \new_[7653]_  | \new_[7650]_ ;
  assign \new_[7655]_  = \new_[7654]_  | \new_[7647]_ ;
  assign \new_[7656]_  = \new_[7655]_  | \new_[7640]_ ;
  assign \new_[7657]_  = \new_[7656]_  | \new_[7627]_ ;
  assign \new_[7658]_  = \new_[7657]_  | \new_[7600]_ ;
  assign \new_[7662]_  = \new_[1826]_  | \new_[1827]_ ;
  assign \new_[7663]_  = \new_[1828]_  | \new_[7662]_ ;
  assign \new_[7666]_  = \new_[1824]_  | \new_[1825]_ ;
  assign \new_[7669]_  = \new_[1822]_  | \new_[1823]_ ;
  assign \new_[7670]_  = \new_[7669]_  | \new_[7666]_ ;
  assign \new_[7671]_  = \new_[7670]_  | \new_[7663]_ ;
  assign \new_[7675]_  = \new_[1819]_  | \new_[1820]_ ;
  assign \new_[7676]_  = \new_[1821]_  | \new_[7675]_ ;
  assign \new_[7679]_  = \new_[1817]_  | \new_[1818]_ ;
  assign \new_[7682]_  = \new_[1815]_  | \new_[1816]_ ;
  assign \new_[7683]_  = \new_[7682]_  | \new_[7679]_ ;
  assign \new_[7684]_  = \new_[7683]_  | \new_[7676]_ ;
  assign \new_[7685]_  = \new_[7684]_  | \new_[7671]_ ;
  assign \new_[7689]_  = \new_[1812]_  | \new_[1813]_ ;
  assign \new_[7690]_  = \new_[1814]_  | \new_[7689]_ ;
  assign \new_[7693]_  = \new_[1810]_  | \new_[1811]_ ;
  assign \new_[7696]_  = \new_[1808]_  | \new_[1809]_ ;
  assign \new_[7697]_  = \new_[7696]_  | \new_[7693]_ ;
  assign \new_[7698]_  = \new_[7697]_  | \new_[7690]_ ;
  assign \new_[7701]_  = \new_[1806]_  | \new_[1807]_ ;
  assign \new_[7704]_  = \new_[1804]_  | \new_[1805]_ ;
  assign \new_[7705]_  = \new_[7704]_  | \new_[7701]_ ;
  assign \new_[7708]_  = \new_[1802]_  | \new_[1803]_ ;
  assign \new_[7711]_  = \new_[1800]_  | \new_[1801]_ ;
  assign \new_[7712]_  = \new_[7711]_  | \new_[7708]_ ;
  assign \new_[7713]_  = \new_[7712]_  | \new_[7705]_ ;
  assign \new_[7714]_  = \new_[7713]_  | \new_[7698]_ ;
  assign \new_[7715]_  = \new_[7714]_  | \new_[7685]_ ;
  assign \new_[7719]_  = \new_[1797]_  | \new_[1798]_ ;
  assign \new_[7720]_  = \new_[1799]_  | \new_[7719]_ ;
  assign \new_[7723]_  = \new_[1795]_  | \new_[1796]_ ;
  assign \new_[7726]_  = \new_[1793]_  | \new_[1794]_ ;
  assign \new_[7727]_  = \new_[7726]_  | \new_[7723]_ ;
  assign \new_[7728]_  = \new_[7727]_  | \new_[7720]_ ;
  assign \new_[7731]_  = \new_[1791]_  | \new_[1792]_ ;
  assign \new_[7734]_  = \new_[1789]_  | \new_[1790]_ ;
  assign \new_[7735]_  = \new_[7734]_  | \new_[7731]_ ;
  assign \new_[7738]_  = \new_[1787]_  | \new_[1788]_ ;
  assign \new_[7741]_  = \new_[1785]_  | \new_[1786]_ ;
  assign \new_[7742]_  = \new_[7741]_  | \new_[7738]_ ;
  assign \new_[7743]_  = \new_[7742]_  | \new_[7735]_ ;
  assign \new_[7744]_  = \new_[7743]_  | \new_[7728]_ ;
  assign \new_[7748]_  = \new_[1782]_  | \new_[1783]_ ;
  assign \new_[7749]_  = \new_[1784]_  | \new_[7748]_ ;
  assign \new_[7752]_  = \new_[1780]_  | \new_[1781]_ ;
  assign \new_[7755]_  = \new_[1778]_  | \new_[1779]_ ;
  assign \new_[7756]_  = \new_[7755]_  | \new_[7752]_ ;
  assign \new_[7757]_  = \new_[7756]_  | \new_[7749]_ ;
  assign \new_[7760]_  = \new_[1776]_  | \new_[1777]_ ;
  assign \new_[7763]_  = \new_[1774]_  | \new_[1775]_ ;
  assign \new_[7764]_  = \new_[7763]_  | \new_[7760]_ ;
  assign \new_[7767]_  = \new_[1772]_  | \new_[1773]_ ;
  assign \new_[7770]_  = \new_[1770]_  | \new_[1771]_ ;
  assign \new_[7771]_  = \new_[7770]_  | \new_[7767]_ ;
  assign \new_[7772]_  = \new_[7771]_  | \new_[7764]_ ;
  assign \new_[7773]_  = \new_[7772]_  | \new_[7757]_ ;
  assign \new_[7774]_  = \new_[7773]_  | \new_[7744]_ ;
  assign \new_[7775]_  = \new_[7774]_  | \new_[7715]_ ;
  assign \new_[7776]_  = \new_[7775]_  | \new_[7658]_ ;
  assign \new_[7780]_  = \new_[1767]_  | \new_[1768]_ ;
  assign \new_[7781]_  = \new_[1769]_  | \new_[7780]_ ;
  assign \new_[7784]_  = \new_[1765]_  | \new_[1766]_ ;
  assign \new_[7787]_  = \new_[1763]_  | \new_[1764]_ ;
  assign \new_[7788]_  = \new_[7787]_  | \new_[7784]_ ;
  assign \new_[7789]_  = \new_[7788]_  | \new_[7781]_ ;
  assign \new_[7793]_  = \new_[1760]_  | \new_[1761]_ ;
  assign \new_[7794]_  = \new_[1762]_  | \new_[7793]_ ;
  assign \new_[7797]_  = \new_[1758]_  | \new_[1759]_ ;
  assign \new_[7800]_  = \new_[1756]_  | \new_[1757]_ ;
  assign \new_[7801]_  = \new_[7800]_  | \new_[7797]_ ;
  assign \new_[7802]_  = \new_[7801]_  | \new_[7794]_ ;
  assign \new_[7803]_  = \new_[7802]_  | \new_[7789]_ ;
  assign \new_[7807]_  = \new_[1753]_  | \new_[1754]_ ;
  assign \new_[7808]_  = \new_[1755]_  | \new_[7807]_ ;
  assign \new_[7811]_  = \new_[1751]_  | \new_[1752]_ ;
  assign \new_[7814]_  = \new_[1749]_  | \new_[1750]_ ;
  assign \new_[7815]_  = \new_[7814]_  | \new_[7811]_ ;
  assign \new_[7816]_  = \new_[7815]_  | \new_[7808]_ ;
  assign \new_[7819]_  = \new_[1747]_  | \new_[1748]_ ;
  assign \new_[7822]_  = \new_[1745]_  | \new_[1746]_ ;
  assign \new_[7823]_  = \new_[7822]_  | \new_[7819]_ ;
  assign \new_[7826]_  = \new_[1743]_  | \new_[1744]_ ;
  assign \new_[7829]_  = \new_[1741]_  | \new_[1742]_ ;
  assign \new_[7830]_  = \new_[7829]_  | \new_[7826]_ ;
  assign \new_[7831]_  = \new_[7830]_  | \new_[7823]_ ;
  assign \new_[7832]_  = \new_[7831]_  | \new_[7816]_ ;
  assign \new_[7833]_  = \new_[7832]_  | \new_[7803]_ ;
  assign \new_[7837]_  = \new_[1738]_  | \new_[1739]_ ;
  assign \new_[7838]_  = \new_[1740]_  | \new_[7837]_ ;
  assign \new_[7841]_  = \new_[1736]_  | \new_[1737]_ ;
  assign \new_[7844]_  = \new_[1734]_  | \new_[1735]_ ;
  assign \new_[7845]_  = \new_[7844]_  | \new_[7841]_ ;
  assign \new_[7846]_  = \new_[7845]_  | \new_[7838]_ ;
  assign \new_[7849]_  = \new_[1732]_  | \new_[1733]_ ;
  assign \new_[7852]_  = \new_[1730]_  | \new_[1731]_ ;
  assign \new_[7853]_  = \new_[7852]_  | \new_[7849]_ ;
  assign \new_[7856]_  = \new_[1728]_  | \new_[1729]_ ;
  assign \new_[7859]_  = \new_[1726]_  | \new_[1727]_ ;
  assign \new_[7860]_  = \new_[7859]_  | \new_[7856]_ ;
  assign \new_[7861]_  = \new_[7860]_  | \new_[7853]_ ;
  assign \new_[7862]_  = \new_[7861]_  | \new_[7846]_ ;
  assign \new_[7866]_  = \new_[1723]_  | \new_[1724]_ ;
  assign \new_[7867]_  = \new_[1725]_  | \new_[7866]_ ;
  assign \new_[7870]_  = \new_[1721]_  | \new_[1722]_ ;
  assign \new_[7873]_  = \new_[1719]_  | \new_[1720]_ ;
  assign \new_[7874]_  = \new_[7873]_  | \new_[7870]_ ;
  assign \new_[7875]_  = \new_[7874]_  | \new_[7867]_ ;
  assign \new_[7878]_  = \new_[1717]_  | \new_[1718]_ ;
  assign \new_[7881]_  = \new_[1715]_  | \new_[1716]_ ;
  assign \new_[7882]_  = \new_[7881]_  | \new_[7878]_ ;
  assign \new_[7885]_  = \new_[1713]_  | \new_[1714]_ ;
  assign \new_[7888]_  = \new_[1711]_  | \new_[1712]_ ;
  assign \new_[7889]_  = \new_[7888]_  | \new_[7885]_ ;
  assign \new_[7890]_  = \new_[7889]_  | \new_[7882]_ ;
  assign \new_[7891]_  = \new_[7890]_  | \new_[7875]_ ;
  assign \new_[7892]_  = \new_[7891]_  | \new_[7862]_ ;
  assign \new_[7893]_  = \new_[7892]_  | \new_[7833]_ ;
  assign \new_[7897]_  = \new_[1708]_  | \new_[1709]_ ;
  assign \new_[7898]_  = \new_[1710]_  | \new_[7897]_ ;
  assign \new_[7901]_  = \new_[1706]_  | \new_[1707]_ ;
  assign \new_[7904]_  = \new_[1704]_  | \new_[1705]_ ;
  assign \new_[7905]_  = \new_[7904]_  | \new_[7901]_ ;
  assign \new_[7906]_  = \new_[7905]_  | \new_[7898]_ ;
  assign \new_[7910]_  = \new_[1701]_  | \new_[1702]_ ;
  assign \new_[7911]_  = \new_[1703]_  | \new_[7910]_ ;
  assign \new_[7914]_  = \new_[1699]_  | \new_[1700]_ ;
  assign \new_[7917]_  = \new_[1697]_  | \new_[1698]_ ;
  assign \new_[7918]_  = \new_[7917]_  | \new_[7914]_ ;
  assign \new_[7919]_  = \new_[7918]_  | \new_[7911]_ ;
  assign \new_[7920]_  = \new_[7919]_  | \new_[7906]_ ;
  assign \new_[7924]_  = \new_[1694]_  | \new_[1695]_ ;
  assign \new_[7925]_  = \new_[1696]_  | \new_[7924]_ ;
  assign \new_[7928]_  = \new_[1692]_  | \new_[1693]_ ;
  assign \new_[7931]_  = \new_[1690]_  | \new_[1691]_ ;
  assign \new_[7932]_  = \new_[7931]_  | \new_[7928]_ ;
  assign \new_[7933]_  = \new_[7932]_  | \new_[7925]_ ;
  assign \new_[7936]_  = \new_[1688]_  | \new_[1689]_ ;
  assign \new_[7939]_  = \new_[1686]_  | \new_[1687]_ ;
  assign \new_[7940]_  = \new_[7939]_  | \new_[7936]_ ;
  assign \new_[7943]_  = \new_[1684]_  | \new_[1685]_ ;
  assign \new_[7946]_  = \new_[1682]_  | \new_[1683]_ ;
  assign \new_[7947]_  = \new_[7946]_  | \new_[7943]_ ;
  assign \new_[7948]_  = \new_[7947]_  | \new_[7940]_ ;
  assign \new_[7949]_  = \new_[7948]_  | \new_[7933]_ ;
  assign \new_[7950]_  = \new_[7949]_  | \new_[7920]_ ;
  assign \new_[7954]_  = \new_[1679]_  | \new_[1680]_ ;
  assign \new_[7955]_  = \new_[1681]_  | \new_[7954]_ ;
  assign \new_[7958]_  = \new_[1677]_  | \new_[1678]_ ;
  assign \new_[7961]_  = \new_[1675]_  | \new_[1676]_ ;
  assign \new_[7962]_  = \new_[7961]_  | \new_[7958]_ ;
  assign \new_[7963]_  = \new_[7962]_  | \new_[7955]_ ;
  assign \new_[7966]_  = \new_[1673]_  | \new_[1674]_ ;
  assign \new_[7969]_  = \new_[1671]_  | \new_[1672]_ ;
  assign \new_[7970]_  = \new_[7969]_  | \new_[7966]_ ;
  assign \new_[7973]_  = \new_[1669]_  | \new_[1670]_ ;
  assign \new_[7976]_  = \new_[1667]_  | \new_[1668]_ ;
  assign \new_[7977]_  = \new_[7976]_  | \new_[7973]_ ;
  assign \new_[7978]_  = \new_[7977]_  | \new_[7970]_ ;
  assign \new_[7979]_  = \new_[7978]_  | \new_[7963]_ ;
  assign \new_[7983]_  = \new_[1664]_  | \new_[1665]_ ;
  assign \new_[7984]_  = \new_[1666]_  | \new_[7983]_ ;
  assign \new_[7987]_  = \new_[1662]_  | \new_[1663]_ ;
  assign \new_[7990]_  = \new_[1660]_  | \new_[1661]_ ;
  assign \new_[7991]_  = \new_[7990]_  | \new_[7987]_ ;
  assign \new_[7992]_  = \new_[7991]_  | \new_[7984]_ ;
  assign \new_[7995]_  = \new_[1658]_  | \new_[1659]_ ;
  assign \new_[7998]_  = \new_[1656]_  | \new_[1657]_ ;
  assign \new_[7999]_  = \new_[7998]_  | \new_[7995]_ ;
  assign \new_[8002]_  = \new_[1654]_  | \new_[1655]_ ;
  assign \new_[8005]_  = \new_[1652]_  | \new_[1653]_ ;
  assign \new_[8006]_  = \new_[8005]_  | \new_[8002]_ ;
  assign \new_[8007]_  = \new_[8006]_  | \new_[7999]_ ;
  assign \new_[8008]_  = \new_[8007]_  | \new_[7992]_ ;
  assign \new_[8009]_  = \new_[8008]_  | \new_[7979]_ ;
  assign \new_[8010]_  = \new_[8009]_  | \new_[7950]_ ;
  assign \new_[8011]_  = \new_[8010]_  | \new_[7893]_ ;
  assign \new_[8012]_  = \new_[8011]_  | \new_[7776]_ ;
  assign \new_[8016]_  = \new_[1649]_  | \new_[1650]_ ;
  assign \new_[8017]_  = \new_[1651]_  | \new_[8016]_ ;
  assign \new_[8020]_  = \new_[1647]_  | \new_[1648]_ ;
  assign \new_[8023]_  = \new_[1645]_  | \new_[1646]_ ;
  assign \new_[8024]_  = \new_[8023]_  | \new_[8020]_ ;
  assign \new_[8025]_  = \new_[8024]_  | \new_[8017]_ ;
  assign \new_[8029]_  = \new_[1642]_  | \new_[1643]_ ;
  assign \new_[8030]_  = \new_[1644]_  | \new_[8029]_ ;
  assign \new_[8033]_  = \new_[1640]_  | \new_[1641]_ ;
  assign \new_[8036]_  = \new_[1638]_  | \new_[1639]_ ;
  assign \new_[8037]_  = \new_[8036]_  | \new_[8033]_ ;
  assign \new_[8038]_  = \new_[8037]_  | \new_[8030]_ ;
  assign \new_[8039]_  = \new_[8038]_  | \new_[8025]_ ;
  assign \new_[8043]_  = \new_[1635]_  | \new_[1636]_ ;
  assign \new_[8044]_  = \new_[1637]_  | \new_[8043]_ ;
  assign \new_[8047]_  = \new_[1633]_  | \new_[1634]_ ;
  assign \new_[8050]_  = \new_[1631]_  | \new_[1632]_ ;
  assign \new_[8051]_  = \new_[8050]_  | \new_[8047]_ ;
  assign \new_[8052]_  = \new_[8051]_  | \new_[8044]_ ;
  assign \new_[8055]_  = \new_[1629]_  | \new_[1630]_ ;
  assign \new_[8058]_  = \new_[1627]_  | \new_[1628]_ ;
  assign \new_[8059]_  = \new_[8058]_  | \new_[8055]_ ;
  assign \new_[8062]_  = \new_[1625]_  | \new_[1626]_ ;
  assign \new_[8065]_  = \new_[1623]_  | \new_[1624]_ ;
  assign \new_[8066]_  = \new_[8065]_  | \new_[8062]_ ;
  assign \new_[8067]_  = \new_[8066]_  | \new_[8059]_ ;
  assign \new_[8068]_  = \new_[8067]_  | \new_[8052]_ ;
  assign \new_[8069]_  = \new_[8068]_  | \new_[8039]_ ;
  assign \new_[8073]_  = \new_[1620]_  | \new_[1621]_ ;
  assign \new_[8074]_  = \new_[1622]_  | \new_[8073]_ ;
  assign \new_[8077]_  = \new_[1618]_  | \new_[1619]_ ;
  assign \new_[8080]_  = \new_[1616]_  | \new_[1617]_ ;
  assign \new_[8081]_  = \new_[8080]_  | \new_[8077]_ ;
  assign \new_[8082]_  = \new_[8081]_  | \new_[8074]_ ;
  assign \new_[8085]_  = \new_[1614]_  | \new_[1615]_ ;
  assign \new_[8088]_  = \new_[1612]_  | \new_[1613]_ ;
  assign \new_[8089]_  = \new_[8088]_  | \new_[8085]_ ;
  assign \new_[8092]_  = \new_[1610]_  | \new_[1611]_ ;
  assign \new_[8095]_  = \new_[1608]_  | \new_[1609]_ ;
  assign \new_[8096]_  = \new_[8095]_  | \new_[8092]_ ;
  assign \new_[8097]_  = \new_[8096]_  | \new_[8089]_ ;
  assign \new_[8098]_  = \new_[8097]_  | \new_[8082]_ ;
  assign \new_[8102]_  = \new_[1605]_  | \new_[1606]_ ;
  assign \new_[8103]_  = \new_[1607]_  | \new_[8102]_ ;
  assign \new_[8106]_  = \new_[1603]_  | \new_[1604]_ ;
  assign \new_[8109]_  = \new_[1601]_  | \new_[1602]_ ;
  assign \new_[8110]_  = \new_[8109]_  | \new_[8106]_ ;
  assign \new_[8111]_  = \new_[8110]_  | \new_[8103]_ ;
  assign \new_[8114]_  = \new_[1599]_  | \new_[1600]_ ;
  assign \new_[8117]_  = \new_[1597]_  | \new_[1598]_ ;
  assign \new_[8118]_  = \new_[8117]_  | \new_[8114]_ ;
  assign \new_[8121]_  = \new_[1595]_  | \new_[1596]_ ;
  assign \new_[8124]_  = \new_[1593]_  | \new_[1594]_ ;
  assign \new_[8125]_  = \new_[8124]_  | \new_[8121]_ ;
  assign \new_[8126]_  = \new_[8125]_  | \new_[8118]_ ;
  assign \new_[8127]_  = \new_[8126]_  | \new_[8111]_ ;
  assign \new_[8128]_  = \new_[8127]_  | \new_[8098]_ ;
  assign \new_[8129]_  = \new_[8128]_  | \new_[8069]_ ;
  assign \new_[8133]_  = \new_[1590]_  | \new_[1591]_ ;
  assign \new_[8134]_  = \new_[1592]_  | \new_[8133]_ ;
  assign \new_[8137]_  = \new_[1588]_  | \new_[1589]_ ;
  assign \new_[8140]_  = \new_[1586]_  | \new_[1587]_ ;
  assign \new_[8141]_  = \new_[8140]_  | \new_[8137]_ ;
  assign \new_[8142]_  = \new_[8141]_  | \new_[8134]_ ;
  assign \new_[8146]_  = \new_[1583]_  | \new_[1584]_ ;
  assign \new_[8147]_  = \new_[1585]_  | \new_[8146]_ ;
  assign \new_[8150]_  = \new_[1581]_  | \new_[1582]_ ;
  assign \new_[8153]_  = \new_[1579]_  | \new_[1580]_ ;
  assign \new_[8154]_  = \new_[8153]_  | \new_[8150]_ ;
  assign \new_[8155]_  = \new_[8154]_  | \new_[8147]_ ;
  assign \new_[8156]_  = \new_[8155]_  | \new_[8142]_ ;
  assign \new_[8160]_  = \new_[1576]_  | \new_[1577]_ ;
  assign \new_[8161]_  = \new_[1578]_  | \new_[8160]_ ;
  assign \new_[8164]_  = \new_[1574]_  | \new_[1575]_ ;
  assign \new_[8167]_  = \new_[1572]_  | \new_[1573]_ ;
  assign \new_[8168]_  = \new_[8167]_  | \new_[8164]_ ;
  assign \new_[8169]_  = \new_[8168]_  | \new_[8161]_ ;
  assign \new_[8172]_  = \new_[1570]_  | \new_[1571]_ ;
  assign \new_[8175]_  = \new_[1568]_  | \new_[1569]_ ;
  assign \new_[8176]_  = \new_[8175]_  | \new_[8172]_ ;
  assign \new_[8179]_  = \new_[1566]_  | \new_[1567]_ ;
  assign \new_[8182]_  = \new_[1564]_  | \new_[1565]_ ;
  assign \new_[8183]_  = \new_[8182]_  | \new_[8179]_ ;
  assign \new_[8184]_  = \new_[8183]_  | \new_[8176]_ ;
  assign \new_[8185]_  = \new_[8184]_  | \new_[8169]_ ;
  assign \new_[8186]_  = \new_[8185]_  | \new_[8156]_ ;
  assign \new_[8190]_  = \new_[1561]_  | \new_[1562]_ ;
  assign \new_[8191]_  = \new_[1563]_  | \new_[8190]_ ;
  assign \new_[8194]_  = \new_[1559]_  | \new_[1560]_ ;
  assign \new_[8197]_  = \new_[1557]_  | \new_[1558]_ ;
  assign \new_[8198]_  = \new_[8197]_  | \new_[8194]_ ;
  assign \new_[8199]_  = \new_[8198]_  | \new_[8191]_ ;
  assign \new_[8202]_  = \new_[1555]_  | \new_[1556]_ ;
  assign \new_[8205]_  = \new_[1553]_  | \new_[1554]_ ;
  assign \new_[8206]_  = \new_[8205]_  | \new_[8202]_ ;
  assign \new_[8209]_  = \new_[1551]_  | \new_[1552]_ ;
  assign \new_[8212]_  = \new_[1549]_  | \new_[1550]_ ;
  assign \new_[8213]_  = \new_[8212]_  | \new_[8209]_ ;
  assign \new_[8214]_  = \new_[8213]_  | \new_[8206]_ ;
  assign \new_[8215]_  = \new_[8214]_  | \new_[8199]_ ;
  assign \new_[8219]_  = \new_[1546]_  | \new_[1547]_ ;
  assign \new_[8220]_  = \new_[1548]_  | \new_[8219]_ ;
  assign \new_[8223]_  = \new_[1544]_  | \new_[1545]_ ;
  assign \new_[8226]_  = \new_[1542]_  | \new_[1543]_ ;
  assign \new_[8227]_  = \new_[8226]_  | \new_[8223]_ ;
  assign \new_[8228]_  = \new_[8227]_  | \new_[8220]_ ;
  assign \new_[8231]_  = \new_[1540]_  | \new_[1541]_ ;
  assign \new_[8234]_  = \new_[1538]_  | \new_[1539]_ ;
  assign \new_[8235]_  = \new_[8234]_  | \new_[8231]_ ;
  assign \new_[8238]_  = \new_[1536]_  | \new_[1537]_ ;
  assign \new_[8241]_  = \new_[1534]_  | \new_[1535]_ ;
  assign \new_[8242]_  = \new_[8241]_  | \new_[8238]_ ;
  assign \new_[8243]_  = \new_[8242]_  | \new_[8235]_ ;
  assign \new_[8244]_  = \new_[8243]_  | \new_[8228]_ ;
  assign \new_[8245]_  = \new_[8244]_  | \new_[8215]_ ;
  assign \new_[8246]_  = \new_[8245]_  | \new_[8186]_ ;
  assign \new_[8247]_  = \new_[8246]_  | \new_[8129]_ ;
  assign \new_[8251]_  = \new_[1531]_  | \new_[1532]_ ;
  assign \new_[8252]_  = \new_[1533]_  | \new_[8251]_ ;
  assign \new_[8255]_  = \new_[1529]_  | \new_[1530]_ ;
  assign \new_[8258]_  = \new_[1527]_  | \new_[1528]_ ;
  assign \new_[8259]_  = \new_[8258]_  | \new_[8255]_ ;
  assign \new_[8260]_  = \new_[8259]_  | \new_[8252]_ ;
  assign \new_[8264]_  = \new_[1524]_  | \new_[1525]_ ;
  assign \new_[8265]_  = \new_[1526]_  | \new_[8264]_ ;
  assign \new_[8268]_  = \new_[1522]_  | \new_[1523]_ ;
  assign \new_[8271]_  = \new_[1520]_  | \new_[1521]_ ;
  assign \new_[8272]_  = \new_[8271]_  | \new_[8268]_ ;
  assign \new_[8273]_  = \new_[8272]_  | \new_[8265]_ ;
  assign \new_[8274]_  = \new_[8273]_  | \new_[8260]_ ;
  assign \new_[8278]_  = \new_[1517]_  | \new_[1518]_ ;
  assign \new_[8279]_  = \new_[1519]_  | \new_[8278]_ ;
  assign \new_[8282]_  = \new_[1515]_  | \new_[1516]_ ;
  assign \new_[8285]_  = \new_[1513]_  | \new_[1514]_ ;
  assign \new_[8286]_  = \new_[8285]_  | \new_[8282]_ ;
  assign \new_[8287]_  = \new_[8286]_  | \new_[8279]_ ;
  assign \new_[8290]_  = \new_[1511]_  | \new_[1512]_ ;
  assign \new_[8293]_  = \new_[1509]_  | \new_[1510]_ ;
  assign \new_[8294]_  = \new_[8293]_  | \new_[8290]_ ;
  assign \new_[8297]_  = \new_[1507]_  | \new_[1508]_ ;
  assign \new_[8300]_  = \new_[1505]_  | \new_[1506]_ ;
  assign \new_[8301]_  = \new_[8300]_  | \new_[8297]_ ;
  assign \new_[8302]_  = \new_[8301]_  | \new_[8294]_ ;
  assign \new_[8303]_  = \new_[8302]_  | \new_[8287]_ ;
  assign \new_[8304]_  = \new_[8303]_  | \new_[8274]_ ;
  assign \new_[8308]_  = \new_[1502]_  | \new_[1503]_ ;
  assign \new_[8309]_  = \new_[1504]_  | \new_[8308]_ ;
  assign \new_[8312]_  = \new_[1500]_  | \new_[1501]_ ;
  assign \new_[8315]_  = \new_[1498]_  | \new_[1499]_ ;
  assign \new_[8316]_  = \new_[8315]_  | \new_[8312]_ ;
  assign \new_[8317]_  = \new_[8316]_  | \new_[8309]_ ;
  assign \new_[8320]_  = \new_[1496]_  | \new_[1497]_ ;
  assign \new_[8323]_  = \new_[1494]_  | \new_[1495]_ ;
  assign \new_[8324]_  = \new_[8323]_  | \new_[8320]_ ;
  assign \new_[8327]_  = \new_[1492]_  | \new_[1493]_ ;
  assign \new_[8330]_  = \new_[1490]_  | \new_[1491]_ ;
  assign \new_[8331]_  = \new_[8330]_  | \new_[8327]_ ;
  assign \new_[8332]_  = \new_[8331]_  | \new_[8324]_ ;
  assign \new_[8333]_  = \new_[8332]_  | \new_[8317]_ ;
  assign \new_[8337]_  = \new_[1487]_  | \new_[1488]_ ;
  assign \new_[8338]_  = \new_[1489]_  | \new_[8337]_ ;
  assign \new_[8341]_  = \new_[1485]_  | \new_[1486]_ ;
  assign \new_[8344]_  = \new_[1483]_  | \new_[1484]_ ;
  assign \new_[8345]_  = \new_[8344]_  | \new_[8341]_ ;
  assign \new_[8346]_  = \new_[8345]_  | \new_[8338]_ ;
  assign \new_[8349]_  = \new_[1481]_  | \new_[1482]_ ;
  assign \new_[8352]_  = \new_[1479]_  | \new_[1480]_ ;
  assign \new_[8353]_  = \new_[8352]_  | \new_[8349]_ ;
  assign \new_[8356]_  = \new_[1477]_  | \new_[1478]_ ;
  assign \new_[8359]_  = \new_[1475]_  | \new_[1476]_ ;
  assign \new_[8360]_  = \new_[8359]_  | \new_[8356]_ ;
  assign \new_[8361]_  = \new_[8360]_  | \new_[8353]_ ;
  assign \new_[8362]_  = \new_[8361]_  | \new_[8346]_ ;
  assign \new_[8363]_  = \new_[8362]_  | \new_[8333]_ ;
  assign \new_[8364]_  = \new_[8363]_  | \new_[8304]_ ;
  assign \new_[8368]_  = \new_[1472]_  | \new_[1473]_ ;
  assign \new_[8369]_  = \new_[1474]_  | \new_[8368]_ ;
  assign \new_[8372]_  = \new_[1470]_  | \new_[1471]_ ;
  assign \new_[8375]_  = \new_[1468]_  | \new_[1469]_ ;
  assign \new_[8376]_  = \new_[8375]_  | \new_[8372]_ ;
  assign \new_[8377]_  = \new_[8376]_  | \new_[8369]_ ;
  assign \new_[8381]_  = \new_[1465]_  | \new_[1466]_ ;
  assign \new_[8382]_  = \new_[1467]_  | \new_[8381]_ ;
  assign \new_[8385]_  = \new_[1463]_  | \new_[1464]_ ;
  assign \new_[8388]_  = \new_[1461]_  | \new_[1462]_ ;
  assign \new_[8389]_  = \new_[8388]_  | \new_[8385]_ ;
  assign \new_[8390]_  = \new_[8389]_  | \new_[8382]_ ;
  assign \new_[8391]_  = \new_[8390]_  | \new_[8377]_ ;
  assign \new_[8395]_  = \new_[1458]_  | \new_[1459]_ ;
  assign \new_[8396]_  = \new_[1460]_  | \new_[8395]_ ;
  assign \new_[8399]_  = \new_[1456]_  | \new_[1457]_ ;
  assign \new_[8402]_  = \new_[1454]_  | \new_[1455]_ ;
  assign \new_[8403]_  = \new_[8402]_  | \new_[8399]_ ;
  assign \new_[8404]_  = \new_[8403]_  | \new_[8396]_ ;
  assign \new_[8407]_  = \new_[1452]_  | \new_[1453]_ ;
  assign \new_[8410]_  = \new_[1450]_  | \new_[1451]_ ;
  assign \new_[8411]_  = \new_[8410]_  | \new_[8407]_ ;
  assign \new_[8414]_  = \new_[1448]_  | \new_[1449]_ ;
  assign \new_[8417]_  = \new_[1446]_  | \new_[1447]_ ;
  assign \new_[8418]_  = \new_[8417]_  | \new_[8414]_ ;
  assign \new_[8419]_  = \new_[8418]_  | \new_[8411]_ ;
  assign \new_[8420]_  = \new_[8419]_  | \new_[8404]_ ;
  assign \new_[8421]_  = \new_[8420]_  | \new_[8391]_ ;
  assign \new_[8425]_  = \new_[1443]_  | \new_[1444]_ ;
  assign \new_[8426]_  = \new_[1445]_  | \new_[8425]_ ;
  assign \new_[8429]_  = \new_[1441]_  | \new_[1442]_ ;
  assign \new_[8432]_  = \new_[1439]_  | \new_[1440]_ ;
  assign \new_[8433]_  = \new_[8432]_  | \new_[8429]_ ;
  assign \new_[8434]_  = \new_[8433]_  | \new_[8426]_ ;
  assign \new_[8437]_  = \new_[1437]_  | \new_[1438]_ ;
  assign \new_[8440]_  = \new_[1435]_  | \new_[1436]_ ;
  assign \new_[8441]_  = \new_[8440]_  | \new_[8437]_ ;
  assign \new_[8444]_  = \new_[1433]_  | \new_[1434]_ ;
  assign \new_[8447]_  = \new_[1431]_  | \new_[1432]_ ;
  assign \new_[8448]_  = \new_[8447]_  | \new_[8444]_ ;
  assign \new_[8449]_  = \new_[8448]_  | \new_[8441]_ ;
  assign \new_[8450]_  = \new_[8449]_  | \new_[8434]_ ;
  assign \new_[8454]_  = \new_[1428]_  | \new_[1429]_ ;
  assign \new_[8455]_  = \new_[1430]_  | \new_[8454]_ ;
  assign \new_[8458]_  = \new_[1426]_  | \new_[1427]_ ;
  assign \new_[8461]_  = \new_[1424]_  | \new_[1425]_ ;
  assign \new_[8462]_  = \new_[8461]_  | \new_[8458]_ ;
  assign \new_[8463]_  = \new_[8462]_  | \new_[8455]_ ;
  assign \new_[8466]_  = \new_[1422]_  | \new_[1423]_ ;
  assign \new_[8469]_  = \new_[1420]_  | \new_[1421]_ ;
  assign \new_[8470]_  = \new_[8469]_  | \new_[8466]_ ;
  assign \new_[8473]_  = \new_[1418]_  | \new_[1419]_ ;
  assign \new_[8476]_  = \new_[1416]_  | \new_[1417]_ ;
  assign \new_[8477]_  = \new_[8476]_  | \new_[8473]_ ;
  assign \new_[8478]_  = \new_[8477]_  | \new_[8470]_ ;
  assign \new_[8479]_  = \new_[8478]_  | \new_[8463]_ ;
  assign \new_[8480]_  = \new_[8479]_  | \new_[8450]_ ;
  assign \new_[8481]_  = \new_[8480]_  | \new_[8421]_ ;
  assign \new_[8482]_  = \new_[8481]_  | \new_[8364]_ ;
  assign \new_[8483]_  = \new_[8482]_  | \new_[8247]_ ;
  assign \new_[8484]_  = \new_[8483]_  | \new_[8012]_ ;
  assign \new_[8488]_  = \new_[1413]_  | \new_[1414]_ ;
  assign \new_[8489]_  = \new_[1415]_  | \new_[8488]_ ;
  assign \new_[8492]_  = \new_[1411]_  | \new_[1412]_ ;
  assign \new_[8495]_  = \new_[1409]_  | \new_[1410]_ ;
  assign \new_[8496]_  = \new_[8495]_  | \new_[8492]_ ;
  assign \new_[8497]_  = \new_[8496]_  | \new_[8489]_ ;
  assign \new_[8501]_  = \new_[1406]_  | \new_[1407]_ ;
  assign \new_[8502]_  = \new_[1408]_  | \new_[8501]_ ;
  assign \new_[8505]_  = \new_[1404]_  | \new_[1405]_ ;
  assign \new_[8508]_  = \new_[1402]_  | \new_[1403]_ ;
  assign \new_[8509]_  = \new_[8508]_  | \new_[8505]_ ;
  assign \new_[8510]_  = \new_[8509]_  | \new_[8502]_ ;
  assign \new_[8511]_  = \new_[8510]_  | \new_[8497]_ ;
  assign \new_[8515]_  = \new_[1399]_  | \new_[1400]_ ;
  assign \new_[8516]_  = \new_[1401]_  | \new_[8515]_ ;
  assign \new_[8519]_  = \new_[1397]_  | \new_[1398]_ ;
  assign \new_[8522]_  = \new_[1395]_  | \new_[1396]_ ;
  assign \new_[8523]_  = \new_[8522]_  | \new_[8519]_ ;
  assign \new_[8524]_  = \new_[8523]_  | \new_[8516]_ ;
  assign \new_[8527]_  = \new_[1393]_  | \new_[1394]_ ;
  assign \new_[8530]_  = \new_[1391]_  | \new_[1392]_ ;
  assign \new_[8531]_  = \new_[8530]_  | \new_[8527]_ ;
  assign \new_[8534]_  = \new_[1389]_  | \new_[1390]_ ;
  assign \new_[8537]_  = \new_[1387]_  | \new_[1388]_ ;
  assign \new_[8538]_  = \new_[8537]_  | \new_[8534]_ ;
  assign \new_[8539]_  = \new_[8538]_  | \new_[8531]_ ;
  assign \new_[8540]_  = \new_[8539]_  | \new_[8524]_ ;
  assign \new_[8541]_  = \new_[8540]_  | \new_[8511]_ ;
  assign \new_[8545]_  = \new_[1384]_  | \new_[1385]_ ;
  assign \new_[8546]_  = \new_[1386]_  | \new_[8545]_ ;
  assign \new_[8549]_  = \new_[1382]_  | \new_[1383]_ ;
  assign \new_[8552]_  = \new_[1380]_  | \new_[1381]_ ;
  assign \new_[8553]_  = \new_[8552]_  | \new_[8549]_ ;
  assign \new_[8554]_  = \new_[8553]_  | \new_[8546]_ ;
  assign \new_[8557]_  = \new_[1378]_  | \new_[1379]_ ;
  assign \new_[8560]_  = \new_[1376]_  | \new_[1377]_ ;
  assign \new_[8561]_  = \new_[8560]_  | \new_[8557]_ ;
  assign \new_[8564]_  = \new_[1374]_  | \new_[1375]_ ;
  assign \new_[8567]_  = \new_[1372]_  | \new_[1373]_ ;
  assign \new_[8568]_  = \new_[8567]_  | \new_[8564]_ ;
  assign \new_[8569]_  = \new_[8568]_  | \new_[8561]_ ;
  assign \new_[8570]_  = \new_[8569]_  | \new_[8554]_ ;
  assign \new_[8574]_  = \new_[1369]_  | \new_[1370]_ ;
  assign \new_[8575]_  = \new_[1371]_  | \new_[8574]_ ;
  assign \new_[8578]_  = \new_[1367]_  | \new_[1368]_ ;
  assign \new_[8581]_  = \new_[1365]_  | \new_[1366]_ ;
  assign \new_[8582]_  = \new_[8581]_  | \new_[8578]_ ;
  assign \new_[8583]_  = \new_[8582]_  | \new_[8575]_ ;
  assign \new_[8586]_  = \new_[1363]_  | \new_[1364]_ ;
  assign \new_[8589]_  = \new_[1361]_  | \new_[1362]_ ;
  assign \new_[8590]_  = \new_[8589]_  | \new_[8586]_ ;
  assign \new_[8593]_  = \new_[1359]_  | \new_[1360]_ ;
  assign \new_[8596]_  = \new_[1357]_  | \new_[1358]_ ;
  assign \new_[8597]_  = \new_[8596]_  | \new_[8593]_ ;
  assign \new_[8598]_  = \new_[8597]_  | \new_[8590]_ ;
  assign \new_[8599]_  = \new_[8598]_  | \new_[8583]_ ;
  assign \new_[8600]_  = \new_[8599]_  | \new_[8570]_ ;
  assign \new_[8601]_  = \new_[8600]_  | \new_[8541]_ ;
  assign \new_[8605]_  = \new_[1354]_  | \new_[1355]_ ;
  assign \new_[8606]_  = \new_[1356]_  | \new_[8605]_ ;
  assign \new_[8609]_  = \new_[1352]_  | \new_[1353]_ ;
  assign \new_[8612]_  = \new_[1350]_  | \new_[1351]_ ;
  assign \new_[8613]_  = \new_[8612]_  | \new_[8609]_ ;
  assign \new_[8614]_  = \new_[8613]_  | \new_[8606]_ ;
  assign \new_[8618]_  = \new_[1347]_  | \new_[1348]_ ;
  assign \new_[8619]_  = \new_[1349]_  | \new_[8618]_ ;
  assign \new_[8622]_  = \new_[1345]_  | \new_[1346]_ ;
  assign \new_[8625]_  = \new_[1343]_  | \new_[1344]_ ;
  assign \new_[8626]_  = \new_[8625]_  | \new_[8622]_ ;
  assign \new_[8627]_  = \new_[8626]_  | \new_[8619]_ ;
  assign \new_[8628]_  = \new_[8627]_  | \new_[8614]_ ;
  assign \new_[8632]_  = \new_[1340]_  | \new_[1341]_ ;
  assign \new_[8633]_  = \new_[1342]_  | \new_[8632]_ ;
  assign \new_[8636]_  = \new_[1338]_  | \new_[1339]_ ;
  assign \new_[8639]_  = \new_[1336]_  | \new_[1337]_ ;
  assign \new_[8640]_  = \new_[8639]_  | \new_[8636]_ ;
  assign \new_[8641]_  = \new_[8640]_  | \new_[8633]_ ;
  assign \new_[8644]_  = \new_[1334]_  | \new_[1335]_ ;
  assign \new_[8647]_  = \new_[1332]_  | \new_[1333]_ ;
  assign \new_[8648]_  = \new_[8647]_  | \new_[8644]_ ;
  assign \new_[8651]_  = \new_[1330]_  | \new_[1331]_ ;
  assign \new_[8654]_  = \new_[1328]_  | \new_[1329]_ ;
  assign \new_[8655]_  = \new_[8654]_  | \new_[8651]_ ;
  assign \new_[8656]_  = \new_[8655]_  | \new_[8648]_ ;
  assign \new_[8657]_  = \new_[8656]_  | \new_[8641]_ ;
  assign \new_[8658]_  = \new_[8657]_  | \new_[8628]_ ;
  assign \new_[8662]_  = \new_[1325]_  | \new_[1326]_ ;
  assign \new_[8663]_  = \new_[1327]_  | \new_[8662]_ ;
  assign \new_[8666]_  = \new_[1323]_  | \new_[1324]_ ;
  assign \new_[8669]_  = \new_[1321]_  | \new_[1322]_ ;
  assign \new_[8670]_  = \new_[8669]_  | \new_[8666]_ ;
  assign \new_[8671]_  = \new_[8670]_  | \new_[8663]_ ;
  assign \new_[8674]_  = \new_[1319]_  | \new_[1320]_ ;
  assign \new_[8677]_  = \new_[1317]_  | \new_[1318]_ ;
  assign \new_[8678]_  = \new_[8677]_  | \new_[8674]_ ;
  assign \new_[8681]_  = \new_[1315]_  | \new_[1316]_ ;
  assign \new_[8684]_  = \new_[1313]_  | \new_[1314]_ ;
  assign \new_[8685]_  = \new_[8684]_  | \new_[8681]_ ;
  assign \new_[8686]_  = \new_[8685]_  | \new_[8678]_ ;
  assign \new_[8687]_  = \new_[8686]_  | \new_[8671]_ ;
  assign \new_[8691]_  = \new_[1310]_  | \new_[1311]_ ;
  assign \new_[8692]_  = \new_[1312]_  | \new_[8691]_ ;
  assign \new_[8695]_  = \new_[1308]_  | \new_[1309]_ ;
  assign \new_[8698]_  = \new_[1306]_  | \new_[1307]_ ;
  assign \new_[8699]_  = \new_[8698]_  | \new_[8695]_ ;
  assign \new_[8700]_  = \new_[8699]_  | \new_[8692]_ ;
  assign \new_[8703]_  = \new_[1304]_  | \new_[1305]_ ;
  assign \new_[8706]_  = \new_[1302]_  | \new_[1303]_ ;
  assign \new_[8707]_  = \new_[8706]_  | \new_[8703]_ ;
  assign \new_[8710]_  = \new_[1300]_  | \new_[1301]_ ;
  assign \new_[8713]_  = \new_[1298]_  | \new_[1299]_ ;
  assign \new_[8714]_  = \new_[8713]_  | \new_[8710]_ ;
  assign \new_[8715]_  = \new_[8714]_  | \new_[8707]_ ;
  assign \new_[8716]_  = \new_[8715]_  | \new_[8700]_ ;
  assign \new_[8717]_  = \new_[8716]_  | \new_[8687]_ ;
  assign \new_[8718]_  = \new_[8717]_  | \new_[8658]_ ;
  assign \new_[8719]_  = \new_[8718]_  | \new_[8601]_ ;
  assign \new_[8723]_  = \new_[1295]_  | \new_[1296]_ ;
  assign \new_[8724]_  = \new_[1297]_  | \new_[8723]_ ;
  assign \new_[8727]_  = \new_[1293]_  | \new_[1294]_ ;
  assign \new_[8730]_  = \new_[1291]_  | \new_[1292]_ ;
  assign \new_[8731]_  = \new_[8730]_  | \new_[8727]_ ;
  assign \new_[8732]_  = \new_[8731]_  | \new_[8724]_ ;
  assign \new_[8736]_  = \new_[1288]_  | \new_[1289]_ ;
  assign \new_[8737]_  = \new_[1290]_  | \new_[8736]_ ;
  assign \new_[8740]_  = \new_[1286]_  | \new_[1287]_ ;
  assign \new_[8743]_  = \new_[1284]_  | \new_[1285]_ ;
  assign \new_[8744]_  = \new_[8743]_  | \new_[8740]_ ;
  assign \new_[8745]_  = \new_[8744]_  | \new_[8737]_ ;
  assign \new_[8746]_  = \new_[8745]_  | \new_[8732]_ ;
  assign \new_[8750]_  = \new_[1281]_  | \new_[1282]_ ;
  assign \new_[8751]_  = \new_[1283]_  | \new_[8750]_ ;
  assign \new_[8754]_  = \new_[1279]_  | \new_[1280]_ ;
  assign \new_[8757]_  = \new_[1277]_  | \new_[1278]_ ;
  assign \new_[8758]_  = \new_[8757]_  | \new_[8754]_ ;
  assign \new_[8759]_  = \new_[8758]_  | \new_[8751]_ ;
  assign \new_[8762]_  = \new_[1275]_  | \new_[1276]_ ;
  assign \new_[8765]_  = \new_[1273]_  | \new_[1274]_ ;
  assign \new_[8766]_  = \new_[8765]_  | \new_[8762]_ ;
  assign \new_[8769]_  = \new_[1271]_  | \new_[1272]_ ;
  assign \new_[8772]_  = \new_[1269]_  | \new_[1270]_ ;
  assign \new_[8773]_  = \new_[8772]_  | \new_[8769]_ ;
  assign \new_[8774]_  = \new_[8773]_  | \new_[8766]_ ;
  assign \new_[8775]_  = \new_[8774]_  | \new_[8759]_ ;
  assign \new_[8776]_  = \new_[8775]_  | \new_[8746]_ ;
  assign \new_[8780]_  = \new_[1266]_  | \new_[1267]_ ;
  assign \new_[8781]_  = \new_[1268]_  | \new_[8780]_ ;
  assign \new_[8784]_  = \new_[1264]_  | \new_[1265]_ ;
  assign \new_[8787]_  = \new_[1262]_  | \new_[1263]_ ;
  assign \new_[8788]_  = \new_[8787]_  | \new_[8784]_ ;
  assign \new_[8789]_  = \new_[8788]_  | \new_[8781]_ ;
  assign \new_[8792]_  = \new_[1260]_  | \new_[1261]_ ;
  assign \new_[8795]_  = \new_[1258]_  | \new_[1259]_ ;
  assign \new_[8796]_  = \new_[8795]_  | \new_[8792]_ ;
  assign \new_[8799]_  = \new_[1256]_  | \new_[1257]_ ;
  assign \new_[8802]_  = \new_[1254]_  | \new_[1255]_ ;
  assign \new_[8803]_  = \new_[8802]_  | \new_[8799]_ ;
  assign \new_[8804]_  = \new_[8803]_  | \new_[8796]_ ;
  assign \new_[8805]_  = \new_[8804]_  | \new_[8789]_ ;
  assign \new_[8809]_  = \new_[1251]_  | \new_[1252]_ ;
  assign \new_[8810]_  = \new_[1253]_  | \new_[8809]_ ;
  assign \new_[8813]_  = \new_[1249]_  | \new_[1250]_ ;
  assign \new_[8816]_  = \new_[1247]_  | \new_[1248]_ ;
  assign \new_[8817]_  = \new_[8816]_  | \new_[8813]_ ;
  assign \new_[8818]_  = \new_[8817]_  | \new_[8810]_ ;
  assign \new_[8821]_  = \new_[1245]_  | \new_[1246]_ ;
  assign \new_[8824]_  = \new_[1243]_  | \new_[1244]_ ;
  assign \new_[8825]_  = \new_[8824]_  | \new_[8821]_ ;
  assign \new_[8828]_  = \new_[1241]_  | \new_[1242]_ ;
  assign \new_[8831]_  = \new_[1239]_  | \new_[1240]_ ;
  assign \new_[8832]_  = \new_[8831]_  | \new_[8828]_ ;
  assign \new_[8833]_  = \new_[8832]_  | \new_[8825]_ ;
  assign \new_[8834]_  = \new_[8833]_  | \new_[8818]_ ;
  assign \new_[8835]_  = \new_[8834]_  | \new_[8805]_ ;
  assign \new_[8836]_  = \new_[8835]_  | \new_[8776]_ ;
  assign \new_[8840]_  = \new_[1236]_  | \new_[1237]_ ;
  assign \new_[8841]_  = \new_[1238]_  | \new_[8840]_ ;
  assign \new_[8844]_  = \new_[1234]_  | \new_[1235]_ ;
  assign \new_[8847]_  = \new_[1232]_  | \new_[1233]_ ;
  assign \new_[8848]_  = \new_[8847]_  | \new_[8844]_ ;
  assign \new_[8849]_  = \new_[8848]_  | \new_[8841]_ ;
  assign \new_[8853]_  = \new_[1229]_  | \new_[1230]_ ;
  assign \new_[8854]_  = \new_[1231]_  | \new_[8853]_ ;
  assign \new_[8857]_  = \new_[1227]_  | \new_[1228]_ ;
  assign \new_[8860]_  = \new_[1225]_  | \new_[1226]_ ;
  assign \new_[8861]_  = \new_[8860]_  | \new_[8857]_ ;
  assign \new_[8862]_  = \new_[8861]_  | \new_[8854]_ ;
  assign \new_[8863]_  = \new_[8862]_  | \new_[8849]_ ;
  assign \new_[8867]_  = \new_[1222]_  | \new_[1223]_ ;
  assign \new_[8868]_  = \new_[1224]_  | \new_[8867]_ ;
  assign \new_[8871]_  = \new_[1220]_  | \new_[1221]_ ;
  assign \new_[8874]_  = \new_[1218]_  | \new_[1219]_ ;
  assign \new_[8875]_  = \new_[8874]_  | \new_[8871]_ ;
  assign \new_[8876]_  = \new_[8875]_  | \new_[8868]_ ;
  assign \new_[8879]_  = \new_[1216]_  | \new_[1217]_ ;
  assign \new_[8882]_  = \new_[1214]_  | \new_[1215]_ ;
  assign \new_[8883]_  = \new_[8882]_  | \new_[8879]_ ;
  assign \new_[8886]_  = \new_[1212]_  | \new_[1213]_ ;
  assign \new_[8889]_  = \new_[1210]_  | \new_[1211]_ ;
  assign \new_[8890]_  = \new_[8889]_  | \new_[8886]_ ;
  assign \new_[8891]_  = \new_[8890]_  | \new_[8883]_ ;
  assign \new_[8892]_  = \new_[8891]_  | \new_[8876]_ ;
  assign \new_[8893]_  = \new_[8892]_  | \new_[8863]_ ;
  assign \new_[8897]_  = \new_[1207]_  | \new_[1208]_ ;
  assign \new_[8898]_  = \new_[1209]_  | \new_[8897]_ ;
  assign \new_[8901]_  = \new_[1205]_  | \new_[1206]_ ;
  assign \new_[8904]_  = \new_[1203]_  | \new_[1204]_ ;
  assign \new_[8905]_  = \new_[8904]_  | \new_[8901]_ ;
  assign \new_[8906]_  = \new_[8905]_  | \new_[8898]_ ;
  assign \new_[8909]_  = \new_[1201]_  | \new_[1202]_ ;
  assign \new_[8912]_  = \new_[1199]_  | \new_[1200]_ ;
  assign \new_[8913]_  = \new_[8912]_  | \new_[8909]_ ;
  assign \new_[8916]_  = \new_[1197]_  | \new_[1198]_ ;
  assign \new_[8919]_  = \new_[1195]_  | \new_[1196]_ ;
  assign \new_[8920]_  = \new_[8919]_  | \new_[8916]_ ;
  assign \new_[8921]_  = \new_[8920]_  | \new_[8913]_ ;
  assign \new_[8922]_  = \new_[8921]_  | \new_[8906]_ ;
  assign \new_[8926]_  = \new_[1192]_  | \new_[1193]_ ;
  assign \new_[8927]_  = \new_[1194]_  | \new_[8926]_ ;
  assign \new_[8930]_  = \new_[1190]_  | \new_[1191]_ ;
  assign \new_[8933]_  = \new_[1188]_  | \new_[1189]_ ;
  assign \new_[8934]_  = \new_[8933]_  | \new_[8930]_ ;
  assign \new_[8935]_  = \new_[8934]_  | \new_[8927]_ ;
  assign \new_[8938]_  = \new_[1186]_  | \new_[1187]_ ;
  assign \new_[8941]_  = \new_[1184]_  | \new_[1185]_ ;
  assign \new_[8942]_  = \new_[8941]_  | \new_[8938]_ ;
  assign \new_[8945]_  = \new_[1182]_  | \new_[1183]_ ;
  assign \new_[8948]_  = \new_[1180]_  | \new_[1181]_ ;
  assign \new_[8949]_  = \new_[8948]_  | \new_[8945]_ ;
  assign \new_[8950]_  = \new_[8949]_  | \new_[8942]_ ;
  assign \new_[8951]_  = \new_[8950]_  | \new_[8935]_ ;
  assign \new_[8952]_  = \new_[8951]_  | \new_[8922]_ ;
  assign \new_[8953]_  = \new_[8952]_  | \new_[8893]_ ;
  assign \new_[8954]_  = \new_[8953]_  | \new_[8836]_ ;
  assign \new_[8955]_  = \new_[8954]_  | \new_[8719]_ ;
  assign \new_[8959]_  = \new_[1177]_  | \new_[1178]_ ;
  assign \new_[8960]_  = \new_[1179]_  | \new_[8959]_ ;
  assign \new_[8963]_  = \new_[1175]_  | \new_[1176]_ ;
  assign \new_[8966]_  = \new_[1173]_  | \new_[1174]_ ;
  assign \new_[8967]_  = \new_[8966]_  | \new_[8963]_ ;
  assign \new_[8968]_  = \new_[8967]_  | \new_[8960]_ ;
  assign \new_[8972]_  = \new_[1170]_  | \new_[1171]_ ;
  assign \new_[8973]_  = \new_[1172]_  | \new_[8972]_ ;
  assign \new_[8976]_  = \new_[1168]_  | \new_[1169]_ ;
  assign \new_[8979]_  = \new_[1166]_  | \new_[1167]_ ;
  assign \new_[8980]_  = \new_[8979]_  | \new_[8976]_ ;
  assign \new_[8981]_  = \new_[8980]_  | \new_[8973]_ ;
  assign \new_[8982]_  = \new_[8981]_  | \new_[8968]_ ;
  assign \new_[8986]_  = \new_[1163]_  | \new_[1164]_ ;
  assign \new_[8987]_  = \new_[1165]_  | \new_[8986]_ ;
  assign \new_[8990]_  = \new_[1161]_  | \new_[1162]_ ;
  assign \new_[8993]_  = \new_[1159]_  | \new_[1160]_ ;
  assign \new_[8994]_  = \new_[8993]_  | \new_[8990]_ ;
  assign \new_[8995]_  = \new_[8994]_  | \new_[8987]_ ;
  assign \new_[8998]_  = \new_[1157]_  | \new_[1158]_ ;
  assign \new_[9001]_  = \new_[1155]_  | \new_[1156]_ ;
  assign \new_[9002]_  = \new_[9001]_  | \new_[8998]_ ;
  assign \new_[9005]_  = \new_[1153]_  | \new_[1154]_ ;
  assign \new_[9008]_  = \new_[1151]_  | \new_[1152]_ ;
  assign \new_[9009]_  = \new_[9008]_  | \new_[9005]_ ;
  assign \new_[9010]_  = \new_[9009]_  | \new_[9002]_ ;
  assign \new_[9011]_  = \new_[9010]_  | \new_[8995]_ ;
  assign \new_[9012]_  = \new_[9011]_  | \new_[8982]_ ;
  assign \new_[9016]_  = \new_[1148]_  | \new_[1149]_ ;
  assign \new_[9017]_  = \new_[1150]_  | \new_[9016]_ ;
  assign \new_[9020]_  = \new_[1146]_  | \new_[1147]_ ;
  assign \new_[9023]_  = \new_[1144]_  | \new_[1145]_ ;
  assign \new_[9024]_  = \new_[9023]_  | \new_[9020]_ ;
  assign \new_[9025]_  = \new_[9024]_  | \new_[9017]_ ;
  assign \new_[9028]_  = \new_[1142]_  | \new_[1143]_ ;
  assign \new_[9031]_  = \new_[1140]_  | \new_[1141]_ ;
  assign \new_[9032]_  = \new_[9031]_  | \new_[9028]_ ;
  assign \new_[9035]_  = \new_[1138]_  | \new_[1139]_ ;
  assign \new_[9038]_  = \new_[1136]_  | \new_[1137]_ ;
  assign \new_[9039]_  = \new_[9038]_  | \new_[9035]_ ;
  assign \new_[9040]_  = \new_[9039]_  | \new_[9032]_ ;
  assign \new_[9041]_  = \new_[9040]_  | \new_[9025]_ ;
  assign \new_[9045]_  = \new_[1133]_  | \new_[1134]_ ;
  assign \new_[9046]_  = \new_[1135]_  | \new_[9045]_ ;
  assign \new_[9049]_  = \new_[1131]_  | \new_[1132]_ ;
  assign \new_[9052]_  = \new_[1129]_  | \new_[1130]_ ;
  assign \new_[9053]_  = \new_[9052]_  | \new_[9049]_ ;
  assign \new_[9054]_  = \new_[9053]_  | \new_[9046]_ ;
  assign \new_[9057]_  = \new_[1127]_  | \new_[1128]_ ;
  assign \new_[9060]_  = \new_[1125]_  | \new_[1126]_ ;
  assign \new_[9061]_  = \new_[9060]_  | \new_[9057]_ ;
  assign \new_[9064]_  = \new_[1123]_  | \new_[1124]_ ;
  assign \new_[9067]_  = \new_[1121]_  | \new_[1122]_ ;
  assign \new_[9068]_  = \new_[9067]_  | \new_[9064]_ ;
  assign \new_[9069]_  = \new_[9068]_  | \new_[9061]_ ;
  assign \new_[9070]_  = \new_[9069]_  | \new_[9054]_ ;
  assign \new_[9071]_  = \new_[9070]_  | \new_[9041]_ ;
  assign \new_[9072]_  = \new_[9071]_  | \new_[9012]_ ;
  assign \new_[9076]_  = \new_[1118]_  | \new_[1119]_ ;
  assign \new_[9077]_  = \new_[1120]_  | \new_[9076]_ ;
  assign \new_[9080]_  = \new_[1116]_  | \new_[1117]_ ;
  assign \new_[9083]_  = \new_[1114]_  | \new_[1115]_ ;
  assign \new_[9084]_  = \new_[9083]_  | \new_[9080]_ ;
  assign \new_[9085]_  = \new_[9084]_  | \new_[9077]_ ;
  assign \new_[9089]_  = \new_[1111]_  | \new_[1112]_ ;
  assign \new_[9090]_  = \new_[1113]_  | \new_[9089]_ ;
  assign \new_[9093]_  = \new_[1109]_  | \new_[1110]_ ;
  assign \new_[9096]_  = \new_[1107]_  | \new_[1108]_ ;
  assign \new_[9097]_  = \new_[9096]_  | \new_[9093]_ ;
  assign \new_[9098]_  = \new_[9097]_  | \new_[9090]_ ;
  assign \new_[9099]_  = \new_[9098]_  | \new_[9085]_ ;
  assign \new_[9103]_  = \new_[1104]_  | \new_[1105]_ ;
  assign \new_[9104]_  = \new_[1106]_  | \new_[9103]_ ;
  assign \new_[9107]_  = \new_[1102]_  | \new_[1103]_ ;
  assign \new_[9110]_  = \new_[1100]_  | \new_[1101]_ ;
  assign \new_[9111]_  = \new_[9110]_  | \new_[9107]_ ;
  assign \new_[9112]_  = \new_[9111]_  | \new_[9104]_ ;
  assign \new_[9115]_  = \new_[1098]_  | \new_[1099]_ ;
  assign \new_[9118]_  = \new_[1096]_  | \new_[1097]_ ;
  assign \new_[9119]_  = \new_[9118]_  | \new_[9115]_ ;
  assign \new_[9122]_  = \new_[1094]_  | \new_[1095]_ ;
  assign \new_[9125]_  = \new_[1092]_  | \new_[1093]_ ;
  assign \new_[9126]_  = \new_[9125]_  | \new_[9122]_ ;
  assign \new_[9127]_  = \new_[9126]_  | \new_[9119]_ ;
  assign \new_[9128]_  = \new_[9127]_  | \new_[9112]_ ;
  assign \new_[9129]_  = \new_[9128]_  | \new_[9099]_ ;
  assign \new_[9133]_  = \new_[1089]_  | \new_[1090]_ ;
  assign \new_[9134]_  = \new_[1091]_  | \new_[9133]_ ;
  assign \new_[9137]_  = \new_[1087]_  | \new_[1088]_ ;
  assign \new_[9140]_  = \new_[1085]_  | \new_[1086]_ ;
  assign \new_[9141]_  = \new_[9140]_  | \new_[9137]_ ;
  assign \new_[9142]_  = \new_[9141]_  | \new_[9134]_ ;
  assign \new_[9145]_  = \new_[1083]_  | \new_[1084]_ ;
  assign \new_[9148]_  = \new_[1081]_  | \new_[1082]_ ;
  assign \new_[9149]_  = \new_[9148]_  | \new_[9145]_ ;
  assign \new_[9152]_  = \new_[1079]_  | \new_[1080]_ ;
  assign \new_[9155]_  = \new_[1077]_  | \new_[1078]_ ;
  assign \new_[9156]_  = \new_[9155]_  | \new_[9152]_ ;
  assign \new_[9157]_  = \new_[9156]_  | \new_[9149]_ ;
  assign \new_[9158]_  = \new_[9157]_  | \new_[9142]_ ;
  assign \new_[9162]_  = \new_[1074]_  | \new_[1075]_ ;
  assign \new_[9163]_  = \new_[1076]_  | \new_[9162]_ ;
  assign \new_[9166]_  = \new_[1072]_  | \new_[1073]_ ;
  assign \new_[9169]_  = \new_[1070]_  | \new_[1071]_ ;
  assign \new_[9170]_  = \new_[9169]_  | \new_[9166]_ ;
  assign \new_[9171]_  = \new_[9170]_  | \new_[9163]_ ;
  assign \new_[9174]_  = \new_[1068]_  | \new_[1069]_ ;
  assign \new_[9177]_  = \new_[1066]_  | \new_[1067]_ ;
  assign \new_[9178]_  = \new_[9177]_  | \new_[9174]_ ;
  assign \new_[9181]_  = \new_[1064]_  | \new_[1065]_ ;
  assign \new_[9184]_  = \new_[1062]_  | \new_[1063]_ ;
  assign \new_[9185]_  = \new_[9184]_  | \new_[9181]_ ;
  assign \new_[9186]_  = \new_[9185]_  | \new_[9178]_ ;
  assign \new_[9187]_  = \new_[9186]_  | \new_[9171]_ ;
  assign \new_[9188]_  = \new_[9187]_  | \new_[9158]_ ;
  assign \new_[9189]_  = \new_[9188]_  | \new_[9129]_ ;
  assign \new_[9190]_  = \new_[9189]_  | \new_[9072]_ ;
  assign \new_[9194]_  = \new_[1059]_  | \new_[1060]_ ;
  assign \new_[9195]_  = \new_[1061]_  | \new_[9194]_ ;
  assign \new_[9198]_  = \new_[1057]_  | \new_[1058]_ ;
  assign \new_[9201]_  = \new_[1055]_  | \new_[1056]_ ;
  assign \new_[9202]_  = \new_[9201]_  | \new_[9198]_ ;
  assign \new_[9203]_  = \new_[9202]_  | \new_[9195]_ ;
  assign \new_[9207]_  = \new_[1052]_  | \new_[1053]_ ;
  assign \new_[9208]_  = \new_[1054]_  | \new_[9207]_ ;
  assign \new_[9211]_  = \new_[1050]_  | \new_[1051]_ ;
  assign \new_[9214]_  = \new_[1048]_  | \new_[1049]_ ;
  assign \new_[9215]_  = \new_[9214]_  | \new_[9211]_ ;
  assign \new_[9216]_  = \new_[9215]_  | \new_[9208]_ ;
  assign \new_[9217]_  = \new_[9216]_  | \new_[9203]_ ;
  assign \new_[9221]_  = \new_[1045]_  | \new_[1046]_ ;
  assign \new_[9222]_  = \new_[1047]_  | \new_[9221]_ ;
  assign \new_[9225]_  = \new_[1043]_  | \new_[1044]_ ;
  assign \new_[9228]_  = \new_[1041]_  | \new_[1042]_ ;
  assign \new_[9229]_  = \new_[9228]_  | \new_[9225]_ ;
  assign \new_[9230]_  = \new_[9229]_  | \new_[9222]_ ;
  assign \new_[9233]_  = \new_[1039]_  | \new_[1040]_ ;
  assign \new_[9236]_  = \new_[1037]_  | \new_[1038]_ ;
  assign \new_[9237]_  = \new_[9236]_  | \new_[9233]_ ;
  assign \new_[9240]_  = \new_[1035]_  | \new_[1036]_ ;
  assign \new_[9243]_  = \new_[1033]_  | \new_[1034]_ ;
  assign \new_[9244]_  = \new_[9243]_  | \new_[9240]_ ;
  assign \new_[9245]_  = \new_[9244]_  | \new_[9237]_ ;
  assign \new_[9246]_  = \new_[9245]_  | \new_[9230]_ ;
  assign \new_[9247]_  = \new_[9246]_  | \new_[9217]_ ;
  assign \new_[9251]_  = \new_[1030]_  | \new_[1031]_ ;
  assign \new_[9252]_  = \new_[1032]_  | \new_[9251]_ ;
  assign \new_[9255]_  = \new_[1028]_  | \new_[1029]_ ;
  assign \new_[9258]_  = \new_[1026]_  | \new_[1027]_ ;
  assign \new_[9259]_  = \new_[9258]_  | \new_[9255]_ ;
  assign \new_[9260]_  = \new_[9259]_  | \new_[9252]_ ;
  assign \new_[9263]_  = \new_[1024]_  | \new_[1025]_ ;
  assign \new_[9266]_  = \new_[1022]_  | \new_[1023]_ ;
  assign \new_[9267]_  = \new_[9266]_  | \new_[9263]_ ;
  assign \new_[9270]_  = \new_[1020]_  | \new_[1021]_ ;
  assign \new_[9273]_  = \new_[1018]_  | \new_[1019]_ ;
  assign \new_[9274]_  = \new_[9273]_  | \new_[9270]_ ;
  assign \new_[9275]_  = \new_[9274]_  | \new_[9267]_ ;
  assign \new_[9276]_  = \new_[9275]_  | \new_[9260]_ ;
  assign \new_[9280]_  = \new_[1015]_  | \new_[1016]_ ;
  assign \new_[9281]_  = \new_[1017]_  | \new_[9280]_ ;
  assign \new_[9284]_  = \new_[1013]_  | \new_[1014]_ ;
  assign \new_[9287]_  = \new_[1011]_  | \new_[1012]_ ;
  assign \new_[9288]_  = \new_[9287]_  | \new_[9284]_ ;
  assign \new_[9289]_  = \new_[9288]_  | \new_[9281]_ ;
  assign \new_[9292]_  = \new_[1009]_  | \new_[1010]_ ;
  assign \new_[9295]_  = \new_[1007]_  | \new_[1008]_ ;
  assign \new_[9296]_  = \new_[9295]_  | \new_[9292]_ ;
  assign \new_[9299]_  = \new_[1005]_  | \new_[1006]_ ;
  assign \new_[9302]_  = \new_[1003]_  | \new_[1004]_ ;
  assign \new_[9303]_  = \new_[9302]_  | \new_[9299]_ ;
  assign \new_[9304]_  = \new_[9303]_  | \new_[9296]_ ;
  assign \new_[9305]_  = \new_[9304]_  | \new_[9289]_ ;
  assign \new_[9306]_  = \new_[9305]_  | \new_[9276]_ ;
  assign \new_[9307]_  = \new_[9306]_  | \new_[9247]_ ;
  assign \new_[9311]_  = \new_[1000]_  | \new_[1001]_ ;
  assign \new_[9312]_  = \new_[1002]_  | \new_[9311]_ ;
  assign \new_[9315]_  = \new_[998]_  | \new_[999]_ ;
  assign \new_[9318]_  = \new_[996]_  | \new_[997]_ ;
  assign \new_[9319]_  = \new_[9318]_  | \new_[9315]_ ;
  assign \new_[9320]_  = \new_[9319]_  | \new_[9312]_ ;
  assign \new_[9324]_  = \new_[993]_  | \new_[994]_ ;
  assign \new_[9325]_  = \new_[995]_  | \new_[9324]_ ;
  assign \new_[9328]_  = \new_[991]_  | \new_[992]_ ;
  assign \new_[9331]_  = \new_[989]_  | \new_[990]_ ;
  assign \new_[9332]_  = \new_[9331]_  | \new_[9328]_ ;
  assign \new_[9333]_  = \new_[9332]_  | \new_[9325]_ ;
  assign \new_[9334]_  = \new_[9333]_  | \new_[9320]_ ;
  assign \new_[9338]_  = \new_[986]_  | \new_[987]_ ;
  assign \new_[9339]_  = \new_[988]_  | \new_[9338]_ ;
  assign \new_[9342]_  = \new_[984]_  | \new_[985]_ ;
  assign \new_[9345]_  = \new_[982]_  | \new_[983]_ ;
  assign \new_[9346]_  = \new_[9345]_  | \new_[9342]_ ;
  assign \new_[9347]_  = \new_[9346]_  | \new_[9339]_ ;
  assign \new_[9350]_  = \new_[980]_  | \new_[981]_ ;
  assign \new_[9353]_  = \new_[978]_  | \new_[979]_ ;
  assign \new_[9354]_  = \new_[9353]_  | \new_[9350]_ ;
  assign \new_[9357]_  = \new_[976]_  | \new_[977]_ ;
  assign \new_[9360]_  = \new_[974]_  | \new_[975]_ ;
  assign \new_[9361]_  = \new_[9360]_  | \new_[9357]_ ;
  assign \new_[9362]_  = \new_[9361]_  | \new_[9354]_ ;
  assign \new_[9363]_  = \new_[9362]_  | \new_[9347]_ ;
  assign \new_[9364]_  = \new_[9363]_  | \new_[9334]_ ;
  assign \new_[9368]_  = \new_[971]_  | \new_[972]_ ;
  assign \new_[9369]_  = \new_[973]_  | \new_[9368]_ ;
  assign \new_[9372]_  = \new_[969]_  | \new_[970]_ ;
  assign \new_[9375]_  = \new_[967]_  | \new_[968]_ ;
  assign \new_[9376]_  = \new_[9375]_  | \new_[9372]_ ;
  assign \new_[9377]_  = \new_[9376]_  | \new_[9369]_ ;
  assign \new_[9380]_  = \new_[965]_  | \new_[966]_ ;
  assign \new_[9383]_  = \new_[963]_  | \new_[964]_ ;
  assign \new_[9384]_  = \new_[9383]_  | \new_[9380]_ ;
  assign \new_[9387]_  = \new_[961]_  | \new_[962]_ ;
  assign \new_[9390]_  = \new_[959]_  | \new_[960]_ ;
  assign \new_[9391]_  = \new_[9390]_  | \new_[9387]_ ;
  assign \new_[9392]_  = \new_[9391]_  | \new_[9384]_ ;
  assign \new_[9393]_  = \new_[9392]_  | \new_[9377]_ ;
  assign \new_[9397]_  = \new_[956]_  | \new_[957]_ ;
  assign \new_[9398]_  = \new_[958]_  | \new_[9397]_ ;
  assign \new_[9401]_  = \new_[954]_  | \new_[955]_ ;
  assign \new_[9404]_  = \new_[952]_  | \new_[953]_ ;
  assign \new_[9405]_  = \new_[9404]_  | \new_[9401]_ ;
  assign \new_[9406]_  = \new_[9405]_  | \new_[9398]_ ;
  assign \new_[9409]_  = \new_[950]_  | \new_[951]_ ;
  assign \new_[9412]_  = \new_[948]_  | \new_[949]_ ;
  assign \new_[9413]_  = \new_[9412]_  | \new_[9409]_ ;
  assign \new_[9416]_  = \new_[946]_  | \new_[947]_ ;
  assign \new_[9419]_  = \new_[944]_  | \new_[945]_ ;
  assign \new_[9420]_  = \new_[9419]_  | \new_[9416]_ ;
  assign \new_[9421]_  = \new_[9420]_  | \new_[9413]_ ;
  assign \new_[9422]_  = \new_[9421]_  | \new_[9406]_ ;
  assign \new_[9423]_  = \new_[9422]_  | \new_[9393]_ ;
  assign \new_[9424]_  = \new_[9423]_  | \new_[9364]_ ;
  assign \new_[9425]_  = \new_[9424]_  | \new_[9307]_ ;
  assign \new_[9426]_  = \new_[9425]_  | \new_[9190]_ ;
  assign \new_[9427]_  = \new_[9426]_  | \new_[8955]_ ;
  assign \new_[9428]_  = \new_[9427]_  | \new_[8484]_ ;
  assign \new_[9432]_  = \new_[941]_  | \new_[942]_ ;
  assign \new_[9433]_  = \new_[943]_  | \new_[9432]_ ;
  assign \new_[9436]_  = \new_[939]_  | \new_[940]_ ;
  assign \new_[9439]_  = \new_[937]_  | \new_[938]_ ;
  assign \new_[9440]_  = \new_[9439]_  | \new_[9436]_ ;
  assign \new_[9441]_  = \new_[9440]_  | \new_[9433]_ ;
  assign \new_[9445]_  = \new_[934]_  | \new_[935]_ ;
  assign \new_[9446]_  = \new_[936]_  | \new_[9445]_ ;
  assign \new_[9449]_  = \new_[932]_  | \new_[933]_ ;
  assign \new_[9452]_  = \new_[930]_  | \new_[931]_ ;
  assign \new_[9453]_  = \new_[9452]_  | \new_[9449]_ ;
  assign \new_[9454]_  = \new_[9453]_  | \new_[9446]_ ;
  assign \new_[9455]_  = \new_[9454]_  | \new_[9441]_ ;
  assign \new_[9459]_  = \new_[927]_  | \new_[928]_ ;
  assign \new_[9460]_  = \new_[929]_  | \new_[9459]_ ;
  assign \new_[9463]_  = \new_[925]_  | \new_[926]_ ;
  assign \new_[9466]_  = \new_[923]_  | \new_[924]_ ;
  assign \new_[9467]_  = \new_[9466]_  | \new_[9463]_ ;
  assign \new_[9468]_  = \new_[9467]_  | \new_[9460]_ ;
  assign \new_[9471]_  = \new_[921]_  | \new_[922]_ ;
  assign \new_[9474]_  = \new_[919]_  | \new_[920]_ ;
  assign \new_[9475]_  = \new_[9474]_  | \new_[9471]_ ;
  assign \new_[9478]_  = \new_[917]_  | \new_[918]_ ;
  assign \new_[9481]_  = \new_[915]_  | \new_[916]_ ;
  assign \new_[9482]_  = \new_[9481]_  | \new_[9478]_ ;
  assign \new_[9483]_  = \new_[9482]_  | \new_[9475]_ ;
  assign \new_[9484]_  = \new_[9483]_  | \new_[9468]_ ;
  assign \new_[9485]_  = \new_[9484]_  | \new_[9455]_ ;
  assign \new_[9489]_  = \new_[912]_  | \new_[913]_ ;
  assign \new_[9490]_  = \new_[914]_  | \new_[9489]_ ;
  assign \new_[9493]_  = \new_[910]_  | \new_[911]_ ;
  assign \new_[9496]_  = \new_[908]_  | \new_[909]_ ;
  assign \new_[9497]_  = \new_[9496]_  | \new_[9493]_ ;
  assign \new_[9498]_  = \new_[9497]_  | \new_[9490]_ ;
  assign \new_[9502]_  = \new_[905]_  | \new_[906]_ ;
  assign \new_[9503]_  = \new_[907]_  | \new_[9502]_ ;
  assign \new_[9506]_  = \new_[903]_  | \new_[904]_ ;
  assign \new_[9509]_  = \new_[901]_  | \new_[902]_ ;
  assign \new_[9510]_  = \new_[9509]_  | \new_[9506]_ ;
  assign \new_[9511]_  = \new_[9510]_  | \new_[9503]_ ;
  assign \new_[9512]_  = \new_[9511]_  | \new_[9498]_ ;
  assign \new_[9516]_  = \new_[898]_  | \new_[899]_ ;
  assign \new_[9517]_  = \new_[900]_  | \new_[9516]_ ;
  assign \new_[9520]_  = \new_[896]_  | \new_[897]_ ;
  assign \new_[9523]_  = \new_[894]_  | \new_[895]_ ;
  assign \new_[9524]_  = \new_[9523]_  | \new_[9520]_ ;
  assign \new_[9525]_  = \new_[9524]_  | \new_[9517]_ ;
  assign \new_[9528]_  = \new_[892]_  | \new_[893]_ ;
  assign \new_[9531]_  = \new_[890]_  | \new_[891]_ ;
  assign \new_[9532]_  = \new_[9531]_  | \new_[9528]_ ;
  assign \new_[9535]_  = \new_[888]_  | \new_[889]_ ;
  assign \new_[9538]_  = \new_[886]_  | \new_[887]_ ;
  assign \new_[9539]_  = \new_[9538]_  | \new_[9535]_ ;
  assign \new_[9540]_  = \new_[9539]_  | \new_[9532]_ ;
  assign \new_[9541]_  = \new_[9540]_  | \new_[9525]_ ;
  assign \new_[9542]_  = \new_[9541]_  | \new_[9512]_ ;
  assign \new_[9543]_  = \new_[9542]_  | \new_[9485]_ ;
  assign \new_[9547]_  = \new_[883]_  | \new_[884]_ ;
  assign \new_[9548]_  = \new_[885]_  | \new_[9547]_ ;
  assign \new_[9551]_  = \new_[881]_  | \new_[882]_ ;
  assign \new_[9554]_  = \new_[879]_  | \new_[880]_ ;
  assign \new_[9555]_  = \new_[9554]_  | \new_[9551]_ ;
  assign \new_[9556]_  = \new_[9555]_  | \new_[9548]_ ;
  assign \new_[9560]_  = \new_[876]_  | \new_[877]_ ;
  assign \new_[9561]_  = \new_[878]_  | \new_[9560]_ ;
  assign \new_[9564]_  = \new_[874]_  | \new_[875]_ ;
  assign \new_[9567]_  = \new_[872]_  | \new_[873]_ ;
  assign \new_[9568]_  = \new_[9567]_  | \new_[9564]_ ;
  assign \new_[9569]_  = \new_[9568]_  | \new_[9561]_ ;
  assign \new_[9570]_  = \new_[9569]_  | \new_[9556]_ ;
  assign \new_[9574]_  = \new_[869]_  | \new_[870]_ ;
  assign \new_[9575]_  = \new_[871]_  | \new_[9574]_ ;
  assign \new_[9578]_  = \new_[867]_  | \new_[868]_ ;
  assign \new_[9581]_  = \new_[865]_  | \new_[866]_ ;
  assign \new_[9582]_  = \new_[9581]_  | \new_[9578]_ ;
  assign \new_[9583]_  = \new_[9582]_  | \new_[9575]_ ;
  assign \new_[9586]_  = \new_[863]_  | \new_[864]_ ;
  assign \new_[9589]_  = \new_[861]_  | \new_[862]_ ;
  assign \new_[9590]_  = \new_[9589]_  | \new_[9586]_ ;
  assign \new_[9593]_  = \new_[859]_  | \new_[860]_ ;
  assign \new_[9596]_  = \new_[857]_  | \new_[858]_ ;
  assign \new_[9597]_  = \new_[9596]_  | \new_[9593]_ ;
  assign \new_[9598]_  = \new_[9597]_  | \new_[9590]_ ;
  assign \new_[9599]_  = \new_[9598]_  | \new_[9583]_ ;
  assign \new_[9600]_  = \new_[9599]_  | \new_[9570]_ ;
  assign \new_[9604]_  = \new_[854]_  | \new_[855]_ ;
  assign \new_[9605]_  = \new_[856]_  | \new_[9604]_ ;
  assign \new_[9608]_  = \new_[852]_  | \new_[853]_ ;
  assign \new_[9611]_  = \new_[850]_  | \new_[851]_ ;
  assign \new_[9612]_  = \new_[9611]_  | \new_[9608]_ ;
  assign \new_[9613]_  = \new_[9612]_  | \new_[9605]_ ;
  assign \new_[9616]_  = \new_[848]_  | \new_[849]_ ;
  assign \new_[9619]_  = \new_[846]_  | \new_[847]_ ;
  assign \new_[9620]_  = \new_[9619]_  | \new_[9616]_ ;
  assign \new_[9623]_  = \new_[844]_  | \new_[845]_ ;
  assign \new_[9626]_  = \new_[842]_  | \new_[843]_ ;
  assign \new_[9627]_  = \new_[9626]_  | \new_[9623]_ ;
  assign \new_[9628]_  = \new_[9627]_  | \new_[9620]_ ;
  assign \new_[9629]_  = \new_[9628]_  | \new_[9613]_ ;
  assign \new_[9633]_  = \new_[839]_  | \new_[840]_ ;
  assign \new_[9634]_  = \new_[841]_  | \new_[9633]_ ;
  assign \new_[9637]_  = \new_[837]_  | \new_[838]_ ;
  assign \new_[9640]_  = \new_[835]_  | \new_[836]_ ;
  assign \new_[9641]_  = \new_[9640]_  | \new_[9637]_ ;
  assign \new_[9642]_  = \new_[9641]_  | \new_[9634]_ ;
  assign \new_[9645]_  = \new_[833]_  | \new_[834]_ ;
  assign \new_[9648]_  = \new_[831]_  | \new_[832]_ ;
  assign \new_[9649]_  = \new_[9648]_  | \new_[9645]_ ;
  assign \new_[9652]_  = \new_[829]_  | \new_[830]_ ;
  assign \new_[9655]_  = \new_[827]_  | \new_[828]_ ;
  assign \new_[9656]_  = \new_[9655]_  | \new_[9652]_ ;
  assign \new_[9657]_  = \new_[9656]_  | \new_[9649]_ ;
  assign \new_[9658]_  = \new_[9657]_  | \new_[9642]_ ;
  assign \new_[9659]_  = \new_[9658]_  | \new_[9629]_ ;
  assign \new_[9660]_  = \new_[9659]_  | \new_[9600]_ ;
  assign \new_[9661]_  = \new_[9660]_  | \new_[9543]_ ;
  assign \new_[9665]_  = \new_[824]_  | \new_[825]_ ;
  assign \new_[9666]_  = \new_[826]_  | \new_[9665]_ ;
  assign \new_[9669]_  = \new_[822]_  | \new_[823]_ ;
  assign \new_[9672]_  = \new_[820]_  | \new_[821]_ ;
  assign \new_[9673]_  = \new_[9672]_  | \new_[9669]_ ;
  assign \new_[9674]_  = \new_[9673]_  | \new_[9666]_ ;
  assign \new_[9678]_  = \new_[817]_  | \new_[818]_ ;
  assign \new_[9679]_  = \new_[819]_  | \new_[9678]_ ;
  assign \new_[9682]_  = \new_[815]_  | \new_[816]_ ;
  assign \new_[9685]_  = \new_[813]_  | \new_[814]_ ;
  assign \new_[9686]_  = \new_[9685]_  | \new_[9682]_ ;
  assign \new_[9687]_  = \new_[9686]_  | \new_[9679]_ ;
  assign \new_[9688]_  = \new_[9687]_  | \new_[9674]_ ;
  assign \new_[9692]_  = \new_[810]_  | \new_[811]_ ;
  assign \new_[9693]_  = \new_[812]_  | \new_[9692]_ ;
  assign \new_[9696]_  = \new_[808]_  | \new_[809]_ ;
  assign \new_[9699]_  = \new_[806]_  | \new_[807]_ ;
  assign \new_[9700]_  = \new_[9699]_  | \new_[9696]_ ;
  assign \new_[9701]_  = \new_[9700]_  | \new_[9693]_ ;
  assign \new_[9704]_  = \new_[804]_  | \new_[805]_ ;
  assign \new_[9707]_  = \new_[802]_  | \new_[803]_ ;
  assign \new_[9708]_  = \new_[9707]_  | \new_[9704]_ ;
  assign \new_[9711]_  = \new_[800]_  | \new_[801]_ ;
  assign \new_[9714]_  = \new_[798]_  | \new_[799]_ ;
  assign \new_[9715]_  = \new_[9714]_  | \new_[9711]_ ;
  assign \new_[9716]_  = \new_[9715]_  | \new_[9708]_ ;
  assign \new_[9717]_  = \new_[9716]_  | \new_[9701]_ ;
  assign \new_[9718]_  = \new_[9717]_  | \new_[9688]_ ;
  assign \new_[9722]_  = \new_[795]_  | \new_[796]_ ;
  assign \new_[9723]_  = \new_[797]_  | \new_[9722]_ ;
  assign \new_[9726]_  = \new_[793]_  | \new_[794]_ ;
  assign \new_[9729]_  = \new_[791]_  | \new_[792]_ ;
  assign \new_[9730]_  = \new_[9729]_  | \new_[9726]_ ;
  assign \new_[9731]_  = \new_[9730]_  | \new_[9723]_ ;
  assign \new_[9734]_  = \new_[789]_  | \new_[790]_ ;
  assign \new_[9737]_  = \new_[787]_  | \new_[788]_ ;
  assign \new_[9738]_  = \new_[9737]_  | \new_[9734]_ ;
  assign \new_[9741]_  = \new_[785]_  | \new_[786]_ ;
  assign \new_[9744]_  = \new_[783]_  | \new_[784]_ ;
  assign \new_[9745]_  = \new_[9744]_  | \new_[9741]_ ;
  assign \new_[9746]_  = \new_[9745]_  | \new_[9738]_ ;
  assign \new_[9747]_  = \new_[9746]_  | \new_[9731]_ ;
  assign \new_[9751]_  = \new_[780]_  | \new_[781]_ ;
  assign \new_[9752]_  = \new_[782]_  | \new_[9751]_ ;
  assign \new_[9755]_  = \new_[778]_  | \new_[779]_ ;
  assign \new_[9758]_  = \new_[776]_  | \new_[777]_ ;
  assign \new_[9759]_  = \new_[9758]_  | \new_[9755]_ ;
  assign \new_[9760]_  = \new_[9759]_  | \new_[9752]_ ;
  assign \new_[9763]_  = \new_[774]_  | \new_[775]_ ;
  assign \new_[9766]_  = \new_[772]_  | \new_[773]_ ;
  assign \new_[9767]_  = \new_[9766]_  | \new_[9763]_ ;
  assign \new_[9770]_  = \new_[770]_  | \new_[771]_ ;
  assign \new_[9773]_  = \new_[768]_  | \new_[769]_ ;
  assign \new_[9774]_  = \new_[9773]_  | \new_[9770]_ ;
  assign \new_[9775]_  = \new_[9774]_  | \new_[9767]_ ;
  assign \new_[9776]_  = \new_[9775]_  | \new_[9760]_ ;
  assign \new_[9777]_  = \new_[9776]_  | \new_[9747]_ ;
  assign \new_[9778]_  = \new_[9777]_  | \new_[9718]_ ;
  assign \new_[9782]_  = \new_[765]_  | \new_[766]_ ;
  assign \new_[9783]_  = \new_[767]_  | \new_[9782]_ ;
  assign \new_[9786]_  = \new_[763]_  | \new_[764]_ ;
  assign \new_[9789]_  = \new_[761]_  | \new_[762]_ ;
  assign \new_[9790]_  = \new_[9789]_  | \new_[9786]_ ;
  assign \new_[9791]_  = \new_[9790]_  | \new_[9783]_ ;
  assign \new_[9795]_  = \new_[758]_  | \new_[759]_ ;
  assign \new_[9796]_  = \new_[760]_  | \new_[9795]_ ;
  assign \new_[9799]_  = \new_[756]_  | \new_[757]_ ;
  assign \new_[9802]_  = \new_[754]_  | \new_[755]_ ;
  assign \new_[9803]_  = \new_[9802]_  | \new_[9799]_ ;
  assign \new_[9804]_  = \new_[9803]_  | \new_[9796]_ ;
  assign \new_[9805]_  = \new_[9804]_  | \new_[9791]_ ;
  assign \new_[9809]_  = \new_[751]_  | \new_[752]_ ;
  assign \new_[9810]_  = \new_[753]_  | \new_[9809]_ ;
  assign \new_[9813]_  = \new_[749]_  | \new_[750]_ ;
  assign \new_[9816]_  = \new_[747]_  | \new_[748]_ ;
  assign \new_[9817]_  = \new_[9816]_  | \new_[9813]_ ;
  assign \new_[9818]_  = \new_[9817]_  | \new_[9810]_ ;
  assign \new_[9821]_  = \new_[745]_  | \new_[746]_ ;
  assign \new_[9824]_  = \new_[743]_  | \new_[744]_ ;
  assign \new_[9825]_  = \new_[9824]_  | \new_[9821]_ ;
  assign \new_[9828]_  = \new_[741]_  | \new_[742]_ ;
  assign \new_[9831]_  = \new_[739]_  | \new_[740]_ ;
  assign \new_[9832]_  = \new_[9831]_  | \new_[9828]_ ;
  assign \new_[9833]_  = \new_[9832]_  | \new_[9825]_ ;
  assign \new_[9834]_  = \new_[9833]_  | \new_[9818]_ ;
  assign \new_[9835]_  = \new_[9834]_  | \new_[9805]_ ;
  assign \new_[9839]_  = \new_[736]_  | \new_[737]_ ;
  assign \new_[9840]_  = \new_[738]_  | \new_[9839]_ ;
  assign \new_[9843]_  = \new_[734]_  | \new_[735]_ ;
  assign \new_[9846]_  = \new_[732]_  | \new_[733]_ ;
  assign \new_[9847]_  = \new_[9846]_  | \new_[9843]_ ;
  assign \new_[9848]_  = \new_[9847]_  | \new_[9840]_ ;
  assign \new_[9851]_  = \new_[730]_  | \new_[731]_ ;
  assign \new_[9854]_  = \new_[728]_  | \new_[729]_ ;
  assign \new_[9855]_  = \new_[9854]_  | \new_[9851]_ ;
  assign \new_[9858]_  = \new_[726]_  | \new_[727]_ ;
  assign \new_[9861]_  = \new_[724]_  | \new_[725]_ ;
  assign \new_[9862]_  = \new_[9861]_  | \new_[9858]_ ;
  assign \new_[9863]_  = \new_[9862]_  | \new_[9855]_ ;
  assign \new_[9864]_  = \new_[9863]_  | \new_[9848]_ ;
  assign \new_[9868]_  = \new_[721]_  | \new_[722]_ ;
  assign \new_[9869]_  = \new_[723]_  | \new_[9868]_ ;
  assign \new_[9872]_  = \new_[719]_  | \new_[720]_ ;
  assign \new_[9875]_  = \new_[717]_  | \new_[718]_ ;
  assign \new_[9876]_  = \new_[9875]_  | \new_[9872]_ ;
  assign \new_[9877]_  = \new_[9876]_  | \new_[9869]_ ;
  assign \new_[9880]_  = \new_[715]_  | \new_[716]_ ;
  assign \new_[9883]_  = \new_[713]_  | \new_[714]_ ;
  assign \new_[9884]_  = \new_[9883]_  | \new_[9880]_ ;
  assign \new_[9887]_  = \new_[711]_  | \new_[712]_ ;
  assign \new_[9890]_  = \new_[709]_  | \new_[710]_ ;
  assign \new_[9891]_  = \new_[9890]_  | \new_[9887]_ ;
  assign \new_[9892]_  = \new_[9891]_  | \new_[9884]_ ;
  assign \new_[9893]_  = \new_[9892]_  | \new_[9877]_ ;
  assign \new_[9894]_  = \new_[9893]_  | \new_[9864]_ ;
  assign \new_[9895]_  = \new_[9894]_  | \new_[9835]_ ;
  assign \new_[9896]_  = \new_[9895]_  | \new_[9778]_ ;
  assign \new_[9897]_  = \new_[9896]_  | \new_[9661]_ ;
  assign \new_[9901]_  = \new_[706]_  | \new_[707]_ ;
  assign \new_[9902]_  = \new_[708]_  | \new_[9901]_ ;
  assign \new_[9905]_  = \new_[704]_  | \new_[705]_ ;
  assign \new_[9908]_  = \new_[702]_  | \new_[703]_ ;
  assign \new_[9909]_  = \new_[9908]_  | \new_[9905]_ ;
  assign \new_[9910]_  = \new_[9909]_  | \new_[9902]_ ;
  assign \new_[9914]_  = \new_[699]_  | \new_[700]_ ;
  assign \new_[9915]_  = \new_[701]_  | \new_[9914]_ ;
  assign \new_[9918]_  = \new_[697]_  | \new_[698]_ ;
  assign \new_[9921]_  = \new_[695]_  | \new_[696]_ ;
  assign \new_[9922]_  = \new_[9921]_  | \new_[9918]_ ;
  assign \new_[9923]_  = \new_[9922]_  | \new_[9915]_ ;
  assign \new_[9924]_  = \new_[9923]_  | \new_[9910]_ ;
  assign \new_[9928]_  = \new_[692]_  | \new_[693]_ ;
  assign \new_[9929]_  = \new_[694]_  | \new_[9928]_ ;
  assign \new_[9932]_  = \new_[690]_  | \new_[691]_ ;
  assign \new_[9935]_  = \new_[688]_  | \new_[689]_ ;
  assign \new_[9936]_  = \new_[9935]_  | \new_[9932]_ ;
  assign \new_[9937]_  = \new_[9936]_  | \new_[9929]_ ;
  assign \new_[9940]_  = \new_[686]_  | \new_[687]_ ;
  assign \new_[9943]_  = \new_[684]_  | \new_[685]_ ;
  assign \new_[9944]_  = \new_[9943]_  | \new_[9940]_ ;
  assign \new_[9947]_  = \new_[682]_  | \new_[683]_ ;
  assign \new_[9950]_  = \new_[680]_  | \new_[681]_ ;
  assign \new_[9951]_  = \new_[9950]_  | \new_[9947]_ ;
  assign \new_[9952]_  = \new_[9951]_  | \new_[9944]_ ;
  assign \new_[9953]_  = \new_[9952]_  | \new_[9937]_ ;
  assign \new_[9954]_  = \new_[9953]_  | \new_[9924]_ ;
  assign \new_[9958]_  = \new_[677]_  | \new_[678]_ ;
  assign \new_[9959]_  = \new_[679]_  | \new_[9958]_ ;
  assign \new_[9962]_  = \new_[675]_  | \new_[676]_ ;
  assign \new_[9965]_  = \new_[673]_  | \new_[674]_ ;
  assign \new_[9966]_  = \new_[9965]_  | \new_[9962]_ ;
  assign \new_[9967]_  = \new_[9966]_  | \new_[9959]_ ;
  assign \new_[9970]_  = \new_[671]_  | \new_[672]_ ;
  assign \new_[9973]_  = \new_[669]_  | \new_[670]_ ;
  assign \new_[9974]_  = \new_[9973]_  | \new_[9970]_ ;
  assign \new_[9977]_  = \new_[667]_  | \new_[668]_ ;
  assign \new_[9980]_  = \new_[665]_  | \new_[666]_ ;
  assign \new_[9981]_  = \new_[9980]_  | \new_[9977]_ ;
  assign \new_[9982]_  = \new_[9981]_  | \new_[9974]_ ;
  assign \new_[9983]_  = \new_[9982]_  | \new_[9967]_ ;
  assign \new_[9987]_  = \new_[662]_  | \new_[663]_ ;
  assign \new_[9988]_  = \new_[664]_  | \new_[9987]_ ;
  assign \new_[9991]_  = \new_[660]_  | \new_[661]_ ;
  assign \new_[9994]_  = \new_[658]_  | \new_[659]_ ;
  assign \new_[9995]_  = \new_[9994]_  | \new_[9991]_ ;
  assign \new_[9996]_  = \new_[9995]_  | \new_[9988]_ ;
  assign \new_[9999]_  = \new_[656]_  | \new_[657]_ ;
  assign \new_[10002]_  = \new_[654]_  | \new_[655]_ ;
  assign \new_[10003]_  = \new_[10002]_  | \new_[9999]_ ;
  assign \new_[10006]_  = \new_[652]_  | \new_[653]_ ;
  assign \new_[10009]_  = \new_[650]_  | \new_[651]_ ;
  assign \new_[10010]_  = \new_[10009]_  | \new_[10006]_ ;
  assign \new_[10011]_  = \new_[10010]_  | \new_[10003]_ ;
  assign \new_[10012]_  = \new_[10011]_  | \new_[9996]_ ;
  assign \new_[10013]_  = \new_[10012]_  | \new_[9983]_ ;
  assign \new_[10014]_  = \new_[10013]_  | \new_[9954]_ ;
  assign \new_[10018]_  = \new_[647]_  | \new_[648]_ ;
  assign \new_[10019]_  = \new_[649]_  | \new_[10018]_ ;
  assign \new_[10022]_  = \new_[645]_  | \new_[646]_ ;
  assign \new_[10025]_  = \new_[643]_  | \new_[644]_ ;
  assign \new_[10026]_  = \new_[10025]_  | \new_[10022]_ ;
  assign \new_[10027]_  = \new_[10026]_  | \new_[10019]_ ;
  assign \new_[10031]_  = \new_[640]_  | \new_[641]_ ;
  assign \new_[10032]_  = \new_[642]_  | \new_[10031]_ ;
  assign \new_[10035]_  = \new_[638]_  | \new_[639]_ ;
  assign \new_[10038]_  = \new_[636]_  | \new_[637]_ ;
  assign \new_[10039]_  = \new_[10038]_  | \new_[10035]_ ;
  assign \new_[10040]_  = \new_[10039]_  | \new_[10032]_ ;
  assign \new_[10041]_  = \new_[10040]_  | \new_[10027]_ ;
  assign \new_[10045]_  = \new_[633]_  | \new_[634]_ ;
  assign \new_[10046]_  = \new_[635]_  | \new_[10045]_ ;
  assign \new_[10049]_  = \new_[631]_  | \new_[632]_ ;
  assign \new_[10052]_  = \new_[629]_  | \new_[630]_ ;
  assign \new_[10053]_  = \new_[10052]_  | \new_[10049]_ ;
  assign \new_[10054]_  = \new_[10053]_  | \new_[10046]_ ;
  assign \new_[10057]_  = \new_[627]_  | \new_[628]_ ;
  assign \new_[10060]_  = \new_[625]_  | \new_[626]_ ;
  assign \new_[10061]_  = \new_[10060]_  | \new_[10057]_ ;
  assign \new_[10064]_  = \new_[623]_  | \new_[624]_ ;
  assign \new_[10067]_  = \new_[621]_  | \new_[622]_ ;
  assign \new_[10068]_  = \new_[10067]_  | \new_[10064]_ ;
  assign \new_[10069]_  = \new_[10068]_  | \new_[10061]_ ;
  assign \new_[10070]_  = \new_[10069]_  | \new_[10054]_ ;
  assign \new_[10071]_  = \new_[10070]_  | \new_[10041]_ ;
  assign \new_[10075]_  = \new_[618]_  | \new_[619]_ ;
  assign \new_[10076]_  = \new_[620]_  | \new_[10075]_ ;
  assign \new_[10079]_  = \new_[616]_  | \new_[617]_ ;
  assign \new_[10082]_  = \new_[614]_  | \new_[615]_ ;
  assign \new_[10083]_  = \new_[10082]_  | \new_[10079]_ ;
  assign \new_[10084]_  = \new_[10083]_  | \new_[10076]_ ;
  assign \new_[10087]_  = \new_[612]_  | \new_[613]_ ;
  assign \new_[10090]_  = \new_[610]_  | \new_[611]_ ;
  assign \new_[10091]_  = \new_[10090]_  | \new_[10087]_ ;
  assign \new_[10094]_  = \new_[608]_  | \new_[609]_ ;
  assign \new_[10097]_  = \new_[606]_  | \new_[607]_ ;
  assign \new_[10098]_  = \new_[10097]_  | \new_[10094]_ ;
  assign \new_[10099]_  = \new_[10098]_  | \new_[10091]_ ;
  assign \new_[10100]_  = \new_[10099]_  | \new_[10084]_ ;
  assign \new_[10104]_  = \new_[603]_  | \new_[604]_ ;
  assign \new_[10105]_  = \new_[605]_  | \new_[10104]_ ;
  assign \new_[10108]_  = \new_[601]_  | \new_[602]_ ;
  assign \new_[10111]_  = \new_[599]_  | \new_[600]_ ;
  assign \new_[10112]_  = \new_[10111]_  | \new_[10108]_ ;
  assign \new_[10113]_  = \new_[10112]_  | \new_[10105]_ ;
  assign \new_[10116]_  = \new_[597]_  | \new_[598]_ ;
  assign \new_[10119]_  = \new_[595]_  | \new_[596]_ ;
  assign \new_[10120]_  = \new_[10119]_  | \new_[10116]_ ;
  assign \new_[10123]_  = \new_[593]_  | \new_[594]_ ;
  assign \new_[10126]_  = \new_[591]_  | \new_[592]_ ;
  assign \new_[10127]_  = \new_[10126]_  | \new_[10123]_ ;
  assign \new_[10128]_  = \new_[10127]_  | \new_[10120]_ ;
  assign \new_[10129]_  = \new_[10128]_  | \new_[10113]_ ;
  assign \new_[10130]_  = \new_[10129]_  | \new_[10100]_ ;
  assign \new_[10131]_  = \new_[10130]_  | \new_[10071]_ ;
  assign \new_[10132]_  = \new_[10131]_  | \new_[10014]_ ;
  assign \new_[10136]_  = \new_[588]_  | \new_[589]_ ;
  assign \new_[10137]_  = \new_[590]_  | \new_[10136]_ ;
  assign \new_[10140]_  = \new_[586]_  | \new_[587]_ ;
  assign \new_[10143]_  = \new_[584]_  | \new_[585]_ ;
  assign \new_[10144]_  = \new_[10143]_  | \new_[10140]_ ;
  assign \new_[10145]_  = \new_[10144]_  | \new_[10137]_ ;
  assign \new_[10149]_  = \new_[581]_  | \new_[582]_ ;
  assign \new_[10150]_  = \new_[583]_  | \new_[10149]_ ;
  assign \new_[10153]_  = \new_[579]_  | \new_[580]_ ;
  assign \new_[10156]_  = \new_[577]_  | \new_[578]_ ;
  assign \new_[10157]_  = \new_[10156]_  | \new_[10153]_ ;
  assign \new_[10158]_  = \new_[10157]_  | \new_[10150]_ ;
  assign \new_[10159]_  = \new_[10158]_  | \new_[10145]_ ;
  assign \new_[10163]_  = \new_[574]_  | \new_[575]_ ;
  assign \new_[10164]_  = \new_[576]_  | \new_[10163]_ ;
  assign \new_[10167]_  = \new_[572]_  | \new_[573]_ ;
  assign \new_[10170]_  = \new_[570]_  | \new_[571]_ ;
  assign \new_[10171]_  = \new_[10170]_  | \new_[10167]_ ;
  assign \new_[10172]_  = \new_[10171]_  | \new_[10164]_ ;
  assign \new_[10175]_  = \new_[568]_  | \new_[569]_ ;
  assign \new_[10178]_  = \new_[566]_  | \new_[567]_ ;
  assign \new_[10179]_  = \new_[10178]_  | \new_[10175]_ ;
  assign \new_[10182]_  = \new_[564]_  | \new_[565]_ ;
  assign \new_[10185]_  = \new_[562]_  | \new_[563]_ ;
  assign \new_[10186]_  = \new_[10185]_  | \new_[10182]_ ;
  assign \new_[10187]_  = \new_[10186]_  | \new_[10179]_ ;
  assign \new_[10188]_  = \new_[10187]_  | \new_[10172]_ ;
  assign \new_[10189]_  = \new_[10188]_  | \new_[10159]_ ;
  assign \new_[10193]_  = \new_[559]_  | \new_[560]_ ;
  assign \new_[10194]_  = \new_[561]_  | \new_[10193]_ ;
  assign \new_[10197]_  = \new_[557]_  | \new_[558]_ ;
  assign \new_[10200]_  = \new_[555]_  | \new_[556]_ ;
  assign \new_[10201]_  = \new_[10200]_  | \new_[10197]_ ;
  assign \new_[10202]_  = \new_[10201]_  | \new_[10194]_ ;
  assign \new_[10205]_  = \new_[553]_  | \new_[554]_ ;
  assign \new_[10208]_  = \new_[551]_  | \new_[552]_ ;
  assign \new_[10209]_  = \new_[10208]_  | \new_[10205]_ ;
  assign \new_[10212]_  = \new_[549]_  | \new_[550]_ ;
  assign \new_[10215]_  = \new_[547]_  | \new_[548]_ ;
  assign \new_[10216]_  = \new_[10215]_  | \new_[10212]_ ;
  assign \new_[10217]_  = \new_[10216]_  | \new_[10209]_ ;
  assign \new_[10218]_  = \new_[10217]_  | \new_[10202]_ ;
  assign \new_[10222]_  = \new_[544]_  | \new_[545]_ ;
  assign \new_[10223]_  = \new_[546]_  | \new_[10222]_ ;
  assign \new_[10226]_  = \new_[542]_  | \new_[543]_ ;
  assign \new_[10229]_  = \new_[540]_  | \new_[541]_ ;
  assign \new_[10230]_  = \new_[10229]_  | \new_[10226]_ ;
  assign \new_[10231]_  = \new_[10230]_  | \new_[10223]_ ;
  assign \new_[10234]_  = \new_[538]_  | \new_[539]_ ;
  assign \new_[10237]_  = \new_[536]_  | \new_[537]_ ;
  assign \new_[10238]_  = \new_[10237]_  | \new_[10234]_ ;
  assign \new_[10241]_  = \new_[534]_  | \new_[535]_ ;
  assign \new_[10244]_  = \new_[532]_  | \new_[533]_ ;
  assign \new_[10245]_  = \new_[10244]_  | \new_[10241]_ ;
  assign \new_[10246]_  = \new_[10245]_  | \new_[10238]_ ;
  assign \new_[10247]_  = \new_[10246]_  | \new_[10231]_ ;
  assign \new_[10248]_  = \new_[10247]_  | \new_[10218]_ ;
  assign \new_[10249]_  = \new_[10248]_  | \new_[10189]_ ;
  assign \new_[10253]_  = \new_[529]_  | \new_[530]_ ;
  assign \new_[10254]_  = \new_[531]_  | \new_[10253]_ ;
  assign \new_[10257]_  = \new_[527]_  | \new_[528]_ ;
  assign \new_[10260]_  = \new_[525]_  | \new_[526]_ ;
  assign \new_[10261]_  = \new_[10260]_  | \new_[10257]_ ;
  assign \new_[10262]_  = \new_[10261]_  | \new_[10254]_ ;
  assign \new_[10266]_  = \new_[522]_  | \new_[523]_ ;
  assign \new_[10267]_  = \new_[524]_  | \new_[10266]_ ;
  assign \new_[10270]_  = \new_[520]_  | \new_[521]_ ;
  assign \new_[10273]_  = \new_[518]_  | \new_[519]_ ;
  assign \new_[10274]_  = \new_[10273]_  | \new_[10270]_ ;
  assign \new_[10275]_  = \new_[10274]_  | \new_[10267]_ ;
  assign \new_[10276]_  = \new_[10275]_  | \new_[10262]_ ;
  assign \new_[10280]_  = \new_[515]_  | \new_[516]_ ;
  assign \new_[10281]_  = \new_[517]_  | \new_[10280]_ ;
  assign \new_[10284]_  = \new_[513]_  | \new_[514]_ ;
  assign \new_[10287]_  = \new_[511]_  | \new_[512]_ ;
  assign \new_[10288]_  = \new_[10287]_  | \new_[10284]_ ;
  assign \new_[10289]_  = \new_[10288]_  | \new_[10281]_ ;
  assign \new_[10292]_  = \new_[509]_  | \new_[510]_ ;
  assign \new_[10295]_  = \new_[507]_  | \new_[508]_ ;
  assign \new_[10296]_  = \new_[10295]_  | \new_[10292]_ ;
  assign \new_[10299]_  = \new_[505]_  | \new_[506]_ ;
  assign \new_[10302]_  = \new_[503]_  | \new_[504]_ ;
  assign \new_[10303]_  = \new_[10302]_  | \new_[10299]_ ;
  assign \new_[10304]_  = \new_[10303]_  | \new_[10296]_ ;
  assign \new_[10305]_  = \new_[10304]_  | \new_[10289]_ ;
  assign \new_[10306]_  = \new_[10305]_  | \new_[10276]_ ;
  assign \new_[10310]_  = \new_[500]_  | \new_[501]_ ;
  assign \new_[10311]_  = \new_[502]_  | \new_[10310]_ ;
  assign \new_[10314]_  = \new_[498]_  | \new_[499]_ ;
  assign \new_[10317]_  = \new_[496]_  | \new_[497]_ ;
  assign \new_[10318]_  = \new_[10317]_  | \new_[10314]_ ;
  assign \new_[10319]_  = \new_[10318]_  | \new_[10311]_ ;
  assign \new_[10322]_  = \new_[494]_  | \new_[495]_ ;
  assign \new_[10325]_  = \new_[492]_  | \new_[493]_ ;
  assign \new_[10326]_  = \new_[10325]_  | \new_[10322]_ ;
  assign \new_[10329]_  = \new_[490]_  | \new_[491]_ ;
  assign \new_[10332]_  = \new_[488]_  | \new_[489]_ ;
  assign \new_[10333]_  = \new_[10332]_  | \new_[10329]_ ;
  assign \new_[10334]_  = \new_[10333]_  | \new_[10326]_ ;
  assign \new_[10335]_  = \new_[10334]_  | \new_[10319]_ ;
  assign \new_[10339]_  = \new_[485]_  | \new_[486]_ ;
  assign \new_[10340]_  = \new_[487]_  | \new_[10339]_ ;
  assign \new_[10343]_  = \new_[483]_  | \new_[484]_ ;
  assign \new_[10346]_  = \new_[481]_  | \new_[482]_ ;
  assign \new_[10347]_  = \new_[10346]_  | \new_[10343]_ ;
  assign \new_[10348]_  = \new_[10347]_  | \new_[10340]_ ;
  assign \new_[10351]_  = \new_[479]_  | \new_[480]_ ;
  assign \new_[10354]_  = \new_[477]_  | \new_[478]_ ;
  assign \new_[10355]_  = \new_[10354]_  | \new_[10351]_ ;
  assign \new_[10358]_  = \new_[475]_  | \new_[476]_ ;
  assign \new_[10361]_  = \new_[473]_  | \new_[474]_ ;
  assign \new_[10362]_  = \new_[10361]_  | \new_[10358]_ ;
  assign \new_[10363]_  = \new_[10362]_  | \new_[10355]_ ;
  assign \new_[10364]_  = \new_[10363]_  | \new_[10348]_ ;
  assign \new_[10365]_  = \new_[10364]_  | \new_[10335]_ ;
  assign \new_[10366]_  = \new_[10365]_  | \new_[10306]_ ;
  assign \new_[10367]_  = \new_[10366]_  | \new_[10249]_ ;
  assign \new_[10368]_  = \new_[10367]_  | \new_[10132]_ ;
  assign \new_[10369]_  = \new_[10368]_  | \new_[9897]_ ;
  assign \new_[10373]_  = \new_[470]_  | \new_[471]_ ;
  assign \new_[10374]_  = \new_[472]_  | \new_[10373]_ ;
  assign \new_[10377]_  = \new_[468]_  | \new_[469]_ ;
  assign \new_[10380]_  = \new_[466]_  | \new_[467]_ ;
  assign \new_[10381]_  = \new_[10380]_  | \new_[10377]_ ;
  assign \new_[10382]_  = \new_[10381]_  | \new_[10374]_ ;
  assign \new_[10386]_  = \new_[463]_  | \new_[464]_ ;
  assign \new_[10387]_  = \new_[465]_  | \new_[10386]_ ;
  assign \new_[10390]_  = \new_[461]_  | \new_[462]_ ;
  assign \new_[10393]_  = \new_[459]_  | \new_[460]_ ;
  assign \new_[10394]_  = \new_[10393]_  | \new_[10390]_ ;
  assign \new_[10395]_  = \new_[10394]_  | \new_[10387]_ ;
  assign \new_[10396]_  = \new_[10395]_  | \new_[10382]_ ;
  assign \new_[10400]_  = \new_[456]_  | \new_[457]_ ;
  assign \new_[10401]_  = \new_[458]_  | \new_[10400]_ ;
  assign \new_[10404]_  = \new_[454]_  | \new_[455]_ ;
  assign \new_[10407]_  = \new_[452]_  | \new_[453]_ ;
  assign \new_[10408]_  = \new_[10407]_  | \new_[10404]_ ;
  assign \new_[10409]_  = \new_[10408]_  | \new_[10401]_ ;
  assign \new_[10412]_  = \new_[450]_  | \new_[451]_ ;
  assign \new_[10415]_  = \new_[448]_  | \new_[449]_ ;
  assign \new_[10416]_  = \new_[10415]_  | \new_[10412]_ ;
  assign \new_[10419]_  = \new_[446]_  | \new_[447]_ ;
  assign \new_[10422]_  = \new_[444]_  | \new_[445]_ ;
  assign \new_[10423]_  = \new_[10422]_  | \new_[10419]_ ;
  assign \new_[10424]_  = \new_[10423]_  | \new_[10416]_ ;
  assign \new_[10425]_  = \new_[10424]_  | \new_[10409]_ ;
  assign \new_[10426]_  = \new_[10425]_  | \new_[10396]_ ;
  assign \new_[10430]_  = \new_[441]_  | \new_[442]_ ;
  assign \new_[10431]_  = \new_[443]_  | \new_[10430]_ ;
  assign \new_[10434]_  = \new_[439]_  | \new_[440]_ ;
  assign \new_[10437]_  = \new_[437]_  | \new_[438]_ ;
  assign \new_[10438]_  = \new_[10437]_  | \new_[10434]_ ;
  assign \new_[10439]_  = \new_[10438]_  | \new_[10431]_ ;
  assign \new_[10442]_  = \new_[435]_  | \new_[436]_ ;
  assign \new_[10445]_  = \new_[433]_  | \new_[434]_ ;
  assign \new_[10446]_  = \new_[10445]_  | \new_[10442]_ ;
  assign \new_[10449]_  = \new_[431]_  | \new_[432]_ ;
  assign \new_[10452]_  = \new_[429]_  | \new_[430]_ ;
  assign \new_[10453]_  = \new_[10452]_  | \new_[10449]_ ;
  assign \new_[10454]_  = \new_[10453]_  | \new_[10446]_ ;
  assign \new_[10455]_  = \new_[10454]_  | \new_[10439]_ ;
  assign \new_[10459]_  = \new_[426]_  | \new_[427]_ ;
  assign \new_[10460]_  = \new_[428]_  | \new_[10459]_ ;
  assign \new_[10463]_  = \new_[424]_  | \new_[425]_ ;
  assign \new_[10466]_  = \new_[422]_  | \new_[423]_ ;
  assign \new_[10467]_  = \new_[10466]_  | \new_[10463]_ ;
  assign \new_[10468]_  = \new_[10467]_  | \new_[10460]_ ;
  assign \new_[10471]_  = \new_[420]_  | \new_[421]_ ;
  assign \new_[10474]_  = \new_[418]_  | \new_[419]_ ;
  assign \new_[10475]_  = \new_[10474]_  | \new_[10471]_ ;
  assign \new_[10478]_  = \new_[416]_  | \new_[417]_ ;
  assign \new_[10481]_  = \new_[414]_  | \new_[415]_ ;
  assign \new_[10482]_  = \new_[10481]_  | \new_[10478]_ ;
  assign \new_[10483]_  = \new_[10482]_  | \new_[10475]_ ;
  assign \new_[10484]_  = \new_[10483]_  | \new_[10468]_ ;
  assign \new_[10485]_  = \new_[10484]_  | \new_[10455]_ ;
  assign \new_[10486]_  = \new_[10485]_  | \new_[10426]_ ;
  assign \new_[10490]_  = \new_[411]_  | \new_[412]_ ;
  assign \new_[10491]_  = \new_[413]_  | \new_[10490]_ ;
  assign \new_[10494]_  = \new_[409]_  | \new_[410]_ ;
  assign \new_[10497]_  = \new_[407]_  | \new_[408]_ ;
  assign \new_[10498]_  = \new_[10497]_  | \new_[10494]_ ;
  assign \new_[10499]_  = \new_[10498]_  | \new_[10491]_ ;
  assign \new_[10503]_  = \new_[404]_  | \new_[405]_ ;
  assign \new_[10504]_  = \new_[406]_  | \new_[10503]_ ;
  assign \new_[10507]_  = \new_[402]_  | \new_[403]_ ;
  assign \new_[10510]_  = \new_[400]_  | \new_[401]_ ;
  assign \new_[10511]_  = \new_[10510]_  | \new_[10507]_ ;
  assign \new_[10512]_  = \new_[10511]_  | \new_[10504]_ ;
  assign \new_[10513]_  = \new_[10512]_  | \new_[10499]_ ;
  assign \new_[10517]_  = \new_[397]_  | \new_[398]_ ;
  assign \new_[10518]_  = \new_[399]_  | \new_[10517]_ ;
  assign \new_[10521]_  = \new_[395]_  | \new_[396]_ ;
  assign \new_[10524]_  = \new_[393]_  | \new_[394]_ ;
  assign \new_[10525]_  = \new_[10524]_  | \new_[10521]_ ;
  assign \new_[10526]_  = \new_[10525]_  | \new_[10518]_ ;
  assign \new_[10529]_  = \new_[391]_  | \new_[392]_ ;
  assign \new_[10532]_  = \new_[389]_  | \new_[390]_ ;
  assign \new_[10533]_  = \new_[10532]_  | \new_[10529]_ ;
  assign \new_[10536]_  = \new_[387]_  | \new_[388]_ ;
  assign \new_[10539]_  = \new_[385]_  | \new_[386]_ ;
  assign \new_[10540]_  = \new_[10539]_  | \new_[10536]_ ;
  assign \new_[10541]_  = \new_[10540]_  | \new_[10533]_ ;
  assign \new_[10542]_  = \new_[10541]_  | \new_[10526]_ ;
  assign \new_[10543]_  = \new_[10542]_  | \new_[10513]_ ;
  assign \new_[10547]_  = \new_[382]_  | \new_[383]_ ;
  assign \new_[10548]_  = \new_[384]_  | \new_[10547]_ ;
  assign \new_[10551]_  = \new_[380]_  | \new_[381]_ ;
  assign \new_[10554]_  = \new_[378]_  | \new_[379]_ ;
  assign \new_[10555]_  = \new_[10554]_  | \new_[10551]_ ;
  assign \new_[10556]_  = \new_[10555]_  | \new_[10548]_ ;
  assign \new_[10559]_  = \new_[376]_  | \new_[377]_ ;
  assign \new_[10562]_  = \new_[374]_  | \new_[375]_ ;
  assign \new_[10563]_  = \new_[10562]_  | \new_[10559]_ ;
  assign \new_[10566]_  = \new_[372]_  | \new_[373]_ ;
  assign \new_[10569]_  = \new_[370]_  | \new_[371]_ ;
  assign \new_[10570]_  = \new_[10569]_  | \new_[10566]_ ;
  assign \new_[10571]_  = \new_[10570]_  | \new_[10563]_ ;
  assign \new_[10572]_  = \new_[10571]_  | \new_[10556]_ ;
  assign \new_[10576]_  = \new_[367]_  | \new_[368]_ ;
  assign \new_[10577]_  = \new_[369]_  | \new_[10576]_ ;
  assign \new_[10580]_  = \new_[365]_  | \new_[366]_ ;
  assign \new_[10583]_  = \new_[363]_  | \new_[364]_ ;
  assign \new_[10584]_  = \new_[10583]_  | \new_[10580]_ ;
  assign \new_[10585]_  = \new_[10584]_  | \new_[10577]_ ;
  assign \new_[10588]_  = \new_[361]_  | \new_[362]_ ;
  assign \new_[10591]_  = \new_[359]_  | \new_[360]_ ;
  assign \new_[10592]_  = \new_[10591]_  | \new_[10588]_ ;
  assign \new_[10595]_  = \new_[357]_  | \new_[358]_ ;
  assign \new_[10598]_  = \new_[355]_  | \new_[356]_ ;
  assign \new_[10599]_  = \new_[10598]_  | \new_[10595]_ ;
  assign \new_[10600]_  = \new_[10599]_  | \new_[10592]_ ;
  assign \new_[10601]_  = \new_[10600]_  | \new_[10585]_ ;
  assign \new_[10602]_  = \new_[10601]_  | \new_[10572]_ ;
  assign \new_[10603]_  = \new_[10602]_  | \new_[10543]_ ;
  assign \new_[10604]_  = \new_[10603]_  | \new_[10486]_ ;
  assign \new_[10608]_  = \new_[352]_  | \new_[353]_ ;
  assign \new_[10609]_  = \new_[354]_  | \new_[10608]_ ;
  assign \new_[10612]_  = \new_[350]_  | \new_[351]_ ;
  assign \new_[10615]_  = \new_[348]_  | \new_[349]_ ;
  assign \new_[10616]_  = \new_[10615]_  | \new_[10612]_ ;
  assign \new_[10617]_  = \new_[10616]_  | \new_[10609]_ ;
  assign \new_[10621]_  = \new_[345]_  | \new_[346]_ ;
  assign \new_[10622]_  = \new_[347]_  | \new_[10621]_ ;
  assign \new_[10625]_  = \new_[343]_  | \new_[344]_ ;
  assign \new_[10628]_  = \new_[341]_  | \new_[342]_ ;
  assign \new_[10629]_  = \new_[10628]_  | \new_[10625]_ ;
  assign \new_[10630]_  = \new_[10629]_  | \new_[10622]_ ;
  assign \new_[10631]_  = \new_[10630]_  | \new_[10617]_ ;
  assign \new_[10635]_  = \new_[338]_  | \new_[339]_ ;
  assign \new_[10636]_  = \new_[340]_  | \new_[10635]_ ;
  assign \new_[10639]_  = \new_[336]_  | \new_[337]_ ;
  assign \new_[10642]_  = \new_[334]_  | \new_[335]_ ;
  assign \new_[10643]_  = \new_[10642]_  | \new_[10639]_ ;
  assign \new_[10644]_  = \new_[10643]_  | \new_[10636]_ ;
  assign \new_[10647]_  = \new_[332]_  | \new_[333]_ ;
  assign \new_[10650]_  = \new_[330]_  | \new_[331]_ ;
  assign \new_[10651]_  = \new_[10650]_  | \new_[10647]_ ;
  assign \new_[10654]_  = \new_[328]_  | \new_[329]_ ;
  assign \new_[10657]_  = \new_[326]_  | \new_[327]_ ;
  assign \new_[10658]_  = \new_[10657]_  | \new_[10654]_ ;
  assign \new_[10659]_  = \new_[10658]_  | \new_[10651]_ ;
  assign \new_[10660]_  = \new_[10659]_  | \new_[10644]_ ;
  assign \new_[10661]_  = \new_[10660]_  | \new_[10631]_ ;
  assign \new_[10665]_  = \new_[323]_  | \new_[324]_ ;
  assign \new_[10666]_  = \new_[325]_  | \new_[10665]_ ;
  assign \new_[10669]_  = \new_[321]_  | \new_[322]_ ;
  assign \new_[10672]_  = \new_[319]_  | \new_[320]_ ;
  assign \new_[10673]_  = \new_[10672]_  | \new_[10669]_ ;
  assign \new_[10674]_  = \new_[10673]_  | \new_[10666]_ ;
  assign \new_[10677]_  = \new_[317]_  | \new_[318]_ ;
  assign \new_[10680]_  = \new_[315]_  | \new_[316]_ ;
  assign \new_[10681]_  = \new_[10680]_  | \new_[10677]_ ;
  assign \new_[10684]_  = \new_[313]_  | \new_[314]_ ;
  assign \new_[10687]_  = \new_[311]_  | \new_[312]_ ;
  assign \new_[10688]_  = \new_[10687]_  | \new_[10684]_ ;
  assign \new_[10689]_  = \new_[10688]_  | \new_[10681]_ ;
  assign \new_[10690]_  = \new_[10689]_  | \new_[10674]_ ;
  assign \new_[10694]_  = \new_[308]_  | \new_[309]_ ;
  assign \new_[10695]_  = \new_[310]_  | \new_[10694]_ ;
  assign \new_[10698]_  = \new_[306]_  | \new_[307]_ ;
  assign \new_[10701]_  = \new_[304]_  | \new_[305]_ ;
  assign \new_[10702]_  = \new_[10701]_  | \new_[10698]_ ;
  assign \new_[10703]_  = \new_[10702]_  | \new_[10695]_ ;
  assign \new_[10706]_  = \new_[302]_  | \new_[303]_ ;
  assign \new_[10709]_  = \new_[300]_  | \new_[301]_ ;
  assign \new_[10710]_  = \new_[10709]_  | \new_[10706]_ ;
  assign \new_[10713]_  = \new_[298]_  | \new_[299]_ ;
  assign \new_[10716]_  = \new_[296]_  | \new_[297]_ ;
  assign \new_[10717]_  = \new_[10716]_  | \new_[10713]_ ;
  assign \new_[10718]_  = \new_[10717]_  | \new_[10710]_ ;
  assign \new_[10719]_  = \new_[10718]_  | \new_[10703]_ ;
  assign \new_[10720]_  = \new_[10719]_  | \new_[10690]_ ;
  assign \new_[10721]_  = \new_[10720]_  | \new_[10661]_ ;
  assign \new_[10725]_  = \new_[293]_  | \new_[294]_ ;
  assign \new_[10726]_  = \new_[295]_  | \new_[10725]_ ;
  assign \new_[10729]_  = \new_[291]_  | \new_[292]_ ;
  assign \new_[10732]_  = \new_[289]_  | \new_[290]_ ;
  assign \new_[10733]_  = \new_[10732]_  | \new_[10729]_ ;
  assign \new_[10734]_  = \new_[10733]_  | \new_[10726]_ ;
  assign \new_[10738]_  = \new_[286]_  | \new_[287]_ ;
  assign \new_[10739]_  = \new_[288]_  | \new_[10738]_ ;
  assign \new_[10742]_  = \new_[284]_  | \new_[285]_ ;
  assign \new_[10745]_  = \new_[282]_  | \new_[283]_ ;
  assign \new_[10746]_  = \new_[10745]_  | \new_[10742]_ ;
  assign \new_[10747]_  = \new_[10746]_  | \new_[10739]_ ;
  assign \new_[10748]_  = \new_[10747]_  | \new_[10734]_ ;
  assign \new_[10752]_  = \new_[279]_  | \new_[280]_ ;
  assign \new_[10753]_  = \new_[281]_  | \new_[10752]_ ;
  assign \new_[10756]_  = \new_[277]_  | \new_[278]_ ;
  assign \new_[10759]_  = \new_[275]_  | \new_[276]_ ;
  assign \new_[10760]_  = \new_[10759]_  | \new_[10756]_ ;
  assign \new_[10761]_  = \new_[10760]_  | \new_[10753]_ ;
  assign \new_[10764]_  = \new_[273]_  | \new_[274]_ ;
  assign \new_[10767]_  = \new_[271]_  | \new_[272]_ ;
  assign \new_[10768]_  = \new_[10767]_  | \new_[10764]_ ;
  assign \new_[10771]_  = \new_[269]_  | \new_[270]_ ;
  assign \new_[10774]_  = \new_[267]_  | \new_[268]_ ;
  assign \new_[10775]_  = \new_[10774]_  | \new_[10771]_ ;
  assign \new_[10776]_  = \new_[10775]_  | \new_[10768]_ ;
  assign \new_[10777]_  = \new_[10776]_  | \new_[10761]_ ;
  assign \new_[10778]_  = \new_[10777]_  | \new_[10748]_ ;
  assign \new_[10782]_  = \new_[264]_  | \new_[265]_ ;
  assign \new_[10783]_  = \new_[266]_  | \new_[10782]_ ;
  assign \new_[10786]_  = \new_[262]_  | \new_[263]_ ;
  assign \new_[10789]_  = \new_[260]_  | \new_[261]_ ;
  assign \new_[10790]_  = \new_[10789]_  | \new_[10786]_ ;
  assign \new_[10791]_  = \new_[10790]_  | \new_[10783]_ ;
  assign \new_[10794]_  = \new_[258]_  | \new_[259]_ ;
  assign \new_[10797]_  = \new_[256]_  | \new_[257]_ ;
  assign \new_[10798]_  = \new_[10797]_  | \new_[10794]_ ;
  assign \new_[10801]_  = \new_[254]_  | \new_[255]_ ;
  assign \new_[10804]_  = \new_[252]_  | \new_[253]_ ;
  assign \new_[10805]_  = \new_[10804]_  | \new_[10801]_ ;
  assign \new_[10806]_  = \new_[10805]_  | \new_[10798]_ ;
  assign \new_[10807]_  = \new_[10806]_  | \new_[10791]_ ;
  assign \new_[10811]_  = \new_[249]_  | \new_[250]_ ;
  assign \new_[10812]_  = \new_[251]_  | \new_[10811]_ ;
  assign \new_[10815]_  = \new_[247]_  | \new_[248]_ ;
  assign \new_[10818]_  = \new_[245]_  | \new_[246]_ ;
  assign \new_[10819]_  = \new_[10818]_  | \new_[10815]_ ;
  assign \new_[10820]_  = \new_[10819]_  | \new_[10812]_ ;
  assign \new_[10823]_  = \new_[243]_  | \new_[244]_ ;
  assign \new_[10826]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[10827]_  = \new_[10826]_  | \new_[10823]_ ;
  assign \new_[10830]_  = \new_[239]_  | \new_[240]_ ;
  assign \new_[10833]_  = \new_[237]_  | \new_[238]_ ;
  assign \new_[10834]_  = \new_[10833]_  | \new_[10830]_ ;
  assign \new_[10835]_  = \new_[10834]_  | \new_[10827]_ ;
  assign \new_[10836]_  = \new_[10835]_  | \new_[10820]_ ;
  assign \new_[10837]_  = \new_[10836]_  | \new_[10807]_ ;
  assign \new_[10838]_  = \new_[10837]_  | \new_[10778]_ ;
  assign \new_[10839]_  = \new_[10838]_  | \new_[10721]_ ;
  assign \new_[10840]_  = \new_[10839]_  | \new_[10604]_ ;
  assign \new_[10844]_  = \new_[234]_  | \new_[235]_ ;
  assign \new_[10845]_  = \new_[236]_  | \new_[10844]_ ;
  assign \new_[10848]_  = \new_[232]_  | \new_[233]_ ;
  assign \new_[10851]_  = \new_[230]_  | \new_[231]_ ;
  assign \new_[10852]_  = \new_[10851]_  | \new_[10848]_ ;
  assign \new_[10853]_  = \new_[10852]_  | \new_[10845]_ ;
  assign \new_[10857]_  = \new_[227]_  | \new_[228]_ ;
  assign \new_[10858]_  = \new_[229]_  | \new_[10857]_ ;
  assign \new_[10861]_  = \new_[225]_  | \new_[226]_ ;
  assign \new_[10864]_  = \new_[223]_  | \new_[224]_ ;
  assign \new_[10865]_  = \new_[10864]_  | \new_[10861]_ ;
  assign \new_[10866]_  = \new_[10865]_  | \new_[10858]_ ;
  assign \new_[10867]_  = \new_[10866]_  | \new_[10853]_ ;
  assign \new_[10871]_  = \new_[220]_  | \new_[221]_ ;
  assign \new_[10872]_  = \new_[222]_  | \new_[10871]_ ;
  assign \new_[10875]_  = \new_[218]_  | \new_[219]_ ;
  assign \new_[10878]_  = \new_[216]_  | \new_[217]_ ;
  assign \new_[10879]_  = \new_[10878]_  | \new_[10875]_ ;
  assign \new_[10880]_  = \new_[10879]_  | \new_[10872]_ ;
  assign \new_[10883]_  = \new_[214]_  | \new_[215]_ ;
  assign \new_[10886]_  = \new_[212]_  | \new_[213]_ ;
  assign \new_[10887]_  = \new_[10886]_  | \new_[10883]_ ;
  assign \new_[10890]_  = \new_[210]_  | \new_[211]_ ;
  assign \new_[10893]_  = \new_[208]_  | \new_[209]_ ;
  assign \new_[10894]_  = \new_[10893]_  | \new_[10890]_ ;
  assign \new_[10895]_  = \new_[10894]_  | \new_[10887]_ ;
  assign \new_[10896]_  = \new_[10895]_  | \new_[10880]_ ;
  assign \new_[10897]_  = \new_[10896]_  | \new_[10867]_ ;
  assign \new_[10901]_  = \new_[205]_  | \new_[206]_ ;
  assign \new_[10902]_  = \new_[207]_  | \new_[10901]_ ;
  assign \new_[10905]_  = \new_[203]_  | \new_[204]_ ;
  assign \new_[10908]_  = \new_[201]_  | \new_[202]_ ;
  assign \new_[10909]_  = \new_[10908]_  | \new_[10905]_ ;
  assign \new_[10910]_  = \new_[10909]_  | \new_[10902]_ ;
  assign \new_[10913]_  = \new_[199]_  | \new_[200]_ ;
  assign \new_[10916]_  = \new_[197]_  | \new_[198]_ ;
  assign \new_[10917]_  = \new_[10916]_  | \new_[10913]_ ;
  assign \new_[10920]_  = \new_[195]_  | \new_[196]_ ;
  assign \new_[10923]_  = \new_[193]_  | \new_[194]_ ;
  assign \new_[10924]_  = \new_[10923]_  | \new_[10920]_ ;
  assign \new_[10925]_  = \new_[10924]_  | \new_[10917]_ ;
  assign \new_[10926]_  = \new_[10925]_  | \new_[10910]_ ;
  assign \new_[10930]_  = \new_[190]_  | \new_[191]_ ;
  assign \new_[10931]_  = \new_[192]_  | \new_[10930]_ ;
  assign \new_[10934]_  = \new_[188]_  | \new_[189]_ ;
  assign \new_[10937]_  = \new_[186]_  | \new_[187]_ ;
  assign \new_[10938]_  = \new_[10937]_  | \new_[10934]_ ;
  assign \new_[10939]_  = \new_[10938]_  | \new_[10931]_ ;
  assign \new_[10942]_  = \new_[184]_  | \new_[185]_ ;
  assign \new_[10945]_  = \new_[182]_  | \new_[183]_ ;
  assign \new_[10946]_  = \new_[10945]_  | \new_[10942]_ ;
  assign \new_[10949]_  = \new_[180]_  | \new_[181]_ ;
  assign \new_[10952]_  = \new_[178]_  | \new_[179]_ ;
  assign \new_[10953]_  = \new_[10952]_  | \new_[10949]_ ;
  assign \new_[10954]_  = \new_[10953]_  | \new_[10946]_ ;
  assign \new_[10955]_  = \new_[10954]_  | \new_[10939]_ ;
  assign \new_[10956]_  = \new_[10955]_  | \new_[10926]_ ;
  assign \new_[10957]_  = \new_[10956]_  | \new_[10897]_ ;
  assign \new_[10961]_  = \new_[175]_  | \new_[176]_ ;
  assign \new_[10962]_  = \new_[177]_  | \new_[10961]_ ;
  assign \new_[10965]_  = \new_[173]_  | \new_[174]_ ;
  assign \new_[10968]_  = \new_[171]_  | \new_[172]_ ;
  assign \new_[10969]_  = \new_[10968]_  | \new_[10965]_ ;
  assign \new_[10970]_  = \new_[10969]_  | \new_[10962]_ ;
  assign \new_[10974]_  = \new_[168]_  | \new_[169]_ ;
  assign \new_[10975]_  = \new_[170]_  | \new_[10974]_ ;
  assign \new_[10978]_  = \new_[166]_  | \new_[167]_ ;
  assign \new_[10981]_  = \new_[164]_  | \new_[165]_ ;
  assign \new_[10982]_  = \new_[10981]_  | \new_[10978]_ ;
  assign \new_[10983]_  = \new_[10982]_  | \new_[10975]_ ;
  assign \new_[10984]_  = \new_[10983]_  | \new_[10970]_ ;
  assign \new_[10988]_  = \new_[161]_  | \new_[162]_ ;
  assign \new_[10989]_  = \new_[163]_  | \new_[10988]_ ;
  assign \new_[10992]_  = \new_[159]_  | \new_[160]_ ;
  assign \new_[10995]_  = \new_[157]_  | \new_[158]_ ;
  assign \new_[10996]_  = \new_[10995]_  | \new_[10992]_ ;
  assign \new_[10997]_  = \new_[10996]_  | \new_[10989]_ ;
  assign \new_[11000]_  = \new_[155]_  | \new_[156]_ ;
  assign \new_[11003]_  = \new_[153]_  | \new_[154]_ ;
  assign \new_[11004]_  = \new_[11003]_  | \new_[11000]_ ;
  assign \new_[11007]_  = \new_[151]_  | \new_[152]_ ;
  assign \new_[11010]_  = \new_[149]_  | \new_[150]_ ;
  assign \new_[11011]_  = \new_[11010]_  | \new_[11007]_ ;
  assign \new_[11012]_  = \new_[11011]_  | \new_[11004]_ ;
  assign \new_[11013]_  = \new_[11012]_  | \new_[10997]_ ;
  assign \new_[11014]_  = \new_[11013]_  | \new_[10984]_ ;
  assign \new_[11018]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[11019]_  = \new_[148]_  | \new_[11018]_ ;
  assign \new_[11022]_  = \new_[144]_  | \new_[145]_ ;
  assign \new_[11025]_  = \new_[142]_  | \new_[143]_ ;
  assign \new_[11026]_  = \new_[11025]_  | \new_[11022]_ ;
  assign \new_[11027]_  = \new_[11026]_  | \new_[11019]_ ;
  assign \new_[11030]_  = \new_[140]_  | \new_[141]_ ;
  assign \new_[11033]_  = \new_[138]_  | \new_[139]_ ;
  assign \new_[11034]_  = \new_[11033]_  | \new_[11030]_ ;
  assign \new_[11037]_  = \new_[136]_  | \new_[137]_ ;
  assign \new_[11040]_  = \new_[134]_  | \new_[135]_ ;
  assign \new_[11041]_  = \new_[11040]_  | \new_[11037]_ ;
  assign \new_[11042]_  = \new_[11041]_  | \new_[11034]_ ;
  assign \new_[11043]_  = \new_[11042]_  | \new_[11027]_ ;
  assign \new_[11047]_  = \new_[131]_  | \new_[132]_ ;
  assign \new_[11048]_  = \new_[133]_  | \new_[11047]_ ;
  assign \new_[11051]_  = \new_[129]_  | \new_[130]_ ;
  assign \new_[11054]_  = \new_[127]_  | \new_[128]_ ;
  assign \new_[11055]_  = \new_[11054]_  | \new_[11051]_ ;
  assign \new_[11056]_  = \new_[11055]_  | \new_[11048]_ ;
  assign \new_[11059]_  = \new_[125]_  | \new_[126]_ ;
  assign \new_[11062]_  = \new_[123]_  | \new_[124]_ ;
  assign \new_[11063]_  = \new_[11062]_  | \new_[11059]_ ;
  assign \new_[11066]_  = \new_[121]_  | \new_[122]_ ;
  assign \new_[11069]_  = \new_[119]_  | \new_[120]_ ;
  assign \new_[11070]_  = \new_[11069]_  | \new_[11066]_ ;
  assign \new_[11071]_  = \new_[11070]_  | \new_[11063]_ ;
  assign \new_[11072]_  = \new_[11071]_  | \new_[11056]_ ;
  assign \new_[11073]_  = \new_[11072]_  | \new_[11043]_ ;
  assign \new_[11074]_  = \new_[11073]_  | \new_[11014]_ ;
  assign \new_[11075]_  = \new_[11074]_  | \new_[10957]_ ;
  assign \new_[11079]_  = \new_[116]_  | \new_[117]_ ;
  assign \new_[11080]_  = \new_[118]_  | \new_[11079]_ ;
  assign \new_[11083]_  = \new_[114]_  | \new_[115]_ ;
  assign \new_[11086]_  = \new_[112]_  | \new_[113]_ ;
  assign \new_[11087]_  = \new_[11086]_  | \new_[11083]_ ;
  assign \new_[11088]_  = \new_[11087]_  | \new_[11080]_ ;
  assign \new_[11092]_  = \new_[109]_  | \new_[110]_ ;
  assign \new_[11093]_  = \new_[111]_  | \new_[11092]_ ;
  assign \new_[11096]_  = \new_[107]_  | \new_[108]_ ;
  assign \new_[11099]_  = \new_[105]_  | \new_[106]_ ;
  assign \new_[11100]_  = \new_[11099]_  | \new_[11096]_ ;
  assign \new_[11101]_  = \new_[11100]_  | \new_[11093]_ ;
  assign \new_[11102]_  = \new_[11101]_  | \new_[11088]_ ;
  assign \new_[11106]_  = \new_[102]_  | \new_[103]_ ;
  assign \new_[11107]_  = \new_[104]_  | \new_[11106]_ ;
  assign \new_[11110]_  = \new_[100]_  | \new_[101]_ ;
  assign \new_[11113]_  = \new_[98]_  | \new_[99]_ ;
  assign \new_[11114]_  = \new_[11113]_  | \new_[11110]_ ;
  assign \new_[11115]_  = \new_[11114]_  | \new_[11107]_ ;
  assign \new_[11118]_  = \new_[96]_  | \new_[97]_ ;
  assign \new_[11121]_  = \new_[94]_  | \new_[95]_ ;
  assign \new_[11122]_  = \new_[11121]_  | \new_[11118]_ ;
  assign \new_[11125]_  = \new_[92]_  | \new_[93]_ ;
  assign \new_[11128]_  = \new_[90]_  | \new_[91]_ ;
  assign \new_[11129]_  = \new_[11128]_  | \new_[11125]_ ;
  assign \new_[11130]_  = \new_[11129]_  | \new_[11122]_ ;
  assign \new_[11131]_  = \new_[11130]_  | \new_[11115]_ ;
  assign \new_[11132]_  = \new_[11131]_  | \new_[11102]_ ;
  assign \new_[11136]_  = \new_[87]_  | \new_[88]_ ;
  assign \new_[11137]_  = \new_[89]_  | \new_[11136]_ ;
  assign \new_[11140]_  = \new_[85]_  | \new_[86]_ ;
  assign \new_[11143]_  = \new_[83]_  | \new_[84]_ ;
  assign \new_[11144]_  = \new_[11143]_  | \new_[11140]_ ;
  assign \new_[11145]_  = \new_[11144]_  | \new_[11137]_ ;
  assign \new_[11148]_  = \new_[81]_  | \new_[82]_ ;
  assign \new_[11151]_  = \new_[79]_  | \new_[80]_ ;
  assign \new_[11152]_  = \new_[11151]_  | \new_[11148]_ ;
  assign \new_[11155]_  = \new_[77]_  | \new_[78]_ ;
  assign \new_[11158]_  = \new_[75]_  | \new_[76]_ ;
  assign \new_[11159]_  = \new_[11158]_  | \new_[11155]_ ;
  assign \new_[11160]_  = \new_[11159]_  | \new_[11152]_ ;
  assign \new_[11161]_  = \new_[11160]_  | \new_[11145]_ ;
  assign \new_[11165]_  = \new_[72]_  | \new_[73]_ ;
  assign \new_[11166]_  = \new_[74]_  | \new_[11165]_ ;
  assign \new_[11169]_  = \new_[70]_  | \new_[71]_ ;
  assign \new_[11172]_  = \new_[68]_  | \new_[69]_ ;
  assign \new_[11173]_  = \new_[11172]_  | \new_[11169]_ ;
  assign \new_[11174]_  = \new_[11173]_  | \new_[11166]_ ;
  assign \new_[11177]_  = \new_[66]_  | \new_[67]_ ;
  assign \new_[11180]_  = \new_[64]_  | \new_[65]_ ;
  assign \new_[11181]_  = \new_[11180]_  | \new_[11177]_ ;
  assign \new_[11184]_  = \new_[62]_  | \new_[63]_ ;
  assign \new_[11187]_  = \new_[60]_  | \new_[61]_ ;
  assign \new_[11188]_  = \new_[11187]_  | \new_[11184]_ ;
  assign \new_[11189]_  = \new_[11188]_  | \new_[11181]_ ;
  assign \new_[11190]_  = \new_[11189]_  | \new_[11174]_ ;
  assign \new_[11191]_  = \new_[11190]_  | \new_[11161]_ ;
  assign \new_[11192]_  = \new_[11191]_  | \new_[11132]_ ;
  assign \new_[11196]_  = \new_[57]_  | \new_[58]_ ;
  assign \new_[11197]_  = \new_[59]_  | \new_[11196]_ ;
  assign \new_[11200]_  = \new_[55]_  | \new_[56]_ ;
  assign \new_[11203]_  = \new_[53]_  | \new_[54]_ ;
  assign \new_[11204]_  = \new_[11203]_  | \new_[11200]_ ;
  assign \new_[11205]_  = \new_[11204]_  | \new_[11197]_ ;
  assign \new_[11209]_  = \new_[50]_  | \new_[51]_ ;
  assign \new_[11210]_  = \new_[52]_  | \new_[11209]_ ;
  assign \new_[11213]_  = \new_[48]_  | \new_[49]_ ;
  assign \new_[11216]_  = \new_[46]_  | \new_[47]_ ;
  assign \new_[11217]_  = \new_[11216]_  | \new_[11213]_ ;
  assign \new_[11218]_  = \new_[11217]_  | \new_[11210]_ ;
  assign \new_[11219]_  = \new_[11218]_  | \new_[11205]_ ;
  assign \new_[11223]_  = \new_[43]_  | \new_[44]_ ;
  assign \new_[11224]_  = \new_[45]_  | \new_[11223]_ ;
  assign \new_[11227]_  = \new_[41]_  | \new_[42]_ ;
  assign \new_[11230]_  = \new_[39]_  | \new_[40]_ ;
  assign \new_[11231]_  = \new_[11230]_  | \new_[11227]_ ;
  assign \new_[11232]_  = \new_[11231]_  | \new_[11224]_ ;
  assign \new_[11235]_  = \new_[37]_  | \new_[38]_ ;
  assign \new_[11238]_  = \new_[35]_  | \new_[36]_ ;
  assign \new_[11239]_  = \new_[11238]_  | \new_[11235]_ ;
  assign \new_[11242]_  = \new_[33]_  | \new_[34]_ ;
  assign \new_[11245]_  = \new_[31]_  | \new_[32]_ ;
  assign \new_[11246]_  = \new_[11245]_  | \new_[11242]_ ;
  assign \new_[11247]_  = \new_[11246]_  | \new_[11239]_ ;
  assign \new_[11248]_  = \new_[11247]_  | \new_[11232]_ ;
  assign \new_[11249]_  = \new_[11248]_  | \new_[11219]_ ;
  assign \new_[11253]_  = \new_[28]_  | \new_[29]_ ;
  assign \new_[11254]_  = \new_[30]_  | \new_[11253]_ ;
  assign \new_[11257]_  = \new_[26]_  | \new_[27]_ ;
  assign \new_[11260]_  = \new_[24]_  | \new_[25]_ ;
  assign \new_[11261]_  = \new_[11260]_  | \new_[11257]_ ;
  assign \new_[11262]_  = \new_[11261]_  | \new_[11254]_ ;
  assign \new_[11265]_  = \new_[22]_  | \new_[23]_ ;
  assign \new_[11268]_  = \new_[20]_  | \new_[21]_ ;
  assign \new_[11269]_  = \new_[11268]_  | \new_[11265]_ ;
  assign \new_[11272]_  = \new_[18]_  | \new_[19]_ ;
  assign \new_[11275]_  = \new_[16]_  | \new_[17]_ ;
  assign \new_[11276]_  = \new_[11275]_  | \new_[11272]_ ;
  assign \new_[11277]_  = \new_[11276]_  | \new_[11269]_ ;
  assign \new_[11278]_  = \new_[11277]_  | \new_[11262]_ ;
  assign \new_[11282]_  = \new_[13]_  | \new_[14]_ ;
  assign \new_[11283]_  = \new_[15]_  | \new_[11282]_ ;
  assign \new_[11286]_  = \new_[11]_  | \new_[12]_ ;
  assign \new_[11289]_  = \new_[9]_  | \new_[10]_ ;
  assign \new_[11290]_  = \new_[11289]_  | \new_[11286]_ ;
  assign \new_[11291]_  = \new_[11290]_  | \new_[11283]_ ;
  assign \new_[11294]_  = \new_[7]_  | \new_[8]_ ;
  assign \new_[11297]_  = \new_[5]_  | \new_[6]_ ;
  assign \new_[11298]_  = \new_[11297]_  | \new_[11294]_ ;
  assign \new_[11301]_  = \new_[3]_  | \new_[4]_ ;
  assign \new_[11304]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[11305]_  = \new_[11304]_  | \new_[11301]_ ;
  assign \new_[11306]_  = \new_[11305]_  | \new_[11298]_ ;
  assign \new_[11307]_  = \new_[11306]_  | \new_[11291]_ ;
  assign \new_[11308]_  = \new_[11307]_  | \new_[11278]_ ;
  assign \new_[11309]_  = \new_[11308]_  | \new_[11249]_ ;
  assign \new_[11310]_  = \new_[11309]_  | \new_[11192]_ ;
  assign \new_[11311]_  = \new_[11310]_  | \new_[11075]_ ;
  assign \new_[11312]_  = \new_[11311]_  | \new_[10840]_ ;
  assign \new_[11313]_  = \new_[11312]_  | \new_[10369]_ ;
  assign \new_[11314]_  = \new_[11313]_  | \new_[9428]_ ;
  assign \new_[11317]_  = A166 & A168;
  assign \new_[11320]_  = A200 & A199;
  assign \new_[11321]_  = \new_[11320]_  & \new_[11317]_ ;
  assign \new_[11324]_  = A233 & ~A232;
  assign \new_[11327]_  = A299 & ~A298;
  assign \new_[11328]_  = \new_[11327]_  & \new_[11324]_ ;
  assign \new_[11331]_  = A166 & A168;
  assign \new_[11334]_  = A200 & A199;
  assign \new_[11335]_  = \new_[11334]_  & \new_[11331]_ ;
  assign \new_[11338]_  = A233 & ~A232;
  assign \new_[11341]_  = A266 & ~A265;
  assign \new_[11342]_  = \new_[11341]_  & \new_[11338]_ ;
  assign \new_[11345]_  = A166 & A168;
  assign \new_[11348]_  = ~A201 & ~A200;
  assign \new_[11349]_  = \new_[11348]_  & \new_[11345]_ ;
  assign \new_[11352]_  = A233 & ~A232;
  assign \new_[11355]_  = A299 & ~A298;
  assign \new_[11356]_  = \new_[11355]_  & \new_[11352]_ ;
  assign \new_[11359]_  = A166 & A168;
  assign \new_[11362]_  = ~A201 & ~A200;
  assign \new_[11363]_  = \new_[11362]_  & \new_[11359]_ ;
  assign \new_[11366]_  = A233 & ~A232;
  assign \new_[11369]_  = A266 & ~A265;
  assign \new_[11370]_  = \new_[11369]_  & \new_[11366]_ ;
  assign \new_[11373]_  = A166 & A168;
  assign \new_[11376]_  = ~A200 & ~A199;
  assign \new_[11377]_  = \new_[11376]_  & \new_[11373]_ ;
  assign \new_[11380]_  = A233 & ~A232;
  assign \new_[11383]_  = A299 & ~A298;
  assign \new_[11384]_  = \new_[11383]_  & \new_[11380]_ ;
  assign \new_[11387]_  = A166 & A168;
  assign \new_[11390]_  = ~A200 & ~A199;
  assign \new_[11391]_  = \new_[11390]_  & \new_[11387]_ ;
  assign \new_[11394]_  = A233 & ~A232;
  assign \new_[11397]_  = A266 & ~A265;
  assign \new_[11398]_  = \new_[11397]_  & \new_[11394]_ ;
  assign \new_[11401]_  = A167 & A168;
  assign \new_[11404]_  = A200 & A199;
  assign \new_[11405]_  = \new_[11404]_  & \new_[11401]_ ;
  assign \new_[11408]_  = A233 & ~A232;
  assign \new_[11411]_  = A299 & ~A298;
  assign \new_[11412]_  = \new_[11411]_  & \new_[11408]_ ;
  assign \new_[11415]_  = A167 & A168;
  assign \new_[11418]_  = A200 & A199;
  assign \new_[11419]_  = \new_[11418]_  & \new_[11415]_ ;
  assign \new_[11422]_  = A233 & ~A232;
  assign \new_[11425]_  = A266 & ~A265;
  assign \new_[11426]_  = \new_[11425]_  & \new_[11422]_ ;
  assign \new_[11429]_  = A167 & A168;
  assign \new_[11432]_  = ~A201 & ~A200;
  assign \new_[11433]_  = \new_[11432]_  & \new_[11429]_ ;
  assign \new_[11436]_  = A233 & ~A232;
  assign \new_[11439]_  = A299 & ~A298;
  assign \new_[11440]_  = \new_[11439]_  & \new_[11436]_ ;
  assign \new_[11443]_  = A167 & A168;
  assign \new_[11446]_  = ~A201 & ~A200;
  assign \new_[11447]_  = \new_[11446]_  & \new_[11443]_ ;
  assign \new_[11450]_  = A233 & ~A232;
  assign \new_[11453]_  = A266 & ~A265;
  assign \new_[11454]_  = \new_[11453]_  & \new_[11450]_ ;
  assign \new_[11457]_  = A167 & A168;
  assign \new_[11460]_  = ~A200 & ~A199;
  assign \new_[11461]_  = \new_[11460]_  & \new_[11457]_ ;
  assign \new_[11464]_  = A233 & ~A232;
  assign \new_[11467]_  = A299 & ~A298;
  assign \new_[11468]_  = \new_[11467]_  & \new_[11464]_ ;
  assign \new_[11471]_  = A167 & A168;
  assign \new_[11474]_  = ~A200 & ~A199;
  assign \new_[11475]_  = \new_[11474]_  & \new_[11471]_ ;
  assign \new_[11478]_  = A233 & ~A232;
  assign \new_[11481]_  = A266 & ~A265;
  assign \new_[11482]_  = \new_[11481]_  & \new_[11478]_ ;
  assign \new_[11485]_  = A166 & A168;
  assign \new_[11488]_  = ~A202 & ~A200;
  assign \new_[11489]_  = \new_[11488]_  & \new_[11485]_ ;
  assign \new_[11492]_  = ~A232 & ~A203;
  assign \new_[11496]_  = A299 & ~A298;
  assign \new_[11497]_  = A233 & \new_[11496]_ ;
  assign \new_[11498]_  = \new_[11497]_  & \new_[11492]_ ;
  assign \new_[11501]_  = A166 & A168;
  assign \new_[11504]_  = ~A202 & ~A200;
  assign \new_[11505]_  = \new_[11504]_  & \new_[11501]_ ;
  assign \new_[11508]_  = ~A232 & ~A203;
  assign \new_[11512]_  = A266 & ~A265;
  assign \new_[11513]_  = A233 & \new_[11512]_ ;
  assign \new_[11514]_  = \new_[11513]_  & \new_[11508]_ ;
  assign \new_[11517]_  = A167 & A168;
  assign \new_[11520]_  = ~A202 & ~A200;
  assign \new_[11521]_  = \new_[11520]_  & \new_[11517]_ ;
  assign \new_[11524]_  = ~A232 & ~A203;
  assign \new_[11528]_  = A299 & ~A298;
  assign \new_[11529]_  = A233 & \new_[11528]_ ;
  assign \new_[11530]_  = \new_[11529]_  & \new_[11524]_ ;
  assign \new_[11533]_  = A167 & A168;
  assign \new_[11536]_  = ~A202 & ~A200;
  assign \new_[11537]_  = \new_[11536]_  & \new_[11533]_ ;
  assign \new_[11540]_  = ~A232 & ~A203;
  assign \new_[11544]_  = A266 & ~A265;
  assign \new_[11545]_  = A233 & \new_[11544]_ ;
  assign \new_[11546]_  = \new_[11545]_  & \new_[11540]_ ;
  assign \new_[11549]_  = ~A167 & A170;
  assign \new_[11552]_  = ~A199 & ~A166;
  assign \new_[11553]_  = \new_[11552]_  & \new_[11549]_ ;
  assign \new_[11556]_  = ~A232 & A200;
  assign \new_[11560]_  = A299 & ~A298;
  assign \new_[11561]_  = A233 & \new_[11560]_ ;
  assign \new_[11562]_  = \new_[11561]_  & \new_[11556]_ ;
  assign \new_[11565]_  = ~A167 & A170;
  assign \new_[11568]_  = ~A199 & ~A166;
  assign \new_[11569]_  = \new_[11568]_  & \new_[11565]_ ;
  assign \new_[11572]_  = ~A232 & A200;
  assign \new_[11576]_  = A266 & ~A265;
  assign \new_[11577]_  = A233 & \new_[11576]_ ;
  assign \new_[11578]_  = \new_[11577]_  & \new_[11572]_ ;
  assign \new_[11581]_  = ~A167 & ~A169;
  assign \new_[11584]_  = ~A199 & ~A166;
  assign \new_[11585]_  = \new_[11584]_  & \new_[11581]_ ;
  assign \new_[11588]_  = ~A232 & A200;
  assign \new_[11592]_  = A299 & ~A298;
  assign \new_[11593]_  = A233 & \new_[11592]_ ;
  assign \new_[11594]_  = \new_[11593]_  & \new_[11588]_ ;
  assign \new_[11597]_  = ~A167 & ~A169;
  assign \new_[11600]_  = ~A199 & ~A166;
  assign \new_[11601]_  = \new_[11600]_  & \new_[11597]_ ;
  assign \new_[11604]_  = ~A232 & A200;
  assign \new_[11608]_  = A266 & ~A265;
  assign \new_[11609]_  = A233 & \new_[11608]_ ;
  assign \new_[11610]_  = \new_[11609]_  & \new_[11604]_ ;
  assign \new_[11613]_  = A166 & A168;
  assign \new_[11617]_  = A232 & A200;
  assign \new_[11618]_  = A199 & \new_[11617]_ ;
  assign \new_[11619]_  = \new_[11618]_  & \new_[11613]_ ;
  assign \new_[11622]_  = A265 & A233;
  assign \new_[11626]_  = ~A300 & ~A299;
  assign \new_[11627]_  = ~A267 & \new_[11626]_ ;
  assign \new_[11628]_  = \new_[11627]_  & \new_[11622]_ ;
  assign \new_[11631]_  = A166 & A168;
  assign \new_[11635]_  = A232 & A200;
  assign \new_[11636]_  = A199 & \new_[11635]_ ;
  assign \new_[11637]_  = \new_[11636]_  & \new_[11631]_ ;
  assign \new_[11640]_  = A265 & A233;
  assign \new_[11644]_  = A299 & A298;
  assign \new_[11645]_  = ~A267 & \new_[11644]_ ;
  assign \new_[11646]_  = \new_[11645]_  & \new_[11640]_ ;
  assign \new_[11649]_  = A166 & A168;
  assign \new_[11653]_  = A232 & A200;
  assign \new_[11654]_  = A199 & \new_[11653]_ ;
  assign \new_[11655]_  = \new_[11654]_  & \new_[11649]_ ;
  assign \new_[11658]_  = A265 & A233;
  assign \new_[11662]_  = ~A299 & ~A298;
  assign \new_[11663]_  = ~A267 & \new_[11662]_ ;
  assign \new_[11664]_  = \new_[11663]_  & \new_[11658]_ ;
  assign \new_[11667]_  = A166 & A168;
  assign \new_[11671]_  = A232 & A200;
  assign \new_[11672]_  = A199 & \new_[11671]_ ;
  assign \new_[11673]_  = \new_[11672]_  & \new_[11667]_ ;
  assign \new_[11676]_  = A265 & A233;
  assign \new_[11680]_  = ~A300 & ~A299;
  assign \new_[11681]_  = A266 & \new_[11680]_ ;
  assign \new_[11682]_  = \new_[11681]_  & \new_[11676]_ ;
  assign \new_[11685]_  = A166 & A168;
  assign \new_[11689]_  = A232 & A200;
  assign \new_[11690]_  = A199 & \new_[11689]_ ;
  assign \new_[11691]_  = \new_[11690]_  & \new_[11685]_ ;
  assign \new_[11694]_  = A265 & A233;
  assign \new_[11698]_  = A299 & A298;
  assign \new_[11699]_  = A266 & \new_[11698]_ ;
  assign \new_[11700]_  = \new_[11699]_  & \new_[11694]_ ;
  assign \new_[11703]_  = A166 & A168;
  assign \new_[11707]_  = A232 & A200;
  assign \new_[11708]_  = A199 & \new_[11707]_ ;
  assign \new_[11709]_  = \new_[11708]_  & \new_[11703]_ ;
  assign \new_[11712]_  = A265 & A233;
  assign \new_[11716]_  = ~A299 & ~A298;
  assign \new_[11717]_  = A266 & \new_[11716]_ ;
  assign \new_[11718]_  = \new_[11717]_  & \new_[11712]_ ;
  assign \new_[11721]_  = A166 & A168;
  assign \new_[11725]_  = A232 & A200;
  assign \new_[11726]_  = A199 & \new_[11725]_ ;
  assign \new_[11727]_  = \new_[11726]_  & \new_[11721]_ ;
  assign \new_[11730]_  = ~A265 & A233;
  assign \new_[11734]_  = ~A300 & ~A299;
  assign \new_[11735]_  = ~A266 & \new_[11734]_ ;
  assign \new_[11736]_  = \new_[11735]_  & \new_[11730]_ ;
  assign \new_[11739]_  = A166 & A168;
  assign \new_[11743]_  = A232 & A200;
  assign \new_[11744]_  = A199 & \new_[11743]_ ;
  assign \new_[11745]_  = \new_[11744]_  & \new_[11739]_ ;
  assign \new_[11748]_  = ~A265 & A233;
  assign \new_[11752]_  = A299 & A298;
  assign \new_[11753]_  = ~A266 & \new_[11752]_ ;
  assign \new_[11754]_  = \new_[11753]_  & \new_[11748]_ ;
  assign \new_[11757]_  = A166 & A168;
  assign \new_[11761]_  = A232 & A200;
  assign \new_[11762]_  = A199 & \new_[11761]_ ;
  assign \new_[11763]_  = \new_[11762]_  & \new_[11757]_ ;
  assign \new_[11766]_  = ~A265 & A233;
  assign \new_[11770]_  = ~A299 & ~A298;
  assign \new_[11771]_  = ~A266 & \new_[11770]_ ;
  assign \new_[11772]_  = \new_[11771]_  & \new_[11766]_ ;
  assign \new_[11775]_  = A166 & A168;
  assign \new_[11779]_  = ~A232 & A200;
  assign \new_[11780]_  = A199 & \new_[11779]_ ;
  assign \new_[11781]_  = \new_[11780]_  & \new_[11775]_ ;
  assign \new_[11784]_  = A298 & A233;
  assign \new_[11788]_  = A301 & A300;
  assign \new_[11789]_  = ~A299 & \new_[11788]_ ;
  assign \new_[11790]_  = \new_[11789]_  & \new_[11784]_ ;
  assign \new_[11793]_  = A166 & A168;
  assign \new_[11797]_  = ~A232 & A200;
  assign \new_[11798]_  = A199 & \new_[11797]_ ;
  assign \new_[11799]_  = \new_[11798]_  & \new_[11793]_ ;
  assign \new_[11802]_  = A298 & A233;
  assign \new_[11806]_  = A302 & A300;
  assign \new_[11807]_  = ~A299 & \new_[11806]_ ;
  assign \new_[11808]_  = \new_[11807]_  & \new_[11802]_ ;
  assign \new_[11811]_  = A166 & A168;
  assign \new_[11815]_  = ~A232 & A200;
  assign \new_[11816]_  = A199 & \new_[11815]_ ;
  assign \new_[11817]_  = \new_[11816]_  & \new_[11811]_ ;
  assign \new_[11820]_  = A265 & A233;
  assign \new_[11824]_  = A268 & A267;
  assign \new_[11825]_  = ~A266 & \new_[11824]_ ;
  assign \new_[11826]_  = \new_[11825]_  & \new_[11820]_ ;
  assign \new_[11829]_  = A166 & A168;
  assign \new_[11833]_  = ~A232 & A200;
  assign \new_[11834]_  = A199 & \new_[11833]_ ;
  assign \new_[11835]_  = \new_[11834]_  & \new_[11829]_ ;
  assign \new_[11838]_  = A265 & A233;
  assign \new_[11842]_  = A269 & A267;
  assign \new_[11843]_  = ~A266 & \new_[11842]_ ;
  assign \new_[11844]_  = \new_[11843]_  & \new_[11838]_ ;
  assign \new_[11847]_  = A166 & A168;
  assign \new_[11851]_  = ~A233 & A200;
  assign \new_[11852]_  = A199 & \new_[11851]_ ;
  assign \new_[11853]_  = \new_[11852]_  & \new_[11847]_ ;
  assign \new_[11856]_  = A265 & ~A234;
  assign \new_[11860]_  = ~A300 & A298;
  assign \new_[11861]_  = A266 & \new_[11860]_ ;
  assign \new_[11862]_  = \new_[11861]_  & \new_[11856]_ ;
  assign \new_[11865]_  = A166 & A168;
  assign \new_[11869]_  = ~A233 & A200;
  assign \new_[11870]_  = A199 & \new_[11869]_ ;
  assign \new_[11871]_  = \new_[11870]_  & \new_[11865]_ ;
  assign \new_[11874]_  = A265 & ~A234;
  assign \new_[11878]_  = A299 & A298;
  assign \new_[11879]_  = A266 & \new_[11878]_ ;
  assign \new_[11880]_  = \new_[11879]_  & \new_[11874]_ ;
  assign \new_[11883]_  = A166 & A168;
  assign \new_[11887]_  = ~A233 & A200;
  assign \new_[11888]_  = A199 & \new_[11887]_ ;
  assign \new_[11889]_  = \new_[11888]_  & \new_[11883]_ ;
  assign \new_[11892]_  = A265 & ~A234;
  assign \new_[11896]_  = ~A299 & ~A298;
  assign \new_[11897]_  = A266 & \new_[11896]_ ;
  assign \new_[11898]_  = \new_[11897]_  & \new_[11892]_ ;
  assign \new_[11901]_  = A166 & A168;
  assign \new_[11905]_  = ~A233 & A200;
  assign \new_[11906]_  = A199 & \new_[11905]_ ;
  assign \new_[11907]_  = \new_[11906]_  & \new_[11901]_ ;
  assign \new_[11910]_  = ~A266 & ~A234;
  assign \new_[11914]_  = ~A300 & A298;
  assign \new_[11915]_  = ~A267 & \new_[11914]_ ;
  assign \new_[11916]_  = \new_[11915]_  & \new_[11910]_ ;
  assign \new_[11919]_  = A166 & A168;
  assign \new_[11923]_  = ~A233 & A200;
  assign \new_[11924]_  = A199 & \new_[11923]_ ;
  assign \new_[11925]_  = \new_[11924]_  & \new_[11919]_ ;
  assign \new_[11928]_  = ~A266 & ~A234;
  assign \new_[11932]_  = A299 & A298;
  assign \new_[11933]_  = ~A267 & \new_[11932]_ ;
  assign \new_[11934]_  = \new_[11933]_  & \new_[11928]_ ;
  assign \new_[11937]_  = A166 & A168;
  assign \new_[11941]_  = ~A233 & A200;
  assign \new_[11942]_  = A199 & \new_[11941]_ ;
  assign \new_[11943]_  = \new_[11942]_  & \new_[11937]_ ;
  assign \new_[11946]_  = ~A266 & ~A234;
  assign \new_[11950]_  = ~A299 & ~A298;
  assign \new_[11951]_  = ~A267 & \new_[11950]_ ;
  assign \new_[11952]_  = \new_[11951]_  & \new_[11946]_ ;
  assign \new_[11955]_  = A166 & A168;
  assign \new_[11959]_  = ~A233 & A200;
  assign \new_[11960]_  = A199 & \new_[11959]_ ;
  assign \new_[11961]_  = \new_[11960]_  & \new_[11955]_ ;
  assign \new_[11964]_  = ~A265 & ~A234;
  assign \new_[11968]_  = ~A300 & A298;
  assign \new_[11969]_  = ~A266 & \new_[11968]_ ;
  assign \new_[11970]_  = \new_[11969]_  & \new_[11964]_ ;
  assign \new_[11973]_  = A166 & A168;
  assign \new_[11977]_  = ~A233 & A200;
  assign \new_[11978]_  = A199 & \new_[11977]_ ;
  assign \new_[11979]_  = \new_[11978]_  & \new_[11973]_ ;
  assign \new_[11982]_  = ~A265 & ~A234;
  assign \new_[11986]_  = A299 & A298;
  assign \new_[11987]_  = ~A266 & \new_[11986]_ ;
  assign \new_[11988]_  = \new_[11987]_  & \new_[11982]_ ;
  assign \new_[11991]_  = A166 & A168;
  assign \new_[11995]_  = ~A233 & A200;
  assign \new_[11996]_  = A199 & \new_[11995]_ ;
  assign \new_[11997]_  = \new_[11996]_  & \new_[11991]_ ;
  assign \new_[12000]_  = ~A265 & ~A234;
  assign \new_[12004]_  = ~A299 & ~A298;
  assign \new_[12005]_  = ~A266 & \new_[12004]_ ;
  assign \new_[12006]_  = \new_[12005]_  & \new_[12000]_ ;
  assign \new_[12009]_  = A166 & A168;
  assign \new_[12013]_  = A232 & A200;
  assign \new_[12014]_  = A199 & \new_[12013]_ ;
  assign \new_[12015]_  = \new_[12014]_  & \new_[12009]_ ;
  assign \new_[12018]_  = A234 & ~A233;
  assign \new_[12022]_  = A299 & ~A298;
  assign \new_[12023]_  = A235 & \new_[12022]_ ;
  assign \new_[12024]_  = \new_[12023]_  & \new_[12018]_ ;
  assign \new_[12027]_  = A166 & A168;
  assign \new_[12031]_  = A232 & A200;
  assign \new_[12032]_  = A199 & \new_[12031]_ ;
  assign \new_[12033]_  = \new_[12032]_  & \new_[12027]_ ;
  assign \new_[12036]_  = A234 & ~A233;
  assign \new_[12040]_  = A266 & ~A265;
  assign \new_[12041]_  = A235 & \new_[12040]_ ;
  assign \new_[12042]_  = \new_[12041]_  & \new_[12036]_ ;
  assign \new_[12045]_  = A166 & A168;
  assign \new_[12049]_  = A232 & A200;
  assign \new_[12050]_  = A199 & \new_[12049]_ ;
  assign \new_[12051]_  = \new_[12050]_  & \new_[12045]_ ;
  assign \new_[12054]_  = A234 & ~A233;
  assign \new_[12058]_  = A299 & ~A298;
  assign \new_[12059]_  = A236 & \new_[12058]_ ;
  assign \new_[12060]_  = \new_[12059]_  & \new_[12054]_ ;
  assign \new_[12063]_  = A166 & A168;
  assign \new_[12067]_  = A232 & A200;
  assign \new_[12068]_  = A199 & \new_[12067]_ ;
  assign \new_[12069]_  = \new_[12068]_  & \new_[12063]_ ;
  assign \new_[12072]_  = A234 & ~A233;
  assign \new_[12076]_  = A266 & ~A265;
  assign \new_[12077]_  = A236 & \new_[12076]_ ;
  assign \new_[12078]_  = \new_[12077]_  & \new_[12072]_ ;
  assign \new_[12081]_  = A166 & A168;
  assign \new_[12085]_  = ~A232 & A200;
  assign \new_[12086]_  = A199 & \new_[12085]_ ;
  assign \new_[12087]_  = \new_[12086]_  & \new_[12081]_ ;
  assign \new_[12090]_  = A265 & ~A233;
  assign \new_[12094]_  = ~A300 & A298;
  assign \new_[12095]_  = A266 & \new_[12094]_ ;
  assign \new_[12096]_  = \new_[12095]_  & \new_[12090]_ ;
  assign \new_[12099]_  = A166 & A168;
  assign \new_[12103]_  = ~A232 & A200;
  assign \new_[12104]_  = A199 & \new_[12103]_ ;
  assign \new_[12105]_  = \new_[12104]_  & \new_[12099]_ ;
  assign \new_[12108]_  = A265 & ~A233;
  assign \new_[12112]_  = A299 & A298;
  assign \new_[12113]_  = A266 & \new_[12112]_ ;
  assign \new_[12114]_  = \new_[12113]_  & \new_[12108]_ ;
  assign \new_[12117]_  = A166 & A168;
  assign \new_[12121]_  = ~A232 & A200;
  assign \new_[12122]_  = A199 & \new_[12121]_ ;
  assign \new_[12123]_  = \new_[12122]_  & \new_[12117]_ ;
  assign \new_[12126]_  = A265 & ~A233;
  assign \new_[12130]_  = ~A299 & ~A298;
  assign \new_[12131]_  = A266 & \new_[12130]_ ;
  assign \new_[12132]_  = \new_[12131]_  & \new_[12126]_ ;
  assign \new_[12135]_  = A166 & A168;
  assign \new_[12139]_  = ~A232 & A200;
  assign \new_[12140]_  = A199 & \new_[12139]_ ;
  assign \new_[12141]_  = \new_[12140]_  & \new_[12135]_ ;
  assign \new_[12144]_  = ~A266 & ~A233;
  assign \new_[12148]_  = ~A300 & A298;
  assign \new_[12149]_  = ~A267 & \new_[12148]_ ;
  assign \new_[12150]_  = \new_[12149]_  & \new_[12144]_ ;
  assign \new_[12153]_  = A166 & A168;
  assign \new_[12157]_  = ~A232 & A200;
  assign \new_[12158]_  = A199 & \new_[12157]_ ;
  assign \new_[12159]_  = \new_[12158]_  & \new_[12153]_ ;
  assign \new_[12162]_  = ~A266 & ~A233;
  assign \new_[12166]_  = A299 & A298;
  assign \new_[12167]_  = ~A267 & \new_[12166]_ ;
  assign \new_[12168]_  = \new_[12167]_  & \new_[12162]_ ;
  assign \new_[12171]_  = A166 & A168;
  assign \new_[12175]_  = ~A232 & A200;
  assign \new_[12176]_  = A199 & \new_[12175]_ ;
  assign \new_[12177]_  = \new_[12176]_  & \new_[12171]_ ;
  assign \new_[12180]_  = ~A266 & ~A233;
  assign \new_[12184]_  = ~A299 & ~A298;
  assign \new_[12185]_  = ~A267 & \new_[12184]_ ;
  assign \new_[12186]_  = \new_[12185]_  & \new_[12180]_ ;
  assign \new_[12189]_  = A166 & A168;
  assign \new_[12193]_  = ~A232 & A200;
  assign \new_[12194]_  = A199 & \new_[12193]_ ;
  assign \new_[12195]_  = \new_[12194]_  & \new_[12189]_ ;
  assign \new_[12198]_  = ~A265 & ~A233;
  assign \new_[12202]_  = ~A300 & A298;
  assign \new_[12203]_  = ~A266 & \new_[12202]_ ;
  assign \new_[12204]_  = \new_[12203]_  & \new_[12198]_ ;
  assign \new_[12207]_  = A166 & A168;
  assign \new_[12211]_  = ~A232 & A200;
  assign \new_[12212]_  = A199 & \new_[12211]_ ;
  assign \new_[12213]_  = \new_[12212]_  & \new_[12207]_ ;
  assign \new_[12216]_  = ~A265 & ~A233;
  assign \new_[12220]_  = A299 & A298;
  assign \new_[12221]_  = ~A266 & \new_[12220]_ ;
  assign \new_[12222]_  = \new_[12221]_  & \new_[12216]_ ;
  assign \new_[12225]_  = A166 & A168;
  assign \new_[12229]_  = ~A232 & A200;
  assign \new_[12230]_  = A199 & \new_[12229]_ ;
  assign \new_[12231]_  = \new_[12230]_  & \new_[12225]_ ;
  assign \new_[12234]_  = ~A265 & ~A233;
  assign \new_[12238]_  = ~A299 & ~A298;
  assign \new_[12239]_  = ~A266 & \new_[12238]_ ;
  assign \new_[12240]_  = \new_[12239]_  & \new_[12234]_ ;
  assign \new_[12243]_  = A166 & A168;
  assign \new_[12247]_  = A232 & ~A201;
  assign \new_[12248]_  = ~A200 & \new_[12247]_ ;
  assign \new_[12249]_  = \new_[12248]_  & \new_[12243]_ ;
  assign \new_[12252]_  = A265 & A233;
  assign \new_[12256]_  = ~A300 & ~A299;
  assign \new_[12257]_  = ~A267 & \new_[12256]_ ;
  assign \new_[12258]_  = \new_[12257]_  & \new_[12252]_ ;
  assign \new_[12261]_  = A166 & A168;
  assign \new_[12265]_  = A232 & ~A201;
  assign \new_[12266]_  = ~A200 & \new_[12265]_ ;
  assign \new_[12267]_  = \new_[12266]_  & \new_[12261]_ ;
  assign \new_[12270]_  = A265 & A233;
  assign \new_[12274]_  = A299 & A298;
  assign \new_[12275]_  = ~A267 & \new_[12274]_ ;
  assign \new_[12276]_  = \new_[12275]_  & \new_[12270]_ ;
  assign \new_[12279]_  = A166 & A168;
  assign \new_[12283]_  = A232 & ~A201;
  assign \new_[12284]_  = ~A200 & \new_[12283]_ ;
  assign \new_[12285]_  = \new_[12284]_  & \new_[12279]_ ;
  assign \new_[12288]_  = A265 & A233;
  assign \new_[12292]_  = ~A299 & ~A298;
  assign \new_[12293]_  = ~A267 & \new_[12292]_ ;
  assign \new_[12294]_  = \new_[12293]_  & \new_[12288]_ ;
  assign \new_[12297]_  = A166 & A168;
  assign \new_[12301]_  = A232 & ~A201;
  assign \new_[12302]_  = ~A200 & \new_[12301]_ ;
  assign \new_[12303]_  = \new_[12302]_  & \new_[12297]_ ;
  assign \new_[12306]_  = A265 & A233;
  assign \new_[12310]_  = ~A300 & ~A299;
  assign \new_[12311]_  = A266 & \new_[12310]_ ;
  assign \new_[12312]_  = \new_[12311]_  & \new_[12306]_ ;
  assign \new_[12315]_  = A166 & A168;
  assign \new_[12319]_  = A232 & ~A201;
  assign \new_[12320]_  = ~A200 & \new_[12319]_ ;
  assign \new_[12321]_  = \new_[12320]_  & \new_[12315]_ ;
  assign \new_[12324]_  = A265 & A233;
  assign \new_[12328]_  = A299 & A298;
  assign \new_[12329]_  = A266 & \new_[12328]_ ;
  assign \new_[12330]_  = \new_[12329]_  & \new_[12324]_ ;
  assign \new_[12333]_  = A166 & A168;
  assign \new_[12337]_  = A232 & ~A201;
  assign \new_[12338]_  = ~A200 & \new_[12337]_ ;
  assign \new_[12339]_  = \new_[12338]_  & \new_[12333]_ ;
  assign \new_[12342]_  = A265 & A233;
  assign \new_[12346]_  = ~A299 & ~A298;
  assign \new_[12347]_  = A266 & \new_[12346]_ ;
  assign \new_[12348]_  = \new_[12347]_  & \new_[12342]_ ;
  assign \new_[12351]_  = A166 & A168;
  assign \new_[12355]_  = A232 & ~A201;
  assign \new_[12356]_  = ~A200 & \new_[12355]_ ;
  assign \new_[12357]_  = \new_[12356]_  & \new_[12351]_ ;
  assign \new_[12360]_  = ~A265 & A233;
  assign \new_[12364]_  = ~A300 & ~A299;
  assign \new_[12365]_  = ~A266 & \new_[12364]_ ;
  assign \new_[12366]_  = \new_[12365]_  & \new_[12360]_ ;
  assign \new_[12369]_  = A166 & A168;
  assign \new_[12373]_  = A232 & ~A201;
  assign \new_[12374]_  = ~A200 & \new_[12373]_ ;
  assign \new_[12375]_  = \new_[12374]_  & \new_[12369]_ ;
  assign \new_[12378]_  = ~A265 & A233;
  assign \new_[12382]_  = A299 & A298;
  assign \new_[12383]_  = ~A266 & \new_[12382]_ ;
  assign \new_[12384]_  = \new_[12383]_  & \new_[12378]_ ;
  assign \new_[12387]_  = A166 & A168;
  assign \new_[12391]_  = A232 & ~A201;
  assign \new_[12392]_  = ~A200 & \new_[12391]_ ;
  assign \new_[12393]_  = \new_[12392]_  & \new_[12387]_ ;
  assign \new_[12396]_  = ~A265 & A233;
  assign \new_[12400]_  = ~A299 & ~A298;
  assign \new_[12401]_  = ~A266 & \new_[12400]_ ;
  assign \new_[12402]_  = \new_[12401]_  & \new_[12396]_ ;
  assign \new_[12405]_  = A166 & A168;
  assign \new_[12409]_  = ~A232 & ~A201;
  assign \new_[12410]_  = ~A200 & \new_[12409]_ ;
  assign \new_[12411]_  = \new_[12410]_  & \new_[12405]_ ;
  assign \new_[12414]_  = A298 & A233;
  assign \new_[12418]_  = A301 & A300;
  assign \new_[12419]_  = ~A299 & \new_[12418]_ ;
  assign \new_[12420]_  = \new_[12419]_  & \new_[12414]_ ;
  assign \new_[12423]_  = A166 & A168;
  assign \new_[12427]_  = ~A232 & ~A201;
  assign \new_[12428]_  = ~A200 & \new_[12427]_ ;
  assign \new_[12429]_  = \new_[12428]_  & \new_[12423]_ ;
  assign \new_[12432]_  = A298 & A233;
  assign \new_[12436]_  = A302 & A300;
  assign \new_[12437]_  = ~A299 & \new_[12436]_ ;
  assign \new_[12438]_  = \new_[12437]_  & \new_[12432]_ ;
  assign \new_[12441]_  = A166 & A168;
  assign \new_[12445]_  = ~A232 & ~A201;
  assign \new_[12446]_  = ~A200 & \new_[12445]_ ;
  assign \new_[12447]_  = \new_[12446]_  & \new_[12441]_ ;
  assign \new_[12450]_  = A265 & A233;
  assign \new_[12454]_  = A268 & A267;
  assign \new_[12455]_  = ~A266 & \new_[12454]_ ;
  assign \new_[12456]_  = \new_[12455]_  & \new_[12450]_ ;
  assign \new_[12459]_  = A166 & A168;
  assign \new_[12463]_  = ~A232 & ~A201;
  assign \new_[12464]_  = ~A200 & \new_[12463]_ ;
  assign \new_[12465]_  = \new_[12464]_  & \new_[12459]_ ;
  assign \new_[12468]_  = A265 & A233;
  assign \new_[12472]_  = A269 & A267;
  assign \new_[12473]_  = ~A266 & \new_[12472]_ ;
  assign \new_[12474]_  = \new_[12473]_  & \new_[12468]_ ;
  assign \new_[12477]_  = A166 & A168;
  assign \new_[12481]_  = ~A233 & ~A201;
  assign \new_[12482]_  = ~A200 & \new_[12481]_ ;
  assign \new_[12483]_  = \new_[12482]_  & \new_[12477]_ ;
  assign \new_[12486]_  = A265 & ~A234;
  assign \new_[12490]_  = ~A300 & A298;
  assign \new_[12491]_  = A266 & \new_[12490]_ ;
  assign \new_[12492]_  = \new_[12491]_  & \new_[12486]_ ;
  assign \new_[12495]_  = A166 & A168;
  assign \new_[12499]_  = ~A233 & ~A201;
  assign \new_[12500]_  = ~A200 & \new_[12499]_ ;
  assign \new_[12501]_  = \new_[12500]_  & \new_[12495]_ ;
  assign \new_[12504]_  = A265 & ~A234;
  assign \new_[12508]_  = A299 & A298;
  assign \new_[12509]_  = A266 & \new_[12508]_ ;
  assign \new_[12510]_  = \new_[12509]_  & \new_[12504]_ ;
  assign \new_[12513]_  = A166 & A168;
  assign \new_[12517]_  = ~A233 & ~A201;
  assign \new_[12518]_  = ~A200 & \new_[12517]_ ;
  assign \new_[12519]_  = \new_[12518]_  & \new_[12513]_ ;
  assign \new_[12522]_  = A265 & ~A234;
  assign \new_[12526]_  = ~A299 & ~A298;
  assign \new_[12527]_  = A266 & \new_[12526]_ ;
  assign \new_[12528]_  = \new_[12527]_  & \new_[12522]_ ;
  assign \new_[12531]_  = A166 & A168;
  assign \new_[12535]_  = ~A233 & ~A201;
  assign \new_[12536]_  = ~A200 & \new_[12535]_ ;
  assign \new_[12537]_  = \new_[12536]_  & \new_[12531]_ ;
  assign \new_[12540]_  = ~A266 & ~A234;
  assign \new_[12544]_  = ~A300 & A298;
  assign \new_[12545]_  = ~A267 & \new_[12544]_ ;
  assign \new_[12546]_  = \new_[12545]_  & \new_[12540]_ ;
  assign \new_[12549]_  = A166 & A168;
  assign \new_[12553]_  = ~A233 & ~A201;
  assign \new_[12554]_  = ~A200 & \new_[12553]_ ;
  assign \new_[12555]_  = \new_[12554]_  & \new_[12549]_ ;
  assign \new_[12558]_  = ~A266 & ~A234;
  assign \new_[12562]_  = A299 & A298;
  assign \new_[12563]_  = ~A267 & \new_[12562]_ ;
  assign \new_[12564]_  = \new_[12563]_  & \new_[12558]_ ;
  assign \new_[12567]_  = A166 & A168;
  assign \new_[12571]_  = ~A233 & ~A201;
  assign \new_[12572]_  = ~A200 & \new_[12571]_ ;
  assign \new_[12573]_  = \new_[12572]_  & \new_[12567]_ ;
  assign \new_[12576]_  = ~A266 & ~A234;
  assign \new_[12580]_  = ~A299 & ~A298;
  assign \new_[12581]_  = ~A267 & \new_[12580]_ ;
  assign \new_[12582]_  = \new_[12581]_  & \new_[12576]_ ;
  assign \new_[12585]_  = A166 & A168;
  assign \new_[12589]_  = ~A233 & ~A201;
  assign \new_[12590]_  = ~A200 & \new_[12589]_ ;
  assign \new_[12591]_  = \new_[12590]_  & \new_[12585]_ ;
  assign \new_[12594]_  = ~A265 & ~A234;
  assign \new_[12598]_  = ~A300 & A298;
  assign \new_[12599]_  = ~A266 & \new_[12598]_ ;
  assign \new_[12600]_  = \new_[12599]_  & \new_[12594]_ ;
  assign \new_[12603]_  = A166 & A168;
  assign \new_[12607]_  = ~A233 & ~A201;
  assign \new_[12608]_  = ~A200 & \new_[12607]_ ;
  assign \new_[12609]_  = \new_[12608]_  & \new_[12603]_ ;
  assign \new_[12612]_  = ~A265 & ~A234;
  assign \new_[12616]_  = A299 & A298;
  assign \new_[12617]_  = ~A266 & \new_[12616]_ ;
  assign \new_[12618]_  = \new_[12617]_  & \new_[12612]_ ;
  assign \new_[12621]_  = A166 & A168;
  assign \new_[12625]_  = ~A233 & ~A201;
  assign \new_[12626]_  = ~A200 & \new_[12625]_ ;
  assign \new_[12627]_  = \new_[12626]_  & \new_[12621]_ ;
  assign \new_[12630]_  = ~A265 & ~A234;
  assign \new_[12634]_  = ~A299 & ~A298;
  assign \new_[12635]_  = ~A266 & \new_[12634]_ ;
  assign \new_[12636]_  = \new_[12635]_  & \new_[12630]_ ;
  assign \new_[12639]_  = A166 & A168;
  assign \new_[12643]_  = A232 & ~A201;
  assign \new_[12644]_  = ~A200 & \new_[12643]_ ;
  assign \new_[12645]_  = \new_[12644]_  & \new_[12639]_ ;
  assign \new_[12648]_  = A234 & ~A233;
  assign \new_[12652]_  = A299 & ~A298;
  assign \new_[12653]_  = A235 & \new_[12652]_ ;
  assign \new_[12654]_  = \new_[12653]_  & \new_[12648]_ ;
  assign \new_[12657]_  = A166 & A168;
  assign \new_[12661]_  = A232 & ~A201;
  assign \new_[12662]_  = ~A200 & \new_[12661]_ ;
  assign \new_[12663]_  = \new_[12662]_  & \new_[12657]_ ;
  assign \new_[12666]_  = A234 & ~A233;
  assign \new_[12670]_  = A266 & ~A265;
  assign \new_[12671]_  = A235 & \new_[12670]_ ;
  assign \new_[12672]_  = \new_[12671]_  & \new_[12666]_ ;
  assign \new_[12675]_  = A166 & A168;
  assign \new_[12679]_  = A232 & ~A201;
  assign \new_[12680]_  = ~A200 & \new_[12679]_ ;
  assign \new_[12681]_  = \new_[12680]_  & \new_[12675]_ ;
  assign \new_[12684]_  = A234 & ~A233;
  assign \new_[12688]_  = A299 & ~A298;
  assign \new_[12689]_  = A236 & \new_[12688]_ ;
  assign \new_[12690]_  = \new_[12689]_  & \new_[12684]_ ;
  assign \new_[12693]_  = A166 & A168;
  assign \new_[12697]_  = A232 & ~A201;
  assign \new_[12698]_  = ~A200 & \new_[12697]_ ;
  assign \new_[12699]_  = \new_[12698]_  & \new_[12693]_ ;
  assign \new_[12702]_  = A234 & ~A233;
  assign \new_[12706]_  = A266 & ~A265;
  assign \new_[12707]_  = A236 & \new_[12706]_ ;
  assign \new_[12708]_  = \new_[12707]_  & \new_[12702]_ ;
  assign \new_[12711]_  = A166 & A168;
  assign \new_[12715]_  = ~A232 & ~A201;
  assign \new_[12716]_  = ~A200 & \new_[12715]_ ;
  assign \new_[12717]_  = \new_[12716]_  & \new_[12711]_ ;
  assign \new_[12720]_  = A265 & ~A233;
  assign \new_[12724]_  = ~A300 & A298;
  assign \new_[12725]_  = A266 & \new_[12724]_ ;
  assign \new_[12726]_  = \new_[12725]_  & \new_[12720]_ ;
  assign \new_[12729]_  = A166 & A168;
  assign \new_[12733]_  = ~A232 & ~A201;
  assign \new_[12734]_  = ~A200 & \new_[12733]_ ;
  assign \new_[12735]_  = \new_[12734]_  & \new_[12729]_ ;
  assign \new_[12738]_  = A265 & ~A233;
  assign \new_[12742]_  = A299 & A298;
  assign \new_[12743]_  = A266 & \new_[12742]_ ;
  assign \new_[12744]_  = \new_[12743]_  & \new_[12738]_ ;
  assign \new_[12747]_  = A166 & A168;
  assign \new_[12751]_  = ~A232 & ~A201;
  assign \new_[12752]_  = ~A200 & \new_[12751]_ ;
  assign \new_[12753]_  = \new_[12752]_  & \new_[12747]_ ;
  assign \new_[12756]_  = A265 & ~A233;
  assign \new_[12760]_  = ~A299 & ~A298;
  assign \new_[12761]_  = A266 & \new_[12760]_ ;
  assign \new_[12762]_  = \new_[12761]_  & \new_[12756]_ ;
  assign \new_[12765]_  = A166 & A168;
  assign \new_[12769]_  = ~A232 & ~A201;
  assign \new_[12770]_  = ~A200 & \new_[12769]_ ;
  assign \new_[12771]_  = \new_[12770]_  & \new_[12765]_ ;
  assign \new_[12774]_  = ~A266 & ~A233;
  assign \new_[12778]_  = ~A300 & A298;
  assign \new_[12779]_  = ~A267 & \new_[12778]_ ;
  assign \new_[12780]_  = \new_[12779]_  & \new_[12774]_ ;
  assign \new_[12783]_  = A166 & A168;
  assign \new_[12787]_  = ~A232 & ~A201;
  assign \new_[12788]_  = ~A200 & \new_[12787]_ ;
  assign \new_[12789]_  = \new_[12788]_  & \new_[12783]_ ;
  assign \new_[12792]_  = ~A266 & ~A233;
  assign \new_[12796]_  = A299 & A298;
  assign \new_[12797]_  = ~A267 & \new_[12796]_ ;
  assign \new_[12798]_  = \new_[12797]_  & \new_[12792]_ ;
  assign \new_[12801]_  = A166 & A168;
  assign \new_[12805]_  = ~A232 & ~A201;
  assign \new_[12806]_  = ~A200 & \new_[12805]_ ;
  assign \new_[12807]_  = \new_[12806]_  & \new_[12801]_ ;
  assign \new_[12810]_  = ~A266 & ~A233;
  assign \new_[12814]_  = ~A299 & ~A298;
  assign \new_[12815]_  = ~A267 & \new_[12814]_ ;
  assign \new_[12816]_  = \new_[12815]_  & \new_[12810]_ ;
  assign \new_[12819]_  = A166 & A168;
  assign \new_[12823]_  = ~A232 & ~A201;
  assign \new_[12824]_  = ~A200 & \new_[12823]_ ;
  assign \new_[12825]_  = \new_[12824]_  & \new_[12819]_ ;
  assign \new_[12828]_  = ~A265 & ~A233;
  assign \new_[12832]_  = ~A300 & A298;
  assign \new_[12833]_  = ~A266 & \new_[12832]_ ;
  assign \new_[12834]_  = \new_[12833]_  & \new_[12828]_ ;
  assign \new_[12837]_  = A166 & A168;
  assign \new_[12841]_  = ~A232 & ~A201;
  assign \new_[12842]_  = ~A200 & \new_[12841]_ ;
  assign \new_[12843]_  = \new_[12842]_  & \new_[12837]_ ;
  assign \new_[12846]_  = ~A265 & ~A233;
  assign \new_[12850]_  = A299 & A298;
  assign \new_[12851]_  = ~A266 & \new_[12850]_ ;
  assign \new_[12852]_  = \new_[12851]_  & \new_[12846]_ ;
  assign \new_[12855]_  = A166 & A168;
  assign \new_[12859]_  = ~A232 & ~A201;
  assign \new_[12860]_  = ~A200 & \new_[12859]_ ;
  assign \new_[12861]_  = \new_[12860]_  & \new_[12855]_ ;
  assign \new_[12864]_  = ~A265 & ~A233;
  assign \new_[12868]_  = ~A299 & ~A298;
  assign \new_[12869]_  = ~A266 & \new_[12868]_ ;
  assign \new_[12870]_  = \new_[12869]_  & \new_[12864]_ ;
  assign \new_[12873]_  = A166 & A168;
  assign \new_[12877]_  = A232 & ~A200;
  assign \new_[12878]_  = ~A199 & \new_[12877]_ ;
  assign \new_[12879]_  = \new_[12878]_  & \new_[12873]_ ;
  assign \new_[12882]_  = A265 & A233;
  assign \new_[12886]_  = ~A300 & ~A299;
  assign \new_[12887]_  = ~A267 & \new_[12886]_ ;
  assign \new_[12888]_  = \new_[12887]_  & \new_[12882]_ ;
  assign \new_[12891]_  = A166 & A168;
  assign \new_[12895]_  = A232 & ~A200;
  assign \new_[12896]_  = ~A199 & \new_[12895]_ ;
  assign \new_[12897]_  = \new_[12896]_  & \new_[12891]_ ;
  assign \new_[12900]_  = A265 & A233;
  assign \new_[12904]_  = A299 & A298;
  assign \new_[12905]_  = ~A267 & \new_[12904]_ ;
  assign \new_[12906]_  = \new_[12905]_  & \new_[12900]_ ;
  assign \new_[12909]_  = A166 & A168;
  assign \new_[12913]_  = A232 & ~A200;
  assign \new_[12914]_  = ~A199 & \new_[12913]_ ;
  assign \new_[12915]_  = \new_[12914]_  & \new_[12909]_ ;
  assign \new_[12918]_  = A265 & A233;
  assign \new_[12922]_  = ~A299 & ~A298;
  assign \new_[12923]_  = ~A267 & \new_[12922]_ ;
  assign \new_[12924]_  = \new_[12923]_  & \new_[12918]_ ;
  assign \new_[12927]_  = A166 & A168;
  assign \new_[12931]_  = A232 & ~A200;
  assign \new_[12932]_  = ~A199 & \new_[12931]_ ;
  assign \new_[12933]_  = \new_[12932]_  & \new_[12927]_ ;
  assign \new_[12936]_  = A265 & A233;
  assign \new_[12940]_  = ~A300 & ~A299;
  assign \new_[12941]_  = A266 & \new_[12940]_ ;
  assign \new_[12942]_  = \new_[12941]_  & \new_[12936]_ ;
  assign \new_[12945]_  = A166 & A168;
  assign \new_[12949]_  = A232 & ~A200;
  assign \new_[12950]_  = ~A199 & \new_[12949]_ ;
  assign \new_[12951]_  = \new_[12950]_  & \new_[12945]_ ;
  assign \new_[12954]_  = A265 & A233;
  assign \new_[12958]_  = A299 & A298;
  assign \new_[12959]_  = A266 & \new_[12958]_ ;
  assign \new_[12960]_  = \new_[12959]_  & \new_[12954]_ ;
  assign \new_[12963]_  = A166 & A168;
  assign \new_[12967]_  = A232 & ~A200;
  assign \new_[12968]_  = ~A199 & \new_[12967]_ ;
  assign \new_[12969]_  = \new_[12968]_  & \new_[12963]_ ;
  assign \new_[12972]_  = A265 & A233;
  assign \new_[12976]_  = ~A299 & ~A298;
  assign \new_[12977]_  = A266 & \new_[12976]_ ;
  assign \new_[12978]_  = \new_[12977]_  & \new_[12972]_ ;
  assign \new_[12981]_  = A166 & A168;
  assign \new_[12985]_  = A232 & ~A200;
  assign \new_[12986]_  = ~A199 & \new_[12985]_ ;
  assign \new_[12987]_  = \new_[12986]_  & \new_[12981]_ ;
  assign \new_[12990]_  = ~A265 & A233;
  assign \new_[12994]_  = ~A300 & ~A299;
  assign \new_[12995]_  = ~A266 & \new_[12994]_ ;
  assign \new_[12996]_  = \new_[12995]_  & \new_[12990]_ ;
  assign \new_[12999]_  = A166 & A168;
  assign \new_[13003]_  = A232 & ~A200;
  assign \new_[13004]_  = ~A199 & \new_[13003]_ ;
  assign \new_[13005]_  = \new_[13004]_  & \new_[12999]_ ;
  assign \new_[13008]_  = ~A265 & A233;
  assign \new_[13012]_  = A299 & A298;
  assign \new_[13013]_  = ~A266 & \new_[13012]_ ;
  assign \new_[13014]_  = \new_[13013]_  & \new_[13008]_ ;
  assign \new_[13017]_  = A166 & A168;
  assign \new_[13021]_  = A232 & ~A200;
  assign \new_[13022]_  = ~A199 & \new_[13021]_ ;
  assign \new_[13023]_  = \new_[13022]_  & \new_[13017]_ ;
  assign \new_[13026]_  = ~A265 & A233;
  assign \new_[13030]_  = ~A299 & ~A298;
  assign \new_[13031]_  = ~A266 & \new_[13030]_ ;
  assign \new_[13032]_  = \new_[13031]_  & \new_[13026]_ ;
  assign \new_[13035]_  = A166 & A168;
  assign \new_[13039]_  = ~A232 & ~A200;
  assign \new_[13040]_  = ~A199 & \new_[13039]_ ;
  assign \new_[13041]_  = \new_[13040]_  & \new_[13035]_ ;
  assign \new_[13044]_  = A298 & A233;
  assign \new_[13048]_  = A301 & A300;
  assign \new_[13049]_  = ~A299 & \new_[13048]_ ;
  assign \new_[13050]_  = \new_[13049]_  & \new_[13044]_ ;
  assign \new_[13053]_  = A166 & A168;
  assign \new_[13057]_  = ~A232 & ~A200;
  assign \new_[13058]_  = ~A199 & \new_[13057]_ ;
  assign \new_[13059]_  = \new_[13058]_  & \new_[13053]_ ;
  assign \new_[13062]_  = A298 & A233;
  assign \new_[13066]_  = A302 & A300;
  assign \new_[13067]_  = ~A299 & \new_[13066]_ ;
  assign \new_[13068]_  = \new_[13067]_  & \new_[13062]_ ;
  assign \new_[13071]_  = A166 & A168;
  assign \new_[13075]_  = ~A232 & ~A200;
  assign \new_[13076]_  = ~A199 & \new_[13075]_ ;
  assign \new_[13077]_  = \new_[13076]_  & \new_[13071]_ ;
  assign \new_[13080]_  = A265 & A233;
  assign \new_[13084]_  = A268 & A267;
  assign \new_[13085]_  = ~A266 & \new_[13084]_ ;
  assign \new_[13086]_  = \new_[13085]_  & \new_[13080]_ ;
  assign \new_[13089]_  = A166 & A168;
  assign \new_[13093]_  = ~A232 & ~A200;
  assign \new_[13094]_  = ~A199 & \new_[13093]_ ;
  assign \new_[13095]_  = \new_[13094]_  & \new_[13089]_ ;
  assign \new_[13098]_  = A265 & A233;
  assign \new_[13102]_  = A269 & A267;
  assign \new_[13103]_  = ~A266 & \new_[13102]_ ;
  assign \new_[13104]_  = \new_[13103]_  & \new_[13098]_ ;
  assign \new_[13107]_  = A166 & A168;
  assign \new_[13111]_  = ~A233 & ~A200;
  assign \new_[13112]_  = ~A199 & \new_[13111]_ ;
  assign \new_[13113]_  = \new_[13112]_  & \new_[13107]_ ;
  assign \new_[13116]_  = A265 & ~A234;
  assign \new_[13120]_  = ~A300 & A298;
  assign \new_[13121]_  = A266 & \new_[13120]_ ;
  assign \new_[13122]_  = \new_[13121]_  & \new_[13116]_ ;
  assign \new_[13125]_  = A166 & A168;
  assign \new_[13129]_  = ~A233 & ~A200;
  assign \new_[13130]_  = ~A199 & \new_[13129]_ ;
  assign \new_[13131]_  = \new_[13130]_  & \new_[13125]_ ;
  assign \new_[13134]_  = A265 & ~A234;
  assign \new_[13138]_  = A299 & A298;
  assign \new_[13139]_  = A266 & \new_[13138]_ ;
  assign \new_[13140]_  = \new_[13139]_  & \new_[13134]_ ;
  assign \new_[13143]_  = A166 & A168;
  assign \new_[13147]_  = ~A233 & ~A200;
  assign \new_[13148]_  = ~A199 & \new_[13147]_ ;
  assign \new_[13149]_  = \new_[13148]_  & \new_[13143]_ ;
  assign \new_[13152]_  = A265 & ~A234;
  assign \new_[13156]_  = ~A299 & ~A298;
  assign \new_[13157]_  = A266 & \new_[13156]_ ;
  assign \new_[13158]_  = \new_[13157]_  & \new_[13152]_ ;
  assign \new_[13161]_  = A166 & A168;
  assign \new_[13165]_  = ~A233 & ~A200;
  assign \new_[13166]_  = ~A199 & \new_[13165]_ ;
  assign \new_[13167]_  = \new_[13166]_  & \new_[13161]_ ;
  assign \new_[13170]_  = ~A266 & ~A234;
  assign \new_[13174]_  = ~A300 & A298;
  assign \new_[13175]_  = ~A267 & \new_[13174]_ ;
  assign \new_[13176]_  = \new_[13175]_  & \new_[13170]_ ;
  assign \new_[13179]_  = A166 & A168;
  assign \new_[13183]_  = ~A233 & ~A200;
  assign \new_[13184]_  = ~A199 & \new_[13183]_ ;
  assign \new_[13185]_  = \new_[13184]_  & \new_[13179]_ ;
  assign \new_[13188]_  = ~A266 & ~A234;
  assign \new_[13192]_  = A299 & A298;
  assign \new_[13193]_  = ~A267 & \new_[13192]_ ;
  assign \new_[13194]_  = \new_[13193]_  & \new_[13188]_ ;
  assign \new_[13197]_  = A166 & A168;
  assign \new_[13201]_  = ~A233 & ~A200;
  assign \new_[13202]_  = ~A199 & \new_[13201]_ ;
  assign \new_[13203]_  = \new_[13202]_  & \new_[13197]_ ;
  assign \new_[13206]_  = ~A266 & ~A234;
  assign \new_[13210]_  = ~A299 & ~A298;
  assign \new_[13211]_  = ~A267 & \new_[13210]_ ;
  assign \new_[13212]_  = \new_[13211]_  & \new_[13206]_ ;
  assign \new_[13215]_  = A166 & A168;
  assign \new_[13219]_  = ~A233 & ~A200;
  assign \new_[13220]_  = ~A199 & \new_[13219]_ ;
  assign \new_[13221]_  = \new_[13220]_  & \new_[13215]_ ;
  assign \new_[13224]_  = ~A265 & ~A234;
  assign \new_[13228]_  = ~A300 & A298;
  assign \new_[13229]_  = ~A266 & \new_[13228]_ ;
  assign \new_[13230]_  = \new_[13229]_  & \new_[13224]_ ;
  assign \new_[13233]_  = A166 & A168;
  assign \new_[13237]_  = ~A233 & ~A200;
  assign \new_[13238]_  = ~A199 & \new_[13237]_ ;
  assign \new_[13239]_  = \new_[13238]_  & \new_[13233]_ ;
  assign \new_[13242]_  = ~A265 & ~A234;
  assign \new_[13246]_  = A299 & A298;
  assign \new_[13247]_  = ~A266 & \new_[13246]_ ;
  assign \new_[13248]_  = \new_[13247]_  & \new_[13242]_ ;
  assign \new_[13251]_  = A166 & A168;
  assign \new_[13255]_  = ~A233 & ~A200;
  assign \new_[13256]_  = ~A199 & \new_[13255]_ ;
  assign \new_[13257]_  = \new_[13256]_  & \new_[13251]_ ;
  assign \new_[13260]_  = ~A265 & ~A234;
  assign \new_[13264]_  = ~A299 & ~A298;
  assign \new_[13265]_  = ~A266 & \new_[13264]_ ;
  assign \new_[13266]_  = \new_[13265]_  & \new_[13260]_ ;
  assign \new_[13269]_  = A166 & A168;
  assign \new_[13273]_  = A232 & ~A200;
  assign \new_[13274]_  = ~A199 & \new_[13273]_ ;
  assign \new_[13275]_  = \new_[13274]_  & \new_[13269]_ ;
  assign \new_[13278]_  = A234 & ~A233;
  assign \new_[13282]_  = A299 & ~A298;
  assign \new_[13283]_  = A235 & \new_[13282]_ ;
  assign \new_[13284]_  = \new_[13283]_  & \new_[13278]_ ;
  assign \new_[13287]_  = A166 & A168;
  assign \new_[13291]_  = A232 & ~A200;
  assign \new_[13292]_  = ~A199 & \new_[13291]_ ;
  assign \new_[13293]_  = \new_[13292]_  & \new_[13287]_ ;
  assign \new_[13296]_  = A234 & ~A233;
  assign \new_[13300]_  = A266 & ~A265;
  assign \new_[13301]_  = A235 & \new_[13300]_ ;
  assign \new_[13302]_  = \new_[13301]_  & \new_[13296]_ ;
  assign \new_[13305]_  = A166 & A168;
  assign \new_[13309]_  = A232 & ~A200;
  assign \new_[13310]_  = ~A199 & \new_[13309]_ ;
  assign \new_[13311]_  = \new_[13310]_  & \new_[13305]_ ;
  assign \new_[13314]_  = A234 & ~A233;
  assign \new_[13318]_  = A299 & ~A298;
  assign \new_[13319]_  = A236 & \new_[13318]_ ;
  assign \new_[13320]_  = \new_[13319]_  & \new_[13314]_ ;
  assign \new_[13323]_  = A166 & A168;
  assign \new_[13327]_  = A232 & ~A200;
  assign \new_[13328]_  = ~A199 & \new_[13327]_ ;
  assign \new_[13329]_  = \new_[13328]_  & \new_[13323]_ ;
  assign \new_[13332]_  = A234 & ~A233;
  assign \new_[13336]_  = A266 & ~A265;
  assign \new_[13337]_  = A236 & \new_[13336]_ ;
  assign \new_[13338]_  = \new_[13337]_  & \new_[13332]_ ;
  assign \new_[13341]_  = A166 & A168;
  assign \new_[13345]_  = ~A232 & ~A200;
  assign \new_[13346]_  = ~A199 & \new_[13345]_ ;
  assign \new_[13347]_  = \new_[13346]_  & \new_[13341]_ ;
  assign \new_[13350]_  = A265 & ~A233;
  assign \new_[13354]_  = ~A300 & A298;
  assign \new_[13355]_  = A266 & \new_[13354]_ ;
  assign \new_[13356]_  = \new_[13355]_  & \new_[13350]_ ;
  assign \new_[13359]_  = A166 & A168;
  assign \new_[13363]_  = ~A232 & ~A200;
  assign \new_[13364]_  = ~A199 & \new_[13363]_ ;
  assign \new_[13365]_  = \new_[13364]_  & \new_[13359]_ ;
  assign \new_[13368]_  = A265 & ~A233;
  assign \new_[13372]_  = A299 & A298;
  assign \new_[13373]_  = A266 & \new_[13372]_ ;
  assign \new_[13374]_  = \new_[13373]_  & \new_[13368]_ ;
  assign \new_[13377]_  = A166 & A168;
  assign \new_[13381]_  = ~A232 & ~A200;
  assign \new_[13382]_  = ~A199 & \new_[13381]_ ;
  assign \new_[13383]_  = \new_[13382]_  & \new_[13377]_ ;
  assign \new_[13386]_  = A265 & ~A233;
  assign \new_[13390]_  = ~A299 & ~A298;
  assign \new_[13391]_  = A266 & \new_[13390]_ ;
  assign \new_[13392]_  = \new_[13391]_  & \new_[13386]_ ;
  assign \new_[13395]_  = A166 & A168;
  assign \new_[13399]_  = ~A232 & ~A200;
  assign \new_[13400]_  = ~A199 & \new_[13399]_ ;
  assign \new_[13401]_  = \new_[13400]_  & \new_[13395]_ ;
  assign \new_[13404]_  = ~A266 & ~A233;
  assign \new_[13408]_  = ~A300 & A298;
  assign \new_[13409]_  = ~A267 & \new_[13408]_ ;
  assign \new_[13410]_  = \new_[13409]_  & \new_[13404]_ ;
  assign \new_[13413]_  = A166 & A168;
  assign \new_[13417]_  = ~A232 & ~A200;
  assign \new_[13418]_  = ~A199 & \new_[13417]_ ;
  assign \new_[13419]_  = \new_[13418]_  & \new_[13413]_ ;
  assign \new_[13422]_  = ~A266 & ~A233;
  assign \new_[13426]_  = A299 & A298;
  assign \new_[13427]_  = ~A267 & \new_[13426]_ ;
  assign \new_[13428]_  = \new_[13427]_  & \new_[13422]_ ;
  assign \new_[13431]_  = A166 & A168;
  assign \new_[13435]_  = ~A232 & ~A200;
  assign \new_[13436]_  = ~A199 & \new_[13435]_ ;
  assign \new_[13437]_  = \new_[13436]_  & \new_[13431]_ ;
  assign \new_[13440]_  = ~A266 & ~A233;
  assign \new_[13444]_  = ~A299 & ~A298;
  assign \new_[13445]_  = ~A267 & \new_[13444]_ ;
  assign \new_[13446]_  = \new_[13445]_  & \new_[13440]_ ;
  assign \new_[13449]_  = A166 & A168;
  assign \new_[13453]_  = ~A232 & ~A200;
  assign \new_[13454]_  = ~A199 & \new_[13453]_ ;
  assign \new_[13455]_  = \new_[13454]_  & \new_[13449]_ ;
  assign \new_[13458]_  = ~A265 & ~A233;
  assign \new_[13462]_  = ~A300 & A298;
  assign \new_[13463]_  = ~A266 & \new_[13462]_ ;
  assign \new_[13464]_  = \new_[13463]_  & \new_[13458]_ ;
  assign \new_[13467]_  = A166 & A168;
  assign \new_[13471]_  = ~A232 & ~A200;
  assign \new_[13472]_  = ~A199 & \new_[13471]_ ;
  assign \new_[13473]_  = \new_[13472]_  & \new_[13467]_ ;
  assign \new_[13476]_  = ~A265 & ~A233;
  assign \new_[13480]_  = A299 & A298;
  assign \new_[13481]_  = ~A266 & \new_[13480]_ ;
  assign \new_[13482]_  = \new_[13481]_  & \new_[13476]_ ;
  assign \new_[13485]_  = A166 & A168;
  assign \new_[13489]_  = ~A232 & ~A200;
  assign \new_[13490]_  = ~A199 & \new_[13489]_ ;
  assign \new_[13491]_  = \new_[13490]_  & \new_[13485]_ ;
  assign \new_[13494]_  = ~A265 & ~A233;
  assign \new_[13498]_  = ~A299 & ~A298;
  assign \new_[13499]_  = ~A266 & \new_[13498]_ ;
  assign \new_[13500]_  = \new_[13499]_  & \new_[13494]_ ;
  assign \new_[13503]_  = A167 & A168;
  assign \new_[13507]_  = A232 & A200;
  assign \new_[13508]_  = A199 & \new_[13507]_ ;
  assign \new_[13509]_  = \new_[13508]_  & \new_[13503]_ ;
  assign \new_[13512]_  = A265 & A233;
  assign \new_[13516]_  = ~A300 & ~A299;
  assign \new_[13517]_  = ~A267 & \new_[13516]_ ;
  assign \new_[13518]_  = \new_[13517]_  & \new_[13512]_ ;
  assign \new_[13521]_  = A167 & A168;
  assign \new_[13525]_  = A232 & A200;
  assign \new_[13526]_  = A199 & \new_[13525]_ ;
  assign \new_[13527]_  = \new_[13526]_  & \new_[13521]_ ;
  assign \new_[13530]_  = A265 & A233;
  assign \new_[13534]_  = A299 & A298;
  assign \new_[13535]_  = ~A267 & \new_[13534]_ ;
  assign \new_[13536]_  = \new_[13535]_  & \new_[13530]_ ;
  assign \new_[13539]_  = A167 & A168;
  assign \new_[13543]_  = A232 & A200;
  assign \new_[13544]_  = A199 & \new_[13543]_ ;
  assign \new_[13545]_  = \new_[13544]_  & \new_[13539]_ ;
  assign \new_[13548]_  = A265 & A233;
  assign \new_[13552]_  = ~A299 & ~A298;
  assign \new_[13553]_  = ~A267 & \new_[13552]_ ;
  assign \new_[13554]_  = \new_[13553]_  & \new_[13548]_ ;
  assign \new_[13557]_  = A167 & A168;
  assign \new_[13561]_  = A232 & A200;
  assign \new_[13562]_  = A199 & \new_[13561]_ ;
  assign \new_[13563]_  = \new_[13562]_  & \new_[13557]_ ;
  assign \new_[13566]_  = A265 & A233;
  assign \new_[13570]_  = ~A300 & ~A299;
  assign \new_[13571]_  = A266 & \new_[13570]_ ;
  assign \new_[13572]_  = \new_[13571]_  & \new_[13566]_ ;
  assign \new_[13575]_  = A167 & A168;
  assign \new_[13579]_  = A232 & A200;
  assign \new_[13580]_  = A199 & \new_[13579]_ ;
  assign \new_[13581]_  = \new_[13580]_  & \new_[13575]_ ;
  assign \new_[13584]_  = A265 & A233;
  assign \new_[13588]_  = A299 & A298;
  assign \new_[13589]_  = A266 & \new_[13588]_ ;
  assign \new_[13590]_  = \new_[13589]_  & \new_[13584]_ ;
  assign \new_[13593]_  = A167 & A168;
  assign \new_[13597]_  = A232 & A200;
  assign \new_[13598]_  = A199 & \new_[13597]_ ;
  assign \new_[13599]_  = \new_[13598]_  & \new_[13593]_ ;
  assign \new_[13602]_  = A265 & A233;
  assign \new_[13606]_  = ~A299 & ~A298;
  assign \new_[13607]_  = A266 & \new_[13606]_ ;
  assign \new_[13608]_  = \new_[13607]_  & \new_[13602]_ ;
  assign \new_[13611]_  = A167 & A168;
  assign \new_[13615]_  = A232 & A200;
  assign \new_[13616]_  = A199 & \new_[13615]_ ;
  assign \new_[13617]_  = \new_[13616]_  & \new_[13611]_ ;
  assign \new_[13620]_  = ~A265 & A233;
  assign \new_[13624]_  = ~A300 & ~A299;
  assign \new_[13625]_  = ~A266 & \new_[13624]_ ;
  assign \new_[13626]_  = \new_[13625]_  & \new_[13620]_ ;
  assign \new_[13629]_  = A167 & A168;
  assign \new_[13633]_  = A232 & A200;
  assign \new_[13634]_  = A199 & \new_[13633]_ ;
  assign \new_[13635]_  = \new_[13634]_  & \new_[13629]_ ;
  assign \new_[13638]_  = ~A265 & A233;
  assign \new_[13642]_  = A299 & A298;
  assign \new_[13643]_  = ~A266 & \new_[13642]_ ;
  assign \new_[13644]_  = \new_[13643]_  & \new_[13638]_ ;
  assign \new_[13647]_  = A167 & A168;
  assign \new_[13651]_  = A232 & A200;
  assign \new_[13652]_  = A199 & \new_[13651]_ ;
  assign \new_[13653]_  = \new_[13652]_  & \new_[13647]_ ;
  assign \new_[13656]_  = ~A265 & A233;
  assign \new_[13660]_  = ~A299 & ~A298;
  assign \new_[13661]_  = ~A266 & \new_[13660]_ ;
  assign \new_[13662]_  = \new_[13661]_  & \new_[13656]_ ;
  assign \new_[13665]_  = A167 & A168;
  assign \new_[13669]_  = ~A232 & A200;
  assign \new_[13670]_  = A199 & \new_[13669]_ ;
  assign \new_[13671]_  = \new_[13670]_  & \new_[13665]_ ;
  assign \new_[13674]_  = A298 & A233;
  assign \new_[13678]_  = A301 & A300;
  assign \new_[13679]_  = ~A299 & \new_[13678]_ ;
  assign \new_[13680]_  = \new_[13679]_  & \new_[13674]_ ;
  assign \new_[13683]_  = A167 & A168;
  assign \new_[13687]_  = ~A232 & A200;
  assign \new_[13688]_  = A199 & \new_[13687]_ ;
  assign \new_[13689]_  = \new_[13688]_  & \new_[13683]_ ;
  assign \new_[13692]_  = A298 & A233;
  assign \new_[13696]_  = A302 & A300;
  assign \new_[13697]_  = ~A299 & \new_[13696]_ ;
  assign \new_[13698]_  = \new_[13697]_  & \new_[13692]_ ;
  assign \new_[13701]_  = A167 & A168;
  assign \new_[13705]_  = ~A232 & A200;
  assign \new_[13706]_  = A199 & \new_[13705]_ ;
  assign \new_[13707]_  = \new_[13706]_  & \new_[13701]_ ;
  assign \new_[13710]_  = A265 & A233;
  assign \new_[13714]_  = A268 & A267;
  assign \new_[13715]_  = ~A266 & \new_[13714]_ ;
  assign \new_[13716]_  = \new_[13715]_  & \new_[13710]_ ;
  assign \new_[13719]_  = A167 & A168;
  assign \new_[13723]_  = ~A232 & A200;
  assign \new_[13724]_  = A199 & \new_[13723]_ ;
  assign \new_[13725]_  = \new_[13724]_  & \new_[13719]_ ;
  assign \new_[13728]_  = A265 & A233;
  assign \new_[13732]_  = A269 & A267;
  assign \new_[13733]_  = ~A266 & \new_[13732]_ ;
  assign \new_[13734]_  = \new_[13733]_  & \new_[13728]_ ;
  assign \new_[13737]_  = A167 & A168;
  assign \new_[13741]_  = ~A233 & A200;
  assign \new_[13742]_  = A199 & \new_[13741]_ ;
  assign \new_[13743]_  = \new_[13742]_  & \new_[13737]_ ;
  assign \new_[13746]_  = A265 & ~A234;
  assign \new_[13750]_  = ~A300 & A298;
  assign \new_[13751]_  = A266 & \new_[13750]_ ;
  assign \new_[13752]_  = \new_[13751]_  & \new_[13746]_ ;
  assign \new_[13755]_  = A167 & A168;
  assign \new_[13759]_  = ~A233 & A200;
  assign \new_[13760]_  = A199 & \new_[13759]_ ;
  assign \new_[13761]_  = \new_[13760]_  & \new_[13755]_ ;
  assign \new_[13764]_  = A265 & ~A234;
  assign \new_[13768]_  = A299 & A298;
  assign \new_[13769]_  = A266 & \new_[13768]_ ;
  assign \new_[13770]_  = \new_[13769]_  & \new_[13764]_ ;
  assign \new_[13773]_  = A167 & A168;
  assign \new_[13777]_  = ~A233 & A200;
  assign \new_[13778]_  = A199 & \new_[13777]_ ;
  assign \new_[13779]_  = \new_[13778]_  & \new_[13773]_ ;
  assign \new_[13782]_  = A265 & ~A234;
  assign \new_[13786]_  = ~A299 & ~A298;
  assign \new_[13787]_  = A266 & \new_[13786]_ ;
  assign \new_[13788]_  = \new_[13787]_  & \new_[13782]_ ;
  assign \new_[13791]_  = A167 & A168;
  assign \new_[13795]_  = ~A233 & A200;
  assign \new_[13796]_  = A199 & \new_[13795]_ ;
  assign \new_[13797]_  = \new_[13796]_  & \new_[13791]_ ;
  assign \new_[13800]_  = ~A266 & ~A234;
  assign \new_[13804]_  = ~A300 & A298;
  assign \new_[13805]_  = ~A267 & \new_[13804]_ ;
  assign \new_[13806]_  = \new_[13805]_  & \new_[13800]_ ;
  assign \new_[13809]_  = A167 & A168;
  assign \new_[13813]_  = ~A233 & A200;
  assign \new_[13814]_  = A199 & \new_[13813]_ ;
  assign \new_[13815]_  = \new_[13814]_  & \new_[13809]_ ;
  assign \new_[13818]_  = ~A266 & ~A234;
  assign \new_[13822]_  = A299 & A298;
  assign \new_[13823]_  = ~A267 & \new_[13822]_ ;
  assign \new_[13824]_  = \new_[13823]_  & \new_[13818]_ ;
  assign \new_[13827]_  = A167 & A168;
  assign \new_[13831]_  = ~A233 & A200;
  assign \new_[13832]_  = A199 & \new_[13831]_ ;
  assign \new_[13833]_  = \new_[13832]_  & \new_[13827]_ ;
  assign \new_[13836]_  = ~A266 & ~A234;
  assign \new_[13840]_  = ~A299 & ~A298;
  assign \new_[13841]_  = ~A267 & \new_[13840]_ ;
  assign \new_[13842]_  = \new_[13841]_  & \new_[13836]_ ;
  assign \new_[13845]_  = A167 & A168;
  assign \new_[13849]_  = ~A233 & A200;
  assign \new_[13850]_  = A199 & \new_[13849]_ ;
  assign \new_[13851]_  = \new_[13850]_  & \new_[13845]_ ;
  assign \new_[13854]_  = ~A265 & ~A234;
  assign \new_[13858]_  = ~A300 & A298;
  assign \new_[13859]_  = ~A266 & \new_[13858]_ ;
  assign \new_[13860]_  = \new_[13859]_  & \new_[13854]_ ;
  assign \new_[13863]_  = A167 & A168;
  assign \new_[13867]_  = ~A233 & A200;
  assign \new_[13868]_  = A199 & \new_[13867]_ ;
  assign \new_[13869]_  = \new_[13868]_  & \new_[13863]_ ;
  assign \new_[13872]_  = ~A265 & ~A234;
  assign \new_[13876]_  = A299 & A298;
  assign \new_[13877]_  = ~A266 & \new_[13876]_ ;
  assign \new_[13878]_  = \new_[13877]_  & \new_[13872]_ ;
  assign \new_[13881]_  = A167 & A168;
  assign \new_[13885]_  = ~A233 & A200;
  assign \new_[13886]_  = A199 & \new_[13885]_ ;
  assign \new_[13887]_  = \new_[13886]_  & \new_[13881]_ ;
  assign \new_[13890]_  = ~A265 & ~A234;
  assign \new_[13894]_  = ~A299 & ~A298;
  assign \new_[13895]_  = ~A266 & \new_[13894]_ ;
  assign \new_[13896]_  = \new_[13895]_  & \new_[13890]_ ;
  assign \new_[13899]_  = A167 & A168;
  assign \new_[13903]_  = A232 & A200;
  assign \new_[13904]_  = A199 & \new_[13903]_ ;
  assign \new_[13905]_  = \new_[13904]_  & \new_[13899]_ ;
  assign \new_[13908]_  = A234 & ~A233;
  assign \new_[13912]_  = A299 & ~A298;
  assign \new_[13913]_  = A235 & \new_[13912]_ ;
  assign \new_[13914]_  = \new_[13913]_  & \new_[13908]_ ;
  assign \new_[13917]_  = A167 & A168;
  assign \new_[13921]_  = A232 & A200;
  assign \new_[13922]_  = A199 & \new_[13921]_ ;
  assign \new_[13923]_  = \new_[13922]_  & \new_[13917]_ ;
  assign \new_[13926]_  = A234 & ~A233;
  assign \new_[13930]_  = A266 & ~A265;
  assign \new_[13931]_  = A235 & \new_[13930]_ ;
  assign \new_[13932]_  = \new_[13931]_  & \new_[13926]_ ;
  assign \new_[13935]_  = A167 & A168;
  assign \new_[13939]_  = A232 & A200;
  assign \new_[13940]_  = A199 & \new_[13939]_ ;
  assign \new_[13941]_  = \new_[13940]_  & \new_[13935]_ ;
  assign \new_[13944]_  = A234 & ~A233;
  assign \new_[13948]_  = A299 & ~A298;
  assign \new_[13949]_  = A236 & \new_[13948]_ ;
  assign \new_[13950]_  = \new_[13949]_  & \new_[13944]_ ;
  assign \new_[13953]_  = A167 & A168;
  assign \new_[13957]_  = A232 & A200;
  assign \new_[13958]_  = A199 & \new_[13957]_ ;
  assign \new_[13959]_  = \new_[13958]_  & \new_[13953]_ ;
  assign \new_[13962]_  = A234 & ~A233;
  assign \new_[13966]_  = A266 & ~A265;
  assign \new_[13967]_  = A236 & \new_[13966]_ ;
  assign \new_[13968]_  = \new_[13967]_  & \new_[13962]_ ;
  assign \new_[13971]_  = A167 & A168;
  assign \new_[13975]_  = ~A232 & A200;
  assign \new_[13976]_  = A199 & \new_[13975]_ ;
  assign \new_[13977]_  = \new_[13976]_  & \new_[13971]_ ;
  assign \new_[13980]_  = A265 & ~A233;
  assign \new_[13984]_  = ~A300 & A298;
  assign \new_[13985]_  = A266 & \new_[13984]_ ;
  assign \new_[13986]_  = \new_[13985]_  & \new_[13980]_ ;
  assign \new_[13989]_  = A167 & A168;
  assign \new_[13993]_  = ~A232 & A200;
  assign \new_[13994]_  = A199 & \new_[13993]_ ;
  assign \new_[13995]_  = \new_[13994]_  & \new_[13989]_ ;
  assign \new_[13998]_  = A265 & ~A233;
  assign \new_[14002]_  = A299 & A298;
  assign \new_[14003]_  = A266 & \new_[14002]_ ;
  assign \new_[14004]_  = \new_[14003]_  & \new_[13998]_ ;
  assign \new_[14007]_  = A167 & A168;
  assign \new_[14011]_  = ~A232 & A200;
  assign \new_[14012]_  = A199 & \new_[14011]_ ;
  assign \new_[14013]_  = \new_[14012]_  & \new_[14007]_ ;
  assign \new_[14016]_  = A265 & ~A233;
  assign \new_[14020]_  = ~A299 & ~A298;
  assign \new_[14021]_  = A266 & \new_[14020]_ ;
  assign \new_[14022]_  = \new_[14021]_  & \new_[14016]_ ;
  assign \new_[14025]_  = A167 & A168;
  assign \new_[14029]_  = ~A232 & A200;
  assign \new_[14030]_  = A199 & \new_[14029]_ ;
  assign \new_[14031]_  = \new_[14030]_  & \new_[14025]_ ;
  assign \new_[14034]_  = ~A266 & ~A233;
  assign \new_[14038]_  = ~A300 & A298;
  assign \new_[14039]_  = ~A267 & \new_[14038]_ ;
  assign \new_[14040]_  = \new_[14039]_  & \new_[14034]_ ;
  assign \new_[14043]_  = A167 & A168;
  assign \new_[14047]_  = ~A232 & A200;
  assign \new_[14048]_  = A199 & \new_[14047]_ ;
  assign \new_[14049]_  = \new_[14048]_  & \new_[14043]_ ;
  assign \new_[14052]_  = ~A266 & ~A233;
  assign \new_[14056]_  = A299 & A298;
  assign \new_[14057]_  = ~A267 & \new_[14056]_ ;
  assign \new_[14058]_  = \new_[14057]_  & \new_[14052]_ ;
  assign \new_[14061]_  = A167 & A168;
  assign \new_[14065]_  = ~A232 & A200;
  assign \new_[14066]_  = A199 & \new_[14065]_ ;
  assign \new_[14067]_  = \new_[14066]_  & \new_[14061]_ ;
  assign \new_[14070]_  = ~A266 & ~A233;
  assign \new_[14074]_  = ~A299 & ~A298;
  assign \new_[14075]_  = ~A267 & \new_[14074]_ ;
  assign \new_[14076]_  = \new_[14075]_  & \new_[14070]_ ;
  assign \new_[14079]_  = A167 & A168;
  assign \new_[14083]_  = ~A232 & A200;
  assign \new_[14084]_  = A199 & \new_[14083]_ ;
  assign \new_[14085]_  = \new_[14084]_  & \new_[14079]_ ;
  assign \new_[14088]_  = ~A265 & ~A233;
  assign \new_[14092]_  = ~A300 & A298;
  assign \new_[14093]_  = ~A266 & \new_[14092]_ ;
  assign \new_[14094]_  = \new_[14093]_  & \new_[14088]_ ;
  assign \new_[14097]_  = A167 & A168;
  assign \new_[14101]_  = ~A232 & A200;
  assign \new_[14102]_  = A199 & \new_[14101]_ ;
  assign \new_[14103]_  = \new_[14102]_  & \new_[14097]_ ;
  assign \new_[14106]_  = ~A265 & ~A233;
  assign \new_[14110]_  = A299 & A298;
  assign \new_[14111]_  = ~A266 & \new_[14110]_ ;
  assign \new_[14112]_  = \new_[14111]_  & \new_[14106]_ ;
  assign \new_[14115]_  = A167 & A168;
  assign \new_[14119]_  = ~A232 & A200;
  assign \new_[14120]_  = A199 & \new_[14119]_ ;
  assign \new_[14121]_  = \new_[14120]_  & \new_[14115]_ ;
  assign \new_[14124]_  = ~A265 & ~A233;
  assign \new_[14128]_  = ~A299 & ~A298;
  assign \new_[14129]_  = ~A266 & \new_[14128]_ ;
  assign \new_[14130]_  = \new_[14129]_  & \new_[14124]_ ;
  assign \new_[14133]_  = A167 & A168;
  assign \new_[14137]_  = A232 & ~A201;
  assign \new_[14138]_  = ~A200 & \new_[14137]_ ;
  assign \new_[14139]_  = \new_[14138]_  & \new_[14133]_ ;
  assign \new_[14142]_  = A265 & A233;
  assign \new_[14146]_  = ~A300 & ~A299;
  assign \new_[14147]_  = ~A267 & \new_[14146]_ ;
  assign \new_[14148]_  = \new_[14147]_  & \new_[14142]_ ;
  assign \new_[14151]_  = A167 & A168;
  assign \new_[14155]_  = A232 & ~A201;
  assign \new_[14156]_  = ~A200 & \new_[14155]_ ;
  assign \new_[14157]_  = \new_[14156]_  & \new_[14151]_ ;
  assign \new_[14160]_  = A265 & A233;
  assign \new_[14164]_  = A299 & A298;
  assign \new_[14165]_  = ~A267 & \new_[14164]_ ;
  assign \new_[14166]_  = \new_[14165]_  & \new_[14160]_ ;
  assign \new_[14169]_  = A167 & A168;
  assign \new_[14173]_  = A232 & ~A201;
  assign \new_[14174]_  = ~A200 & \new_[14173]_ ;
  assign \new_[14175]_  = \new_[14174]_  & \new_[14169]_ ;
  assign \new_[14178]_  = A265 & A233;
  assign \new_[14182]_  = ~A299 & ~A298;
  assign \new_[14183]_  = ~A267 & \new_[14182]_ ;
  assign \new_[14184]_  = \new_[14183]_  & \new_[14178]_ ;
  assign \new_[14187]_  = A167 & A168;
  assign \new_[14191]_  = A232 & ~A201;
  assign \new_[14192]_  = ~A200 & \new_[14191]_ ;
  assign \new_[14193]_  = \new_[14192]_  & \new_[14187]_ ;
  assign \new_[14196]_  = A265 & A233;
  assign \new_[14200]_  = ~A300 & ~A299;
  assign \new_[14201]_  = A266 & \new_[14200]_ ;
  assign \new_[14202]_  = \new_[14201]_  & \new_[14196]_ ;
  assign \new_[14205]_  = A167 & A168;
  assign \new_[14209]_  = A232 & ~A201;
  assign \new_[14210]_  = ~A200 & \new_[14209]_ ;
  assign \new_[14211]_  = \new_[14210]_  & \new_[14205]_ ;
  assign \new_[14214]_  = A265 & A233;
  assign \new_[14218]_  = A299 & A298;
  assign \new_[14219]_  = A266 & \new_[14218]_ ;
  assign \new_[14220]_  = \new_[14219]_  & \new_[14214]_ ;
  assign \new_[14223]_  = A167 & A168;
  assign \new_[14227]_  = A232 & ~A201;
  assign \new_[14228]_  = ~A200 & \new_[14227]_ ;
  assign \new_[14229]_  = \new_[14228]_  & \new_[14223]_ ;
  assign \new_[14232]_  = A265 & A233;
  assign \new_[14236]_  = ~A299 & ~A298;
  assign \new_[14237]_  = A266 & \new_[14236]_ ;
  assign \new_[14238]_  = \new_[14237]_  & \new_[14232]_ ;
  assign \new_[14241]_  = A167 & A168;
  assign \new_[14245]_  = A232 & ~A201;
  assign \new_[14246]_  = ~A200 & \new_[14245]_ ;
  assign \new_[14247]_  = \new_[14246]_  & \new_[14241]_ ;
  assign \new_[14250]_  = ~A265 & A233;
  assign \new_[14254]_  = ~A300 & ~A299;
  assign \new_[14255]_  = ~A266 & \new_[14254]_ ;
  assign \new_[14256]_  = \new_[14255]_  & \new_[14250]_ ;
  assign \new_[14259]_  = A167 & A168;
  assign \new_[14263]_  = A232 & ~A201;
  assign \new_[14264]_  = ~A200 & \new_[14263]_ ;
  assign \new_[14265]_  = \new_[14264]_  & \new_[14259]_ ;
  assign \new_[14268]_  = ~A265 & A233;
  assign \new_[14272]_  = A299 & A298;
  assign \new_[14273]_  = ~A266 & \new_[14272]_ ;
  assign \new_[14274]_  = \new_[14273]_  & \new_[14268]_ ;
  assign \new_[14277]_  = A167 & A168;
  assign \new_[14281]_  = A232 & ~A201;
  assign \new_[14282]_  = ~A200 & \new_[14281]_ ;
  assign \new_[14283]_  = \new_[14282]_  & \new_[14277]_ ;
  assign \new_[14286]_  = ~A265 & A233;
  assign \new_[14290]_  = ~A299 & ~A298;
  assign \new_[14291]_  = ~A266 & \new_[14290]_ ;
  assign \new_[14292]_  = \new_[14291]_  & \new_[14286]_ ;
  assign \new_[14295]_  = A167 & A168;
  assign \new_[14299]_  = ~A232 & ~A201;
  assign \new_[14300]_  = ~A200 & \new_[14299]_ ;
  assign \new_[14301]_  = \new_[14300]_  & \new_[14295]_ ;
  assign \new_[14304]_  = A298 & A233;
  assign \new_[14308]_  = A301 & A300;
  assign \new_[14309]_  = ~A299 & \new_[14308]_ ;
  assign \new_[14310]_  = \new_[14309]_  & \new_[14304]_ ;
  assign \new_[14313]_  = A167 & A168;
  assign \new_[14317]_  = ~A232 & ~A201;
  assign \new_[14318]_  = ~A200 & \new_[14317]_ ;
  assign \new_[14319]_  = \new_[14318]_  & \new_[14313]_ ;
  assign \new_[14322]_  = A298 & A233;
  assign \new_[14326]_  = A302 & A300;
  assign \new_[14327]_  = ~A299 & \new_[14326]_ ;
  assign \new_[14328]_  = \new_[14327]_  & \new_[14322]_ ;
  assign \new_[14331]_  = A167 & A168;
  assign \new_[14335]_  = ~A232 & ~A201;
  assign \new_[14336]_  = ~A200 & \new_[14335]_ ;
  assign \new_[14337]_  = \new_[14336]_  & \new_[14331]_ ;
  assign \new_[14340]_  = A265 & A233;
  assign \new_[14344]_  = A268 & A267;
  assign \new_[14345]_  = ~A266 & \new_[14344]_ ;
  assign \new_[14346]_  = \new_[14345]_  & \new_[14340]_ ;
  assign \new_[14349]_  = A167 & A168;
  assign \new_[14353]_  = ~A232 & ~A201;
  assign \new_[14354]_  = ~A200 & \new_[14353]_ ;
  assign \new_[14355]_  = \new_[14354]_  & \new_[14349]_ ;
  assign \new_[14358]_  = A265 & A233;
  assign \new_[14362]_  = A269 & A267;
  assign \new_[14363]_  = ~A266 & \new_[14362]_ ;
  assign \new_[14364]_  = \new_[14363]_  & \new_[14358]_ ;
  assign \new_[14367]_  = A167 & A168;
  assign \new_[14371]_  = ~A233 & ~A201;
  assign \new_[14372]_  = ~A200 & \new_[14371]_ ;
  assign \new_[14373]_  = \new_[14372]_  & \new_[14367]_ ;
  assign \new_[14376]_  = A265 & ~A234;
  assign \new_[14380]_  = ~A300 & A298;
  assign \new_[14381]_  = A266 & \new_[14380]_ ;
  assign \new_[14382]_  = \new_[14381]_  & \new_[14376]_ ;
  assign \new_[14385]_  = A167 & A168;
  assign \new_[14389]_  = ~A233 & ~A201;
  assign \new_[14390]_  = ~A200 & \new_[14389]_ ;
  assign \new_[14391]_  = \new_[14390]_  & \new_[14385]_ ;
  assign \new_[14394]_  = A265 & ~A234;
  assign \new_[14398]_  = A299 & A298;
  assign \new_[14399]_  = A266 & \new_[14398]_ ;
  assign \new_[14400]_  = \new_[14399]_  & \new_[14394]_ ;
  assign \new_[14403]_  = A167 & A168;
  assign \new_[14407]_  = ~A233 & ~A201;
  assign \new_[14408]_  = ~A200 & \new_[14407]_ ;
  assign \new_[14409]_  = \new_[14408]_  & \new_[14403]_ ;
  assign \new_[14412]_  = A265 & ~A234;
  assign \new_[14416]_  = ~A299 & ~A298;
  assign \new_[14417]_  = A266 & \new_[14416]_ ;
  assign \new_[14418]_  = \new_[14417]_  & \new_[14412]_ ;
  assign \new_[14421]_  = A167 & A168;
  assign \new_[14425]_  = ~A233 & ~A201;
  assign \new_[14426]_  = ~A200 & \new_[14425]_ ;
  assign \new_[14427]_  = \new_[14426]_  & \new_[14421]_ ;
  assign \new_[14430]_  = ~A266 & ~A234;
  assign \new_[14434]_  = ~A300 & A298;
  assign \new_[14435]_  = ~A267 & \new_[14434]_ ;
  assign \new_[14436]_  = \new_[14435]_  & \new_[14430]_ ;
  assign \new_[14439]_  = A167 & A168;
  assign \new_[14443]_  = ~A233 & ~A201;
  assign \new_[14444]_  = ~A200 & \new_[14443]_ ;
  assign \new_[14445]_  = \new_[14444]_  & \new_[14439]_ ;
  assign \new_[14448]_  = ~A266 & ~A234;
  assign \new_[14452]_  = A299 & A298;
  assign \new_[14453]_  = ~A267 & \new_[14452]_ ;
  assign \new_[14454]_  = \new_[14453]_  & \new_[14448]_ ;
  assign \new_[14457]_  = A167 & A168;
  assign \new_[14461]_  = ~A233 & ~A201;
  assign \new_[14462]_  = ~A200 & \new_[14461]_ ;
  assign \new_[14463]_  = \new_[14462]_  & \new_[14457]_ ;
  assign \new_[14466]_  = ~A266 & ~A234;
  assign \new_[14470]_  = ~A299 & ~A298;
  assign \new_[14471]_  = ~A267 & \new_[14470]_ ;
  assign \new_[14472]_  = \new_[14471]_  & \new_[14466]_ ;
  assign \new_[14475]_  = A167 & A168;
  assign \new_[14479]_  = ~A233 & ~A201;
  assign \new_[14480]_  = ~A200 & \new_[14479]_ ;
  assign \new_[14481]_  = \new_[14480]_  & \new_[14475]_ ;
  assign \new_[14484]_  = ~A265 & ~A234;
  assign \new_[14488]_  = ~A300 & A298;
  assign \new_[14489]_  = ~A266 & \new_[14488]_ ;
  assign \new_[14490]_  = \new_[14489]_  & \new_[14484]_ ;
  assign \new_[14493]_  = A167 & A168;
  assign \new_[14497]_  = ~A233 & ~A201;
  assign \new_[14498]_  = ~A200 & \new_[14497]_ ;
  assign \new_[14499]_  = \new_[14498]_  & \new_[14493]_ ;
  assign \new_[14502]_  = ~A265 & ~A234;
  assign \new_[14506]_  = A299 & A298;
  assign \new_[14507]_  = ~A266 & \new_[14506]_ ;
  assign \new_[14508]_  = \new_[14507]_  & \new_[14502]_ ;
  assign \new_[14511]_  = A167 & A168;
  assign \new_[14515]_  = ~A233 & ~A201;
  assign \new_[14516]_  = ~A200 & \new_[14515]_ ;
  assign \new_[14517]_  = \new_[14516]_  & \new_[14511]_ ;
  assign \new_[14520]_  = ~A265 & ~A234;
  assign \new_[14524]_  = ~A299 & ~A298;
  assign \new_[14525]_  = ~A266 & \new_[14524]_ ;
  assign \new_[14526]_  = \new_[14525]_  & \new_[14520]_ ;
  assign \new_[14529]_  = A167 & A168;
  assign \new_[14533]_  = A232 & ~A201;
  assign \new_[14534]_  = ~A200 & \new_[14533]_ ;
  assign \new_[14535]_  = \new_[14534]_  & \new_[14529]_ ;
  assign \new_[14538]_  = A234 & ~A233;
  assign \new_[14542]_  = A299 & ~A298;
  assign \new_[14543]_  = A235 & \new_[14542]_ ;
  assign \new_[14544]_  = \new_[14543]_  & \new_[14538]_ ;
  assign \new_[14547]_  = A167 & A168;
  assign \new_[14551]_  = A232 & ~A201;
  assign \new_[14552]_  = ~A200 & \new_[14551]_ ;
  assign \new_[14553]_  = \new_[14552]_  & \new_[14547]_ ;
  assign \new_[14556]_  = A234 & ~A233;
  assign \new_[14560]_  = A266 & ~A265;
  assign \new_[14561]_  = A235 & \new_[14560]_ ;
  assign \new_[14562]_  = \new_[14561]_  & \new_[14556]_ ;
  assign \new_[14565]_  = A167 & A168;
  assign \new_[14569]_  = A232 & ~A201;
  assign \new_[14570]_  = ~A200 & \new_[14569]_ ;
  assign \new_[14571]_  = \new_[14570]_  & \new_[14565]_ ;
  assign \new_[14574]_  = A234 & ~A233;
  assign \new_[14578]_  = A299 & ~A298;
  assign \new_[14579]_  = A236 & \new_[14578]_ ;
  assign \new_[14580]_  = \new_[14579]_  & \new_[14574]_ ;
  assign \new_[14583]_  = A167 & A168;
  assign \new_[14587]_  = A232 & ~A201;
  assign \new_[14588]_  = ~A200 & \new_[14587]_ ;
  assign \new_[14589]_  = \new_[14588]_  & \new_[14583]_ ;
  assign \new_[14592]_  = A234 & ~A233;
  assign \new_[14596]_  = A266 & ~A265;
  assign \new_[14597]_  = A236 & \new_[14596]_ ;
  assign \new_[14598]_  = \new_[14597]_  & \new_[14592]_ ;
  assign \new_[14601]_  = A167 & A168;
  assign \new_[14605]_  = ~A232 & ~A201;
  assign \new_[14606]_  = ~A200 & \new_[14605]_ ;
  assign \new_[14607]_  = \new_[14606]_  & \new_[14601]_ ;
  assign \new_[14610]_  = A265 & ~A233;
  assign \new_[14614]_  = ~A300 & A298;
  assign \new_[14615]_  = A266 & \new_[14614]_ ;
  assign \new_[14616]_  = \new_[14615]_  & \new_[14610]_ ;
  assign \new_[14619]_  = A167 & A168;
  assign \new_[14623]_  = ~A232 & ~A201;
  assign \new_[14624]_  = ~A200 & \new_[14623]_ ;
  assign \new_[14625]_  = \new_[14624]_  & \new_[14619]_ ;
  assign \new_[14628]_  = A265 & ~A233;
  assign \new_[14632]_  = A299 & A298;
  assign \new_[14633]_  = A266 & \new_[14632]_ ;
  assign \new_[14634]_  = \new_[14633]_  & \new_[14628]_ ;
  assign \new_[14637]_  = A167 & A168;
  assign \new_[14641]_  = ~A232 & ~A201;
  assign \new_[14642]_  = ~A200 & \new_[14641]_ ;
  assign \new_[14643]_  = \new_[14642]_  & \new_[14637]_ ;
  assign \new_[14646]_  = A265 & ~A233;
  assign \new_[14650]_  = ~A299 & ~A298;
  assign \new_[14651]_  = A266 & \new_[14650]_ ;
  assign \new_[14652]_  = \new_[14651]_  & \new_[14646]_ ;
  assign \new_[14655]_  = A167 & A168;
  assign \new_[14659]_  = ~A232 & ~A201;
  assign \new_[14660]_  = ~A200 & \new_[14659]_ ;
  assign \new_[14661]_  = \new_[14660]_  & \new_[14655]_ ;
  assign \new_[14664]_  = ~A266 & ~A233;
  assign \new_[14668]_  = ~A300 & A298;
  assign \new_[14669]_  = ~A267 & \new_[14668]_ ;
  assign \new_[14670]_  = \new_[14669]_  & \new_[14664]_ ;
  assign \new_[14673]_  = A167 & A168;
  assign \new_[14677]_  = ~A232 & ~A201;
  assign \new_[14678]_  = ~A200 & \new_[14677]_ ;
  assign \new_[14679]_  = \new_[14678]_  & \new_[14673]_ ;
  assign \new_[14682]_  = ~A266 & ~A233;
  assign \new_[14686]_  = A299 & A298;
  assign \new_[14687]_  = ~A267 & \new_[14686]_ ;
  assign \new_[14688]_  = \new_[14687]_  & \new_[14682]_ ;
  assign \new_[14691]_  = A167 & A168;
  assign \new_[14695]_  = ~A232 & ~A201;
  assign \new_[14696]_  = ~A200 & \new_[14695]_ ;
  assign \new_[14697]_  = \new_[14696]_  & \new_[14691]_ ;
  assign \new_[14700]_  = ~A266 & ~A233;
  assign \new_[14704]_  = ~A299 & ~A298;
  assign \new_[14705]_  = ~A267 & \new_[14704]_ ;
  assign \new_[14706]_  = \new_[14705]_  & \new_[14700]_ ;
  assign \new_[14709]_  = A167 & A168;
  assign \new_[14713]_  = ~A232 & ~A201;
  assign \new_[14714]_  = ~A200 & \new_[14713]_ ;
  assign \new_[14715]_  = \new_[14714]_  & \new_[14709]_ ;
  assign \new_[14718]_  = ~A265 & ~A233;
  assign \new_[14722]_  = ~A300 & A298;
  assign \new_[14723]_  = ~A266 & \new_[14722]_ ;
  assign \new_[14724]_  = \new_[14723]_  & \new_[14718]_ ;
  assign \new_[14727]_  = A167 & A168;
  assign \new_[14731]_  = ~A232 & ~A201;
  assign \new_[14732]_  = ~A200 & \new_[14731]_ ;
  assign \new_[14733]_  = \new_[14732]_  & \new_[14727]_ ;
  assign \new_[14736]_  = ~A265 & ~A233;
  assign \new_[14740]_  = A299 & A298;
  assign \new_[14741]_  = ~A266 & \new_[14740]_ ;
  assign \new_[14742]_  = \new_[14741]_  & \new_[14736]_ ;
  assign \new_[14745]_  = A167 & A168;
  assign \new_[14749]_  = ~A232 & ~A201;
  assign \new_[14750]_  = ~A200 & \new_[14749]_ ;
  assign \new_[14751]_  = \new_[14750]_  & \new_[14745]_ ;
  assign \new_[14754]_  = ~A265 & ~A233;
  assign \new_[14758]_  = ~A299 & ~A298;
  assign \new_[14759]_  = ~A266 & \new_[14758]_ ;
  assign \new_[14760]_  = \new_[14759]_  & \new_[14754]_ ;
  assign \new_[14763]_  = A167 & A168;
  assign \new_[14767]_  = A232 & ~A200;
  assign \new_[14768]_  = ~A199 & \new_[14767]_ ;
  assign \new_[14769]_  = \new_[14768]_  & \new_[14763]_ ;
  assign \new_[14772]_  = A265 & A233;
  assign \new_[14776]_  = ~A300 & ~A299;
  assign \new_[14777]_  = ~A267 & \new_[14776]_ ;
  assign \new_[14778]_  = \new_[14777]_  & \new_[14772]_ ;
  assign \new_[14781]_  = A167 & A168;
  assign \new_[14785]_  = A232 & ~A200;
  assign \new_[14786]_  = ~A199 & \new_[14785]_ ;
  assign \new_[14787]_  = \new_[14786]_  & \new_[14781]_ ;
  assign \new_[14790]_  = A265 & A233;
  assign \new_[14794]_  = A299 & A298;
  assign \new_[14795]_  = ~A267 & \new_[14794]_ ;
  assign \new_[14796]_  = \new_[14795]_  & \new_[14790]_ ;
  assign \new_[14799]_  = A167 & A168;
  assign \new_[14803]_  = A232 & ~A200;
  assign \new_[14804]_  = ~A199 & \new_[14803]_ ;
  assign \new_[14805]_  = \new_[14804]_  & \new_[14799]_ ;
  assign \new_[14808]_  = A265 & A233;
  assign \new_[14812]_  = ~A299 & ~A298;
  assign \new_[14813]_  = ~A267 & \new_[14812]_ ;
  assign \new_[14814]_  = \new_[14813]_  & \new_[14808]_ ;
  assign \new_[14817]_  = A167 & A168;
  assign \new_[14821]_  = A232 & ~A200;
  assign \new_[14822]_  = ~A199 & \new_[14821]_ ;
  assign \new_[14823]_  = \new_[14822]_  & \new_[14817]_ ;
  assign \new_[14826]_  = A265 & A233;
  assign \new_[14830]_  = ~A300 & ~A299;
  assign \new_[14831]_  = A266 & \new_[14830]_ ;
  assign \new_[14832]_  = \new_[14831]_  & \new_[14826]_ ;
  assign \new_[14835]_  = A167 & A168;
  assign \new_[14839]_  = A232 & ~A200;
  assign \new_[14840]_  = ~A199 & \new_[14839]_ ;
  assign \new_[14841]_  = \new_[14840]_  & \new_[14835]_ ;
  assign \new_[14844]_  = A265 & A233;
  assign \new_[14848]_  = A299 & A298;
  assign \new_[14849]_  = A266 & \new_[14848]_ ;
  assign \new_[14850]_  = \new_[14849]_  & \new_[14844]_ ;
  assign \new_[14853]_  = A167 & A168;
  assign \new_[14857]_  = A232 & ~A200;
  assign \new_[14858]_  = ~A199 & \new_[14857]_ ;
  assign \new_[14859]_  = \new_[14858]_  & \new_[14853]_ ;
  assign \new_[14862]_  = A265 & A233;
  assign \new_[14866]_  = ~A299 & ~A298;
  assign \new_[14867]_  = A266 & \new_[14866]_ ;
  assign \new_[14868]_  = \new_[14867]_  & \new_[14862]_ ;
  assign \new_[14871]_  = A167 & A168;
  assign \new_[14875]_  = A232 & ~A200;
  assign \new_[14876]_  = ~A199 & \new_[14875]_ ;
  assign \new_[14877]_  = \new_[14876]_  & \new_[14871]_ ;
  assign \new_[14880]_  = ~A265 & A233;
  assign \new_[14884]_  = ~A300 & ~A299;
  assign \new_[14885]_  = ~A266 & \new_[14884]_ ;
  assign \new_[14886]_  = \new_[14885]_  & \new_[14880]_ ;
  assign \new_[14889]_  = A167 & A168;
  assign \new_[14893]_  = A232 & ~A200;
  assign \new_[14894]_  = ~A199 & \new_[14893]_ ;
  assign \new_[14895]_  = \new_[14894]_  & \new_[14889]_ ;
  assign \new_[14898]_  = ~A265 & A233;
  assign \new_[14902]_  = A299 & A298;
  assign \new_[14903]_  = ~A266 & \new_[14902]_ ;
  assign \new_[14904]_  = \new_[14903]_  & \new_[14898]_ ;
  assign \new_[14907]_  = A167 & A168;
  assign \new_[14911]_  = A232 & ~A200;
  assign \new_[14912]_  = ~A199 & \new_[14911]_ ;
  assign \new_[14913]_  = \new_[14912]_  & \new_[14907]_ ;
  assign \new_[14916]_  = ~A265 & A233;
  assign \new_[14920]_  = ~A299 & ~A298;
  assign \new_[14921]_  = ~A266 & \new_[14920]_ ;
  assign \new_[14922]_  = \new_[14921]_  & \new_[14916]_ ;
  assign \new_[14925]_  = A167 & A168;
  assign \new_[14929]_  = ~A232 & ~A200;
  assign \new_[14930]_  = ~A199 & \new_[14929]_ ;
  assign \new_[14931]_  = \new_[14930]_  & \new_[14925]_ ;
  assign \new_[14934]_  = A298 & A233;
  assign \new_[14938]_  = A301 & A300;
  assign \new_[14939]_  = ~A299 & \new_[14938]_ ;
  assign \new_[14940]_  = \new_[14939]_  & \new_[14934]_ ;
  assign \new_[14943]_  = A167 & A168;
  assign \new_[14947]_  = ~A232 & ~A200;
  assign \new_[14948]_  = ~A199 & \new_[14947]_ ;
  assign \new_[14949]_  = \new_[14948]_  & \new_[14943]_ ;
  assign \new_[14952]_  = A298 & A233;
  assign \new_[14956]_  = A302 & A300;
  assign \new_[14957]_  = ~A299 & \new_[14956]_ ;
  assign \new_[14958]_  = \new_[14957]_  & \new_[14952]_ ;
  assign \new_[14961]_  = A167 & A168;
  assign \new_[14965]_  = ~A232 & ~A200;
  assign \new_[14966]_  = ~A199 & \new_[14965]_ ;
  assign \new_[14967]_  = \new_[14966]_  & \new_[14961]_ ;
  assign \new_[14970]_  = A265 & A233;
  assign \new_[14974]_  = A268 & A267;
  assign \new_[14975]_  = ~A266 & \new_[14974]_ ;
  assign \new_[14976]_  = \new_[14975]_  & \new_[14970]_ ;
  assign \new_[14979]_  = A167 & A168;
  assign \new_[14983]_  = ~A232 & ~A200;
  assign \new_[14984]_  = ~A199 & \new_[14983]_ ;
  assign \new_[14985]_  = \new_[14984]_  & \new_[14979]_ ;
  assign \new_[14988]_  = A265 & A233;
  assign \new_[14992]_  = A269 & A267;
  assign \new_[14993]_  = ~A266 & \new_[14992]_ ;
  assign \new_[14994]_  = \new_[14993]_  & \new_[14988]_ ;
  assign \new_[14997]_  = A167 & A168;
  assign \new_[15001]_  = ~A233 & ~A200;
  assign \new_[15002]_  = ~A199 & \new_[15001]_ ;
  assign \new_[15003]_  = \new_[15002]_  & \new_[14997]_ ;
  assign \new_[15006]_  = A265 & ~A234;
  assign \new_[15010]_  = ~A300 & A298;
  assign \new_[15011]_  = A266 & \new_[15010]_ ;
  assign \new_[15012]_  = \new_[15011]_  & \new_[15006]_ ;
  assign \new_[15015]_  = A167 & A168;
  assign \new_[15019]_  = ~A233 & ~A200;
  assign \new_[15020]_  = ~A199 & \new_[15019]_ ;
  assign \new_[15021]_  = \new_[15020]_  & \new_[15015]_ ;
  assign \new_[15024]_  = A265 & ~A234;
  assign \new_[15028]_  = A299 & A298;
  assign \new_[15029]_  = A266 & \new_[15028]_ ;
  assign \new_[15030]_  = \new_[15029]_  & \new_[15024]_ ;
  assign \new_[15033]_  = A167 & A168;
  assign \new_[15037]_  = ~A233 & ~A200;
  assign \new_[15038]_  = ~A199 & \new_[15037]_ ;
  assign \new_[15039]_  = \new_[15038]_  & \new_[15033]_ ;
  assign \new_[15042]_  = A265 & ~A234;
  assign \new_[15046]_  = ~A299 & ~A298;
  assign \new_[15047]_  = A266 & \new_[15046]_ ;
  assign \new_[15048]_  = \new_[15047]_  & \new_[15042]_ ;
  assign \new_[15051]_  = A167 & A168;
  assign \new_[15055]_  = ~A233 & ~A200;
  assign \new_[15056]_  = ~A199 & \new_[15055]_ ;
  assign \new_[15057]_  = \new_[15056]_  & \new_[15051]_ ;
  assign \new_[15060]_  = ~A266 & ~A234;
  assign \new_[15064]_  = ~A300 & A298;
  assign \new_[15065]_  = ~A267 & \new_[15064]_ ;
  assign \new_[15066]_  = \new_[15065]_  & \new_[15060]_ ;
  assign \new_[15069]_  = A167 & A168;
  assign \new_[15073]_  = ~A233 & ~A200;
  assign \new_[15074]_  = ~A199 & \new_[15073]_ ;
  assign \new_[15075]_  = \new_[15074]_  & \new_[15069]_ ;
  assign \new_[15078]_  = ~A266 & ~A234;
  assign \new_[15082]_  = A299 & A298;
  assign \new_[15083]_  = ~A267 & \new_[15082]_ ;
  assign \new_[15084]_  = \new_[15083]_  & \new_[15078]_ ;
  assign \new_[15087]_  = A167 & A168;
  assign \new_[15091]_  = ~A233 & ~A200;
  assign \new_[15092]_  = ~A199 & \new_[15091]_ ;
  assign \new_[15093]_  = \new_[15092]_  & \new_[15087]_ ;
  assign \new_[15096]_  = ~A266 & ~A234;
  assign \new_[15100]_  = ~A299 & ~A298;
  assign \new_[15101]_  = ~A267 & \new_[15100]_ ;
  assign \new_[15102]_  = \new_[15101]_  & \new_[15096]_ ;
  assign \new_[15105]_  = A167 & A168;
  assign \new_[15109]_  = ~A233 & ~A200;
  assign \new_[15110]_  = ~A199 & \new_[15109]_ ;
  assign \new_[15111]_  = \new_[15110]_  & \new_[15105]_ ;
  assign \new_[15114]_  = ~A265 & ~A234;
  assign \new_[15118]_  = ~A300 & A298;
  assign \new_[15119]_  = ~A266 & \new_[15118]_ ;
  assign \new_[15120]_  = \new_[15119]_  & \new_[15114]_ ;
  assign \new_[15123]_  = A167 & A168;
  assign \new_[15127]_  = ~A233 & ~A200;
  assign \new_[15128]_  = ~A199 & \new_[15127]_ ;
  assign \new_[15129]_  = \new_[15128]_  & \new_[15123]_ ;
  assign \new_[15132]_  = ~A265 & ~A234;
  assign \new_[15136]_  = A299 & A298;
  assign \new_[15137]_  = ~A266 & \new_[15136]_ ;
  assign \new_[15138]_  = \new_[15137]_  & \new_[15132]_ ;
  assign \new_[15141]_  = A167 & A168;
  assign \new_[15145]_  = ~A233 & ~A200;
  assign \new_[15146]_  = ~A199 & \new_[15145]_ ;
  assign \new_[15147]_  = \new_[15146]_  & \new_[15141]_ ;
  assign \new_[15150]_  = ~A265 & ~A234;
  assign \new_[15154]_  = ~A299 & ~A298;
  assign \new_[15155]_  = ~A266 & \new_[15154]_ ;
  assign \new_[15156]_  = \new_[15155]_  & \new_[15150]_ ;
  assign \new_[15159]_  = A167 & A168;
  assign \new_[15163]_  = A232 & ~A200;
  assign \new_[15164]_  = ~A199 & \new_[15163]_ ;
  assign \new_[15165]_  = \new_[15164]_  & \new_[15159]_ ;
  assign \new_[15168]_  = A234 & ~A233;
  assign \new_[15172]_  = A299 & ~A298;
  assign \new_[15173]_  = A235 & \new_[15172]_ ;
  assign \new_[15174]_  = \new_[15173]_  & \new_[15168]_ ;
  assign \new_[15177]_  = A167 & A168;
  assign \new_[15181]_  = A232 & ~A200;
  assign \new_[15182]_  = ~A199 & \new_[15181]_ ;
  assign \new_[15183]_  = \new_[15182]_  & \new_[15177]_ ;
  assign \new_[15186]_  = A234 & ~A233;
  assign \new_[15190]_  = A266 & ~A265;
  assign \new_[15191]_  = A235 & \new_[15190]_ ;
  assign \new_[15192]_  = \new_[15191]_  & \new_[15186]_ ;
  assign \new_[15195]_  = A167 & A168;
  assign \new_[15199]_  = A232 & ~A200;
  assign \new_[15200]_  = ~A199 & \new_[15199]_ ;
  assign \new_[15201]_  = \new_[15200]_  & \new_[15195]_ ;
  assign \new_[15204]_  = A234 & ~A233;
  assign \new_[15208]_  = A299 & ~A298;
  assign \new_[15209]_  = A236 & \new_[15208]_ ;
  assign \new_[15210]_  = \new_[15209]_  & \new_[15204]_ ;
  assign \new_[15213]_  = A167 & A168;
  assign \new_[15217]_  = A232 & ~A200;
  assign \new_[15218]_  = ~A199 & \new_[15217]_ ;
  assign \new_[15219]_  = \new_[15218]_  & \new_[15213]_ ;
  assign \new_[15222]_  = A234 & ~A233;
  assign \new_[15226]_  = A266 & ~A265;
  assign \new_[15227]_  = A236 & \new_[15226]_ ;
  assign \new_[15228]_  = \new_[15227]_  & \new_[15222]_ ;
  assign \new_[15231]_  = A167 & A168;
  assign \new_[15235]_  = ~A232 & ~A200;
  assign \new_[15236]_  = ~A199 & \new_[15235]_ ;
  assign \new_[15237]_  = \new_[15236]_  & \new_[15231]_ ;
  assign \new_[15240]_  = A265 & ~A233;
  assign \new_[15244]_  = ~A300 & A298;
  assign \new_[15245]_  = A266 & \new_[15244]_ ;
  assign \new_[15246]_  = \new_[15245]_  & \new_[15240]_ ;
  assign \new_[15249]_  = A167 & A168;
  assign \new_[15253]_  = ~A232 & ~A200;
  assign \new_[15254]_  = ~A199 & \new_[15253]_ ;
  assign \new_[15255]_  = \new_[15254]_  & \new_[15249]_ ;
  assign \new_[15258]_  = A265 & ~A233;
  assign \new_[15262]_  = A299 & A298;
  assign \new_[15263]_  = A266 & \new_[15262]_ ;
  assign \new_[15264]_  = \new_[15263]_  & \new_[15258]_ ;
  assign \new_[15267]_  = A167 & A168;
  assign \new_[15271]_  = ~A232 & ~A200;
  assign \new_[15272]_  = ~A199 & \new_[15271]_ ;
  assign \new_[15273]_  = \new_[15272]_  & \new_[15267]_ ;
  assign \new_[15276]_  = A265 & ~A233;
  assign \new_[15280]_  = ~A299 & ~A298;
  assign \new_[15281]_  = A266 & \new_[15280]_ ;
  assign \new_[15282]_  = \new_[15281]_  & \new_[15276]_ ;
  assign \new_[15285]_  = A167 & A168;
  assign \new_[15289]_  = ~A232 & ~A200;
  assign \new_[15290]_  = ~A199 & \new_[15289]_ ;
  assign \new_[15291]_  = \new_[15290]_  & \new_[15285]_ ;
  assign \new_[15294]_  = ~A266 & ~A233;
  assign \new_[15298]_  = ~A300 & A298;
  assign \new_[15299]_  = ~A267 & \new_[15298]_ ;
  assign \new_[15300]_  = \new_[15299]_  & \new_[15294]_ ;
  assign \new_[15303]_  = A167 & A168;
  assign \new_[15307]_  = ~A232 & ~A200;
  assign \new_[15308]_  = ~A199 & \new_[15307]_ ;
  assign \new_[15309]_  = \new_[15308]_  & \new_[15303]_ ;
  assign \new_[15312]_  = ~A266 & ~A233;
  assign \new_[15316]_  = A299 & A298;
  assign \new_[15317]_  = ~A267 & \new_[15316]_ ;
  assign \new_[15318]_  = \new_[15317]_  & \new_[15312]_ ;
  assign \new_[15321]_  = A167 & A168;
  assign \new_[15325]_  = ~A232 & ~A200;
  assign \new_[15326]_  = ~A199 & \new_[15325]_ ;
  assign \new_[15327]_  = \new_[15326]_  & \new_[15321]_ ;
  assign \new_[15330]_  = ~A266 & ~A233;
  assign \new_[15334]_  = ~A299 & ~A298;
  assign \new_[15335]_  = ~A267 & \new_[15334]_ ;
  assign \new_[15336]_  = \new_[15335]_  & \new_[15330]_ ;
  assign \new_[15339]_  = A167 & A168;
  assign \new_[15343]_  = ~A232 & ~A200;
  assign \new_[15344]_  = ~A199 & \new_[15343]_ ;
  assign \new_[15345]_  = \new_[15344]_  & \new_[15339]_ ;
  assign \new_[15348]_  = ~A265 & ~A233;
  assign \new_[15352]_  = ~A300 & A298;
  assign \new_[15353]_  = ~A266 & \new_[15352]_ ;
  assign \new_[15354]_  = \new_[15353]_  & \new_[15348]_ ;
  assign \new_[15357]_  = A167 & A168;
  assign \new_[15361]_  = ~A232 & ~A200;
  assign \new_[15362]_  = ~A199 & \new_[15361]_ ;
  assign \new_[15363]_  = \new_[15362]_  & \new_[15357]_ ;
  assign \new_[15366]_  = ~A265 & ~A233;
  assign \new_[15370]_  = A299 & A298;
  assign \new_[15371]_  = ~A266 & \new_[15370]_ ;
  assign \new_[15372]_  = \new_[15371]_  & \new_[15366]_ ;
  assign \new_[15375]_  = A167 & A168;
  assign \new_[15379]_  = ~A232 & ~A200;
  assign \new_[15380]_  = ~A199 & \new_[15379]_ ;
  assign \new_[15381]_  = \new_[15380]_  & \new_[15375]_ ;
  assign \new_[15384]_  = ~A265 & ~A233;
  assign \new_[15388]_  = ~A299 & ~A298;
  assign \new_[15389]_  = ~A266 & \new_[15388]_ ;
  assign \new_[15390]_  = \new_[15389]_  & \new_[15384]_ ;
  assign \new_[15393]_  = ~A168 & A170;
  assign \new_[15397]_  = ~A199 & A166;
  assign \new_[15398]_  = A167 & \new_[15397]_ ;
  assign \new_[15399]_  = \new_[15398]_  & \new_[15393]_ ;
  assign \new_[15402]_  = ~A232 & A200;
  assign \new_[15406]_  = A299 & ~A298;
  assign \new_[15407]_  = A233 & \new_[15406]_ ;
  assign \new_[15408]_  = \new_[15407]_  & \new_[15402]_ ;
  assign \new_[15411]_  = ~A168 & A170;
  assign \new_[15415]_  = ~A199 & A166;
  assign \new_[15416]_  = A167 & \new_[15415]_ ;
  assign \new_[15417]_  = \new_[15416]_  & \new_[15411]_ ;
  assign \new_[15420]_  = ~A232 & A200;
  assign \new_[15424]_  = A266 & ~A265;
  assign \new_[15425]_  = A233 & \new_[15424]_ ;
  assign \new_[15426]_  = \new_[15425]_  & \new_[15420]_ ;
  assign \new_[15429]_  = ~A168 & ~A170;
  assign \new_[15433]_  = ~A199 & ~A166;
  assign \new_[15434]_  = A167 & \new_[15433]_ ;
  assign \new_[15435]_  = \new_[15434]_  & \new_[15429]_ ;
  assign \new_[15438]_  = ~A232 & A200;
  assign \new_[15442]_  = A299 & ~A298;
  assign \new_[15443]_  = A233 & \new_[15442]_ ;
  assign \new_[15444]_  = \new_[15443]_  & \new_[15438]_ ;
  assign \new_[15447]_  = ~A168 & ~A170;
  assign \new_[15451]_  = ~A199 & ~A166;
  assign \new_[15452]_  = A167 & \new_[15451]_ ;
  assign \new_[15453]_  = \new_[15452]_  & \new_[15447]_ ;
  assign \new_[15456]_  = ~A232 & A200;
  assign \new_[15460]_  = A266 & ~A265;
  assign \new_[15461]_  = A233 & \new_[15460]_ ;
  assign \new_[15462]_  = \new_[15461]_  & \new_[15456]_ ;
  assign \new_[15465]_  = ~A168 & ~A170;
  assign \new_[15469]_  = ~A199 & A166;
  assign \new_[15470]_  = ~A167 & \new_[15469]_ ;
  assign \new_[15471]_  = \new_[15470]_  & \new_[15465]_ ;
  assign \new_[15474]_  = ~A232 & A200;
  assign \new_[15478]_  = A299 & ~A298;
  assign \new_[15479]_  = A233 & \new_[15478]_ ;
  assign \new_[15480]_  = \new_[15479]_  & \new_[15474]_ ;
  assign \new_[15483]_  = ~A168 & ~A170;
  assign \new_[15487]_  = ~A199 & A166;
  assign \new_[15488]_  = ~A167 & \new_[15487]_ ;
  assign \new_[15489]_  = \new_[15488]_  & \new_[15483]_ ;
  assign \new_[15492]_  = ~A232 & A200;
  assign \new_[15496]_  = A266 & ~A265;
  assign \new_[15497]_  = A233 & \new_[15496]_ ;
  assign \new_[15498]_  = \new_[15497]_  & \new_[15492]_ ;
  assign \new_[15501]_  = ~A168 & A169;
  assign \new_[15505]_  = ~A199 & ~A166;
  assign \new_[15506]_  = A167 & \new_[15505]_ ;
  assign \new_[15507]_  = \new_[15506]_  & \new_[15501]_ ;
  assign \new_[15510]_  = ~A232 & A200;
  assign \new_[15514]_  = A299 & ~A298;
  assign \new_[15515]_  = A233 & \new_[15514]_ ;
  assign \new_[15516]_  = \new_[15515]_  & \new_[15510]_ ;
  assign \new_[15519]_  = ~A168 & A169;
  assign \new_[15523]_  = ~A199 & ~A166;
  assign \new_[15524]_  = A167 & \new_[15523]_ ;
  assign \new_[15525]_  = \new_[15524]_  & \new_[15519]_ ;
  assign \new_[15528]_  = ~A232 & A200;
  assign \new_[15532]_  = A266 & ~A265;
  assign \new_[15533]_  = A233 & \new_[15532]_ ;
  assign \new_[15534]_  = \new_[15533]_  & \new_[15528]_ ;
  assign \new_[15537]_  = ~A168 & A169;
  assign \new_[15541]_  = ~A199 & A166;
  assign \new_[15542]_  = ~A167 & \new_[15541]_ ;
  assign \new_[15543]_  = \new_[15542]_  & \new_[15537]_ ;
  assign \new_[15546]_  = ~A232 & A200;
  assign \new_[15550]_  = A299 & ~A298;
  assign \new_[15551]_  = A233 & \new_[15550]_ ;
  assign \new_[15552]_  = \new_[15551]_  & \new_[15546]_ ;
  assign \new_[15555]_  = ~A168 & A169;
  assign \new_[15559]_  = ~A199 & A166;
  assign \new_[15560]_  = ~A167 & \new_[15559]_ ;
  assign \new_[15561]_  = \new_[15560]_  & \new_[15555]_ ;
  assign \new_[15564]_  = ~A232 & A200;
  assign \new_[15568]_  = A266 & ~A265;
  assign \new_[15569]_  = A233 & \new_[15568]_ ;
  assign \new_[15570]_  = \new_[15569]_  & \new_[15564]_ ;
  assign \new_[15573]_  = A169 & ~A170;
  assign \new_[15577]_  = A199 & A166;
  assign \new_[15578]_  = A167 & \new_[15577]_ ;
  assign \new_[15579]_  = \new_[15578]_  & \new_[15573]_ ;
  assign \new_[15582]_  = ~A232 & A200;
  assign \new_[15586]_  = A299 & ~A298;
  assign \new_[15587]_  = A233 & \new_[15586]_ ;
  assign \new_[15588]_  = \new_[15587]_  & \new_[15582]_ ;
  assign \new_[15591]_  = A169 & ~A170;
  assign \new_[15595]_  = A199 & A166;
  assign \new_[15596]_  = A167 & \new_[15595]_ ;
  assign \new_[15597]_  = \new_[15596]_  & \new_[15591]_ ;
  assign \new_[15600]_  = ~A232 & A200;
  assign \new_[15604]_  = A266 & ~A265;
  assign \new_[15605]_  = A233 & \new_[15604]_ ;
  assign \new_[15606]_  = \new_[15605]_  & \new_[15600]_ ;
  assign \new_[15609]_  = A169 & ~A170;
  assign \new_[15613]_  = ~A200 & A166;
  assign \new_[15614]_  = A167 & \new_[15613]_ ;
  assign \new_[15615]_  = \new_[15614]_  & \new_[15609]_ ;
  assign \new_[15618]_  = ~A232 & ~A201;
  assign \new_[15622]_  = A299 & ~A298;
  assign \new_[15623]_  = A233 & \new_[15622]_ ;
  assign \new_[15624]_  = \new_[15623]_  & \new_[15618]_ ;
  assign \new_[15627]_  = A169 & ~A170;
  assign \new_[15631]_  = ~A200 & A166;
  assign \new_[15632]_  = A167 & \new_[15631]_ ;
  assign \new_[15633]_  = \new_[15632]_  & \new_[15627]_ ;
  assign \new_[15636]_  = ~A232 & ~A201;
  assign \new_[15640]_  = A266 & ~A265;
  assign \new_[15641]_  = A233 & \new_[15640]_ ;
  assign \new_[15642]_  = \new_[15641]_  & \new_[15636]_ ;
  assign \new_[15645]_  = A169 & ~A170;
  assign \new_[15649]_  = ~A199 & A166;
  assign \new_[15650]_  = A167 & \new_[15649]_ ;
  assign \new_[15651]_  = \new_[15650]_  & \new_[15645]_ ;
  assign \new_[15654]_  = ~A232 & ~A200;
  assign \new_[15658]_  = A299 & ~A298;
  assign \new_[15659]_  = A233 & \new_[15658]_ ;
  assign \new_[15660]_  = \new_[15659]_  & \new_[15654]_ ;
  assign \new_[15663]_  = A169 & ~A170;
  assign \new_[15667]_  = ~A199 & A166;
  assign \new_[15668]_  = A167 & \new_[15667]_ ;
  assign \new_[15669]_  = \new_[15668]_  & \new_[15663]_ ;
  assign \new_[15672]_  = ~A232 & ~A200;
  assign \new_[15676]_  = A266 & ~A265;
  assign \new_[15677]_  = A233 & \new_[15676]_ ;
  assign \new_[15678]_  = \new_[15677]_  & \new_[15672]_ ;
  assign \new_[15681]_  = A169 & ~A170;
  assign \new_[15685]_  = A199 & ~A166;
  assign \new_[15686]_  = ~A167 & \new_[15685]_ ;
  assign \new_[15687]_  = \new_[15686]_  & \new_[15681]_ ;
  assign \new_[15690]_  = ~A232 & A200;
  assign \new_[15694]_  = A299 & ~A298;
  assign \new_[15695]_  = A233 & \new_[15694]_ ;
  assign \new_[15696]_  = \new_[15695]_  & \new_[15690]_ ;
  assign \new_[15699]_  = A169 & ~A170;
  assign \new_[15703]_  = A199 & ~A166;
  assign \new_[15704]_  = ~A167 & \new_[15703]_ ;
  assign \new_[15705]_  = \new_[15704]_  & \new_[15699]_ ;
  assign \new_[15708]_  = ~A232 & A200;
  assign \new_[15712]_  = A266 & ~A265;
  assign \new_[15713]_  = A233 & \new_[15712]_ ;
  assign \new_[15714]_  = \new_[15713]_  & \new_[15708]_ ;
  assign \new_[15717]_  = A169 & ~A170;
  assign \new_[15721]_  = ~A200 & ~A166;
  assign \new_[15722]_  = ~A167 & \new_[15721]_ ;
  assign \new_[15723]_  = \new_[15722]_  & \new_[15717]_ ;
  assign \new_[15726]_  = ~A232 & ~A201;
  assign \new_[15730]_  = A299 & ~A298;
  assign \new_[15731]_  = A233 & \new_[15730]_ ;
  assign \new_[15732]_  = \new_[15731]_  & \new_[15726]_ ;
  assign \new_[15735]_  = A169 & ~A170;
  assign \new_[15739]_  = ~A200 & ~A166;
  assign \new_[15740]_  = ~A167 & \new_[15739]_ ;
  assign \new_[15741]_  = \new_[15740]_  & \new_[15735]_ ;
  assign \new_[15744]_  = ~A232 & ~A201;
  assign \new_[15748]_  = A266 & ~A265;
  assign \new_[15749]_  = A233 & \new_[15748]_ ;
  assign \new_[15750]_  = \new_[15749]_  & \new_[15744]_ ;
  assign \new_[15753]_  = A169 & ~A170;
  assign \new_[15757]_  = ~A199 & ~A166;
  assign \new_[15758]_  = ~A167 & \new_[15757]_ ;
  assign \new_[15759]_  = \new_[15758]_  & \new_[15753]_ ;
  assign \new_[15762]_  = ~A232 & ~A200;
  assign \new_[15766]_  = A299 & ~A298;
  assign \new_[15767]_  = A233 & \new_[15766]_ ;
  assign \new_[15768]_  = \new_[15767]_  & \new_[15762]_ ;
  assign \new_[15771]_  = A169 & ~A170;
  assign \new_[15775]_  = ~A199 & ~A166;
  assign \new_[15776]_  = ~A167 & \new_[15775]_ ;
  assign \new_[15777]_  = \new_[15776]_  & \new_[15771]_ ;
  assign \new_[15780]_  = ~A232 & ~A200;
  assign \new_[15784]_  = A266 & ~A265;
  assign \new_[15785]_  = A233 & \new_[15784]_ ;
  assign \new_[15786]_  = \new_[15785]_  & \new_[15780]_ ;
  assign \new_[15789]_  = ~A168 & ~A169;
  assign \new_[15793]_  = ~A199 & A166;
  assign \new_[15794]_  = A167 & \new_[15793]_ ;
  assign \new_[15795]_  = \new_[15794]_  & \new_[15789]_ ;
  assign \new_[15798]_  = ~A232 & A200;
  assign \new_[15802]_  = A299 & ~A298;
  assign \new_[15803]_  = A233 & \new_[15802]_ ;
  assign \new_[15804]_  = \new_[15803]_  & \new_[15798]_ ;
  assign \new_[15807]_  = ~A168 & ~A169;
  assign \new_[15811]_  = ~A199 & A166;
  assign \new_[15812]_  = A167 & \new_[15811]_ ;
  assign \new_[15813]_  = \new_[15812]_  & \new_[15807]_ ;
  assign \new_[15816]_  = ~A232 & A200;
  assign \new_[15820]_  = A266 & ~A265;
  assign \new_[15821]_  = A233 & \new_[15820]_ ;
  assign \new_[15822]_  = \new_[15821]_  & \new_[15816]_ ;
  assign \new_[15825]_  = ~A169 & A170;
  assign \new_[15829]_  = A199 & ~A166;
  assign \new_[15830]_  = A167 & \new_[15829]_ ;
  assign \new_[15831]_  = \new_[15830]_  & \new_[15825]_ ;
  assign \new_[15834]_  = ~A232 & A200;
  assign \new_[15838]_  = A299 & ~A298;
  assign \new_[15839]_  = A233 & \new_[15838]_ ;
  assign \new_[15840]_  = \new_[15839]_  & \new_[15834]_ ;
  assign \new_[15843]_  = ~A169 & A170;
  assign \new_[15847]_  = A199 & ~A166;
  assign \new_[15848]_  = A167 & \new_[15847]_ ;
  assign \new_[15849]_  = \new_[15848]_  & \new_[15843]_ ;
  assign \new_[15852]_  = ~A232 & A200;
  assign \new_[15856]_  = A266 & ~A265;
  assign \new_[15857]_  = A233 & \new_[15856]_ ;
  assign \new_[15858]_  = \new_[15857]_  & \new_[15852]_ ;
  assign \new_[15861]_  = ~A169 & A170;
  assign \new_[15865]_  = ~A200 & ~A166;
  assign \new_[15866]_  = A167 & \new_[15865]_ ;
  assign \new_[15867]_  = \new_[15866]_  & \new_[15861]_ ;
  assign \new_[15870]_  = ~A232 & ~A201;
  assign \new_[15874]_  = A299 & ~A298;
  assign \new_[15875]_  = A233 & \new_[15874]_ ;
  assign \new_[15876]_  = \new_[15875]_  & \new_[15870]_ ;
  assign \new_[15879]_  = ~A169 & A170;
  assign \new_[15883]_  = ~A200 & ~A166;
  assign \new_[15884]_  = A167 & \new_[15883]_ ;
  assign \new_[15885]_  = \new_[15884]_  & \new_[15879]_ ;
  assign \new_[15888]_  = ~A232 & ~A201;
  assign \new_[15892]_  = A266 & ~A265;
  assign \new_[15893]_  = A233 & \new_[15892]_ ;
  assign \new_[15894]_  = \new_[15893]_  & \new_[15888]_ ;
  assign \new_[15897]_  = ~A169 & A170;
  assign \new_[15901]_  = ~A199 & ~A166;
  assign \new_[15902]_  = A167 & \new_[15901]_ ;
  assign \new_[15903]_  = \new_[15902]_  & \new_[15897]_ ;
  assign \new_[15906]_  = ~A232 & ~A200;
  assign \new_[15910]_  = A299 & ~A298;
  assign \new_[15911]_  = A233 & \new_[15910]_ ;
  assign \new_[15912]_  = \new_[15911]_  & \new_[15906]_ ;
  assign \new_[15915]_  = ~A169 & A170;
  assign \new_[15919]_  = ~A199 & ~A166;
  assign \new_[15920]_  = A167 & \new_[15919]_ ;
  assign \new_[15921]_  = \new_[15920]_  & \new_[15915]_ ;
  assign \new_[15924]_  = ~A232 & ~A200;
  assign \new_[15928]_  = A266 & ~A265;
  assign \new_[15929]_  = A233 & \new_[15928]_ ;
  assign \new_[15930]_  = \new_[15929]_  & \new_[15924]_ ;
  assign \new_[15933]_  = ~A169 & A170;
  assign \new_[15937]_  = A199 & A166;
  assign \new_[15938]_  = ~A167 & \new_[15937]_ ;
  assign \new_[15939]_  = \new_[15938]_  & \new_[15933]_ ;
  assign \new_[15942]_  = ~A232 & A200;
  assign \new_[15946]_  = A299 & ~A298;
  assign \new_[15947]_  = A233 & \new_[15946]_ ;
  assign \new_[15948]_  = \new_[15947]_  & \new_[15942]_ ;
  assign \new_[15951]_  = ~A169 & A170;
  assign \new_[15955]_  = A199 & A166;
  assign \new_[15956]_  = ~A167 & \new_[15955]_ ;
  assign \new_[15957]_  = \new_[15956]_  & \new_[15951]_ ;
  assign \new_[15960]_  = ~A232 & A200;
  assign \new_[15964]_  = A266 & ~A265;
  assign \new_[15965]_  = A233 & \new_[15964]_ ;
  assign \new_[15966]_  = \new_[15965]_  & \new_[15960]_ ;
  assign \new_[15969]_  = ~A169 & A170;
  assign \new_[15973]_  = ~A200 & A166;
  assign \new_[15974]_  = ~A167 & \new_[15973]_ ;
  assign \new_[15975]_  = \new_[15974]_  & \new_[15969]_ ;
  assign \new_[15978]_  = ~A232 & ~A201;
  assign \new_[15982]_  = A299 & ~A298;
  assign \new_[15983]_  = A233 & \new_[15982]_ ;
  assign \new_[15984]_  = \new_[15983]_  & \new_[15978]_ ;
  assign \new_[15987]_  = ~A169 & A170;
  assign \new_[15991]_  = ~A200 & A166;
  assign \new_[15992]_  = ~A167 & \new_[15991]_ ;
  assign \new_[15993]_  = \new_[15992]_  & \new_[15987]_ ;
  assign \new_[15996]_  = ~A232 & ~A201;
  assign \new_[16000]_  = A266 & ~A265;
  assign \new_[16001]_  = A233 & \new_[16000]_ ;
  assign \new_[16002]_  = \new_[16001]_  & \new_[15996]_ ;
  assign \new_[16005]_  = ~A169 & A170;
  assign \new_[16009]_  = ~A199 & A166;
  assign \new_[16010]_  = ~A167 & \new_[16009]_ ;
  assign \new_[16011]_  = \new_[16010]_  & \new_[16005]_ ;
  assign \new_[16014]_  = ~A232 & ~A200;
  assign \new_[16018]_  = A299 & ~A298;
  assign \new_[16019]_  = A233 & \new_[16018]_ ;
  assign \new_[16020]_  = \new_[16019]_  & \new_[16014]_ ;
  assign \new_[16023]_  = ~A169 & A170;
  assign \new_[16027]_  = ~A199 & A166;
  assign \new_[16028]_  = ~A167 & \new_[16027]_ ;
  assign \new_[16029]_  = \new_[16028]_  & \new_[16023]_ ;
  assign \new_[16032]_  = ~A232 & ~A200;
  assign \new_[16036]_  = A266 & ~A265;
  assign \new_[16037]_  = A233 & \new_[16036]_ ;
  assign \new_[16038]_  = \new_[16037]_  & \new_[16032]_ ;
  assign \new_[16041]_  = A166 & A168;
  assign \new_[16045]_  = A232 & A200;
  assign \new_[16046]_  = A199 & \new_[16045]_ ;
  assign \new_[16047]_  = \new_[16046]_  & \new_[16041]_ ;
  assign \new_[16051]_  = ~A268 & A265;
  assign \new_[16052]_  = A233 & \new_[16051]_ ;
  assign \new_[16056]_  = ~A300 & ~A299;
  assign \new_[16057]_  = ~A269 & \new_[16056]_ ;
  assign \new_[16058]_  = \new_[16057]_  & \new_[16052]_ ;
  assign \new_[16061]_  = A166 & A168;
  assign \new_[16065]_  = A232 & A200;
  assign \new_[16066]_  = A199 & \new_[16065]_ ;
  assign \new_[16067]_  = \new_[16066]_  & \new_[16061]_ ;
  assign \new_[16071]_  = ~A268 & A265;
  assign \new_[16072]_  = A233 & \new_[16071]_ ;
  assign \new_[16076]_  = A299 & A298;
  assign \new_[16077]_  = ~A269 & \new_[16076]_ ;
  assign \new_[16078]_  = \new_[16077]_  & \new_[16072]_ ;
  assign \new_[16081]_  = A166 & A168;
  assign \new_[16085]_  = A232 & A200;
  assign \new_[16086]_  = A199 & \new_[16085]_ ;
  assign \new_[16087]_  = \new_[16086]_  & \new_[16081]_ ;
  assign \new_[16091]_  = ~A268 & A265;
  assign \new_[16092]_  = A233 & \new_[16091]_ ;
  assign \new_[16096]_  = ~A299 & ~A298;
  assign \new_[16097]_  = ~A269 & \new_[16096]_ ;
  assign \new_[16098]_  = \new_[16097]_  & \new_[16092]_ ;
  assign \new_[16101]_  = A166 & A168;
  assign \new_[16105]_  = A232 & A200;
  assign \new_[16106]_  = A199 & \new_[16105]_ ;
  assign \new_[16107]_  = \new_[16106]_  & \new_[16101]_ ;
  assign \new_[16111]_  = ~A267 & A265;
  assign \new_[16112]_  = A233 & \new_[16111]_ ;
  assign \new_[16116]_  = ~A302 & ~A301;
  assign \new_[16117]_  = ~A299 & \new_[16116]_ ;
  assign \new_[16118]_  = \new_[16117]_  & \new_[16112]_ ;
  assign \new_[16121]_  = A166 & A168;
  assign \new_[16125]_  = A232 & A200;
  assign \new_[16126]_  = A199 & \new_[16125]_ ;
  assign \new_[16127]_  = \new_[16126]_  & \new_[16121]_ ;
  assign \new_[16131]_  = A266 & A265;
  assign \new_[16132]_  = A233 & \new_[16131]_ ;
  assign \new_[16136]_  = ~A302 & ~A301;
  assign \new_[16137]_  = ~A299 & \new_[16136]_ ;
  assign \new_[16138]_  = \new_[16137]_  & \new_[16132]_ ;
  assign \new_[16141]_  = A166 & A168;
  assign \new_[16145]_  = A232 & A200;
  assign \new_[16146]_  = A199 & \new_[16145]_ ;
  assign \new_[16147]_  = \new_[16146]_  & \new_[16141]_ ;
  assign \new_[16151]_  = ~A266 & ~A265;
  assign \new_[16152]_  = A233 & \new_[16151]_ ;
  assign \new_[16156]_  = ~A302 & ~A301;
  assign \new_[16157]_  = ~A299 & \new_[16156]_ ;
  assign \new_[16158]_  = \new_[16157]_  & \new_[16152]_ ;
  assign \new_[16161]_  = A166 & A168;
  assign \new_[16165]_  = ~A233 & A200;
  assign \new_[16166]_  = A199 & \new_[16165]_ ;
  assign \new_[16167]_  = \new_[16166]_  & \new_[16161]_ ;
  assign \new_[16171]_  = A265 & ~A236;
  assign \new_[16172]_  = ~A235 & \new_[16171]_ ;
  assign \new_[16176]_  = ~A300 & A298;
  assign \new_[16177]_  = A266 & \new_[16176]_ ;
  assign \new_[16178]_  = \new_[16177]_  & \new_[16172]_ ;
  assign \new_[16181]_  = A166 & A168;
  assign \new_[16185]_  = ~A233 & A200;
  assign \new_[16186]_  = A199 & \new_[16185]_ ;
  assign \new_[16187]_  = \new_[16186]_  & \new_[16181]_ ;
  assign \new_[16191]_  = A265 & ~A236;
  assign \new_[16192]_  = ~A235 & \new_[16191]_ ;
  assign \new_[16196]_  = A299 & A298;
  assign \new_[16197]_  = A266 & \new_[16196]_ ;
  assign \new_[16198]_  = \new_[16197]_  & \new_[16192]_ ;
  assign \new_[16201]_  = A166 & A168;
  assign \new_[16205]_  = ~A233 & A200;
  assign \new_[16206]_  = A199 & \new_[16205]_ ;
  assign \new_[16207]_  = \new_[16206]_  & \new_[16201]_ ;
  assign \new_[16211]_  = A265 & ~A236;
  assign \new_[16212]_  = ~A235 & \new_[16211]_ ;
  assign \new_[16216]_  = ~A299 & ~A298;
  assign \new_[16217]_  = A266 & \new_[16216]_ ;
  assign \new_[16218]_  = \new_[16217]_  & \new_[16212]_ ;
  assign \new_[16221]_  = A166 & A168;
  assign \new_[16225]_  = ~A233 & A200;
  assign \new_[16226]_  = A199 & \new_[16225]_ ;
  assign \new_[16227]_  = \new_[16226]_  & \new_[16221]_ ;
  assign \new_[16231]_  = ~A266 & ~A236;
  assign \new_[16232]_  = ~A235 & \new_[16231]_ ;
  assign \new_[16236]_  = ~A300 & A298;
  assign \new_[16237]_  = ~A267 & \new_[16236]_ ;
  assign \new_[16238]_  = \new_[16237]_  & \new_[16232]_ ;
  assign \new_[16241]_  = A166 & A168;
  assign \new_[16245]_  = ~A233 & A200;
  assign \new_[16246]_  = A199 & \new_[16245]_ ;
  assign \new_[16247]_  = \new_[16246]_  & \new_[16241]_ ;
  assign \new_[16251]_  = ~A266 & ~A236;
  assign \new_[16252]_  = ~A235 & \new_[16251]_ ;
  assign \new_[16256]_  = A299 & A298;
  assign \new_[16257]_  = ~A267 & \new_[16256]_ ;
  assign \new_[16258]_  = \new_[16257]_  & \new_[16252]_ ;
  assign \new_[16261]_  = A166 & A168;
  assign \new_[16265]_  = ~A233 & A200;
  assign \new_[16266]_  = A199 & \new_[16265]_ ;
  assign \new_[16267]_  = \new_[16266]_  & \new_[16261]_ ;
  assign \new_[16271]_  = ~A266 & ~A236;
  assign \new_[16272]_  = ~A235 & \new_[16271]_ ;
  assign \new_[16276]_  = ~A299 & ~A298;
  assign \new_[16277]_  = ~A267 & \new_[16276]_ ;
  assign \new_[16278]_  = \new_[16277]_  & \new_[16272]_ ;
  assign \new_[16281]_  = A166 & A168;
  assign \new_[16285]_  = ~A233 & A200;
  assign \new_[16286]_  = A199 & \new_[16285]_ ;
  assign \new_[16287]_  = \new_[16286]_  & \new_[16281]_ ;
  assign \new_[16291]_  = ~A265 & ~A236;
  assign \new_[16292]_  = ~A235 & \new_[16291]_ ;
  assign \new_[16296]_  = ~A300 & A298;
  assign \new_[16297]_  = ~A266 & \new_[16296]_ ;
  assign \new_[16298]_  = \new_[16297]_  & \new_[16292]_ ;
  assign \new_[16301]_  = A166 & A168;
  assign \new_[16305]_  = ~A233 & A200;
  assign \new_[16306]_  = A199 & \new_[16305]_ ;
  assign \new_[16307]_  = \new_[16306]_  & \new_[16301]_ ;
  assign \new_[16311]_  = ~A265 & ~A236;
  assign \new_[16312]_  = ~A235 & \new_[16311]_ ;
  assign \new_[16316]_  = A299 & A298;
  assign \new_[16317]_  = ~A266 & \new_[16316]_ ;
  assign \new_[16318]_  = \new_[16317]_  & \new_[16312]_ ;
  assign \new_[16321]_  = A166 & A168;
  assign \new_[16325]_  = ~A233 & A200;
  assign \new_[16326]_  = A199 & \new_[16325]_ ;
  assign \new_[16327]_  = \new_[16326]_  & \new_[16321]_ ;
  assign \new_[16331]_  = ~A265 & ~A236;
  assign \new_[16332]_  = ~A235 & \new_[16331]_ ;
  assign \new_[16336]_  = ~A299 & ~A298;
  assign \new_[16337]_  = ~A266 & \new_[16336]_ ;
  assign \new_[16338]_  = \new_[16337]_  & \new_[16332]_ ;
  assign \new_[16341]_  = A166 & A168;
  assign \new_[16345]_  = ~A233 & A200;
  assign \new_[16346]_  = A199 & \new_[16345]_ ;
  assign \new_[16347]_  = \new_[16346]_  & \new_[16341]_ ;
  assign \new_[16351]_  = A266 & A265;
  assign \new_[16352]_  = ~A234 & \new_[16351]_ ;
  assign \new_[16356]_  = ~A302 & ~A301;
  assign \new_[16357]_  = A298 & \new_[16356]_ ;
  assign \new_[16358]_  = \new_[16357]_  & \new_[16352]_ ;
  assign \new_[16361]_  = A166 & A168;
  assign \new_[16365]_  = ~A233 & A200;
  assign \new_[16366]_  = A199 & \new_[16365]_ ;
  assign \new_[16367]_  = \new_[16366]_  & \new_[16361]_ ;
  assign \new_[16371]_  = ~A268 & ~A266;
  assign \new_[16372]_  = ~A234 & \new_[16371]_ ;
  assign \new_[16376]_  = ~A300 & A298;
  assign \new_[16377]_  = ~A269 & \new_[16376]_ ;
  assign \new_[16378]_  = \new_[16377]_  & \new_[16372]_ ;
  assign \new_[16381]_  = A166 & A168;
  assign \new_[16385]_  = ~A233 & A200;
  assign \new_[16386]_  = A199 & \new_[16385]_ ;
  assign \new_[16387]_  = \new_[16386]_  & \new_[16381]_ ;
  assign \new_[16391]_  = ~A268 & ~A266;
  assign \new_[16392]_  = ~A234 & \new_[16391]_ ;
  assign \new_[16396]_  = A299 & A298;
  assign \new_[16397]_  = ~A269 & \new_[16396]_ ;
  assign \new_[16398]_  = \new_[16397]_  & \new_[16392]_ ;
  assign \new_[16401]_  = A166 & A168;
  assign \new_[16405]_  = ~A233 & A200;
  assign \new_[16406]_  = A199 & \new_[16405]_ ;
  assign \new_[16407]_  = \new_[16406]_  & \new_[16401]_ ;
  assign \new_[16411]_  = ~A268 & ~A266;
  assign \new_[16412]_  = ~A234 & \new_[16411]_ ;
  assign \new_[16416]_  = ~A299 & ~A298;
  assign \new_[16417]_  = ~A269 & \new_[16416]_ ;
  assign \new_[16418]_  = \new_[16417]_  & \new_[16412]_ ;
  assign \new_[16421]_  = A166 & A168;
  assign \new_[16425]_  = ~A233 & A200;
  assign \new_[16426]_  = A199 & \new_[16425]_ ;
  assign \new_[16427]_  = \new_[16426]_  & \new_[16421]_ ;
  assign \new_[16431]_  = ~A267 & ~A266;
  assign \new_[16432]_  = ~A234 & \new_[16431]_ ;
  assign \new_[16436]_  = ~A302 & ~A301;
  assign \new_[16437]_  = A298 & \new_[16436]_ ;
  assign \new_[16438]_  = \new_[16437]_  & \new_[16432]_ ;
  assign \new_[16441]_  = A166 & A168;
  assign \new_[16445]_  = ~A233 & A200;
  assign \new_[16446]_  = A199 & \new_[16445]_ ;
  assign \new_[16447]_  = \new_[16446]_  & \new_[16441]_ ;
  assign \new_[16451]_  = ~A266 & ~A265;
  assign \new_[16452]_  = ~A234 & \new_[16451]_ ;
  assign \new_[16456]_  = ~A302 & ~A301;
  assign \new_[16457]_  = A298 & \new_[16456]_ ;
  assign \new_[16458]_  = \new_[16457]_  & \new_[16452]_ ;
  assign \new_[16461]_  = A166 & A168;
  assign \new_[16465]_  = ~A232 & A200;
  assign \new_[16466]_  = A199 & \new_[16465]_ ;
  assign \new_[16467]_  = \new_[16466]_  & \new_[16461]_ ;
  assign \new_[16471]_  = A266 & A265;
  assign \new_[16472]_  = ~A233 & \new_[16471]_ ;
  assign \new_[16476]_  = ~A302 & ~A301;
  assign \new_[16477]_  = A298 & \new_[16476]_ ;
  assign \new_[16478]_  = \new_[16477]_  & \new_[16472]_ ;
  assign \new_[16481]_  = A166 & A168;
  assign \new_[16485]_  = ~A232 & A200;
  assign \new_[16486]_  = A199 & \new_[16485]_ ;
  assign \new_[16487]_  = \new_[16486]_  & \new_[16481]_ ;
  assign \new_[16491]_  = ~A268 & ~A266;
  assign \new_[16492]_  = ~A233 & \new_[16491]_ ;
  assign \new_[16496]_  = ~A300 & A298;
  assign \new_[16497]_  = ~A269 & \new_[16496]_ ;
  assign \new_[16498]_  = \new_[16497]_  & \new_[16492]_ ;
  assign \new_[16501]_  = A166 & A168;
  assign \new_[16505]_  = ~A232 & A200;
  assign \new_[16506]_  = A199 & \new_[16505]_ ;
  assign \new_[16507]_  = \new_[16506]_  & \new_[16501]_ ;
  assign \new_[16511]_  = ~A268 & ~A266;
  assign \new_[16512]_  = ~A233 & \new_[16511]_ ;
  assign \new_[16516]_  = A299 & A298;
  assign \new_[16517]_  = ~A269 & \new_[16516]_ ;
  assign \new_[16518]_  = \new_[16517]_  & \new_[16512]_ ;
  assign \new_[16521]_  = A166 & A168;
  assign \new_[16525]_  = ~A232 & A200;
  assign \new_[16526]_  = A199 & \new_[16525]_ ;
  assign \new_[16527]_  = \new_[16526]_  & \new_[16521]_ ;
  assign \new_[16531]_  = ~A268 & ~A266;
  assign \new_[16532]_  = ~A233 & \new_[16531]_ ;
  assign \new_[16536]_  = ~A299 & ~A298;
  assign \new_[16537]_  = ~A269 & \new_[16536]_ ;
  assign \new_[16538]_  = \new_[16537]_  & \new_[16532]_ ;
  assign \new_[16541]_  = A166 & A168;
  assign \new_[16545]_  = ~A232 & A200;
  assign \new_[16546]_  = A199 & \new_[16545]_ ;
  assign \new_[16547]_  = \new_[16546]_  & \new_[16541]_ ;
  assign \new_[16551]_  = ~A267 & ~A266;
  assign \new_[16552]_  = ~A233 & \new_[16551]_ ;
  assign \new_[16556]_  = ~A302 & ~A301;
  assign \new_[16557]_  = A298 & \new_[16556]_ ;
  assign \new_[16558]_  = \new_[16557]_  & \new_[16552]_ ;
  assign \new_[16561]_  = A166 & A168;
  assign \new_[16565]_  = ~A232 & A200;
  assign \new_[16566]_  = A199 & \new_[16565]_ ;
  assign \new_[16567]_  = \new_[16566]_  & \new_[16561]_ ;
  assign \new_[16571]_  = ~A266 & ~A265;
  assign \new_[16572]_  = ~A233 & \new_[16571]_ ;
  assign \new_[16576]_  = ~A302 & ~A301;
  assign \new_[16577]_  = A298 & \new_[16576]_ ;
  assign \new_[16578]_  = \new_[16577]_  & \new_[16572]_ ;
  assign \new_[16581]_  = A166 & A168;
  assign \new_[16585]_  = ~A203 & ~A202;
  assign \new_[16586]_  = ~A200 & \new_[16585]_ ;
  assign \new_[16587]_  = \new_[16586]_  & \new_[16581]_ ;
  assign \new_[16591]_  = A265 & A233;
  assign \new_[16592]_  = A232 & \new_[16591]_ ;
  assign \new_[16596]_  = ~A300 & ~A299;
  assign \new_[16597]_  = ~A267 & \new_[16596]_ ;
  assign \new_[16598]_  = \new_[16597]_  & \new_[16592]_ ;
  assign \new_[16601]_  = A166 & A168;
  assign \new_[16605]_  = ~A203 & ~A202;
  assign \new_[16606]_  = ~A200 & \new_[16605]_ ;
  assign \new_[16607]_  = \new_[16606]_  & \new_[16601]_ ;
  assign \new_[16611]_  = A265 & A233;
  assign \new_[16612]_  = A232 & \new_[16611]_ ;
  assign \new_[16616]_  = A299 & A298;
  assign \new_[16617]_  = ~A267 & \new_[16616]_ ;
  assign \new_[16618]_  = \new_[16617]_  & \new_[16612]_ ;
  assign \new_[16621]_  = A166 & A168;
  assign \new_[16625]_  = ~A203 & ~A202;
  assign \new_[16626]_  = ~A200 & \new_[16625]_ ;
  assign \new_[16627]_  = \new_[16626]_  & \new_[16621]_ ;
  assign \new_[16631]_  = A265 & A233;
  assign \new_[16632]_  = A232 & \new_[16631]_ ;
  assign \new_[16636]_  = ~A299 & ~A298;
  assign \new_[16637]_  = ~A267 & \new_[16636]_ ;
  assign \new_[16638]_  = \new_[16637]_  & \new_[16632]_ ;
  assign \new_[16641]_  = A166 & A168;
  assign \new_[16645]_  = ~A203 & ~A202;
  assign \new_[16646]_  = ~A200 & \new_[16645]_ ;
  assign \new_[16647]_  = \new_[16646]_  & \new_[16641]_ ;
  assign \new_[16651]_  = A265 & A233;
  assign \new_[16652]_  = A232 & \new_[16651]_ ;
  assign \new_[16656]_  = ~A300 & ~A299;
  assign \new_[16657]_  = A266 & \new_[16656]_ ;
  assign \new_[16658]_  = \new_[16657]_  & \new_[16652]_ ;
  assign \new_[16661]_  = A166 & A168;
  assign \new_[16665]_  = ~A203 & ~A202;
  assign \new_[16666]_  = ~A200 & \new_[16665]_ ;
  assign \new_[16667]_  = \new_[16666]_  & \new_[16661]_ ;
  assign \new_[16671]_  = A265 & A233;
  assign \new_[16672]_  = A232 & \new_[16671]_ ;
  assign \new_[16676]_  = A299 & A298;
  assign \new_[16677]_  = A266 & \new_[16676]_ ;
  assign \new_[16678]_  = \new_[16677]_  & \new_[16672]_ ;
  assign \new_[16681]_  = A166 & A168;
  assign \new_[16685]_  = ~A203 & ~A202;
  assign \new_[16686]_  = ~A200 & \new_[16685]_ ;
  assign \new_[16687]_  = \new_[16686]_  & \new_[16681]_ ;
  assign \new_[16691]_  = A265 & A233;
  assign \new_[16692]_  = A232 & \new_[16691]_ ;
  assign \new_[16696]_  = ~A299 & ~A298;
  assign \new_[16697]_  = A266 & \new_[16696]_ ;
  assign \new_[16698]_  = \new_[16697]_  & \new_[16692]_ ;
  assign \new_[16701]_  = A166 & A168;
  assign \new_[16705]_  = ~A203 & ~A202;
  assign \new_[16706]_  = ~A200 & \new_[16705]_ ;
  assign \new_[16707]_  = \new_[16706]_  & \new_[16701]_ ;
  assign \new_[16711]_  = ~A265 & A233;
  assign \new_[16712]_  = A232 & \new_[16711]_ ;
  assign \new_[16716]_  = ~A300 & ~A299;
  assign \new_[16717]_  = ~A266 & \new_[16716]_ ;
  assign \new_[16718]_  = \new_[16717]_  & \new_[16712]_ ;
  assign \new_[16721]_  = A166 & A168;
  assign \new_[16725]_  = ~A203 & ~A202;
  assign \new_[16726]_  = ~A200 & \new_[16725]_ ;
  assign \new_[16727]_  = \new_[16726]_  & \new_[16721]_ ;
  assign \new_[16731]_  = ~A265 & A233;
  assign \new_[16732]_  = A232 & \new_[16731]_ ;
  assign \new_[16736]_  = A299 & A298;
  assign \new_[16737]_  = ~A266 & \new_[16736]_ ;
  assign \new_[16738]_  = \new_[16737]_  & \new_[16732]_ ;
  assign \new_[16741]_  = A166 & A168;
  assign \new_[16745]_  = ~A203 & ~A202;
  assign \new_[16746]_  = ~A200 & \new_[16745]_ ;
  assign \new_[16747]_  = \new_[16746]_  & \new_[16741]_ ;
  assign \new_[16751]_  = ~A265 & A233;
  assign \new_[16752]_  = A232 & \new_[16751]_ ;
  assign \new_[16756]_  = ~A299 & ~A298;
  assign \new_[16757]_  = ~A266 & \new_[16756]_ ;
  assign \new_[16758]_  = \new_[16757]_  & \new_[16752]_ ;
  assign \new_[16761]_  = A166 & A168;
  assign \new_[16765]_  = ~A203 & ~A202;
  assign \new_[16766]_  = ~A200 & \new_[16765]_ ;
  assign \new_[16767]_  = \new_[16766]_  & \new_[16761]_ ;
  assign \new_[16771]_  = A298 & A233;
  assign \new_[16772]_  = ~A232 & \new_[16771]_ ;
  assign \new_[16776]_  = A301 & A300;
  assign \new_[16777]_  = ~A299 & \new_[16776]_ ;
  assign \new_[16778]_  = \new_[16777]_  & \new_[16772]_ ;
  assign \new_[16781]_  = A166 & A168;
  assign \new_[16785]_  = ~A203 & ~A202;
  assign \new_[16786]_  = ~A200 & \new_[16785]_ ;
  assign \new_[16787]_  = \new_[16786]_  & \new_[16781]_ ;
  assign \new_[16791]_  = A298 & A233;
  assign \new_[16792]_  = ~A232 & \new_[16791]_ ;
  assign \new_[16796]_  = A302 & A300;
  assign \new_[16797]_  = ~A299 & \new_[16796]_ ;
  assign \new_[16798]_  = \new_[16797]_  & \new_[16792]_ ;
  assign \new_[16801]_  = A166 & A168;
  assign \new_[16805]_  = ~A203 & ~A202;
  assign \new_[16806]_  = ~A200 & \new_[16805]_ ;
  assign \new_[16807]_  = \new_[16806]_  & \new_[16801]_ ;
  assign \new_[16811]_  = A265 & A233;
  assign \new_[16812]_  = ~A232 & \new_[16811]_ ;
  assign \new_[16816]_  = A268 & A267;
  assign \new_[16817]_  = ~A266 & \new_[16816]_ ;
  assign \new_[16818]_  = \new_[16817]_  & \new_[16812]_ ;
  assign \new_[16821]_  = A166 & A168;
  assign \new_[16825]_  = ~A203 & ~A202;
  assign \new_[16826]_  = ~A200 & \new_[16825]_ ;
  assign \new_[16827]_  = \new_[16826]_  & \new_[16821]_ ;
  assign \new_[16831]_  = A265 & A233;
  assign \new_[16832]_  = ~A232 & \new_[16831]_ ;
  assign \new_[16836]_  = A269 & A267;
  assign \new_[16837]_  = ~A266 & \new_[16836]_ ;
  assign \new_[16838]_  = \new_[16837]_  & \new_[16832]_ ;
  assign \new_[16841]_  = A166 & A168;
  assign \new_[16845]_  = ~A203 & ~A202;
  assign \new_[16846]_  = ~A200 & \new_[16845]_ ;
  assign \new_[16847]_  = \new_[16846]_  & \new_[16841]_ ;
  assign \new_[16851]_  = A265 & ~A234;
  assign \new_[16852]_  = ~A233 & \new_[16851]_ ;
  assign \new_[16856]_  = ~A300 & A298;
  assign \new_[16857]_  = A266 & \new_[16856]_ ;
  assign \new_[16858]_  = \new_[16857]_  & \new_[16852]_ ;
  assign \new_[16861]_  = A166 & A168;
  assign \new_[16865]_  = ~A203 & ~A202;
  assign \new_[16866]_  = ~A200 & \new_[16865]_ ;
  assign \new_[16867]_  = \new_[16866]_  & \new_[16861]_ ;
  assign \new_[16871]_  = A265 & ~A234;
  assign \new_[16872]_  = ~A233 & \new_[16871]_ ;
  assign \new_[16876]_  = A299 & A298;
  assign \new_[16877]_  = A266 & \new_[16876]_ ;
  assign \new_[16878]_  = \new_[16877]_  & \new_[16872]_ ;
  assign \new_[16881]_  = A166 & A168;
  assign \new_[16885]_  = ~A203 & ~A202;
  assign \new_[16886]_  = ~A200 & \new_[16885]_ ;
  assign \new_[16887]_  = \new_[16886]_  & \new_[16881]_ ;
  assign \new_[16891]_  = A265 & ~A234;
  assign \new_[16892]_  = ~A233 & \new_[16891]_ ;
  assign \new_[16896]_  = ~A299 & ~A298;
  assign \new_[16897]_  = A266 & \new_[16896]_ ;
  assign \new_[16898]_  = \new_[16897]_  & \new_[16892]_ ;
  assign \new_[16901]_  = A166 & A168;
  assign \new_[16905]_  = ~A203 & ~A202;
  assign \new_[16906]_  = ~A200 & \new_[16905]_ ;
  assign \new_[16907]_  = \new_[16906]_  & \new_[16901]_ ;
  assign \new_[16911]_  = ~A266 & ~A234;
  assign \new_[16912]_  = ~A233 & \new_[16911]_ ;
  assign \new_[16916]_  = ~A300 & A298;
  assign \new_[16917]_  = ~A267 & \new_[16916]_ ;
  assign \new_[16918]_  = \new_[16917]_  & \new_[16912]_ ;
  assign \new_[16921]_  = A166 & A168;
  assign \new_[16925]_  = ~A203 & ~A202;
  assign \new_[16926]_  = ~A200 & \new_[16925]_ ;
  assign \new_[16927]_  = \new_[16926]_  & \new_[16921]_ ;
  assign \new_[16931]_  = ~A266 & ~A234;
  assign \new_[16932]_  = ~A233 & \new_[16931]_ ;
  assign \new_[16936]_  = A299 & A298;
  assign \new_[16937]_  = ~A267 & \new_[16936]_ ;
  assign \new_[16938]_  = \new_[16937]_  & \new_[16932]_ ;
  assign \new_[16941]_  = A166 & A168;
  assign \new_[16945]_  = ~A203 & ~A202;
  assign \new_[16946]_  = ~A200 & \new_[16945]_ ;
  assign \new_[16947]_  = \new_[16946]_  & \new_[16941]_ ;
  assign \new_[16951]_  = ~A266 & ~A234;
  assign \new_[16952]_  = ~A233 & \new_[16951]_ ;
  assign \new_[16956]_  = ~A299 & ~A298;
  assign \new_[16957]_  = ~A267 & \new_[16956]_ ;
  assign \new_[16958]_  = \new_[16957]_  & \new_[16952]_ ;
  assign \new_[16961]_  = A166 & A168;
  assign \new_[16965]_  = ~A203 & ~A202;
  assign \new_[16966]_  = ~A200 & \new_[16965]_ ;
  assign \new_[16967]_  = \new_[16966]_  & \new_[16961]_ ;
  assign \new_[16971]_  = ~A265 & ~A234;
  assign \new_[16972]_  = ~A233 & \new_[16971]_ ;
  assign \new_[16976]_  = ~A300 & A298;
  assign \new_[16977]_  = ~A266 & \new_[16976]_ ;
  assign \new_[16978]_  = \new_[16977]_  & \new_[16972]_ ;
  assign \new_[16981]_  = A166 & A168;
  assign \new_[16985]_  = ~A203 & ~A202;
  assign \new_[16986]_  = ~A200 & \new_[16985]_ ;
  assign \new_[16987]_  = \new_[16986]_  & \new_[16981]_ ;
  assign \new_[16991]_  = ~A265 & ~A234;
  assign \new_[16992]_  = ~A233 & \new_[16991]_ ;
  assign \new_[16996]_  = A299 & A298;
  assign \new_[16997]_  = ~A266 & \new_[16996]_ ;
  assign \new_[16998]_  = \new_[16997]_  & \new_[16992]_ ;
  assign \new_[17001]_  = A166 & A168;
  assign \new_[17005]_  = ~A203 & ~A202;
  assign \new_[17006]_  = ~A200 & \new_[17005]_ ;
  assign \new_[17007]_  = \new_[17006]_  & \new_[17001]_ ;
  assign \new_[17011]_  = ~A265 & ~A234;
  assign \new_[17012]_  = ~A233 & \new_[17011]_ ;
  assign \new_[17016]_  = ~A299 & ~A298;
  assign \new_[17017]_  = ~A266 & \new_[17016]_ ;
  assign \new_[17018]_  = \new_[17017]_  & \new_[17012]_ ;
  assign \new_[17021]_  = A166 & A168;
  assign \new_[17025]_  = ~A203 & ~A202;
  assign \new_[17026]_  = ~A200 & \new_[17025]_ ;
  assign \new_[17027]_  = \new_[17026]_  & \new_[17021]_ ;
  assign \new_[17031]_  = A234 & ~A233;
  assign \new_[17032]_  = A232 & \new_[17031]_ ;
  assign \new_[17036]_  = A299 & ~A298;
  assign \new_[17037]_  = A235 & \new_[17036]_ ;
  assign \new_[17038]_  = \new_[17037]_  & \new_[17032]_ ;
  assign \new_[17041]_  = A166 & A168;
  assign \new_[17045]_  = ~A203 & ~A202;
  assign \new_[17046]_  = ~A200 & \new_[17045]_ ;
  assign \new_[17047]_  = \new_[17046]_  & \new_[17041]_ ;
  assign \new_[17051]_  = A234 & ~A233;
  assign \new_[17052]_  = A232 & \new_[17051]_ ;
  assign \new_[17056]_  = A266 & ~A265;
  assign \new_[17057]_  = A235 & \new_[17056]_ ;
  assign \new_[17058]_  = \new_[17057]_  & \new_[17052]_ ;
  assign \new_[17061]_  = A166 & A168;
  assign \new_[17065]_  = ~A203 & ~A202;
  assign \new_[17066]_  = ~A200 & \new_[17065]_ ;
  assign \new_[17067]_  = \new_[17066]_  & \new_[17061]_ ;
  assign \new_[17071]_  = A234 & ~A233;
  assign \new_[17072]_  = A232 & \new_[17071]_ ;
  assign \new_[17076]_  = A299 & ~A298;
  assign \new_[17077]_  = A236 & \new_[17076]_ ;
  assign \new_[17078]_  = \new_[17077]_  & \new_[17072]_ ;
  assign \new_[17081]_  = A166 & A168;
  assign \new_[17085]_  = ~A203 & ~A202;
  assign \new_[17086]_  = ~A200 & \new_[17085]_ ;
  assign \new_[17087]_  = \new_[17086]_  & \new_[17081]_ ;
  assign \new_[17091]_  = A234 & ~A233;
  assign \new_[17092]_  = A232 & \new_[17091]_ ;
  assign \new_[17096]_  = A266 & ~A265;
  assign \new_[17097]_  = A236 & \new_[17096]_ ;
  assign \new_[17098]_  = \new_[17097]_  & \new_[17092]_ ;
  assign \new_[17101]_  = A166 & A168;
  assign \new_[17105]_  = ~A203 & ~A202;
  assign \new_[17106]_  = ~A200 & \new_[17105]_ ;
  assign \new_[17107]_  = \new_[17106]_  & \new_[17101]_ ;
  assign \new_[17111]_  = A265 & ~A233;
  assign \new_[17112]_  = ~A232 & \new_[17111]_ ;
  assign \new_[17116]_  = ~A300 & A298;
  assign \new_[17117]_  = A266 & \new_[17116]_ ;
  assign \new_[17118]_  = \new_[17117]_  & \new_[17112]_ ;
  assign \new_[17121]_  = A166 & A168;
  assign \new_[17125]_  = ~A203 & ~A202;
  assign \new_[17126]_  = ~A200 & \new_[17125]_ ;
  assign \new_[17127]_  = \new_[17126]_  & \new_[17121]_ ;
  assign \new_[17131]_  = A265 & ~A233;
  assign \new_[17132]_  = ~A232 & \new_[17131]_ ;
  assign \new_[17136]_  = A299 & A298;
  assign \new_[17137]_  = A266 & \new_[17136]_ ;
  assign \new_[17138]_  = \new_[17137]_  & \new_[17132]_ ;
  assign \new_[17141]_  = A166 & A168;
  assign \new_[17145]_  = ~A203 & ~A202;
  assign \new_[17146]_  = ~A200 & \new_[17145]_ ;
  assign \new_[17147]_  = \new_[17146]_  & \new_[17141]_ ;
  assign \new_[17151]_  = A265 & ~A233;
  assign \new_[17152]_  = ~A232 & \new_[17151]_ ;
  assign \new_[17156]_  = ~A299 & ~A298;
  assign \new_[17157]_  = A266 & \new_[17156]_ ;
  assign \new_[17158]_  = \new_[17157]_  & \new_[17152]_ ;
  assign \new_[17161]_  = A166 & A168;
  assign \new_[17165]_  = ~A203 & ~A202;
  assign \new_[17166]_  = ~A200 & \new_[17165]_ ;
  assign \new_[17167]_  = \new_[17166]_  & \new_[17161]_ ;
  assign \new_[17171]_  = ~A266 & ~A233;
  assign \new_[17172]_  = ~A232 & \new_[17171]_ ;
  assign \new_[17176]_  = ~A300 & A298;
  assign \new_[17177]_  = ~A267 & \new_[17176]_ ;
  assign \new_[17178]_  = \new_[17177]_  & \new_[17172]_ ;
  assign \new_[17181]_  = A166 & A168;
  assign \new_[17185]_  = ~A203 & ~A202;
  assign \new_[17186]_  = ~A200 & \new_[17185]_ ;
  assign \new_[17187]_  = \new_[17186]_  & \new_[17181]_ ;
  assign \new_[17191]_  = ~A266 & ~A233;
  assign \new_[17192]_  = ~A232 & \new_[17191]_ ;
  assign \new_[17196]_  = A299 & A298;
  assign \new_[17197]_  = ~A267 & \new_[17196]_ ;
  assign \new_[17198]_  = \new_[17197]_  & \new_[17192]_ ;
  assign \new_[17201]_  = A166 & A168;
  assign \new_[17205]_  = ~A203 & ~A202;
  assign \new_[17206]_  = ~A200 & \new_[17205]_ ;
  assign \new_[17207]_  = \new_[17206]_  & \new_[17201]_ ;
  assign \new_[17211]_  = ~A266 & ~A233;
  assign \new_[17212]_  = ~A232 & \new_[17211]_ ;
  assign \new_[17216]_  = ~A299 & ~A298;
  assign \new_[17217]_  = ~A267 & \new_[17216]_ ;
  assign \new_[17218]_  = \new_[17217]_  & \new_[17212]_ ;
  assign \new_[17221]_  = A166 & A168;
  assign \new_[17225]_  = ~A203 & ~A202;
  assign \new_[17226]_  = ~A200 & \new_[17225]_ ;
  assign \new_[17227]_  = \new_[17226]_  & \new_[17221]_ ;
  assign \new_[17231]_  = ~A265 & ~A233;
  assign \new_[17232]_  = ~A232 & \new_[17231]_ ;
  assign \new_[17236]_  = ~A300 & A298;
  assign \new_[17237]_  = ~A266 & \new_[17236]_ ;
  assign \new_[17238]_  = \new_[17237]_  & \new_[17232]_ ;
  assign \new_[17241]_  = A166 & A168;
  assign \new_[17245]_  = ~A203 & ~A202;
  assign \new_[17246]_  = ~A200 & \new_[17245]_ ;
  assign \new_[17247]_  = \new_[17246]_  & \new_[17241]_ ;
  assign \new_[17251]_  = ~A265 & ~A233;
  assign \new_[17252]_  = ~A232 & \new_[17251]_ ;
  assign \new_[17256]_  = A299 & A298;
  assign \new_[17257]_  = ~A266 & \new_[17256]_ ;
  assign \new_[17258]_  = \new_[17257]_  & \new_[17252]_ ;
  assign \new_[17261]_  = A166 & A168;
  assign \new_[17265]_  = ~A203 & ~A202;
  assign \new_[17266]_  = ~A200 & \new_[17265]_ ;
  assign \new_[17267]_  = \new_[17266]_  & \new_[17261]_ ;
  assign \new_[17271]_  = ~A265 & ~A233;
  assign \new_[17272]_  = ~A232 & \new_[17271]_ ;
  assign \new_[17276]_  = ~A299 & ~A298;
  assign \new_[17277]_  = ~A266 & \new_[17276]_ ;
  assign \new_[17278]_  = \new_[17277]_  & \new_[17272]_ ;
  assign \new_[17281]_  = A166 & A168;
  assign \new_[17285]_  = A232 & ~A201;
  assign \new_[17286]_  = ~A200 & \new_[17285]_ ;
  assign \new_[17287]_  = \new_[17286]_  & \new_[17281]_ ;
  assign \new_[17291]_  = ~A268 & A265;
  assign \new_[17292]_  = A233 & \new_[17291]_ ;
  assign \new_[17296]_  = ~A300 & ~A299;
  assign \new_[17297]_  = ~A269 & \new_[17296]_ ;
  assign \new_[17298]_  = \new_[17297]_  & \new_[17292]_ ;
  assign \new_[17301]_  = A166 & A168;
  assign \new_[17305]_  = A232 & ~A201;
  assign \new_[17306]_  = ~A200 & \new_[17305]_ ;
  assign \new_[17307]_  = \new_[17306]_  & \new_[17301]_ ;
  assign \new_[17311]_  = ~A268 & A265;
  assign \new_[17312]_  = A233 & \new_[17311]_ ;
  assign \new_[17316]_  = A299 & A298;
  assign \new_[17317]_  = ~A269 & \new_[17316]_ ;
  assign \new_[17318]_  = \new_[17317]_  & \new_[17312]_ ;
  assign \new_[17321]_  = A166 & A168;
  assign \new_[17325]_  = A232 & ~A201;
  assign \new_[17326]_  = ~A200 & \new_[17325]_ ;
  assign \new_[17327]_  = \new_[17326]_  & \new_[17321]_ ;
  assign \new_[17331]_  = ~A268 & A265;
  assign \new_[17332]_  = A233 & \new_[17331]_ ;
  assign \new_[17336]_  = ~A299 & ~A298;
  assign \new_[17337]_  = ~A269 & \new_[17336]_ ;
  assign \new_[17338]_  = \new_[17337]_  & \new_[17332]_ ;
  assign \new_[17341]_  = A166 & A168;
  assign \new_[17345]_  = A232 & ~A201;
  assign \new_[17346]_  = ~A200 & \new_[17345]_ ;
  assign \new_[17347]_  = \new_[17346]_  & \new_[17341]_ ;
  assign \new_[17351]_  = ~A267 & A265;
  assign \new_[17352]_  = A233 & \new_[17351]_ ;
  assign \new_[17356]_  = ~A302 & ~A301;
  assign \new_[17357]_  = ~A299 & \new_[17356]_ ;
  assign \new_[17358]_  = \new_[17357]_  & \new_[17352]_ ;
  assign \new_[17361]_  = A166 & A168;
  assign \new_[17365]_  = A232 & ~A201;
  assign \new_[17366]_  = ~A200 & \new_[17365]_ ;
  assign \new_[17367]_  = \new_[17366]_  & \new_[17361]_ ;
  assign \new_[17371]_  = A266 & A265;
  assign \new_[17372]_  = A233 & \new_[17371]_ ;
  assign \new_[17376]_  = ~A302 & ~A301;
  assign \new_[17377]_  = ~A299 & \new_[17376]_ ;
  assign \new_[17378]_  = \new_[17377]_  & \new_[17372]_ ;
  assign \new_[17381]_  = A166 & A168;
  assign \new_[17385]_  = A232 & ~A201;
  assign \new_[17386]_  = ~A200 & \new_[17385]_ ;
  assign \new_[17387]_  = \new_[17386]_  & \new_[17381]_ ;
  assign \new_[17391]_  = ~A266 & ~A265;
  assign \new_[17392]_  = A233 & \new_[17391]_ ;
  assign \new_[17396]_  = ~A302 & ~A301;
  assign \new_[17397]_  = ~A299 & \new_[17396]_ ;
  assign \new_[17398]_  = \new_[17397]_  & \new_[17392]_ ;
  assign \new_[17401]_  = A166 & A168;
  assign \new_[17405]_  = ~A233 & ~A201;
  assign \new_[17406]_  = ~A200 & \new_[17405]_ ;
  assign \new_[17407]_  = \new_[17406]_  & \new_[17401]_ ;
  assign \new_[17411]_  = A265 & ~A236;
  assign \new_[17412]_  = ~A235 & \new_[17411]_ ;
  assign \new_[17416]_  = ~A300 & A298;
  assign \new_[17417]_  = A266 & \new_[17416]_ ;
  assign \new_[17418]_  = \new_[17417]_  & \new_[17412]_ ;
  assign \new_[17421]_  = A166 & A168;
  assign \new_[17425]_  = ~A233 & ~A201;
  assign \new_[17426]_  = ~A200 & \new_[17425]_ ;
  assign \new_[17427]_  = \new_[17426]_  & \new_[17421]_ ;
  assign \new_[17431]_  = A265 & ~A236;
  assign \new_[17432]_  = ~A235 & \new_[17431]_ ;
  assign \new_[17436]_  = A299 & A298;
  assign \new_[17437]_  = A266 & \new_[17436]_ ;
  assign \new_[17438]_  = \new_[17437]_  & \new_[17432]_ ;
  assign \new_[17441]_  = A166 & A168;
  assign \new_[17445]_  = ~A233 & ~A201;
  assign \new_[17446]_  = ~A200 & \new_[17445]_ ;
  assign \new_[17447]_  = \new_[17446]_  & \new_[17441]_ ;
  assign \new_[17451]_  = A265 & ~A236;
  assign \new_[17452]_  = ~A235 & \new_[17451]_ ;
  assign \new_[17456]_  = ~A299 & ~A298;
  assign \new_[17457]_  = A266 & \new_[17456]_ ;
  assign \new_[17458]_  = \new_[17457]_  & \new_[17452]_ ;
  assign \new_[17461]_  = A166 & A168;
  assign \new_[17465]_  = ~A233 & ~A201;
  assign \new_[17466]_  = ~A200 & \new_[17465]_ ;
  assign \new_[17467]_  = \new_[17466]_  & \new_[17461]_ ;
  assign \new_[17471]_  = ~A266 & ~A236;
  assign \new_[17472]_  = ~A235 & \new_[17471]_ ;
  assign \new_[17476]_  = ~A300 & A298;
  assign \new_[17477]_  = ~A267 & \new_[17476]_ ;
  assign \new_[17478]_  = \new_[17477]_  & \new_[17472]_ ;
  assign \new_[17481]_  = A166 & A168;
  assign \new_[17485]_  = ~A233 & ~A201;
  assign \new_[17486]_  = ~A200 & \new_[17485]_ ;
  assign \new_[17487]_  = \new_[17486]_  & \new_[17481]_ ;
  assign \new_[17491]_  = ~A266 & ~A236;
  assign \new_[17492]_  = ~A235 & \new_[17491]_ ;
  assign \new_[17496]_  = A299 & A298;
  assign \new_[17497]_  = ~A267 & \new_[17496]_ ;
  assign \new_[17498]_  = \new_[17497]_  & \new_[17492]_ ;
  assign \new_[17501]_  = A166 & A168;
  assign \new_[17505]_  = ~A233 & ~A201;
  assign \new_[17506]_  = ~A200 & \new_[17505]_ ;
  assign \new_[17507]_  = \new_[17506]_  & \new_[17501]_ ;
  assign \new_[17511]_  = ~A266 & ~A236;
  assign \new_[17512]_  = ~A235 & \new_[17511]_ ;
  assign \new_[17516]_  = ~A299 & ~A298;
  assign \new_[17517]_  = ~A267 & \new_[17516]_ ;
  assign \new_[17518]_  = \new_[17517]_  & \new_[17512]_ ;
  assign \new_[17521]_  = A166 & A168;
  assign \new_[17525]_  = ~A233 & ~A201;
  assign \new_[17526]_  = ~A200 & \new_[17525]_ ;
  assign \new_[17527]_  = \new_[17526]_  & \new_[17521]_ ;
  assign \new_[17531]_  = ~A265 & ~A236;
  assign \new_[17532]_  = ~A235 & \new_[17531]_ ;
  assign \new_[17536]_  = ~A300 & A298;
  assign \new_[17537]_  = ~A266 & \new_[17536]_ ;
  assign \new_[17538]_  = \new_[17537]_  & \new_[17532]_ ;
  assign \new_[17541]_  = A166 & A168;
  assign \new_[17545]_  = ~A233 & ~A201;
  assign \new_[17546]_  = ~A200 & \new_[17545]_ ;
  assign \new_[17547]_  = \new_[17546]_  & \new_[17541]_ ;
  assign \new_[17551]_  = ~A265 & ~A236;
  assign \new_[17552]_  = ~A235 & \new_[17551]_ ;
  assign \new_[17556]_  = A299 & A298;
  assign \new_[17557]_  = ~A266 & \new_[17556]_ ;
  assign \new_[17558]_  = \new_[17557]_  & \new_[17552]_ ;
  assign \new_[17561]_  = A166 & A168;
  assign \new_[17565]_  = ~A233 & ~A201;
  assign \new_[17566]_  = ~A200 & \new_[17565]_ ;
  assign \new_[17567]_  = \new_[17566]_  & \new_[17561]_ ;
  assign \new_[17571]_  = ~A265 & ~A236;
  assign \new_[17572]_  = ~A235 & \new_[17571]_ ;
  assign \new_[17576]_  = ~A299 & ~A298;
  assign \new_[17577]_  = ~A266 & \new_[17576]_ ;
  assign \new_[17578]_  = \new_[17577]_  & \new_[17572]_ ;
  assign \new_[17581]_  = A166 & A168;
  assign \new_[17585]_  = ~A233 & ~A201;
  assign \new_[17586]_  = ~A200 & \new_[17585]_ ;
  assign \new_[17587]_  = \new_[17586]_  & \new_[17581]_ ;
  assign \new_[17591]_  = A266 & A265;
  assign \new_[17592]_  = ~A234 & \new_[17591]_ ;
  assign \new_[17596]_  = ~A302 & ~A301;
  assign \new_[17597]_  = A298 & \new_[17596]_ ;
  assign \new_[17598]_  = \new_[17597]_  & \new_[17592]_ ;
  assign \new_[17601]_  = A166 & A168;
  assign \new_[17605]_  = ~A233 & ~A201;
  assign \new_[17606]_  = ~A200 & \new_[17605]_ ;
  assign \new_[17607]_  = \new_[17606]_  & \new_[17601]_ ;
  assign \new_[17611]_  = ~A268 & ~A266;
  assign \new_[17612]_  = ~A234 & \new_[17611]_ ;
  assign \new_[17616]_  = ~A300 & A298;
  assign \new_[17617]_  = ~A269 & \new_[17616]_ ;
  assign \new_[17618]_  = \new_[17617]_  & \new_[17612]_ ;
  assign \new_[17621]_  = A166 & A168;
  assign \new_[17625]_  = ~A233 & ~A201;
  assign \new_[17626]_  = ~A200 & \new_[17625]_ ;
  assign \new_[17627]_  = \new_[17626]_  & \new_[17621]_ ;
  assign \new_[17631]_  = ~A268 & ~A266;
  assign \new_[17632]_  = ~A234 & \new_[17631]_ ;
  assign \new_[17636]_  = A299 & A298;
  assign \new_[17637]_  = ~A269 & \new_[17636]_ ;
  assign \new_[17638]_  = \new_[17637]_  & \new_[17632]_ ;
  assign \new_[17641]_  = A166 & A168;
  assign \new_[17645]_  = ~A233 & ~A201;
  assign \new_[17646]_  = ~A200 & \new_[17645]_ ;
  assign \new_[17647]_  = \new_[17646]_  & \new_[17641]_ ;
  assign \new_[17651]_  = ~A268 & ~A266;
  assign \new_[17652]_  = ~A234 & \new_[17651]_ ;
  assign \new_[17656]_  = ~A299 & ~A298;
  assign \new_[17657]_  = ~A269 & \new_[17656]_ ;
  assign \new_[17658]_  = \new_[17657]_  & \new_[17652]_ ;
  assign \new_[17661]_  = A166 & A168;
  assign \new_[17665]_  = ~A233 & ~A201;
  assign \new_[17666]_  = ~A200 & \new_[17665]_ ;
  assign \new_[17667]_  = \new_[17666]_  & \new_[17661]_ ;
  assign \new_[17671]_  = ~A267 & ~A266;
  assign \new_[17672]_  = ~A234 & \new_[17671]_ ;
  assign \new_[17676]_  = ~A302 & ~A301;
  assign \new_[17677]_  = A298 & \new_[17676]_ ;
  assign \new_[17678]_  = \new_[17677]_  & \new_[17672]_ ;
  assign \new_[17681]_  = A166 & A168;
  assign \new_[17685]_  = ~A233 & ~A201;
  assign \new_[17686]_  = ~A200 & \new_[17685]_ ;
  assign \new_[17687]_  = \new_[17686]_  & \new_[17681]_ ;
  assign \new_[17691]_  = ~A266 & ~A265;
  assign \new_[17692]_  = ~A234 & \new_[17691]_ ;
  assign \new_[17696]_  = ~A302 & ~A301;
  assign \new_[17697]_  = A298 & \new_[17696]_ ;
  assign \new_[17698]_  = \new_[17697]_  & \new_[17692]_ ;
  assign \new_[17701]_  = A166 & A168;
  assign \new_[17705]_  = ~A232 & ~A201;
  assign \new_[17706]_  = ~A200 & \new_[17705]_ ;
  assign \new_[17707]_  = \new_[17706]_  & \new_[17701]_ ;
  assign \new_[17711]_  = A266 & A265;
  assign \new_[17712]_  = ~A233 & \new_[17711]_ ;
  assign \new_[17716]_  = ~A302 & ~A301;
  assign \new_[17717]_  = A298 & \new_[17716]_ ;
  assign \new_[17718]_  = \new_[17717]_  & \new_[17712]_ ;
  assign \new_[17721]_  = A166 & A168;
  assign \new_[17725]_  = ~A232 & ~A201;
  assign \new_[17726]_  = ~A200 & \new_[17725]_ ;
  assign \new_[17727]_  = \new_[17726]_  & \new_[17721]_ ;
  assign \new_[17731]_  = ~A268 & ~A266;
  assign \new_[17732]_  = ~A233 & \new_[17731]_ ;
  assign \new_[17736]_  = ~A300 & A298;
  assign \new_[17737]_  = ~A269 & \new_[17736]_ ;
  assign \new_[17738]_  = \new_[17737]_  & \new_[17732]_ ;
  assign \new_[17741]_  = A166 & A168;
  assign \new_[17745]_  = ~A232 & ~A201;
  assign \new_[17746]_  = ~A200 & \new_[17745]_ ;
  assign \new_[17747]_  = \new_[17746]_  & \new_[17741]_ ;
  assign \new_[17751]_  = ~A268 & ~A266;
  assign \new_[17752]_  = ~A233 & \new_[17751]_ ;
  assign \new_[17756]_  = A299 & A298;
  assign \new_[17757]_  = ~A269 & \new_[17756]_ ;
  assign \new_[17758]_  = \new_[17757]_  & \new_[17752]_ ;
  assign \new_[17761]_  = A166 & A168;
  assign \new_[17765]_  = ~A232 & ~A201;
  assign \new_[17766]_  = ~A200 & \new_[17765]_ ;
  assign \new_[17767]_  = \new_[17766]_  & \new_[17761]_ ;
  assign \new_[17771]_  = ~A268 & ~A266;
  assign \new_[17772]_  = ~A233 & \new_[17771]_ ;
  assign \new_[17776]_  = ~A299 & ~A298;
  assign \new_[17777]_  = ~A269 & \new_[17776]_ ;
  assign \new_[17778]_  = \new_[17777]_  & \new_[17772]_ ;
  assign \new_[17781]_  = A166 & A168;
  assign \new_[17785]_  = ~A232 & ~A201;
  assign \new_[17786]_  = ~A200 & \new_[17785]_ ;
  assign \new_[17787]_  = \new_[17786]_  & \new_[17781]_ ;
  assign \new_[17791]_  = ~A267 & ~A266;
  assign \new_[17792]_  = ~A233 & \new_[17791]_ ;
  assign \new_[17796]_  = ~A302 & ~A301;
  assign \new_[17797]_  = A298 & \new_[17796]_ ;
  assign \new_[17798]_  = \new_[17797]_  & \new_[17792]_ ;
  assign \new_[17801]_  = A166 & A168;
  assign \new_[17805]_  = ~A232 & ~A201;
  assign \new_[17806]_  = ~A200 & \new_[17805]_ ;
  assign \new_[17807]_  = \new_[17806]_  & \new_[17801]_ ;
  assign \new_[17811]_  = ~A266 & ~A265;
  assign \new_[17812]_  = ~A233 & \new_[17811]_ ;
  assign \new_[17816]_  = ~A302 & ~A301;
  assign \new_[17817]_  = A298 & \new_[17816]_ ;
  assign \new_[17818]_  = \new_[17817]_  & \new_[17812]_ ;
  assign \new_[17821]_  = A166 & A168;
  assign \new_[17825]_  = A232 & ~A200;
  assign \new_[17826]_  = ~A199 & \new_[17825]_ ;
  assign \new_[17827]_  = \new_[17826]_  & \new_[17821]_ ;
  assign \new_[17831]_  = ~A268 & A265;
  assign \new_[17832]_  = A233 & \new_[17831]_ ;
  assign \new_[17836]_  = ~A300 & ~A299;
  assign \new_[17837]_  = ~A269 & \new_[17836]_ ;
  assign \new_[17838]_  = \new_[17837]_  & \new_[17832]_ ;
  assign \new_[17841]_  = A166 & A168;
  assign \new_[17845]_  = A232 & ~A200;
  assign \new_[17846]_  = ~A199 & \new_[17845]_ ;
  assign \new_[17847]_  = \new_[17846]_  & \new_[17841]_ ;
  assign \new_[17851]_  = ~A268 & A265;
  assign \new_[17852]_  = A233 & \new_[17851]_ ;
  assign \new_[17856]_  = A299 & A298;
  assign \new_[17857]_  = ~A269 & \new_[17856]_ ;
  assign \new_[17858]_  = \new_[17857]_  & \new_[17852]_ ;
  assign \new_[17861]_  = A166 & A168;
  assign \new_[17865]_  = A232 & ~A200;
  assign \new_[17866]_  = ~A199 & \new_[17865]_ ;
  assign \new_[17867]_  = \new_[17866]_  & \new_[17861]_ ;
  assign \new_[17871]_  = ~A268 & A265;
  assign \new_[17872]_  = A233 & \new_[17871]_ ;
  assign \new_[17876]_  = ~A299 & ~A298;
  assign \new_[17877]_  = ~A269 & \new_[17876]_ ;
  assign \new_[17878]_  = \new_[17877]_  & \new_[17872]_ ;
  assign \new_[17881]_  = A166 & A168;
  assign \new_[17885]_  = A232 & ~A200;
  assign \new_[17886]_  = ~A199 & \new_[17885]_ ;
  assign \new_[17887]_  = \new_[17886]_  & \new_[17881]_ ;
  assign \new_[17891]_  = ~A267 & A265;
  assign \new_[17892]_  = A233 & \new_[17891]_ ;
  assign \new_[17896]_  = ~A302 & ~A301;
  assign \new_[17897]_  = ~A299 & \new_[17896]_ ;
  assign \new_[17898]_  = \new_[17897]_  & \new_[17892]_ ;
  assign \new_[17901]_  = A166 & A168;
  assign \new_[17905]_  = A232 & ~A200;
  assign \new_[17906]_  = ~A199 & \new_[17905]_ ;
  assign \new_[17907]_  = \new_[17906]_  & \new_[17901]_ ;
  assign \new_[17911]_  = A266 & A265;
  assign \new_[17912]_  = A233 & \new_[17911]_ ;
  assign \new_[17916]_  = ~A302 & ~A301;
  assign \new_[17917]_  = ~A299 & \new_[17916]_ ;
  assign \new_[17918]_  = \new_[17917]_  & \new_[17912]_ ;
  assign \new_[17921]_  = A166 & A168;
  assign \new_[17925]_  = A232 & ~A200;
  assign \new_[17926]_  = ~A199 & \new_[17925]_ ;
  assign \new_[17927]_  = \new_[17926]_  & \new_[17921]_ ;
  assign \new_[17931]_  = ~A266 & ~A265;
  assign \new_[17932]_  = A233 & \new_[17931]_ ;
  assign \new_[17936]_  = ~A302 & ~A301;
  assign \new_[17937]_  = ~A299 & \new_[17936]_ ;
  assign \new_[17938]_  = \new_[17937]_  & \new_[17932]_ ;
  assign \new_[17941]_  = A166 & A168;
  assign \new_[17945]_  = ~A233 & ~A200;
  assign \new_[17946]_  = ~A199 & \new_[17945]_ ;
  assign \new_[17947]_  = \new_[17946]_  & \new_[17941]_ ;
  assign \new_[17951]_  = A265 & ~A236;
  assign \new_[17952]_  = ~A235 & \new_[17951]_ ;
  assign \new_[17956]_  = ~A300 & A298;
  assign \new_[17957]_  = A266 & \new_[17956]_ ;
  assign \new_[17958]_  = \new_[17957]_  & \new_[17952]_ ;
  assign \new_[17961]_  = A166 & A168;
  assign \new_[17965]_  = ~A233 & ~A200;
  assign \new_[17966]_  = ~A199 & \new_[17965]_ ;
  assign \new_[17967]_  = \new_[17966]_  & \new_[17961]_ ;
  assign \new_[17971]_  = A265 & ~A236;
  assign \new_[17972]_  = ~A235 & \new_[17971]_ ;
  assign \new_[17976]_  = A299 & A298;
  assign \new_[17977]_  = A266 & \new_[17976]_ ;
  assign \new_[17978]_  = \new_[17977]_  & \new_[17972]_ ;
  assign \new_[17981]_  = A166 & A168;
  assign \new_[17985]_  = ~A233 & ~A200;
  assign \new_[17986]_  = ~A199 & \new_[17985]_ ;
  assign \new_[17987]_  = \new_[17986]_  & \new_[17981]_ ;
  assign \new_[17991]_  = A265 & ~A236;
  assign \new_[17992]_  = ~A235 & \new_[17991]_ ;
  assign \new_[17996]_  = ~A299 & ~A298;
  assign \new_[17997]_  = A266 & \new_[17996]_ ;
  assign \new_[17998]_  = \new_[17997]_  & \new_[17992]_ ;
  assign \new_[18001]_  = A166 & A168;
  assign \new_[18005]_  = ~A233 & ~A200;
  assign \new_[18006]_  = ~A199 & \new_[18005]_ ;
  assign \new_[18007]_  = \new_[18006]_  & \new_[18001]_ ;
  assign \new_[18011]_  = ~A266 & ~A236;
  assign \new_[18012]_  = ~A235 & \new_[18011]_ ;
  assign \new_[18016]_  = ~A300 & A298;
  assign \new_[18017]_  = ~A267 & \new_[18016]_ ;
  assign \new_[18018]_  = \new_[18017]_  & \new_[18012]_ ;
  assign \new_[18021]_  = A166 & A168;
  assign \new_[18025]_  = ~A233 & ~A200;
  assign \new_[18026]_  = ~A199 & \new_[18025]_ ;
  assign \new_[18027]_  = \new_[18026]_  & \new_[18021]_ ;
  assign \new_[18031]_  = ~A266 & ~A236;
  assign \new_[18032]_  = ~A235 & \new_[18031]_ ;
  assign \new_[18036]_  = A299 & A298;
  assign \new_[18037]_  = ~A267 & \new_[18036]_ ;
  assign \new_[18038]_  = \new_[18037]_  & \new_[18032]_ ;
  assign \new_[18041]_  = A166 & A168;
  assign \new_[18045]_  = ~A233 & ~A200;
  assign \new_[18046]_  = ~A199 & \new_[18045]_ ;
  assign \new_[18047]_  = \new_[18046]_  & \new_[18041]_ ;
  assign \new_[18051]_  = ~A266 & ~A236;
  assign \new_[18052]_  = ~A235 & \new_[18051]_ ;
  assign \new_[18056]_  = ~A299 & ~A298;
  assign \new_[18057]_  = ~A267 & \new_[18056]_ ;
  assign \new_[18058]_  = \new_[18057]_  & \new_[18052]_ ;
  assign \new_[18061]_  = A166 & A168;
  assign \new_[18065]_  = ~A233 & ~A200;
  assign \new_[18066]_  = ~A199 & \new_[18065]_ ;
  assign \new_[18067]_  = \new_[18066]_  & \new_[18061]_ ;
  assign \new_[18071]_  = ~A265 & ~A236;
  assign \new_[18072]_  = ~A235 & \new_[18071]_ ;
  assign \new_[18076]_  = ~A300 & A298;
  assign \new_[18077]_  = ~A266 & \new_[18076]_ ;
  assign \new_[18078]_  = \new_[18077]_  & \new_[18072]_ ;
  assign \new_[18081]_  = A166 & A168;
  assign \new_[18085]_  = ~A233 & ~A200;
  assign \new_[18086]_  = ~A199 & \new_[18085]_ ;
  assign \new_[18087]_  = \new_[18086]_  & \new_[18081]_ ;
  assign \new_[18091]_  = ~A265 & ~A236;
  assign \new_[18092]_  = ~A235 & \new_[18091]_ ;
  assign \new_[18096]_  = A299 & A298;
  assign \new_[18097]_  = ~A266 & \new_[18096]_ ;
  assign \new_[18098]_  = \new_[18097]_  & \new_[18092]_ ;
  assign \new_[18101]_  = A166 & A168;
  assign \new_[18105]_  = ~A233 & ~A200;
  assign \new_[18106]_  = ~A199 & \new_[18105]_ ;
  assign \new_[18107]_  = \new_[18106]_  & \new_[18101]_ ;
  assign \new_[18111]_  = ~A265 & ~A236;
  assign \new_[18112]_  = ~A235 & \new_[18111]_ ;
  assign \new_[18116]_  = ~A299 & ~A298;
  assign \new_[18117]_  = ~A266 & \new_[18116]_ ;
  assign \new_[18118]_  = \new_[18117]_  & \new_[18112]_ ;
  assign \new_[18121]_  = A166 & A168;
  assign \new_[18125]_  = ~A233 & ~A200;
  assign \new_[18126]_  = ~A199 & \new_[18125]_ ;
  assign \new_[18127]_  = \new_[18126]_  & \new_[18121]_ ;
  assign \new_[18131]_  = A266 & A265;
  assign \new_[18132]_  = ~A234 & \new_[18131]_ ;
  assign \new_[18136]_  = ~A302 & ~A301;
  assign \new_[18137]_  = A298 & \new_[18136]_ ;
  assign \new_[18138]_  = \new_[18137]_  & \new_[18132]_ ;
  assign \new_[18141]_  = A166 & A168;
  assign \new_[18145]_  = ~A233 & ~A200;
  assign \new_[18146]_  = ~A199 & \new_[18145]_ ;
  assign \new_[18147]_  = \new_[18146]_  & \new_[18141]_ ;
  assign \new_[18151]_  = ~A268 & ~A266;
  assign \new_[18152]_  = ~A234 & \new_[18151]_ ;
  assign \new_[18156]_  = ~A300 & A298;
  assign \new_[18157]_  = ~A269 & \new_[18156]_ ;
  assign \new_[18158]_  = \new_[18157]_  & \new_[18152]_ ;
  assign \new_[18161]_  = A166 & A168;
  assign \new_[18165]_  = ~A233 & ~A200;
  assign \new_[18166]_  = ~A199 & \new_[18165]_ ;
  assign \new_[18167]_  = \new_[18166]_  & \new_[18161]_ ;
  assign \new_[18171]_  = ~A268 & ~A266;
  assign \new_[18172]_  = ~A234 & \new_[18171]_ ;
  assign \new_[18176]_  = A299 & A298;
  assign \new_[18177]_  = ~A269 & \new_[18176]_ ;
  assign \new_[18178]_  = \new_[18177]_  & \new_[18172]_ ;
  assign \new_[18181]_  = A166 & A168;
  assign \new_[18185]_  = ~A233 & ~A200;
  assign \new_[18186]_  = ~A199 & \new_[18185]_ ;
  assign \new_[18187]_  = \new_[18186]_  & \new_[18181]_ ;
  assign \new_[18191]_  = ~A268 & ~A266;
  assign \new_[18192]_  = ~A234 & \new_[18191]_ ;
  assign \new_[18196]_  = ~A299 & ~A298;
  assign \new_[18197]_  = ~A269 & \new_[18196]_ ;
  assign \new_[18198]_  = \new_[18197]_  & \new_[18192]_ ;
  assign \new_[18201]_  = A166 & A168;
  assign \new_[18205]_  = ~A233 & ~A200;
  assign \new_[18206]_  = ~A199 & \new_[18205]_ ;
  assign \new_[18207]_  = \new_[18206]_  & \new_[18201]_ ;
  assign \new_[18211]_  = ~A267 & ~A266;
  assign \new_[18212]_  = ~A234 & \new_[18211]_ ;
  assign \new_[18216]_  = ~A302 & ~A301;
  assign \new_[18217]_  = A298 & \new_[18216]_ ;
  assign \new_[18218]_  = \new_[18217]_  & \new_[18212]_ ;
  assign \new_[18221]_  = A166 & A168;
  assign \new_[18225]_  = ~A233 & ~A200;
  assign \new_[18226]_  = ~A199 & \new_[18225]_ ;
  assign \new_[18227]_  = \new_[18226]_  & \new_[18221]_ ;
  assign \new_[18231]_  = ~A266 & ~A265;
  assign \new_[18232]_  = ~A234 & \new_[18231]_ ;
  assign \new_[18236]_  = ~A302 & ~A301;
  assign \new_[18237]_  = A298 & \new_[18236]_ ;
  assign \new_[18238]_  = \new_[18237]_  & \new_[18232]_ ;
  assign \new_[18241]_  = A166 & A168;
  assign \new_[18245]_  = ~A232 & ~A200;
  assign \new_[18246]_  = ~A199 & \new_[18245]_ ;
  assign \new_[18247]_  = \new_[18246]_  & \new_[18241]_ ;
  assign \new_[18251]_  = A266 & A265;
  assign \new_[18252]_  = ~A233 & \new_[18251]_ ;
  assign \new_[18256]_  = ~A302 & ~A301;
  assign \new_[18257]_  = A298 & \new_[18256]_ ;
  assign \new_[18258]_  = \new_[18257]_  & \new_[18252]_ ;
  assign \new_[18261]_  = A166 & A168;
  assign \new_[18265]_  = ~A232 & ~A200;
  assign \new_[18266]_  = ~A199 & \new_[18265]_ ;
  assign \new_[18267]_  = \new_[18266]_  & \new_[18261]_ ;
  assign \new_[18271]_  = ~A268 & ~A266;
  assign \new_[18272]_  = ~A233 & \new_[18271]_ ;
  assign \new_[18276]_  = ~A300 & A298;
  assign \new_[18277]_  = ~A269 & \new_[18276]_ ;
  assign \new_[18278]_  = \new_[18277]_  & \new_[18272]_ ;
  assign \new_[18281]_  = A166 & A168;
  assign \new_[18285]_  = ~A232 & ~A200;
  assign \new_[18286]_  = ~A199 & \new_[18285]_ ;
  assign \new_[18287]_  = \new_[18286]_  & \new_[18281]_ ;
  assign \new_[18291]_  = ~A268 & ~A266;
  assign \new_[18292]_  = ~A233 & \new_[18291]_ ;
  assign \new_[18296]_  = A299 & A298;
  assign \new_[18297]_  = ~A269 & \new_[18296]_ ;
  assign \new_[18298]_  = \new_[18297]_  & \new_[18292]_ ;
  assign \new_[18301]_  = A166 & A168;
  assign \new_[18305]_  = ~A232 & ~A200;
  assign \new_[18306]_  = ~A199 & \new_[18305]_ ;
  assign \new_[18307]_  = \new_[18306]_  & \new_[18301]_ ;
  assign \new_[18311]_  = ~A268 & ~A266;
  assign \new_[18312]_  = ~A233 & \new_[18311]_ ;
  assign \new_[18316]_  = ~A299 & ~A298;
  assign \new_[18317]_  = ~A269 & \new_[18316]_ ;
  assign \new_[18318]_  = \new_[18317]_  & \new_[18312]_ ;
  assign \new_[18321]_  = A166 & A168;
  assign \new_[18325]_  = ~A232 & ~A200;
  assign \new_[18326]_  = ~A199 & \new_[18325]_ ;
  assign \new_[18327]_  = \new_[18326]_  & \new_[18321]_ ;
  assign \new_[18331]_  = ~A267 & ~A266;
  assign \new_[18332]_  = ~A233 & \new_[18331]_ ;
  assign \new_[18336]_  = ~A302 & ~A301;
  assign \new_[18337]_  = A298 & \new_[18336]_ ;
  assign \new_[18338]_  = \new_[18337]_  & \new_[18332]_ ;
  assign \new_[18341]_  = A166 & A168;
  assign \new_[18345]_  = ~A232 & ~A200;
  assign \new_[18346]_  = ~A199 & \new_[18345]_ ;
  assign \new_[18347]_  = \new_[18346]_  & \new_[18341]_ ;
  assign \new_[18351]_  = ~A266 & ~A265;
  assign \new_[18352]_  = ~A233 & \new_[18351]_ ;
  assign \new_[18356]_  = ~A302 & ~A301;
  assign \new_[18357]_  = A298 & \new_[18356]_ ;
  assign \new_[18358]_  = \new_[18357]_  & \new_[18352]_ ;
  assign \new_[18361]_  = A167 & A168;
  assign \new_[18365]_  = A232 & A200;
  assign \new_[18366]_  = A199 & \new_[18365]_ ;
  assign \new_[18367]_  = \new_[18366]_  & \new_[18361]_ ;
  assign \new_[18371]_  = ~A268 & A265;
  assign \new_[18372]_  = A233 & \new_[18371]_ ;
  assign \new_[18376]_  = ~A300 & ~A299;
  assign \new_[18377]_  = ~A269 & \new_[18376]_ ;
  assign \new_[18378]_  = \new_[18377]_  & \new_[18372]_ ;
  assign \new_[18381]_  = A167 & A168;
  assign \new_[18385]_  = A232 & A200;
  assign \new_[18386]_  = A199 & \new_[18385]_ ;
  assign \new_[18387]_  = \new_[18386]_  & \new_[18381]_ ;
  assign \new_[18391]_  = ~A268 & A265;
  assign \new_[18392]_  = A233 & \new_[18391]_ ;
  assign \new_[18396]_  = A299 & A298;
  assign \new_[18397]_  = ~A269 & \new_[18396]_ ;
  assign \new_[18398]_  = \new_[18397]_  & \new_[18392]_ ;
  assign \new_[18401]_  = A167 & A168;
  assign \new_[18405]_  = A232 & A200;
  assign \new_[18406]_  = A199 & \new_[18405]_ ;
  assign \new_[18407]_  = \new_[18406]_  & \new_[18401]_ ;
  assign \new_[18411]_  = ~A268 & A265;
  assign \new_[18412]_  = A233 & \new_[18411]_ ;
  assign \new_[18416]_  = ~A299 & ~A298;
  assign \new_[18417]_  = ~A269 & \new_[18416]_ ;
  assign \new_[18418]_  = \new_[18417]_  & \new_[18412]_ ;
  assign \new_[18421]_  = A167 & A168;
  assign \new_[18425]_  = A232 & A200;
  assign \new_[18426]_  = A199 & \new_[18425]_ ;
  assign \new_[18427]_  = \new_[18426]_  & \new_[18421]_ ;
  assign \new_[18431]_  = ~A267 & A265;
  assign \new_[18432]_  = A233 & \new_[18431]_ ;
  assign \new_[18436]_  = ~A302 & ~A301;
  assign \new_[18437]_  = ~A299 & \new_[18436]_ ;
  assign \new_[18438]_  = \new_[18437]_  & \new_[18432]_ ;
  assign \new_[18441]_  = A167 & A168;
  assign \new_[18445]_  = A232 & A200;
  assign \new_[18446]_  = A199 & \new_[18445]_ ;
  assign \new_[18447]_  = \new_[18446]_  & \new_[18441]_ ;
  assign \new_[18451]_  = A266 & A265;
  assign \new_[18452]_  = A233 & \new_[18451]_ ;
  assign \new_[18456]_  = ~A302 & ~A301;
  assign \new_[18457]_  = ~A299 & \new_[18456]_ ;
  assign \new_[18458]_  = \new_[18457]_  & \new_[18452]_ ;
  assign \new_[18461]_  = A167 & A168;
  assign \new_[18465]_  = A232 & A200;
  assign \new_[18466]_  = A199 & \new_[18465]_ ;
  assign \new_[18467]_  = \new_[18466]_  & \new_[18461]_ ;
  assign \new_[18471]_  = ~A266 & ~A265;
  assign \new_[18472]_  = A233 & \new_[18471]_ ;
  assign \new_[18476]_  = ~A302 & ~A301;
  assign \new_[18477]_  = ~A299 & \new_[18476]_ ;
  assign \new_[18478]_  = \new_[18477]_  & \new_[18472]_ ;
  assign \new_[18481]_  = A167 & A168;
  assign \new_[18485]_  = ~A233 & A200;
  assign \new_[18486]_  = A199 & \new_[18485]_ ;
  assign \new_[18487]_  = \new_[18486]_  & \new_[18481]_ ;
  assign \new_[18491]_  = A265 & ~A236;
  assign \new_[18492]_  = ~A235 & \new_[18491]_ ;
  assign \new_[18496]_  = ~A300 & A298;
  assign \new_[18497]_  = A266 & \new_[18496]_ ;
  assign \new_[18498]_  = \new_[18497]_  & \new_[18492]_ ;
  assign \new_[18501]_  = A167 & A168;
  assign \new_[18505]_  = ~A233 & A200;
  assign \new_[18506]_  = A199 & \new_[18505]_ ;
  assign \new_[18507]_  = \new_[18506]_  & \new_[18501]_ ;
  assign \new_[18511]_  = A265 & ~A236;
  assign \new_[18512]_  = ~A235 & \new_[18511]_ ;
  assign \new_[18516]_  = A299 & A298;
  assign \new_[18517]_  = A266 & \new_[18516]_ ;
  assign \new_[18518]_  = \new_[18517]_  & \new_[18512]_ ;
  assign \new_[18521]_  = A167 & A168;
  assign \new_[18525]_  = ~A233 & A200;
  assign \new_[18526]_  = A199 & \new_[18525]_ ;
  assign \new_[18527]_  = \new_[18526]_  & \new_[18521]_ ;
  assign \new_[18531]_  = A265 & ~A236;
  assign \new_[18532]_  = ~A235 & \new_[18531]_ ;
  assign \new_[18536]_  = ~A299 & ~A298;
  assign \new_[18537]_  = A266 & \new_[18536]_ ;
  assign \new_[18538]_  = \new_[18537]_  & \new_[18532]_ ;
  assign \new_[18541]_  = A167 & A168;
  assign \new_[18545]_  = ~A233 & A200;
  assign \new_[18546]_  = A199 & \new_[18545]_ ;
  assign \new_[18547]_  = \new_[18546]_  & \new_[18541]_ ;
  assign \new_[18551]_  = ~A266 & ~A236;
  assign \new_[18552]_  = ~A235 & \new_[18551]_ ;
  assign \new_[18556]_  = ~A300 & A298;
  assign \new_[18557]_  = ~A267 & \new_[18556]_ ;
  assign \new_[18558]_  = \new_[18557]_  & \new_[18552]_ ;
  assign \new_[18561]_  = A167 & A168;
  assign \new_[18565]_  = ~A233 & A200;
  assign \new_[18566]_  = A199 & \new_[18565]_ ;
  assign \new_[18567]_  = \new_[18566]_  & \new_[18561]_ ;
  assign \new_[18571]_  = ~A266 & ~A236;
  assign \new_[18572]_  = ~A235 & \new_[18571]_ ;
  assign \new_[18576]_  = A299 & A298;
  assign \new_[18577]_  = ~A267 & \new_[18576]_ ;
  assign \new_[18578]_  = \new_[18577]_  & \new_[18572]_ ;
  assign \new_[18581]_  = A167 & A168;
  assign \new_[18585]_  = ~A233 & A200;
  assign \new_[18586]_  = A199 & \new_[18585]_ ;
  assign \new_[18587]_  = \new_[18586]_  & \new_[18581]_ ;
  assign \new_[18591]_  = ~A266 & ~A236;
  assign \new_[18592]_  = ~A235 & \new_[18591]_ ;
  assign \new_[18596]_  = ~A299 & ~A298;
  assign \new_[18597]_  = ~A267 & \new_[18596]_ ;
  assign \new_[18598]_  = \new_[18597]_  & \new_[18592]_ ;
  assign \new_[18601]_  = A167 & A168;
  assign \new_[18605]_  = ~A233 & A200;
  assign \new_[18606]_  = A199 & \new_[18605]_ ;
  assign \new_[18607]_  = \new_[18606]_  & \new_[18601]_ ;
  assign \new_[18611]_  = ~A265 & ~A236;
  assign \new_[18612]_  = ~A235 & \new_[18611]_ ;
  assign \new_[18616]_  = ~A300 & A298;
  assign \new_[18617]_  = ~A266 & \new_[18616]_ ;
  assign \new_[18618]_  = \new_[18617]_  & \new_[18612]_ ;
  assign \new_[18621]_  = A167 & A168;
  assign \new_[18625]_  = ~A233 & A200;
  assign \new_[18626]_  = A199 & \new_[18625]_ ;
  assign \new_[18627]_  = \new_[18626]_  & \new_[18621]_ ;
  assign \new_[18631]_  = ~A265 & ~A236;
  assign \new_[18632]_  = ~A235 & \new_[18631]_ ;
  assign \new_[18636]_  = A299 & A298;
  assign \new_[18637]_  = ~A266 & \new_[18636]_ ;
  assign \new_[18638]_  = \new_[18637]_  & \new_[18632]_ ;
  assign \new_[18641]_  = A167 & A168;
  assign \new_[18645]_  = ~A233 & A200;
  assign \new_[18646]_  = A199 & \new_[18645]_ ;
  assign \new_[18647]_  = \new_[18646]_  & \new_[18641]_ ;
  assign \new_[18651]_  = ~A265 & ~A236;
  assign \new_[18652]_  = ~A235 & \new_[18651]_ ;
  assign \new_[18656]_  = ~A299 & ~A298;
  assign \new_[18657]_  = ~A266 & \new_[18656]_ ;
  assign \new_[18658]_  = \new_[18657]_  & \new_[18652]_ ;
  assign \new_[18661]_  = A167 & A168;
  assign \new_[18665]_  = ~A233 & A200;
  assign \new_[18666]_  = A199 & \new_[18665]_ ;
  assign \new_[18667]_  = \new_[18666]_  & \new_[18661]_ ;
  assign \new_[18671]_  = A266 & A265;
  assign \new_[18672]_  = ~A234 & \new_[18671]_ ;
  assign \new_[18676]_  = ~A302 & ~A301;
  assign \new_[18677]_  = A298 & \new_[18676]_ ;
  assign \new_[18678]_  = \new_[18677]_  & \new_[18672]_ ;
  assign \new_[18681]_  = A167 & A168;
  assign \new_[18685]_  = ~A233 & A200;
  assign \new_[18686]_  = A199 & \new_[18685]_ ;
  assign \new_[18687]_  = \new_[18686]_  & \new_[18681]_ ;
  assign \new_[18691]_  = ~A268 & ~A266;
  assign \new_[18692]_  = ~A234 & \new_[18691]_ ;
  assign \new_[18696]_  = ~A300 & A298;
  assign \new_[18697]_  = ~A269 & \new_[18696]_ ;
  assign \new_[18698]_  = \new_[18697]_  & \new_[18692]_ ;
  assign \new_[18701]_  = A167 & A168;
  assign \new_[18705]_  = ~A233 & A200;
  assign \new_[18706]_  = A199 & \new_[18705]_ ;
  assign \new_[18707]_  = \new_[18706]_  & \new_[18701]_ ;
  assign \new_[18711]_  = ~A268 & ~A266;
  assign \new_[18712]_  = ~A234 & \new_[18711]_ ;
  assign \new_[18716]_  = A299 & A298;
  assign \new_[18717]_  = ~A269 & \new_[18716]_ ;
  assign \new_[18718]_  = \new_[18717]_  & \new_[18712]_ ;
  assign \new_[18721]_  = A167 & A168;
  assign \new_[18725]_  = ~A233 & A200;
  assign \new_[18726]_  = A199 & \new_[18725]_ ;
  assign \new_[18727]_  = \new_[18726]_  & \new_[18721]_ ;
  assign \new_[18731]_  = ~A268 & ~A266;
  assign \new_[18732]_  = ~A234 & \new_[18731]_ ;
  assign \new_[18736]_  = ~A299 & ~A298;
  assign \new_[18737]_  = ~A269 & \new_[18736]_ ;
  assign \new_[18738]_  = \new_[18737]_  & \new_[18732]_ ;
  assign \new_[18741]_  = A167 & A168;
  assign \new_[18745]_  = ~A233 & A200;
  assign \new_[18746]_  = A199 & \new_[18745]_ ;
  assign \new_[18747]_  = \new_[18746]_  & \new_[18741]_ ;
  assign \new_[18751]_  = ~A267 & ~A266;
  assign \new_[18752]_  = ~A234 & \new_[18751]_ ;
  assign \new_[18756]_  = ~A302 & ~A301;
  assign \new_[18757]_  = A298 & \new_[18756]_ ;
  assign \new_[18758]_  = \new_[18757]_  & \new_[18752]_ ;
  assign \new_[18761]_  = A167 & A168;
  assign \new_[18765]_  = ~A233 & A200;
  assign \new_[18766]_  = A199 & \new_[18765]_ ;
  assign \new_[18767]_  = \new_[18766]_  & \new_[18761]_ ;
  assign \new_[18771]_  = ~A266 & ~A265;
  assign \new_[18772]_  = ~A234 & \new_[18771]_ ;
  assign \new_[18776]_  = ~A302 & ~A301;
  assign \new_[18777]_  = A298 & \new_[18776]_ ;
  assign \new_[18778]_  = \new_[18777]_  & \new_[18772]_ ;
  assign \new_[18781]_  = A167 & A168;
  assign \new_[18785]_  = ~A232 & A200;
  assign \new_[18786]_  = A199 & \new_[18785]_ ;
  assign \new_[18787]_  = \new_[18786]_  & \new_[18781]_ ;
  assign \new_[18791]_  = A266 & A265;
  assign \new_[18792]_  = ~A233 & \new_[18791]_ ;
  assign \new_[18796]_  = ~A302 & ~A301;
  assign \new_[18797]_  = A298 & \new_[18796]_ ;
  assign \new_[18798]_  = \new_[18797]_  & \new_[18792]_ ;
  assign \new_[18801]_  = A167 & A168;
  assign \new_[18805]_  = ~A232 & A200;
  assign \new_[18806]_  = A199 & \new_[18805]_ ;
  assign \new_[18807]_  = \new_[18806]_  & \new_[18801]_ ;
  assign \new_[18811]_  = ~A268 & ~A266;
  assign \new_[18812]_  = ~A233 & \new_[18811]_ ;
  assign \new_[18816]_  = ~A300 & A298;
  assign \new_[18817]_  = ~A269 & \new_[18816]_ ;
  assign \new_[18818]_  = \new_[18817]_  & \new_[18812]_ ;
  assign \new_[18821]_  = A167 & A168;
  assign \new_[18825]_  = ~A232 & A200;
  assign \new_[18826]_  = A199 & \new_[18825]_ ;
  assign \new_[18827]_  = \new_[18826]_  & \new_[18821]_ ;
  assign \new_[18831]_  = ~A268 & ~A266;
  assign \new_[18832]_  = ~A233 & \new_[18831]_ ;
  assign \new_[18836]_  = A299 & A298;
  assign \new_[18837]_  = ~A269 & \new_[18836]_ ;
  assign \new_[18838]_  = \new_[18837]_  & \new_[18832]_ ;
  assign \new_[18841]_  = A167 & A168;
  assign \new_[18845]_  = ~A232 & A200;
  assign \new_[18846]_  = A199 & \new_[18845]_ ;
  assign \new_[18847]_  = \new_[18846]_  & \new_[18841]_ ;
  assign \new_[18851]_  = ~A268 & ~A266;
  assign \new_[18852]_  = ~A233 & \new_[18851]_ ;
  assign \new_[18856]_  = ~A299 & ~A298;
  assign \new_[18857]_  = ~A269 & \new_[18856]_ ;
  assign \new_[18858]_  = \new_[18857]_  & \new_[18852]_ ;
  assign \new_[18861]_  = A167 & A168;
  assign \new_[18865]_  = ~A232 & A200;
  assign \new_[18866]_  = A199 & \new_[18865]_ ;
  assign \new_[18867]_  = \new_[18866]_  & \new_[18861]_ ;
  assign \new_[18871]_  = ~A267 & ~A266;
  assign \new_[18872]_  = ~A233 & \new_[18871]_ ;
  assign \new_[18876]_  = ~A302 & ~A301;
  assign \new_[18877]_  = A298 & \new_[18876]_ ;
  assign \new_[18878]_  = \new_[18877]_  & \new_[18872]_ ;
  assign \new_[18881]_  = A167 & A168;
  assign \new_[18885]_  = ~A232 & A200;
  assign \new_[18886]_  = A199 & \new_[18885]_ ;
  assign \new_[18887]_  = \new_[18886]_  & \new_[18881]_ ;
  assign \new_[18891]_  = ~A266 & ~A265;
  assign \new_[18892]_  = ~A233 & \new_[18891]_ ;
  assign \new_[18896]_  = ~A302 & ~A301;
  assign \new_[18897]_  = A298 & \new_[18896]_ ;
  assign \new_[18898]_  = \new_[18897]_  & \new_[18892]_ ;
  assign \new_[18901]_  = A167 & A168;
  assign \new_[18905]_  = ~A203 & ~A202;
  assign \new_[18906]_  = ~A200 & \new_[18905]_ ;
  assign \new_[18907]_  = \new_[18906]_  & \new_[18901]_ ;
  assign \new_[18911]_  = A265 & A233;
  assign \new_[18912]_  = A232 & \new_[18911]_ ;
  assign \new_[18916]_  = ~A300 & ~A299;
  assign \new_[18917]_  = ~A267 & \new_[18916]_ ;
  assign \new_[18918]_  = \new_[18917]_  & \new_[18912]_ ;
  assign \new_[18921]_  = A167 & A168;
  assign \new_[18925]_  = ~A203 & ~A202;
  assign \new_[18926]_  = ~A200 & \new_[18925]_ ;
  assign \new_[18927]_  = \new_[18926]_  & \new_[18921]_ ;
  assign \new_[18931]_  = A265 & A233;
  assign \new_[18932]_  = A232 & \new_[18931]_ ;
  assign \new_[18936]_  = A299 & A298;
  assign \new_[18937]_  = ~A267 & \new_[18936]_ ;
  assign \new_[18938]_  = \new_[18937]_  & \new_[18932]_ ;
  assign \new_[18941]_  = A167 & A168;
  assign \new_[18945]_  = ~A203 & ~A202;
  assign \new_[18946]_  = ~A200 & \new_[18945]_ ;
  assign \new_[18947]_  = \new_[18946]_  & \new_[18941]_ ;
  assign \new_[18951]_  = A265 & A233;
  assign \new_[18952]_  = A232 & \new_[18951]_ ;
  assign \new_[18956]_  = ~A299 & ~A298;
  assign \new_[18957]_  = ~A267 & \new_[18956]_ ;
  assign \new_[18958]_  = \new_[18957]_  & \new_[18952]_ ;
  assign \new_[18961]_  = A167 & A168;
  assign \new_[18965]_  = ~A203 & ~A202;
  assign \new_[18966]_  = ~A200 & \new_[18965]_ ;
  assign \new_[18967]_  = \new_[18966]_  & \new_[18961]_ ;
  assign \new_[18971]_  = A265 & A233;
  assign \new_[18972]_  = A232 & \new_[18971]_ ;
  assign \new_[18976]_  = ~A300 & ~A299;
  assign \new_[18977]_  = A266 & \new_[18976]_ ;
  assign \new_[18978]_  = \new_[18977]_  & \new_[18972]_ ;
  assign \new_[18981]_  = A167 & A168;
  assign \new_[18985]_  = ~A203 & ~A202;
  assign \new_[18986]_  = ~A200 & \new_[18985]_ ;
  assign \new_[18987]_  = \new_[18986]_  & \new_[18981]_ ;
  assign \new_[18991]_  = A265 & A233;
  assign \new_[18992]_  = A232 & \new_[18991]_ ;
  assign \new_[18996]_  = A299 & A298;
  assign \new_[18997]_  = A266 & \new_[18996]_ ;
  assign \new_[18998]_  = \new_[18997]_  & \new_[18992]_ ;
  assign \new_[19001]_  = A167 & A168;
  assign \new_[19005]_  = ~A203 & ~A202;
  assign \new_[19006]_  = ~A200 & \new_[19005]_ ;
  assign \new_[19007]_  = \new_[19006]_  & \new_[19001]_ ;
  assign \new_[19011]_  = A265 & A233;
  assign \new_[19012]_  = A232 & \new_[19011]_ ;
  assign \new_[19016]_  = ~A299 & ~A298;
  assign \new_[19017]_  = A266 & \new_[19016]_ ;
  assign \new_[19018]_  = \new_[19017]_  & \new_[19012]_ ;
  assign \new_[19021]_  = A167 & A168;
  assign \new_[19025]_  = ~A203 & ~A202;
  assign \new_[19026]_  = ~A200 & \new_[19025]_ ;
  assign \new_[19027]_  = \new_[19026]_  & \new_[19021]_ ;
  assign \new_[19031]_  = ~A265 & A233;
  assign \new_[19032]_  = A232 & \new_[19031]_ ;
  assign \new_[19036]_  = ~A300 & ~A299;
  assign \new_[19037]_  = ~A266 & \new_[19036]_ ;
  assign \new_[19038]_  = \new_[19037]_  & \new_[19032]_ ;
  assign \new_[19041]_  = A167 & A168;
  assign \new_[19045]_  = ~A203 & ~A202;
  assign \new_[19046]_  = ~A200 & \new_[19045]_ ;
  assign \new_[19047]_  = \new_[19046]_  & \new_[19041]_ ;
  assign \new_[19051]_  = ~A265 & A233;
  assign \new_[19052]_  = A232 & \new_[19051]_ ;
  assign \new_[19056]_  = A299 & A298;
  assign \new_[19057]_  = ~A266 & \new_[19056]_ ;
  assign \new_[19058]_  = \new_[19057]_  & \new_[19052]_ ;
  assign \new_[19061]_  = A167 & A168;
  assign \new_[19065]_  = ~A203 & ~A202;
  assign \new_[19066]_  = ~A200 & \new_[19065]_ ;
  assign \new_[19067]_  = \new_[19066]_  & \new_[19061]_ ;
  assign \new_[19071]_  = ~A265 & A233;
  assign \new_[19072]_  = A232 & \new_[19071]_ ;
  assign \new_[19076]_  = ~A299 & ~A298;
  assign \new_[19077]_  = ~A266 & \new_[19076]_ ;
  assign \new_[19078]_  = \new_[19077]_  & \new_[19072]_ ;
  assign \new_[19081]_  = A167 & A168;
  assign \new_[19085]_  = ~A203 & ~A202;
  assign \new_[19086]_  = ~A200 & \new_[19085]_ ;
  assign \new_[19087]_  = \new_[19086]_  & \new_[19081]_ ;
  assign \new_[19091]_  = A298 & A233;
  assign \new_[19092]_  = ~A232 & \new_[19091]_ ;
  assign \new_[19096]_  = A301 & A300;
  assign \new_[19097]_  = ~A299 & \new_[19096]_ ;
  assign \new_[19098]_  = \new_[19097]_  & \new_[19092]_ ;
  assign \new_[19101]_  = A167 & A168;
  assign \new_[19105]_  = ~A203 & ~A202;
  assign \new_[19106]_  = ~A200 & \new_[19105]_ ;
  assign \new_[19107]_  = \new_[19106]_  & \new_[19101]_ ;
  assign \new_[19111]_  = A298 & A233;
  assign \new_[19112]_  = ~A232 & \new_[19111]_ ;
  assign \new_[19116]_  = A302 & A300;
  assign \new_[19117]_  = ~A299 & \new_[19116]_ ;
  assign \new_[19118]_  = \new_[19117]_  & \new_[19112]_ ;
  assign \new_[19121]_  = A167 & A168;
  assign \new_[19125]_  = ~A203 & ~A202;
  assign \new_[19126]_  = ~A200 & \new_[19125]_ ;
  assign \new_[19127]_  = \new_[19126]_  & \new_[19121]_ ;
  assign \new_[19131]_  = A265 & A233;
  assign \new_[19132]_  = ~A232 & \new_[19131]_ ;
  assign \new_[19136]_  = A268 & A267;
  assign \new_[19137]_  = ~A266 & \new_[19136]_ ;
  assign \new_[19138]_  = \new_[19137]_  & \new_[19132]_ ;
  assign \new_[19141]_  = A167 & A168;
  assign \new_[19145]_  = ~A203 & ~A202;
  assign \new_[19146]_  = ~A200 & \new_[19145]_ ;
  assign \new_[19147]_  = \new_[19146]_  & \new_[19141]_ ;
  assign \new_[19151]_  = A265 & A233;
  assign \new_[19152]_  = ~A232 & \new_[19151]_ ;
  assign \new_[19156]_  = A269 & A267;
  assign \new_[19157]_  = ~A266 & \new_[19156]_ ;
  assign \new_[19158]_  = \new_[19157]_  & \new_[19152]_ ;
  assign \new_[19161]_  = A167 & A168;
  assign \new_[19165]_  = ~A203 & ~A202;
  assign \new_[19166]_  = ~A200 & \new_[19165]_ ;
  assign \new_[19167]_  = \new_[19166]_  & \new_[19161]_ ;
  assign \new_[19171]_  = A265 & ~A234;
  assign \new_[19172]_  = ~A233 & \new_[19171]_ ;
  assign \new_[19176]_  = ~A300 & A298;
  assign \new_[19177]_  = A266 & \new_[19176]_ ;
  assign \new_[19178]_  = \new_[19177]_  & \new_[19172]_ ;
  assign \new_[19181]_  = A167 & A168;
  assign \new_[19185]_  = ~A203 & ~A202;
  assign \new_[19186]_  = ~A200 & \new_[19185]_ ;
  assign \new_[19187]_  = \new_[19186]_  & \new_[19181]_ ;
  assign \new_[19191]_  = A265 & ~A234;
  assign \new_[19192]_  = ~A233 & \new_[19191]_ ;
  assign \new_[19196]_  = A299 & A298;
  assign \new_[19197]_  = A266 & \new_[19196]_ ;
  assign \new_[19198]_  = \new_[19197]_  & \new_[19192]_ ;
  assign \new_[19201]_  = A167 & A168;
  assign \new_[19205]_  = ~A203 & ~A202;
  assign \new_[19206]_  = ~A200 & \new_[19205]_ ;
  assign \new_[19207]_  = \new_[19206]_  & \new_[19201]_ ;
  assign \new_[19211]_  = A265 & ~A234;
  assign \new_[19212]_  = ~A233 & \new_[19211]_ ;
  assign \new_[19216]_  = ~A299 & ~A298;
  assign \new_[19217]_  = A266 & \new_[19216]_ ;
  assign \new_[19218]_  = \new_[19217]_  & \new_[19212]_ ;
  assign \new_[19221]_  = A167 & A168;
  assign \new_[19225]_  = ~A203 & ~A202;
  assign \new_[19226]_  = ~A200 & \new_[19225]_ ;
  assign \new_[19227]_  = \new_[19226]_  & \new_[19221]_ ;
  assign \new_[19231]_  = ~A266 & ~A234;
  assign \new_[19232]_  = ~A233 & \new_[19231]_ ;
  assign \new_[19236]_  = ~A300 & A298;
  assign \new_[19237]_  = ~A267 & \new_[19236]_ ;
  assign \new_[19238]_  = \new_[19237]_  & \new_[19232]_ ;
  assign \new_[19241]_  = A167 & A168;
  assign \new_[19245]_  = ~A203 & ~A202;
  assign \new_[19246]_  = ~A200 & \new_[19245]_ ;
  assign \new_[19247]_  = \new_[19246]_  & \new_[19241]_ ;
  assign \new_[19251]_  = ~A266 & ~A234;
  assign \new_[19252]_  = ~A233 & \new_[19251]_ ;
  assign \new_[19256]_  = A299 & A298;
  assign \new_[19257]_  = ~A267 & \new_[19256]_ ;
  assign \new_[19258]_  = \new_[19257]_  & \new_[19252]_ ;
  assign \new_[19261]_  = A167 & A168;
  assign \new_[19265]_  = ~A203 & ~A202;
  assign \new_[19266]_  = ~A200 & \new_[19265]_ ;
  assign \new_[19267]_  = \new_[19266]_  & \new_[19261]_ ;
  assign \new_[19271]_  = ~A266 & ~A234;
  assign \new_[19272]_  = ~A233 & \new_[19271]_ ;
  assign \new_[19276]_  = ~A299 & ~A298;
  assign \new_[19277]_  = ~A267 & \new_[19276]_ ;
  assign \new_[19278]_  = \new_[19277]_  & \new_[19272]_ ;
  assign \new_[19281]_  = A167 & A168;
  assign \new_[19285]_  = ~A203 & ~A202;
  assign \new_[19286]_  = ~A200 & \new_[19285]_ ;
  assign \new_[19287]_  = \new_[19286]_  & \new_[19281]_ ;
  assign \new_[19291]_  = ~A265 & ~A234;
  assign \new_[19292]_  = ~A233 & \new_[19291]_ ;
  assign \new_[19296]_  = ~A300 & A298;
  assign \new_[19297]_  = ~A266 & \new_[19296]_ ;
  assign \new_[19298]_  = \new_[19297]_  & \new_[19292]_ ;
  assign \new_[19301]_  = A167 & A168;
  assign \new_[19305]_  = ~A203 & ~A202;
  assign \new_[19306]_  = ~A200 & \new_[19305]_ ;
  assign \new_[19307]_  = \new_[19306]_  & \new_[19301]_ ;
  assign \new_[19311]_  = ~A265 & ~A234;
  assign \new_[19312]_  = ~A233 & \new_[19311]_ ;
  assign \new_[19316]_  = A299 & A298;
  assign \new_[19317]_  = ~A266 & \new_[19316]_ ;
  assign \new_[19318]_  = \new_[19317]_  & \new_[19312]_ ;
  assign \new_[19321]_  = A167 & A168;
  assign \new_[19325]_  = ~A203 & ~A202;
  assign \new_[19326]_  = ~A200 & \new_[19325]_ ;
  assign \new_[19327]_  = \new_[19326]_  & \new_[19321]_ ;
  assign \new_[19331]_  = ~A265 & ~A234;
  assign \new_[19332]_  = ~A233 & \new_[19331]_ ;
  assign \new_[19336]_  = ~A299 & ~A298;
  assign \new_[19337]_  = ~A266 & \new_[19336]_ ;
  assign \new_[19338]_  = \new_[19337]_  & \new_[19332]_ ;
  assign \new_[19341]_  = A167 & A168;
  assign \new_[19345]_  = ~A203 & ~A202;
  assign \new_[19346]_  = ~A200 & \new_[19345]_ ;
  assign \new_[19347]_  = \new_[19346]_  & \new_[19341]_ ;
  assign \new_[19351]_  = A234 & ~A233;
  assign \new_[19352]_  = A232 & \new_[19351]_ ;
  assign \new_[19356]_  = A299 & ~A298;
  assign \new_[19357]_  = A235 & \new_[19356]_ ;
  assign \new_[19358]_  = \new_[19357]_  & \new_[19352]_ ;
  assign \new_[19361]_  = A167 & A168;
  assign \new_[19365]_  = ~A203 & ~A202;
  assign \new_[19366]_  = ~A200 & \new_[19365]_ ;
  assign \new_[19367]_  = \new_[19366]_  & \new_[19361]_ ;
  assign \new_[19371]_  = A234 & ~A233;
  assign \new_[19372]_  = A232 & \new_[19371]_ ;
  assign \new_[19376]_  = A266 & ~A265;
  assign \new_[19377]_  = A235 & \new_[19376]_ ;
  assign \new_[19378]_  = \new_[19377]_  & \new_[19372]_ ;
  assign \new_[19381]_  = A167 & A168;
  assign \new_[19385]_  = ~A203 & ~A202;
  assign \new_[19386]_  = ~A200 & \new_[19385]_ ;
  assign \new_[19387]_  = \new_[19386]_  & \new_[19381]_ ;
  assign \new_[19391]_  = A234 & ~A233;
  assign \new_[19392]_  = A232 & \new_[19391]_ ;
  assign \new_[19396]_  = A299 & ~A298;
  assign \new_[19397]_  = A236 & \new_[19396]_ ;
  assign \new_[19398]_  = \new_[19397]_  & \new_[19392]_ ;
  assign \new_[19401]_  = A167 & A168;
  assign \new_[19405]_  = ~A203 & ~A202;
  assign \new_[19406]_  = ~A200 & \new_[19405]_ ;
  assign \new_[19407]_  = \new_[19406]_  & \new_[19401]_ ;
  assign \new_[19411]_  = A234 & ~A233;
  assign \new_[19412]_  = A232 & \new_[19411]_ ;
  assign \new_[19416]_  = A266 & ~A265;
  assign \new_[19417]_  = A236 & \new_[19416]_ ;
  assign \new_[19418]_  = \new_[19417]_  & \new_[19412]_ ;
  assign \new_[19421]_  = A167 & A168;
  assign \new_[19425]_  = ~A203 & ~A202;
  assign \new_[19426]_  = ~A200 & \new_[19425]_ ;
  assign \new_[19427]_  = \new_[19426]_  & \new_[19421]_ ;
  assign \new_[19431]_  = A265 & ~A233;
  assign \new_[19432]_  = ~A232 & \new_[19431]_ ;
  assign \new_[19436]_  = ~A300 & A298;
  assign \new_[19437]_  = A266 & \new_[19436]_ ;
  assign \new_[19438]_  = \new_[19437]_  & \new_[19432]_ ;
  assign \new_[19441]_  = A167 & A168;
  assign \new_[19445]_  = ~A203 & ~A202;
  assign \new_[19446]_  = ~A200 & \new_[19445]_ ;
  assign \new_[19447]_  = \new_[19446]_  & \new_[19441]_ ;
  assign \new_[19451]_  = A265 & ~A233;
  assign \new_[19452]_  = ~A232 & \new_[19451]_ ;
  assign \new_[19456]_  = A299 & A298;
  assign \new_[19457]_  = A266 & \new_[19456]_ ;
  assign \new_[19458]_  = \new_[19457]_  & \new_[19452]_ ;
  assign \new_[19461]_  = A167 & A168;
  assign \new_[19465]_  = ~A203 & ~A202;
  assign \new_[19466]_  = ~A200 & \new_[19465]_ ;
  assign \new_[19467]_  = \new_[19466]_  & \new_[19461]_ ;
  assign \new_[19471]_  = A265 & ~A233;
  assign \new_[19472]_  = ~A232 & \new_[19471]_ ;
  assign \new_[19476]_  = ~A299 & ~A298;
  assign \new_[19477]_  = A266 & \new_[19476]_ ;
  assign \new_[19478]_  = \new_[19477]_  & \new_[19472]_ ;
  assign \new_[19481]_  = A167 & A168;
  assign \new_[19485]_  = ~A203 & ~A202;
  assign \new_[19486]_  = ~A200 & \new_[19485]_ ;
  assign \new_[19487]_  = \new_[19486]_  & \new_[19481]_ ;
  assign \new_[19491]_  = ~A266 & ~A233;
  assign \new_[19492]_  = ~A232 & \new_[19491]_ ;
  assign \new_[19496]_  = ~A300 & A298;
  assign \new_[19497]_  = ~A267 & \new_[19496]_ ;
  assign \new_[19498]_  = \new_[19497]_  & \new_[19492]_ ;
  assign \new_[19501]_  = A167 & A168;
  assign \new_[19505]_  = ~A203 & ~A202;
  assign \new_[19506]_  = ~A200 & \new_[19505]_ ;
  assign \new_[19507]_  = \new_[19506]_  & \new_[19501]_ ;
  assign \new_[19511]_  = ~A266 & ~A233;
  assign \new_[19512]_  = ~A232 & \new_[19511]_ ;
  assign \new_[19516]_  = A299 & A298;
  assign \new_[19517]_  = ~A267 & \new_[19516]_ ;
  assign \new_[19518]_  = \new_[19517]_  & \new_[19512]_ ;
  assign \new_[19521]_  = A167 & A168;
  assign \new_[19525]_  = ~A203 & ~A202;
  assign \new_[19526]_  = ~A200 & \new_[19525]_ ;
  assign \new_[19527]_  = \new_[19526]_  & \new_[19521]_ ;
  assign \new_[19531]_  = ~A266 & ~A233;
  assign \new_[19532]_  = ~A232 & \new_[19531]_ ;
  assign \new_[19536]_  = ~A299 & ~A298;
  assign \new_[19537]_  = ~A267 & \new_[19536]_ ;
  assign \new_[19538]_  = \new_[19537]_  & \new_[19532]_ ;
  assign \new_[19541]_  = A167 & A168;
  assign \new_[19545]_  = ~A203 & ~A202;
  assign \new_[19546]_  = ~A200 & \new_[19545]_ ;
  assign \new_[19547]_  = \new_[19546]_  & \new_[19541]_ ;
  assign \new_[19551]_  = ~A265 & ~A233;
  assign \new_[19552]_  = ~A232 & \new_[19551]_ ;
  assign \new_[19556]_  = ~A300 & A298;
  assign \new_[19557]_  = ~A266 & \new_[19556]_ ;
  assign \new_[19558]_  = \new_[19557]_  & \new_[19552]_ ;
  assign \new_[19561]_  = A167 & A168;
  assign \new_[19565]_  = ~A203 & ~A202;
  assign \new_[19566]_  = ~A200 & \new_[19565]_ ;
  assign \new_[19567]_  = \new_[19566]_  & \new_[19561]_ ;
  assign \new_[19571]_  = ~A265 & ~A233;
  assign \new_[19572]_  = ~A232 & \new_[19571]_ ;
  assign \new_[19576]_  = A299 & A298;
  assign \new_[19577]_  = ~A266 & \new_[19576]_ ;
  assign \new_[19578]_  = \new_[19577]_  & \new_[19572]_ ;
  assign \new_[19581]_  = A167 & A168;
  assign \new_[19585]_  = ~A203 & ~A202;
  assign \new_[19586]_  = ~A200 & \new_[19585]_ ;
  assign \new_[19587]_  = \new_[19586]_  & \new_[19581]_ ;
  assign \new_[19591]_  = ~A265 & ~A233;
  assign \new_[19592]_  = ~A232 & \new_[19591]_ ;
  assign \new_[19596]_  = ~A299 & ~A298;
  assign \new_[19597]_  = ~A266 & \new_[19596]_ ;
  assign \new_[19598]_  = \new_[19597]_  & \new_[19592]_ ;
  assign \new_[19601]_  = A167 & A168;
  assign \new_[19605]_  = A232 & ~A201;
  assign \new_[19606]_  = ~A200 & \new_[19605]_ ;
  assign \new_[19607]_  = \new_[19606]_  & \new_[19601]_ ;
  assign \new_[19611]_  = ~A268 & A265;
  assign \new_[19612]_  = A233 & \new_[19611]_ ;
  assign \new_[19616]_  = ~A300 & ~A299;
  assign \new_[19617]_  = ~A269 & \new_[19616]_ ;
  assign \new_[19618]_  = \new_[19617]_  & \new_[19612]_ ;
  assign \new_[19621]_  = A167 & A168;
  assign \new_[19625]_  = A232 & ~A201;
  assign \new_[19626]_  = ~A200 & \new_[19625]_ ;
  assign \new_[19627]_  = \new_[19626]_  & \new_[19621]_ ;
  assign \new_[19631]_  = ~A268 & A265;
  assign \new_[19632]_  = A233 & \new_[19631]_ ;
  assign \new_[19636]_  = A299 & A298;
  assign \new_[19637]_  = ~A269 & \new_[19636]_ ;
  assign \new_[19638]_  = \new_[19637]_  & \new_[19632]_ ;
  assign \new_[19641]_  = A167 & A168;
  assign \new_[19645]_  = A232 & ~A201;
  assign \new_[19646]_  = ~A200 & \new_[19645]_ ;
  assign \new_[19647]_  = \new_[19646]_  & \new_[19641]_ ;
  assign \new_[19651]_  = ~A268 & A265;
  assign \new_[19652]_  = A233 & \new_[19651]_ ;
  assign \new_[19656]_  = ~A299 & ~A298;
  assign \new_[19657]_  = ~A269 & \new_[19656]_ ;
  assign \new_[19658]_  = \new_[19657]_  & \new_[19652]_ ;
  assign \new_[19661]_  = A167 & A168;
  assign \new_[19665]_  = A232 & ~A201;
  assign \new_[19666]_  = ~A200 & \new_[19665]_ ;
  assign \new_[19667]_  = \new_[19666]_  & \new_[19661]_ ;
  assign \new_[19671]_  = ~A267 & A265;
  assign \new_[19672]_  = A233 & \new_[19671]_ ;
  assign \new_[19676]_  = ~A302 & ~A301;
  assign \new_[19677]_  = ~A299 & \new_[19676]_ ;
  assign \new_[19678]_  = \new_[19677]_  & \new_[19672]_ ;
  assign \new_[19681]_  = A167 & A168;
  assign \new_[19685]_  = A232 & ~A201;
  assign \new_[19686]_  = ~A200 & \new_[19685]_ ;
  assign \new_[19687]_  = \new_[19686]_  & \new_[19681]_ ;
  assign \new_[19691]_  = A266 & A265;
  assign \new_[19692]_  = A233 & \new_[19691]_ ;
  assign \new_[19696]_  = ~A302 & ~A301;
  assign \new_[19697]_  = ~A299 & \new_[19696]_ ;
  assign \new_[19698]_  = \new_[19697]_  & \new_[19692]_ ;
  assign \new_[19701]_  = A167 & A168;
  assign \new_[19705]_  = A232 & ~A201;
  assign \new_[19706]_  = ~A200 & \new_[19705]_ ;
  assign \new_[19707]_  = \new_[19706]_  & \new_[19701]_ ;
  assign \new_[19711]_  = ~A266 & ~A265;
  assign \new_[19712]_  = A233 & \new_[19711]_ ;
  assign \new_[19716]_  = ~A302 & ~A301;
  assign \new_[19717]_  = ~A299 & \new_[19716]_ ;
  assign \new_[19718]_  = \new_[19717]_  & \new_[19712]_ ;
  assign \new_[19721]_  = A167 & A168;
  assign \new_[19725]_  = ~A233 & ~A201;
  assign \new_[19726]_  = ~A200 & \new_[19725]_ ;
  assign \new_[19727]_  = \new_[19726]_  & \new_[19721]_ ;
  assign \new_[19731]_  = A265 & ~A236;
  assign \new_[19732]_  = ~A235 & \new_[19731]_ ;
  assign \new_[19736]_  = ~A300 & A298;
  assign \new_[19737]_  = A266 & \new_[19736]_ ;
  assign \new_[19738]_  = \new_[19737]_  & \new_[19732]_ ;
  assign \new_[19741]_  = A167 & A168;
  assign \new_[19745]_  = ~A233 & ~A201;
  assign \new_[19746]_  = ~A200 & \new_[19745]_ ;
  assign \new_[19747]_  = \new_[19746]_  & \new_[19741]_ ;
  assign \new_[19751]_  = A265 & ~A236;
  assign \new_[19752]_  = ~A235 & \new_[19751]_ ;
  assign \new_[19756]_  = A299 & A298;
  assign \new_[19757]_  = A266 & \new_[19756]_ ;
  assign \new_[19758]_  = \new_[19757]_  & \new_[19752]_ ;
  assign \new_[19761]_  = A167 & A168;
  assign \new_[19765]_  = ~A233 & ~A201;
  assign \new_[19766]_  = ~A200 & \new_[19765]_ ;
  assign \new_[19767]_  = \new_[19766]_  & \new_[19761]_ ;
  assign \new_[19771]_  = A265 & ~A236;
  assign \new_[19772]_  = ~A235 & \new_[19771]_ ;
  assign \new_[19776]_  = ~A299 & ~A298;
  assign \new_[19777]_  = A266 & \new_[19776]_ ;
  assign \new_[19778]_  = \new_[19777]_  & \new_[19772]_ ;
  assign \new_[19781]_  = A167 & A168;
  assign \new_[19785]_  = ~A233 & ~A201;
  assign \new_[19786]_  = ~A200 & \new_[19785]_ ;
  assign \new_[19787]_  = \new_[19786]_  & \new_[19781]_ ;
  assign \new_[19791]_  = ~A266 & ~A236;
  assign \new_[19792]_  = ~A235 & \new_[19791]_ ;
  assign \new_[19796]_  = ~A300 & A298;
  assign \new_[19797]_  = ~A267 & \new_[19796]_ ;
  assign \new_[19798]_  = \new_[19797]_  & \new_[19792]_ ;
  assign \new_[19801]_  = A167 & A168;
  assign \new_[19805]_  = ~A233 & ~A201;
  assign \new_[19806]_  = ~A200 & \new_[19805]_ ;
  assign \new_[19807]_  = \new_[19806]_  & \new_[19801]_ ;
  assign \new_[19811]_  = ~A266 & ~A236;
  assign \new_[19812]_  = ~A235 & \new_[19811]_ ;
  assign \new_[19816]_  = A299 & A298;
  assign \new_[19817]_  = ~A267 & \new_[19816]_ ;
  assign \new_[19818]_  = \new_[19817]_  & \new_[19812]_ ;
  assign \new_[19821]_  = A167 & A168;
  assign \new_[19825]_  = ~A233 & ~A201;
  assign \new_[19826]_  = ~A200 & \new_[19825]_ ;
  assign \new_[19827]_  = \new_[19826]_  & \new_[19821]_ ;
  assign \new_[19831]_  = ~A266 & ~A236;
  assign \new_[19832]_  = ~A235 & \new_[19831]_ ;
  assign \new_[19836]_  = ~A299 & ~A298;
  assign \new_[19837]_  = ~A267 & \new_[19836]_ ;
  assign \new_[19838]_  = \new_[19837]_  & \new_[19832]_ ;
  assign \new_[19841]_  = A167 & A168;
  assign \new_[19845]_  = ~A233 & ~A201;
  assign \new_[19846]_  = ~A200 & \new_[19845]_ ;
  assign \new_[19847]_  = \new_[19846]_  & \new_[19841]_ ;
  assign \new_[19851]_  = ~A265 & ~A236;
  assign \new_[19852]_  = ~A235 & \new_[19851]_ ;
  assign \new_[19856]_  = ~A300 & A298;
  assign \new_[19857]_  = ~A266 & \new_[19856]_ ;
  assign \new_[19858]_  = \new_[19857]_  & \new_[19852]_ ;
  assign \new_[19861]_  = A167 & A168;
  assign \new_[19865]_  = ~A233 & ~A201;
  assign \new_[19866]_  = ~A200 & \new_[19865]_ ;
  assign \new_[19867]_  = \new_[19866]_  & \new_[19861]_ ;
  assign \new_[19871]_  = ~A265 & ~A236;
  assign \new_[19872]_  = ~A235 & \new_[19871]_ ;
  assign \new_[19876]_  = A299 & A298;
  assign \new_[19877]_  = ~A266 & \new_[19876]_ ;
  assign \new_[19878]_  = \new_[19877]_  & \new_[19872]_ ;
  assign \new_[19881]_  = A167 & A168;
  assign \new_[19885]_  = ~A233 & ~A201;
  assign \new_[19886]_  = ~A200 & \new_[19885]_ ;
  assign \new_[19887]_  = \new_[19886]_  & \new_[19881]_ ;
  assign \new_[19891]_  = ~A265 & ~A236;
  assign \new_[19892]_  = ~A235 & \new_[19891]_ ;
  assign \new_[19896]_  = ~A299 & ~A298;
  assign \new_[19897]_  = ~A266 & \new_[19896]_ ;
  assign \new_[19898]_  = \new_[19897]_  & \new_[19892]_ ;
  assign \new_[19901]_  = A167 & A168;
  assign \new_[19905]_  = ~A233 & ~A201;
  assign \new_[19906]_  = ~A200 & \new_[19905]_ ;
  assign \new_[19907]_  = \new_[19906]_  & \new_[19901]_ ;
  assign \new_[19911]_  = A266 & A265;
  assign \new_[19912]_  = ~A234 & \new_[19911]_ ;
  assign \new_[19916]_  = ~A302 & ~A301;
  assign \new_[19917]_  = A298 & \new_[19916]_ ;
  assign \new_[19918]_  = \new_[19917]_  & \new_[19912]_ ;
  assign \new_[19921]_  = A167 & A168;
  assign \new_[19925]_  = ~A233 & ~A201;
  assign \new_[19926]_  = ~A200 & \new_[19925]_ ;
  assign \new_[19927]_  = \new_[19926]_  & \new_[19921]_ ;
  assign \new_[19931]_  = ~A268 & ~A266;
  assign \new_[19932]_  = ~A234 & \new_[19931]_ ;
  assign \new_[19936]_  = ~A300 & A298;
  assign \new_[19937]_  = ~A269 & \new_[19936]_ ;
  assign \new_[19938]_  = \new_[19937]_  & \new_[19932]_ ;
  assign \new_[19941]_  = A167 & A168;
  assign \new_[19945]_  = ~A233 & ~A201;
  assign \new_[19946]_  = ~A200 & \new_[19945]_ ;
  assign \new_[19947]_  = \new_[19946]_  & \new_[19941]_ ;
  assign \new_[19951]_  = ~A268 & ~A266;
  assign \new_[19952]_  = ~A234 & \new_[19951]_ ;
  assign \new_[19956]_  = A299 & A298;
  assign \new_[19957]_  = ~A269 & \new_[19956]_ ;
  assign \new_[19958]_  = \new_[19957]_  & \new_[19952]_ ;
  assign \new_[19961]_  = A167 & A168;
  assign \new_[19965]_  = ~A233 & ~A201;
  assign \new_[19966]_  = ~A200 & \new_[19965]_ ;
  assign \new_[19967]_  = \new_[19966]_  & \new_[19961]_ ;
  assign \new_[19971]_  = ~A268 & ~A266;
  assign \new_[19972]_  = ~A234 & \new_[19971]_ ;
  assign \new_[19976]_  = ~A299 & ~A298;
  assign \new_[19977]_  = ~A269 & \new_[19976]_ ;
  assign \new_[19978]_  = \new_[19977]_  & \new_[19972]_ ;
  assign \new_[19981]_  = A167 & A168;
  assign \new_[19985]_  = ~A233 & ~A201;
  assign \new_[19986]_  = ~A200 & \new_[19985]_ ;
  assign \new_[19987]_  = \new_[19986]_  & \new_[19981]_ ;
  assign \new_[19991]_  = ~A267 & ~A266;
  assign \new_[19992]_  = ~A234 & \new_[19991]_ ;
  assign \new_[19996]_  = ~A302 & ~A301;
  assign \new_[19997]_  = A298 & \new_[19996]_ ;
  assign \new_[19998]_  = \new_[19997]_  & \new_[19992]_ ;
  assign \new_[20001]_  = A167 & A168;
  assign \new_[20005]_  = ~A233 & ~A201;
  assign \new_[20006]_  = ~A200 & \new_[20005]_ ;
  assign \new_[20007]_  = \new_[20006]_  & \new_[20001]_ ;
  assign \new_[20011]_  = ~A266 & ~A265;
  assign \new_[20012]_  = ~A234 & \new_[20011]_ ;
  assign \new_[20016]_  = ~A302 & ~A301;
  assign \new_[20017]_  = A298 & \new_[20016]_ ;
  assign \new_[20018]_  = \new_[20017]_  & \new_[20012]_ ;
  assign \new_[20021]_  = A167 & A168;
  assign \new_[20025]_  = ~A232 & ~A201;
  assign \new_[20026]_  = ~A200 & \new_[20025]_ ;
  assign \new_[20027]_  = \new_[20026]_  & \new_[20021]_ ;
  assign \new_[20031]_  = A266 & A265;
  assign \new_[20032]_  = ~A233 & \new_[20031]_ ;
  assign \new_[20036]_  = ~A302 & ~A301;
  assign \new_[20037]_  = A298 & \new_[20036]_ ;
  assign \new_[20038]_  = \new_[20037]_  & \new_[20032]_ ;
  assign \new_[20041]_  = A167 & A168;
  assign \new_[20045]_  = ~A232 & ~A201;
  assign \new_[20046]_  = ~A200 & \new_[20045]_ ;
  assign \new_[20047]_  = \new_[20046]_  & \new_[20041]_ ;
  assign \new_[20051]_  = ~A268 & ~A266;
  assign \new_[20052]_  = ~A233 & \new_[20051]_ ;
  assign \new_[20056]_  = ~A300 & A298;
  assign \new_[20057]_  = ~A269 & \new_[20056]_ ;
  assign \new_[20058]_  = \new_[20057]_  & \new_[20052]_ ;
  assign \new_[20061]_  = A167 & A168;
  assign \new_[20065]_  = ~A232 & ~A201;
  assign \new_[20066]_  = ~A200 & \new_[20065]_ ;
  assign \new_[20067]_  = \new_[20066]_  & \new_[20061]_ ;
  assign \new_[20071]_  = ~A268 & ~A266;
  assign \new_[20072]_  = ~A233 & \new_[20071]_ ;
  assign \new_[20076]_  = A299 & A298;
  assign \new_[20077]_  = ~A269 & \new_[20076]_ ;
  assign \new_[20078]_  = \new_[20077]_  & \new_[20072]_ ;
  assign \new_[20081]_  = A167 & A168;
  assign \new_[20085]_  = ~A232 & ~A201;
  assign \new_[20086]_  = ~A200 & \new_[20085]_ ;
  assign \new_[20087]_  = \new_[20086]_  & \new_[20081]_ ;
  assign \new_[20091]_  = ~A268 & ~A266;
  assign \new_[20092]_  = ~A233 & \new_[20091]_ ;
  assign \new_[20096]_  = ~A299 & ~A298;
  assign \new_[20097]_  = ~A269 & \new_[20096]_ ;
  assign \new_[20098]_  = \new_[20097]_  & \new_[20092]_ ;
  assign \new_[20101]_  = A167 & A168;
  assign \new_[20105]_  = ~A232 & ~A201;
  assign \new_[20106]_  = ~A200 & \new_[20105]_ ;
  assign \new_[20107]_  = \new_[20106]_  & \new_[20101]_ ;
  assign \new_[20111]_  = ~A267 & ~A266;
  assign \new_[20112]_  = ~A233 & \new_[20111]_ ;
  assign \new_[20116]_  = ~A302 & ~A301;
  assign \new_[20117]_  = A298 & \new_[20116]_ ;
  assign \new_[20118]_  = \new_[20117]_  & \new_[20112]_ ;
  assign \new_[20121]_  = A167 & A168;
  assign \new_[20125]_  = ~A232 & ~A201;
  assign \new_[20126]_  = ~A200 & \new_[20125]_ ;
  assign \new_[20127]_  = \new_[20126]_  & \new_[20121]_ ;
  assign \new_[20131]_  = ~A266 & ~A265;
  assign \new_[20132]_  = ~A233 & \new_[20131]_ ;
  assign \new_[20136]_  = ~A302 & ~A301;
  assign \new_[20137]_  = A298 & \new_[20136]_ ;
  assign \new_[20138]_  = \new_[20137]_  & \new_[20132]_ ;
  assign \new_[20141]_  = A167 & A168;
  assign \new_[20145]_  = A232 & ~A200;
  assign \new_[20146]_  = ~A199 & \new_[20145]_ ;
  assign \new_[20147]_  = \new_[20146]_  & \new_[20141]_ ;
  assign \new_[20151]_  = ~A268 & A265;
  assign \new_[20152]_  = A233 & \new_[20151]_ ;
  assign \new_[20156]_  = ~A300 & ~A299;
  assign \new_[20157]_  = ~A269 & \new_[20156]_ ;
  assign \new_[20158]_  = \new_[20157]_  & \new_[20152]_ ;
  assign \new_[20161]_  = A167 & A168;
  assign \new_[20165]_  = A232 & ~A200;
  assign \new_[20166]_  = ~A199 & \new_[20165]_ ;
  assign \new_[20167]_  = \new_[20166]_  & \new_[20161]_ ;
  assign \new_[20171]_  = ~A268 & A265;
  assign \new_[20172]_  = A233 & \new_[20171]_ ;
  assign \new_[20176]_  = A299 & A298;
  assign \new_[20177]_  = ~A269 & \new_[20176]_ ;
  assign \new_[20178]_  = \new_[20177]_  & \new_[20172]_ ;
  assign \new_[20181]_  = A167 & A168;
  assign \new_[20185]_  = A232 & ~A200;
  assign \new_[20186]_  = ~A199 & \new_[20185]_ ;
  assign \new_[20187]_  = \new_[20186]_  & \new_[20181]_ ;
  assign \new_[20191]_  = ~A268 & A265;
  assign \new_[20192]_  = A233 & \new_[20191]_ ;
  assign \new_[20196]_  = ~A299 & ~A298;
  assign \new_[20197]_  = ~A269 & \new_[20196]_ ;
  assign \new_[20198]_  = \new_[20197]_  & \new_[20192]_ ;
  assign \new_[20201]_  = A167 & A168;
  assign \new_[20205]_  = A232 & ~A200;
  assign \new_[20206]_  = ~A199 & \new_[20205]_ ;
  assign \new_[20207]_  = \new_[20206]_  & \new_[20201]_ ;
  assign \new_[20211]_  = ~A267 & A265;
  assign \new_[20212]_  = A233 & \new_[20211]_ ;
  assign \new_[20216]_  = ~A302 & ~A301;
  assign \new_[20217]_  = ~A299 & \new_[20216]_ ;
  assign \new_[20218]_  = \new_[20217]_  & \new_[20212]_ ;
  assign \new_[20221]_  = A167 & A168;
  assign \new_[20225]_  = A232 & ~A200;
  assign \new_[20226]_  = ~A199 & \new_[20225]_ ;
  assign \new_[20227]_  = \new_[20226]_  & \new_[20221]_ ;
  assign \new_[20231]_  = A266 & A265;
  assign \new_[20232]_  = A233 & \new_[20231]_ ;
  assign \new_[20236]_  = ~A302 & ~A301;
  assign \new_[20237]_  = ~A299 & \new_[20236]_ ;
  assign \new_[20238]_  = \new_[20237]_  & \new_[20232]_ ;
  assign \new_[20241]_  = A167 & A168;
  assign \new_[20245]_  = A232 & ~A200;
  assign \new_[20246]_  = ~A199 & \new_[20245]_ ;
  assign \new_[20247]_  = \new_[20246]_  & \new_[20241]_ ;
  assign \new_[20251]_  = ~A266 & ~A265;
  assign \new_[20252]_  = A233 & \new_[20251]_ ;
  assign \new_[20256]_  = ~A302 & ~A301;
  assign \new_[20257]_  = ~A299 & \new_[20256]_ ;
  assign \new_[20258]_  = \new_[20257]_  & \new_[20252]_ ;
  assign \new_[20261]_  = A167 & A168;
  assign \new_[20265]_  = ~A233 & ~A200;
  assign \new_[20266]_  = ~A199 & \new_[20265]_ ;
  assign \new_[20267]_  = \new_[20266]_  & \new_[20261]_ ;
  assign \new_[20271]_  = A265 & ~A236;
  assign \new_[20272]_  = ~A235 & \new_[20271]_ ;
  assign \new_[20276]_  = ~A300 & A298;
  assign \new_[20277]_  = A266 & \new_[20276]_ ;
  assign \new_[20278]_  = \new_[20277]_  & \new_[20272]_ ;
  assign \new_[20281]_  = A167 & A168;
  assign \new_[20285]_  = ~A233 & ~A200;
  assign \new_[20286]_  = ~A199 & \new_[20285]_ ;
  assign \new_[20287]_  = \new_[20286]_  & \new_[20281]_ ;
  assign \new_[20291]_  = A265 & ~A236;
  assign \new_[20292]_  = ~A235 & \new_[20291]_ ;
  assign \new_[20296]_  = A299 & A298;
  assign \new_[20297]_  = A266 & \new_[20296]_ ;
  assign \new_[20298]_  = \new_[20297]_  & \new_[20292]_ ;
  assign \new_[20301]_  = A167 & A168;
  assign \new_[20305]_  = ~A233 & ~A200;
  assign \new_[20306]_  = ~A199 & \new_[20305]_ ;
  assign \new_[20307]_  = \new_[20306]_  & \new_[20301]_ ;
  assign \new_[20311]_  = A265 & ~A236;
  assign \new_[20312]_  = ~A235 & \new_[20311]_ ;
  assign \new_[20316]_  = ~A299 & ~A298;
  assign \new_[20317]_  = A266 & \new_[20316]_ ;
  assign \new_[20318]_  = \new_[20317]_  & \new_[20312]_ ;
  assign \new_[20321]_  = A167 & A168;
  assign \new_[20325]_  = ~A233 & ~A200;
  assign \new_[20326]_  = ~A199 & \new_[20325]_ ;
  assign \new_[20327]_  = \new_[20326]_  & \new_[20321]_ ;
  assign \new_[20331]_  = ~A266 & ~A236;
  assign \new_[20332]_  = ~A235 & \new_[20331]_ ;
  assign \new_[20336]_  = ~A300 & A298;
  assign \new_[20337]_  = ~A267 & \new_[20336]_ ;
  assign \new_[20338]_  = \new_[20337]_  & \new_[20332]_ ;
  assign \new_[20341]_  = A167 & A168;
  assign \new_[20345]_  = ~A233 & ~A200;
  assign \new_[20346]_  = ~A199 & \new_[20345]_ ;
  assign \new_[20347]_  = \new_[20346]_  & \new_[20341]_ ;
  assign \new_[20351]_  = ~A266 & ~A236;
  assign \new_[20352]_  = ~A235 & \new_[20351]_ ;
  assign \new_[20356]_  = A299 & A298;
  assign \new_[20357]_  = ~A267 & \new_[20356]_ ;
  assign \new_[20358]_  = \new_[20357]_  & \new_[20352]_ ;
  assign \new_[20361]_  = A167 & A168;
  assign \new_[20365]_  = ~A233 & ~A200;
  assign \new_[20366]_  = ~A199 & \new_[20365]_ ;
  assign \new_[20367]_  = \new_[20366]_  & \new_[20361]_ ;
  assign \new_[20371]_  = ~A266 & ~A236;
  assign \new_[20372]_  = ~A235 & \new_[20371]_ ;
  assign \new_[20376]_  = ~A299 & ~A298;
  assign \new_[20377]_  = ~A267 & \new_[20376]_ ;
  assign \new_[20378]_  = \new_[20377]_  & \new_[20372]_ ;
  assign \new_[20381]_  = A167 & A168;
  assign \new_[20385]_  = ~A233 & ~A200;
  assign \new_[20386]_  = ~A199 & \new_[20385]_ ;
  assign \new_[20387]_  = \new_[20386]_  & \new_[20381]_ ;
  assign \new_[20391]_  = ~A265 & ~A236;
  assign \new_[20392]_  = ~A235 & \new_[20391]_ ;
  assign \new_[20396]_  = ~A300 & A298;
  assign \new_[20397]_  = ~A266 & \new_[20396]_ ;
  assign \new_[20398]_  = \new_[20397]_  & \new_[20392]_ ;
  assign \new_[20401]_  = A167 & A168;
  assign \new_[20405]_  = ~A233 & ~A200;
  assign \new_[20406]_  = ~A199 & \new_[20405]_ ;
  assign \new_[20407]_  = \new_[20406]_  & \new_[20401]_ ;
  assign \new_[20411]_  = ~A265 & ~A236;
  assign \new_[20412]_  = ~A235 & \new_[20411]_ ;
  assign \new_[20416]_  = A299 & A298;
  assign \new_[20417]_  = ~A266 & \new_[20416]_ ;
  assign \new_[20418]_  = \new_[20417]_  & \new_[20412]_ ;
  assign \new_[20421]_  = A167 & A168;
  assign \new_[20425]_  = ~A233 & ~A200;
  assign \new_[20426]_  = ~A199 & \new_[20425]_ ;
  assign \new_[20427]_  = \new_[20426]_  & \new_[20421]_ ;
  assign \new_[20431]_  = ~A265 & ~A236;
  assign \new_[20432]_  = ~A235 & \new_[20431]_ ;
  assign \new_[20436]_  = ~A299 & ~A298;
  assign \new_[20437]_  = ~A266 & \new_[20436]_ ;
  assign \new_[20438]_  = \new_[20437]_  & \new_[20432]_ ;
  assign \new_[20441]_  = A167 & A168;
  assign \new_[20445]_  = ~A233 & ~A200;
  assign \new_[20446]_  = ~A199 & \new_[20445]_ ;
  assign \new_[20447]_  = \new_[20446]_  & \new_[20441]_ ;
  assign \new_[20451]_  = A266 & A265;
  assign \new_[20452]_  = ~A234 & \new_[20451]_ ;
  assign \new_[20456]_  = ~A302 & ~A301;
  assign \new_[20457]_  = A298 & \new_[20456]_ ;
  assign \new_[20458]_  = \new_[20457]_  & \new_[20452]_ ;
  assign \new_[20461]_  = A167 & A168;
  assign \new_[20465]_  = ~A233 & ~A200;
  assign \new_[20466]_  = ~A199 & \new_[20465]_ ;
  assign \new_[20467]_  = \new_[20466]_  & \new_[20461]_ ;
  assign \new_[20471]_  = ~A268 & ~A266;
  assign \new_[20472]_  = ~A234 & \new_[20471]_ ;
  assign \new_[20476]_  = ~A300 & A298;
  assign \new_[20477]_  = ~A269 & \new_[20476]_ ;
  assign \new_[20478]_  = \new_[20477]_  & \new_[20472]_ ;
  assign \new_[20481]_  = A167 & A168;
  assign \new_[20485]_  = ~A233 & ~A200;
  assign \new_[20486]_  = ~A199 & \new_[20485]_ ;
  assign \new_[20487]_  = \new_[20486]_  & \new_[20481]_ ;
  assign \new_[20491]_  = ~A268 & ~A266;
  assign \new_[20492]_  = ~A234 & \new_[20491]_ ;
  assign \new_[20496]_  = A299 & A298;
  assign \new_[20497]_  = ~A269 & \new_[20496]_ ;
  assign \new_[20498]_  = \new_[20497]_  & \new_[20492]_ ;
  assign \new_[20501]_  = A167 & A168;
  assign \new_[20505]_  = ~A233 & ~A200;
  assign \new_[20506]_  = ~A199 & \new_[20505]_ ;
  assign \new_[20507]_  = \new_[20506]_  & \new_[20501]_ ;
  assign \new_[20511]_  = ~A268 & ~A266;
  assign \new_[20512]_  = ~A234 & \new_[20511]_ ;
  assign \new_[20516]_  = ~A299 & ~A298;
  assign \new_[20517]_  = ~A269 & \new_[20516]_ ;
  assign \new_[20518]_  = \new_[20517]_  & \new_[20512]_ ;
  assign \new_[20521]_  = A167 & A168;
  assign \new_[20525]_  = ~A233 & ~A200;
  assign \new_[20526]_  = ~A199 & \new_[20525]_ ;
  assign \new_[20527]_  = \new_[20526]_  & \new_[20521]_ ;
  assign \new_[20531]_  = ~A267 & ~A266;
  assign \new_[20532]_  = ~A234 & \new_[20531]_ ;
  assign \new_[20536]_  = ~A302 & ~A301;
  assign \new_[20537]_  = A298 & \new_[20536]_ ;
  assign \new_[20538]_  = \new_[20537]_  & \new_[20532]_ ;
  assign \new_[20541]_  = A167 & A168;
  assign \new_[20545]_  = ~A233 & ~A200;
  assign \new_[20546]_  = ~A199 & \new_[20545]_ ;
  assign \new_[20547]_  = \new_[20546]_  & \new_[20541]_ ;
  assign \new_[20551]_  = ~A266 & ~A265;
  assign \new_[20552]_  = ~A234 & \new_[20551]_ ;
  assign \new_[20556]_  = ~A302 & ~A301;
  assign \new_[20557]_  = A298 & \new_[20556]_ ;
  assign \new_[20558]_  = \new_[20557]_  & \new_[20552]_ ;
  assign \new_[20561]_  = A167 & A168;
  assign \new_[20565]_  = ~A232 & ~A200;
  assign \new_[20566]_  = ~A199 & \new_[20565]_ ;
  assign \new_[20567]_  = \new_[20566]_  & \new_[20561]_ ;
  assign \new_[20571]_  = A266 & A265;
  assign \new_[20572]_  = ~A233 & \new_[20571]_ ;
  assign \new_[20576]_  = ~A302 & ~A301;
  assign \new_[20577]_  = A298 & \new_[20576]_ ;
  assign \new_[20578]_  = \new_[20577]_  & \new_[20572]_ ;
  assign \new_[20581]_  = A167 & A168;
  assign \new_[20585]_  = ~A232 & ~A200;
  assign \new_[20586]_  = ~A199 & \new_[20585]_ ;
  assign \new_[20587]_  = \new_[20586]_  & \new_[20581]_ ;
  assign \new_[20591]_  = ~A268 & ~A266;
  assign \new_[20592]_  = ~A233 & \new_[20591]_ ;
  assign \new_[20596]_  = ~A300 & A298;
  assign \new_[20597]_  = ~A269 & \new_[20596]_ ;
  assign \new_[20598]_  = \new_[20597]_  & \new_[20592]_ ;
  assign \new_[20601]_  = A167 & A168;
  assign \new_[20605]_  = ~A232 & ~A200;
  assign \new_[20606]_  = ~A199 & \new_[20605]_ ;
  assign \new_[20607]_  = \new_[20606]_  & \new_[20601]_ ;
  assign \new_[20611]_  = ~A268 & ~A266;
  assign \new_[20612]_  = ~A233 & \new_[20611]_ ;
  assign \new_[20616]_  = A299 & A298;
  assign \new_[20617]_  = ~A269 & \new_[20616]_ ;
  assign \new_[20618]_  = \new_[20617]_  & \new_[20612]_ ;
  assign \new_[20621]_  = A167 & A168;
  assign \new_[20625]_  = ~A232 & ~A200;
  assign \new_[20626]_  = ~A199 & \new_[20625]_ ;
  assign \new_[20627]_  = \new_[20626]_  & \new_[20621]_ ;
  assign \new_[20631]_  = ~A268 & ~A266;
  assign \new_[20632]_  = ~A233 & \new_[20631]_ ;
  assign \new_[20636]_  = ~A299 & ~A298;
  assign \new_[20637]_  = ~A269 & \new_[20636]_ ;
  assign \new_[20638]_  = \new_[20637]_  & \new_[20632]_ ;
  assign \new_[20641]_  = A167 & A168;
  assign \new_[20645]_  = ~A232 & ~A200;
  assign \new_[20646]_  = ~A199 & \new_[20645]_ ;
  assign \new_[20647]_  = \new_[20646]_  & \new_[20641]_ ;
  assign \new_[20651]_  = ~A267 & ~A266;
  assign \new_[20652]_  = ~A233 & \new_[20651]_ ;
  assign \new_[20656]_  = ~A302 & ~A301;
  assign \new_[20657]_  = A298 & \new_[20656]_ ;
  assign \new_[20658]_  = \new_[20657]_  & \new_[20652]_ ;
  assign \new_[20661]_  = A167 & A168;
  assign \new_[20665]_  = ~A232 & ~A200;
  assign \new_[20666]_  = ~A199 & \new_[20665]_ ;
  assign \new_[20667]_  = \new_[20666]_  & \new_[20661]_ ;
  assign \new_[20671]_  = ~A266 & ~A265;
  assign \new_[20672]_  = ~A233 & \new_[20671]_ ;
  assign \new_[20676]_  = ~A302 & ~A301;
  assign \new_[20677]_  = A298 & \new_[20676]_ ;
  assign \new_[20678]_  = \new_[20677]_  & \new_[20672]_ ;
  assign \new_[20681]_  = ~A167 & A170;
  assign \new_[20685]_  = A200 & ~A199;
  assign \new_[20686]_  = ~A166 & \new_[20685]_ ;
  assign \new_[20687]_  = \new_[20686]_  & \new_[20681]_ ;
  assign \new_[20691]_  = A265 & A233;
  assign \new_[20692]_  = A232 & \new_[20691]_ ;
  assign \new_[20696]_  = ~A300 & ~A299;
  assign \new_[20697]_  = ~A267 & \new_[20696]_ ;
  assign \new_[20698]_  = \new_[20697]_  & \new_[20692]_ ;
  assign \new_[20701]_  = ~A167 & A170;
  assign \new_[20705]_  = A200 & ~A199;
  assign \new_[20706]_  = ~A166 & \new_[20705]_ ;
  assign \new_[20707]_  = \new_[20706]_  & \new_[20701]_ ;
  assign \new_[20711]_  = A265 & A233;
  assign \new_[20712]_  = A232 & \new_[20711]_ ;
  assign \new_[20716]_  = A299 & A298;
  assign \new_[20717]_  = ~A267 & \new_[20716]_ ;
  assign \new_[20718]_  = \new_[20717]_  & \new_[20712]_ ;
  assign \new_[20721]_  = ~A167 & A170;
  assign \new_[20725]_  = A200 & ~A199;
  assign \new_[20726]_  = ~A166 & \new_[20725]_ ;
  assign \new_[20727]_  = \new_[20726]_  & \new_[20721]_ ;
  assign \new_[20731]_  = A265 & A233;
  assign \new_[20732]_  = A232 & \new_[20731]_ ;
  assign \new_[20736]_  = ~A299 & ~A298;
  assign \new_[20737]_  = ~A267 & \new_[20736]_ ;
  assign \new_[20738]_  = \new_[20737]_  & \new_[20732]_ ;
  assign \new_[20741]_  = ~A167 & A170;
  assign \new_[20745]_  = A200 & ~A199;
  assign \new_[20746]_  = ~A166 & \new_[20745]_ ;
  assign \new_[20747]_  = \new_[20746]_  & \new_[20741]_ ;
  assign \new_[20751]_  = A265 & A233;
  assign \new_[20752]_  = A232 & \new_[20751]_ ;
  assign \new_[20756]_  = ~A300 & ~A299;
  assign \new_[20757]_  = A266 & \new_[20756]_ ;
  assign \new_[20758]_  = \new_[20757]_  & \new_[20752]_ ;
  assign \new_[20761]_  = ~A167 & A170;
  assign \new_[20765]_  = A200 & ~A199;
  assign \new_[20766]_  = ~A166 & \new_[20765]_ ;
  assign \new_[20767]_  = \new_[20766]_  & \new_[20761]_ ;
  assign \new_[20771]_  = A265 & A233;
  assign \new_[20772]_  = A232 & \new_[20771]_ ;
  assign \new_[20776]_  = A299 & A298;
  assign \new_[20777]_  = A266 & \new_[20776]_ ;
  assign \new_[20778]_  = \new_[20777]_  & \new_[20772]_ ;
  assign \new_[20781]_  = ~A167 & A170;
  assign \new_[20785]_  = A200 & ~A199;
  assign \new_[20786]_  = ~A166 & \new_[20785]_ ;
  assign \new_[20787]_  = \new_[20786]_  & \new_[20781]_ ;
  assign \new_[20791]_  = A265 & A233;
  assign \new_[20792]_  = A232 & \new_[20791]_ ;
  assign \new_[20796]_  = ~A299 & ~A298;
  assign \new_[20797]_  = A266 & \new_[20796]_ ;
  assign \new_[20798]_  = \new_[20797]_  & \new_[20792]_ ;
  assign \new_[20801]_  = ~A167 & A170;
  assign \new_[20805]_  = A200 & ~A199;
  assign \new_[20806]_  = ~A166 & \new_[20805]_ ;
  assign \new_[20807]_  = \new_[20806]_  & \new_[20801]_ ;
  assign \new_[20811]_  = ~A265 & A233;
  assign \new_[20812]_  = A232 & \new_[20811]_ ;
  assign \new_[20816]_  = ~A300 & ~A299;
  assign \new_[20817]_  = ~A266 & \new_[20816]_ ;
  assign \new_[20818]_  = \new_[20817]_  & \new_[20812]_ ;
  assign \new_[20821]_  = ~A167 & A170;
  assign \new_[20825]_  = A200 & ~A199;
  assign \new_[20826]_  = ~A166 & \new_[20825]_ ;
  assign \new_[20827]_  = \new_[20826]_  & \new_[20821]_ ;
  assign \new_[20831]_  = ~A265 & A233;
  assign \new_[20832]_  = A232 & \new_[20831]_ ;
  assign \new_[20836]_  = A299 & A298;
  assign \new_[20837]_  = ~A266 & \new_[20836]_ ;
  assign \new_[20838]_  = \new_[20837]_  & \new_[20832]_ ;
  assign \new_[20841]_  = ~A167 & A170;
  assign \new_[20845]_  = A200 & ~A199;
  assign \new_[20846]_  = ~A166 & \new_[20845]_ ;
  assign \new_[20847]_  = \new_[20846]_  & \new_[20841]_ ;
  assign \new_[20851]_  = ~A265 & A233;
  assign \new_[20852]_  = A232 & \new_[20851]_ ;
  assign \new_[20856]_  = ~A299 & ~A298;
  assign \new_[20857]_  = ~A266 & \new_[20856]_ ;
  assign \new_[20858]_  = \new_[20857]_  & \new_[20852]_ ;
  assign \new_[20861]_  = ~A167 & A170;
  assign \new_[20865]_  = A200 & ~A199;
  assign \new_[20866]_  = ~A166 & \new_[20865]_ ;
  assign \new_[20867]_  = \new_[20866]_  & \new_[20861]_ ;
  assign \new_[20871]_  = A298 & A233;
  assign \new_[20872]_  = ~A232 & \new_[20871]_ ;
  assign \new_[20876]_  = A301 & A300;
  assign \new_[20877]_  = ~A299 & \new_[20876]_ ;
  assign \new_[20878]_  = \new_[20877]_  & \new_[20872]_ ;
  assign \new_[20881]_  = ~A167 & A170;
  assign \new_[20885]_  = A200 & ~A199;
  assign \new_[20886]_  = ~A166 & \new_[20885]_ ;
  assign \new_[20887]_  = \new_[20886]_  & \new_[20881]_ ;
  assign \new_[20891]_  = A298 & A233;
  assign \new_[20892]_  = ~A232 & \new_[20891]_ ;
  assign \new_[20896]_  = A302 & A300;
  assign \new_[20897]_  = ~A299 & \new_[20896]_ ;
  assign \new_[20898]_  = \new_[20897]_  & \new_[20892]_ ;
  assign \new_[20901]_  = ~A167 & A170;
  assign \new_[20905]_  = A200 & ~A199;
  assign \new_[20906]_  = ~A166 & \new_[20905]_ ;
  assign \new_[20907]_  = \new_[20906]_  & \new_[20901]_ ;
  assign \new_[20911]_  = A265 & A233;
  assign \new_[20912]_  = ~A232 & \new_[20911]_ ;
  assign \new_[20916]_  = A268 & A267;
  assign \new_[20917]_  = ~A266 & \new_[20916]_ ;
  assign \new_[20918]_  = \new_[20917]_  & \new_[20912]_ ;
  assign \new_[20921]_  = ~A167 & A170;
  assign \new_[20925]_  = A200 & ~A199;
  assign \new_[20926]_  = ~A166 & \new_[20925]_ ;
  assign \new_[20927]_  = \new_[20926]_  & \new_[20921]_ ;
  assign \new_[20931]_  = A265 & A233;
  assign \new_[20932]_  = ~A232 & \new_[20931]_ ;
  assign \new_[20936]_  = A269 & A267;
  assign \new_[20937]_  = ~A266 & \new_[20936]_ ;
  assign \new_[20938]_  = \new_[20937]_  & \new_[20932]_ ;
  assign \new_[20941]_  = ~A167 & A170;
  assign \new_[20945]_  = A200 & ~A199;
  assign \new_[20946]_  = ~A166 & \new_[20945]_ ;
  assign \new_[20947]_  = \new_[20946]_  & \new_[20941]_ ;
  assign \new_[20951]_  = A265 & ~A234;
  assign \new_[20952]_  = ~A233 & \new_[20951]_ ;
  assign \new_[20956]_  = ~A300 & A298;
  assign \new_[20957]_  = A266 & \new_[20956]_ ;
  assign \new_[20958]_  = \new_[20957]_  & \new_[20952]_ ;
  assign \new_[20961]_  = ~A167 & A170;
  assign \new_[20965]_  = A200 & ~A199;
  assign \new_[20966]_  = ~A166 & \new_[20965]_ ;
  assign \new_[20967]_  = \new_[20966]_  & \new_[20961]_ ;
  assign \new_[20971]_  = A265 & ~A234;
  assign \new_[20972]_  = ~A233 & \new_[20971]_ ;
  assign \new_[20976]_  = A299 & A298;
  assign \new_[20977]_  = A266 & \new_[20976]_ ;
  assign \new_[20978]_  = \new_[20977]_  & \new_[20972]_ ;
  assign \new_[20981]_  = ~A167 & A170;
  assign \new_[20985]_  = A200 & ~A199;
  assign \new_[20986]_  = ~A166 & \new_[20985]_ ;
  assign \new_[20987]_  = \new_[20986]_  & \new_[20981]_ ;
  assign \new_[20991]_  = A265 & ~A234;
  assign \new_[20992]_  = ~A233 & \new_[20991]_ ;
  assign \new_[20996]_  = ~A299 & ~A298;
  assign \new_[20997]_  = A266 & \new_[20996]_ ;
  assign \new_[20998]_  = \new_[20997]_  & \new_[20992]_ ;
  assign \new_[21001]_  = ~A167 & A170;
  assign \new_[21005]_  = A200 & ~A199;
  assign \new_[21006]_  = ~A166 & \new_[21005]_ ;
  assign \new_[21007]_  = \new_[21006]_  & \new_[21001]_ ;
  assign \new_[21011]_  = ~A266 & ~A234;
  assign \new_[21012]_  = ~A233 & \new_[21011]_ ;
  assign \new_[21016]_  = ~A300 & A298;
  assign \new_[21017]_  = ~A267 & \new_[21016]_ ;
  assign \new_[21018]_  = \new_[21017]_  & \new_[21012]_ ;
  assign \new_[21021]_  = ~A167 & A170;
  assign \new_[21025]_  = A200 & ~A199;
  assign \new_[21026]_  = ~A166 & \new_[21025]_ ;
  assign \new_[21027]_  = \new_[21026]_  & \new_[21021]_ ;
  assign \new_[21031]_  = ~A266 & ~A234;
  assign \new_[21032]_  = ~A233 & \new_[21031]_ ;
  assign \new_[21036]_  = A299 & A298;
  assign \new_[21037]_  = ~A267 & \new_[21036]_ ;
  assign \new_[21038]_  = \new_[21037]_  & \new_[21032]_ ;
  assign \new_[21041]_  = ~A167 & A170;
  assign \new_[21045]_  = A200 & ~A199;
  assign \new_[21046]_  = ~A166 & \new_[21045]_ ;
  assign \new_[21047]_  = \new_[21046]_  & \new_[21041]_ ;
  assign \new_[21051]_  = ~A266 & ~A234;
  assign \new_[21052]_  = ~A233 & \new_[21051]_ ;
  assign \new_[21056]_  = ~A299 & ~A298;
  assign \new_[21057]_  = ~A267 & \new_[21056]_ ;
  assign \new_[21058]_  = \new_[21057]_  & \new_[21052]_ ;
  assign \new_[21061]_  = ~A167 & A170;
  assign \new_[21065]_  = A200 & ~A199;
  assign \new_[21066]_  = ~A166 & \new_[21065]_ ;
  assign \new_[21067]_  = \new_[21066]_  & \new_[21061]_ ;
  assign \new_[21071]_  = ~A265 & ~A234;
  assign \new_[21072]_  = ~A233 & \new_[21071]_ ;
  assign \new_[21076]_  = ~A300 & A298;
  assign \new_[21077]_  = ~A266 & \new_[21076]_ ;
  assign \new_[21078]_  = \new_[21077]_  & \new_[21072]_ ;
  assign \new_[21081]_  = ~A167 & A170;
  assign \new_[21085]_  = A200 & ~A199;
  assign \new_[21086]_  = ~A166 & \new_[21085]_ ;
  assign \new_[21087]_  = \new_[21086]_  & \new_[21081]_ ;
  assign \new_[21091]_  = ~A265 & ~A234;
  assign \new_[21092]_  = ~A233 & \new_[21091]_ ;
  assign \new_[21096]_  = A299 & A298;
  assign \new_[21097]_  = ~A266 & \new_[21096]_ ;
  assign \new_[21098]_  = \new_[21097]_  & \new_[21092]_ ;
  assign \new_[21101]_  = ~A167 & A170;
  assign \new_[21105]_  = A200 & ~A199;
  assign \new_[21106]_  = ~A166 & \new_[21105]_ ;
  assign \new_[21107]_  = \new_[21106]_  & \new_[21101]_ ;
  assign \new_[21111]_  = ~A265 & ~A234;
  assign \new_[21112]_  = ~A233 & \new_[21111]_ ;
  assign \new_[21116]_  = ~A299 & ~A298;
  assign \new_[21117]_  = ~A266 & \new_[21116]_ ;
  assign \new_[21118]_  = \new_[21117]_  & \new_[21112]_ ;
  assign \new_[21121]_  = ~A167 & A170;
  assign \new_[21125]_  = A200 & ~A199;
  assign \new_[21126]_  = ~A166 & \new_[21125]_ ;
  assign \new_[21127]_  = \new_[21126]_  & \new_[21121]_ ;
  assign \new_[21131]_  = A234 & ~A233;
  assign \new_[21132]_  = A232 & \new_[21131]_ ;
  assign \new_[21136]_  = A299 & ~A298;
  assign \new_[21137]_  = A235 & \new_[21136]_ ;
  assign \new_[21138]_  = \new_[21137]_  & \new_[21132]_ ;
  assign \new_[21141]_  = ~A167 & A170;
  assign \new_[21145]_  = A200 & ~A199;
  assign \new_[21146]_  = ~A166 & \new_[21145]_ ;
  assign \new_[21147]_  = \new_[21146]_  & \new_[21141]_ ;
  assign \new_[21151]_  = A234 & ~A233;
  assign \new_[21152]_  = A232 & \new_[21151]_ ;
  assign \new_[21156]_  = A266 & ~A265;
  assign \new_[21157]_  = A235 & \new_[21156]_ ;
  assign \new_[21158]_  = \new_[21157]_  & \new_[21152]_ ;
  assign \new_[21161]_  = ~A167 & A170;
  assign \new_[21165]_  = A200 & ~A199;
  assign \new_[21166]_  = ~A166 & \new_[21165]_ ;
  assign \new_[21167]_  = \new_[21166]_  & \new_[21161]_ ;
  assign \new_[21171]_  = A234 & ~A233;
  assign \new_[21172]_  = A232 & \new_[21171]_ ;
  assign \new_[21176]_  = A299 & ~A298;
  assign \new_[21177]_  = A236 & \new_[21176]_ ;
  assign \new_[21178]_  = \new_[21177]_  & \new_[21172]_ ;
  assign \new_[21181]_  = ~A167 & A170;
  assign \new_[21185]_  = A200 & ~A199;
  assign \new_[21186]_  = ~A166 & \new_[21185]_ ;
  assign \new_[21187]_  = \new_[21186]_  & \new_[21181]_ ;
  assign \new_[21191]_  = A234 & ~A233;
  assign \new_[21192]_  = A232 & \new_[21191]_ ;
  assign \new_[21196]_  = A266 & ~A265;
  assign \new_[21197]_  = A236 & \new_[21196]_ ;
  assign \new_[21198]_  = \new_[21197]_  & \new_[21192]_ ;
  assign \new_[21201]_  = ~A167 & A170;
  assign \new_[21205]_  = A200 & ~A199;
  assign \new_[21206]_  = ~A166 & \new_[21205]_ ;
  assign \new_[21207]_  = \new_[21206]_  & \new_[21201]_ ;
  assign \new_[21211]_  = A265 & ~A233;
  assign \new_[21212]_  = ~A232 & \new_[21211]_ ;
  assign \new_[21216]_  = ~A300 & A298;
  assign \new_[21217]_  = A266 & \new_[21216]_ ;
  assign \new_[21218]_  = \new_[21217]_  & \new_[21212]_ ;
  assign \new_[21221]_  = ~A167 & A170;
  assign \new_[21225]_  = A200 & ~A199;
  assign \new_[21226]_  = ~A166 & \new_[21225]_ ;
  assign \new_[21227]_  = \new_[21226]_  & \new_[21221]_ ;
  assign \new_[21231]_  = A265 & ~A233;
  assign \new_[21232]_  = ~A232 & \new_[21231]_ ;
  assign \new_[21236]_  = A299 & A298;
  assign \new_[21237]_  = A266 & \new_[21236]_ ;
  assign \new_[21238]_  = \new_[21237]_  & \new_[21232]_ ;
  assign \new_[21241]_  = ~A167 & A170;
  assign \new_[21245]_  = A200 & ~A199;
  assign \new_[21246]_  = ~A166 & \new_[21245]_ ;
  assign \new_[21247]_  = \new_[21246]_  & \new_[21241]_ ;
  assign \new_[21251]_  = A265 & ~A233;
  assign \new_[21252]_  = ~A232 & \new_[21251]_ ;
  assign \new_[21256]_  = ~A299 & ~A298;
  assign \new_[21257]_  = A266 & \new_[21256]_ ;
  assign \new_[21258]_  = \new_[21257]_  & \new_[21252]_ ;
  assign \new_[21261]_  = ~A167 & A170;
  assign \new_[21265]_  = A200 & ~A199;
  assign \new_[21266]_  = ~A166 & \new_[21265]_ ;
  assign \new_[21267]_  = \new_[21266]_  & \new_[21261]_ ;
  assign \new_[21271]_  = ~A266 & ~A233;
  assign \new_[21272]_  = ~A232 & \new_[21271]_ ;
  assign \new_[21276]_  = ~A300 & A298;
  assign \new_[21277]_  = ~A267 & \new_[21276]_ ;
  assign \new_[21278]_  = \new_[21277]_  & \new_[21272]_ ;
  assign \new_[21281]_  = ~A167 & A170;
  assign \new_[21285]_  = A200 & ~A199;
  assign \new_[21286]_  = ~A166 & \new_[21285]_ ;
  assign \new_[21287]_  = \new_[21286]_  & \new_[21281]_ ;
  assign \new_[21291]_  = ~A266 & ~A233;
  assign \new_[21292]_  = ~A232 & \new_[21291]_ ;
  assign \new_[21296]_  = A299 & A298;
  assign \new_[21297]_  = ~A267 & \new_[21296]_ ;
  assign \new_[21298]_  = \new_[21297]_  & \new_[21292]_ ;
  assign \new_[21301]_  = ~A167 & A170;
  assign \new_[21305]_  = A200 & ~A199;
  assign \new_[21306]_  = ~A166 & \new_[21305]_ ;
  assign \new_[21307]_  = \new_[21306]_  & \new_[21301]_ ;
  assign \new_[21311]_  = ~A266 & ~A233;
  assign \new_[21312]_  = ~A232 & \new_[21311]_ ;
  assign \new_[21316]_  = ~A299 & ~A298;
  assign \new_[21317]_  = ~A267 & \new_[21316]_ ;
  assign \new_[21318]_  = \new_[21317]_  & \new_[21312]_ ;
  assign \new_[21321]_  = ~A167 & A170;
  assign \new_[21325]_  = A200 & ~A199;
  assign \new_[21326]_  = ~A166 & \new_[21325]_ ;
  assign \new_[21327]_  = \new_[21326]_  & \new_[21321]_ ;
  assign \new_[21331]_  = ~A265 & ~A233;
  assign \new_[21332]_  = ~A232 & \new_[21331]_ ;
  assign \new_[21336]_  = ~A300 & A298;
  assign \new_[21337]_  = ~A266 & \new_[21336]_ ;
  assign \new_[21338]_  = \new_[21337]_  & \new_[21332]_ ;
  assign \new_[21341]_  = ~A167 & A170;
  assign \new_[21345]_  = A200 & ~A199;
  assign \new_[21346]_  = ~A166 & \new_[21345]_ ;
  assign \new_[21347]_  = \new_[21346]_  & \new_[21341]_ ;
  assign \new_[21351]_  = ~A265 & ~A233;
  assign \new_[21352]_  = ~A232 & \new_[21351]_ ;
  assign \new_[21356]_  = A299 & A298;
  assign \new_[21357]_  = ~A266 & \new_[21356]_ ;
  assign \new_[21358]_  = \new_[21357]_  & \new_[21352]_ ;
  assign \new_[21361]_  = ~A167 & A170;
  assign \new_[21365]_  = A200 & ~A199;
  assign \new_[21366]_  = ~A166 & \new_[21365]_ ;
  assign \new_[21367]_  = \new_[21366]_  & \new_[21361]_ ;
  assign \new_[21371]_  = ~A265 & ~A233;
  assign \new_[21372]_  = ~A232 & \new_[21371]_ ;
  assign \new_[21376]_  = ~A299 & ~A298;
  assign \new_[21377]_  = ~A266 & \new_[21376]_ ;
  assign \new_[21378]_  = \new_[21377]_  & \new_[21372]_ ;
  assign \new_[21381]_  = ~A167 & A170;
  assign \new_[21385]_  = ~A200 & A199;
  assign \new_[21386]_  = ~A166 & \new_[21385]_ ;
  assign \new_[21387]_  = \new_[21386]_  & \new_[21381]_ ;
  assign \new_[21391]_  = ~A232 & A202;
  assign \new_[21392]_  = A201 & \new_[21391]_ ;
  assign \new_[21396]_  = A299 & ~A298;
  assign \new_[21397]_  = A233 & \new_[21396]_ ;
  assign \new_[21398]_  = \new_[21397]_  & \new_[21392]_ ;
  assign \new_[21401]_  = ~A167 & A170;
  assign \new_[21405]_  = ~A200 & A199;
  assign \new_[21406]_  = ~A166 & \new_[21405]_ ;
  assign \new_[21407]_  = \new_[21406]_  & \new_[21401]_ ;
  assign \new_[21411]_  = ~A232 & A202;
  assign \new_[21412]_  = A201 & \new_[21411]_ ;
  assign \new_[21416]_  = A266 & ~A265;
  assign \new_[21417]_  = A233 & \new_[21416]_ ;
  assign \new_[21418]_  = \new_[21417]_  & \new_[21412]_ ;
  assign \new_[21421]_  = ~A167 & A170;
  assign \new_[21425]_  = ~A200 & A199;
  assign \new_[21426]_  = ~A166 & \new_[21425]_ ;
  assign \new_[21427]_  = \new_[21426]_  & \new_[21421]_ ;
  assign \new_[21431]_  = ~A232 & A203;
  assign \new_[21432]_  = A201 & \new_[21431]_ ;
  assign \new_[21436]_  = A299 & ~A298;
  assign \new_[21437]_  = A233 & \new_[21436]_ ;
  assign \new_[21438]_  = \new_[21437]_  & \new_[21432]_ ;
  assign \new_[21441]_  = ~A167 & A170;
  assign \new_[21445]_  = ~A200 & A199;
  assign \new_[21446]_  = ~A166 & \new_[21445]_ ;
  assign \new_[21447]_  = \new_[21446]_  & \new_[21441]_ ;
  assign \new_[21451]_  = ~A232 & A203;
  assign \new_[21452]_  = A201 & \new_[21451]_ ;
  assign \new_[21456]_  = A266 & ~A265;
  assign \new_[21457]_  = A233 & \new_[21456]_ ;
  assign \new_[21458]_  = \new_[21457]_  & \new_[21452]_ ;
  assign \new_[21461]_  = A169 & ~A170;
  assign \new_[21465]_  = ~A200 & A166;
  assign \new_[21466]_  = A167 & \new_[21465]_ ;
  assign \new_[21467]_  = \new_[21466]_  & \new_[21461]_ ;
  assign \new_[21471]_  = ~A232 & ~A203;
  assign \new_[21472]_  = ~A202 & \new_[21471]_ ;
  assign \new_[21476]_  = A299 & ~A298;
  assign \new_[21477]_  = A233 & \new_[21476]_ ;
  assign \new_[21478]_  = \new_[21477]_  & \new_[21472]_ ;
  assign \new_[21481]_  = A169 & ~A170;
  assign \new_[21485]_  = ~A200 & A166;
  assign \new_[21486]_  = A167 & \new_[21485]_ ;
  assign \new_[21487]_  = \new_[21486]_  & \new_[21481]_ ;
  assign \new_[21491]_  = ~A232 & ~A203;
  assign \new_[21492]_  = ~A202 & \new_[21491]_ ;
  assign \new_[21496]_  = A266 & ~A265;
  assign \new_[21497]_  = A233 & \new_[21496]_ ;
  assign \new_[21498]_  = \new_[21497]_  & \new_[21492]_ ;
  assign \new_[21501]_  = A169 & ~A170;
  assign \new_[21505]_  = ~A200 & ~A166;
  assign \new_[21506]_  = ~A167 & \new_[21505]_ ;
  assign \new_[21507]_  = \new_[21506]_  & \new_[21501]_ ;
  assign \new_[21511]_  = ~A232 & ~A203;
  assign \new_[21512]_  = ~A202 & \new_[21511]_ ;
  assign \new_[21516]_  = A299 & ~A298;
  assign \new_[21517]_  = A233 & \new_[21516]_ ;
  assign \new_[21518]_  = \new_[21517]_  & \new_[21512]_ ;
  assign \new_[21521]_  = A169 & ~A170;
  assign \new_[21525]_  = ~A200 & ~A166;
  assign \new_[21526]_  = ~A167 & \new_[21525]_ ;
  assign \new_[21527]_  = \new_[21526]_  & \new_[21521]_ ;
  assign \new_[21531]_  = ~A232 & ~A203;
  assign \new_[21532]_  = ~A202 & \new_[21531]_ ;
  assign \new_[21536]_  = A266 & ~A265;
  assign \new_[21537]_  = A233 & \new_[21536]_ ;
  assign \new_[21538]_  = \new_[21537]_  & \new_[21532]_ ;
  assign \new_[21541]_  = ~A167 & ~A169;
  assign \new_[21545]_  = A200 & ~A199;
  assign \new_[21546]_  = ~A166 & \new_[21545]_ ;
  assign \new_[21547]_  = \new_[21546]_  & \new_[21541]_ ;
  assign \new_[21551]_  = A265 & A233;
  assign \new_[21552]_  = A232 & \new_[21551]_ ;
  assign \new_[21556]_  = ~A300 & ~A299;
  assign \new_[21557]_  = ~A267 & \new_[21556]_ ;
  assign \new_[21558]_  = \new_[21557]_  & \new_[21552]_ ;
  assign \new_[21561]_  = ~A167 & ~A169;
  assign \new_[21565]_  = A200 & ~A199;
  assign \new_[21566]_  = ~A166 & \new_[21565]_ ;
  assign \new_[21567]_  = \new_[21566]_  & \new_[21561]_ ;
  assign \new_[21571]_  = A265 & A233;
  assign \new_[21572]_  = A232 & \new_[21571]_ ;
  assign \new_[21576]_  = A299 & A298;
  assign \new_[21577]_  = ~A267 & \new_[21576]_ ;
  assign \new_[21578]_  = \new_[21577]_  & \new_[21572]_ ;
  assign \new_[21581]_  = ~A167 & ~A169;
  assign \new_[21585]_  = A200 & ~A199;
  assign \new_[21586]_  = ~A166 & \new_[21585]_ ;
  assign \new_[21587]_  = \new_[21586]_  & \new_[21581]_ ;
  assign \new_[21591]_  = A265 & A233;
  assign \new_[21592]_  = A232 & \new_[21591]_ ;
  assign \new_[21596]_  = ~A299 & ~A298;
  assign \new_[21597]_  = ~A267 & \new_[21596]_ ;
  assign \new_[21598]_  = \new_[21597]_  & \new_[21592]_ ;
  assign \new_[21601]_  = ~A167 & ~A169;
  assign \new_[21605]_  = A200 & ~A199;
  assign \new_[21606]_  = ~A166 & \new_[21605]_ ;
  assign \new_[21607]_  = \new_[21606]_  & \new_[21601]_ ;
  assign \new_[21611]_  = A265 & A233;
  assign \new_[21612]_  = A232 & \new_[21611]_ ;
  assign \new_[21616]_  = ~A300 & ~A299;
  assign \new_[21617]_  = A266 & \new_[21616]_ ;
  assign \new_[21618]_  = \new_[21617]_  & \new_[21612]_ ;
  assign \new_[21621]_  = ~A167 & ~A169;
  assign \new_[21625]_  = A200 & ~A199;
  assign \new_[21626]_  = ~A166 & \new_[21625]_ ;
  assign \new_[21627]_  = \new_[21626]_  & \new_[21621]_ ;
  assign \new_[21631]_  = A265 & A233;
  assign \new_[21632]_  = A232 & \new_[21631]_ ;
  assign \new_[21636]_  = A299 & A298;
  assign \new_[21637]_  = A266 & \new_[21636]_ ;
  assign \new_[21638]_  = \new_[21637]_  & \new_[21632]_ ;
  assign \new_[21641]_  = ~A167 & ~A169;
  assign \new_[21645]_  = A200 & ~A199;
  assign \new_[21646]_  = ~A166 & \new_[21645]_ ;
  assign \new_[21647]_  = \new_[21646]_  & \new_[21641]_ ;
  assign \new_[21651]_  = A265 & A233;
  assign \new_[21652]_  = A232 & \new_[21651]_ ;
  assign \new_[21656]_  = ~A299 & ~A298;
  assign \new_[21657]_  = A266 & \new_[21656]_ ;
  assign \new_[21658]_  = \new_[21657]_  & \new_[21652]_ ;
  assign \new_[21661]_  = ~A167 & ~A169;
  assign \new_[21665]_  = A200 & ~A199;
  assign \new_[21666]_  = ~A166 & \new_[21665]_ ;
  assign \new_[21667]_  = \new_[21666]_  & \new_[21661]_ ;
  assign \new_[21671]_  = ~A265 & A233;
  assign \new_[21672]_  = A232 & \new_[21671]_ ;
  assign \new_[21676]_  = ~A300 & ~A299;
  assign \new_[21677]_  = ~A266 & \new_[21676]_ ;
  assign \new_[21678]_  = \new_[21677]_  & \new_[21672]_ ;
  assign \new_[21681]_  = ~A167 & ~A169;
  assign \new_[21685]_  = A200 & ~A199;
  assign \new_[21686]_  = ~A166 & \new_[21685]_ ;
  assign \new_[21687]_  = \new_[21686]_  & \new_[21681]_ ;
  assign \new_[21691]_  = ~A265 & A233;
  assign \new_[21692]_  = A232 & \new_[21691]_ ;
  assign \new_[21696]_  = A299 & A298;
  assign \new_[21697]_  = ~A266 & \new_[21696]_ ;
  assign \new_[21698]_  = \new_[21697]_  & \new_[21692]_ ;
  assign \new_[21701]_  = ~A167 & ~A169;
  assign \new_[21705]_  = A200 & ~A199;
  assign \new_[21706]_  = ~A166 & \new_[21705]_ ;
  assign \new_[21707]_  = \new_[21706]_  & \new_[21701]_ ;
  assign \new_[21711]_  = ~A265 & A233;
  assign \new_[21712]_  = A232 & \new_[21711]_ ;
  assign \new_[21716]_  = ~A299 & ~A298;
  assign \new_[21717]_  = ~A266 & \new_[21716]_ ;
  assign \new_[21718]_  = \new_[21717]_  & \new_[21712]_ ;
  assign \new_[21721]_  = ~A167 & ~A169;
  assign \new_[21725]_  = A200 & ~A199;
  assign \new_[21726]_  = ~A166 & \new_[21725]_ ;
  assign \new_[21727]_  = \new_[21726]_  & \new_[21721]_ ;
  assign \new_[21731]_  = A298 & A233;
  assign \new_[21732]_  = ~A232 & \new_[21731]_ ;
  assign \new_[21736]_  = A301 & A300;
  assign \new_[21737]_  = ~A299 & \new_[21736]_ ;
  assign \new_[21738]_  = \new_[21737]_  & \new_[21732]_ ;
  assign \new_[21741]_  = ~A167 & ~A169;
  assign \new_[21745]_  = A200 & ~A199;
  assign \new_[21746]_  = ~A166 & \new_[21745]_ ;
  assign \new_[21747]_  = \new_[21746]_  & \new_[21741]_ ;
  assign \new_[21751]_  = A298 & A233;
  assign \new_[21752]_  = ~A232 & \new_[21751]_ ;
  assign \new_[21756]_  = A302 & A300;
  assign \new_[21757]_  = ~A299 & \new_[21756]_ ;
  assign \new_[21758]_  = \new_[21757]_  & \new_[21752]_ ;
  assign \new_[21761]_  = ~A167 & ~A169;
  assign \new_[21765]_  = A200 & ~A199;
  assign \new_[21766]_  = ~A166 & \new_[21765]_ ;
  assign \new_[21767]_  = \new_[21766]_  & \new_[21761]_ ;
  assign \new_[21771]_  = A265 & A233;
  assign \new_[21772]_  = ~A232 & \new_[21771]_ ;
  assign \new_[21776]_  = A268 & A267;
  assign \new_[21777]_  = ~A266 & \new_[21776]_ ;
  assign \new_[21778]_  = \new_[21777]_  & \new_[21772]_ ;
  assign \new_[21781]_  = ~A167 & ~A169;
  assign \new_[21785]_  = A200 & ~A199;
  assign \new_[21786]_  = ~A166 & \new_[21785]_ ;
  assign \new_[21787]_  = \new_[21786]_  & \new_[21781]_ ;
  assign \new_[21791]_  = A265 & A233;
  assign \new_[21792]_  = ~A232 & \new_[21791]_ ;
  assign \new_[21796]_  = A269 & A267;
  assign \new_[21797]_  = ~A266 & \new_[21796]_ ;
  assign \new_[21798]_  = \new_[21797]_  & \new_[21792]_ ;
  assign \new_[21801]_  = ~A167 & ~A169;
  assign \new_[21805]_  = A200 & ~A199;
  assign \new_[21806]_  = ~A166 & \new_[21805]_ ;
  assign \new_[21807]_  = \new_[21806]_  & \new_[21801]_ ;
  assign \new_[21811]_  = A265 & ~A234;
  assign \new_[21812]_  = ~A233 & \new_[21811]_ ;
  assign \new_[21816]_  = ~A300 & A298;
  assign \new_[21817]_  = A266 & \new_[21816]_ ;
  assign \new_[21818]_  = \new_[21817]_  & \new_[21812]_ ;
  assign \new_[21821]_  = ~A167 & ~A169;
  assign \new_[21825]_  = A200 & ~A199;
  assign \new_[21826]_  = ~A166 & \new_[21825]_ ;
  assign \new_[21827]_  = \new_[21826]_  & \new_[21821]_ ;
  assign \new_[21831]_  = A265 & ~A234;
  assign \new_[21832]_  = ~A233 & \new_[21831]_ ;
  assign \new_[21836]_  = A299 & A298;
  assign \new_[21837]_  = A266 & \new_[21836]_ ;
  assign \new_[21838]_  = \new_[21837]_  & \new_[21832]_ ;
  assign \new_[21841]_  = ~A167 & ~A169;
  assign \new_[21845]_  = A200 & ~A199;
  assign \new_[21846]_  = ~A166 & \new_[21845]_ ;
  assign \new_[21847]_  = \new_[21846]_  & \new_[21841]_ ;
  assign \new_[21851]_  = A265 & ~A234;
  assign \new_[21852]_  = ~A233 & \new_[21851]_ ;
  assign \new_[21856]_  = ~A299 & ~A298;
  assign \new_[21857]_  = A266 & \new_[21856]_ ;
  assign \new_[21858]_  = \new_[21857]_  & \new_[21852]_ ;
  assign \new_[21861]_  = ~A167 & ~A169;
  assign \new_[21865]_  = A200 & ~A199;
  assign \new_[21866]_  = ~A166 & \new_[21865]_ ;
  assign \new_[21867]_  = \new_[21866]_  & \new_[21861]_ ;
  assign \new_[21871]_  = ~A266 & ~A234;
  assign \new_[21872]_  = ~A233 & \new_[21871]_ ;
  assign \new_[21876]_  = ~A300 & A298;
  assign \new_[21877]_  = ~A267 & \new_[21876]_ ;
  assign \new_[21878]_  = \new_[21877]_  & \new_[21872]_ ;
  assign \new_[21881]_  = ~A167 & ~A169;
  assign \new_[21885]_  = A200 & ~A199;
  assign \new_[21886]_  = ~A166 & \new_[21885]_ ;
  assign \new_[21887]_  = \new_[21886]_  & \new_[21881]_ ;
  assign \new_[21891]_  = ~A266 & ~A234;
  assign \new_[21892]_  = ~A233 & \new_[21891]_ ;
  assign \new_[21896]_  = A299 & A298;
  assign \new_[21897]_  = ~A267 & \new_[21896]_ ;
  assign \new_[21898]_  = \new_[21897]_  & \new_[21892]_ ;
  assign \new_[21901]_  = ~A167 & ~A169;
  assign \new_[21905]_  = A200 & ~A199;
  assign \new_[21906]_  = ~A166 & \new_[21905]_ ;
  assign \new_[21907]_  = \new_[21906]_  & \new_[21901]_ ;
  assign \new_[21911]_  = ~A266 & ~A234;
  assign \new_[21912]_  = ~A233 & \new_[21911]_ ;
  assign \new_[21916]_  = ~A299 & ~A298;
  assign \new_[21917]_  = ~A267 & \new_[21916]_ ;
  assign \new_[21918]_  = \new_[21917]_  & \new_[21912]_ ;
  assign \new_[21921]_  = ~A167 & ~A169;
  assign \new_[21925]_  = A200 & ~A199;
  assign \new_[21926]_  = ~A166 & \new_[21925]_ ;
  assign \new_[21927]_  = \new_[21926]_  & \new_[21921]_ ;
  assign \new_[21931]_  = ~A265 & ~A234;
  assign \new_[21932]_  = ~A233 & \new_[21931]_ ;
  assign \new_[21936]_  = ~A300 & A298;
  assign \new_[21937]_  = ~A266 & \new_[21936]_ ;
  assign \new_[21938]_  = \new_[21937]_  & \new_[21932]_ ;
  assign \new_[21941]_  = ~A167 & ~A169;
  assign \new_[21945]_  = A200 & ~A199;
  assign \new_[21946]_  = ~A166 & \new_[21945]_ ;
  assign \new_[21947]_  = \new_[21946]_  & \new_[21941]_ ;
  assign \new_[21951]_  = ~A265 & ~A234;
  assign \new_[21952]_  = ~A233 & \new_[21951]_ ;
  assign \new_[21956]_  = A299 & A298;
  assign \new_[21957]_  = ~A266 & \new_[21956]_ ;
  assign \new_[21958]_  = \new_[21957]_  & \new_[21952]_ ;
  assign \new_[21961]_  = ~A167 & ~A169;
  assign \new_[21965]_  = A200 & ~A199;
  assign \new_[21966]_  = ~A166 & \new_[21965]_ ;
  assign \new_[21967]_  = \new_[21966]_  & \new_[21961]_ ;
  assign \new_[21971]_  = ~A265 & ~A234;
  assign \new_[21972]_  = ~A233 & \new_[21971]_ ;
  assign \new_[21976]_  = ~A299 & ~A298;
  assign \new_[21977]_  = ~A266 & \new_[21976]_ ;
  assign \new_[21978]_  = \new_[21977]_  & \new_[21972]_ ;
  assign \new_[21981]_  = ~A167 & ~A169;
  assign \new_[21985]_  = A200 & ~A199;
  assign \new_[21986]_  = ~A166 & \new_[21985]_ ;
  assign \new_[21987]_  = \new_[21986]_  & \new_[21981]_ ;
  assign \new_[21991]_  = A234 & ~A233;
  assign \new_[21992]_  = A232 & \new_[21991]_ ;
  assign \new_[21996]_  = A299 & ~A298;
  assign \new_[21997]_  = A235 & \new_[21996]_ ;
  assign \new_[21998]_  = \new_[21997]_  & \new_[21992]_ ;
  assign \new_[22001]_  = ~A167 & ~A169;
  assign \new_[22005]_  = A200 & ~A199;
  assign \new_[22006]_  = ~A166 & \new_[22005]_ ;
  assign \new_[22007]_  = \new_[22006]_  & \new_[22001]_ ;
  assign \new_[22011]_  = A234 & ~A233;
  assign \new_[22012]_  = A232 & \new_[22011]_ ;
  assign \new_[22016]_  = A266 & ~A265;
  assign \new_[22017]_  = A235 & \new_[22016]_ ;
  assign \new_[22018]_  = \new_[22017]_  & \new_[22012]_ ;
  assign \new_[22021]_  = ~A167 & ~A169;
  assign \new_[22025]_  = A200 & ~A199;
  assign \new_[22026]_  = ~A166 & \new_[22025]_ ;
  assign \new_[22027]_  = \new_[22026]_  & \new_[22021]_ ;
  assign \new_[22031]_  = A234 & ~A233;
  assign \new_[22032]_  = A232 & \new_[22031]_ ;
  assign \new_[22036]_  = A299 & ~A298;
  assign \new_[22037]_  = A236 & \new_[22036]_ ;
  assign \new_[22038]_  = \new_[22037]_  & \new_[22032]_ ;
  assign \new_[22041]_  = ~A167 & ~A169;
  assign \new_[22045]_  = A200 & ~A199;
  assign \new_[22046]_  = ~A166 & \new_[22045]_ ;
  assign \new_[22047]_  = \new_[22046]_  & \new_[22041]_ ;
  assign \new_[22051]_  = A234 & ~A233;
  assign \new_[22052]_  = A232 & \new_[22051]_ ;
  assign \new_[22056]_  = A266 & ~A265;
  assign \new_[22057]_  = A236 & \new_[22056]_ ;
  assign \new_[22058]_  = \new_[22057]_  & \new_[22052]_ ;
  assign \new_[22061]_  = ~A167 & ~A169;
  assign \new_[22065]_  = A200 & ~A199;
  assign \new_[22066]_  = ~A166 & \new_[22065]_ ;
  assign \new_[22067]_  = \new_[22066]_  & \new_[22061]_ ;
  assign \new_[22071]_  = A265 & ~A233;
  assign \new_[22072]_  = ~A232 & \new_[22071]_ ;
  assign \new_[22076]_  = ~A300 & A298;
  assign \new_[22077]_  = A266 & \new_[22076]_ ;
  assign \new_[22078]_  = \new_[22077]_  & \new_[22072]_ ;
  assign \new_[22081]_  = ~A167 & ~A169;
  assign \new_[22085]_  = A200 & ~A199;
  assign \new_[22086]_  = ~A166 & \new_[22085]_ ;
  assign \new_[22087]_  = \new_[22086]_  & \new_[22081]_ ;
  assign \new_[22091]_  = A265 & ~A233;
  assign \new_[22092]_  = ~A232 & \new_[22091]_ ;
  assign \new_[22096]_  = A299 & A298;
  assign \new_[22097]_  = A266 & \new_[22096]_ ;
  assign \new_[22098]_  = \new_[22097]_  & \new_[22092]_ ;
  assign \new_[22101]_  = ~A167 & ~A169;
  assign \new_[22105]_  = A200 & ~A199;
  assign \new_[22106]_  = ~A166 & \new_[22105]_ ;
  assign \new_[22107]_  = \new_[22106]_  & \new_[22101]_ ;
  assign \new_[22111]_  = A265 & ~A233;
  assign \new_[22112]_  = ~A232 & \new_[22111]_ ;
  assign \new_[22116]_  = ~A299 & ~A298;
  assign \new_[22117]_  = A266 & \new_[22116]_ ;
  assign \new_[22118]_  = \new_[22117]_  & \new_[22112]_ ;
  assign \new_[22121]_  = ~A167 & ~A169;
  assign \new_[22125]_  = A200 & ~A199;
  assign \new_[22126]_  = ~A166 & \new_[22125]_ ;
  assign \new_[22127]_  = \new_[22126]_  & \new_[22121]_ ;
  assign \new_[22131]_  = ~A266 & ~A233;
  assign \new_[22132]_  = ~A232 & \new_[22131]_ ;
  assign \new_[22136]_  = ~A300 & A298;
  assign \new_[22137]_  = ~A267 & \new_[22136]_ ;
  assign \new_[22138]_  = \new_[22137]_  & \new_[22132]_ ;
  assign \new_[22141]_  = ~A167 & ~A169;
  assign \new_[22145]_  = A200 & ~A199;
  assign \new_[22146]_  = ~A166 & \new_[22145]_ ;
  assign \new_[22147]_  = \new_[22146]_  & \new_[22141]_ ;
  assign \new_[22151]_  = ~A266 & ~A233;
  assign \new_[22152]_  = ~A232 & \new_[22151]_ ;
  assign \new_[22156]_  = A299 & A298;
  assign \new_[22157]_  = ~A267 & \new_[22156]_ ;
  assign \new_[22158]_  = \new_[22157]_  & \new_[22152]_ ;
  assign \new_[22161]_  = ~A167 & ~A169;
  assign \new_[22165]_  = A200 & ~A199;
  assign \new_[22166]_  = ~A166 & \new_[22165]_ ;
  assign \new_[22167]_  = \new_[22166]_  & \new_[22161]_ ;
  assign \new_[22171]_  = ~A266 & ~A233;
  assign \new_[22172]_  = ~A232 & \new_[22171]_ ;
  assign \new_[22176]_  = ~A299 & ~A298;
  assign \new_[22177]_  = ~A267 & \new_[22176]_ ;
  assign \new_[22178]_  = \new_[22177]_  & \new_[22172]_ ;
  assign \new_[22181]_  = ~A167 & ~A169;
  assign \new_[22185]_  = A200 & ~A199;
  assign \new_[22186]_  = ~A166 & \new_[22185]_ ;
  assign \new_[22187]_  = \new_[22186]_  & \new_[22181]_ ;
  assign \new_[22191]_  = ~A265 & ~A233;
  assign \new_[22192]_  = ~A232 & \new_[22191]_ ;
  assign \new_[22196]_  = ~A300 & A298;
  assign \new_[22197]_  = ~A266 & \new_[22196]_ ;
  assign \new_[22198]_  = \new_[22197]_  & \new_[22192]_ ;
  assign \new_[22201]_  = ~A167 & ~A169;
  assign \new_[22205]_  = A200 & ~A199;
  assign \new_[22206]_  = ~A166 & \new_[22205]_ ;
  assign \new_[22207]_  = \new_[22206]_  & \new_[22201]_ ;
  assign \new_[22211]_  = ~A265 & ~A233;
  assign \new_[22212]_  = ~A232 & \new_[22211]_ ;
  assign \new_[22216]_  = A299 & A298;
  assign \new_[22217]_  = ~A266 & \new_[22216]_ ;
  assign \new_[22218]_  = \new_[22217]_  & \new_[22212]_ ;
  assign \new_[22221]_  = ~A167 & ~A169;
  assign \new_[22225]_  = A200 & ~A199;
  assign \new_[22226]_  = ~A166 & \new_[22225]_ ;
  assign \new_[22227]_  = \new_[22226]_  & \new_[22221]_ ;
  assign \new_[22231]_  = ~A265 & ~A233;
  assign \new_[22232]_  = ~A232 & \new_[22231]_ ;
  assign \new_[22236]_  = ~A299 & ~A298;
  assign \new_[22237]_  = ~A266 & \new_[22236]_ ;
  assign \new_[22238]_  = \new_[22237]_  & \new_[22232]_ ;
  assign \new_[22241]_  = ~A167 & ~A169;
  assign \new_[22245]_  = ~A200 & A199;
  assign \new_[22246]_  = ~A166 & \new_[22245]_ ;
  assign \new_[22247]_  = \new_[22246]_  & \new_[22241]_ ;
  assign \new_[22251]_  = ~A232 & A202;
  assign \new_[22252]_  = A201 & \new_[22251]_ ;
  assign \new_[22256]_  = A299 & ~A298;
  assign \new_[22257]_  = A233 & \new_[22256]_ ;
  assign \new_[22258]_  = \new_[22257]_  & \new_[22252]_ ;
  assign \new_[22261]_  = ~A167 & ~A169;
  assign \new_[22265]_  = ~A200 & A199;
  assign \new_[22266]_  = ~A166 & \new_[22265]_ ;
  assign \new_[22267]_  = \new_[22266]_  & \new_[22261]_ ;
  assign \new_[22271]_  = ~A232 & A202;
  assign \new_[22272]_  = A201 & \new_[22271]_ ;
  assign \new_[22276]_  = A266 & ~A265;
  assign \new_[22277]_  = A233 & \new_[22276]_ ;
  assign \new_[22278]_  = \new_[22277]_  & \new_[22272]_ ;
  assign \new_[22281]_  = ~A167 & ~A169;
  assign \new_[22285]_  = ~A200 & A199;
  assign \new_[22286]_  = ~A166 & \new_[22285]_ ;
  assign \new_[22287]_  = \new_[22286]_  & \new_[22281]_ ;
  assign \new_[22291]_  = ~A232 & A203;
  assign \new_[22292]_  = A201 & \new_[22291]_ ;
  assign \new_[22296]_  = A299 & ~A298;
  assign \new_[22297]_  = A233 & \new_[22296]_ ;
  assign \new_[22298]_  = \new_[22297]_  & \new_[22292]_ ;
  assign \new_[22301]_  = ~A167 & ~A169;
  assign \new_[22305]_  = ~A200 & A199;
  assign \new_[22306]_  = ~A166 & \new_[22305]_ ;
  assign \new_[22307]_  = \new_[22306]_  & \new_[22301]_ ;
  assign \new_[22311]_  = ~A232 & A203;
  assign \new_[22312]_  = A201 & \new_[22311]_ ;
  assign \new_[22316]_  = A266 & ~A265;
  assign \new_[22317]_  = A233 & \new_[22316]_ ;
  assign \new_[22318]_  = \new_[22317]_  & \new_[22312]_ ;
  assign \new_[22321]_  = ~A169 & A170;
  assign \new_[22325]_  = ~A200 & ~A166;
  assign \new_[22326]_  = A167 & \new_[22325]_ ;
  assign \new_[22327]_  = \new_[22326]_  & \new_[22321]_ ;
  assign \new_[22331]_  = ~A232 & ~A203;
  assign \new_[22332]_  = ~A202 & \new_[22331]_ ;
  assign \new_[22336]_  = A299 & ~A298;
  assign \new_[22337]_  = A233 & \new_[22336]_ ;
  assign \new_[22338]_  = \new_[22337]_  & \new_[22332]_ ;
  assign \new_[22341]_  = ~A169 & A170;
  assign \new_[22345]_  = ~A200 & ~A166;
  assign \new_[22346]_  = A167 & \new_[22345]_ ;
  assign \new_[22347]_  = \new_[22346]_  & \new_[22341]_ ;
  assign \new_[22351]_  = ~A232 & ~A203;
  assign \new_[22352]_  = ~A202 & \new_[22351]_ ;
  assign \new_[22356]_  = A266 & ~A265;
  assign \new_[22357]_  = A233 & \new_[22356]_ ;
  assign \new_[22358]_  = \new_[22357]_  & \new_[22352]_ ;
  assign \new_[22361]_  = ~A169 & A170;
  assign \new_[22365]_  = ~A200 & A166;
  assign \new_[22366]_  = ~A167 & \new_[22365]_ ;
  assign \new_[22367]_  = \new_[22366]_  & \new_[22361]_ ;
  assign \new_[22371]_  = ~A232 & ~A203;
  assign \new_[22372]_  = ~A202 & \new_[22371]_ ;
  assign \new_[22376]_  = A299 & ~A298;
  assign \new_[22377]_  = A233 & \new_[22376]_ ;
  assign \new_[22378]_  = \new_[22377]_  & \new_[22372]_ ;
  assign \new_[22381]_  = ~A169 & A170;
  assign \new_[22385]_  = ~A200 & A166;
  assign \new_[22386]_  = ~A167 & \new_[22385]_ ;
  assign \new_[22387]_  = \new_[22386]_  & \new_[22381]_ ;
  assign \new_[22391]_  = ~A232 & ~A203;
  assign \new_[22392]_  = ~A202 & \new_[22391]_ ;
  assign \new_[22396]_  = A266 & ~A265;
  assign \new_[22397]_  = A233 & \new_[22396]_ ;
  assign \new_[22398]_  = \new_[22397]_  & \new_[22392]_ ;
  assign \new_[22401]_  = ~A169 & ~A170;
  assign \new_[22405]_  = ~A200 & A199;
  assign \new_[22406]_  = ~A168 & \new_[22405]_ ;
  assign \new_[22407]_  = \new_[22406]_  & \new_[22401]_ ;
  assign \new_[22411]_  = ~A232 & A202;
  assign \new_[22412]_  = A201 & \new_[22411]_ ;
  assign \new_[22416]_  = A299 & ~A298;
  assign \new_[22417]_  = A233 & \new_[22416]_ ;
  assign \new_[22418]_  = \new_[22417]_  & \new_[22412]_ ;
  assign \new_[22421]_  = ~A169 & ~A170;
  assign \new_[22425]_  = ~A200 & A199;
  assign \new_[22426]_  = ~A168 & \new_[22425]_ ;
  assign \new_[22427]_  = \new_[22426]_  & \new_[22421]_ ;
  assign \new_[22431]_  = ~A232 & A202;
  assign \new_[22432]_  = A201 & \new_[22431]_ ;
  assign \new_[22436]_  = A266 & ~A265;
  assign \new_[22437]_  = A233 & \new_[22436]_ ;
  assign \new_[22438]_  = \new_[22437]_  & \new_[22432]_ ;
  assign \new_[22441]_  = ~A169 & ~A170;
  assign \new_[22445]_  = ~A200 & A199;
  assign \new_[22446]_  = ~A168 & \new_[22445]_ ;
  assign \new_[22447]_  = \new_[22446]_  & \new_[22441]_ ;
  assign \new_[22451]_  = ~A232 & A203;
  assign \new_[22452]_  = A201 & \new_[22451]_ ;
  assign \new_[22456]_  = A299 & ~A298;
  assign \new_[22457]_  = A233 & \new_[22456]_ ;
  assign \new_[22458]_  = \new_[22457]_  & \new_[22452]_ ;
  assign \new_[22461]_  = ~A169 & ~A170;
  assign \new_[22465]_  = ~A200 & A199;
  assign \new_[22466]_  = ~A168 & \new_[22465]_ ;
  assign \new_[22467]_  = \new_[22466]_  & \new_[22461]_ ;
  assign \new_[22471]_  = ~A232 & A203;
  assign \new_[22472]_  = A201 & \new_[22471]_ ;
  assign \new_[22476]_  = A266 & ~A265;
  assign \new_[22477]_  = A233 & \new_[22476]_ ;
  assign \new_[22478]_  = \new_[22477]_  & \new_[22472]_ ;
  assign \new_[22482]_  = A199 & A166;
  assign \new_[22483]_  = A168 & \new_[22482]_ ;
  assign \new_[22487]_  = A233 & A232;
  assign \new_[22488]_  = A200 & \new_[22487]_ ;
  assign \new_[22489]_  = \new_[22488]_  & \new_[22483]_ ;
  assign \new_[22493]_  = ~A269 & ~A268;
  assign \new_[22494]_  = A265 & \new_[22493]_ ;
  assign \new_[22498]_  = ~A302 & ~A301;
  assign \new_[22499]_  = ~A299 & \new_[22498]_ ;
  assign \new_[22500]_  = \new_[22499]_  & \new_[22494]_ ;
  assign \new_[22504]_  = A199 & A166;
  assign \new_[22505]_  = A168 & \new_[22504]_ ;
  assign \new_[22509]_  = ~A235 & ~A233;
  assign \new_[22510]_  = A200 & \new_[22509]_ ;
  assign \new_[22511]_  = \new_[22510]_  & \new_[22505]_ ;
  assign \new_[22515]_  = A266 & A265;
  assign \new_[22516]_  = ~A236 & \new_[22515]_ ;
  assign \new_[22520]_  = ~A302 & ~A301;
  assign \new_[22521]_  = A298 & \new_[22520]_ ;
  assign \new_[22522]_  = \new_[22521]_  & \new_[22516]_ ;
  assign \new_[22526]_  = A199 & A166;
  assign \new_[22527]_  = A168 & \new_[22526]_ ;
  assign \new_[22531]_  = ~A235 & ~A233;
  assign \new_[22532]_  = A200 & \new_[22531]_ ;
  assign \new_[22533]_  = \new_[22532]_  & \new_[22527]_ ;
  assign \new_[22537]_  = ~A268 & ~A266;
  assign \new_[22538]_  = ~A236 & \new_[22537]_ ;
  assign \new_[22542]_  = ~A300 & A298;
  assign \new_[22543]_  = ~A269 & \new_[22542]_ ;
  assign \new_[22544]_  = \new_[22543]_  & \new_[22538]_ ;
  assign \new_[22548]_  = A199 & A166;
  assign \new_[22549]_  = A168 & \new_[22548]_ ;
  assign \new_[22553]_  = ~A235 & ~A233;
  assign \new_[22554]_  = A200 & \new_[22553]_ ;
  assign \new_[22555]_  = \new_[22554]_  & \new_[22549]_ ;
  assign \new_[22559]_  = ~A268 & ~A266;
  assign \new_[22560]_  = ~A236 & \new_[22559]_ ;
  assign \new_[22564]_  = A299 & A298;
  assign \new_[22565]_  = ~A269 & \new_[22564]_ ;
  assign \new_[22566]_  = \new_[22565]_  & \new_[22560]_ ;
  assign \new_[22570]_  = A199 & A166;
  assign \new_[22571]_  = A168 & \new_[22570]_ ;
  assign \new_[22575]_  = ~A235 & ~A233;
  assign \new_[22576]_  = A200 & \new_[22575]_ ;
  assign \new_[22577]_  = \new_[22576]_  & \new_[22571]_ ;
  assign \new_[22581]_  = ~A268 & ~A266;
  assign \new_[22582]_  = ~A236 & \new_[22581]_ ;
  assign \new_[22586]_  = ~A299 & ~A298;
  assign \new_[22587]_  = ~A269 & \new_[22586]_ ;
  assign \new_[22588]_  = \new_[22587]_  & \new_[22582]_ ;
  assign \new_[22592]_  = A199 & A166;
  assign \new_[22593]_  = A168 & \new_[22592]_ ;
  assign \new_[22597]_  = ~A235 & ~A233;
  assign \new_[22598]_  = A200 & \new_[22597]_ ;
  assign \new_[22599]_  = \new_[22598]_  & \new_[22593]_ ;
  assign \new_[22603]_  = ~A267 & ~A266;
  assign \new_[22604]_  = ~A236 & \new_[22603]_ ;
  assign \new_[22608]_  = ~A302 & ~A301;
  assign \new_[22609]_  = A298 & \new_[22608]_ ;
  assign \new_[22610]_  = \new_[22609]_  & \new_[22604]_ ;
  assign \new_[22614]_  = A199 & A166;
  assign \new_[22615]_  = A168 & \new_[22614]_ ;
  assign \new_[22619]_  = ~A235 & ~A233;
  assign \new_[22620]_  = A200 & \new_[22619]_ ;
  assign \new_[22621]_  = \new_[22620]_  & \new_[22615]_ ;
  assign \new_[22625]_  = ~A266 & ~A265;
  assign \new_[22626]_  = ~A236 & \new_[22625]_ ;
  assign \new_[22630]_  = ~A302 & ~A301;
  assign \new_[22631]_  = A298 & \new_[22630]_ ;
  assign \new_[22632]_  = \new_[22631]_  & \new_[22626]_ ;
  assign \new_[22636]_  = A199 & A166;
  assign \new_[22637]_  = A168 & \new_[22636]_ ;
  assign \new_[22641]_  = ~A234 & ~A233;
  assign \new_[22642]_  = A200 & \new_[22641]_ ;
  assign \new_[22643]_  = \new_[22642]_  & \new_[22637]_ ;
  assign \new_[22647]_  = ~A269 & ~A268;
  assign \new_[22648]_  = ~A266 & \new_[22647]_ ;
  assign \new_[22652]_  = ~A302 & ~A301;
  assign \new_[22653]_  = A298 & \new_[22652]_ ;
  assign \new_[22654]_  = \new_[22653]_  & \new_[22648]_ ;
  assign \new_[22658]_  = A199 & A166;
  assign \new_[22659]_  = A168 & \new_[22658]_ ;
  assign \new_[22663]_  = ~A233 & A232;
  assign \new_[22664]_  = A200 & \new_[22663]_ ;
  assign \new_[22665]_  = \new_[22664]_  & \new_[22659]_ ;
  assign \new_[22669]_  = A298 & A235;
  assign \new_[22670]_  = A234 & \new_[22669]_ ;
  assign \new_[22674]_  = A301 & A300;
  assign \new_[22675]_  = ~A299 & \new_[22674]_ ;
  assign \new_[22676]_  = \new_[22675]_  & \new_[22670]_ ;
  assign \new_[22680]_  = A199 & A166;
  assign \new_[22681]_  = A168 & \new_[22680]_ ;
  assign \new_[22685]_  = ~A233 & A232;
  assign \new_[22686]_  = A200 & \new_[22685]_ ;
  assign \new_[22687]_  = \new_[22686]_  & \new_[22681]_ ;
  assign \new_[22691]_  = A298 & A235;
  assign \new_[22692]_  = A234 & \new_[22691]_ ;
  assign \new_[22696]_  = A302 & A300;
  assign \new_[22697]_  = ~A299 & \new_[22696]_ ;
  assign \new_[22698]_  = \new_[22697]_  & \new_[22692]_ ;
  assign \new_[22702]_  = A199 & A166;
  assign \new_[22703]_  = A168 & \new_[22702]_ ;
  assign \new_[22707]_  = ~A233 & A232;
  assign \new_[22708]_  = A200 & \new_[22707]_ ;
  assign \new_[22709]_  = \new_[22708]_  & \new_[22703]_ ;
  assign \new_[22713]_  = A265 & A235;
  assign \new_[22714]_  = A234 & \new_[22713]_ ;
  assign \new_[22718]_  = A268 & A267;
  assign \new_[22719]_  = ~A266 & \new_[22718]_ ;
  assign \new_[22720]_  = \new_[22719]_  & \new_[22714]_ ;
  assign \new_[22724]_  = A199 & A166;
  assign \new_[22725]_  = A168 & \new_[22724]_ ;
  assign \new_[22729]_  = ~A233 & A232;
  assign \new_[22730]_  = A200 & \new_[22729]_ ;
  assign \new_[22731]_  = \new_[22730]_  & \new_[22725]_ ;
  assign \new_[22735]_  = A265 & A235;
  assign \new_[22736]_  = A234 & \new_[22735]_ ;
  assign \new_[22740]_  = A269 & A267;
  assign \new_[22741]_  = ~A266 & \new_[22740]_ ;
  assign \new_[22742]_  = \new_[22741]_  & \new_[22736]_ ;
  assign \new_[22746]_  = A199 & A166;
  assign \new_[22747]_  = A168 & \new_[22746]_ ;
  assign \new_[22751]_  = ~A233 & A232;
  assign \new_[22752]_  = A200 & \new_[22751]_ ;
  assign \new_[22753]_  = \new_[22752]_  & \new_[22747]_ ;
  assign \new_[22757]_  = A298 & A236;
  assign \new_[22758]_  = A234 & \new_[22757]_ ;
  assign \new_[22762]_  = A301 & A300;
  assign \new_[22763]_  = ~A299 & \new_[22762]_ ;
  assign \new_[22764]_  = \new_[22763]_  & \new_[22758]_ ;
  assign \new_[22768]_  = A199 & A166;
  assign \new_[22769]_  = A168 & \new_[22768]_ ;
  assign \new_[22773]_  = ~A233 & A232;
  assign \new_[22774]_  = A200 & \new_[22773]_ ;
  assign \new_[22775]_  = \new_[22774]_  & \new_[22769]_ ;
  assign \new_[22779]_  = A298 & A236;
  assign \new_[22780]_  = A234 & \new_[22779]_ ;
  assign \new_[22784]_  = A302 & A300;
  assign \new_[22785]_  = ~A299 & \new_[22784]_ ;
  assign \new_[22786]_  = \new_[22785]_  & \new_[22780]_ ;
  assign \new_[22790]_  = A199 & A166;
  assign \new_[22791]_  = A168 & \new_[22790]_ ;
  assign \new_[22795]_  = ~A233 & A232;
  assign \new_[22796]_  = A200 & \new_[22795]_ ;
  assign \new_[22797]_  = \new_[22796]_  & \new_[22791]_ ;
  assign \new_[22801]_  = A265 & A236;
  assign \new_[22802]_  = A234 & \new_[22801]_ ;
  assign \new_[22806]_  = A268 & A267;
  assign \new_[22807]_  = ~A266 & \new_[22806]_ ;
  assign \new_[22808]_  = \new_[22807]_  & \new_[22802]_ ;
  assign \new_[22812]_  = A199 & A166;
  assign \new_[22813]_  = A168 & \new_[22812]_ ;
  assign \new_[22817]_  = ~A233 & A232;
  assign \new_[22818]_  = A200 & \new_[22817]_ ;
  assign \new_[22819]_  = \new_[22818]_  & \new_[22813]_ ;
  assign \new_[22823]_  = A265 & A236;
  assign \new_[22824]_  = A234 & \new_[22823]_ ;
  assign \new_[22828]_  = A269 & A267;
  assign \new_[22829]_  = ~A266 & \new_[22828]_ ;
  assign \new_[22830]_  = \new_[22829]_  & \new_[22824]_ ;
  assign \new_[22834]_  = A199 & A166;
  assign \new_[22835]_  = A168 & \new_[22834]_ ;
  assign \new_[22839]_  = ~A233 & ~A232;
  assign \new_[22840]_  = A200 & \new_[22839]_ ;
  assign \new_[22841]_  = \new_[22840]_  & \new_[22835]_ ;
  assign \new_[22845]_  = ~A269 & ~A268;
  assign \new_[22846]_  = ~A266 & \new_[22845]_ ;
  assign \new_[22850]_  = ~A302 & ~A301;
  assign \new_[22851]_  = A298 & \new_[22850]_ ;
  assign \new_[22852]_  = \new_[22851]_  & \new_[22846]_ ;
  assign \new_[22856]_  = ~A200 & A166;
  assign \new_[22857]_  = A168 & \new_[22856]_ ;
  assign \new_[22861]_  = A232 & ~A203;
  assign \new_[22862]_  = ~A202 & \new_[22861]_ ;
  assign \new_[22863]_  = \new_[22862]_  & \new_[22857]_ ;
  assign \new_[22867]_  = ~A268 & A265;
  assign \new_[22868]_  = A233 & \new_[22867]_ ;
  assign \new_[22872]_  = ~A300 & ~A299;
  assign \new_[22873]_  = ~A269 & \new_[22872]_ ;
  assign \new_[22874]_  = \new_[22873]_  & \new_[22868]_ ;
  assign \new_[22878]_  = ~A200 & A166;
  assign \new_[22879]_  = A168 & \new_[22878]_ ;
  assign \new_[22883]_  = A232 & ~A203;
  assign \new_[22884]_  = ~A202 & \new_[22883]_ ;
  assign \new_[22885]_  = \new_[22884]_  & \new_[22879]_ ;
  assign \new_[22889]_  = ~A268 & A265;
  assign \new_[22890]_  = A233 & \new_[22889]_ ;
  assign \new_[22894]_  = A299 & A298;
  assign \new_[22895]_  = ~A269 & \new_[22894]_ ;
  assign \new_[22896]_  = \new_[22895]_  & \new_[22890]_ ;
  assign \new_[22900]_  = ~A200 & A166;
  assign \new_[22901]_  = A168 & \new_[22900]_ ;
  assign \new_[22905]_  = A232 & ~A203;
  assign \new_[22906]_  = ~A202 & \new_[22905]_ ;
  assign \new_[22907]_  = \new_[22906]_  & \new_[22901]_ ;
  assign \new_[22911]_  = ~A268 & A265;
  assign \new_[22912]_  = A233 & \new_[22911]_ ;
  assign \new_[22916]_  = ~A299 & ~A298;
  assign \new_[22917]_  = ~A269 & \new_[22916]_ ;
  assign \new_[22918]_  = \new_[22917]_  & \new_[22912]_ ;
  assign \new_[22922]_  = ~A200 & A166;
  assign \new_[22923]_  = A168 & \new_[22922]_ ;
  assign \new_[22927]_  = A232 & ~A203;
  assign \new_[22928]_  = ~A202 & \new_[22927]_ ;
  assign \new_[22929]_  = \new_[22928]_  & \new_[22923]_ ;
  assign \new_[22933]_  = ~A267 & A265;
  assign \new_[22934]_  = A233 & \new_[22933]_ ;
  assign \new_[22938]_  = ~A302 & ~A301;
  assign \new_[22939]_  = ~A299 & \new_[22938]_ ;
  assign \new_[22940]_  = \new_[22939]_  & \new_[22934]_ ;
  assign \new_[22944]_  = ~A200 & A166;
  assign \new_[22945]_  = A168 & \new_[22944]_ ;
  assign \new_[22949]_  = A232 & ~A203;
  assign \new_[22950]_  = ~A202 & \new_[22949]_ ;
  assign \new_[22951]_  = \new_[22950]_  & \new_[22945]_ ;
  assign \new_[22955]_  = A266 & A265;
  assign \new_[22956]_  = A233 & \new_[22955]_ ;
  assign \new_[22960]_  = ~A302 & ~A301;
  assign \new_[22961]_  = ~A299 & \new_[22960]_ ;
  assign \new_[22962]_  = \new_[22961]_  & \new_[22956]_ ;
  assign \new_[22966]_  = ~A200 & A166;
  assign \new_[22967]_  = A168 & \new_[22966]_ ;
  assign \new_[22971]_  = A232 & ~A203;
  assign \new_[22972]_  = ~A202 & \new_[22971]_ ;
  assign \new_[22973]_  = \new_[22972]_  & \new_[22967]_ ;
  assign \new_[22977]_  = ~A266 & ~A265;
  assign \new_[22978]_  = A233 & \new_[22977]_ ;
  assign \new_[22982]_  = ~A302 & ~A301;
  assign \new_[22983]_  = ~A299 & \new_[22982]_ ;
  assign \new_[22984]_  = \new_[22983]_  & \new_[22978]_ ;
  assign \new_[22988]_  = ~A200 & A166;
  assign \new_[22989]_  = A168 & \new_[22988]_ ;
  assign \new_[22993]_  = ~A233 & ~A203;
  assign \new_[22994]_  = ~A202 & \new_[22993]_ ;
  assign \new_[22995]_  = \new_[22994]_  & \new_[22989]_ ;
  assign \new_[22999]_  = A265 & ~A236;
  assign \new_[23000]_  = ~A235 & \new_[22999]_ ;
  assign \new_[23004]_  = ~A300 & A298;
  assign \new_[23005]_  = A266 & \new_[23004]_ ;
  assign \new_[23006]_  = \new_[23005]_  & \new_[23000]_ ;
  assign \new_[23010]_  = ~A200 & A166;
  assign \new_[23011]_  = A168 & \new_[23010]_ ;
  assign \new_[23015]_  = ~A233 & ~A203;
  assign \new_[23016]_  = ~A202 & \new_[23015]_ ;
  assign \new_[23017]_  = \new_[23016]_  & \new_[23011]_ ;
  assign \new_[23021]_  = A265 & ~A236;
  assign \new_[23022]_  = ~A235 & \new_[23021]_ ;
  assign \new_[23026]_  = A299 & A298;
  assign \new_[23027]_  = A266 & \new_[23026]_ ;
  assign \new_[23028]_  = \new_[23027]_  & \new_[23022]_ ;
  assign \new_[23032]_  = ~A200 & A166;
  assign \new_[23033]_  = A168 & \new_[23032]_ ;
  assign \new_[23037]_  = ~A233 & ~A203;
  assign \new_[23038]_  = ~A202 & \new_[23037]_ ;
  assign \new_[23039]_  = \new_[23038]_  & \new_[23033]_ ;
  assign \new_[23043]_  = A265 & ~A236;
  assign \new_[23044]_  = ~A235 & \new_[23043]_ ;
  assign \new_[23048]_  = ~A299 & ~A298;
  assign \new_[23049]_  = A266 & \new_[23048]_ ;
  assign \new_[23050]_  = \new_[23049]_  & \new_[23044]_ ;
  assign \new_[23054]_  = ~A200 & A166;
  assign \new_[23055]_  = A168 & \new_[23054]_ ;
  assign \new_[23059]_  = ~A233 & ~A203;
  assign \new_[23060]_  = ~A202 & \new_[23059]_ ;
  assign \new_[23061]_  = \new_[23060]_  & \new_[23055]_ ;
  assign \new_[23065]_  = ~A266 & ~A236;
  assign \new_[23066]_  = ~A235 & \new_[23065]_ ;
  assign \new_[23070]_  = ~A300 & A298;
  assign \new_[23071]_  = ~A267 & \new_[23070]_ ;
  assign \new_[23072]_  = \new_[23071]_  & \new_[23066]_ ;
  assign \new_[23076]_  = ~A200 & A166;
  assign \new_[23077]_  = A168 & \new_[23076]_ ;
  assign \new_[23081]_  = ~A233 & ~A203;
  assign \new_[23082]_  = ~A202 & \new_[23081]_ ;
  assign \new_[23083]_  = \new_[23082]_  & \new_[23077]_ ;
  assign \new_[23087]_  = ~A266 & ~A236;
  assign \new_[23088]_  = ~A235 & \new_[23087]_ ;
  assign \new_[23092]_  = A299 & A298;
  assign \new_[23093]_  = ~A267 & \new_[23092]_ ;
  assign \new_[23094]_  = \new_[23093]_  & \new_[23088]_ ;
  assign \new_[23098]_  = ~A200 & A166;
  assign \new_[23099]_  = A168 & \new_[23098]_ ;
  assign \new_[23103]_  = ~A233 & ~A203;
  assign \new_[23104]_  = ~A202 & \new_[23103]_ ;
  assign \new_[23105]_  = \new_[23104]_  & \new_[23099]_ ;
  assign \new_[23109]_  = ~A266 & ~A236;
  assign \new_[23110]_  = ~A235 & \new_[23109]_ ;
  assign \new_[23114]_  = ~A299 & ~A298;
  assign \new_[23115]_  = ~A267 & \new_[23114]_ ;
  assign \new_[23116]_  = \new_[23115]_  & \new_[23110]_ ;
  assign \new_[23120]_  = ~A200 & A166;
  assign \new_[23121]_  = A168 & \new_[23120]_ ;
  assign \new_[23125]_  = ~A233 & ~A203;
  assign \new_[23126]_  = ~A202 & \new_[23125]_ ;
  assign \new_[23127]_  = \new_[23126]_  & \new_[23121]_ ;
  assign \new_[23131]_  = ~A265 & ~A236;
  assign \new_[23132]_  = ~A235 & \new_[23131]_ ;
  assign \new_[23136]_  = ~A300 & A298;
  assign \new_[23137]_  = ~A266 & \new_[23136]_ ;
  assign \new_[23138]_  = \new_[23137]_  & \new_[23132]_ ;
  assign \new_[23142]_  = ~A200 & A166;
  assign \new_[23143]_  = A168 & \new_[23142]_ ;
  assign \new_[23147]_  = ~A233 & ~A203;
  assign \new_[23148]_  = ~A202 & \new_[23147]_ ;
  assign \new_[23149]_  = \new_[23148]_  & \new_[23143]_ ;
  assign \new_[23153]_  = ~A265 & ~A236;
  assign \new_[23154]_  = ~A235 & \new_[23153]_ ;
  assign \new_[23158]_  = A299 & A298;
  assign \new_[23159]_  = ~A266 & \new_[23158]_ ;
  assign \new_[23160]_  = \new_[23159]_  & \new_[23154]_ ;
  assign \new_[23164]_  = ~A200 & A166;
  assign \new_[23165]_  = A168 & \new_[23164]_ ;
  assign \new_[23169]_  = ~A233 & ~A203;
  assign \new_[23170]_  = ~A202 & \new_[23169]_ ;
  assign \new_[23171]_  = \new_[23170]_  & \new_[23165]_ ;
  assign \new_[23175]_  = ~A265 & ~A236;
  assign \new_[23176]_  = ~A235 & \new_[23175]_ ;
  assign \new_[23180]_  = ~A299 & ~A298;
  assign \new_[23181]_  = ~A266 & \new_[23180]_ ;
  assign \new_[23182]_  = \new_[23181]_  & \new_[23176]_ ;
  assign \new_[23186]_  = ~A200 & A166;
  assign \new_[23187]_  = A168 & \new_[23186]_ ;
  assign \new_[23191]_  = ~A233 & ~A203;
  assign \new_[23192]_  = ~A202 & \new_[23191]_ ;
  assign \new_[23193]_  = \new_[23192]_  & \new_[23187]_ ;
  assign \new_[23197]_  = A266 & A265;
  assign \new_[23198]_  = ~A234 & \new_[23197]_ ;
  assign \new_[23202]_  = ~A302 & ~A301;
  assign \new_[23203]_  = A298 & \new_[23202]_ ;
  assign \new_[23204]_  = \new_[23203]_  & \new_[23198]_ ;
  assign \new_[23208]_  = ~A200 & A166;
  assign \new_[23209]_  = A168 & \new_[23208]_ ;
  assign \new_[23213]_  = ~A233 & ~A203;
  assign \new_[23214]_  = ~A202 & \new_[23213]_ ;
  assign \new_[23215]_  = \new_[23214]_  & \new_[23209]_ ;
  assign \new_[23219]_  = ~A268 & ~A266;
  assign \new_[23220]_  = ~A234 & \new_[23219]_ ;
  assign \new_[23224]_  = ~A300 & A298;
  assign \new_[23225]_  = ~A269 & \new_[23224]_ ;
  assign \new_[23226]_  = \new_[23225]_  & \new_[23220]_ ;
  assign \new_[23230]_  = ~A200 & A166;
  assign \new_[23231]_  = A168 & \new_[23230]_ ;
  assign \new_[23235]_  = ~A233 & ~A203;
  assign \new_[23236]_  = ~A202 & \new_[23235]_ ;
  assign \new_[23237]_  = \new_[23236]_  & \new_[23231]_ ;
  assign \new_[23241]_  = ~A268 & ~A266;
  assign \new_[23242]_  = ~A234 & \new_[23241]_ ;
  assign \new_[23246]_  = A299 & A298;
  assign \new_[23247]_  = ~A269 & \new_[23246]_ ;
  assign \new_[23248]_  = \new_[23247]_  & \new_[23242]_ ;
  assign \new_[23252]_  = ~A200 & A166;
  assign \new_[23253]_  = A168 & \new_[23252]_ ;
  assign \new_[23257]_  = ~A233 & ~A203;
  assign \new_[23258]_  = ~A202 & \new_[23257]_ ;
  assign \new_[23259]_  = \new_[23258]_  & \new_[23253]_ ;
  assign \new_[23263]_  = ~A268 & ~A266;
  assign \new_[23264]_  = ~A234 & \new_[23263]_ ;
  assign \new_[23268]_  = ~A299 & ~A298;
  assign \new_[23269]_  = ~A269 & \new_[23268]_ ;
  assign \new_[23270]_  = \new_[23269]_  & \new_[23264]_ ;
  assign \new_[23274]_  = ~A200 & A166;
  assign \new_[23275]_  = A168 & \new_[23274]_ ;
  assign \new_[23279]_  = ~A233 & ~A203;
  assign \new_[23280]_  = ~A202 & \new_[23279]_ ;
  assign \new_[23281]_  = \new_[23280]_  & \new_[23275]_ ;
  assign \new_[23285]_  = ~A267 & ~A266;
  assign \new_[23286]_  = ~A234 & \new_[23285]_ ;
  assign \new_[23290]_  = ~A302 & ~A301;
  assign \new_[23291]_  = A298 & \new_[23290]_ ;
  assign \new_[23292]_  = \new_[23291]_  & \new_[23286]_ ;
  assign \new_[23296]_  = ~A200 & A166;
  assign \new_[23297]_  = A168 & \new_[23296]_ ;
  assign \new_[23301]_  = ~A233 & ~A203;
  assign \new_[23302]_  = ~A202 & \new_[23301]_ ;
  assign \new_[23303]_  = \new_[23302]_  & \new_[23297]_ ;
  assign \new_[23307]_  = ~A266 & ~A265;
  assign \new_[23308]_  = ~A234 & \new_[23307]_ ;
  assign \new_[23312]_  = ~A302 & ~A301;
  assign \new_[23313]_  = A298 & \new_[23312]_ ;
  assign \new_[23314]_  = \new_[23313]_  & \new_[23308]_ ;
  assign \new_[23318]_  = ~A200 & A166;
  assign \new_[23319]_  = A168 & \new_[23318]_ ;
  assign \new_[23323]_  = ~A232 & ~A203;
  assign \new_[23324]_  = ~A202 & \new_[23323]_ ;
  assign \new_[23325]_  = \new_[23324]_  & \new_[23319]_ ;
  assign \new_[23329]_  = A266 & A265;
  assign \new_[23330]_  = ~A233 & \new_[23329]_ ;
  assign \new_[23334]_  = ~A302 & ~A301;
  assign \new_[23335]_  = A298 & \new_[23334]_ ;
  assign \new_[23336]_  = \new_[23335]_  & \new_[23330]_ ;
  assign \new_[23340]_  = ~A200 & A166;
  assign \new_[23341]_  = A168 & \new_[23340]_ ;
  assign \new_[23345]_  = ~A232 & ~A203;
  assign \new_[23346]_  = ~A202 & \new_[23345]_ ;
  assign \new_[23347]_  = \new_[23346]_  & \new_[23341]_ ;
  assign \new_[23351]_  = ~A268 & ~A266;
  assign \new_[23352]_  = ~A233 & \new_[23351]_ ;
  assign \new_[23356]_  = ~A300 & A298;
  assign \new_[23357]_  = ~A269 & \new_[23356]_ ;
  assign \new_[23358]_  = \new_[23357]_  & \new_[23352]_ ;
  assign \new_[23362]_  = ~A200 & A166;
  assign \new_[23363]_  = A168 & \new_[23362]_ ;
  assign \new_[23367]_  = ~A232 & ~A203;
  assign \new_[23368]_  = ~A202 & \new_[23367]_ ;
  assign \new_[23369]_  = \new_[23368]_  & \new_[23363]_ ;
  assign \new_[23373]_  = ~A268 & ~A266;
  assign \new_[23374]_  = ~A233 & \new_[23373]_ ;
  assign \new_[23378]_  = A299 & A298;
  assign \new_[23379]_  = ~A269 & \new_[23378]_ ;
  assign \new_[23380]_  = \new_[23379]_  & \new_[23374]_ ;
  assign \new_[23384]_  = ~A200 & A166;
  assign \new_[23385]_  = A168 & \new_[23384]_ ;
  assign \new_[23389]_  = ~A232 & ~A203;
  assign \new_[23390]_  = ~A202 & \new_[23389]_ ;
  assign \new_[23391]_  = \new_[23390]_  & \new_[23385]_ ;
  assign \new_[23395]_  = ~A268 & ~A266;
  assign \new_[23396]_  = ~A233 & \new_[23395]_ ;
  assign \new_[23400]_  = ~A299 & ~A298;
  assign \new_[23401]_  = ~A269 & \new_[23400]_ ;
  assign \new_[23402]_  = \new_[23401]_  & \new_[23396]_ ;
  assign \new_[23406]_  = ~A200 & A166;
  assign \new_[23407]_  = A168 & \new_[23406]_ ;
  assign \new_[23411]_  = ~A232 & ~A203;
  assign \new_[23412]_  = ~A202 & \new_[23411]_ ;
  assign \new_[23413]_  = \new_[23412]_  & \new_[23407]_ ;
  assign \new_[23417]_  = ~A267 & ~A266;
  assign \new_[23418]_  = ~A233 & \new_[23417]_ ;
  assign \new_[23422]_  = ~A302 & ~A301;
  assign \new_[23423]_  = A298 & \new_[23422]_ ;
  assign \new_[23424]_  = \new_[23423]_  & \new_[23418]_ ;
  assign \new_[23428]_  = ~A200 & A166;
  assign \new_[23429]_  = A168 & \new_[23428]_ ;
  assign \new_[23433]_  = ~A232 & ~A203;
  assign \new_[23434]_  = ~A202 & \new_[23433]_ ;
  assign \new_[23435]_  = \new_[23434]_  & \new_[23429]_ ;
  assign \new_[23439]_  = ~A266 & ~A265;
  assign \new_[23440]_  = ~A233 & \new_[23439]_ ;
  assign \new_[23444]_  = ~A302 & ~A301;
  assign \new_[23445]_  = A298 & \new_[23444]_ ;
  assign \new_[23446]_  = \new_[23445]_  & \new_[23440]_ ;
  assign \new_[23450]_  = ~A200 & A166;
  assign \new_[23451]_  = A168 & \new_[23450]_ ;
  assign \new_[23455]_  = A233 & A232;
  assign \new_[23456]_  = ~A201 & \new_[23455]_ ;
  assign \new_[23457]_  = \new_[23456]_  & \new_[23451]_ ;
  assign \new_[23461]_  = ~A269 & ~A268;
  assign \new_[23462]_  = A265 & \new_[23461]_ ;
  assign \new_[23466]_  = ~A302 & ~A301;
  assign \new_[23467]_  = ~A299 & \new_[23466]_ ;
  assign \new_[23468]_  = \new_[23467]_  & \new_[23462]_ ;
  assign \new_[23472]_  = ~A200 & A166;
  assign \new_[23473]_  = A168 & \new_[23472]_ ;
  assign \new_[23477]_  = ~A235 & ~A233;
  assign \new_[23478]_  = ~A201 & \new_[23477]_ ;
  assign \new_[23479]_  = \new_[23478]_  & \new_[23473]_ ;
  assign \new_[23483]_  = A266 & A265;
  assign \new_[23484]_  = ~A236 & \new_[23483]_ ;
  assign \new_[23488]_  = ~A302 & ~A301;
  assign \new_[23489]_  = A298 & \new_[23488]_ ;
  assign \new_[23490]_  = \new_[23489]_  & \new_[23484]_ ;
  assign \new_[23494]_  = ~A200 & A166;
  assign \new_[23495]_  = A168 & \new_[23494]_ ;
  assign \new_[23499]_  = ~A235 & ~A233;
  assign \new_[23500]_  = ~A201 & \new_[23499]_ ;
  assign \new_[23501]_  = \new_[23500]_  & \new_[23495]_ ;
  assign \new_[23505]_  = ~A268 & ~A266;
  assign \new_[23506]_  = ~A236 & \new_[23505]_ ;
  assign \new_[23510]_  = ~A300 & A298;
  assign \new_[23511]_  = ~A269 & \new_[23510]_ ;
  assign \new_[23512]_  = \new_[23511]_  & \new_[23506]_ ;
  assign \new_[23516]_  = ~A200 & A166;
  assign \new_[23517]_  = A168 & \new_[23516]_ ;
  assign \new_[23521]_  = ~A235 & ~A233;
  assign \new_[23522]_  = ~A201 & \new_[23521]_ ;
  assign \new_[23523]_  = \new_[23522]_  & \new_[23517]_ ;
  assign \new_[23527]_  = ~A268 & ~A266;
  assign \new_[23528]_  = ~A236 & \new_[23527]_ ;
  assign \new_[23532]_  = A299 & A298;
  assign \new_[23533]_  = ~A269 & \new_[23532]_ ;
  assign \new_[23534]_  = \new_[23533]_  & \new_[23528]_ ;
  assign \new_[23538]_  = ~A200 & A166;
  assign \new_[23539]_  = A168 & \new_[23538]_ ;
  assign \new_[23543]_  = ~A235 & ~A233;
  assign \new_[23544]_  = ~A201 & \new_[23543]_ ;
  assign \new_[23545]_  = \new_[23544]_  & \new_[23539]_ ;
  assign \new_[23549]_  = ~A268 & ~A266;
  assign \new_[23550]_  = ~A236 & \new_[23549]_ ;
  assign \new_[23554]_  = ~A299 & ~A298;
  assign \new_[23555]_  = ~A269 & \new_[23554]_ ;
  assign \new_[23556]_  = \new_[23555]_  & \new_[23550]_ ;
  assign \new_[23560]_  = ~A200 & A166;
  assign \new_[23561]_  = A168 & \new_[23560]_ ;
  assign \new_[23565]_  = ~A235 & ~A233;
  assign \new_[23566]_  = ~A201 & \new_[23565]_ ;
  assign \new_[23567]_  = \new_[23566]_  & \new_[23561]_ ;
  assign \new_[23571]_  = ~A267 & ~A266;
  assign \new_[23572]_  = ~A236 & \new_[23571]_ ;
  assign \new_[23576]_  = ~A302 & ~A301;
  assign \new_[23577]_  = A298 & \new_[23576]_ ;
  assign \new_[23578]_  = \new_[23577]_  & \new_[23572]_ ;
  assign \new_[23582]_  = ~A200 & A166;
  assign \new_[23583]_  = A168 & \new_[23582]_ ;
  assign \new_[23587]_  = ~A235 & ~A233;
  assign \new_[23588]_  = ~A201 & \new_[23587]_ ;
  assign \new_[23589]_  = \new_[23588]_  & \new_[23583]_ ;
  assign \new_[23593]_  = ~A266 & ~A265;
  assign \new_[23594]_  = ~A236 & \new_[23593]_ ;
  assign \new_[23598]_  = ~A302 & ~A301;
  assign \new_[23599]_  = A298 & \new_[23598]_ ;
  assign \new_[23600]_  = \new_[23599]_  & \new_[23594]_ ;
  assign \new_[23604]_  = ~A200 & A166;
  assign \new_[23605]_  = A168 & \new_[23604]_ ;
  assign \new_[23609]_  = ~A234 & ~A233;
  assign \new_[23610]_  = ~A201 & \new_[23609]_ ;
  assign \new_[23611]_  = \new_[23610]_  & \new_[23605]_ ;
  assign \new_[23615]_  = ~A269 & ~A268;
  assign \new_[23616]_  = ~A266 & \new_[23615]_ ;
  assign \new_[23620]_  = ~A302 & ~A301;
  assign \new_[23621]_  = A298 & \new_[23620]_ ;
  assign \new_[23622]_  = \new_[23621]_  & \new_[23616]_ ;
  assign \new_[23626]_  = ~A200 & A166;
  assign \new_[23627]_  = A168 & \new_[23626]_ ;
  assign \new_[23631]_  = ~A233 & A232;
  assign \new_[23632]_  = ~A201 & \new_[23631]_ ;
  assign \new_[23633]_  = \new_[23632]_  & \new_[23627]_ ;
  assign \new_[23637]_  = A298 & A235;
  assign \new_[23638]_  = A234 & \new_[23637]_ ;
  assign \new_[23642]_  = A301 & A300;
  assign \new_[23643]_  = ~A299 & \new_[23642]_ ;
  assign \new_[23644]_  = \new_[23643]_  & \new_[23638]_ ;
  assign \new_[23648]_  = ~A200 & A166;
  assign \new_[23649]_  = A168 & \new_[23648]_ ;
  assign \new_[23653]_  = ~A233 & A232;
  assign \new_[23654]_  = ~A201 & \new_[23653]_ ;
  assign \new_[23655]_  = \new_[23654]_  & \new_[23649]_ ;
  assign \new_[23659]_  = A298 & A235;
  assign \new_[23660]_  = A234 & \new_[23659]_ ;
  assign \new_[23664]_  = A302 & A300;
  assign \new_[23665]_  = ~A299 & \new_[23664]_ ;
  assign \new_[23666]_  = \new_[23665]_  & \new_[23660]_ ;
  assign \new_[23670]_  = ~A200 & A166;
  assign \new_[23671]_  = A168 & \new_[23670]_ ;
  assign \new_[23675]_  = ~A233 & A232;
  assign \new_[23676]_  = ~A201 & \new_[23675]_ ;
  assign \new_[23677]_  = \new_[23676]_  & \new_[23671]_ ;
  assign \new_[23681]_  = A265 & A235;
  assign \new_[23682]_  = A234 & \new_[23681]_ ;
  assign \new_[23686]_  = A268 & A267;
  assign \new_[23687]_  = ~A266 & \new_[23686]_ ;
  assign \new_[23688]_  = \new_[23687]_  & \new_[23682]_ ;
  assign \new_[23692]_  = ~A200 & A166;
  assign \new_[23693]_  = A168 & \new_[23692]_ ;
  assign \new_[23697]_  = ~A233 & A232;
  assign \new_[23698]_  = ~A201 & \new_[23697]_ ;
  assign \new_[23699]_  = \new_[23698]_  & \new_[23693]_ ;
  assign \new_[23703]_  = A265 & A235;
  assign \new_[23704]_  = A234 & \new_[23703]_ ;
  assign \new_[23708]_  = A269 & A267;
  assign \new_[23709]_  = ~A266 & \new_[23708]_ ;
  assign \new_[23710]_  = \new_[23709]_  & \new_[23704]_ ;
  assign \new_[23714]_  = ~A200 & A166;
  assign \new_[23715]_  = A168 & \new_[23714]_ ;
  assign \new_[23719]_  = ~A233 & A232;
  assign \new_[23720]_  = ~A201 & \new_[23719]_ ;
  assign \new_[23721]_  = \new_[23720]_  & \new_[23715]_ ;
  assign \new_[23725]_  = A298 & A236;
  assign \new_[23726]_  = A234 & \new_[23725]_ ;
  assign \new_[23730]_  = A301 & A300;
  assign \new_[23731]_  = ~A299 & \new_[23730]_ ;
  assign \new_[23732]_  = \new_[23731]_  & \new_[23726]_ ;
  assign \new_[23736]_  = ~A200 & A166;
  assign \new_[23737]_  = A168 & \new_[23736]_ ;
  assign \new_[23741]_  = ~A233 & A232;
  assign \new_[23742]_  = ~A201 & \new_[23741]_ ;
  assign \new_[23743]_  = \new_[23742]_  & \new_[23737]_ ;
  assign \new_[23747]_  = A298 & A236;
  assign \new_[23748]_  = A234 & \new_[23747]_ ;
  assign \new_[23752]_  = A302 & A300;
  assign \new_[23753]_  = ~A299 & \new_[23752]_ ;
  assign \new_[23754]_  = \new_[23753]_  & \new_[23748]_ ;
  assign \new_[23758]_  = ~A200 & A166;
  assign \new_[23759]_  = A168 & \new_[23758]_ ;
  assign \new_[23763]_  = ~A233 & A232;
  assign \new_[23764]_  = ~A201 & \new_[23763]_ ;
  assign \new_[23765]_  = \new_[23764]_  & \new_[23759]_ ;
  assign \new_[23769]_  = A265 & A236;
  assign \new_[23770]_  = A234 & \new_[23769]_ ;
  assign \new_[23774]_  = A268 & A267;
  assign \new_[23775]_  = ~A266 & \new_[23774]_ ;
  assign \new_[23776]_  = \new_[23775]_  & \new_[23770]_ ;
  assign \new_[23780]_  = ~A200 & A166;
  assign \new_[23781]_  = A168 & \new_[23780]_ ;
  assign \new_[23785]_  = ~A233 & A232;
  assign \new_[23786]_  = ~A201 & \new_[23785]_ ;
  assign \new_[23787]_  = \new_[23786]_  & \new_[23781]_ ;
  assign \new_[23791]_  = A265 & A236;
  assign \new_[23792]_  = A234 & \new_[23791]_ ;
  assign \new_[23796]_  = A269 & A267;
  assign \new_[23797]_  = ~A266 & \new_[23796]_ ;
  assign \new_[23798]_  = \new_[23797]_  & \new_[23792]_ ;
  assign \new_[23802]_  = ~A200 & A166;
  assign \new_[23803]_  = A168 & \new_[23802]_ ;
  assign \new_[23807]_  = ~A233 & ~A232;
  assign \new_[23808]_  = ~A201 & \new_[23807]_ ;
  assign \new_[23809]_  = \new_[23808]_  & \new_[23803]_ ;
  assign \new_[23813]_  = ~A269 & ~A268;
  assign \new_[23814]_  = ~A266 & \new_[23813]_ ;
  assign \new_[23818]_  = ~A302 & ~A301;
  assign \new_[23819]_  = A298 & \new_[23818]_ ;
  assign \new_[23820]_  = \new_[23819]_  & \new_[23814]_ ;
  assign \new_[23824]_  = ~A199 & A166;
  assign \new_[23825]_  = A168 & \new_[23824]_ ;
  assign \new_[23829]_  = A233 & A232;
  assign \new_[23830]_  = ~A200 & \new_[23829]_ ;
  assign \new_[23831]_  = \new_[23830]_  & \new_[23825]_ ;
  assign \new_[23835]_  = ~A269 & ~A268;
  assign \new_[23836]_  = A265 & \new_[23835]_ ;
  assign \new_[23840]_  = ~A302 & ~A301;
  assign \new_[23841]_  = ~A299 & \new_[23840]_ ;
  assign \new_[23842]_  = \new_[23841]_  & \new_[23836]_ ;
  assign \new_[23846]_  = ~A199 & A166;
  assign \new_[23847]_  = A168 & \new_[23846]_ ;
  assign \new_[23851]_  = ~A235 & ~A233;
  assign \new_[23852]_  = ~A200 & \new_[23851]_ ;
  assign \new_[23853]_  = \new_[23852]_  & \new_[23847]_ ;
  assign \new_[23857]_  = A266 & A265;
  assign \new_[23858]_  = ~A236 & \new_[23857]_ ;
  assign \new_[23862]_  = ~A302 & ~A301;
  assign \new_[23863]_  = A298 & \new_[23862]_ ;
  assign \new_[23864]_  = \new_[23863]_  & \new_[23858]_ ;
  assign \new_[23868]_  = ~A199 & A166;
  assign \new_[23869]_  = A168 & \new_[23868]_ ;
  assign \new_[23873]_  = ~A235 & ~A233;
  assign \new_[23874]_  = ~A200 & \new_[23873]_ ;
  assign \new_[23875]_  = \new_[23874]_  & \new_[23869]_ ;
  assign \new_[23879]_  = ~A268 & ~A266;
  assign \new_[23880]_  = ~A236 & \new_[23879]_ ;
  assign \new_[23884]_  = ~A300 & A298;
  assign \new_[23885]_  = ~A269 & \new_[23884]_ ;
  assign \new_[23886]_  = \new_[23885]_  & \new_[23880]_ ;
  assign \new_[23890]_  = ~A199 & A166;
  assign \new_[23891]_  = A168 & \new_[23890]_ ;
  assign \new_[23895]_  = ~A235 & ~A233;
  assign \new_[23896]_  = ~A200 & \new_[23895]_ ;
  assign \new_[23897]_  = \new_[23896]_  & \new_[23891]_ ;
  assign \new_[23901]_  = ~A268 & ~A266;
  assign \new_[23902]_  = ~A236 & \new_[23901]_ ;
  assign \new_[23906]_  = A299 & A298;
  assign \new_[23907]_  = ~A269 & \new_[23906]_ ;
  assign \new_[23908]_  = \new_[23907]_  & \new_[23902]_ ;
  assign \new_[23912]_  = ~A199 & A166;
  assign \new_[23913]_  = A168 & \new_[23912]_ ;
  assign \new_[23917]_  = ~A235 & ~A233;
  assign \new_[23918]_  = ~A200 & \new_[23917]_ ;
  assign \new_[23919]_  = \new_[23918]_  & \new_[23913]_ ;
  assign \new_[23923]_  = ~A268 & ~A266;
  assign \new_[23924]_  = ~A236 & \new_[23923]_ ;
  assign \new_[23928]_  = ~A299 & ~A298;
  assign \new_[23929]_  = ~A269 & \new_[23928]_ ;
  assign \new_[23930]_  = \new_[23929]_  & \new_[23924]_ ;
  assign \new_[23934]_  = ~A199 & A166;
  assign \new_[23935]_  = A168 & \new_[23934]_ ;
  assign \new_[23939]_  = ~A235 & ~A233;
  assign \new_[23940]_  = ~A200 & \new_[23939]_ ;
  assign \new_[23941]_  = \new_[23940]_  & \new_[23935]_ ;
  assign \new_[23945]_  = ~A267 & ~A266;
  assign \new_[23946]_  = ~A236 & \new_[23945]_ ;
  assign \new_[23950]_  = ~A302 & ~A301;
  assign \new_[23951]_  = A298 & \new_[23950]_ ;
  assign \new_[23952]_  = \new_[23951]_  & \new_[23946]_ ;
  assign \new_[23956]_  = ~A199 & A166;
  assign \new_[23957]_  = A168 & \new_[23956]_ ;
  assign \new_[23961]_  = ~A235 & ~A233;
  assign \new_[23962]_  = ~A200 & \new_[23961]_ ;
  assign \new_[23963]_  = \new_[23962]_  & \new_[23957]_ ;
  assign \new_[23967]_  = ~A266 & ~A265;
  assign \new_[23968]_  = ~A236 & \new_[23967]_ ;
  assign \new_[23972]_  = ~A302 & ~A301;
  assign \new_[23973]_  = A298 & \new_[23972]_ ;
  assign \new_[23974]_  = \new_[23973]_  & \new_[23968]_ ;
  assign \new_[23978]_  = ~A199 & A166;
  assign \new_[23979]_  = A168 & \new_[23978]_ ;
  assign \new_[23983]_  = ~A234 & ~A233;
  assign \new_[23984]_  = ~A200 & \new_[23983]_ ;
  assign \new_[23985]_  = \new_[23984]_  & \new_[23979]_ ;
  assign \new_[23989]_  = ~A269 & ~A268;
  assign \new_[23990]_  = ~A266 & \new_[23989]_ ;
  assign \new_[23994]_  = ~A302 & ~A301;
  assign \new_[23995]_  = A298 & \new_[23994]_ ;
  assign \new_[23996]_  = \new_[23995]_  & \new_[23990]_ ;
  assign \new_[24000]_  = ~A199 & A166;
  assign \new_[24001]_  = A168 & \new_[24000]_ ;
  assign \new_[24005]_  = ~A233 & A232;
  assign \new_[24006]_  = ~A200 & \new_[24005]_ ;
  assign \new_[24007]_  = \new_[24006]_  & \new_[24001]_ ;
  assign \new_[24011]_  = A298 & A235;
  assign \new_[24012]_  = A234 & \new_[24011]_ ;
  assign \new_[24016]_  = A301 & A300;
  assign \new_[24017]_  = ~A299 & \new_[24016]_ ;
  assign \new_[24018]_  = \new_[24017]_  & \new_[24012]_ ;
  assign \new_[24022]_  = ~A199 & A166;
  assign \new_[24023]_  = A168 & \new_[24022]_ ;
  assign \new_[24027]_  = ~A233 & A232;
  assign \new_[24028]_  = ~A200 & \new_[24027]_ ;
  assign \new_[24029]_  = \new_[24028]_  & \new_[24023]_ ;
  assign \new_[24033]_  = A298 & A235;
  assign \new_[24034]_  = A234 & \new_[24033]_ ;
  assign \new_[24038]_  = A302 & A300;
  assign \new_[24039]_  = ~A299 & \new_[24038]_ ;
  assign \new_[24040]_  = \new_[24039]_  & \new_[24034]_ ;
  assign \new_[24044]_  = ~A199 & A166;
  assign \new_[24045]_  = A168 & \new_[24044]_ ;
  assign \new_[24049]_  = ~A233 & A232;
  assign \new_[24050]_  = ~A200 & \new_[24049]_ ;
  assign \new_[24051]_  = \new_[24050]_  & \new_[24045]_ ;
  assign \new_[24055]_  = A265 & A235;
  assign \new_[24056]_  = A234 & \new_[24055]_ ;
  assign \new_[24060]_  = A268 & A267;
  assign \new_[24061]_  = ~A266 & \new_[24060]_ ;
  assign \new_[24062]_  = \new_[24061]_  & \new_[24056]_ ;
  assign \new_[24066]_  = ~A199 & A166;
  assign \new_[24067]_  = A168 & \new_[24066]_ ;
  assign \new_[24071]_  = ~A233 & A232;
  assign \new_[24072]_  = ~A200 & \new_[24071]_ ;
  assign \new_[24073]_  = \new_[24072]_  & \new_[24067]_ ;
  assign \new_[24077]_  = A265 & A235;
  assign \new_[24078]_  = A234 & \new_[24077]_ ;
  assign \new_[24082]_  = A269 & A267;
  assign \new_[24083]_  = ~A266 & \new_[24082]_ ;
  assign \new_[24084]_  = \new_[24083]_  & \new_[24078]_ ;
  assign \new_[24088]_  = ~A199 & A166;
  assign \new_[24089]_  = A168 & \new_[24088]_ ;
  assign \new_[24093]_  = ~A233 & A232;
  assign \new_[24094]_  = ~A200 & \new_[24093]_ ;
  assign \new_[24095]_  = \new_[24094]_  & \new_[24089]_ ;
  assign \new_[24099]_  = A298 & A236;
  assign \new_[24100]_  = A234 & \new_[24099]_ ;
  assign \new_[24104]_  = A301 & A300;
  assign \new_[24105]_  = ~A299 & \new_[24104]_ ;
  assign \new_[24106]_  = \new_[24105]_  & \new_[24100]_ ;
  assign \new_[24110]_  = ~A199 & A166;
  assign \new_[24111]_  = A168 & \new_[24110]_ ;
  assign \new_[24115]_  = ~A233 & A232;
  assign \new_[24116]_  = ~A200 & \new_[24115]_ ;
  assign \new_[24117]_  = \new_[24116]_  & \new_[24111]_ ;
  assign \new_[24121]_  = A298 & A236;
  assign \new_[24122]_  = A234 & \new_[24121]_ ;
  assign \new_[24126]_  = A302 & A300;
  assign \new_[24127]_  = ~A299 & \new_[24126]_ ;
  assign \new_[24128]_  = \new_[24127]_  & \new_[24122]_ ;
  assign \new_[24132]_  = ~A199 & A166;
  assign \new_[24133]_  = A168 & \new_[24132]_ ;
  assign \new_[24137]_  = ~A233 & A232;
  assign \new_[24138]_  = ~A200 & \new_[24137]_ ;
  assign \new_[24139]_  = \new_[24138]_  & \new_[24133]_ ;
  assign \new_[24143]_  = A265 & A236;
  assign \new_[24144]_  = A234 & \new_[24143]_ ;
  assign \new_[24148]_  = A268 & A267;
  assign \new_[24149]_  = ~A266 & \new_[24148]_ ;
  assign \new_[24150]_  = \new_[24149]_  & \new_[24144]_ ;
  assign \new_[24154]_  = ~A199 & A166;
  assign \new_[24155]_  = A168 & \new_[24154]_ ;
  assign \new_[24159]_  = ~A233 & A232;
  assign \new_[24160]_  = ~A200 & \new_[24159]_ ;
  assign \new_[24161]_  = \new_[24160]_  & \new_[24155]_ ;
  assign \new_[24165]_  = A265 & A236;
  assign \new_[24166]_  = A234 & \new_[24165]_ ;
  assign \new_[24170]_  = A269 & A267;
  assign \new_[24171]_  = ~A266 & \new_[24170]_ ;
  assign \new_[24172]_  = \new_[24171]_  & \new_[24166]_ ;
  assign \new_[24176]_  = ~A199 & A166;
  assign \new_[24177]_  = A168 & \new_[24176]_ ;
  assign \new_[24181]_  = ~A233 & ~A232;
  assign \new_[24182]_  = ~A200 & \new_[24181]_ ;
  assign \new_[24183]_  = \new_[24182]_  & \new_[24177]_ ;
  assign \new_[24187]_  = ~A269 & ~A268;
  assign \new_[24188]_  = ~A266 & \new_[24187]_ ;
  assign \new_[24192]_  = ~A302 & ~A301;
  assign \new_[24193]_  = A298 & \new_[24192]_ ;
  assign \new_[24194]_  = \new_[24193]_  & \new_[24188]_ ;
  assign \new_[24198]_  = A199 & A167;
  assign \new_[24199]_  = A168 & \new_[24198]_ ;
  assign \new_[24203]_  = A233 & A232;
  assign \new_[24204]_  = A200 & \new_[24203]_ ;
  assign \new_[24205]_  = \new_[24204]_  & \new_[24199]_ ;
  assign \new_[24209]_  = ~A269 & ~A268;
  assign \new_[24210]_  = A265 & \new_[24209]_ ;
  assign \new_[24214]_  = ~A302 & ~A301;
  assign \new_[24215]_  = ~A299 & \new_[24214]_ ;
  assign \new_[24216]_  = \new_[24215]_  & \new_[24210]_ ;
  assign \new_[24220]_  = A199 & A167;
  assign \new_[24221]_  = A168 & \new_[24220]_ ;
  assign \new_[24225]_  = ~A235 & ~A233;
  assign \new_[24226]_  = A200 & \new_[24225]_ ;
  assign \new_[24227]_  = \new_[24226]_  & \new_[24221]_ ;
  assign \new_[24231]_  = A266 & A265;
  assign \new_[24232]_  = ~A236 & \new_[24231]_ ;
  assign \new_[24236]_  = ~A302 & ~A301;
  assign \new_[24237]_  = A298 & \new_[24236]_ ;
  assign \new_[24238]_  = \new_[24237]_  & \new_[24232]_ ;
  assign \new_[24242]_  = A199 & A167;
  assign \new_[24243]_  = A168 & \new_[24242]_ ;
  assign \new_[24247]_  = ~A235 & ~A233;
  assign \new_[24248]_  = A200 & \new_[24247]_ ;
  assign \new_[24249]_  = \new_[24248]_  & \new_[24243]_ ;
  assign \new_[24253]_  = ~A268 & ~A266;
  assign \new_[24254]_  = ~A236 & \new_[24253]_ ;
  assign \new_[24258]_  = ~A300 & A298;
  assign \new_[24259]_  = ~A269 & \new_[24258]_ ;
  assign \new_[24260]_  = \new_[24259]_  & \new_[24254]_ ;
  assign \new_[24264]_  = A199 & A167;
  assign \new_[24265]_  = A168 & \new_[24264]_ ;
  assign \new_[24269]_  = ~A235 & ~A233;
  assign \new_[24270]_  = A200 & \new_[24269]_ ;
  assign \new_[24271]_  = \new_[24270]_  & \new_[24265]_ ;
  assign \new_[24275]_  = ~A268 & ~A266;
  assign \new_[24276]_  = ~A236 & \new_[24275]_ ;
  assign \new_[24280]_  = A299 & A298;
  assign \new_[24281]_  = ~A269 & \new_[24280]_ ;
  assign \new_[24282]_  = \new_[24281]_  & \new_[24276]_ ;
  assign \new_[24286]_  = A199 & A167;
  assign \new_[24287]_  = A168 & \new_[24286]_ ;
  assign \new_[24291]_  = ~A235 & ~A233;
  assign \new_[24292]_  = A200 & \new_[24291]_ ;
  assign \new_[24293]_  = \new_[24292]_  & \new_[24287]_ ;
  assign \new_[24297]_  = ~A268 & ~A266;
  assign \new_[24298]_  = ~A236 & \new_[24297]_ ;
  assign \new_[24302]_  = ~A299 & ~A298;
  assign \new_[24303]_  = ~A269 & \new_[24302]_ ;
  assign \new_[24304]_  = \new_[24303]_  & \new_[24298]_ ;
  assign \new_[24308]_  = A199 & A167;
  assign \new_[24309]_  = A168 & \new_[24308]_ ;
  assign \new_[24313]_  = ~A235 & ~A233;
  assign \new_[24314]_  = A200 & \new_[24313]_ ;
  assign \new_[24315]_  = \new_[24314]_  & \new_[24309]_ ;
  assign \new_[24319]_  = ~A267 & ~A266;
  assign \new_[24320]_  = ~A236 & \new_[24319]_ ;
  assign \new_[24324]_  = ~A302 & ~A301;
  assign \new_[24325]_  = A298 & \new_[24324]_ ;
  assign \new_[24326]_  = \new_[24325]_  & \new_[24320]_ ;
  assign \new_[24330]_  = A199 & A167;
  assign \new_[24331]_  = A168 & \new_[24330]_ ;
  assign \new_[24335]_  = ~A235 & ~A233;
  assign \new_[24336]_  = A200 & \new_[24335]_ ;
  assign \new_[24337]_  = \new_[24336]_  & \new_[24331]_ ;
  assign \new_[24341]_  = ~A266 & ~A265;
  assign \new_[24342]_  = ~A236 & \new_[24341]_ ;
  assign \new_[24346]_  = ~A302 & ~A301;
  assign \new_[24347]_  = A298 & \new_[24346]_ ;
  assign \new_[24348]_  = \new_[24347]_  & \new_[24342]_ ;
  assign \new_[24352]_  = A199 & A167;
  assign \new_[24353]_  = A168 & \new_[24352]_ ;
  assign \new_[24357]_  = ~A234 & ~A233;
  assign \new_[24358]_  = A200 & \new_[24357]_ ;
  assign \new_[24359]_  = \new_[24358]_  & \new_[24353]_ ;
  assign \new_[24363]_  = ~A269 & ~A268;
  assign \new_[24364]_  = ~A266 & \new_[24363]_ ;
  assign \new_[24368]_  = ~A302 & ~A301;
  assign \new_[24369]_  = A298 & \new_[24368]_ ;
  assign \new_[24370]_  = \new_[24369]_  & \new_[24364]_ ;
  assign \new_[24374]_  = A199 & A167;
  assign \new_[24375]_  = A168 & \new_[24374]_ ;
  assign \new_[24379]_  = ~A233 & A232;
  assign \new_[24380]_  = A200 & \new_[24379]_ ;
  assign \new_[24381]_  = \new_[24380]_  & \new_[24375]_ ;
  assign \new_[24385]_  = A298 & A235;
  assign \new_[24386]_  = A234 & \new_[24385]_ ;
  assign \new_[24390]_  = A301 & A300;
  assign \new_[24391]_  = ~A299 & \new_[24390]_ ;
  assign \new_[24392]_  = \new_[24391]_  & \new_[24386]_ ;
  assign \new_[24396]_  = A199 & A167;
  assign \new_[24397]_  = A168 & \new_[24396]_ ;
  assign \new_[24401]_  = ~A233 & A232;
  assign \new_[24402]_  = A200 & \new_[24401]_ ;
  assign \new_[24403]_  = \new_[24402]_  & \new_[24397]_ ;
  assign \new_[24407]_  = A298 & A235;
  assign \new_[24408]_  = A234 & \new_[24407]_ ;
  assign \new_[24412]_  = A302 & A300;
  assign \new_[24413]_  = ~A299 & \new_[24412]_ ;
  assign \new_[24414]_  = \new_[24413]_  & \new_[24408]_ ;
  assign \new_[24418]_  = A199 & A167;
  assign \new_[24419]_  = A168 & \new_[24418]_ ;
  assign \new_[24423]_  = ~A233 & A232;
  assign \new_[24424]_  = A200 & \new_[24423]_ ;
  assign \new_[24425]_  = \new_[24424]_  & \new_[24419]_ ;
  assign \new_[24429]_  = A265 & A235;
  assign \new_[24430]_  = A234 & \new_[24429]_ ;
  assign \new_[24434]_  = A268 & A267;
  assign \new_[24435]_  = ~A266 & \new_[24434]_ ;
  assign \new_[24436]_  = \new_[24435]_  & \new_[24430]_ ;
  assign \new_[24440]_  = A199 & A167;
  assign \new_[24441]_  = A168 & \new_[24440]_ ;
  assign \new_[24445]_  = ~A233 & A232;
  assign \new_[24446]_  = A200 & \new_[24445]_ ;
  assign \new_[24447]_  = \new_[24446]_  & \new_[24441]_ ;
  assign \new_[24451]_  = A265 & A235;
  assign \new_[24452]_  = A234 & \new_[24451]_ ;
  assign \new_[24456]_  = A269 & A267;
  assign \new_[24457]_  = ~A266 & \new_[24456]_ ;
  assign \new_[24458]_  = \new_[24457]_  & \new_[24452]_ ;
  assign \new_[24462]_  = A199 & A167;
  assign \new_[24463]_  = A168 & \new_[24462]_ ;
  assign \new_[24467]_  = ~A233 & A232;
  assign \new_[24468]_  = A200 & \new_[24467]_ ;
  assign \new_[24469]_  = \new_[24468]_  & \new_[24463]_ ;
  assign \new_[24473]_  = A298 & A236;
  assign \new_[24474]_  = A234 & \new_[24473]_ ;
  assign \new_[24478]_  = A301 & A300;
  assign \new_[24479]_  = ~A299 & \new_[24478]_ ;
  assign \new_[24480]_  = \new_[24479]_  & \new_[24474]_ ;
  assign \new_[24484]_  = A199 & A167;
  assign \new_[24485]_  = A168 & \new_[24484]_ ;
  assign \new_[24489]_  = ~A233 & A232;
  assign \new_[24490]_  = A200 & \new_[24489]_ ;
  assign \new_[24491]_  = \new_[24490]_  & \new_[24485]_ ;
  assign \new_[24495]_  = A298 & A236;
  assign \new_[24496]_  = A234 & \new_[24495]_ ;
  assign \new_[24500]_  = A302 & A300;
  assign \new_[24501]_  = ~A299 & \new_[24500]_ ;
  assign \new_[24502]_  = \new_[24501]_  & \new_[24496]_ ;
  assign \new_[24506]_  = A199 & A167;
  assign \new_[24507]_  = A168 & \new_[24506]_ ;
  assign \new_[24511]_  = ~A233 & A232;
  assign \new_[24512]_  = A200 & \new_[24511]_ ;
  assign \new_[24513]_  = \new_[24512]_  & \new_[24507]_ ;
  assign \new_[24517]_  = A265 & A236;
  assign \new_[24518]_  = A234 & \new_[24517]_ ;
  assign \new_[24522]_  = A268 & A267;
  assign \new_[24523]_  = ~A266 & \new_[24522]_ ;
  assign \new_[24524]_  = \new_[24523]_  & \new_[24518]_ ;
  assign \new_[24528]_  = A199 & A167;
  assign \new_[24529]_  = A168 & \new_[24528]_ ;
  assign \new_[24533]_  = ~A233 & A232;
  assign \new_[24534]_  = A200 & \new_[24533]_ ;
  assign \new_[24535]_  = \new_[24534]_  & \new_[24529]_ ;
  assign \new_[24539]_  = A265 & A236;
  assign \new_[24540]_  = A234 & \new_[24539]_ ;
  assign \new_[24544]_  = A269 & A267;
  assign \new_[24545]_  = ~A266 & \new_[24544]_ ;
  assign \new_[24546]_  = \new_[24545]_  & \new_[24540]_ ;
  assign \new_[24550]_  = A199 & A167;
  assign \new_[24551]_  = A168 & \new_[24550]_ ;
  assign \new_[24555]_  = ~A233 & ~A232;
  assign \new_[24556]_  = A200 & \new_[24555]_ ;
  assign \new_[24557]_  = \new_[24556]_  & \new_[24551]_ ;
  assign \new_[24561]_  = ~A269 & ~A268;
  assign \new_[24562]_  = ~A266 & \new_[24561]_ ;
  assign \new_[24566]_  = ~A302 & ~A301;
  assign \new_[24567]_  = A298 & \new_[24566]_ ;
  assign \new_[24568]_  = \new_[24567]_  & \new_[24562]_ ;
  assign \new_[24572]_  = ~A200 & A167;
  assign \new_[24573]_  = A168 & \new_[24572]_ ;
  assign \new_[24577]_  = A232 & ~A203;
  assign \new_[24578]_  = ~A202 & \new_[24577]_ ;
  assign \new_[24579]_  = \new_[24578]_  & \new_[24573]_ ;
  assign \new_[24583]_  = ~A268 & A265;
  assign \new_[24584]_  = A233 & \new_[24583]_ ;
  assign \new_[24588]_  = ~A300 & ~A299;
  assign \new_[24589]_  = ~A269 & \new_[24588]_ ;
  assign \new_[24590]_  = \new_[24589]_  & \new_[24584]_ ;
  assign \new_[24594]_  = ~A200 & A167;
  assign \new_[24595]_  = A168 & \new_[24594]_ ;
  assign \new_[24599]_  = A232 & ~A203;
  assign \new_[24600]_  = ~A202 & \new_[24599]_ ;
  assign \new_[24601]_  = \new_[24600]_  & \new_[24595]_ ;
  assign \new_[24605]_  = ~A268 & A265;
  assign \new_[24606]_  = A233 & \new_[24605]_ ;
  assign \new_[24610]_  = A299 & A298;
  assign \new_[24611]_  = ~A269 & \new_[24610]_ ;
  assign \new_[24612]_  = \new_[24611]_  & \new_[24606]_ ;
  assign \new_[24616]_  = ~A200 & A167;
  assign \new_[24617]_  = A168 & \new_[24616]_ ;
  assign \new_[24621]_  = A232 & ~A203;
  assign \new_[24622]_  = ~A202 & \new_[24621]_ ;
  assign \new_[24623]_  = \new_[24622]_  & \new_[24617]_ ;
  assign \new_[24627]_  = ~A268 & A265;
  assign \new_[24628]_  = A233 & \new_[24627]_ ;
  assign \new_[24632]_  = ~A299 & ~A298;
  assign \new_[24633]_  = ~A269 & \new_[24632]_ ;
  assign \new_[24634]_  = \new_[24633]_  & \new_[24628]_ ;
  assign \new_[24638]_  = ~A200 & A167;
  assign \new_[24639]_  = A168 & \new_[24638]_ ;
  assign \new_[24643]_  = A232 & ~A203;
  assign \new_[24644]_  = ~A202 & \new_[24643]_ ;
  assign \new_[24645]_  = \new_[24644]_  & \new_[24639]_ ;
  assign \new_[24649]_  = ~A267 & A265;
  assign \new_[24650]_  = A233 & \new_[24649]_ ;
  assign \new_[24654]_  = ~A302 & ~A301;
  assign \new_[24655]_  = ~A299 & \new_[24654]_ ;
  assign \new_[24656]_  = \new_[24655]_  & \new_[24650]_ ;
  assign \new_[24660]_  = ~A200 & A167;
  assign \new_[24661]_  = A168 & \new_[24660]_ ;
  assign \new_[24665]_  = A232 & ~A203;
  assign \new_[24666]_  = ~A202 & \new_[24665]_ ;
  assign \new_[24667]_  = \new_[24666]_  & \new_[24661]_ ;
  assign \new_[24671]_  = A266 & A265;
  assign \new_[24672]_  = A233 & \new_[24671]_ ;
  assign \new_[24676]_  = ~A302 & ~A301;
  assign \new_[24677]_  = ~A299 & \new_[24676]_ ;
  assign \new_[24678]_  = \new_[24677]_  & \new_[24672]_ ;
  assign \new_[24682]_  = ~A200 & A167;
  assign \new_[24683]_  = A168 & \new_[24682]_ ;
  assign \new_[24687]_  = A232 & ~A203;
  assign \new_[24688]_  = ~A202 & \new_[24687]_ ;
  assign \new_[24689]_  = \new_[24688]_  & \new_[24683]_ ;
  assign \new_[24693]_  = ~A266 & ~A265;
  assign \new_[24694]_  = A233 & \new_[24693]_ ;
  assign \new_[24698]_  = ~A302 & ~A301;
  assign \new_[24699]_  = ~A299 & \new_[24698]_ ;
  assign \new_[24700]_  = \new_[24699]_  & \new_[24694]_ ;
  assign \new_[24704]_  = ~A200 & A167;
  assign \new_[24705]_  = A168 & \new_[24704]_ ;
  assign \new_[24709]_  = ~A233 & ~A203;
  assign \new_[24710]_  = ~A202 & \new_[24709]_ ;
  assign \new_[24711]_  = \new_[24710]_  & \new_[24705]_ ;
  assign \new_[24715]_  = A265 & ~A236;
  assign \new_[24716]_  = ~A235 & \new_[24715]_ ;
  assign \new_[24720]_  = ~A300 & A298;
  assign \new_[24721]_  = A266 & \new_[24720]_ ;
  assign \new_[24722]_  = \new_[24721]_  & \new_[24716]_ ;
  assign \new_[24726]_  = ~A200 & A167;
  assign \new_[24727]_  = A168 & \new_[24726]_ ;
  assign \new_[24731]_  = ~A233 & ~A203;
  assign \new_[24732]_  = ~A202 & \new_[24731]_ ;
  assign \new_[24733]_  = \new_[24732]_  & \new_[24727]_ ;
  assign \new_[24737]_  = A265 & ~A236;
  assign \new_[24738]_  = ~A235 & \new_[24737]_ ;
  assign \new_[24742]_  = A299 & A298;
  assign \new_[24743]_  = A266 & \new_[24742]_ ;
  assign \new_[24744]_  = \new_[24743]_  & \new_[24738]_ ;
  assign \new_[24748]_  = ~A200 & A167;
  assign \new_[24749]_  = A168 & \new_[24748]_ ;
  assign \new_[24753]_  = ~A233 & ~A203;
  assign \new_[24754]_  = ~A202 & \new_[24753]_ ;
  assign \new_[24755]_  = \new_[24754]_  & \new_[24749]_ ;
  assign \new_[24759]_  = A265 & ~A236;
  assign \new_[24760]_  = ~A235 & \new_[24759]_ ;
  assign \new_[24764]_  = ~A299 & ~A298;
  assign \new_[24765]_  = A266 & \new_[24764]_ ;
  assign \new_[24766]_  = \new_[24765]_  & \new_[24760]_ ;
  assign \new_[24770]_  = ~A200 & A167;
  assign \new_[24771]_  = A168 & \new_[24770]_ ;
  assign \new_[24775]_  = ~A233 & ~A203;
  assign \new_[24776]_  = ~A202 & \new_[24775]_ ;
  assign \new_[24777]_  = \new_[24776]_  & \new_[24771]_ ;
  assign \new_[24781]_  = ~A266 & ~A236;
  assign \new_[24782]_  = ~A235 & \new_[24781]_ ;
  assign \new_[24786]_  = ~A300 & A298;
  assign \new_[24787]_  = ~A267 & \new_[24786]_ ;
  assign \new_[24788]_  = \new_[24787]_  & \new_[24782]_ ;
  assign \new_[24792]_  = ~A200 & A167;
  assign \new_[24793]_  = A168 & \new_[24792]_ ;
  assign \new_[24797]_  = ~A233 & ~A203;
  assign \new_[24798]_  = ~A202 & \new_[24797]_ ;
  assign \new_[24799]_  = \new_[24798]_  & \new_[24793]_ ;
  assign \new_[24803]_  = ~A266 & ~A236;
  assign \new_[24804]_  = ~A235 & \new_[24803]_ ;
  assign \new_[24808]_  = A299 & A298;
  assign \new_[24809]_  = ~A267 & \new_[24808]_ ;
  assign \new_[24810]_  = \new_[24809]_  & \new_[24804]_ ;
  assign \new_[24814]_  = ~A200 & A167;
  assign \new_[24815]_  = A168 & \new_[24814]_ ;
  assign \new_[24819]_  = ~A233 & ~A203;
  assign \new_[24820]_  = ~A202 & \new_[24819]_ ;
  assign \new_[24821]_  = \new_[24820]_  & \new_[24815]_ ;
  assign \new_[24825]_  = ~A266 & ~A236;
  assign \new_[24826]_  = ~A235 & \new_[24825]_ ;
  assign \new_[24830]_  = ~A299 & ~A298;
  assign \new_[24831]_  = ~A267 & \new_[24830]_ ;
  assign \new_[24832]_  = \new_[24831]_  & \new_[24826]_ ;
  assign \new_[24836]_  = ~A200 & A167;
  assign \new_[24837]_  = A168 & \new_[24836]_ ;
  assign \new_[24841]_  = ~A233 & ~A203;
  assign \new_[24842]_  = ~A202 & \new_[24841]_ ;
  assign \new_[24843]_  = \new_[24842]_  & \new_[24837]_ ;
  assign \new_[24847]_  = ~A265 & ~A236;
  assign \new_[24848]_  = ~A235 & \new_[24847]_ ;
  assign \new_[24852]_  = ~A300 & A298;
  assign \new_[24853]_  = ~A266 & \new_[24852]_ ;
  assign \new_[24854]_  = \new_[24853]_  & \new_[24848]_ ;
  assign \new_[24858]_  = ~A200 & A167;
  assign \new_[24859]_  = A168 & \new_[24858]_ ;
  assign \new_[24863]_  = ~A233 & ~A203;
  assign \new_[24864]_  = ~A202 & \new_[24863]_ ;
  assign \new_[24865]_  = \new_[24864]_  & \new_[24859]_ ;
  assign \new_[24869]_  = ~A265 & ~A236;
  assign \new_[24870]_  = ~A235 & \new_[24869]_ ;
  assign \new_[24874]_  = A299 & A298;
  assign \new_[24875]_  = ~A266 & \new_[24874]_ ;
  assign \new_[24876]_  = \new_[24875]_  & \new_[24870]_ ;
  assign \new_[24880]_  = ~A200 & A167;
  assign \new_[24881]_  = A168 & \new_[24880]_ ;
  assign \new_[24885]_  = ~A233 & ~A203;
  assign \new_[24886]_  = ~A202 & \new_[24885]_ ;
  assign \new_[24887]_  = \new_[24886]_  & \new_[24881]_ ;
  assign \new_[24891]_  = ~A265 & ~A236;
  assign \new_[24892]_  = ~A235 & \new_[24891]_ ;
  assign \new_[24896]_  = ~A299 & ~A298;
  assign \new_[24897]_  = ~A266 & \new_[24896]_ ;
  assign \new_[24898]_  = \new_[24897]_  & \new_[24892]_ ;
  assign \new_[24902]_  = ~A200 & A167;
  assign \new_[24903]_  = A168 & \new_[24902]_ ;
  assign \new_[24907]_  = ~A233 & ~A203;
  assign \new_[24908]_  = ~A202 & \new_[24907]_ ;
  assign \new_[24909]_  = \new_[24908]_  & \new_[24903]_ ;
  assign \new_[24913]_  = A266 & A265;
  assign \new_[24914]_  = ~A234 & \new_[24913]_ ;
  assign \new_[24918]_  = ~A302 & ~A301;
  assign \new_[24919]_  = A298 & \new_[24918]_ ;
  assign \new_[24920]_  = \new_[24919]_  & \new_[24914]_ ;
  assign \new_[24924]_  = ~A200 & A167;
  assign \new_[24925]_  = A168 & \new_[24924]_ ;
  assign \new_[24929]_  = ~A233 & ~A203;
  assign \new_[24930]_  = ~A202 & \new_[24929]_ ;
  assign \new_[24931]_  = \new_[24930]_  & \new_[24925]_ ;
  assign \new_[24935]_  = ~A268 & ~A266;
  assign \new_[24936]_  = ~A234 & \new_[24935]_ ;
  assign \new_[24940]_  = ~A300 & A298;
  assign \new_[24941]_  = ~A269 & \new_[24940]_ ;
  assign \new_[24942]_  = \new_[24941]_  & \new_[24936]_ ;
  assign \new_[24946]_  = ~A200 & A167;
  assign \new_[24947]_  = A168 & \new_[24946]_ ;
  assign \new_[24951]_  = ~A233 & ~A203;
  assign \new_[24952]_  = ~A202 & \new_[24951]_ ;
  assign \new_[24953]_  = \new_[24952]_  & \new_[24947]_ ;
  assign \new_[24957]_  = ~A268 & ~A266;
  assign \new_[24958]_  = ~A234 & \new_[24957]_ ;
  assign \new_[24962]_  = A299 & A298;
  assign \new_[24963]_  = ~A269 & \new_[24962]_ ;
  assign \new_[24964]_  = \new_[24963]_  & \new_[24958]_ ;
  assign \new_[24968]_  = ~A200 & A167;
  assign \new_[24969]_  = A168 & \new_[24968]_ ;
  assign \new_[24973]_  = ~A233 & ~A203;
  assign \new_[24974]_  = ~A202 & \new_[24973]_ ;
  assign \new_[24975]_  = \new_[24974]_  & \new_[24969]_ ;
  assign \new_[24979]_  = ~A268 & ~A266;
  assign \new_[24980]_  = ~A234 & \new_[24979]_ ;
  assign \new_[24984]_  = ~A299 & ~A298;
  assign \new_[24985]_  = ~A269 & \new_[24984]_ ;
  assign \new_[24986]_  = \new_[24985]_  & \new_[24980]_ ;
  assign \new_[24990]_  = ~A200 & A167;
  assign \new_[24991]_  = A168 & \new_[24990]_ ;
  assign \new_[24995]_  = ~A233 & ~A203;
  assign \new_[24996]_  = ~A202 & \new_[24995]_ ;
  assign \new_[24997]_  = \new_[24996]_  & \new_[24991]_ ;
  assign \new_[25001]_  = ~A267 & ~A266;
  assign \new_[25002]_  = ~A234 & \new_[25001]_ ;
  assign \new_[25006]_  = ~A302 & ~A301;
  assign \new_[25007]_  = A298 & \new_[25006]_ ;
  assign \new_[25008]_  = \new_[25007]_  & \new_[25002]_ ;
  assign \new_[25012]_  = ~A200 & A167;
  assign \new_[25013]_  = A168 & \new_[25012]_ ;
  assign \new_[25017]_  = ~A233 & ~A203;
  assign \new_[25018]_  = ~A202 & \new_[25017]_ ;
  assign \new_[25019]_  = \new_[25018]_  & \new_[25013]_ ;
  assign \new_[25023]_  = ~A266 & ~A265;
  assign \new_[25024]_  = ~A234 & \new_[25023]_ ;
  assign \new_[25028]_  = ~A302 & ~A301;
  assign \new_[25029]_  = A298 & \new_[25028]_ ;
  assign \new_[25030]_  = \new_[25029]_  & \new_[25024]_ ;
  assign \new_[25034]_  = ~A200 & A167;
  assign \new_[25035]_  = A168 & \new_[25034]_ ;
  assign \new_[25039]_  = ~A232 & ~A203;
  assign \new_[25040]_  = ~A202 & \new_[25039]_ ;
  assign \new_[25041]_  = \new_[25040]_  & \new_[25035]_ ;
  assign \new_[25045]_  = A266 & A265;
  assign \new_[25046]_  = ~A233 & \new_[25045]_ ;
  assign \new_[25050]_  = ~A302 & ~A301;
  assign \new_[25051]_  = A298 & \new_[25050]_ ;
  assign \new_[25052]_  = \new_[25051]_  & \new_[25046]_ ;
  assign \new_[25056]_  = ~A200 & A167;
  assign \new_[25057]_  = A168 & \new_[25056]_ ;
  assign \new_[25061]_  = ~A232 & ~A203;
  assign \new_[25062]_  = ~A202 & \new_[25061]_ ;
  assign \new_[25063]_  = \new_[25062]_  & \new_[25057]_ ;
  assign \new_[25067]_  = ~A268 & ~A266;
  assign \new_[25068]_  = ~A233 & \new_[25067]_ ;
  assign \new_[25072]_  = ~A300 & A298;
  assign \new_[25073]_  = ~A269 & \new_[25072]_ ;
  assign \new_[25074]_  = \new_[25073]_  & \new_[25068]_ ;
  assign \new_[25078]_  = ~A200 & A167;
  assign \new_[25079]_  = A168 & \new_[25078]_ ;
  assign \new_[25083]_  = ~A232 & ~A203;
  assign \new_[25084]_  = ~A202 & \new_[25083]_ ;
  assign \new_[25085]_  = \new_[25084]_  & \new_[25079]_ ;
  assign \new_[25089]_  = ~A268 & ~A266;
  assign \new_[25090]_  = ~A233 & \new_[25089]_ ;
  assign \new_[25094]_  = A299 & A298;
  assign \new_[25095]_  = ~A269 & \new_[25094]_ ;
  assign \new_[25096]_  = \new_[25095]_  & \new_[25090]_ ;
  assign \new_[25100]_  = ~A200 & A167;
  assign \new_[25101]_  = A168 & \new_[25100]_ ;
  assign \new_[25105]_  = ~A232 & ~A203;
  assign \new_[25106]_  = ~A202 & \new_[25105]_ ;
  assign \new_[25107]_  = \new_[25106]_  & \new_[25101]_ ;
  assign \new_[25111]_  = ~A268 & ~A266;
  assign \new_[25112]_  = ~A233 & \new_[25111]_ ;
  assign \new_[25116]_  = ~A299 & ~A298;
  assign \new_[25117]_  = ~A269 & \new_[25116]_ ;
  assign \new_[25118]_  = \new_[25117]_  & \new_[25112]_ ;
  assign \new_[25122]_  = ~A200 & A167;
  assign \new_[25123]_  = A168 & \new_[25122]_ ;
  assign \new_[25127]_  = ~A232 & ~A203;
  assign \new_[25128]_  = ~A202 & \new_[25127]_ ;
  assign \new_[25129]_  = \new_[25128]_  & \new_[25123]_ ;
  assign \new_[25133]_  = ~A267 & ~A266;
  assign \new_[25134]_  = ~A233 & \new_[25133]_ ;
  assign \new_[25138]_  = ~A302 & ~A301;
  assign \new_[25139]_  = A298 & \new_[25138]_ ;
  assign \new_[25140]_  = \new_[25139]_  & \new_[25134]_ ;
  assign \new_[25144]_  = ~A200 & A167;
  assign \new_[25145]_  = A168 & \new_[25144]_ ;
  assign \new_[25149]_  = ~A232 & ~A203;
  assign \new_[25150]_  = ~A202 & \new_[25149]_ ;
  assign \new_[25151]_  = \new_[25150]_  & \new_[25145]_ ;
  assign \new_[25155]_  = ~A266 & ~A265;
  assign \new_[25156]_  = ~A233 & \new_[25155]_ ;
  assign \new_[25160]_  = ~A302 & ~A301;
  assign \new_[25161]_  = A298 & \new_[25160]_ ;
  assign \new_[25162]_  = \new_[25161]_  & \new_[25156]_ ;
  assign \new_[25166]_  = ~A200 & A167;
  assign \new_[25167]_  = A168 & \new_[25166]_ ;
  assign \new_[25171]_  = A233 & A232;
  assign \new_[25172]_  = ~A201 & \new_[25171]_ ;
  assign \new_[25173]_  = \new_[25172]_  & \new_[25167]_ ;
  assign \new_[25177]_  = ~A269 & ~A268;
  assign \new_[25178]_  = A265 & \new_[25177]_ ;
  assign \new_[25182]_  = ~A302 & ~A301;
  assign \new_[25183]_  = ~A299 & \new_[25182]_ ;
  assign \new_[25184]_  = \new_[25183]_  & \new_[25178]_ ;
  assign \new_[25188]_  = ~A200 & A167;
  assign \new_[25189]_  = A168 & \new_[25188]_ ;
  assign \new_[25193]_  = ~A235 & ~A233;
  assign \new_[25194]_  = ~A201 & \new_[25193]_ ;
  assign \new_[25195]_  = \new_[25194]_  & \new_[25189]_ ;
  assign \new_[25199]_  = A266 & A265;
  assign \new_[25200]_  = ~A236 & \new_[25199]_ ;
  assign \new_[25204]_  = ~A302 & ~A301;
  assign \new_[25205]_  = A298 & \new_[25204]_ ;
  assign \new_[25206]_  = \new_[25205]_  & \new_[25200]_ ;
  assign \new_[25210]_  = ~A200 & A167;
  assign \new_[25211]_  = A168 & \new_[25210]_ ;
  assign \new_[25215]_  = ~A235 & ~A233;
  assign \new_[25216]_  = ~A201 & \new_[25215]_ ;
  assign \new_[25217]_  = \new_[25216]_  & \new_[25211]_ ;
  assign \new_[25221]_  = ~A268 & ~A266;
  assign \new_[25222]_  = ~A236 & \new_[25221]_ ;
  assign \new_[25226]_  = ~A300 & A298;
  assign \new_[25227]_  = ~A269 & \new_[25226]_ ;
  assign \new_[25228]_  = \new_[25227]_  & \new_[25222]_ ;
  assign \new_[25232]_  = ~A200 & A167;
  assign \new_[25233]_  = A168 & \new_[25232]_ ;
  assign \new_[25237]_  = ~A235 & ~A233;
  assign \new_[25238]_  = ~A201 & \new_[25237]_ ;
  assign \new_[25239]_  = \new_[25238]_  & \new_[25233]_ ;
  assign \new_[25243]_  = ~A268 & ~A266;
  assign \new_[25244]_  = ~A236 & \new_[25243]_ ;
  assign \new_[25248]_  = A299 & A298;
  assign \new_[25249]_  = ~A269 & \new_[25248]_ ;
  assign \new_[25250]_  = \new_[25249]_  & \new_[25244]_ ;
  assign \new_[25254]_  = ~A200 & A167;
  assign \new_[25255]_  = A168 & \new_[25254]_ ;
  assign \new_[25259]_  = ~A235 & ~A233;
  assign \new_[25260]_  = ~A201 & \new_[25259]_ ;
  assign \new_[25261]_  = \new_[25260]_  & \new_[25255]_ ;
  assign \new_[25265]_  = ~A268 & ~A266;
  assign \new_[25266]_  = ~A236 & \new_[25265]_ ;
  assign \new_[25270]_  = ~A299 & ~A298;
  assign \new_[25271]_  = ~A269 & \new_[25270]_ ;
  assign \new_[25272]_  = \new_[25271]_  & \new_[25266]_ ;
  assign \new_[25276]_  = ~A200 & A167;
  assign \new_[25277]_  = A168 & \new_[25276]_ ;
  assign \new_[25281]_  = ~A235 & ~A233;
  assign \new_[25282]_  = ~A201 & \new_[25281]_ ;
  assign \new_[25283]_  = \new_[25282]_  & \new_[25277]_ ;
  assign \new_[25287]_  = ~A267 & ~A266;
  assign \new_[25288]_  = ~A236 & \new_[25287]_ ;
  assign \new_[25292]_  = ~A302 & ~A301;
  assign \new_[25293]_  = A298 & \new_[25292]_ ;
  assign \new_[25294]_  = \new_[25293]_  & \new_[25288]_ ;
  assign \new_[25298]_  = ~A200 & A167;
  assign \new_[25299]_  = A168 & \new_[25298]_ ;
  assign \new_[25303]_  = ~A235 & ~A233;
  assign \new_[25304]_  = ~A201 & \new_[25303]_ ;
  assign \new_[25305]_  = \new_[25304]_  & \new_[25299]_ ;
  assign \new_[25309]_  = ~A266 & ~A265;
  assign \new_[25310]_  = ~A236 & \new_[25309]_ ;
  assign \new_[25314]_  = ~A302 & ~A301;
  assign \new_[25315]_  = A298 & \new_[25314]_ ;
  assign \new_[25316]_  = \new_[25315]_  & \new_[25310]_ ;
  assign \new_[25320]_  = ~A200 & A167;
  assign \new_[25321]_  = A168 & \new_[25320]_ ;
  assign \new_[25325]_  = ~A234 & ~A233;
  assign \new_[25326]_  = ~A201 & \new_[25325]_ ;
  assign \new_[25327]_  = \new_[25326]_  & \new_[25321]_ ;
  assign \new_[25331]_  = ~A269 & ~A268;
  assign \new_[25332]_  = ~A266 & \new_[25331]_ ;
  assign \new_[25336]_  = ~A302 & ~A301;
  assign \new_[25337]_  = A298 & \new_[25336]_ ;
  assign \new_[25338]_  = \new_[25337]_  & \new_[25332]_ ;
  assign \new_[25342]_  = ~A200 & A167;
  assign \new_[25343]_  = A168 & \new_[25342]_ ;
  assign \new_[25347]_  = ~A233 & A232;
  assign \new_[25348]_  = ~A201 & \new_[25347]_ ;
  assign \new_[25349]_  = \new_[25348]_  & \new_[25343]_ ;
  assign \new_[25353]_  = A298 & A235;
  assign \new_[25354]_  = A234 & \new_[25353]_ ;
  assign \new_[25358]_  = A301 & A300;
  assign \new_[25359]_  = ~A299 & \new_[25358]_ ;
  assign \new_[25360]_  = \new_[25359]_  & \new_[25354]_ ;
  assign \new_[25364]_  = ~A200 & A167;
  assign \new_[25365]_  = A168 & \new_[25364]_ ;
  assign \new_[25369]_  = ~A233 & A232;
  assign \new_[25370]_  = ~A201 & \new_[25369]_ ;
  assign \new_[25371]_  = \new_[25370]_  & \new_[25365]_ ;
  assign \new_[25375]_  = A298 & A235;
  assign \new_[25376]_  = A234 & \new_[25375]_ ;
  assign \new_[25380]_  = A302 & A300;
  assign \new_[25381]_  = ~A299 & \new_[25380]_ ;
  assign \new_[25382]_  = \new_[25381]_  & \new_[25376]_ ;
  assign \new_[25386]_  = ~A200 & A167;
  assign \new_[25387]_  = A168 & \new_[25386]_ ;
  assign \new_[25391]_  = ~A233 & A232;
  assign \new_[25392]_  = ~A201 & \new_[25391]_ ;
  assign \new_[25393]_  = \new_[25392]_  & \new_[25387]_ ;
  assign \new_[25397]_  = A265 & A235;
  assign \new_[25398]_  = A234 & \new_[25397]_ ;
  assign \new_[25402]_  = A268 & A267;
  assign \new_[25403]_  = ~A266 & \new_[25402]_ ;
  assign \new_[25404]_  = \new_[25403]_  & \new_[25398]_ ;
  assign \new_[25408]_  = ~A200 & A167;
  assign \new_[25409]_  = A168 & \new_[25408]_ ;
  assign \new_[25413]_  = ~A233 & A232;
  assign \new_[25414]_  = ~A201 & \new_[25413]_ ;
  assign \new_[25415]_  = \new_[25414]_  & \new_[25409]_ ;
  assign \new_[25419]_  = A265 & A235;
  assign \new_[25420]_  = A234 & \new_[25419]_ ;
  assign \new_[25424]_  = A269 & A267;
  assign \new_[25425]_  = ~A266 & \new_[25424]_ ;
  assign \new_[25426]_  = \new_[25425]_  & \new_[25420]_ ;
  assign \new_[25430]_  = ~A200 & A167;
  assign \new_[25431]_  = A168 & \new_[25430]_ ;
  assign \new_[25435]_  = ~A233 & A232;
  assign \new_[25436]_  = ~A201 & \new_[25435]_ ;
  assign \new_[25437]_  = \new_[25436]_  & \new_[25431]_ ;
  assign \new_[25441]_  = A298 & A236;
  assign \new_[25442]_  = A234 & \new_[25441]_ ;
  assign \new_[25446]_  = A301 & A300;
  assign \new_[25447]_  = ~A299 & \new_[25446]_ ;
  assign \new_[25448]_  = \new_[25447]_  & \new_[25442]_ ;
  assign \new_[25452]_  = ~A200 & A167;
  assign \new_[25453]_  = A168 & \new_[25452]_ ;
  assign \new_[25457]_  = ~A233 & A232;
  assign \new_[25458]_  = ~A201 & \new_[25457]_ ;
  assign \new_[25459]_  = \new_[25458]_  & \new_[25453]_ ;
  assign \new_[25463]_  = A298 & A236;
  assign \new_[25464]_  = A234 & \new_[25463]_ ;
  assign \new_[25468]_  = A302 & A300;
  assign \new_[25469]_  = ~A299 & \new_[25468]_ ;
  assign \new_[25470]_  = \new_[25469]_  & \new_[25464]_ ;
  assign \new_[25474]_  = ~A200 & A167;
  assign \new_[25475]_  = A168 & \new_[25474]_ ;
  assign \new_[25479]_  = ~A233 & A232;
  assign \new_[25480]_  = ~A201 & \new_[25479]_ ;
  assign \new_[25481]_  = \new_[25480]_  & \new_[25475]_ ;
  assign \new_[25485]_  = A265 & A236;
  assign \new_[25486]_  = A234 & \new_[25485]_ ;
  assign \new_[25490]_  = A268 & A267;
  assign \new_[25491]_  = ~A266 & \new_[25490]_ ;
  assign \new_[25492]_  = \new_[25491]_  & \new_[25486]_ ;
  assign \new_[25496]_  = ~A200 & A167;
  assign \new_[25497]_  = A168 & \new_[25496]_ ;
  assign \new_[25501]_  = ~A233 & A232;
  assign \new_[25502]_  = ~A201 & \new_[25501]_ ;
  assign \new_[25503]_  = \new_[25502]_  & \new_[25497]_ ;
  assign \new_[25507]_  = A265 & A236;
  assign \new_[25508]_  = A234 & \new_[25507]_ ;
  assign \new_[25512]_  = A269 & A267;
  assign \new_[25513]_  = ~A266 & \new_[25512]_ ;
  assign \new_[25514]_  = \new_[25513]_  & \new_[25508]_ ;
  assign \new_[25518]_  = ~A200 & A167;
  assign \new_[25519]_  = A168 & \new_[25518]_ ;
  assign \new_[25523]_  = ~A233 & ~A232;
  assign \new_[25524]_  = ~A201 & \new_[25523]_ ;
  assign \new_[25525]_  = \new_[25524]_  & \new_[25519]_ ;
  assign \new_[25529]_  = ~A269 & ~A268;
  assign \new_[25530]_  = ~A266 & \new_[25529]_ ;
  assign \new_[25534]_  = ~A302 & ~A301;
  assign \new_[25535]_  = A298 & \new_[25534]_ ;
  assign \new_[25536]_  = \new_[25535]_  & \new_[25530]_ ;
  assign \new_[25540]_  = ~A199 & A167;
  assign \new_[25541]_  = A168 & \new_[25540]_ ;
  assign \new_[25545]_  = A233 & A232;
  assign \new_[25546]_  = ~A200 & \new_[25545]_ ;
  assign \new_[25547]_  = \new_[25546]_  & \new_[25541]_ ;
  assign \new_[25551]_  = ~A269 & ~A268;
  assign \new_[25552]_  = A265 & \new_[25551]_ ;
  assign \new_[25556]_  = ~A302 & ~A301;
  assign \new_[25557]_  = ~A299 & \new_[25556]_ ;
  assign \new_[25558]_  = \new_[25557]_  & \new_[25552]_ ;
  assign \new_[25562]_  = ~A199 & A167;
  assign \new_[25563]_  = A168 & \new_[25562]_ ;
  assign \new_[25567]_  = ~A235 & ~A233;
  assign \new_[25568]_  = ~A200 & \new_[25567]_ ;
  assign \new_[25569]_  = \new_[25568]_  & \new_[25563]_ ;
  assign \new_[25573]_  = A266 & A265;
  assign \new_[25574]_  = ~A236 & \new_[25573]_ ;
  assign \new_[25578]_  = ~A302 & ~A301;
  assign \new_[25579]_  = A298 & \new_[25578]_ ;
  assign \new_[25580]_  = \new_[25579]_  & \new_[25574]_ ;
  assign \new_[25584]_  = ~A199 & A167;
  assign \new_[25585]_  = A168 & \new_[25584]_ ;
  assign \new_[25589]_  = ~A235 & ~A233;
  assign \new_[25590]_  = ~A200 & \new_[25589]_ ;
  assign \new_[25591]_  = \new_[25590]_  & \new_[25585]_ ;
  assign \new_[25595]_  = ~A268 & ~A266;
  assign \new_[25596]_  = ~A236 & \new_[25595]_ ;
  assign \new_[25600]_  = ~A300 & A298;
  assign \new_[25601]_  = ~A269 & \new_[25600]_ ;
  assign \new_[25602]_  = \new_[25601]_  & \new_[25596]_ ;
  assign \new_[25606]_  = ~A199 & A167;
  assign \new_[25607]_  = A168 & \new_[25606]_ ;
  assign \new_[25611]_  = ~A235 & ~A233;
  assign \new_[25612]_  = ~A200 & \new_[25611]_ ;
  assign \new_[25613]_  = \new_[25612]_  & \new_[25607]_ ;
  assign \new_[25617]_  = ~A268 & ~A266;
  assign \new_[25618]_  = ~A236 & \new_[25617]_ ;
  assign \new_[25622]_  = A299 & A298;
  assign \new_[25623]_  = ~A269 & \new_[25622]_ ;
  assign \new_[25624]_  = \new_[25623]_  & \new_[25618]_ ;
  assign \new_[25628]_  = ~A199 & A167;
  assign \new_[25629]_  = A168 & \new_[25628]_ ;
  assign \new_[25633]_  = ~A235 & ~A233;
  assign \new_[25634]_  = ~A200 & \new_[25633]_ ;
  assign \new_[25635]_  = \new_[25634]_  & \new_[25629]_ ;
  assign \new_[25639]_  = ~A268 & ~A266;
  assign \new_[25640]_  = ~A236 & \new_[25639]_ ;
  assign \new_[25644]_  = ~A299 & ~A298;
  assign \new_[25645]_  = ~A269 & \new_[25644]_ ;
  assign \new_[25646]_  = \new_[25645]_  & \new_[25640]_ ;
  assign \new_[25650]_  = ~A199 & A167;
  assign \new_[25651]_  = A168 & \new_[25650]_ ;
  assign \new_[25655]_  = ~A235 & ~A233;
  assign \new_[25656]_  = ~A200 & \new_[25655]_ ;
  assign \new_[25657]_  = \new_[25656]_  & \new_[25651]_ ;
  assign \new_[25661]_  = ~A267 & ~A266;
  assign \new_[25662]_  = ~A236 & \new_[25661]_ ;
  assign \new_[25666]_  = ~A302 & ~A301;
  assign \new_[25667]_  = A298 & \new_[25666]_ ;
  assign \new_[25668]_  = \new_[25667]_  & \new_[25662]_ ;
  assign \new_[25672]_  = ~A199 & A167;
  assign \new_[25673]_  = A168 & \new_[25672]_ ;
  assign \new_[25677]_  = ~A235 & ~A233;
  assign \new_[25678]_  = ~A200 & \new_[25677]_ ;
  assign \new_[25679]_  = \new_[25678]_  & \new_[25673]_ ;
  assign \new_[25683]_  = ~A266 & ~A265;
  assign \new_[25684]_  = ~A236 & \new_[25683]_ ;
  assign \new_[25688]_  = ~A302 & ~A301;
  assign \new_[25689]_  = A298 & \new_[25688]_ ;
  assign \new_[25690]_  = \new_[25689]_  & \new_[25684]_ ;
  assign \new_[25694]_  = ~A199 & A167;
  assign \new_[25695]_  = A168 & \new_[25694]_ ;
  assign \new_[25699]_  = ~A234 & ~A233;
  assign \new_[25700]_  = ~A200 & \new_[25699]_ ;
  assign \new_[25701]_  = \new_[25700]_  & \new_[25695]_ ;
  assign \new_[25705]_  = ~A269 & ~A268;
  assign \new_[25706]_  = ~A266 & \new_[25705]_ ;
  assign \new_[25710]_  = ~A302 & ~A301;
  assign \new_[25711]_  = A298 & \new_[25710]_ ;
  assign \new_[25712]_  = \new_[25711]_  & \new_[25706]_ ;
  assign \new_[25716]_  = ~A199 & A167;
  assign \new_[25717]_  = A168 & \new_[25716]_ ;
  assign \new_[25721]_  = ~A233 & A232;
  assign \new_[25722]_  = ~A200 & \new_[25721]_ ;
  assign \new_[25723]_  = \new_[25722]_  & \new_[25717]_ ;
  assign \new_[25727]_  = A298 & A235;
  assign \new_[25728]_  = A234 & \new_[25727]_ ;
  assign \new_[25732]_  = A301 & A300;
  assign \new_[25733]_  = ~A299 & \new_[25732]_ ;
  assign \new_[25734]_  = \new_[25733]_  & \new_[25728]_ ;
  assign \new_[25738]_  = ~A199 & A167;
  assign \new_[25739]_  = A168 & \new_[25738]_ ;
  assign \new_[25743]_  = ~A233 & A232;
  assign \new_[25744]_  = ~A200 & \new_[25743]_ ;
  assign \new_[25745]_  = \new_[25744]_  & \new_[25739]_ ;
  assign \new_[25749]_  = A298 & A235;
  assign \new_[25750]_  = A234 & \new_[25749]_ ;
  assign \new_[25754]_  = A302 & A300;
  assign \new_[25755]_  = ~A299 & \new_[25754]_ ;
  assign \new_[25756]_  = \new_[25755]_  & \new_[25750]_ ;
  assign \new_[25760]_  = ~A199 & A167;
  assign \new_[25761]_  = A168 & \new_[25760]_ ;
  assign \new_[25765]_  = ~A233 & A232;
  assign \new_[25766]_  = ~A200 & \new_[25765]_ ;
  assign \new_[25767]_  = \new_[25766]_  & \new_[25761]_ ;
  assign \new_[25771]_  = A265 & A235;
  assign \new_[25772]_  = A234 & \new_[25771]_ ;
  assign \new_[25776]_  = A268 & A267;
  assign \new_[25777]_  = ~A266 & \new_[25776]_ ;
  assign \new_[25778]_  = \new_[25777]_  & \new_[25772]_ ;
  assign \new_[25782]_  = ~A199 & A167;
  assign \new_[25783]_  = A168 & \new_[25782]_ ;
  assign \new_[25787]_  = ~A233 & A232;
  assign \new_[25788]_  = ~A200 & \new_[25787]_ ;
  assign \new_[25789]_  = \new_[25788]_  & \new_[25783]_ ;
  assign \new_[25793]_  = A265 & A235;
  assign \new_[25794]_  = A234 & \new_[25793]_ ;
  assign \new_[25798]_  = A269 & A267;
  assign \new_[25799]_  = ~A266 & \new_[25798]_ ;
  assign \new_[25800]_  = \new_[25799]_  & \new_[25794]_ ;
  assign \new_[25804]_  = ~A199 & A167;
  assign \new_[25805]_  = A168 & \new_[25804]_ ;
  assign \new_[25809]_  = ~A233 & A232;
  assign \new_[25810]_  = ~A200 & \new_[25809]_ ;
  assign \new_[25811]_  = \new_[25810]_  & \new_[25805]_ ;
  assign \new_[25815]_  = A298 & A236;
  assign \new_[25816]_  = A234 & \new_[25815]_ ;
  assign \new_[25820]_  = A301 & A300;
  assign \new_[25821]_  = ~A299 & \new_[25820]_ ;
  assign \new_[25822]_  = \new_[25821]_  & \new_[25816]_ ;
  assign \new_[25826]_  = ~A199 & A167;
  assign \new_[25827]_  = A168 & \new_[25826]_ ;
  assign \new_[25831]_  = ~A233 & A232;
  assign \new_[25832]_  = ~A200 & \new_[25831]_ ;
  assign \new_[25833]_  = \new_[25832]_  & \new_[25827]_ ;
  assign \new_[25837]_  = A298 & A236;
  assign \new_[25838]_  = A234 & \new_[25837]_ ;
  assign \new_[25842]_  = A302 & A300;
  assign \new_[25843]_  = ~A299 & \new_[25842]_ ;
  assign \new_[25844]_  = \new_[25843]_  & \new_[25838]_ ;
  assign \new_[25848]_  = ~A199 & A167;
  assign \new_[25849]_  = A168 & \new_[25848]_ ;
  assign \new_[25853]_  = ~A233 & A232;
  assign \new_[25854]_  = ~A200 & \new_[25853]_ ;
  assign \new_[25855]_  = \new_[25854]_  & \new_[25849]_ ;
  assign \new_[25859]_  = A265 & A236;
  assign \new_[25860]_  = A234 & \new_[25859]_ ;
  assign \new_[25864]_  = A268 & A267;
  assign \new_[25865]_  = ~A266 & \new_[25864]_ ;
  assign \new_[25866]_  = \new_[25865]_  & \new_[25860]_ ;
  assign \new_[25870]_  = ~A199 & A167;
  assign \new_[25871]_  = A168 & \new_[25870]_ ;
  assign \new_[25875]_  = ~A233 & A232;
  assign \new_[25876]_  = ~A200 & \new_[25875]_ ;
  assign \new_[25877]_  = \new_[25876]_  & \new_[25871]_ ;
  assign \new_[25881]_  = A265 & A236;
  assign \new_[25882]_  = A234 & \new_[25881]_ ;
  assign \new_[25886]_  = A269 & A267;
  assign \new_[25887]_  = ~A266 & \new_[25886]_ ;
  assign \new_[25888]_  = \new_[25887]_  & \new_[25882]_ ;
  assign \new_[25892]_  = ~A199 & A167;
  assign \new_[25893]_  = A168 & \new_[25892]_ ;
  assign \new_[25897]_  = ~A233 & ~A232;
  assign \new_[25898]_  = ~A200 & \new_[25897]_ ;
  assign \new_[25899]_  = \new_[25898]_  & \new_[25893]_ ;
  assign \new_[25903]_  = ~A269 & ~A268;
  assign \new_[25904]_  = ~A266 & \new_[25903]_ ;
  assign \new_[25908]_  = ~A302 & ~A301;
  assign \new_[25909]_  = A298 & \new_[25908]_ ;
  assign \new_[25910]_  = \new_[25909]_  & \new_[25904]_ ;
  assign \new_[25914]_  = ~A166 & ~A167;
  assign \new_[25915]_  = A170 & \new_[25914]_ ;
  assign \new_[25919]_  = A232 & A200;
  assign \new_[25920]_  = ~A199 & \new_[25919]_ ;
  assign \new_[25921]_  = \new_[25920]_  & \new_[25915]_ ;
  assign \new_[25925]_  = ~A268 & A265;
  assign \new_[25926]_  = A233 & \new_[25925]_ ;
  assign \new_[25930]_  = ~A300 & ~A299;
  assign \new_[25931]_  = ~A269 & \new_[25930]_ ;
  assign \new_[25932]_  = \new_[25931]_  & \new_[25926]_ ;
  assign \new_[25936]_  = ~A166 & ~A167;
  assign \new_[25937]_  = A170 & \new_[25936]_ ;
  assign \new_[25941]_  = A232 & A200;
  assign \new_[25942]_  = ~A199 & \new_[25941]_ ;
  assign \new_[25943]_  = \new_[25942]_  & \new_[25937]_ ;
  assign \new_[25947]_  = ~A268 & A265;
  assign \new_[25948]_  = A233 & \new_[25947]_ ;
  assign \new_[25952]_  = A299 & A298;
  assign \new_[25953]_  = ~A269 & \new_[25952]_ ;
  assign \new_[25954]_  = \new_[25953]_  & \new_[25948]_ ;
  assign \new_[25958]_  = ~A166 & ~A167;
  assign \new_[25959]_  = A170 & \new_[25958]_ ;
  assign \new_[25963]_  = A232 & A200;
  assign \new_[25964]_  = ~A199 & \new_[25963]_ ;
  assign \new_[25965]_  = \new_[25964]_  & \new_[25959]_ ;
  assign \new_[25969]_  = ~A268 & A265;
  assign \new_[25970]_  = A233 & \new_[25969]_ ;
  assign \new_[25974]_  = ~A299 & ~A298;
  assign \new_[25975]_  = ~A269 & \new_[25974]_ ;
  assign \new_[25976]_  = \new_[25975]_  & \new_[25970]_ ;
  assign \new_[25980]_  = ~A166 & ~A167;
  assign \new_[25981]_  = A170 & \new_[25980]_ ;
  assign \new_[25985]_  = A232 & A200;
  assign \new_[25986]_  = ~A199 & \new_[25985]_ ;
  assign \new_[25987]_  = \new_[25986]_  & \new_[25981]_ ;
  assign \new_[25991]_  = ~A267 & A265;
  assign \new_[25992]_  = A233 & \new_[25991]_ ;
  assign \new_[25996]_  = ~A302 & ~A301;
  assign \new_[25997]_  = ~A299 & \new_[25996]_ ;
  assign \new_[25998]_  = \new_[25997]_  & \new_[25992]_ ;
  assign \new_[26002]_  = ~A166 & ~A167;
  assign \new_[26003]_  = A170 & \new_[26002]_ ;
  assign \new_[26007]_  = A232 & A200;
  assign \new_[26008]_  = ~A199 & \new_[26007]_ ;
  assign \new_[26009]_  = \new_[26008]_  & \new_[26003]_ ;
  assign \new_[26013]_  = A266 & A265;
  assign \new_[26014]_  = A233 & \new_[26013]_ ;
  assign \new_[26018]_  = ~A302 & ~A301;
  assign \new_[26019]_  = ~A299 & \new_[26018]_ ;
  assign \new_[26020]_  = \new_[26019]_  & \new_[26014]_ ;
  assign \new_[26024]_  = ~A166 & ~A167;
  assign \new_[26025]_  = A170 & \new_[26024]_ ;
  assign \new_[26029]_  = A232 & A200;
  assign \new_[26030]_  = ~A199 & \new_[26029]_ ;
  assign \new_[26031]_  = \new_[26030]_  & \new_[26025]_ ;
  assign \new_[26035]_  = ~A266 & ~A265;
  assign \new_[26036]_  = A233 & \new_[26035]_ ;
  assign \new_[26040]_  = ~A302 & ~A301;
  assign \new_[26041]_  = ~A299 & \new_[26040]_ ;
  assign \new_[26042]_  = \new_[26041]_  & \new_[26036]_ ;
  assign \new_[26046]_  = ~A166 & ~A167;
  assign \new_[26047]_  = A170 & \new_[26046]_ ;
  assign \new_[26051]_  = ~A233 & A200;
  assign \new_[26052]_  = ~A199 & \new_[26051]_ ;
  assign \new_[26053]_  = \new_[26052]_  & \new_[26047]_ ;
  assign \new_[26057]_  = A265 & ~A236;
  assign \new_[26058]_  = ~A235 & \new_[26057]_ ;
  assign \new_[26062]_  = ~A300 & A298;
  assign \new_[26063]_  = A266 & \new_[26062]_ ;
  assign \new_[26064]_  = \new_[26063]_  & \new_[26058]_ ;
  assign \new_[26068]_  = ~A166 & ~A167;
  assign \new_[26069]_  = A170 & \new_[26068]_ ;
  assign \new_[26073]_  = ~A233 & A200;
  assign \new_[26074]_  = ~A199 & \new_[26073]_ ;
  assign \new_[26075]_  = \new_[26074]_  & \new_[26069]_ ;
  assign \new_[26079]_  = A265 & ~A236;
  assign \new_[26080]_  = ~A235 & \new_[26079]_ ;
  assign \new_[26084]_  = A299 & A298;
  assign \new_[26085]_  = A266 & \new_[26084]_ ;
  assign \new_[26086]_  = \new_[26085]_  & \new_[26080]_ ;
  assign \new_[26090]_  = ~A166 & ~A167;
  assign \new_[26091]_  = A170 & \new_[26090]_ ;
  assign \new_[26095]_  = ~A233 & A200;
  assign \new_[26096]_  = ~A199 & \new_[26095]_ ;
  assign \new_[26097]_  = \new_[26096]_  & \new_[26091]_ ;
  assign \new_[26101]_  = A265 & ~A236;
  assign \new_[26102]_  = ~A235 & \new_[26101]_ ;
  assign \new_[26106]_  = ~A299 & ~A298;
  assign \new_[26107]_  = A266 & \new_[26106]_ ;
  assign \new_[26108]_  = \new_[26107]_  & \new_[26102]_ ;
  assign \new_[26112]_  = ~A166 & ~A167;
  assign \new_[26113]_  = A170 & \new_[26112]_ ;
  assign \new_[26117]_  = ~A233 & A200;
  assign \new_[26118]_  = ~A199 & \new_[26117]_ ;
  assign \new_[26119]_  = \new_[26118]_  & \new_[26113]_ ;
  assign \new_[26123]_  = ~A266 & ~A236;
  assign \new_[26124]_  = ~A235 & \new_[26123]_ ;
  assign \new_[26128]_  = ~A300 & A298;
  assign \new_[26129]_  = ~A267 & \new_[26128]_ ;
  assign \new_[26130]_  = \new_[26129]_  & \new_[26124]_ ;
  assign \new_[26134]_  = ~A166 & ~A167;
  assign \new_[26135]_  = A170 & \new_[26134]_ ;
  assign \new_[26139]_  = ~A233 & A200;
  assign \new_[26140]_  = ~A199 & \new_[26139]_ ;
  assign \new_[26141]_  = \new_[26140]_  & \new_[26135]_ ;
  assign \new_[26145]_  = ~A266 & ~A236;
  assign \new_[26146]_  = ~A235 & \new_[26145]_ ;
  assign \new_[26150]_  = A299 & A298;
  assign \new_[26151]_  = ~A267 & \new_[26150]_ ;
  assign \new_[26152]_  = \new_[26151]_  & \new_[26146]_ ;
  assign \new_[26156]_  = ~A166 & ~A167;
  assign \new_[26157]_  = A170 & \new_[26156]_ ;
  assign \new_[26161]_  = ~A233 & A200;
  assign \new_[26162]_  = ~A199 & \new_[26161]_ ;
  assign \new_[26163]_  = \new_[26162]_  & \new_[26157]_ ;
  assign \new_[26167]_  = ~A266 & ~A236;
  assign \new_[26168]_  = ~A235 & \new_[26167]_ ;
  assign \new_[26172]_  = ~A299 & ~A298;
  assign \new_[26173]_  = ~A267 & \new_[26172]_ ;
  assign \new_[26174]_  = \new_[26173]_  & \new_[26168]_ ;
  assign \new_[26178]_  = ~A166 & ~A167;
  assign \new_[26179]_  = A170 & \new_[26178]_ ;
  assign \new_[26183]_  = ~A233 & A200;
  assign \new_[26184]_  = ~A199 & \new_[26183]_ ;
  assign \new_[26185]_  = \new_[26184]_  & \new_[26179]_ ;
  assign \new_[26189]_  = ~A265 & ~A236;
  assign \new_[26190]_  = ~A235 & \new_[26189]_ ;
  assign \new_[26194]_  = ~A300 & A298;
  assign \new_[26195]_  = ~A266 & \new_[26194]_ ;
  assign \new_[26196]_  = \new_[26195]_  & \new_[26190]_ ;
  assign \new_[26200]_  = ~A166 & ~A167;
  assign \new_[26201]_  = A170 & \new_[26200]_ ;
  assign \new_[26205]_  = ~A233 & A200;
  assign \new_[26206]_  = ~A199 & \new_[26205]_ ;
  assign \new_[26207]_  = \new_[26206]_  & \new_[26201]_ ;
  assign \new_[26211]_  = ~A265 & ~A236;
  assign \new_[26212]_  = ~A235 & \new_[26211]_ ;
  assign \new_[26216]_  = A299 & A298;
  assign \new_[26217]_  = ~A266 & \new_[26216]_ ;
  assign \new_[26218]_  = \new_[26217]_  & \new_[26212]_ ;
  assign \new_[26222]_  = ~A166 & ~A167;
  assign \new_[26223]_  = A170 & \new_[26222]_ ;
  assign \new_[26227]_  = ~A233 & A200;
  assign \new_[26228]_  = ~A199 & \new_[26227]_ ;
  assign \new_[26229]_  = \new_[26228]_  & \new_[26223]_ ;
  assign \new_[26233]_  = ~A265 & ~A236;
  assign \new_[26234]_  = ~A235 & \new_[26233]_ ;
  assign \new_[26238]_  = ~A299 & ~A298;
  assign \new_[26239]_  = ~A266 & \new_[26238]_ ;
  assign \new_[26240]_  = \new_[26239]_  & \new_[26234]_ ;
  assign \new_[26244]_  = ~A166 & ~A167;
  assign \new_[26245]_  = A170 & \new_[26244]_ ;
  assign \new_[26249]_  = ~A233 & A200;
  assign \new_[26250]_  = ~A199 & \new_[26249]_ ;
  assign \new_[26251]_  = \new_[26250]_  & \new_[26245]_ ;
  assign \new_[26255]_  = A266 & A265;
  assign \new_[26256]_  = ~A234 & \new_[26255]_ ;
  assign \new_[26260]_  = ~A302 & ~A301;
  assign \new_[26261]_  = A298 & \new_[26260]_ ;
  assign \new_[26262]_  = \new_[26261]_  & \new_[26256]_ ;
  assign \new_[26266]_  = ~A166 & ~A167;
  assign \new_[26267]_  = A170 & \new_[26266]_ ;
  assign \new_[26271]_  = ~A233 & A200;
  assign \new_[26272]_  = ~A199 & \new_[26271]_ ;
  assign \new_[26273]_  = \new_[26272]_  & \new_[26267]_ ;
  assign \new_[26277]_  = ~A268 & ~A266;
  assign \new_[26278]_  = ~A234 & \new_[26277]_ ;
  assign \new_[26282]_  = ~A300 & A298;
  assign \new_[26283]_  = ~A269 & \new_[26282]_ ;
  assign \new_[26284]_  = \new_[26283]_  & \new_[26278]_ ;
  assign \new_[26288]_  = ~A166 & ~A167;
  assign \new_[26289]_  = A170 & \new_[26288]_ ;
  assign \new_[26293]_  = ~A233 & A200;
  assign \new_[26294]_  = ~A199 & \new_[26293]_ ;
  assign \new_[26295]_  = \new_[26294]_  & \new_[26289]_ ;
  assign \new_[26299]_  = ~A268 & ~A266;
  assign \new_[26300]_  = ~A234 & \new_[26299]_ ;
  assign \new_[26304]_  = A299 & A298;
  assign \new_[26305]_  = ~A269 & \new_[26304]_ ;
  assign \new_[26306]_  = \new_[26305]_  & \new_[26300]_ ;
  assign \new_[26310]_  = ~A166 & ~A167;
  assign \new_[26311]_  = A170 & \new_[26310]_ ;
  assign \new_[26315]_  = ~A233 & A200;
  assign \new_[26316]_  = ~A199 & \new_[26315]_ ;
  assign \new_[26317]_  = \new_[26316]_  & \new_[26311]_ ;
  assign \new_[26321]_  = ~A268 & ~A266;
  assign \new_[26322]_  = ~A234 & \new_[26321]_ ;
  assign \new_[26326]_  = ~A299 & ~A298;
  assign \new_[26327]_  = ~A269 & \new_[26326]_ ;
  assign \new_[26328]_  = \new_[26327]_  & \new_[26322]_ ;
  assign \new_[26332]_  = ~A166 & ~A167;
  assign \new_[26333]_  = A170 & \new_[26332]_ ;
  assign \new_[26337]_  = ~A233 & A200;
  assign \new_[26338]_  = ~A199 & \new_[26337]_ ;
  assign \new_[26339]_  = \new_[26338]_  & \new_[26333]_ ;
  assign \new_[26343]_  = ~A267 & ~A266;
  assign \new_[26344]_  = ~A234 & \new_[26343]_ ;
  assign \new_[26348]_  = ~A302 & ~A301;
  assign \new_[26349]_  = A298 & \new_[26348]_ ;
  assign \new_[26350]_  = \new_[26349]_  & \new_[26344]_ ;
  assign \new_[26354]_  = ~A166 & ~A167;
  assign \new_[26355]_  = A170 & \new_[26354]_ ;
  assign \new_[26359]_  = ~A233 & A200;
  assign \new_[26360]_  = ~A199 & \new_[26359]_ ;
  assign \new_[26361]_  = \new_[26360]_  & \new_[26355]_ ;
  assign \new_[26365]_  = ~A266 & ~A265;
  assign \new_[26366]_  = ~A234 & \new_[26365]_ ;
  assign \new_[26370]_  = ~A302 & ~A301;
  assign \new_[26371]_  = A298 & \new_[26370]_ ;
  assign \new_[26372]_  = \new_[26371]_  & \new_[26366]_ ;
  assign \new_[26376]_  = ~A166 & ~A167;
  assign \new_[26377]_  = A170 & \new_[26376]_ ;
  assign \new_[26381]_  = ~A232 & A200;
  assign \new_[26382]_  = ~A199 & \new_[26381]_ ;
  assign \new_[26383]_  = \new_[26382]_  & \new_[26377]_ ;
  assign \new_[26387]_  = A266 & A265;
  assign \new_[26388]_  = ~A233 & \new_[26387]_ ;
  assign \new_[26392]_  = ~A302 & ~A301;
  assign \new_[26393]_  = A298 & \new_[26392]_ ;
  assign \new_[26394]_  = \new_[26393]_  & \new_[26388]_ ;
  assign \new_[26398]_  = ~A166 & ~A167;
  assign \new_[26399]_  = A170 & \new_[26398]_ ;
  assign \new_[26403]_  = ~A232 & A200;
  assign \new_[26404]_  = ~A199 & \new_[26403]_ ;
  assign \new_[26405]_  = \new_[26404]_  & \new_[26399]_ ;
  assign \new_[26409]_  = ~A268 & ~A266;
  assign \new_[26410]_  = ~A233 & \new_[26409]_ ;
  assign \new_[26414]_  = ~A300 & A298;
  assign \new_[26415]_  = ~A269 & \new_[26414]_ ;
  assign \new_[26416]_  = \new_[26415]_  & \new_[26410]_ ;
  assign \new_[26420]_  = ~A166 & ~A167;
  assign \new_[26421]_  = A170 & \new_[26420]_ ;
  assign \new_[26425]_  = ~A232 & A200;
  assign \new_[26426]_  = ~A199 & \new_[26425]_ ;
  assign \new_[26427]_  = \new_[26426]_  & \new_[26421]_ ;
  assign \new_[26431]_  = ~A268 & ~A266;
  assign \new_[26432]_  = ~A233 & \new_[26431]_ ;
  assign \new_[26436]_  = A299 & A298;
  assign \new_[26437]_  = ~A269 & \new_[26436]_ ;
  assign \new_[26438]_  = \new_[26437]_  & \new_[26432]_ ;
  assign \new_[26442]_  = ~A166 & ~A167;
  assign \new_[26443]_  = A170 & \new_[26442]_ ;
  assign \new_[26447]_  = ~A232 & A200;
  assign \new_[26448]_  = ~A199 & \new_[26447]_ ;
  assign \new_[26449]_  = \new_[26448]_  & \new_[26443]_ ;
  assign \new_[26453]_  = ~A268 & ~A266;
  assign \new_[26454]_  = ~A233 & \new_[26453]_ ;
  assign \new_[26458]_  = ~A299 & ~A298;
  assign \new_[26459]_  = ~A269 & \new_[26458]_ ;
  assign \new_[26460]_  = \new_[26459]_  & \new_[26454]_ ;
  assign \new_[26464]_  = ~A166 & ~A167;
  assign \new_[26465]_  = A170 & \new_[26464]_ ;
  assign \new_[26469]_  = ~A232 & A200;
  assign \new_[26470]_  = ~A199 & \new_[26469]_ ;
  assign \new_[26471]_  = \new_[26470]_  & \new_[26465]_ ;
  assign \new_[26475]_  = ~A267 & ~A266;
  assign \new_[26476]_  = ~A233 & \new_[26475]_ ;
  assign \new_[26480]_  = ~A302 & ~A301;
  assign \new_[26481]_  = A298 & \new_[26480]_ ;
  assign \new_[26482]_  = \new_[26481]_  & \new_[26476]_ ;
  assign \new_[26486]_  = ~A166 & ~A167;
  assign \new_[26487]_  = A170 & \new_[26486]_ ;
  assign \new_[26491]_  = ~A232 & A200;
  assign \new_[26492]_  = ~A199 & \new_[26491]_ ;
  assign \new_[26493]_  = \new_[26492]_  & \new_[26487]_ ;
  assign \new_[26497]_  = ~A266 & ~A265;
  assign \new_[26498]_  = ~A233 & \new_[26497]_ ;
  assign \new_[26502]_  = ~A302 & ~A301;
  assign \new_[26503]_  = A298 & \new_[26502]_ ;
  assign \new_[26504]_  = \new_[26503]_  & \new_[26498]_ ;
  assign \new_[26508]_  = A167 & ~A168;
  assign \new_[26509]_  = A170 & \new_[26508]_ ;
  assign \new_[26513]_  = A200 & ~A199;
  assign \new_[26514]_  = A166 & \new_[26513]_ ;
  assign \new_[26515]_  = \new_[26514]_  & \new_[26509]_ ;
  assign \new_[26519]_  = A265 & A233;
  assign \new_[26520]_  = A232 & \new_[26519]_ ;
  assign \new_[26524]_  = ~A300 & ~A299;
  assign \new_[26525]_  = ~A267 & \new_[26524]_ ;
  assign \new_[26526]_  = \new_[26525]_  & \new_[26520]_ ;
  assign \new_[26530]_  = A167 & ~A168;
  assign \new_[26531]_  = A170 & \new_[26530]_ ;
  assign \new_[26535]_  = A200 & ~A199;
  assign \new_[26536]_  = A166 & \new_[26535]_ ;
  assign \new_[26537]_  = \new_[26536]_  & \new_[26531]_ ;
  assign \new_[26541]_  = A265 & A233;
  assign \new_[26542]_  = A232 & \new_[26541]_ ;
  assign \new_[26546]_  = A299 & A298;
  assign \new_[26547]_  = ~A267 & \new_[26546]_ ;
  assign \new_[26548]_  = \new_[26547]_  & \new_[26542]_ ;
  assign \new_[26552]_  = A167 & ~A168;
  assign \new_[26553]_  = A170 & \new_[26552]_ ;
  assign \new_[26557]_  = A200 & ~A199;
  assign \new_[26558]_  = A166 & \new_[26557]_ ;
  assign \new_[26559]_  = \new_[26558]_  & \new_[26553]_ ;
  assign \new_[26563]_  = A265 & A233;
  assign \new_[26564]_  = A232 & \new_[26563]_ ;
  assign \new_[26568]_  = ~A299 & ~A298;
  assign \new_[26569]_  = ~A267 & \new_[26568]_ ;
  assign \new_[26570]_  = \new_[26569]_  & \new_[26564]_ ;
  assign \new_[26574]_  = A167 & ~A168;
  assign \new_[26575]_  = A170 & \new_[26574]_ ;
  assign \new_[26579]_  = A200 & ~A199;
  assign \new_[26580]_  = A166 & \new_[26579]_ ;
  assign \new_[26581]_  = \new_[26580]_  & \new_[26575]_ ;
  assign \new_[26585]_  = A265 & A233;
  assign \new_[26586]_  = A232 & \new_[26585]_ ;
  assign \new_[26590]_  = ~A300 & ~A299;
  assign \new_[26591]_  = A266 & \new_[26590]_ ;
  assign \new_[26592]_  = \new_[26591]_  & \new_[26586]_ ;
  assign \new_[26596]_  = A167 & ~A168;
  assign \new_[26597]_  = A170 & \new_[26596]_ ;
  assign \new_[26601]_  = A200 & ~A199;
  assign \new_[26602]_  = A166 & \new_[26601]_ ;
  assign \new_[26603]_  = \new_[26602]_  & \new_[26597]_ ;
  assign \new_[26607]_  = A265 & A233;
  assign \new_[26608]_  = A232 & \new_[26607]_ ;
  assign \new_[26612]_  = A299 & A298;
  assign \new_[26613]_  = A266 & \new_[26612]_ ;
  assign \new_[26614]_  = \new_[26613]_  & \new_[26608]_ ;
  assign \new_[26618]_  = A167 & ~A168;
  assign \new_[26619]_  = A170 & \new_[26618]_ ;
  assign \new_[26623]_  = A200 & ~A199;
  assign \new_[26624]_  = A166 & \new_[26623]_ ;
  assign \new_[26625]_  = \new_[26624]_  & \new_[26619]_ ;
  assign \new_[26629]_  = A265 & A233;
  assign \new_[26630]_  = A232 & \new_[26629]_ ;
  assign \new_[26634]_  = ~A299 & ~A298;
  assign \new_[26635]_  = A266 & \new_[26634]_ ;
  assign \new_[26636]_  = \new_[26635]_  & \new_[26630]_ ;
  assign \new_[26640]_  = A167 & ~A168;
  assign \new_[26641]_  = A170 & \new_[26640]_ ;
  assign \new_[26645]_  = A200 & ~A199;
  assign \new_[26646]_  = A166 & \new_[26645]_ ;
  assign \new_[26647]_  = \new_[26646]_  & \new_[26641]_ ;
  assign \new_[26651]_  = ~A265 & A233;
  assign \new_[26652]_  = A232 & \new_[26651]_ ;
  assign \new_[26656]_  = ~A300 & ~A299;
  assign \new_[26657]_  = ~A266 & \new_[26656]_ ;
  assign \new_[26658]_  = \new_[26657]_  & \new_[26652]_ ;
  assign \new_[26662]_  = A167 & ~A168;
  assign \new_[26663]_  = A170 & \new_[26662]_ ;
  assign \new_[26667]_  = A200 & ~A199;
  assign \new_[26668]_  = A166 & \new_[26667]_ ;
  assign \new_[26669]_  = \new_[26668]_  & \new_[26663]_ ;
  assign \new_[26673]_  = ~A265 & A233;
  assign \new_[26674]_  = A232 & \new_[26673]_ ;
  assign \new_[26678]_  = A299 & A298;
  assign \new_[26679]_  = ~A266 & \new_[26678]_ ;
  assign \new_[26680]_  = \new_[26679]_  & \new_[26674]_ ;
  assign \new_[26684]_  = A167 & ~A168;
  assign \new_[26685]_  = A170 & \new_[26684]_ ;
  assign \new_[26689]_  = A200 & ~A199;
  assign \new_[26690]_  = A166 & \new_[26689]_ ;
  assign \new_[26691]_  = \new_[26690]_  & \new_[26685]_ ;
  assign \new_[26695]_  = ~A265 & A233;
  assign \new_[26696]_  = A232 & \new_[26695]_ ;
  assign \new_[26700]_  = ~A299 & ~A298;
  assign \new_[26701]_  = ~A266 & \new_[26700]_ ;
  assign \new_[26702]_  = \new_[26701]_  & \new_[26696]_ ;
  assign \new_[26706]_  = A167 & ~A168;
  assign \new_[26707]_  = A170 & \new_[26706]_ ;
  assign \new_[26711]_  = A200 & ~A199;
  assign \new_[26712]_  = A166 & \new_[26711]_ ;
  assign \new_[26713]_  = \new_[26712]_  & \new_[26707]_ ;
  assign \new_[26717]_  = A298 & A233;
  assign \new_[26718]_  = ~A232 & \new_[26717]_ ;
  assign \new_[26722]_  = A301 & A300;
  assign \new_[26723]_  = ~A299 & \new_[26722]_ ;
  assign \new_[26724]_  = \new_[26723]_  & \new_[26718]_ ;
  assign \new_[26728]_  = A167 & ~A168;
  assign \new_[26729]_  = A170 & \new_[26728]_ ;
  assign \new_[26733]_  = A200 & ~A199;
  assign \new_[26734]_  = A166 & \new_[26733]_ ;
  assign \new_[26735]_  = \new_[26734]_  & \new_[26729]_ ;
  assign \new_[26739]_  = A298 & A233;
  assign \new_[26740]_  = ~A232 & \new_[26739]_ ;
  assign \new_[26744]_  = A302 & A300;
  assign \new_[26745]_  = ~A299 & \new_[26744]_ ;
  assign \new_[26746]_  = \new_[26745]_  & \new_[26740]_ ;
  assign \new_[26750]_  = A167 & ~A168;
  assign \new_[26751]_  = A170 & \new_[26750]_ ;
  assign \new_[26755]_  = A200 & ~A199;
  assign \new_[26756]_  = A166 & \new_[26755]_ ;
  assign \new_[26757]_  = \new_[26756]_  & \new_[26751]_ ;
  assign \new_[26761]_  = A265 & A233;
  assign \new_[26762]_  = ~A232 & \new_[26761]_ ;
  assign \new_[26766]_  = A268 & A267;
  assign \new_[26767]_  = ~A266 & \new_[26766]_ ;
  assign \new_[26768]_  = \new_[26767]_  & \new_[26762]_ ;
  assign \new_[26772]_  = A167 & ~A168;
  assign \new_[26773]_  = A170 & \new_[26772]_ ;
  assign \new_[26777]_  = A200 & ~A199;
  assign \new_[26778]_  = A166 & \new_[26777]_ ;
  assign \new_[26779]_  = \new_[26778]_  & \new_[26773]_ ;
  assign \new_[26783]_  = A265 & A233;
  assign \new_[26784]_  = ~A232 & \new_[26783]_ ;
  assign \new_[26788]_  = A269 & A267;
  assign \new_[26789]_  = ~A266 & \new_[26788]_ ;
  assign \new_[26790]_  = \new_[26789]_  & \new_[26784]_ ;
  assign \new_[26794]_  = A167 & ~A168;
  assign \new_[26795]_  = A170 & \new_[26794]_ ;
  assign \new_[26799]_  = A200 & ~A199;
  assign \new_[26800]_  = A166 & \new_[26799]_ ;
  assign \new_[26801]_  = \new_[26800]_  & \new_[26795]_ ;
  assign \new_[26805]_  = A265 & ~A234;
  assign \new_[26806]_  = ~A233 & \new_[26805]_ ;
  assign \new_[26810]_  = ~A300 & A298;
  assign \new_[26811]_  = A266 & \new_[26810]_ ;
  assign \new_[26812]_  = \new_[26811]_  & \new_[26806]_ ;
  assign \new_[26816]_  = A167 & ~A168;
  assign \new_[26817]_  = A170 & \new_[26816]_ ;
  assign \new_[26821]_  = A200 & ~A199;
  assign \new_[26822]_  = A166 & \new_[26821]_ ;
  assign \new_[26823]_  = \new_[26822]_  & \new_[26817]_ ;
  assign \new_[26827]_  = A265 & ~A234;
  assign \new_[26828]_  = ~A233 & \new_[26827]_ ;
  assign \new_[26832]_  = A299 & A298;
  assign \new_[26833]_  = A266 & \new_[26832]_ ;
  assign \new_[26834]_  = \new_[26833]_  & \new_[26828]_ ;
  assign \new_[26838]_  = A167 & ~A168;
  assign \new_[26839]_  = A170 & \new_[26838]_ ;
  assign \new_[26843]_  = A200 & ~A199;
  assign \new_[26844]_  = A166 & \new_[26843]_ ;
  assign \new_[26845]_  = \new_[26844]_  & \new_[26839]_ ;
  assign \new_[26849]_  = A265 & ~A234;
  assign \new_[26850]_  = ~A233 & \new_[26849]_ ;
  assign \new_[26854]_  = ~A299 & ~A298;
  assign \new_[26855]_  = A266 & \new_[26854]_ ;
  assign \new_[26856]_  = \new_[26855]_  & \new_[26850]_ ;
  assign \new_[26860]_  = A167 & ~A168;
  assign \new_[26861]_  = A170 & \new_[26860]_ ;
  assign \new_[26865]_  = A200 & ~A199;
  assign \new_[26866]_  = A166 & \new_[26865]_ ;
  assign \new_[26867]_  = \new_[26866]_  & \new_[26861]_ ;
  assign \new_[26871]_  = ~A266 & ~A234;
  assign \new_[26872]_  = ~A233 & \new_[26871]_ ;
  assign \new_[26876]_  = ~A300 & A298;
  assign \new_[26877]_  = ~A267 & \new_[26876]_ ;
  assign \new_[26878]_  = \new_[26877]_  & \new_[26872]_ ;
  assign \new_[26882]_  = A167 & ~A168;
  assign \new_[26883]_  = A170 & \new_[26882]_ ;
  assign \new_[26887]_  = A200 & ~A199;
  assign \new_[26888]_  = A166 & \new_[26887]_ ;
  assign \new_[26889]_  = \new_[26888]_  & \new_[26883]_ ;
  assign \new_[26893]_  = ~A266 & ~A234;
  assign \new_[26894]_  = ~A233 & \new_[26893]_ ;
  assign \new_[26898]_  = A299 & A298;
  assign \new_[26899]_  = ~A267 & \new_[26898]_ ;
  assign \new_[26900]_  = \new_[26899]_  & \new_[26894]_ ;
  assign \new_[26904]_  = A167 & ~A168;
  assign \new_[26905]_  = A170 & \new_[26904]_ ;
  assign \new_[26909]_  = A200 & ~A199;
  assign \new_[26910]_  = A166 & \new_[26909]_ ;
  assign \new_[26911]_  = \new_[26910]_  & \new_[26905]_ ;
  assign \new_[26915]_  = ~A266 & ~A234;
  assign \new_[26916]_  = ~A233 & \new_[26915]_ ;
  assign \new_[26920]_  = ~A299 & ~A298;
  assign \new_[26921]_  = ~A267 & \new_[26920]_ ;
  assign \new_[26922]_  = \new_[26921]_  & \new_[26916]_ ;
  assign \new_[26926]_  = A167 & ~A168;
  assign \new_[26927]_  = A170 & \new_[26926]_ ;
  assign \new_[26931]_  = A200 & ~A199;
  assign \new_[26932]_  = A166 & \new_[26931]_ ;
  assign \new_[26933]_  = \new_[26932]_  & \new_[26927]_ ;
  assign \new_[26937]_  = ~A265 & ~A234;
  assign \new_[26938]_  = ~A233 & \new_[26937]_ ;
  assign \new_[26942]_  = ~A300 & A298;
  assign \new_[26943]_  = ~A266 & \new_[26942]_ ;
  assign \new_[26944]_  = \new_[26943]_  & \new_[26938]_ ;
  assign \new_[26948]_  = A167 & ~A168;
  assign \new_[26949]_  = A170 & \new_[26948]_ ;
  assign \new_[26953]_  = A200 & ~A199;
  assign \new_[26954]_  = A166 & \new_[26953]_ ;
  assign \new_[26955]_  = \new_[26954]_  & \new_[26949]_ ;
  assign \new_[26959]_  = ~A265 & ~A234;
  assign \new_[26960]_  = ~A233 & \new_[26959]_ ;
  assign \new_[26964]_  = A299 & A298;
  assign \new_[26965]_  = ~A266 & \new_[26964]_ ;
  assign \new_[26966]_  = \new_[26965]_  & \new_[26960]_ ;
  assign \new_[26970]_  = A167 & ~A168;
  assign \new_[26971]_  = A170 & \new_[26970]_ ;
  assign \new_[26975]_  = A200 & ~A199;
  assign \new_[26976]_  = A166 & \new_[26975]_ ;
  assign \new_[26977]_  = \new_[26976]_  & \new_[26971]_ ;
  assign \new_[26981]_  = ~A265 & ~A234;
  assign \new_[26982]_  = ~A233 & \new_[26981]_ ;
  assign \new_[26986]_  = ~A299 & ~A298;
  assign \new_[26987]_  = ~A266 & \new_[26986]_ ;
  assign \new_[26988]_  = \new_[26987]_  & \new_[26982]_ ;
  assign \new_[26992]_  = A167 & ~A168;
  assign \new_[26993]_  = A170 & \new_[26992]_ ;
  assign \new_[26997]_  = A200 & ~A199;
  assign \new_[26998]_  = A166 & \new_[26997]_ ;
  assign \new_[26999]_  = \new_[26998]_  & \new_[26993]_ ;
  assign \new_[27003]_  = A234 & ~A233;
  assign \new_[27004]_  = A232 & \new_[27003]_ ;
  assign \new_[27008]_  = A299 & ~A298;
  assign \new_[27009]_  = A235 & \new_[27008]_ ;
  assign \new_[27010]_  = \new_[27009]_  & \new_[27004]_ ;
  assign \new_[27014]_  = A167 & ~A168;
  assign \new_[27015]_  = A170 & \new_[27014]_ ;
  assign \new_[27019]_  = A200 & ~A199;
  assign \new_[27020]_  = A166 & \new_[27019]_ ;
  assign \new_[27021]_  = \new_[27020]_  & \new_[27015]_ ;
  assign \new_[27025]_  = A234 & ~A233;
  assign \new_[27026]_  = A232 & \new_[27025]_ ;
  assign \new_[27030]_  = A266 & ~A265;
  assign \new_[27031]_  = A235 & \new_[27030]_ ;
  assign \new_[27032]_  = \new_[27031]_  & \new_[27026]_ ;
  assign \new_[27036]_  = A167 & ~A168;
  assign \new_[27037]_  = A170 & \new_[27036]_ ;
  assign \new_[27041]_  = A200 & ~A199;
  assign \new_[27042]_  = A166 & \new_[27041]_ ;
  assign \new_[27043]_  = \new_[27042]_  & \new_[27037]_ ;
  assign \new_[27047]_  = A234 & ~A233;
  assign \new_[27048]_  = A232 & \new_[27047]_ ;
  assign \new_[27052]_  = A299 & ~A298;
  assign \new_[27053]_  = A236 & \new_[27052]_ ;
  assign \new_[27054]_  = \new_[27053]_  & \new_[27048]_ ;
  assign \new_[27058]_  = A167 & ~A168;
  assign \new_[27059]_  = A170 & \new_[27058]_ ;
  assign \new_[27063]_  = A200 & ~A199;
  assign \new_[27064]_  = A166 & \new_[27063]_ ;
  assign \new_[27065]_  = \new_[27064]_  & \new_[27059]_ ;
  assign \new_[27069]_  = A234 & ~A233;
  assign \new_[27070]_  = A232 & \new_[27069]_ ;
  assign \new_[27074]_  = A266 & ~A265;
  assign \new_[27075]_  = A236 & \new_[27074]_ ;
  assign \new_[27076]_  = \new_[27075]_  & \new_[27070]_ ;
  assign \new_[27080]_  = A167 & ~A168;
  assign \new_[27081]_  = A170 & \new_[27080]_ ;
  assign \new_[27085]_  = A200 & ~A199;
  assign \new_[27086]_  = A166 & \new_[27085]_ ;
  assign \new_[27087]_  = \new_[27086]_  & \new_[27081]_ ;
  assign \new_[27091]_  = A265 & ~A233;
  assign \new_[27092]_  = ~A232 & \new_[27091]_ ;
  assign \new_[27096]_  = ~A300 & A298;
  assign \new_[27097]_  = A266 & \new_[27096]_ ;
  assign \new_[27098]_  = \new_[27097]_  & \new_[27092]_ ;
  assign \new_[27102]_  = A167 & ~A168;
  assign \new_[27103]_  = A170 & \new_[27102]_ ;
  assign \new_[27107]_  = A200 & ~A199;
  assign \new_[27108]_  = A166 & \new_[27107]_ ;
  assign \new_[27109]_  = \new_[27108]_  & \new_[27103]_ ;
  assign \new_[27113]_  = A265 & ~A233;
  assign \new_[27114]_  = ~A232 & \new_[27113]_ ;
  assign \new_[27118]_  = A299 & A298;
  assign \new_[27119]_  = A266 & \new_[27118]_ ;
  assign \new_[27120]_  = \new_[27119]_  & \new_[27114]_ ;
  assign \new_[27124]_  = A167 & ~A168;
  assign \new_[27125]_  = A170 & \new_[27124]_ ;
  assign \new_[27129]_  = A200 & ~A199;
  assign \new_[27130]_  = A166 & \new_[27129]_ ;
  assign \new_[27131]_  = \new_[27130]_  & \new_[27125]_ ;
  assign \new_[27135]_  = A265 & ~A233;
  assign \new_[27136]_  = ~A232 & \new_[27135]_ ;
  assign \new_[27140]_  = ~A299 & ~A298;
  assign \new_[27141]_  = A266 & \new_[27140]_ ;
  assign \new_[27142]_  = \new_[27141]_  & \new_[27136]_ ;
  assign \new_[27146]_  = A167 & ~A168;
  assign \new_[27147]_  = A170 & \new_[27146]_ ;
  assign \new_[27151]_  = A200 & ~A199;
  assign \new_[27152]_  = A166 & \new_[27151]_ ;
  assign \new_[27153]_  = \new_[27152]_  & \new_[27147]_ ;
  assign \new_[27157]_  = ~A266 & ~A233;
  assign \new_[27158]_  = ~A232 & \new_[27157]_ ;
  assign \new_[27162]_  = ~A300 & A298;
  assign \new_[27163]_  = ~A267 & \new_[27162]_ ;
  assign \new_[27164]_  = \new_[27163]_  & \new_[27158]_ ;
  assign \new_[27168]_  = A167 & ~A168;
  assign \new_[27169]_  = A170 & \new_[27168]_ ;
  assign \new_[27173]_  = A200 & ~A199;
  assign \new_[27174]_  = A166 & \new_[27173]_ ;
  assign \new_[27175]_  = \new_[27174]_  & \new_[27169]_ ;
  assign \new_[27179]_  = ~A266 & ~A233;
  assign \new_[27180]_  = ~A232 & \new_[27179]_ ;
  assign \new_[27184]_  = A299 & A298;
  assign \new_[27185]_  = ~A267 & \new_[27184]_ ;
  assign \new_[27186]_  = \new_[27185]_  & \new_[27180]_ ;
  assign \new_[27190]_  = A167 & ~A168;
  assign \new_[27191]_  = A170 & \new_[27190]_ ;
  assign \new_[27195]_  = A200 & ~A199;
  assign \new_[27196]_  = A166 & \new_[27195]_ ;
  assign \new_[27197]_  = \new_[27196]_  & \new_[27191]_ ;
  assign \new_[27201]_  = ~A266 & ~A233;
  assign \new_[27202]_  = ~A232 & \new_[27201]_ ;
  assign \new_[27206]_  = ~A299 & ~A298;
  assign \new_[27207]_  = ~A267 & \new_[27206]_ ;
  assign \new_[27208]_  = \new_[27207]_  & \new_[27202]_ ;
  assign \new_[27212]_  = A167 & ~A168;
  assign \new_[27213]_  = A170 & \new_[27212]_ ;
  assign \new_[27217]_  = A200 & ~A199;
  assign \new_[27218]_  = A166 & \new_[27217]_ ;
  assign \new_[27219]_  = \new_[27218]_  & \new_[27213]_ ;
  assign \new_[27223]_  = ~A265 & ~A233;
  assign \new_[27224]_  = ~A232 & \new_[27223]_ ;
  assign \new_[27228]_  = ~A300 & A298;
  assign \new_[27229]_  = ~A266 & \new_[27228]_ ;
  assign \new_[27230]_  = \new_[27229]_  & \new_[27224]_ ;
  assign \new_[27234]_  = A167 & ~A168;
  assign \new_[27235]_  = A170 & \new_[27234]_ ;
  assign \new_[27239]_  = A200 & ~A199;
  assign \new_[27240]_  = A166 & \new_[27239]_ ;
  assign \new_[27241]_  = \new_[27240]_  & \new_[27235]_ ;
  assign \new_[27245]_  = ~A265 & ~A233;
  assign \new_[27246]_  = ~A232 & \new_[27245]_ ;
  assign \new_[27250]_  = A299 & A298;
  assign \new_[27251]_  = ~A266 & \new_[27250]_ ;
  assign \new_[27252]_  = \new_[27251]_  & \new_[27246]_ ;
  assign \new_[27256]_  = A167 & ~A168;
  assign \new_[27257]_  = A170 & \new_[27256]_ ;
  assign \new_[27261]_  = A200 & ~A199;
  assign \new_[27262]_  = A166 & \new_[27261]_ ;
  assign \new_[27263]_  = \new_[27262]_  & \new_[27257]_ ;
  assign \new_[27267]_  = ~A265 & ~A233;
  assign \new_[27268]_  = ~A232 & \new_[27267]_ ;
  assign \new_[27272]_  = ~A299 & ~A298;
  assign \new_[27273]_  = ~A266 & \new_[27272]_ ;
  assign \new_[27274]_  = \new_[27273]_  & \new_[27268]_ ;
  assign \new_[27278]_  = A167 & ~A168;
  assign \new_[27279]_  = ~A170 & \new_[27278]_ ;
  assign \new_[27283]_  = A200 & ~A199;
  assign \new_[27284]_  = ~A166 & \new_[27283]_ ;
  assign \new_[27285]_  = \new_[27284]_  & \new_[27279]_ ;
  assign \new_[27289]_  = A265 & A233;
  assign \new_[27290]_  = A232 & \new_[27289]_ ;
  assign \new_[27294]_  = ~A300 & ~A299;
  assign \new_[27295]_  = ~A267 & \new_[27294]_ ;
  assign \new_[27296]_  = \new_[27295]_  & \new_[27290]_ ;
  assign \new_[27300]_  = A167 & ~A168;
  assign \new_[27301]_  = ~A170 & \new_[27300]_ ;
  assign \new_[27305]_  = A200 & ~A199;
  assign \new_[27306]_  = ~A166 & \new_[27305]_ ;
  assign \new_[27307]_  = \new_[27306]_  & \new_[27301]_ ;
  assign \new_[27311]_  = A265 & A233;
  assign \new_[27312]_  = A232 & \new_[27311]_ ;
  assign \new_[27316]_  = A299 & A298;
  assign \new_[27317]_  = ~A267 & \new_[27316]_ ;
  assign \new_[27318]_  = \new_[27317]_  & \new_[27312]_ ;
  assign \new_[27322]_  = A167 & ~A168;
  assign \new_[27323]_  = ~A170 & \new_[27322]_ ;
  assign \new_[27327]_  = A200 & ~A199;
  assign \new_[27328]_  = ~A166 & \new_[27327]_ ;
  assign \new_[27329]_  = \new_[27328]_  & \new_[27323]_ ;
  assign \new_[27333]_  = A265 & A233;
  assign \new_[27334]_  = A232 & \new_[27333]_ ;
  assign \new_[27338]_  = ~A299 & ~A298;
  assign \new_[27339]_  = ~A267 & \new_[27338]_ ;
  assign \new_[27340]_  = \new_[27339]_  & \new_[27334]_ ;
  assign \new_[27344]_  = A167 & ~A168;
  assign \new_[27345]_  = ~A170 & \new_[27344]_ ;
  assign \new_[27349]_  = A200 & ~A199;
  assign \new_[27350]_  = ~A166 & \new_[27349]_ ;
  assign \new_[27351]_  = \new_[27350]_  & \new_[27345]_ ;
  assign \new_[27355]_  = A265 & A233;
  assign \new_[27356]_  = A232 & \new_[27355]_ ;
  assign \new_[27360]_  = ~A300 & ~A299;
  assign \new_[27361]_  = A266 & \new_[27360]_ ;
  assign \new_[27362]_  = \new_[27361]_  & \new_[27356]_ ;
  assign \new_[27366]_  = A167 & ~A168;
  assign \new_[27367]_  = ~A170 & \new_[27366]_ ;
  assign \new_[27371]_  = A200 & ~A199;
  assign \new_[27372]_  = ~A166 & \new_[27371]_ ;
  assign \new_[27373]_  = \new_[27372]_  & \new_[27367]_ ;
  assign \new_[27377]_  = A265 & A233;
  assign \new_[27378]_  = A232 & \new_[27377]_ ;
  assign \new_[27382]_  = A299 & A298;
  assign \new_[27383]_  = A266 & \new_[27382]_ ;
  assign \new_[27384]_  = \new_[27383]_  & \new_[27378]_ ;
  assign \new_[27388]_  = A167 & ~A168;
  assign \new_[27389]_  = ~A170 & \new_[27388]_ ;
  assign \new_[27393]_  = A200 & ~A199;
  assign \new_[27394]_  = ~A166 & \new_[27393]_ ;
  assign \new_[27395]_  = \new_[27394]_  & \new_[27389]_ ;
  assign \new_[27399]_  = A265 & A233;
  assign \new_[27400]_  = A232 & \new_[27399]_ ;
  assign \new_[27404]_  = ~A299 & ~A298;
  assign \new_[27405]_  = A266 & \new_[27404]_ ;
  assign \new_[27406]_  = \new_[27405]_  & \new_[27400]_ ;
  assign \new_[27410]_  = A167 & ~A168;
  assign \new_[27411]_  = ~A170 & \new_[27410]_ ;
  assign \new_[27415]_  = A200 & ~A199;
  assign \new_[27416]_  = ~A166 & \new_[27415]_ ;
  assign \new_[27417]_  = \new_[27416]_  & \new_[27411]_ ;
  assign \new_[27421]_  = ~A265 & A233;
  assign \new_[27422]_  = A232 & \new_[27421]_ ;
  assign \new_[27426]_  = ~A300 & ~A299;
  assign \new_[27427]_  = ~A266 & \new_[27426]_ ;
  assign \new_[27428]_  = \new_[27427]_  & \new_[27422]_ ;
  assign \new_[27432]_  = A167 & ~A168;
  assign \new_[27433]_  = ~A170 & \new_[27432]_ ;
  assign \new_[27437]_  = A200 & ~A199;
  assign \new_[27438]_  = ~A166 & \new_[27437]_ ;
  assign \new_[27439]_  = \new_[27438]_  & \new_[27433]_ ;
  assign \new_[27443]_  = ~A265 & A233;
  assign \new_[27444]_  = A232 & \new_[27443]_ ;
  assign \new_[27448]_  = A299 & A298;
  assign \new_[27449]_  = ~A266 & \new_[27448]_ ;
  assign \new_[27450]_  = \new_[27449]_  & \new_[27444]_ ;
  assign \new_[27454]_  = A167 & ~A168;
  assign \new_[27455]_  = ~A170 & \new_[27454]_ ;
  assign \new_[27459]_  = A200 & ~A199;
  assign \new_[27460]_  = ~A166 & \new_[27459]_ ;
  assign \new_[27461]_  = \new_[27460]_  & \new_[27455]_ ;
  assign \new_[27465]_  = ~A265 & A233;
  assign \new_[27466]_  = A232 & \new_[27465]_ ;
  assign \new_[27470]_  = ~A299 & ~A298;
  assign \new_[27471]_  = ~A266 & \new_[27470]_ ;
  assign \new_[27472]_  = \new_[27471]_  & \new_[27466]_ ;
  assign \new_[27476]_  = A167 & ~A168;
  assign \new_[27477]_  = ~A170 & \new_[27476]_ ;
  assign \new_[27481]_  = A200 & ~A199;
  assign \new_[27482]_  = ~A166 & \new_[27481]_ ;
  assign \new_[27483]_  = \new_[27482]_  & \new_[27477]_ ;
  assign \new_[27487]_  = A298 & A233;
  assign \new_[27488]_  = ~A232 & \new_[27487]_ ;
  assign \new_[27492]_  = A301 & A300;
  assign \new_[27493]_  = ~A299 & \new_[27492]_ ;
  assign \new_[27494]_  = \new_[27493]_  & \new_[27488]_ ;
  assign \new_[27498]_  = A167 & ~A168;
  assign \new_[27499]_  = ~A170 & \new_[27498]_ ;
  assign \new_[27503]_  = A200 & ~A199;
  assign \new_[27504]_  = ~A166 & \new_[27503]_ ;
  assign \new_[27505]_  = \new_[27504]_  & \new_[27499]_ ;
  assign \new_[27509]_  = A298 & A233;
  assign \new_[27510]_  = ~A232 & \new_[27509]_ ;
  assign \new_[27514]_  = A302 & A300;
  assign \new_[27515]_  = ~A299 & \new_[27514]_ ;
  assign \new_[27516]_  = \new_[27515]_  & \new_[27510]_ ;
  assign \new_[27520]_  = A167 & ~A168;
  assign \new_[27521]_  = ~A170 & \new_[27520]_ ;
  assign \new_[27525]_  = A200 & ~A199;
  assign \new_[27526]_  = ~A166 & \new_[27525]_ ;
  assign \new_[27527]_  = \new_[27526]_  & \new_[27521]_ ;
  assign \new_[27531]_  = A265 & A233;
  assign \new_[27532]_  = ~A232 & \new_[27531]_ ;
  assign \new_[27536]_  = A268 & A267;
  assign \new_[27537]_  = ~A266 & \new_[27536]_ ;
  assign \new_[27538]_  = \new_[27537]_  & \new_[27532]_ ;
  assign \new_[27542]_  = A167 & ~A168;
  assign \new_[27543]_  = ~A170 & \new_[27542]_ ;
  assign \new_[27547]_  = A200 & ~A199;
  assign \new_[27548]_  = ~A166 & \new_[27547]_ ;
  assign \new_[27549]_  = \new_[27548]_  & \new_[27543]_ ;
  assign \new_[27553]_  = A265 & A233;
  assign \new_[27554]_  = ~A232 & \new_[27553]_ ;
  assign \new_[27558]_  = A269 & A267;
  assign \new_[27559]_  = ~A266 & \new_[27558]_ ;
  assign \new_[27560]_  = \new_[27559]_  & \new_[27554]_ ;
  assign \new_[27564]_  = A167 & ~A168;
  assign \new_[27565]_  = ~A170 & \new_[27564]_ ;
  assign \new_[27569]_  = A200 & ~A199;
  assign \new_[27570]_  = ~A166 & \new_[27569]_ ;
  assign \new_[27571]_  = \new_[27570]_  & \new_[27565]_ ;
  assign \new_[27575]_  = A265 & ~A234;
  assign \new_[27576]_  = ~A233 & \new_[27575]_ ;
  assign \new_[27580]_  = ~A300 & A298;
  assign \new_[27581]_  = A266 & \new_[27580]_ ;
  assign \new_[27582]_  = \new_[27581]_  & \new_[27576]_ ;
  assign \new_[27586]_  = A167 & ~A168;
  assign \new_[27587]_  = ~A170 & \new_[27586]_ ;
  assign \new_[27591]_  = A200 & ~A199;
  assign \new_[27592]_  = ~A166 & \new_[27591]_ ;
  assign \new_[27593]_  = \new_[27592]_  & \new_[27587]_ ;
  assign \new_[27597]_  = A265 & ~A234;
  assign \new_[27598]_  = ~A233 & \new_[27597]_ ;
  assign \new_[27602]_  = A299 & A298;
  assign \new_[27603]_  = A266 & \new_[27602]_ ;
  assign \new_[27604]_  = \new_[27603]_  & \new_[27598]_ ;
  assign \new_[27608]_  = A167 & ~A168;
  assign \new_[27609]_  = ~A170 & \new_[27608]_ ;
  assign \new_[27613]_  = A200 & ~A199;
  assign \new_[27614]_  = ~A166 & \new_[27613]_ ;
  assign \new_[27615]_  = \new_[27614]_  & \new_[27609]_ ;
  assign \new_[27619]_  = A265 & ~A234;
  assign \new_[27620]_  = ~A233 & \new_[27619]_ ;
  assign \new_[27624]_  = ~A299 & ~A298;
  assign \new_[27625]_  = A266 & \new_[27624]_ ;
  assign \new_[27626]_  = \new_[27625]_  & \new_[27620]_ ;
  assign \new_[27630]_  = A167 & ~A168;
  assign \new_[27631]_  = ~A170 & \new_[27630]_ ;
  assign \new_[27635]_  = A200 & ~A199;
  assign \new_[27636]_  = ~A166 & \new_[27635]_ ;
  assign \new_[27637]_  = \new_[27636]_  & \new_[27631]_ ;
  assign \new_[27641]_  = ~A266 & ~A234;
  assign \new_[27642]_  = ~A233 & \new_[27641]_ ;
  assign \new_[27646]_  = ~A300 & A298;
  assign \new_[27647]_  = ~A267 & \new_[27646]_ ;
  assign \new_[27648]_  = \new_[27647]_  & \new_[27642]_ ;
  assign \new_[27652]_  = A167 & ~A168;
  assign \new_[27653]_  = ~A170 & \new_[27652]_ ;
  assign \new_[27657]_  = A200 & ~A199;
  assign \new_[27658]_  = ~A166 & \new_[27657]_ ;
  assign \new_[27659]_  = \new_[27658]_  & \new_[27653]_ ;
  assign \new_[27663]_  = ~A266 & ~A234;
  assign \new_[27664]_  = ~A233 & \new_[27663]_ ;
  assign \new_[27668]_  = A299 & A298;
  assign \new_[27669]_  = ~A267 & \new_[27668]_ ;
  assign \new_[27670]_  = \new_[27669]_  & \new_[27664]_ ;
  assign \new_[27674]_  = A167 & ~A168;
  assign \new_[27675]_  = ~A170 & \new_[27674]_ ;
  assign \new_[27679]_  = A200 & ~A199;
  assign \new_[27680]_  = ~A166 & \new_[27679]_ ;
  assign \new_[27681]_  = \new_[27680]_  & \new_[27675]_ ;
  assign \new_[27685]_  = ~A266 & ~A234;
  assign \new_[27686]_  = ~A233 & \new_[27685]_ ;
  assign \new_[27690]_  = ~A299 & ~A298;
  assign \new_[27691]_  = ~A267 & \new_[27690]_ ;
  assign \new_[27692]_  = \new_[27691]_  & \new_[27686]_ ;
  assign \new_[27696]_  = A167 & ~A168;
  assign \new_[27697]_  = ~A170 & \new_[27696]_ ;
  assign \new_[27701]_  = A200 & ~A199;
  assign \new_[27702]_  = ~A166 & \new_[27701]_ ;
  assign \new_[27703]_  = \new_[27702]_  & \new_[27697]_ ;
  assign \new_[27707]_  = ~A265 & ~A234;
  assign \new_[27708]_  = ~A233 & \new_[27707]_ ;
  assign \new_[27712]_  = ~A300 & A298;
  assign \new_[27713]_  = ~A266 & \new_[27712]_ ;
  assign \new_[27714]_  = \new_[27713]_  & \new_[27708]_ ;
  assign \new_[27718]_  = A167 & ~A168;
  assign \new_[27719]_  = ~A170 & \new_[27718]_ ;
  assign \new_[27723]_  = A200 & ~A199;
  assign \new_[27724]_  = ~A166 & \new_[27723]_ ;
  assign \new_[27725]_  = \new_[27724]_  & \new_[27719]_ ;
  assign \new_[27729]_  = ~A265 & ~A234;
  assign \new_[27730]_  = ~A233 & \new_[27729]_ ;
  assign \new_[27734]_  = A299 & A298;
  assign \new_[27735]_  = ~A266 & \new_[27734]_ ;
  assign \new_[27736]_  = \new_[27735]_  & \new_[27730]_ ;
  assign \new_[27740]_  = A167 & ~A168;
  assign \new_[27741]_  = ~A170 & \new_[27740]_ ;
  assign \new_[27745]_  = A200 & ~A199;
  assign \new_[27746]_  = ~A166 & \new_[27745]_ ;
  assign \new_[27747]_  = \new_[27746]_  & \new_[27741]_ ;
  assign \new_[27751]_  = ~A265 & ~A234;
  assign \new_[27752]_  = ~A233 & \new_[27751]_ ;
  assign \new_[27756]_  = ~A299 & ~A298;
  assign \new_[27757]_  = ~A266 & \new_[27756]_ ;
  assign \new_[27758]_  = \new_[27757]_  & \new_[27752]_ ;
  assign \new_[27762]_  = A167 & ~A168;
  assign \new_[27763]_  = ~A170 & \new_[27762]_ ;
  assign \new_[27767]_  = A200 & ~A199;
  assign \new_[27768]_  = ~A166 & \new_[27767]_ ;
  assign \new_[27769]_  = \new_[27768]_  & \new_[27763]_ ;
  assign \new_[27773]_  = A234 & ~A233;
  assign \new_[27774]_  = A232 & \new_[27773]_ ;
  assign \new_[27778]_  = A299 & ~A298;
  assign \new_[27779]_  = A235 & \new_[27778]_ ;
  assign \new_[27780]_  = \new_[27779]_  & \new_[27774]_ ;
  assign \new_[27784]_  = A167 & ~A168;
  assign \new_[27785]_  = ~A170 & \new_[27784]_ ;
  assign \new_[27789]_  = A200 & ~A199;
  assign \new_[27790]_  = ~A166 & \new_[27789]_ ;
  assign \new_[27791]_  = \new_[27790]_  & \new_[27785]_ ;
  assign \new_[27795]_  = A234 & ~A233;
  assign \new_[27796]_  = A232 & \new_[27795]_ ;
  assign \new_[27800]_  = A266 & ~A265;
  assign \new_[27801]_  = A235 & \new_[27800]_ ;
  assign \new_[27802]_  = \new_[27801]_  & \new_[27796]_ ;
  assign \new_[27806]_  = A167 & ~A168;
  assign \new_[27807]_  = ~A170 & \new_[27806]_ ;
  assign \new_[27811]_  = A200 & ~A199;
  assign \new_[27812]_  = ~A166 & \new_[27811]_ ;
  assign \new_[27813]_  = \new_[27812]_  & \new_[27807]_ ;
  assign \new_[27817]_  = A234 & ~A233;
  assign \new_[27818]_  = A232 & \new_[27817]_ ;
  assign \new_[27822]_  = A299 & ~A298;
  assign \new_[27823]_  = A236 & \new_[27822]_ ;
  assign \new_[27824]_  = \new_[27823]_  & \new_[27818]_ ;
  assign \new_[27828]_  = A167 & ~A168;
  assign \new_[27829]_  = ~A170 & \new_[27828]_ ;
  assign \new_[27833]_  = A200 & ~A199;
  assign \new_[27834]_  = ~A166 & \new_[27833]_ ;
  assign \new_[27835]_  = \new_[27834]_  & \new_[27829]_ ;
  assign \new_[27839]_  = A234 & ~A233;
  assign \new_[27840]_  = A232 & \new_[27839]_ ;
  assign \new_[27844]_  = A266 & ~A265;
  assign \new_[27845]_  = A236 & \new_[27844]_ ;
  assign \new_[27846]_  = \new_[27845]_  & \new_[27840]_ ;
  assign \new_[27850]_  = A167 & ~A168;
  assign \new_[27851]_  = ~A170 & \new_[27850]_ ;
  assign \new_[27855]_  = A200 & ~A199;
  assign \new_[27856]_  = ~A166 & \new_[27855]_ ;
  assign \new_[27857]_  = \new_[27856]_  & \new_[27851]_ ;
  assign \new_[27861]_  = A265 & ~A233;
  assign \new_[27862]_  = ~A232 & \new_[27861]_ ;
  assign \new_[27866]_  = ~A300 & A298;
  assign \new_[27867]_  = A266 & \new_[27866]_ ;
  assign \new_[27868]_  = \new_[27867]_  & \new_[27862]_ ;
  assign \new_[27872]_  = A167 & ~A168;
  assign \new_[27873]_  = ~A170 & \new_[27872]_ ;
  assign \new_[27877]_  = A200 & ~A199;
  assign \new_[27878]_  = ~A166 & \new_[27877]_ ;
  assign \new_[27879]_  = \new_[27878]_  & \new_[27873]_ ;
  assign \new_[27883]_  = A265 & ~A233;
  assign \new_[27884]_  = ~A232 & \new_[27883]_ ;
  assign \new_[27888]_  = A299 & A298;
  assign \new_[27889]_  = A266 & \new_[27888]_ ;
  assign \new_[27890]_  = \new_[27889]_  & \new_[27884]_ ;
  assign \new_[27894]_  = A167 & ~A168;
  assign \new_[27895]_  = ~A170 & \new_[27894]_ ;
  assign \new_[27899]_  = A200 & ~A199;
  assign \new_[27900]_  = ~A166 & \new_[27899]_ ;
  assign \new_[27901]_  = \new_[27900]_  & \new_[27895]_ ;
  assign \new_[27905]_  = A265 & ~A233;
  assign \new_[27906]_  = ~A232 & \new_[27905]_ ;
  assign \new_[27910]_  = ~A299 & ~A298;
  assign \new_[27911]_  = A266 & \new_[27910]_ ;
  assign \new_[27912]_  = \new_[27911]_  & \new_[27906]_ ;
  assign \new_[27916]_  = A167 & ~A168;
  assign \new_[27917]_  = ~A170 & \new_[27916]_ ;
  assign \new_[27921]_  = A200 & ~A199;
  assign \new_[27922]_  = ~A166 & \new_[27921]_ ;
  assign \new_[27923]_  = \new_[27922]_  & \new_[27917]_ ;
  assign \new_[27927]_  = ~A266 & ~A233;
  assign \new_[27928]_  = ~A232 & \new_[27927]_ ;
  assign \new_[27932]_  = ~A300 & A298;
  assign \new_[27933]_  = ~A267 & \new_[27932]_ ;
  assign \new_[27934]_  = \new_[27933]_  & \new_[27928]_ ;
  assign \new_[27938]_  = A167 & ~A168;
  assign \new_[27939]_  = ~A170 & \new_[27938]_ ;
  assign \new_[27943]_  = A200 & ~A199;
  assign \new_[27944]_  = ~A166 & \new_[27943]_ ;
  assign \new_[27945]_  = \new_[27944]_  & \new_[27939]_ ;
  assign \new_[27949]_  = ~A266 & ~A233;
  assign \new_[27950]_  = ~A232 & \new_[27949]_ ;
  assign \new_[27954]_  = A299 & A298;
  assign \new_[27955]_  = ~A267 & \new_[27954]_ ;
  assign \new_[27956]_  = \new_[27955]_  & \new_[27950]_ ;
  assign \new_[27960]_  = A167 & ~A168;
  assign \new_[27961]_  = ~A170 & \new_[27960]_ ;
  assign \new_[27965]_  = A200 & ~A199;
  assign \new_[27966]_  = ~A166 & \new_[27965]_ ;
  assign \new_[27967]_  = \new_[27966]_  & \new_[27961]_ ;
  assign \new_[27971]_  = ~A266 & ~A233;
  assign \new_[27972]_  = ~A232 & \new_[27971]_ ;
  assign \new_[27976]_  = ~A299 & ~A298;
  assign \new_[27977]_  = ~A267 & \new_[27976]_ ;
  assign \new_[27978]_  = \new_[27977]_  & \new_[27972]_ ;
  assign \new_[27982]_  = A167 & ~A168;
  assign \new_[27983]_  = ~A170 & \new_[27982]_ ;
  assign \new_[27987]_  = A200 & ~A199;
  assign \new_[27988]_  = ~A166 & \new_[27987]_ ;
  assign \new_[27989]_  = \new_[27988]_  & \new_[27983]_ ;
  assign \new_[27993]_  = ~A265 & ~A233;
  assign \new_[27994]_  = ~A232 & \new_[27993]_ ;
  assign \new_[27998]_  = ~A300 & A298;
  assign \new_[27999]_  = ~A266 & \new_[27998]_ ;
  assign \new_[28000]_  = \new_[27999]_  & \new_[27994]_ ;
  assign \new_[28004]_  = A167 & ~A168;
  assign \new_[28005]_  = ~A170 & \new_[28004]_ ;
  assign \new_[28009]_  = A200 & ~A199;
  assign \new_[28010]_  = ~A166 & \new_[28009]_ ;
  assign \new_[28011]_  = \new_[28010]_  & \new_[28005]_ ;
  assign \new_[28015]_  = ~A265 & ~A233;
  assign \new_[28016]_  = ~A232 & \new_[28015]_ ;
  assign \new_[28020]_  = A299 & A298;
  assign \new_[28021]_  = ~A266 & \new_[28020]_ ;
  assign \new_[28022]_  = \new_[28021]_  & \new_[28016]_ ;
  assign \new_[28026]_  = A167 & ~A168;
  assign \new_[28027]_  = ~A170 & \new_[28026]_ ;
  assign \new_[28031]_  = A200 & ~A199;
  assign \new_[28032]_  = ~A166 & \new_[28031]_ ;
  assign \new_[28033]_  = \new_[28032]_  & \new_[28027]_ ;
  assign \new_[28037]_  = ~A265 & ~A233;
  assign \new_[28038]_  = ~A232 & \new_[28037]_ ;
  assign \new_[28042]_  = ~A299 & ~A298;
  assign \new_[28043]_  = ~A266 & \new_[28042]_ ;
  assign \new_[28044]_  = \new_[28043]_  & \new_[28038]_ ;
  assign \new_[28048]_  = ~A167 & ~A168;
  assign \new_[28049]_  = ~A170 & \new_[28048]_ ;
  assign \new_[28053]_  = A200 & ~A199;
  assign \new_[28054]_  = A166 & \new_[28053]_ ;
  assign \new_[28055]_  = \new_[28054]_  & \new_[28049]_ ;
  assign \new_[28059]_  = A265 & A233;
  assign \new_[28060]_  = A232 & \new_[28059]_ ;
  assign \new_[28064]_  = ~A300 & ~A299;
  assign \new_[28065]_  = ~A267 & \new_[28064]_ ;
  assign \new_[28066]_  = \new_[28065]_  & \new_[28060]_ ;
  assign \new_[28070]_  = ~A167 & ~A168;
  assign \new_[28071]_  = ~A170 & \new_[28070]_ ;
  assign \new_[28075]_  = A200 & ~A199;
  assign \new_[28076]_  = A166 & \new_[28075]_ ;
  assign \new_[28077]_  = \new_[28076]_  & \new_[28071]_ ;
  assign \new_[28081]_  = A265 & A233;
  assign \new_[28082]_  = A232 & \new_[28081]_ ;
  assign \new_[28086]_  = A299 & A298;
  assign \new_[28087]_  = ~A267 & \new_[28086]_ ;
  assign \new_[28088]_  = \new_[28087]_  & \new_[28082]_ ;
  assign \new_[28092]_  = ~A167 & ~A168;
  assign \new_[28093]_  = ~A170 & \new_[28092]_ ;
  assign \new_[28097]_  = A200 & ~A199;
  assign \new_[28098]_  = A166 & \new_[28097]_ ;
  assign \new_[28099]_  = \new_[28098]_  & \new_[28093]_ ;
  assign \new_[28103]_  = A265 & A233;
  assign \new_[28104]_  = A232 & \new_[28103]_ ;
  assign \new_[28108]_  = ~A299 & ~A298;
  assign \new_[28109]_  = ~A267 & \new_[28108]_ ;
  assign \new_[28110]_  = \new_[28109]_  & \new_[28104]_ ;
  assign \new_[28114]_  = ~A167 & ~A168;
  assign \new_[28115]_  = ~A170 & \new_[28114]_ ;
  assign \new_[28119]_  = A200 & ~A199;
  assign \new_[28120]_  = A166 & \new_[28119]_ ;
  assign \new_[28121]_  = \new_[28120]_  & \new_[28115]_ ;
  assign \new_[28125]_  = A265 & A233;
  assign \new_[28126]_  = A232 & \new_[28125]_ ;
  assign \new_[28130]_  = ~A300 & ~A299;
  assign \new_[28131]_  = A266 & \new_[28130]_ ;
  assign \new_[28132]_  = \new_[28131]_  & \new_[28126]_ ;
  assign \new_[28136]_  = ~A167 & ~A168;
  assign \new_[28137]_  = ~A170 & \new_[28136]_ ;
  assign \new_[28141]_  = A200 & ~A199;
  assign \new_[28142]_  = A166 & \new_[28141]_ ;
  assign \new_[28143]_  = \new_[28142]_  & \new_[28137]_ ;
  assign \new_[28147]_  = A265 & A233;
  assign \new_[28148]_  = A232 & \new_[28147]_ ;
  assign \new_[28152]_  = A299 & A298;
  assign \new_[28153]_  = A266 & \new_[28152]_ ;
  assign \new_[28154]_  = \new_[28153]_  & \new_[28148]_ ;
  assign \new_[28158]_  = ~A167 & ~A168;
  assign \new_[28159]_  = ~A170 & \new_[28158]_ ;
  assign \new_[28163]_  = A200 & ~A199;
  assign \new_[28164]_  = A166 & \new_[28163]_ ;
  assign \new_[28165]_  = \new_[28164]_  & \new_[28159]_ ;
  assign \new_[28169]_  = A265 & A233;
  assign \new_[28170]_  = A232 & \new_[28169]_ ;
  assign \new_[28174]_  = ~A299 & ~A298;
  assign \new_[28175]_  = A266 & \new_[28174]_ ;
  assign \new_[28176]_  = \new_[28175]_  & \new_[28170]_ ;
  assign \new_[28180]_  = ~A167 & ~A168;
  assign \new_[28181]_  = ~A170 & \new_[28180]_ ;
  assign \new_[28185]_  = A200 & ~A199;
  assign \new_[28186]_  = A166 & \new_[28185]_ ;
  assign \new_[28187]_  = \new_[28186]_  & \new_[28181]_ ;
  assign \new_[28191]_  = ~A265 & A233;
  assign \new_[28192]_  = A232 & \new_[28191]_ ;
  assign \new_[28196]_  = ~A300 & ~A299;
  assign \new_[28197]_  = ~A266 & \new_[28196]_ ;
  assign \new_[28198]_  = \new_[28197]_  & \new_[28192]_ ;
  assign \new_[28202]_  = ~A167 & ~A168;
  assign \new_[28203]_  = ~A170 & \new_[28202]_ ;
  assign \new_[28207]_  = A200 & ~A199;
  assign \new_[28208]_  = A166 & \new_[28207]_ ;
  assign \new_[28209]_  = \new_[28208]_  & \new_[28203]_ ;
  assign \new_[28213]_  = ~A265 & A233;
  assign \new_[28214]_  = A232 & \new_[28213]_ ;
  assign \new_[28218]_  = A299 & A298;
  assign \new_[28219]_  = ~A266 & \new_[28218]_ ;
  assign \new_[28220]_  = \new_[28219]_  & \new_[28214]_ ;
  assign \new_[28224]_  = ~A167 & ~A168;
  assign \new_[28225]_  = ~A170 & \new_[28224]_ ;
  assign \new_[28229]_  = A200 & ~A199;
  assign \new_[28230]_  = A166 & \new_[28229]_ ;
  assign \new_[28231]_  = \new_[28230]_  & \new_[28225]_ ;
  assign \new_[28235]_  = ~A265 & A233;
  assign \new_[28236]_  = A232 & \new_[28235]_ ;
  assign \new_[28240]_  = ~A299 & ~A298;
  assign \new_[28241]_  = ~A266 & \new_[28240]_ ;
  assign \new_[28242]_  = \new_[28241]_  & \new_[28236]_ ;
  assign \new_[28246]_  = ~A167 & ~A168;
  assign \new_[28247]_  = ~A170 & \new_[28246]_ ;
  assign \new_[28251]_  = A200 & ~A199;
  assign \new_[28252]_  = A166 & \new_[28251]_ ;
  assign \new_[28253]_  = \new_[28252]_  & \new_[28247]_ ;
  assign \new_[28257]_  = A298 & A233;
  assign \new_[28258]_  = ~A232 & \new_[28257]_ ;
  assign \new_[28262]_  = A301 & A300;
  assign \new_[28263]_  = ~A299 & \new_[28262]_ ;
  assign \new_[28264]_  = \new_[28263]_  & \new_[28258]_ ;
  assign \new_[28268]_  = ~A167 & ~A168;
  assign \new_[28269]_  = ~A170 & \new_[28268]_ ;
  assign \new_[28273]_  = A200 & ~A199;
  assign \new_[28274]_  = A166 & \new_[28273]_ ;
  assign \new_[28275]_  = \new_[28274]_  & \new_[28269]_ ;
  assign \new_[28279]_  = A298 & A233;
  assign \new_[28280]_  = ~A232 & \new_[28279]_ ;
  assign \new_[28284]_  = A302 & A300;
  assign \new_[28285]_  = ~A299 & \new_[28284]_ ;
  assign \new_[28286]_  = \new_[28285]_  & \new_[28280]_ ;
  assign \new_[28290]_  = ~A167 & ~A168;
  assign \new_[28291]_  = ~A170 & \new_[28290]_ ;
  assign \new_[28295]_  = A200 & ~A199;
  assign \new_[28296]_  = A166 & \new_[28295]_ ;
  assign \new_[28297]_  = \new_[28296]_  & \new_[28291]_ ;
  assign \new_[28301]_  = A265 & A233;
  assign \new_[28302]_  = ~A232 & \new_[28301]_ ;
  assign \new_[28306]_  = A268 & A267;
  assign \new_[28307]_  = ~A266 & \new_[28306]_ ;
  assign \new_[28308]_  = \new_[28307]_  & \new_[28302]_ ;
  assign \new_[28312]_  = ~A167 & ~A168;
  assign \new_[28313]_  = ~A170 & \new_[28312]_ ;
  assign \new_[28317]_  = A200 & ~A199;
  assign \new_[28318]_  = A166 & \new_[28317]_ ;
  assign \new_[28319]_  = \new_[28318]_  & \new_[28313]_ ;
  assign \new_[28323]_  = A265 & A233;
  assign \new_[28324]_  = ~A232 & \new_[28323]_ ;
  assign \new_[28328]_  = A269 & A267;
  assign \new_[28329]_  = ~A266 & \new_[28328]_ ;
  assign \new_[28330]_  = \new_[28329]_  & \new_[28324]_ ;
  assign \new_[28334]_  = ~A167 & ~A168;
  assign \new_[28335]_  = ~A170 & \new_[28334]_ ;
  assign \new_[28339]_  = A200 & ~A199;
  assign \new_[28340]_  = A166 & \new_[28339]_ ;
  assign \new_[28341]_  = \new_[28340]_  & \new_[28335]_ ;
  assign \new_[28345]_  = A265 & ~A234;
  assign \new_[28346]_  = ~A233 & \new_[28345]_ ;
  assign \new_[28350]_  = ~A300 & A298;
  assign \new_[28351]_  = A266 & \new_[28350]_ ;
  assign \new_[28352]_  = \new_[28351]_  & \new_[28346]_ ;
  assign \new_[28356]_  = ~A167 & ~A168;
  assign \new_[28357]_  = ~A170 & \new_[28356]_ ;
  assign \new_[28361]_  = A200 & ~A199;
  assign \new_[28362]_  = A166 & \new_[28361]_ ;
  assign \new_[28363]_  = \new_[28362]_  & \new_[28357]_ ;
  assign \new_[28367]_  = A265 & ~A234;
  assign \new_[28368]_  = ~A233 & \new_[28367]_ ;
  assign \new_[28372]_  = A299 & A298;
  assign \new_[28373]_  = A266 & \new_[28372]_ ;
  assign \new_[28374]_  = \new_[28373]_  & \new_[28368]_ ;
  assign \new_[28378]_  = ~A167 & ~A168;
  assign \new_[28379]_  = ~A170 & \new_[28378]_ ;
  assign \new_[28383]_  = A200 & ~A199;
  assign \new_[28384]_  = A166 & \new_[28383]_ ;
  assign \new_[28385]_  = \new_[28384]_  & \new_[28379]_ ;
  assign \new_[28389]_  = A265 & ~A234;
  assign \new_[28390]_  = ~A233 & \new_[28389]_ ;
  assign \new_[28394]_  = ~A299 & ~A298;
  assign \new_[28395]_  = A266 & \new_[28394]_ ;
  assign \new_[28396]_  = \new_[28395]_  & \new_[28390]_ ;
  assign \new_[28400]_  = ~A167 & ~A168;
  assign \new_[28401]_  = ~A170 & \new_[28400]_ ;
  assign \new_[28405]_  = A200 & ~A199;
  assign \new_[28406]_  = A166 & \new_[28405]_ ;
  assign \new_[28407]_  = \new_[28406]_  & \new_[28401]_ ;
  assign \new_[28411]_  = ~A266 & ~A234;
  assign \new_[28412]_  = ~A233 & \new_[28411]_ ;
  assign \new_[28416]_  = ~A300 & A298;
  assign \new_[28417]_  = ~A267 & \new_[28416]_ ;
  assign \new_[28418]_  = \new_[28417]_  & \new_[28412]_ ;
  assign \new_[28422]_  = ~A167 & ~A168;
  assign \new_[28423]_  = ~A170 & \new_[28422]_ ;
  assign \new_[28427]_  = A200 & ~A199;
  assign \new_[28428]_  = A166 & \new_[28427]_ ;
  assign \new_[28429]_  = \new_[28428]_  & \new_[28423]_ ;
  assign \new_[28433]_  = ~A266 & ~A234;
  assign \new_[28434]_  = ~A233 & \new_[28433]_ ;
  assign \new_[28438]_  = A299 & A298;
  assign \new_[28439]_  = ~A267 & \new_[28438]_ ;
  assign \new_[28440]_  = \new_[28439]_  & \new_[28434]_ ;
  assign \new_[28444]_  = ~A167 & ~A168;
  assign \new_[28445]_  = ~A170 & \new_[28444]_ ;
  assign \new_[28449]_  = A200 & ~A199;
  assign \new_[28450]_  = A166 & \new_[28449]_ ;
  assign \new_[28451]_  = \new_[28450]_  & \new_[28445]_ ;
  assign \new_[28455]_  = ~A266 & ~A234;
  assign \new_[28456]_  = ~A233 & \new_[28455]_ ;
  assign \new_[28460]_  = ~A299 & ~A298;
  assign \new_[28461]_  = ~A267 & \new_[28460]_ ;
  assign \new_[28462]_  = \new_[28461]_  & \new_[28456]_ ;
  assign \new_[28466]_  = ~A167 & ~A168;
  assign \new_[28467]_  = ~A170 & \new_[28466]_ ;
  assign \new_[28471]_  = A200 & ~A199;
  assign \new_[28472]_  = A166 & \new_[28471]_ ;
  assign \new_[28473]_  = \new_[28472]_  & \new_[28467]_ ;
  assign \new_[28477]_  = ~A265 & ~A234;
  assign \new_[28478]_  = ~A233 & \new_[28477]_ ;
  assign \new_[28482]_  = ~A300 & A298;
  assign \new_[28483]_  = ~A266 & \new_[28482]_ ;
  assign \new_[28484]_  = \new_[28483]_  & \new_[28478]_ ;
  assign \new_[28488]_  = ~A167 & ~A168;
  assign \new_[28489]_  = ~A170 & \new_[28488]_ ;
  assign \new_[28493]_  = A200 & ~A199;
  assign \new_[28494]_  = A166 & \new_[28493]_ ;
  assign \new_[28495]_  = \new_[28494]_  & \new_[28489]_ ;
  assign \new_[28499]_  = ~A265 & ~A234;
  assign \new_[28500]_  = ~A233 & \new_[28499]_ ;
  assign \new_[28504]_  = A299 & A298;
  assign \new_[28505]_  = ~A266 & \new_[28504]_ ;
  assign \new_[28506]_  = \new_[28505]_  & \new_[28500]_ ;
  assign \new_[28510]_  = ~A167 & ~A168;
  assign \new_[28511]_  = ~A170 & \new_[28510]_ ;
  assign \new_[28515]_  = A200 & ~A199;
  assign \new_[28516]_  = A166 & \new_[28515]_ ;
  assign \new_[28517]_  = \new_[28516]_  & \new_[28511]_ ;
  assign \new_[28521]_  = ~A265 & ~A234;
  assign \new_[28522]_  = ~A233 & \new_[28521]_ ;
  assign \new_[28526]_  = ~A299 & ~A298;
  assign \new_[28527]_  = ~A266 & \new_[28526]_ ;
  assign \new_[28528]_  = \new_[28527]_  & \new_[28522]_ ;
  assign \new_[28532]_  = ~A167 & ~A168;
  assign \new_[28533]_  = ~A170 & \new_[28532]_ ;
  assign \new_[28537]_  = A200 & ~A199;
  assign \new_[28538]_  = A166 & \new_[28537]_ ;
  assign \new_[28539]_  = \new_[28538]_  & \new_[28533]_ ;
  assign \new_[28543]_  = A234 & ~A233;
  assign \new_[28544]_  = A232 & \new_[28543]_ ;
  assign \new_[28548]_  = A299 & ~A298;
  assign \new_[28549]_  = A235 & \new_[28548]_ ;
  assign \new_[28550]_  = \new_[28549]_  & \new_[28544]_ ;
  assign \new_[28554]_  = ~A167 & ~A168;
  assign \new_[28555]_  = ~A170 & \new_[28554]_ ;
  assign \new_[28559]_  = A200 & ~A199;
  assign \new_[28560]_  = A166 & \new_[28559]_ ;
  assign \new_[28561]_  = \new_[28560]_  & \new_[28555]_ ;
  assign \new_[28565]_  = A234 & ~A233;
  assign \new_[28566]_  = A232 & \new_[28565]_ ;
  assign \new_[28570]_  = A266 & ~A265;
  assign \new_[28571]_  = A235 & \new_[28570]_ ;
  assign \new_[28572]_  = \new_[28571]_  & \new_[28566]_ ;
  assign \new_[28576]_  = ~A167 & ~A168;
  assign \new_[28577]_  = ~A170 & \new_[28576]_ ;
  assign \new_[28581]_  = A200 & ~A199;
  assign \new_[28582]_  = A166 & \new_[28581]_ ;
  assign \new_[28583]_  = \new_[28582]_  & \new_[28577]_ ;
  assign \new_[28587]_  = A234 & ~A233;
  assign \new_[28588]_  = A232 & \new_[28587]_ ;
  assign \new_[28592]_  = A299 & ~A298;
  assign \new_[28593]_  = A236 & \new_[28592]_ ;
  assign \new_[28594]_  = \new_[28593]_  & \new_[28588]_ ;
  assign \new_[28598]_  = ~A167 & ~A168;
  assign \new_[28599]_  = ~A170 & \new_[28598]_ ;
  assign \new_[28603]_  = A200 & ~A199;
  assign \new_[28604]_  = A166 & \new_[28603]_ ;
  assign \new_[28605]_  = \new_[28604]_  & \new_[28599]_ ;
  assign \new_[28609]_  = A234 & ~A233;
  assign \new_[28610]_  = A232 & \new_[28609]_ ;
  assign \new_[28614]_  = A266 & ~A265;
  assign \new_[28615]_  = A236 & \new_[28614]_ ;
  assign \new_[28616]_  = \new_[28615]_  & \new_[28610]_ ;
  assign \new_[28620]_  = ~A167 & ~A168;
  assign \new_[28621]_  = ~A170 & \new_[28620]_ ;
  assign \new_[28625]_  = A200 & ~A199;
  assign \new_[28626]_  = A166 & \new_[28625]_ ;
  assign \new_[28627]_  = \new_[28626]_  & \new_[28621]_ ;
  assign \new_[28631]_  = A265 & ~A233;
  assign \new_[28632]_  = ~A232 & \new_[28631]_ ;
  assign \new_[28636]_  = ~A300 & A298;
  assign \new_[28637]_  = A266 & \new_[28636]_ ;
  assign \new_[28638]_  = \new_[28637]_  & \new_[28632]_ ;
  assign \new_[28642]_  = ~A167 & ~A168;
  assign \new_[28643]_  = ~A170 & \new_[28642]_ ;
  assign \new_[28647]_  = A200 & ~A199;
  assign \new_[28648]_  = A166 & \new_[28647]_ ;
  assign \new_[28649]_  = \new_[28648]_  & \new_[28643]_ ;
  assign \new_[28653]_  = A265 & ~A233;
  assign \new_[28654]_  = ~A232 & \new_[28653]_ ;
  assign \new_[28658]_  = A299 & A298;
  assign \new_[28659]_  = A266 & \new_[28658]_ ;
  assign \new_[28660]_  = \new_[28659]_  & \new_[28654]_ ;
  assign \new_[28664]_  = ~A167 & ~A168;
  assign \new_[28665]_  = ~A170 & \new_[28664]_ ;
  assign \new_[28669]_  = A200 & ~A199;
  assign \new_[28670]_  = A166 & \new_[28669]_ ;
  assign \new_[28671]_  = \new_[28670]_  & \new_[28665]_ ;
  assign \new_[28675]_  = A265 & ~A233;
  assign \new_[28676]_  = ~A232 & \new_[28675]_ ;
  assign \new_[28680]_  = ~A299 & ~A298;
  assign \new_[28681]_  = A266 & \new_[28680]_ ;
  assign \new_[28682]_  = \new_[28681]_  & \new_[28676]_ ;
  assign \new_[28686]_  = ~A167 & ~A168;
  assign \new_[28687]_  = ~A170 & \new_[28686]_ ;
  assign \new_[28691]_  = A200 & ~A199;
  assign \new_[28692]_  = A166 & \new_[28691]_ ;
  assign \new_[28693]_  = \new_[28692]_  & \new_[28687]_ ;
  assign \new_[28697]_  = ~A266 & ~A233;
  assign \new_[28698]_  = ~A232 & \new_[28697]_ ;
  assign \new_[28702]_  = ~A300 & A298;
  assign \new_[28703]_  = ~A267 & \new_[28702]_ ;
  assign \new_[28704]_  = \new_[28703]_  & \new_[28698]_ ;
  assign \new_[28708]_  = ~A167 & ~A168;
  assign \new_[28709]_  = ~A170 & \new_[28708]_ ;
  assign \new_[28713]_  = A200 & ~A199;
  assign \new_[28714]_  = A166 & \new_[28713]_ ;
  assign \new_[28715]_  = \new_[28714]_  & \new_[28709]_ ;
  assign \new_[28719]_  = ~A266 & ~A233;
  assign \new_[28720]_  = ~A232 & \new_[28719]_ ;
  assign \new_[28724]_  = A299 & A298;
  assign \new_[28725]_  = ~A267 & \new_[28724]_ ;
  assign \new_[28726]_  = \new_[28725]_  & \new_[28720]_ ;
  assign \new_[28730]_  = ~A167 & ~A168;
  assign \new_[28731]_  = ~A170 & \new_[28730]_ ;
  assign \new_[28735]_  = A200 & ~A199;
  assign \new_[28736]_  = A166 & \new_[28735]_ ;
  assign \new_[28737]_  = \new_[28736]_  & \new_[28731]_ ;
  assign \new_[28741]_  = ~A266 & ~A233;
  assign \new_[28742]_  = ~A232 & \new_[28741]_ ;
  assign \new_[28746]_  = ~A299 & ~A298;
  assign \new_[28747]_  = ~A267 & \new_[28746]_ ;
  assign \new_[28748]_  = \new_[28747]_  & \new_[28742]_ ;
  assign \new_[28752]_  = ~A167 & ~A168;
  assign \new_[28753]_  = ~A170 & \new_[28752]_ ;
  assign \new_[28757]_  = A200 & ~A199;
  assign \new_[28758]_  = A166 & \new_[28757]_ ;
  assign \new_[28759]_  = \new_[28758]_  & \new_[28753]_ ;
  assign \new_[28763]_  = ~A265 & ~A233;
  assign \new_[28764]_  = ~A232 & \new_[28763]_ ;
  assign \new_[28768]_  = ~A300 & A298;
  assign \new_[28769]_  = ~A266 & \new_[28768]_ ;
  assign \new_[28770]_  = \new_[28769]_  & \new_[28764]_ ;
  assign \new_[28774]_  = ~A167 & ~A168;
  assign \new_[28775]_  = ~A170 & \new_[28774]_ ;
  assign \new_[28779]_  = A200 & ~A199;
  assign \new_[28780]_  = A166 & \new_[28779]_ ;
  assign \new_[28781]_  = \new_[28780]_  & \new_[28775]_ ;
  assign \new_[28785]_  = ~A265 & ~A233;
  assign \new_[28786]_  = ~A232 & \new_[28785]_ ;
  assign \new_[28790]_  = A299 & A298;
  assign \new_[28791]_  = ~A266 & \new_[28790]_ ;
  assign \new_[28792]_  = \new_[28791]_  & \new_[28786]_ ;
  assign \new_[28796]_  = ~A167 & ~A168;
  assign \new_[28797]_  = ~A170 & \new_[28796]_ ;
  assign \new_[28801]_  = A200 & ~A199;
  assign \new_[28802]_  = A166 & \new_[28801]_ ;
  assign \new_[28803]_  = \new_[28802]_  & \new_[28797]_ ;
  assign \new_[28807]_  = ~A265 & ~A233;
  assign \new_[28808]_  = ~A232 & \new_[28807]_ ;
  assign \new_[28812]_  = ~A299 & ~A298;
  assign \new_[28813]_  = ~A266 & \new_[28812]_ ;
  assign \new_[28814]_  = \new_[28813]_  & \new_[28808]_ ;
  assign \new_[28818]_  = A167 & ~A168;
  assign \new_[28819]_  = A169 & \new_[28818]_ ;
  assign \new_[28823]_  = A200 & ~A199;
  assign \new_[28824]_  = ~A166 & \new_[28823]_ ;
  assign \new_[28825]_  = \new_[28824]_  & \new_[28819]_ ;
  assign \new_[28829]_  = A265 & A233;
  assign \new_[28830]_  = A232 & \new_[28829]_ ;
  assign \new_[28834]_  = ~A300 & ~A299;
  assign \new_[28835]_  = ~A267 & \new_[28834]_ ;
  assign \new_[28836]_  = \new_[28835]_  & \new_[28830]_ ;
  assign \new_[28840]_  = A167 & ~A168;
  assign \new_[28841]_  = A169 & \new_[28840]_ ;
  assign \new_[28845]_  = A200 & ~A199;
  assign \new_[28846]_  = ~A166 & \new_[28845]_ ;
  assign \new_[28847]_  = \new_[28846]_  & \new_[28841]_ ;
  assign \new_[28851]_  = A265 & A233;
  assign \new_[28852]_  = A232 & \new_[28851]_ ;
  assign \new_[28856]_  = A299 & A298;
  assign \new_[28857]_  = ~A267 & \new_[28856]_ ;
  assign \new_[28858]_  = \new_[28857]_  & \new_[28852]_ ;
  assign \new_[28862]_  = A167 & ~A168;
  assign \new_[28863]_  = A169 & \new_[28862]_ ;
  assign \new_[28867]_  = A200 & ~A199;
  assign \new_[28868]_  = ~A166 & \new_[28867]_ ;
  assign \new_[28869]_  = \new_[28868]_  & \new_[28863]_ ;
  assign \new_[28873]_  = A265 & A233;
  assign \new_[28874]_  = A232 & \new_[28873]_ ;
  assign \new_[28878]_  = ~A299 & ~A298;
  assign \new_[28879]_  = ~A267 & \new_[28878]_ ;
  assign \new_[28880]_  = \new_[28879]_  & \new_[28874]_ ;
  assign \new_[28884]_  = A167 & ~A168;
  assign \new_[28885]_  = A169 & \new_[28884]_ ;
  assign \new_[28889]_  = A200 & ~A199;
  assign \new_[28890]_  = ~A166 & \new_[28889]_ ;
  assign \new_[28891]_  = \new_[28890]_  & \new_[28885]_ ;
  assign \new_[28895]_  = A265 & A233;
  assign \new_[28896]_  = A232 & \new_[28895]_ ;
  assign \new_[28900]_  = ~A300 & ~A299;
  assign \new_[28901]_  = A266 & \new_[28900]_ ;
  assign \new_[28902]_  = \new_[28901]_  & \new_[28896]_ ;
  assign \new_[28906]_  = A167 & ~A168;
  assign \new_[28907]_  = A169 & \new_[28906]_ ;
  assign \new_[28911]_  = A200 & ~A199;
  assign \new_[28912]_  = ~A166 & \new_[28911]_ ;
  assign \new_[28913]_  = \new_[28912]_  & \new_[28907]_ ;
  assign \new_[28917]_  = A265 & A233;
  assign \new_[28918]_  = A232 & \new_[28917]_ ;
  assign \new_[28922]_  = A299 & A298;
  assign \new_[28923]_  = A266 & \new_[28922]_ ;
  assign \new_[28924]_  = \new_[28923]_  & \new_[28918]_ ;
  assign \new_[28928]_  = A167 & ~A168;
  assign \new_[28929]_  = A169 & \new_[28928]_ ;
  assign \new_[28933]_  = A200 & ~A199;
  assign \new_[28934]_  = ~A166 & \new_[28933]_ ;
  assign \new_[28935]_  = \new_[28934]_  & \new_[28929]_ ;
  assign \new_[28939]_  = A265 & A233;
  assign \new_[28940]_  = A232 & \new_[28939]_ ;
  assign \new_[28944]_  = ~A299 & ~A298;
  assign \new_[28945]_  = A266 & \new_[28944]_ ;
  assign \new_[28946]_  = \new_[28945]_  & \new_[28940]_ ;
  assign \new_[28950]_  = A167 & ~A168;
  assign \new_[28951]_  = A169 & \new_[28950]_ ;
  assign \new_[28955]_  = A200 & ~A199;
  assign \new_[28956]_  = ~A166 & \new_[28955]_ ;
  assign \new_[28957]_  = \new_[28956]_  & \new_[28951]_ ;
  assign \new_[28961]_  = ~A265 & A233;
  assign \new_[28962]_  = A232 & \new_[28961]_ ;
  assign \new_[28966]_  = ~A300 & ~A299;
  assign \new_[28967]_  = ~A266 & \new_[28966]_ ;
  assign \new_[28968]_  = \new_[28967]_  & \new_[28962]_ ;
  assign \new_[28972]_  = A167 & ~A168;
  assign \new_[28973]_  = A169 & \new_[28972]_ ;
  assign \new_[28977]_  = A200 & ~A199;
  assign \new_[28978]_  = ~A166 & \new_[28977]_ ;
  assign \new_[28979]_  = \new_[28978]_  & \new_[28973]_ ;
  assign \new_[28983]_  = ~A265 & A233;
  assign \new_[28984]_  = A232 & \new_[28983]_ ;
  assign \new_[28988]_  = A299 & A298;
  assign \new_[28989]_  = ~A266 & \new_[28988]_ ;
  assign \new_[28990]_  = \new_[28989]_  & \new_[28984]_ ;
  assign \new_[28994]_  = A167 & ~A168;
  assign \new_[28995]_  = A169 & \new_[28994]_ ;
  assign \new_[28999]_  = A200 & ~A199;
  assign \new_[29000]_  = ~A166 & \new_[28999]_ ;
  assign \new_[29001]_  = \new_[29000]_  & \new_[28995]_ ;
  assign \new_[29005]_  = ~A265 & A233;
  assign \new_[29006]_  = A232 & \new_[29005]_ ;
  assign \new_[29010]_  = ~A299 & ~A298;
  assign \new_[29011]_  = ~A266 & \new_[29010]_ ;
  assign \new_[29012]_  = \new_[29011]_  & \new_[29006]_ ;
  assign \new_[29016]_  = A167 & ~A168;
  assign \new_[29017]_  = A169 & \new_[29016]_ ;
  assign \new_[29021]_  = A200 & ~A199;
  assign \new_[29022]_  = ~A166 & \new_[29021]_ ;
  assign \new_[29023]_  = \new_[29022]_  & \new_[29017]_ ;
  assign \new_[29027]_  = A298 & A233;
  assign \new_[29028]_  = ~A232 & \new_[29027]_ ;
  assign \new_[29032]_  = A301 & A300;
  assign \new_[29033]_  = ~A299 & \new_[29032]_ ;
  assign \new_[29034]_  = \new_[29033]_  & \new_[29028]_ ;
  assign \new_[29038]_  = A167 & ~A168;
  assign \new_[29039]_  = A169 & \new_[29038]_ ;
  assign \new_[29043]_  = A200 & ~A199;
  assign \new_[29044]_  = ~A166 & \new_[29043]_ ;
  assign \new_[29045]_  = \new_[29044]_  & \new_[29039]_ ;
  assign \new_[29049]_  = A298 & A233;
  assign \new_[29050]_  = ~A232 & \new_[29049]_ ;
  assign \new_[29054]_  = A302 & A300;
  assign \new_[29055]_  = ~A299 & \new_[29054]_ ;
  assign \new_[29056]_  = \new_[29055]_  & \new_[29050]_ ;
  assign \new_[29060]_  = A167 & ~A168;
  assign \new_[29061]_  = A169 & \new_[29060]_ ;
  assign \new_[29065]_  = A200 & ~A199;
  assign \new_[29066]_  = ~A166 & \new_[29065]_ ;
  assign \new_[29067]_  = \new_[29066]_  & \new_[29061]_ ;
  assign \new_[29071]_  = A265 & A233;
  assign \new_[29072]_  = ~A232 & \new_[29071]_ ;
  assign \new_[29076]_  = A268 & A267;
  assign \new_[29077]_  = ~A266 & \new_[29076]_ ;
  assign \new_[29078]_  = \new_[29077]_  & \new_[29072]_ ;
  assign \new_[29082]_  = A167 & ~A168;
  assign \new_[29083]_  = A169 & \new_[29082]_ ;
  assign \new_[29087]_  = A200 & ~A199;
  assign \new_[29088]_  = ~A166 & \new_[29087]_ ;
  assign \new_[29089]_  = \new_[29088]_  & \new_[29083]_ ;
  assign \new_[29093]_  = A265 & A233;
  assign \new_[29094]_  = ~A232 & \new_[29093]_ ;
  assign \new_[29098]_  = A269 & A267;
  assign \new_[29099]_  = ~A266 & \new_[29098]_ ;
  assign \new_[29100]_  = \new_[29099]_  & \new_[29094]_ ;
  assign \new_[29104]_  = A167 & ~A168;
  assign \new_[29105]_  = A169 & \new_[29104]_ ;
  assign \new_[29109]_  = A200 & ~A199;
  assign \new_[29110]_  = ~A166 & \new_[29109]_ ;
  assign \new_[29111]_  = \new_[29110]_  & \new_[29105]_ ;
  assign \new_[29115]_  = A265 & ~A234;
  assign \new_[29116]_  = ~A233 & \new_[29115]_ ;
  assign \new_[29120]_  = ~A300 & A298;
  assign \new_[29121]_  = A266 & \new_[29120]_ ;
  assign \new_[29122]_  = \new_[29121]_  & \new_[29116]_ ;
  assign \new_[29126]_  = A167 & ~A168;
  assign \new_[29127]_  = A169 & \new_[29126]_ ;
  assign \new_[29131]_  = A200 & ~A199;
  assign \new_[29132]_  = ~A166 & \new_[29131]_ ;
  assign \new_[29133]_  = \new_[29132]_  & \new_[29127]_ ;
  assign \new_[29137]_  = A265 & ~A234;
  assign \new_[29138]_  = ~A233 & \new_[29137]_ ;
  assign \new_[29142]_  = A299 & A298;
  assign \new_[29143]_  = A266 & \new_[29142]_ ;
  assign \new_[29144]_  = \new_[29143]_  & \new_[29138]_ ;
  assign \new_[29148]_  = A167 & ~A168;
  assign \new_[29149]_  = A169 & \new_[29148]_ ;
  assign \new_[29153]_  = A200 & ~A199;
  assign \new_[29154]_  = ~A166 & \new_[29153]_ ;
  assign \new_[29155]_  = \new_[29154]_  & \new_[29149]_ ;
  assign \new_[29159]_  = A265 & ~A234;
  assign \new_[29160]_  = ~A233 & \new_[29159]_ ;
  assign \new_[29164]_  = ~A299 & ~A298;
  assign \new_[29165]_  = A266 & \new_[29164]_ ;
  assign \new_[29166]_  = \new_[29165]_  & \new_[29160]_ ;
  assign \new_[29170]_  = A167 & ~A168;
  assign \new_[29171]_  = A169 & \new_[29170]_ ;
  assign \new_[29175]_  = A200 & ~A199;
  assign \new_[29176]_  = ~A166 & \new_[29175]_ ;
  assign \new_[29177]_  = \new_[29176]_  & \new_[29171]_ ;
  assign \new_[29181]_  = ~A266 & ~A234;
  assign \new_[29182]_  = ~A233 & \new_[29181]_ ;
  assign \new_[29186]_  = ~A300 & A298;
  assign \new_[29187]_  = ~A267 & \new_[29186]_ ;
  assign \new_[29188]_  = \new_[29187]_  & \new_[29182]_ ;
  assign \new_[29192]_  = A167 & ~A168;
  assign \new_[29193]_  = A169 & \new_[29192]_ ;
  assign \new_[29197]_  = A200 & ~A199;
  assign \new_[29198]_  = ~A166 & \new_[29197]_ ;
  assign \new_[29199]_  = \new_[29198]_  & \new_[29193]_ ;
  assign \new_[29203]_  = ~A266 & ~A234;
  assign \new_[29204]_  = ~A233 & \new_[29203]_ ;
  assign \new_[29208]_  = A299 & A298;
  assign \new_[29209]_  = ~A267 & \new_[29208]_ ;
  assign \new_[29210]_  = \new_[29209]_  & \new_[29204]_ ;
  assign \new_[29214]_  = A167 & ~A168;
  assign \new_[29215]_  = A169 & \new_[29214]_ ;
  assign \new_[29219]_  = A200 & ~A199;
  assign \new_[29220]_  = ~A166 & \new_[29219]_ ;
  assign \new_[29221]_  = \new_[29220]_  & \new_[29215]_ ;
  assign \new_[29225]_  = ~A266 & ~A234;
  assign \new_[29226]_  = ~A233 & \new_[29225]_ ;
  assign \new_[29230]_  = ~A299 & ~A298;
  assign \new_[29231]_  = ~A267 & \new_[29230]_ ;
  assign \new_[29232]_  = \new_[29231]_  & \new_[29226]_ ;
  assign \new_[29236]_  = A167 & ~A168;
  assign \new_[29237]_  = A169 & \new_[29236]_ ;
  assign \new_[29241]_  = A200 & ~A199;
  assign \new_[29242]_  = ~A166 & \new_[29241]_ ;
  assign \new_[29243]_  = \new_[29242]_  & \new_[29237]_ ;
  assign \new_[29247]_  = ~A265 & ~A234;
  assign \new_[29248]_  = ~A233 & \new_[29247]_ ;
  assign \new_[29252]_  = ~A300 & A298;
  assign \new_[29253]_  = ~A266 & \new_[29252]_ ;
  assign \new_[29254]_  = \new_[29253]_  & \new_[29248]_ ;
  assign \new_[29258]_  = A167 & ~A168;
  assign \new_[29259]_  = A169 & \new_[29258]_ ;
  assign \new_[29263]_  = A200 & ~A199;
  assign \new_[29264]_  = ~A166 & \new_[29263]_ ;
  assign \new_[29265]_  = \new_[29264]_  & \new_[29259]_ ;
  assign \new_[29269]_  = ~A265 & ~A234;
  assign \new_[29270]_  = ~A233 & \new_[29269]_ ;
  assign \new_[29274]_  = A299 & A298;
  assign \new_[29275]_  = ~A266 & \new_[29274]_ ;
  assign \new_[29276]_  = \new_[29275]_  & \new_[29270]_ ;
  assign \new_[29280]_  = A167 & ~A168;
  assign \new_[29281]_  = A169 & \new_[29280]_ ;
  assign \new_[29285]_  = A200 & ~A199;
  assign \new_[29286]_  = ~A166 & \new_[29285]_ ;
  assign \new_[29287]_  = \new_[29286]_  & \new_[29281]_ ;
  assign \new_[29291]_  = ~A265 & ~A234;
  assign \new_[29292]_  = ~A233 & \new_[29291]_ ;
  assign \new_[29296]_  = ~A299 & ~A298;
  assign \new_[29297]_  = ~A266 & \new_[29296]_ ;
  assign \new_[29298]_  = \new_[29297]_  & \new_[29292]_ ;
  assign \new_[29302]_  = A167 & ~A168;
  assign \new_[29303]_  = A169 & \new_[29302]_ ;
  assign \new_[29307]_  = A200 & ~A199;
  assign \new_[29308]_  = ~A166 & \new_[29307]_ ;
  assign \new_[29309]_  = \new_[29308]_  & \new_[29303]_ ;
  assign \new_[29313]_  = A234 & ~A233;
  assign \new_[29314]_  = A232 & \new_[29313]_ ;
  assign \new_[29318]_  = A299 & ~A298;
  assign \new_[29319]_  = A235 & \new_[29318]_ ;
  assign \new_[29320]_  = \new_[29319]_  & \new_[29314]_ ;
  assign \new_[29324]_  = A167 & ~A168;
  assign \new_[29325]_  = A169 & \new_[29324]_ ;
  assign \new_[29329]_  = A200 & ~A199;
  assign \new_[29330]_  = ~A166 & \new_[29329]_ ;
  assign \new_[29331]_  = \new_[29330]_  & \new_[29325]_ ;
  assign \new_[29335]_  = A234 & ~A233;
  assign \new_[29336]_  = A232 & \new_[29335]_ ;
  assign \new_[29340]_  = A266 & ~A265;
  assign \new_[29341]_  = A235 & \new_[29340]_ ;
  assign \new_[29342]_  = \new_[29341]_  & \new_[29336]_ ;
  assign \new_[29346]_  = A167 & ~A168;
  assign \new_[29347]_  = A169 & \new_[29346]_ ;
  assign \new_[29351]_  = A200 & ~A199;
  assign \new_[29352]_  = ~A166 & \new_[29351]_ ;
  assign \new_[29353]_  = \new_[29352]_  & \new_[29347]_ ;
  assign \new_[29357]_  = A234 & ~A233;
  assign \new_[29358]_  = A232 & \new_[29357]_ ;
  assign \new_[29362]_  = A299 & ~A298;
  assign \new_[29363]_  = A236 & \new_[29362]_ ;
  assign \new_[29364]_  = \new_[29363]_  & \new_[29358]_ ;
  assign \new_[29368]_  = A167 & ~A168;
  assign \new_[29369]_  = A169 & \new_[29368]_ ;
  assign \new_[29373]_  = A200 & ~A199;
  assign \new_[29374]_  = ~A166 & \new_[29373]_ ;
  assign \new_[29375]_  = \new_[29374]_  & \new_[29369]_ ;
  assign \new_[29379]_  = A234 & ~A233;
  assign \new_[29380]_  = A232 & \new_[29379]_ ;
  assign \new_[29384]_  = A266 & ~A265;
  assign \new_[29385]_  = A236 & \new_[29384]_ ;
  assign \new_[29386]_  = \new_[29385]_  & \new_[29380]_ ;
  assign \new_[29390]_  = A167 & ~A168;
  assign \new_[29391]_  = A169 & \new_[29390]_ ;
  assign \new_[29395]_  = A200 & ~A199;
  assign \new_[29396]_  = ~A166 & \new_[29395]_ ;
  assign \new_[29397]_  = \new_[29396]_  & \new_[29391]_ ;
  assign \new_[29401]_  = A265 & ~A233;
  assign \new_[29402]_  = ~A232 & \new_[29401]_ ;
  assign \new_[29406]_  = ~A300 & A298;
  assign \new_[29407]_  = A266 & \new_[29406]_ ;
  assign \new_[29408]_  = \new_[29407]_  & \new_[29402]_ ;
  assign \new_[29412]_  = A167 & ~A168;
  assign \new_[29413]_  = A169 & \new_[29412]_ ;
  assign \new_[29417]_  = A200 & ~A199;
  assign \new_[29418]_  = ~A166 & \new_[29417]_ ;
  assign \new_[29419]_  = \new_[29418]_  & \new_[29413]_ ;
  assign \new_[29423]_  = A265 & ~A233;
  assign \new_[29424]_  = ~A232 & \new_[29423]_ ;
  assign \new_[29428]_  = A299 & A298;
  assign \new_[29429]_  = A266 & \new_[29428]_ ;
  assign \new_[29430]_  = \new_[29429]_  & \new_[29424]_ ;
  assign \new_[29434]_  = A167 & ~A168;
  assign \new_[29435]_  = A169 & \new_[29434]_ ;
  assign \new_[29439]_  = A200 & ~A199;
  assign \new_[29440]_  = ~A166 & \new_[29439]_ ;
  assign \new_[29441]_  = \new_[29440]_  & \new_[29435]_ ;
  assign \new_[29445]_  = A265 & ~A233;
  assign \new_[29446]_  = ~A232 & \new_[29445]_ ;
  assign \new_[29450]_  = ~A299 & ~A298;
  assign \new_[29451]_  = A266 & \new_[29450]_ ;
  assign \new_[29452]_  = \new_[29451]_  & \new_[29446]_ ;
  assign \new_[29456]_  = A167 & ~A168;
  assign \new_[29457]_  = A169 & \new_[29456]_ ;
  assign \new_[29461]_  = A200 & ~A199;
  assign \new_[29462]_  = ~A166 & \new_[29461]_ ;
  assign \new_[29463]_  = \new_[29462]_  & \new_[29457]_ ;
  assign \new_[29467]_  = ~A266 & ~A233;
  assign \new_[29468]_  = ~A232 & \new_[29467]_ ;
  assign \new_[29472]_  = ~A300 & A298;
  assign \new_[29473]_  = ~A267 & \new_[29472]_ ;
  assign \new_[29474]_  = \new_[29473]_  & \new_[29468]_ ;
  assign \new_[29478]_  = A167 & ~A168;
  assign \new_[29479]_  = A169 & \new_[29478]_ ;
  assign \new_[29483]_  = A200 & ~A199;
  assign \new_[29484]_  = ~A166 & \new_[29483]_ ;
  assign \new_[29485]_  = \new_[29484]_  & \new_[29479]_ ;
  assign \new_[29489]_  = ~A266 & ~A233;
  assign \new_[29490]_  = ~A232 & \new_[29489]_ ;
  assign \new_[29494]_  = A299 & A298;
  assign \new_[29495]_  = ~A267 & \new_[29494]_ ;
  assign \new_[29496]_  = \new_[29495]_  & \new_[29490]_ ;
  assign \new_[29500]_  = A167 & ~A168;
  assign \new_[29501]_  = A169 & \new_[29500]_ ;
  assign \new_[29505]_  = A200 & ~A199;
  assign \new_[29506]_  = ~A166 & \new_[29505]_ ;
  assign \new_[29507]_  = \new_[29506]_  & \new_[29501]_ ;
  assign \new_[29511]_  = ~A266 & ~A233;
  assign \new_[29512]_  = ~A232 & \new_[29511]_ ;
  assign \new_[29516]_  = ~A299 & ~A298;
  assign \new_[29517]_  = ~A267 & \new_[29516]_ ;
  assign \new_[29518]_  = \new_[29517]_  & \new_[29512]_ ;
  assign \new_[29522]_  = A167 & ~A168;
  assign \new_[29523]_  = A169 & \new_[29522]_ ;
  assign \new_[29527]_  = A200 & ~A199;
  assign \new_[29528]_  = ~A166 & \new_[29527]_ ;
  assign \new_[29529]_  = \new_[29528]_  & \new_[29523]_ ;
  assign \new_[29533]_  = ~A265 & ~A233;
  assign \new_[29534]_  = ~A232 & \new_[29533]_ ;
  assign \new_[29538]_  = ~A300 & A298;
  assign \new_[29539]_  = ~A266 & \new_[29538]_ ;
  assign \new_[29540]_  = \new_[29539]_  & \new_[29534]_ ;
  assign \new_[29544]_  = A167 & ~A168;
  assign \new_[29545]_  = A169 & \new_[29544]_ ;
  assign \new_[29549]_  = A200 & ~A199;
  assign \new_[29550]_  = ~A166 & \new_[29549]_ ;
  assign \new_[29551]_  = \new_[29550]_  & \new_[29545]_ ;
  assign \new_[29555]_  = ~A265 & ~A233;
  assign \new_[29556]_  = ~A232 & \new_[29555]_ ;
  assign \new_[29560]_  = A299 & A298;
  assign \new_[29561]_  = ~A266 & \new_[29560]_ ;
  assign \new_[29562]_  = \new_[29561]_  & \new_[29556]_ ;
  assign \new_[29566]_  = A167 & ~A168;
  assign \new_[29567]_  = A169 & \new_[29566]_ ;
  assign \new_[29571]_  = A200 & ~A199;
  assign \new_[29572]_  = ~A166 & \new_[29571]_ ;
  assign \new_[29573]_  = \new_[29572]_  & \new_[29567]_ ;
  assign \new_[29577]_  = ~A265 & ~A233;
  assign \new_[29578]_  = ~A232 & \new_[29577]_ ;
  assign \new_[29582]_  = ~A299 & ~A298;
  assign \new_[29583]_  = ~A266 & \new_[29582]_ ;
  assign \new_[29584]_  = \new_[29583]_  & \new_[29578]_ ;
  assign \new_[29588]_  = A167 & ~A168;
  assign \new_[29589]_  = A169 & \new_[29588]_ ;
  assign \new_[29593]_  = ~A200 & A199;
  assign \new_[29594]_  = ~A166 & \new_[29593]_ ;
  assign \new_[29595]_  = \new_[29594]_  & \new_[29589]_ ;
  assign \new_[29599]_  = ~A232 & A202;
  assign \new_[29600]_  = A201 & \new_[29599]_ ;
  assign \new_[29604]_  = A299 & ~A298;
  assign \new_[29605]_  = A233 & \new_[29604]_ ;
  assign \new_[29606]_  = \new_[29605]_  & \new_[29600]_ ;
  assign \new_[29610]_  = A167 & ~A168;
  assign \new_[29611]_  = A169 & \new_[29610]_ ;
  assign \new_[29615]_  = ~A200 & A199;
  assign \new_[29616]_  = ~A166 & \new_[29615]_ ;
  assign \new_[29617]_  = \new_[29616]_  & \new_[29611]_ ;
  assign \new_[29621]_  = ~A232 & A202;
  assign \new_[29622]_  = A201 & \new_[29621]_ ;
  assign \new_[29626]_  = A266 & ~A265;
  assign \new_[29627]_  = A233 & \new_[29626]_ ;
  assign \new_[29628]_  = \new_[29627]_  & \new_[29622]_ ;
  assign \new_[29632]_  = A167 & ~A168;
  assign \new_[29633]_  = A169 & \new_[29632]_ ;
  assign \new_[29637]_  = ~A200 & A199;
  assign \new_[29638]_  = ~A166 & \new_[29637]_ ;
  assign \new_[29639]_  = \new_[29638]_  & \new_[29633]_ ;
  assign \new_[29643]_  = ~A232 & A203;
  assign \new_[29644]_  = A201 & \new_[29643]_ ;
  assign \new_[29648]_  = A299 & ~A298;
  assign \new_[29649]_  = A233 & \new_[29648]_ ;
  assign \new_[29650]_  = \new_[29649]_  & \new_[29644]_ ;
  assign \new_[29654]_  = A167 & ~A168;
  assign \new_[29655]_  = A169 & \new_[29654]_ ;
  assign \new_[29659]_  = ~A200 & A199;
  assign \new_[29660]_  = ~A166 & \new_[29659]_ ;
  assign \new_[29661]_  = \new_[29660]_  & \new_[29655]_ ;
  assign \new_[29665]_  = ~A232 & A203;
  assign \new_[29666]_  = A201 & \new_[29665]_ ;
  assign \new_[29670]_  = A266 & ~A265;
  assign \new_[29671]_  = A233 & \new_[29670]_ ;
  assign \new_[29672]_  = \new_[29671]_  & \new_[29666]_ ;
  assign \new_[29676]_  = ~A167 & ~A168;
  assign \new_[29677]_  = A169 & \new_[29676]_ ;
  assign \new_[29681]_  = A200 & ~A199;
  assign \new_[29682]_  = A166 & \new_[29681]_ ;
  assign \new_[29683]_  = \new_[29682]_  & \new_[29677]_ ;
  assign \new_[29687]_  = A265 & A233;
  assign \new_[29688]_  = A232 & \new_[29687]_ ;
  assign \new_[29692]_  = ~A300 & ~A299;
  assign \new_[29693]_  = ~A267 & \new_[29692]_ ;
  assign \new_[29694]_  = \new_[29693]_  & \new_[29688]_ ;
  assign \new_[29698]_  = ~A167 & ~A168;
  assign \new_[29699]_  = A169 & \new_[29698]_ ;
  assign \new_[29703]_  = A200 & ~A199;
  assign \new_[29704]_  = A166 & \new_[29703]_ ;
  assign \new_[29705]_  = \new_[29704]_  & \new_[29699]_ ;
  assign \new_[29709]_  = A265 & A233;
  assign \new_[29710]_  = A232 & \new_[29709]_ ;
  assign \new_[29714]_  = A299 & A298;
  assign \new_[29715]_  = ~A267 & \new_[29714]_ ;
  assign \new_[29716]_  = \new_[29715]_  & \new_[29710]_ ;
  assign \new_[29720]_  = ~A167 & ~A168;
  assign \new_[29721]_  = A169 & \new_[29720]_ ;
  assign \new_[29725]_  = A200 & ~A199;
  assign \new_[29726]_  = A166 & \new_[29725]_ ;
  assign \new_[29727]_  = \new_[29726]_  & \new_[29721]_ ;
  assign \new_[29731]_  = A265 & A233;
  assign \new_[29732]_  = A232 & \new_[29731]_ ;
  assign \new_[29736]_  = ~A299 & ~A298;
  assign \new_[29737]_  = ~A267 & \new_[29736]_ ;
  assign \new_[29738]_  = \new_[29737]_  & \new_[29732]_ ;
  assign \new_[29742]_  = ~A167 & ~A168;
  assign \new_[29743]_  = A169 & \new_[29742]_ ;
  assign \new_[29747]_  = A200 & ~A199;
  assign \new_[29748]_  = A166 & \new_[29747]_ ;
  assign \new_[29749]_  = \new_[29748]_  & \new_[29743]_ ;
  assign \new_[29753]_  = A265 & A233;
  assign \new_[29754]_  = A232 & \new_[29753]_ ;
  assign \new_[29758]_  = ~A300 & ~A299;
  assign \new_[29759]_  = A266 & \new_[29758]_ ;
  assign \new_[29760]_  = \new_[29759]_  & \new_[29754]_ ;
  assign \new_[29764]_  = ~A167 & ~A168;
  assign \new_[29765]_  = A169 & \new_[29764]_ ;
  assign \new_[29769]_  = A200 & ~A199;
  assign \new_[29770]_  = A166 & \new_[29769]_ ;
  assign \new_[29771]_  = \new_[29770]_  & \new_[29765]_ ;
  assign \new_[29775]_  = A265 & A233;
  assign \new_[29776]_  = A232 & \new_[29775]_ ;
  assign \new_[29780]_  = A299 & A298;
  assign \new_[29781]_  = A266 & \new_[29780]_ ;
  assign \new_[29782]_  = \new_[29781]_  & \new_[29776]_ ;
  assign \new_[29786]_  = ~A167 & ~A168;
  assign \new_[29787]_  = A169 & \new_[29786]_ ;
  assign \new_[29791]_  = A200 & ~A199;
  assign \new_[29792]_  = A166 & \new_[29791]_ ;
  assign \new_[29793]_  = \new_[29792]_  & \new_[29787]_ ;
  assign \new_[29797]_  = A265 & A233;
  assign \new_[29798]_  = A232 & \new_[29797]_ ;
  assign \new_[29802]_  = ~A299 & ~A298;
  assign \new_[29803]_  = A266 & \new_[29802]_ ;
  assign \new_[29804]_  = \new_[29803]_  & \new_[29798]_ ;
  assign \new_[29808]_  = ~A167 & ~A168;
  assign \new_[29809]_  = A169 & \new_[29808]_ ;
  assign \new_[29813]_  = A200 & ~A199;
  assign \new_[29814]_  = A166 & \new_[29813]_ ;
  assign \new_[29815]_  = \new_[29814]_  & \new_[29809]_ ;
  assign \new_[29819]_  = ~A265 & A233;
  assign \new_[29820]_  = A232 & \new_[29819]_ ;
  assign \new_[29824]_  = ~A300 & ~A299;
  assign \new_[29825]_  = ~A266 & \new_[29824]_ ;
  assign \new_[29826]_  = \new_[29825]_  & \new_[29820]_ ;
  assign \new_[29830]_  = ~A167 & ~A168;
  assign \new_[29831]_  = A169 & \new_[29830]_ ;
  assign \new_[29835]_  = A200 & ~A199;
  assign \new_[29836]_  = A166 & \new_[29835]_ ;
  assign \new_[29837]_  = \new_[29836]_  & \new_[29831]_ ;
  assign \new_[29841]_  = ~A265 & A233;
  assign \new_[29842]_  = A232 & \new_[29841]_ ;
  assign \new_[29846]_  = A299 & A298;
  assign \new_[29847]_  = ~A266 & \new_[29846]_ ;
  assign \new_[29848]_  = \new_[29847]_  & \new_[29842]_ ;
  assign \new_[29852]_  = ~A167 & ~A168;
  assign \new_[29853]_  = A169 & \new_[29852]_ ;
  assign \new_[29857]_  = A200 & ~A199;
  assign \new_[29858]_  = A166 & \new_[29857]_ ;
  assign \new_[29859]_  = \new_[29858]_  & \new_[29853]_ ;
  assign \new_[29863]_  = ~A265 & A233;
  assign \new_[29864]_  = A232 & \new_[29863]_ ;
  assign \new_[29868]_  = ~A299 & ~A298;
  assign \new_[29869]_  = ~A266 & \new_[29868]_ ;
  assign \new_[29870]_  = \new_[29869]_  & \new_[29864]_ ;
  assign \new_[29874]_  = ~A167 & ~A168;
  assign \new_[29875]_  = A169 & \new_[29874]_ ;
  assign \new_[29879]_  = A200 & ~A199;
  assign \new_[29880]_  = A166 & \new_[29879]_ ;
  assign \new_[29881]_  = \new_[29880]_  & \new_[29875]_ ;
  assign \new_[29885]_  = A298 & A233;
  assign \new_[29886]_  = ~A232 & \new_[29885]_ ;
  assign \new_[29890]_  = A301 & A300;
  assign \new_[29891]_  = ~A299 & \new_[29890]_ ;
  assign \new_[29892]_  = \new_[29891]_  & \new_[29886]_ ;
  assign \new_[29896]_  = ~A167 & ~A168;
  assign \new_[29897]_  = A169 & \new_[29896]_ ;
  assign \new_[29901]_  = A200 & ~A199;
  assign \new_[29902]_  = A166 & \new_[29901]_ ;
  assign \new_[29903]_  = \new_[29902]_  & \new_[29897]_ ;
  assign \new_[29907]_  = A298 & A233;
  assign \new_[29908]_  = ~A232 & \new_[29907]_ ;
  assign \new_[29912]_  = A302 & A300;
  assign \new_[29913]_  = ~A299 & \new_[29912]_ ;
  assign \new_[29914]_  = \new_[29913]_  & \new_[29908]_ ;
  assign \new_[29918]_  = ~A167 & ~A168;
  assign \new_[29919]_  = A169 & \new_[29918]_ ;
  assign \new_[29923]_  = A200 & ~A199;
  assign \new_[29924]_  = A166 & \new_[29923]_ ;
  assign \new_[29925]_  = \new_[29924]_  & \new_[29919]_ ;
  assign \new_[29929]_  = A265 & A233;
  assign \new_[29930]_  = ~A232 & \new_[29929]_ ;
  assign \new_[29934]_  = A268 & A267;
  assign \new_[29935]_  = ~A266 & \new_[29934]_ ;
  assign \new_[29936]_  = \new_[29935]_  & \new_[29930]_ ;
  assign \new_[29940]_  = ~A167 & ~A168;
  assign \new_[29941]_  = A169 & \new_[29940]_ ;
  assign \new_[29945]_  = A200 & ~A199;
  assign \new_[29946]_  = A166 & \new_[29945]_ ;
  assign \new_[29947]_  = \new_[29946]_  & \new_[29941]_ ;
  assign \new_[29951]_  = A265 & A233;
  assign \new_[29952]_  = ~A232 & \new_[29951]_ ;
  assign \new_[29956]_  = A269 & A267;
  assign \new_[29957]_  = ~A266 & \new_[29956]_ ;
  assign \new_[29958]_  = \new_[29957]_  & \new_[29952]_ ;
  assign \new_[29962]_  = ~A167 & ~A168;
  assign \new_[29963]_  = A169 & \new_[29962]_ ;
  assign \new_[29967]_  = A200 & ~A199;
  assign \new_[29968]_  = A166 & \new_[29967]_ ;
  assign \new_[29969]_  = \new_[29968]_  & \new_[29963]_ ;
  assign \new_[29973]_  = A265 & ~A234;
  assign \new_[29974]_  = ~A233 & \new_[29973]_ ;
  assign \new_[29978]_  = ~A300 & A298;
  assign \new_[29979]_  = A266 & \new_[29978]_ ;
  assign \new_[29980]_  = \new_[29979]_  & \new_[29974]_ ;
  assign \new_[29984]_  = ~A167 & ~A168;
  assign \new_[29985]_  = A169 & \new_[29984]_ ;
  assign \new_[29989]_  = A200 & ~A199;
  assign \new_[29990]_  = A166 & \new_[29989]_ ;
  assign \new_[29991]_  = \new_[29990]_  & \new_[29985]_ ;
  assign \new_[29995]_  = A265 & ~A234;
  assign \new_[29996]_  = ~A233 & \new_[29995]_ ;
  assign \new_[30000]_  = A299 & A298;
  assign \new_[30001]_  = A266 & \new_[30000]_ ;
  assign \new_[30002]_  = \new_[30001]_  & \new_[29996]_ ;
  assign \new_[30006]_  = ~A167 & ~A168;
  assign \new_[30007]_  = A169 & \new_[30006]_ ;
  assign \new_[30011]_  = A200 & ~A199;
  assign \new_[30012]_  = A166 & \new_[30011]_ ;
  assign \new_[30013]_  = \new_[30012]_  & \new_[30007]_ ;
  assign \new_[30017]_  = A265 & ~A234;
  assign \new_[30018]_  = ~A233 & \new_[30017]_ ;
  assign \new_[30022]_  = ~A299 & ~A298;
  assign \new_[30023]_  = A266 & \new_[30022]_ ;
  assign \new_[30024]_  = \new_[30023]_  & \new_[30018]_ ;
  assign \new_[30028]_  = ~A167 & ~A168;
  assign \new_[30029]_  = A169 & \new_[30028]_ ;
  assign \new_[30033]_  = A200 & ~A199;
  assign \new_[30034]_  = A166 & \new_[30033]_ ;
  assign \new_[30035]_  = \new_[30034]_  & \new_[30029]_ ;
  assign \new_[30039]_  = ~A266 & ~A234;
  assign \new_[30040]_  = ~A233 & \new_[30039]_ ;
  assign \new_[30044]_  = ~A300 & A298;
  assign \new_[30045]_  = ~A267 & \new_[30044]_ ;
  assign \new_[30046]_  = \new_[30045]_  & \new_[30040]_ ;
  assign \new_[30050]_  = ~A167 & ~A168;
  assign \new_[30051]_  = A169 & \new_[30050]_ ;
  assign \new_[30055]_  = A200 & ~A199;
  assign \new_[30056]_  = A166 & \new_[30055]_ ;
  assign \new_[30057]_  = \new_[30056]_  & \new_[30051]_ ;
  assign \new_[30061]_  = ~A266 & ~A234;
  assign \new_[30062]_  = ~A233 & \new_[30061]_ ;
  assign \new_[30066]_  = A299 & A298;
  assign \new_[30067]_  = ~A267 & \new_[30066]_ ;
  assign \new_[30068]_  = \new_[30067]_  & \new_[30062]_ ;
  assign \new_[30072]_  = ~A167 & ~A168;
  assign \new_[30073]_  = A169 & \new_[30072]_ ;
  assign \new_[30077]_  = A200 & ~A199;
  assign \new_[30078]_  = A166 & \new_[30077]_ ;
  assign \new_[30079]_  = \new_[30078]_  & \new_[30073]_ ;
  assign \new_[30083]_  = ~A266 & ~A234;
  assign \new_[30084]_  = ~A233 & \new_[30083]_ ;
  assign \new_[30088]_  = ~A299 & ~A298;
  assign \new_[30089]_  = ~A267 & \new_[30088]_ ;
  assign \new_[30090]_  = \new_[30089]_  & \new_[30084]_ ;
  assign \new_[30094]_  = ~A167 & ~A168;
  assign \new_[30095]_  = A169 & \new_[30094]_ ;
  assign \new_[30099]_  = A200 & ~A199;
  assign \new_[30100]_  = A166 & \new_[30099]_ ;
  assign \new_[30101]_  = \new_[30100]_  & \new_[30095]_ ;
  assign \new_[30105]_  = ~A265 & ~A234;
  assign \new_[30106]_  = ~A233 & \new_[30105]_ ;
  assign \new_[30110]_  = ~A300 & A298;
  assign \new_[30111]_  = ~A266 & \new_[30110]_ ;
  assign \new_[30112]_  = \new_[30111]_  & \new_[30106]_ ;
  assign \new_[30116]_  = ~A167 & ~A168;
  assign \new_[30117]_  = A169 & \new_[30116]_ ;
  assign \new_[30121]_  = A200 & ~A199;
  assign \new_[30122]_  = A166 & \new_[30121]_ ;
  assign \new_[30123]_  = \new_[30122]_  & \new_[30117]_ ;
  assign \new_[30127]_  = ~A265 & ~A234;
  assign \new_[30128]_  = ~A233 & \new_[30127]_ ;
  assign \new_[30132]_  = A299 & A298;
  assign \new_[30133]_  = ~A266 & \new_[30132]_ ;
  assign \new_[30134]_  = \new_[30133]_  & \new_[30128]_ ;
  assign \new_[30138]_  = ~A167 & ~A168;
  assign \new_[30139]_  = A169 & \new_[30138]_ ;
  assign \new_[30143]_  = A200 & ~A199;
  assign \new_[30144]_  = A166 & \new_[30143]_ ;
  assign \new_[30145]_  = \new_[30144]_  & \new_[30139]_ ;
  assign \new_[30149]_  = ~A265 & ~A234;
  assign \new_[30150]_  = ~A233 & \new_[30149]_ ;
  assign \new_[30154]_  = ~A299 & ~A298;
  assign \new_[30155]_  = ~A266 & \new_[30154]_ ;
  assign \new_[30156]_  = \new_[30155]_  & \new_[30150]_ ;
  assign \new_[30160]_  = ~A167 & ~A168;
  assign \new_[30161]_  = A169 & \new_[30160]_ ;
  assign \new_[30165]_  = A200 & ~A199;
  assign \new_[30166]_  = A166 & \new_[30165]_ ;
  assign \new_[30167]_  = \new_[30166]_  & \new_[30161]_ ;
  assign \new_[30171]_  = A234 & ~A233;
  assign \new_[30172]_  = A232 & \new_[30171]_ ;
  assign \new_[30176]_  = A299 & ~A298;
  assign \new_[30177]_  = A235 & \new_[30176]_ ;
  assign \new_[30178]_  = \new_[30177]_  & \new_[30172]_ ;
  assign \new_[30182]_  = ~A167 & ~A168;
  assign \new_[30183]_  = A169 & \new_[30182]_ ;
  assign \new_[30187]_  = A200 & ~A199;
  assign \new_[30188]_  = A166 & \new_[30187]_ ;
  assign \new_[30189]_  = \new_[30188]_  & \new_[30183]_ ;
  assign \new_[30193]_  = A234 & ~A233;
  assign \new_[30194]_  = A232 & \new_[30193]_ ;
  assign \new_[30198]_  = A266 & ~A265;
  assign \new_[30199]_  = A235 & \new_[30198]_ ;
  assign \new_[30200]_  = \new_[30199]_  & \new_[30194]_ ;
  assign \new_[30204]_  = ~A167 & ~A168;
  assign \new_[30205]_  = A169 & \new_[30204]_ ;
  assign \new_[30209]_  = A200 & ~A199;
  assign \new_[30210]_  = A166 & \new_[30209]_ ;
  assign \new_[30211]_  = \new_[30210]_  & \new_[30205]_ ;
  assign \new_[30215]_  = A234 & ~A233;
  assign \new_[30216]_  = A232 & \new_[30215]_ ;
  assign \new_[30220]_  = A299 & ~A298;
  assign \new_[30221]_  = A236 & \new_[30220]_ ;
  assign \new_[30222]_  = \new_[30221]_  & \new_[30216]_ ;
  assign \new_[30226]_  = ~A167 & ~A168;
  assign \new_[30227]_  = A169 & \new_[30226]_ ;
  assign \new_[30231]_  = A200 & ~A199;
  assign \new_[30232]_  = A166 & \new_[30231]_ ;
  assign \new_[30233]_  = \new_[30232]_  & \new_[30227]_ ;
  assign \new_[30237]_  = A234 & ~A233;
  assign \new_[30238]_  = A232 & \new_[30237]_ ;
  assign \new_[30242]_  = A266 & ~A265;
  assign \new_[30243]_  = A236 & \new_[30242]_ ;
  assign \new_[30244]_  = \new_[30243]_  & \new_[30238]_ ;
  assign \new_[30248]_  = ~A167 & ~A168;
  assign \new_[30249]_  = A169 & \new_[30248]_ ;
  assign \new_[30253]_  = A200 & ~A199;
  assign \new_[30254]_  = A166 & \new_[30253]_ ;
  assign \new_[30255]_  = \new_[30254]_  & \new_[30249]_ ;
  assign \new_[30259]_  = A265 & ~A233;
  assign \new_[30260]_  = ~A232 & \new_[30259]_ ;
  assign \new_[30264]_  = ~A300 & A298;
  assign \new_[30265]_  = A266 & \new_[30264]_ ;
  assign \new_[30266]_  = \new_[30265]_  & \new_[30260]_ ;
  assign \new_[30270]_  = ~A167 & ~A168;
  assign \new_[30271]_  = A169 & \new_[30270]_ ;
  assign \new_[30275]_  = A200 & ~A199;
  assign \new_[30276]_  = A166 & \new_[30275]_ ;
  assign \new_[30277]_  = \new_[30276]_  & \new_[30271]_ ;
  assign \new_[30281]_  = A265 & ~A233;
  assign \new_[30282]_  = ~A232 & \new_[30281]_ ;
  assign \new_[30286]_  = A299 & A298;
  assign \new_[30287]_  = A266 & \new_[30286]_ ;
  assign \new_[30288]_  = \new_[30287]_  & \new_[30282]_ ;
  assign \new_[30292]_  = ~A167 & ~A168;
  assign \new_[30293]_  = A169 & \new_[30292]_ ;
  assign \new_[30297]_  = A200 & ~A199;
  assign \new_[30298]_  = A166 & \new_[30297]_ ;
  assign \new_[30299]_  = \new_[30298]_  & \new_[30293]_ ;
  assign \new_[30303]_  = A265 & ~A233;
  assign \new_[30304]_  = ~A232 & \new_[30303]_ ;
  assign \new_[30308]_  = ~A299 & ~A298;
  assign \new_[30309]_  = A266 & \new_[30308]_ ;
  assign \new_[30310]_  = \new_[30309]_  & \new_[30304]_ ;
  assign \new_[30314]_  = ~A167 & ~A168;
  assign \new_[30315]_  = A169 & \new_[30314]_ ;
  assign \new_[30319]_  = A200 & ~A199;
  assign \new_[30320]_  = A166 & \new_[30319]_ ;
  assign \new_[30321]_  = \new_[30320]_  & \new_[30315]_ ;
  assign \new_[30325]_  = ~A266 & ~A233;
  assign \new_[30326]_  = ~A232 & \new_[30325]_ ;
  assign \new_[30330]_  = ~A300 & A298;
  assign \new_[30331]_  = ~A267 & \new_[30330]_ ;
  assign \new_[30332]_  = \new_[30331]_  & \new_[30326]_ ;
  assign \new_[30336]_  = ~A167 & ~A168;
  assign \new_[30337]_  = A169 & \new_[30336]_ ;
  assign \new_[30341]_  = A200 & ~A199;
  assign \new_[30342]_  = A166 & \new_[30341]_ ;
  assign \new_[30343]_  = \new_[30342]_  & \new_[30337]_ ;
  assign \new_[30347]_  = ~A266 & ~A233;
  assign \new_[30348]_  = ~A232 & \new_[30347]_ ;
  assign \new_[30352]_  = A299 & A298;
  assign \new_[30353]_  = ~A267 & \new_[30352]_ ;
  assign \new_[30354]_  = \new_[30353]_  & \new_[30348]_ ;
  assign \new_[30358]_  = ~A167 & ~A168;
  assign \new_[30359]_  = A169 & \new_[30358]_ ;
  assign \new_[30363]_  = A200 & ~A199;
  assign \new_[30364]_  = A166 & \new_[30363]_ ;
  assign \new_[30365]_  = \new_[30364]_  & \new_[30359]_ ;
  assign \new_[30369]_  = ~A266 & ~A233;
  assign \new_[30370]_  = ~A232 & \new_[30369]_ ;
  assign \new_[30374]_  = ~A299 & ~A298;
  assign \new_[30375]_  = ~A267 & \new_[30374]_ ;
  assign \new_[30376]_  = \new_[30375]_  & \new_[30370]_ ;
  assign \new_[30380]_  = ~A167 & ~A168;
  assign \new_[30381]_  = A169 & \new_[30380]_ ;
  assign \new_[30385]_  = A200 & ~A199;
  assign \new_[30386]_  = A166 & \new_[30385]_ ;
  assign \new_[30387]_  = \new_[30386]_  & \new_[30381]_ ;
  assign \new_[30391]_  = ~A265 & ~A233;
  assign \new_[30392]_  = ~A232 & \new_[30391]_ ;
  assign \new_[30396]_  = ~A300 & A298;
  assign \new_[30397]_  = ~A266 & \new_[30396]_ ;
  assign \new_[30398]_  = \new_[30397]_  & \new_[30392]_ ;
  assign \new_[30402]_  = ~A167 & ~A168;
  assign \new_[30403]_  = A169 & \new_[30402]_ ;
  assign \new_[30407]_  = A200 & ~A199;
  assign \new_[30408]_  = A166 & \new_[30407]_ ;
  assign \new_[30409]_  = \new_[30408]_  & \new_[30403]_ ;
  assign \new_[30413]_  = ~A265 & ~A233;
  assign \new_[30414]_  = ~A232 & \new_[30413]_ ;
  assign \new_[30418]_  = A299 & A298;
  assign \new_[30419]_  = ~A266 & \new_[30418]_ ;
  assign \new_[30420]_  = \new_[30419]_  & \new_[30414]_ ;
  assign \new_[30424]_  = ~A167 & ~A168;
  assign \new_[30425]_  = A169 & \new_[30424]_ ;
  assign \new_[30429]_  = A200 & ~A199;
  assign \new_[30430]_  = A166 & \new_[30429]_ ;
  assign \new_[30431]_  = \new_[30430]_  & \new_[30425]_ ;
  assign \new_[30435]_  = ~A265 & ~A233;
  assign \new_[30436]_  = ~A232 & \new_[30435]_ ;
  assign \new_[30440]_  = ~A299 & ~A298;
  assign \new_[30441]_  = ~A266 & \new_[30440]_ ;
  assign \new_[30442]_  = \new_[30441]_  & \new_[30436]_ ;
  assign \new_[30446]_  = ~A167 & ~A168;
  assign \new_[30447]_  = A169 & \new_[30446]_ ;
  assign \new_[30451]_  = ~A200 & A199;
  assign \new_[30452]_  = A166 & \new_[30451]_ ;
  assign \new_[30453]_  = \new_[30452]_  & \new_[30447]_ ;
  assign \new_[30457]_  = ~A232 & A202;
  assign \new_[30458]_  = A201 & \new_[30457]_ ;
  assign \new_[30462]_  = A299 & ~A298;
  assign \new_[30463]_  = A233 & \new_[30462]_ ;
  assign \new_[30464]_  = \new_[30463]_  & \new_[30458]_ ;
  assign \new_[30468]_  = ~A167 & ~A168;
  assign \new_[30469]_  = A169 & \new_[30468]_ ;
  assign \new_[30473]_  = ~A200 & A199;
  assign \new_[30474]_  = A166 & \new_[30473]_ ;
  assign \new_[30475]_  = \new_[30474]_  & \new_[30469]_ ;
  assign \new_[30479]_  = ~A232 & A202;
  assign \new_[30480]_  = A201 & \new_[30479]_ ;
  assign \new_[30484]_  = A266 & ~A265;
  assign \new_[30485]_  = A233 & \new_[30484]_ ;
  assign \new_[30486]_  = \new_[30485]_  & \new_[30480]_ ;
  assign \new_[30490]_  = ~A167 & ~A168;
  assign \new_[30491]_  = A169 & \new_[30490]_ ;
  assign \new_[30495]_  = ~A200 & A199;
  assign \new_[30496]_  = A166 & \new_[30495]_ ;
  assign \new_[30497]_  = \new_[30496]_  & \new_[30491]_ ;
  assign \new_[30501]_  = ~A232 & A203;
  assign \new_[30502]_  = A201 & \new_[30501]_ ;
  assign \new_[30506]_  = A299 & ~A298;
  assign \new_[30507]_  = A233 & \new_[30506]_ ;
  assign \new_[30508]_  = \new_[30507]_  & \new_[30502]_ ;
  assign \new_[30512]_  = ~A167 & ~A168;
  assign \new_[30513]_  = A169 & \new_[30512]_ ;
  assign \new_[30517]_  = ~A200 & A199;
  assign \new_[30518]_  = A166 & \new_[30517]_ ;
  assign \new_[30519]_  = \new_[30518]_  & \new_[30513]_ ;
  assign \new_[30523]_  = ~A232 & A203;
  assign \new_[30524]_  = A201 & \new_[30523]_ ;
  assign \new_[30528]_  = A266 & ~A265;
  assign \new_[30529]_  = A233 & \new_[30528]_ ;
  assign \new_[30530]_  = \new_[30529]_  & \new_[30524]_ ;
  assign \new_[30534]_  = ~A168 & A169;
  assign \new_[30535]_  = A170 & \new_[30534]_ ;
  assign \new_[30539]_  = ~A200 & A199;
  assign \new_[30540]_  = A166 & \new_[30539]_ ;
  assign \new_[30541]_  = \new_[30540]_  & \new_[30535]_ ;
  assign \new_[30545]_  = ~A232 & A202;
  assign \new_[30546]_  = A201 & \new_[30545]_ ;
  assign \new_[30550]_  = A299 & ~A298;
  assign \new_[30551]_  = A233 & \new_[30550]_ ;
  assign \new_[30552]_  = \new_[30551]_  & \new_[30546]_ ;
  assign \new_[30556]_  = ~A168 & A169;
  assign \new_[30557]_  = A170 & \new_[30556]_ ;
  assign \new_[30561]_  = ~A200 & A199;
  assign \new_[30562]_  = A166 & \new_[30561]_ ;
  assign \new_[30563]_  = \new_[30562]_  & \new_[30557]_ ;
  assign \new_[30567]_  = ~A232 & A202;
  assign \new_[30568]_  = A201 & \new_[30567]_ ;
  assign \new_[30572]_  = A266 & ~A265;
  assign \new_[30573]_  = A233 & \new_[30572]_ ;
  assign \new_[30574]_  = \new_[30573]_  & \new_[30568]_ ;
  assign \new_[30578]_  = ~A168 & A169;
  assign \new_[30579]_  = A170 & \new_[30578]_ ;
  assign \new_[30583]_  = ~A200 & A199;
  assign \new_[30584]_  = A166 & \new_[30583]_ ;
  assign \new_[30585]_  = \new_[30584]_  & \new_[30579]_ ;
  assign \new_[30589]_  = ~A232 & A203;
  assign \new_[30590]_  = A201 & \new_[30589]_ ;
  assign \new_[30594]_  = A299 & ~A298;
  assign \new_[30595]_  = A233 & \new_[30594]_ ;
  assign \new_[30596]_  = \new_[30595]_  & \new_[30590]_ ;
  assign \new_[30600]_  = ~A168 & A169;
  assign \new_[30601]_  = A170 & \new_[30600]_ ;
  assign \new_[30605]_  = ~A200 & A199;
  assign \new_[30606]_  = A166 & \new_[30605]_ ;
  assign \new_[30607]_  = \new_[30606]_  & \new_[30601]_ ;
  assign \new_[30611]_  = ~A232 & A203;
  assign \new_[30612]_  = A201 & \new_[30611]_ ;
  assign \new_[30616]_  = A266 & ~A265;
  assign \new_[30617]_  = A233 & \new_[30616]_ ;
  assign \new_[30618]_  = \new_[30617]_  & \new_[30612]_ ;
  assign \new_[30622]_  = A167 & A169;
  assign \new_[30623]_  = ~A170 & \new_[30622]_ ;
  assign \new_[30627]_  = A200 & A199;
  assign \new_[30628]_  = A166 & \new_[30627]_ ;
  assign \new_[30629]_  = \new_[30628]_  & \new_[30623]_ ;
  assign \new_[30633]_  = A265 & A233;
  assign \new_[30634]_  = A232 & \new_[30633]_ ;
  assign \new_[30638]_  = ~A300 & ~A299;
  assign \new_[30639]_  = ~A267 & \new_[30638]_ ;
  assign \new_[30640]_  = \new_[30639]_  & \new_[30634]_ ;
  assign \new_[30644]_  = A167 & A169;
  assign \new_[30645]_  = ~A170 & \new_[30644]_ ;
  assign \new_[30649]_  = A200 & A199;
  assign \new_[30650]_  = A166 & \new_[30649]_ ;
  assign \new_[30651]_  = \new_[30650]_  & \new_[30645]_ ;
  assign \new_[30655]_  = A265 & A233;
  assign \new_[30656]_  = A232 & \new_[30655]_ ;
  assign \new_[30660]_  = A299 & A298;
  assign \new_[30661]_  = ~A267 & \new_[30660]_ ;
  assign \new_[30662]_  = \new_[30661]_  & \new_[30656]_ ;
  assign \new_[30666]_  = A167 & A169;
  assign \new_[30667]_  = ~A170 & \new_[30666]_ ;
  assign \new_[30671]_  = A200 & A199;
  assign \new_[30672]_  = A166 & \new_[30671]_ ;
  assign \new_[30673]_  = \new_[30672]_  & \new_[30667]_ ;
  assign \new_[30677]_  = A265 & A233;
  assign \new_[30678]_  = A232 & \new_[30677]_ ;
  assign \new_[30682]_  = ~A299 & ~A298;
  assign \new_[30683]_  = ~A267 & \new_[30682]_ ;
  assign \new_[30684]_  = \new_[30683]_  & \new_[30678]_ ;
  assign \new_[30688]_  = A167 & A169;
  assign \new_[30689]_  = ~A170 & \new_[30688]_ ;
  assign \new_[30693]_  = A200 & A199;
  assign \new_[30694]_  = A166 & \new_[30693]_ ;
  assign \new_[30695]_  = \new_[30694]_  & \new_[30689]_ ;
  assign \new_[30699]_  = A265 & A233;
  assign \new_[30700]_  = A232 & \new_[30699]_ ;
  assign \new_[30704]_  = ~A300 & ~A299;
  assign \new_[30705]_  = A266 & \new_[30704]_ ;
  assign \new_[30706]_  = \new_[30705]_  & \new_[30700]_ ;
  assign \new_[30710]_  = A167 & A169;
  assign \new_[30711]_  = ~A170 & \new_[30710]_ ;
  assign \new_[30715]_  = A200 & A199;
  assign \new_[30716]_  = A166 & \new_[30715]_ ;
  assign \new_[30717]_  = \new_[30716]_  & \new_[30711]_ ;
  assign \new_[30721]_  = A265 & A233;
  assign \new_[30722]_  = A232 & \new_[30721]_ ;
  assign \new_[30726]_  = A299 & A298;
  assign \new_[30727]_  = A266 & \new_[30726]_ ;
  assign \new_[30728]_  = \new_[30727]_  & \new_[30722]_ ;
  assign \new_[30732]_  = A167 & A169;
  assign \new_[30733]_  = ~A170 & \new_[30732]_ ;
  assign \new_[30737]_  = A200 & A199;
  assign \new_[30738]_  = A166 & \new_[30737]_ ;
  assign \new_[30739]_  = \new_[30738]_  & \new_[30733]_ ;
  assign \new_[30743]_  = A265 & A233;
  assign \new_[30744]_  = A232 & \new_[30743]_ ;
  assign \new_[30748]_  = ~A299 & ~A298;
  assign \new_[30749]_  = A266 & \new_[30748]_ ;
  assign \new_[30750]_  = \new_[30749]_  & \new_[30744]_ ;
  assign \new_[30754]_  = A167 & A169;
  assign \new_[30755]_  = ~A170 & \new_[30754]_ ;
  assign \new_[30759]_  = A200 & A199;
  assign \new_[30760]_  = A166 & \new_[30759]_ ;
  assign \new_[30761]_  = \new_[30760]_  & \new_[30755]_ ;
  assign \new_[30765]_  = ~A265 & A233;
  assign \new_[30766]_  = A232 & \new_[30765]_ ;
  assign \new_[30770]_  = ~A300 & ~A299;
  assign \new_[30771]_  = ~A266 & \new_[30770]_ ;
  assign \new_[30772]_  = \new_[30771]_  & \new_[30766]_ ;
  assign \new_[30776]_  = A167 & A169;
  assign \new_[30777]_  = ~A170 & \new_[30776]_ ;
  assign \new_[30781]_  = A200 & A199;
  assign \new_[30782]_  = A166 & \new_[30781]_ ;
  assign \new_[30783]_  = \new_[30782]_  & \new_[30777]_ ;
  assign \new_[30787]_  = ~A265 & A233;
  assign \new_[30788]_  = A232 & \new_[30787]_ ;
  assign \new_[30792]_  = A299 & A298;
  assign \new_[30793]_  = ~A266 & \new_[30792]_ ;
  assign \new_[30794]_  = \new_[30793]_  & \new_[30788]_ ;
  assign \new_[30798]_  = A167 & A169;
  assign \new_[30799]_  = ~A170 & \new_[30798]_ ;
  assign \new_[30803]_  = A200 & A199;
  assign \new_[30804]_  = A166 & \new_[30803]_ ;
  assign \new_[30805]_  = \new_[30804]_  & \new_[30799]_ ;
  assign \new_[30809]_  = ~A265 & A233;
  assign \new_[30810]_  = A232 & \new_[30809]_ ;
  assign \new_[30814]_  = ~A299 & ~A298;
  assign \new_[30815]_  = ~A266 & \new_[30814]_ ;
  assign \new_[30816]_  = \new_[30815]_  & \new_[30810]_ ;
  assign \new_[30820]_  = A167 & A169;
  assign \new_[30821]_  = ~A170 & \new_[30820]_ ;
  assign \new_[30825]_  = A200 & A199;
  assign \new_[30826]_  = A166 & \new_[30825]_ ;
  assign \new_[30827]_  = \new_[30826]_  & \new_[30821]_ ;
  assign \new_[30831]_  = A298 & A233;
  assign \new_[30832]_  = ~A232 & \new_[30831]_ ;
  assign \new_[30836]_  = A301 & A300;
  assign \new_[30837]_  = ~A299 & \new_[30836]_ ;
  assign \new_[30838]_  = \new_[30837]_  & \new_[30832]_ ;
  assign \new_[30842]_  = A167 & A169;
  assign \new_[30843]_  = ~A170 & \new_[30842]_ ;
  assign \new_[30847]_  = A200 & A199;
  assign \new_[30848]_  = A166 & \new_[30847]_ ;
  assign \new_[30849]_  = \new_[30848]_  & \new_[30843]_ ;
  assign \new_[30853]_  = A298 & A233;
  assign \new_[30854]_  = ~A232 & \new_[30853]_ ;
  assign \new_[30858]_  = A302 & A300;
  assign \new_[30859]_  = ~A299 & \new_[30858]_ ;
  assign \new_[30860]_  = \new_[30859]_  & \new_[30854]_ ;
  assign \new_[30864]_  = A167 & A169;
  assign \new_[30865]_  = ~A170 & \new_[30864]_ ;
  assign \new_[30869]_  = A200 & A199;
  assign \new_[30870]_  = A166 & \new_[30869]_ ;
  assign \new_[30871]_  = \new_[30870]_  & \new_[30865]_ ;
  assign \new_[30875]_  = A265 & A233;
  assign \new_[30876]_  = ~A232 & \new_[30875]_ ;
  assign \new_[30880]_  = A268 & A267;
  assign \new_[30881]_  = ~A266 & \new_[30880]_ ;
  assign \new_[30882]_  = \new_[30881]_  & \new_[30876]_ ;
  assign \new_[30886]_  = A167 & A169;
  assign \new_[30887]_  = ~A170 & \new_[30886]_ ;
  assign \new_[30891]_  = A200 & A199;
  assign \new_[30892]_  = A166 & \new_[30891]_ ;
  assign \new_[30893]_  = \new_[30892]_  & \new_[30887]_ ;
  assign \new_[30897]_  = A265 & A233;
  assign \new_[30898]_  = ~A232 & \new_[30897]_ ;
  assign \new_[30902]_  = A269 & A267;
  assign \new_[30903]_  = ~A266 & \new_[30902]_ ;
  assign \new_[30904]_  = \new_[30903]_  & \new_[30898]_ ;
  assign \new_[30908]_  = A167 & A169;
  assign \new_[30909]_  = ~A170 & \new_[30908]_ ;
  assign \new_[30913]_  = A200 & A199;
  assign \new_[30914]_  = A166 & \new_[30913]_ ;
  assign \new_[30915]_  = \new_[30914]_  & \new_[30909]_ ;
  assign \new_[30919]_  = A265 & ~A234;
  assign \new_[30920]_  = ~A233 & \new_[30919]_ ;
  assign \new_[30924]_  = ~A300 & A298;
  assign \new_[30925]_  = A266 & \new_[30924]_ ;
  assign \new_[30926]_  = \new_[30925]_  & \new_[30920]_ ;
  assign \new_[30930]_  = A167 & A169;
  assign \new_[30931]_  = ~A170 & \new_[30930]_ ;
  assign \new_[30935]_  = A200 & A199;
  assign \new_[30936]_  = A166 & \new_[30935]_ ;
  assign \new_[30937]_  = \new_[30936]_  & \new_[30931]_ ;
  assign \new_[30941]_  = A265 & ~A234;
  assign \new_[30942]_  = ~A233 & \new_[30941]_ ;
  assign \new_[30946]_  = A299 & A298;
  assign \new_[30947]_  = A266 & \new_[30946]_ ;
  assign \new_[30948]_  = \new_[30947]_  & \new_[30942]_ ;
  assign \new_[30952]_  = A167 & A169;
  assign \new_[30953]_  = ~A170 & \new_[30952]_ ;
  assign \new_[30957]_  = A200 & A199;
  assign \new_[30958]_  = A166 & \new_[30957]_ ;
  assign \new_[30959]_  = \new_[30958]_  & \new_[30953]_ ;
  assign \new_[30963]_  = A265 & ~A234;
  assign \new_[30964]_  = ~A233 & \new_[30963]_ ;
  assign \new_[30968]_  = ~A299 & ~A298;
  assign \new_[30969]_  = A266 & \new_[30968]_ ;
  assign \new_[30970]_  = \new_[30969]_  & \new_[30964]_ ;
  assign \new_[30974]_  = A167 & A169;
  assign \new_[30975]_  = ~A170 & \new_[30974]_ ;
  assign \new_[30979]_  = A200 & A199;
  assign \new_[30980]_  = A166 & \new_[30979]_ ;
  assign \new_[30981]_  = \new_[30980]_  & \new_[30975]_ ;
  assign \new_[30985]_  = ~A266 & ~A234;
  assign \new_[30986]_  = ~A233 & \new_[30985]_ ;
  assign \new_[30990]_  = ~A300 & A298;
  assign \new_[30991]_  = ~A267 & \new_[30990]_ ;
  assign \new_[30992]_  = \new_[30991]_  & \new_[30986]_ ;
  assign \new_[30996]_  = A167 & A169;
  assign \new_[30997]_  = ~A170 & \new_[30996]_ ;
  assign \new_[31001]_  = A200 & A199;
  assign \new_[31002]_  = A166 & \new_[31001]_ ;
  assign \new_[31003]_  = \new_[31002]_  & \new_[30997]_ ;
  assign \new_[31007]_  = ~A266 & ~A234;
  assign \new_[31008]_  = ~A233 & \new_[31007]_ ;
  assign \new_[31012]_  = A299 & A298;
  assign \new_[31013]_  = ~A267 & \new_[31012]_ ;
  assign \new_[31014]_  = \new_[31013]_  & \new_[31008]_ ;
  assign \new_[31018]_  = A167 & A169;
  assign \new_[31019]_  = ~A170 & \new_[31018]_ ;
  assign \new_[31023]_  = A200 & A199;
  assign \new_[31024]_  = A166 & \new_[31023]_ ;
  assign \new_[31025]_  = \new_[31024]_  & \new_[31019]_ ;
  assign \new_[31029]_  = ~A266 & ~A234;
  assign \new_[31030]_  = ~A233 & \new_[31029]_ ;
  assign \new_[31034]_  = ~A299 & ~A298;
  assign \new_[31035]_  = ~A267 & \new_[31034]_ ;
  assign \new_[31036]_  = \new_[31035]_  & \new_[31030]_ ;
  assign \new_[31040]_  = A167 & A169;
  assign \new_[31041]_  = ~A170 & \new_[31040]_ ;
  assign \new_[31045]_  = A200 & A199;
  assign \new_[31046]_  = A166 & \new_[31045]_ ;
  assign \new_[31047]_  = \new_[31046]_  & \new_[31041]_ ;
  assign \new_[31051]_  = ~A265 & ~A234;
  assign \new_[31052]_  = ~A233 & \new_[31051]_ ;
  assign \new_[31056]_  = ~A300 & A298;
  assign \new_[31057]_  = ~A266 & \new_[31056]_ ;
  assign \new_[31058]_  = \new_[31057]_  & \new_[31052]_ ;
  assign \new_[31062]_  = A167 & A169;
  assign \new_[31063]_  = ~A170 & \new_[31062]_ ;
  assign \new_[31067]_  = A200 & A199;
  assign \new_[31068]_  = A166 & \new_[31067]_ ;
  assign \new_[31069]_  = \new_[31068]_  & \new_[31063]_ ;
  assign \new_[31073]_  = ~A265 & ~A234;
  assign \new_[31074]_  = ~A233 & \new_[31073]_ ;
  assign \new_[31078]_  = A299 & A298;
  assign \new_[31079]_  = ~A266 & \new_[31078]_ ;
  assign \new_[31080]_  = \new_[31079]_  & \new_[31074]_ ;
  assign \new_[31084]_  = A167 & A169;
  assign \new_[31085]_  = ~A170 & \new_[31084]_ ;
  assign \new_[31089]_  = A200 & A199;
  assign \new_[31090]_  = A166 & \new_[31089]_ ;
  assign \new_[31091]_  = \new_[31090]_  & \new_[31085]_ ;
  assign \new_[31095]_  = ~A265 & ~A234;
  assign \new_[31096]_  = ~A233 & \new_[31095]_ ;
  assign \new_[31100]_  = ~A299 & ~A298;
  assign \new_[31101]_  = ~A266 & \new_[31100]_ ;
  assign \new_[31102]_  = \new_[31101]_  & \new_[31096]_ ;
  assign \new_[31106]_  = A167 & A169;
  assign \new_[31107]_  = ~A170 & \new_[31106]_ ;
  assign \new_[31111]_  = A200 & A199;
  assign \new_[31112]_  = A166 & \new_[31111]_ ;
  assign \new_[31113]_  = \new_[31112]_  & \new_[31107]_ ;
  assign \new_[31117]_  = A234 & ~A233;
  assign \new_[31118]_  = A232 & \new_[31117]_ ;
  assign \new_[31122]_  = A299 & ~A298;
  assign \new_[31123]_  = A235 & \new_[31122]_ ;
  assign \new_[31124]_  = \new_[31123]_  & \new_[31118]_ ;
  assign \new_[31128]_  = A167 & A169;
  assign \new_[31129]_  = ~A170 & \new_[31128]_ ;
  assign \new_[31133]_  = A200 & A199;
  assign \new_[31134]_  = A166 & \new_[31133]_ ;
  assign \new_[31135]_  = \new_[31134]_  & \new_[31129]_ ;
  assign \new_[31139]_  = A234 & ~A233;
  assign \new_[31140]_  = A232 & \new_[31139]_ ;
  assign \new_[31144]_  = A266 & ~A265;
  assign \new_[31145]_  = A235 & \new_[31144]_ ;
  assign \new_[31146]_  = \new_[31145]_  & \new_[31140]_ ;
  assign \new_[31150]_  = A167 & A169;
  assign \new_[31151]_  = ~A170 & \new_[31150]_ ;
  assign \new_[31155]_  = A200 & A199;
  assign \new_[31156]_  = A166 & \new_[31155]_ ;
  assign \new_[31157]_  = \new_[31156]_  & \new_[31151]_ ;
  assign \new_[31161]_  = A234 & ~A233;
  assign \new_[31162]_  = A232 & \new_[31161]_ ;
  assign \new_[31166]_  = A299 & ~A298;
  assign \new_[31167]_  = A236 & \new_[31166]_ ;
  assign \new_[31168]_  = \new_[31167]_  & \new_[31162]_ ;
  assign \new_[31172]_  = A167 & A169;
  assign \new_[31173]_  = ~A170 & \new_[31172]_ ;
  assign \new_[31177]_  = A200 & A199;
  assign \new_[31178]_  = A166 & \new_[31177]_ ;
  assign \new_[31179]_  = \new_[31178]_  & \new_[31173]_ ;
  assign \new_[31183]_  = A234 & ~A233;
  assign \new_[31184]_  = A232 & \new_[31183]_ ;
  assign \new_[31188]_  = A266 & ~A265;
  assign \new_[31189]_  = A236 & \new_[31188]_ ;
  assign \new_[31190]_  = \new_[31189]_  & \new_[31184]_ ;
  assign \new_[31194]_  = A167 & A169;
  assign \new_[31195]_  = ~A170 & \new_[31194]_ ;
  assign \new_[31199]_  = A200 & A199;
  assign \new_[31200]_  = A166 & \new_[31199]_ ;
  assign \new_[31201]_  = \new_[31200]_  & \new_[31195]_ ;
  assign \new_[31205]_  = A265 & ~A233;
  assign \new_[31206]_  = ~A232 & \new_[31205]_ ;
  assign \new_[31210]_  = ~A300 & A298;
  assign \new_[31211]_  = A266 & \new_[31210]_ ;
  assign \new_[31212]_  = \new_[31211]_  & \new_[31206]_ ;
  assign \new_[31216]_  = A167 & A169;
  assign \new_[31217]_  = ~A170 & \new_[31216]_ ;
  assign \new_[31221]_  = A200 & A199;
  assign \new_[31222]_  = A166 & \new_[31221]_ ;
  assign \new_[31223]_  = \new_[31222]_  & \new_[31217]_ ;
  assign \new_[31227]_  = A265 & ~A233;
  assign \new_[31228]_  = ~A232 & \new_[31227]_ ;
  assign \new_[31232]_  = A299 & A298;
  assign \new_[31233]_  = A266 & \new_[31232]_ ;
  assign \new_[31234]_  = \new_[31233]_  & \new_[31228]_ ;
  assign \new_[31238]_  = A167 & A169;
  assign \new_[31239]_  = ~A170 & \new_[31238]_ ;
  assign \new_[31243]_  = A200 & A199;
  assign \new_[31244]_  = A166 & \new_[31243]_ ;
  assign \new_[31245]_  = \new_[31244]_  & \new_[31239]_ ;
  assign \new_[31249]_  = A265 & ~A233;
  assign \new_[31250]_  = ~A232 & \new_[31249]_ ;
  assign \new_[31254]_  = ~A299 & ~A298;
  assign \new_[31255]_  = A266 & \new_[31254]_ ;
  assign \new_[31256]_  = \new_[31255]_  & \new_[31250]_ ;
  assign \new_[31260]_  = A167 & A169;
  assign \new_[31261]_  = ~A170 & \new_[31260]_ ;
  assign \new_[31265]_  = A200 & A199;
  assign \new_[31266]_  = A166 & \new_[31265]_ ;
  assign \new_[31267]_  = \new_[31266]_  & \new_[31261]_ ;
  assign \new_[31271]_  = ~A266 & ~A233;
  assign \new_[31272]_  = ~A232 & \new_[31271]_ ;
  assign \new_[31276]_  = ~A300 & A298;
  assign \new_[31277]_  = ~A267 & \new_[31276]_ ;
  assign \new_[31278]_  = \new_[31277]_  & \new_[31272]_ ;
  assign \new_[31282]_  = A167 & A169;
  assign \new_[31283]_  = ~A170 & \new_[31282]_ ;
  assign \new_[31287]_  = A200 & A199;
  assign \new_[31288]_  = A166 & \new_[31287]_ ;
  assign \new_[31289]_  = \new_[31288]_  & \new_[31283]_ ;
  assign \new_[31293]_  = ~A266 & ~A233;
  assign \new_[31294]_  = ~A232 & \new_[31293]_ ;
  assign \new_[31298]_  = A299 & A298;
  assign \new_[31299]_  = ~A267 & \new_[31298]_ ;
  assign \new_[31300]_  = \new_[31299]_  & \new_[31294]_ ;
  assign \new_[31304]_  = A167 & A169;
  assign \new_[31305]_  = ~A170 & \new_[31304]_ ;
  assign \new_[31309]_  = A200 & A199;
  assign \new_[31310]_  = A166 & \new_[31309]_ ;
  assign \new_[31311]_  = \new_[31310]_  & \new_[31305]_ ;
  assign \new_[31315]_  = ~A266 & ~A233;
  assign \new_[31316]_  = ~A232 & \new_[31315]_ ;
  assign \new_[31320]_  = ~A299 & ~A298;
  assign \new_[31321]_  = ~A267 & \new_[31320]_ ;
  assign \new_[31322]_  = \new_[31321]_  & \new_[31316]_ ;
  assign \new_[31326]_  = A167 & A169;
  assign \new_[31327]_  = ~A170 & \new_[31326]_ ;
  assign \new_[31331]_  = A200 & A199;
  assign \new_[31332]_  = A166 & \new_[31331]_ ;
  assign \new_[31333]_  = \new_[31332]_  & \new_[31327]_ ;
  assign \new_[31337]_  = ~A265 & ~A233;
  assign \new_[31338]_  = ~A232 & \new_[31337]_ ;
  assign \new_[31342]_  = ~A300 & A298;
  assign \new_[31343]_  = ~A266 & \new_[31342]_ ;
  assign \new_[31344]_  = \new_[31343]_  & \new_[31338]_ ;
  assign \new_[31348]_  = A167 & A169;
  assign \new_[31349]_  = ~A170 & \new_[31348]_ ;
  assign \new_[31353]_  = A200 & A199;
  assign \new_[31354]_  = A166 & \new_[31353]_ ;
  assign \new_[31355]_  = \new_[31354]_  & \new_[31349]_ ;
  assign \new_[31359]_  = ~A265 & ~A233;
  assign \new_[31360]_  = ~A232 & \new_[31359]_ ;
  assign \new_[31364]_  = A299 & A298;
  assign \new_[31365]_  = ~A266 & \new_[31364]_ ;
  assign \new_[31366]_  = \new_[31365]_  & \new_[31360]_ ;
  assign \new_[31370]_  = A167 & A169;
  assign \new_[31371]_  = ~A170 & \new_[31370]_ ;
  assign \new_[31375]_  = A200 & A199;
  assign \new_[31376]_  = A166 & \new_[31375]_ ;
  assign \new_[31377]_  = \new_[31376]_  & \new_[31371]_ ;
  assign \new_[31381]_  = ~A265 & ~A233;
  assign \new_[31382]_  = ~A232 & \new_[31381]_ ;
  assign \new_[31386]_  = ~A299 & ~A298;
  assign \new_[31387]_  = ~A266 & \new_[31386]_ ;
  assign \new_[31388]_  = \new_[31387]_  & \new_[31382]_ ;
  assign \new_[31392]_  = A167 & A169;
  assign \new_[31393]_  = ~A170 & \new_[31392]_ ;
  assign \new_[31397]_  = ~A201 & ~A200;
  assign \new_[31398]_  = A166 & \new_[31397]_ ;
  assign \new_[31399]_  = \new_[31398]_  & \new_[31393]_ ;
  assign \new_[31403]_  = A265 & A233;
  assign \new_[31404]_  = A232 & \new_[31403]_ ;
  assign \new_[31408]_  = ~A300 & ~A299;
  assign \new_[31409]_  = ~A267 & \new_[31408]_ ;
  assign \new_[31410]_  = \new_[31409]_  & \new_[31404]_ ;
  assign \new_[31414]_  = A167 & A169;
  assign \new_[31415]_  = ~A170 & \new_[31414]_ ;
  assign \new_[31419]_  = ~A201 & ~A200;
  assign \new_[31420]_  = A166 & \new_[31419]_ ;
  assign \new_[31421]_  = \new_[31420]_  & \new_[31415]_ ;
  assign \new_[31425]_  = A265 & A233;
  assign \new_[31426]_  = A232 & \new_[31425]_ ;
  assign \new_[31430]_  = A299 & A298;
  assign \new_[31431]_  = ~A267 & \new_[31430]_ ;
  assign \new_[31432]_  = \new_[31431]_  & \new_[31426]_ ;
  assign \new_[31436]_  = A167 & A169;
  assign \new_[31437]_  = ~A170 & \new_[31436]_ ;
  assign \new_[31441]_  = ~A201 & ~A200;
  assign \new_[31442]_  = A166 & \new_[31441]_ ;
  assign \new_[31443]_  = \new_[31442]_  & \new_[31437]_ ;
  assign \new_[31447]_  = A265 & A233;
  assign \new_[31448]_  = A232 & \new_[31447]_ ;
  assign \new_[31452]_  = ~A299 & ~A298;
  assign \new_[31453]_  = ~A267 & \new_[31452]_ ;
  assign \new_[31454]_  = \new_[31453]_  & \new_[31448]_ ;
  assign \new_[31458]_  = A167 & A169;
  assign \new_[31459]_  = ~A170 & \new_[31458]_ ;
  assign \new_[31463]_  = ~A201 & ~A200;
  assign \new_[31464]_  = A166 & \new_[31463]_ ;
  assign \new_[31465]_  = \new_[31464]_  & \new_[31459]_ ;
  assign \new_[31469]_  = A265 & A233;
  assign \new_[31470]_  = A232 & \new_[31469]_ ;
  assign \new_[31474]_  = ~A300 & ~A299;
  assign \new_[31475]_  = A266 & \new_[31474]_ ;
  assign \new_[31476]_  = \new_[31475]_  & \new_[31470]_ ;
  assign \new_[31480]_  = A167 & A169;
  assign \new_[31481]_  = ~A170 & \new_[31480]_ ;
  assign \new_[31485]_  = ~A201 & ~A200;
  assign \new_[31486]_  = A166 & \new_[31485]_ ;
  assign \new_[31487]_  = \new_[31486]_  & \new_[31481]_ ;
  assign \new_[31491]_  = A265 & A233;
  assign \new_[31492]_  = A232 & \new_[31491]_ ;
  assign \new_[31496]_  = A299 & A298;
  assign \new_[31497]_  = A266 & \new_[31496]_ ;
  assign \new_[31498]_  = \new_[31497]_  & \new_[31492]_ ;
  assign \new_[31502]_  = A167 & A169;
  assign \new_[31503]_  = ~A170 & \new_[31502]_ ;
  assign \new_[31507]_  = ~A201 & ~A200;
  assign \new_[31508]_  = A166 & \new_[31507]_ ;
  assign \new_[31509]_  = \new_[31508]_  & \new_[31503]_ ;
  assign \new_[31513]_  = A265 & A233;
  assign \new_[31514]_  = A232 & \new_[31513]_ ;
  assign \new_[31518]_  = ~A299 & ~A298;
  assign \new_[31519]_  = A266 & \new_[31518]_ ;
  assign \new_[31520]_  = \new_[31519]_  & \new_[31514]_ ;
  assign \new_[31524]_  = A167 & A169;
  assign \new_[31525]_  = ~A170 & \new_[31524]_ ;
  assign \new_[31529]_  = ~A201 & ~A200;
  assign \new_[31530]_  = A166 & \new_[31529]_ ;
  assign \new_[31531]_  = \new_[31530]_  & \new_[31525]_ ;
  assign \new_[31535]_  = ~A265 & A233;
  assign \new_[31536]_  = A232 & \new_[31535]_ ;
  assign \new_[31540]_  = ~A300 & ~A299;
  assign \new_[31541]_  = ~A266 & \new_[31540]_ ;
  assign \new_[31542]_  = \new_[31541]_  & \new_[31536]_ ;
  assign \new_[31546]_  = A167 & A169;
  assign \new_[31547]_  = ~A170 & \new_[31546]_ ;
  assign \new_[31551]_  = ~A201 & ~A200;
  assign \new_[31552]_  = A166 & \new_[31551]_ ;
  assign \new_[31553]_  = \new_[31552]_  & \new_[31547]_ ;
  assign \new_[31557]_  = ~A265 & A233;
  assign \new_[31558]_  = A232 & \new_[31557]_ ;
  assign \new_[31562]_  = A299 & A298;
  assign \new_[31563]_  = ~A266 & \new_[31562]_ ;
  assign \new_[31564]_  = \new_[31563]_  & \new_[31558]_ ;
  assign \new_[31568]_  = A167 & A169;
  assign \new_[31569]_  = ~A170 & \new_[31568]_ ;
  assign \new_[31573]_  = ~A201 & ~A200;
  assign \new_[31574]_  = A166 & \new_[31573]_ ;
  assign \new_[31575]_  = \new_[31574]_  & \new_[31569]_ ;
  assign \new_[31579]_  = ~A265 & A233;
  assign \new_[31580]_  = A232 & \new_[31579]_ ;
  assign \new_[31584]_  = ~A299 & ~A298;
  assign \new_[31585]_  = ~A266 & \new_[31584]_ ;
  assign \new_[31586]_  = \new_[31585]_  & \new_[31580]_ ;
  assign \new_[31590]_  = A167 & A169;
  assign \new_[31591]_  = ~A170 & \new_[31590]_ ;
  assign \new_[31595]_  = ~A201 & ~A200;
  assign \new_[31596]_  = A166 & \new_[31595]_ ;
  assign \new_[31597]_  = \new_[31596]_  & \new_[31591]_ ;
  assign \new_[31601]_  = A298 & A233;
  assign \new_[31602]_  = ~A232 & \new_[31601]_ ;
  assign \new_[31606]_  = A301 & A300;
  assign \new_[31607]_  = ~A299 & \new_[31606]_ ;
  assign \new_[31608]_  = \new_[31607]_  & \new_[31602]_ ;
  assign \new_[31612]_  = A167 & A169;
  assign \new_[31613]_  = ~A170 & \new_[31612]_ ;
  assign \new_[31617]_  = ~A201 & ~A200;
  assign \new_[31618]_  = A166 & \new_[31617]_ ;
  assign \new_[31619]_  = \new_[31618]_  & \new_[31613]_ ;
  assign \new_[31623]_  = A298 & A233;
  assign \new_[31624]_  = ~A232 & \new_[31623]_ ;
  assign \new_[31628]_  = A302 & A300;
  assign \new_[31629]_  = ~A299 & \new_[31628]_ ;
  assign \new_[31630]_  = \new_[31629]_  & \new_[31624]_ ;
  assign \new_[31634]_  = A167 & A169;
  assign \new_[31635]_  = ~A170 & \new_[31634]_ ;
  assign \new_[31639]_  = ~A201 & ~A200;
  assign \new_[31640]_  = A166 & \new_[31639]_ ;
  assign \new_[31641]_  = \new_[31640]_  & \new_[31635]_ ;
  assign \new_[31645]_  = A265 & A233;
  assign \new_[31646]_  = ~A232 & \new_[31645]_ ;
  assign \new_[31650]_  = A268 & A267;
  assign \new_[31651]_  = ~A266 & \new_[31650]_ ;
  assign \new_[31652]_  = \new_[31651]_  & \new_[31646]_ ;
  assign \new_[31656]_  = A167 & A169;
  assign \new_[31657]_  = ~A170 & \new_[31656]_ ;
  assign \new_[31661]_  = ~A201 & ~A200;
  assign \new_[31662]_  = A166 & \new_[31661]_ ;
  assign \new_[31663]_  = \new_[31662]_  & \new_[31657]_ ;
  assign \new_[31667]_  = A265 & A233;
  assign \new_[31668]_  = ~A232 & \new_[31667]_ ;
  assign \new_[31672]_  = A269 & A267;
  assign \new_[31673]_  = ~A266 & \new_[31672]_ ;
  assign \new_[31674]_  = \new_[31673]_  & \new_[31668]_ ;
  assign \new_[31678]_  = A167 & A169;
  assign \new_[31679]_  = ~A170 & \new_[31678]_ ;
  assign \new_[31683]_  = ~A201 & ~A200;
  assign \new_[31684]_  = A166 & \new_[31683]_ ;
  assign \new_[31685]_  = \new_[31684]_  & \new_[31679]_ ;
  assign \new_[31689]_  = A265 & ~A234;
  assign \new_[31690]_  = ~A233 & \new_[31689]_ ;
  assign \new_[31694]_  = ~A300 & A298;
  assign \new_[31695]_  = A266 & \new_[31694]_ ;
  assign \new_[31696]_  = \new_[31695]_  & \new_[31690]_ ;
  assign \new_[31700]_  = A167 & A169;
  assign \new_[31701]_  = ~A170 & \new_[31700]_ ;
  assign \new_[31705]_  = ~A201 & ~A200;
  assign \new_[31706]_  = A166 & \new_[31705]_ ;
  assign \new_[31707]_  = \new_[31706]_  & \new_[31701]_ ;
  assign \new_[31711]_  = A265 & ~A234;
  assign \new_[31712]_  = ~A233 & \new_[31711]_ ;
  assign \new_[31716]_  = A299 & A298;
  assign \new_[31717]_  = A266 & \new_[31716]_ ;
  assign \new_[31718]_  = \new_[31717]_  & \new_[31712]_ ;
  assign \new_[31722]_  = A167 & A169;
  assign \new_[31723]_  = ~A170 & \new_[31722]_ ;
  assign \new_[31727]_  = ~A201 & ~A200;
  assign \new_[31728]_  = A166 & \new_[31727]_ ;
  assign \new_[31729]_  = \new_[31728]_  & \new_[31723]_ ;
  assign \new_[31733]_  = A265 & ~A234;
  assign \new_[31734]_  = ~A233 & \new_[31733]_ ;
  assign \new_[31738]_  = ~A299 & ~A298;
  assign \new_[31739]_  = A266 & \new_[31738]_ ;
  assign \new_[31740]_  = \new_[31739]_  & \new_[31734]_ ;
  assign \new_[31744]_  = A167 & A169;
  assign \new_[31745]_  = ~A170 & \new_[31744]_ ;
  assign \new_[31749]_  = ~A201 & ~A200;
  assign \new_[31750]_  = A166 & \new_[31749]_ ;
  assign \new_[31751]_  = \new_[31750]_  & \new_[31745]_ ;
  assign \new_[31755]_  = ~A266 & ~A234;
  assign \new_[31756]_  = ~A233 & \new_[31755]_ ;
  assign \new_[31760]_  = ~A300 & A298;
  assign \new_[31761]_  = ~A267 & \new_[31760]_ ;
  assign \new_[31762]_  = \new_[31761]_  & \new_[31756]_ ;
  assign \new_[31766]_  = A167 & A169;
  assign \new_[31767]_  = ~A170 & \new_[31766]_ ;
  assign \new_[31771]_  = ~A201 & ~A200;
  assign \new_[31772]_  = A166 & \new_[31771]_ ;
  assign \new_[31773]_  = \new_[31772]_  & \new_[31767]_ ;
  assign \new_[31777]_  = ~A266 & ~A234;
  assign \new_[31778]_  = ~A233 & \new_[31777]_ ;
  assign \new_[31782]_  = A299 & A298;
  assign \new_[31783]_  = ~A267 & \new_[31782]_ ;
  assign \new_[31784]_  = \new_[31783]_  & \new_[31778]_ ;
  assign \new_[31788]_  = A167 & A169;
  assign \new_[31789]_  = ~A170 & \new_[31788]_ ;
  assign \new_[31793]_  = ~A201 & ~A200;
  assign \new_[31794]_  = A166 & \new_[31793]_ ;
  assign \new_[31795]_  = \new_[31794]_  & \new_[31789]_ ;
  assign \new_[31799]_  = ~A266 & ~A234;
  assign \new_[31800]_  = ~A233 & \new_[31799]_ ;
  assign \new_[31804]_  = ~A299 & ~A298;
  assign \new_[31805]_  = ~A267 & \new_[31804]_ ;
  assign \new_[31806]_  = \new_[31805]_  & \new_[31800]_ ;
  assign \new_[31810]_  = A167 & A169;
  assign \new_[31811]_  = ~A170 & \new_[31810]_ ;
  assign \new_[31815]_  = ~A201 & ~A200;
  assign \new_[31816]_  = A166 & \new_[31815]_ ;
  assign \new_[31817]_  = \new_[31816]_  & \new_[31811]_ ;
  assign \new_[31821]_  = ~A265 & ~A234;
  assign \new_[31822]_  = ~A233 & \new_[31821]_ ;
  assign \new_[31826]_  = ~A300 & A298;
  assign \new_[31827]_  = ~A266 & \new_[31826]_ ;
  assign \new_[31828]_  = \new_[31827]_  & \new_[31822]_ ;
  assign \new_[31832]_  = A167 & A169;
  assign \new_[31833]_  = ~A170 & \new_[31832]_ ;
  assign \new_[31837]_  = ~A201 & ~A200;
  assign \new_[31838]_  = A166 & \new_[31837]_ ;
  assign \new_[31839]_  = \new_[31838]_  & \new_[31833]_ ;
  assign \new_[31843]_  = ~A265 & ~A234;
  assign \new_[31844]_  = ~A233 & \new_[31843]_ ;
  assign \new_[31848]_  = A299 & A298;
  assign \new_[31849]_  = ~A266 & \new_[31848]_ ;
  assign \new_[31850]_  = \new_[31849]_  & \new_[31844]_ ;
  assign \new_[31854]_  = A167 & A169;
  assign \new_[31855]_  = ~A170 & \new_[31854]_ ;
  assign \new_[31859]_  = ~A201 & ~A200;
  assign \new_[31860]_  = A166 & \new_[31859]_ ;
  assign \new_[31861]_  = \new_[31860]_  & \new_[31855]_ ;
  assign \new_[31865]_  = ~A265 & ~A234;
  assign \new_[31866]_  = ~A233 & \new_[31865]_ ;
  assign \new_[31870]_  = ~A299 & ~A298;
  assign \new_[31871]_  = ~A266 & \new_[31870]_ ;
  assign \new_[31872]_  = \new_[31871]_  & \new_[31866]_ ;
  assign \new_[31876]_  = A167 & A169;
  assign \new_[31877]_  = ~A170 & \new_[31876]_ ;
  assign \new_[31881]_  = ~A201 & ~A200;
  assign \new_[31882]_  = A166 & \new_[31881]_ ;
  assign \new_[31883]_  = \new_[31882]_  & \new_[31877]_ ;
  assign \new_[31887]_  = A234 & ~A233;
  assign \new_[31888]_  = A232 & \new_[31887]_ ;
  assign \new_[31892]_  = A299 & ~A298;
  assign \new_[31893]_  = A235 & \new_[31892]_ ;
  assign \new_[31894]_  = \new_[31893]_  & \new_[31888]_ ;
  assign \new_[31898]_  = A167 & A169;
  assign \new_[31899]_  = ~A170 & \new_[31898]_ ;
  assign \new_[31903]_  = ~A201 & ~A200;
  assign \new_[31904]_  = A166 & \new_[31903]_ ;
  assign \new_[31905]_  = \new_[31904]_  & \new_[31899]_ ;
  assign \new_[31909]_  = A234 & ~A233;
  assign \new_[31910]_  = A232 & \new_[31909]_ ;
  assign \new_[31914]_  = A266 & ~A265;
  assign \new_[31915]_  = A235 & \new_[31914]_ ;
  assign \new_[31916]_  = \new_[31915]_  & \new_[31910]_ ;
  assign \new_[31920]_  = A167 & A169;
  assign \new_[31921]_  = ~A170 & \new_[31920]_ ;
  assign \new_[31925]_  = ~A201 & ~A200;
  assign \new_[31926]_  = A166 & \new_[31925]_ ;
  assign \new_[31927]_  = \new_[31926]_  & \new_[31921]_ ;
  assign \new_[31931]_  = A234 & ~A233;
  assign \new_[31932]_  = A232 & \new_[31931]_ ;
  assign \new_[31936]_  = A299 & ~A298;
  assign \new_[31937]_  = A236 & \new_[31936]_ ;
  assign \new_[31938]_  = \new_[31937]_  & \new_[31932]_ ;
  assign \new_[31942]_  = A167 & A169;
  assign \new_[31943]_  = ~A170 & \new_[31942]_ ;
  assign \new_[31947]_  = ~A201 & ~A200;
  assign \new_[31948]_  = A166 & \new_[31947]_ ;
  assign \new_[31949]_  = \new_[31948]_  & \new_[31943]_ ;
  assign \new_[31953]_  = A234 & ~A233;
  assign \new_[31954]_  = A232 & \new_[31953]_ ;
  assign \new_[31958]_  = A266 & ~A265;
  assign \new_[31959]_  = A236 & \new_[31958]_ ;
  assign \new_[31960]_  = \new_[31959]_  & \new_[31954]_ ;
  assign \new_[31964]_  = A167 & A169;
  assign \new_[31965]_  = ~A170 & \new_[31964]_ ;
  assign \new_[31969]_  = ~A201 & ~A200;
  assign \new_[31970]_  = A166 & \new_[31969]_ ;
  assign \new_[31971]_  = \new_[31970]_  & \new_[31965]_ ;
  assign \new_[31975]_  = A265 & ~A233;
  assign \new_[31976]_  = ~A232 & \new_[31975]_ ;
  assign \new_[31980]_  = ~A300 & A298;
  assign \new_[31981]_  = A266 & \new_[31980]_ ;
  assign \new_[31982]_  = \new_[31981]_  & \new_[31976]_ ;
  assign \new_[31986]_  = A167 & A169;
  assign \new_[31987]_  = ~A170 & \new_[31986]_ ;
  assign \new_[31991]_  = ~A201 & ~A200;
  assign \new_[31992]_  = A166 & \new_[31991]_ ;
  assign \new_[31993]_  = \new_[31992]_  & \new_[31987]_ ;
  assign \new_[31997]_  = A265 & ~A233;
  assign \new_[31998]_  = ~A232 & \new_[31997]_ ;
  assign \new_[32002]_  = A299 & A298;
  assign \new_[32003]_  = A266 & \new_[32002]_ ;
  assign \new_[32004]_  = \new_[32003]_  & \new_[31998]_ ;
  assign \new_[32008]_  = A167 & A169;
  assign \new_[32009]_  = ~A170 & \new_[32008]_ ;
  assign \new_[32013]_  = ~A201 & ~A200;
  assign \new_[32014]_  = A166 & \new_[32013]_ ;
  assign \new_[32015]_  = \new_[32014]_  & \new_[32009]_ ;
  assign \new_[32019]_  = A265 & ~A233;
  assign \new_[32020]_  = ~A232 & \new_[32019]_ ;
  assign \new_[32024]_  = ~A299 & ~A298;
  assign \new_[32025]_  = A266 & \new_[32024]_ ;
  assign \new_[32026]_  = \new_[32025]_  & \new_[32020]_ ;
  assign \new_[32030]_  = A167 & A169;
  assign \new_[32031]_  = ~A170 & \new_[32030]_ ;
  assign \new_[32035]_  = ~A201 & ~A200;
  assign \new_[32036]_  = A166 & \new_[32035]_ ;
  assign \new_[32037]_  = \new_[32036]_  & \new_[32031]_ ;
  assign \new_[32041]_  = ~A266 & ~A233;
  assign \new_[32042]_  = ~A232 & \new_[32041]_ ;
  assign \new_[32046]_  = ~A300 & A298;
  assign \new_[32047]_  = ~A267 & \new_[32046]_ ;
  assign \new_[32048]_  = \new_[32047]_  & \new_[32042]_ ;
  assign \new_[32052]_  = A167 & A169;
  assign \new_[32053]_  = ~A170 & \new_[32052]_ ;
  assign \new_[32057]_  = ~A201 & ~A200;
  assign \new_[32058]_  = A166 & \new_[32057]_ ;
  assign \new_[32059]_  = \new_[32058]_  & \new_[32053]_ ;
  assign \new_[32063]_  = ~A266 & ~A233;
  assign \new_[32064]_  = ~A232 & \new_[32063]_ ;
  assign \new_[32068]_  = A299 & A298;
  assign \new_[32069]_  = ~A267 & \new_[32068]_ ;
  assign \new_[32070]_  = \new_[32069]_  & \new_[32064]_ ;
  assign \new_[32074]_  = A167 & A169;
  assign \new_[32075]_  = ~A170 & \new_[32074]_ ;
  assign \new_[32079]_  = ~A201 & ~A200;
  assign \new_[32080]_  = A166 & \new_[32079]_ ;
  assign \new_[32081]_  = \new_[32080]_  & \new_[32075]_ ;
  assign \new_[32085]_  = ~A266 & ~A233;
  assign \new_[32086]_  = ~A232 & \new_[32085]_ ;
  assign \new_[32090]_  = ~A299 & ~A298;
  assign \new_[32091]_  = ~A267 & \new_[32090]_ ;
  assign \new_[32092]_  = \new_[32091]_  & \new_[32086]_ ;
  assign \new_[32096]_  = A167 & A169;
  assign \new_[32097]_  = ~A170 & \new_[32096]_ ;
  assign \new_[32101]_  = ~A201 & ~A200;
  assign \new_[32102]_  = A166 & \new_[32101]_ ;
  assign \new_[32103]_  = \new_[32102]_  & \new_[32097]_ ;
  assign \new_[32107]_  = ~A265 & ~A233;
  assign \new_[32108]_  = ~A232 & \new_[32107]_ ;
  assign \new_[32112]_  = ~A300 & A298;
  assign \new_[32113]_  = ~A266 & \new_[32112]_ ;
  assign \new_[32114]_  = \new_[32113]_  & \new_[32108]_ ;
  assign \new_[32118]_  = A167 & A169;
  assign \new_[32119]_  = ~A170 & \new_[32118]_ ;
  assign \new_[32123]_  = ~A201 & ~A200;
  assign \new_[32124]_  = A166 & \new_[32123]_ ;
  assign \new_[32125]_  = \new_[32124]_  & \new_[32119]_ ;
  assign \new_[32129]_  = ~A265 & ~A233;
  assign \new_[32130]_  = ~A232 & \new_[32129]_ ;
  assign \new_[32134]_  = A299 & A298;
  assign \new_[32135]_  = ~A266 & \new_[32134]_ ;
  assign \new_[32136]_  = \new_[32135]_  & \new_[32130]_ ;
  assign \new_[32140]_  = A167 & A169;
  assign \new_[32141]_  = ~A170 & \new_[32140]_ ;
  assign \new_[32145]_  = ~A201 & ~A200;
  assign \new_[32146]_  = A166 & \new_[32145]_ ;
  assign \new_[32147]_  = \new_[32146]_  & \new_[32141]_ ;
  assign \new_[32151]_  = ~A265 & ~A233;
  assign \new_[32152]_  = ~A232 & \new_[32151]_ ;
  assign \new_[32156]_  = ~A299 & ~A298;
  assign \new_[32157]_  = ~A266 & \new_[32156]_ ;
  assign \new_[32158]_  = \new_[32157]_  & \new_[32152]_ ;
  assign \new_[32162]_  = A167 & A169;
  assign \new_[32163]_  = ~A170 & \new_[32162]_ ;
  assign \new_[32167]_  = ~A200 & ~A199;
  assign \new_[32168]_  = A166 & \new_[32167]_ ;
  assign \new_[32169]_  = \new_[32168]_  & \new_[32163]_ ;
  assign \new_[32173]_  = A265 & A233;
  assign \new_[32174]_  = A232 & \new_[32173]_ ;
  assign \new_[32178]_  = ~A300 & ~A299;
  assign \new_[32179]_  = ~A267 & \new_[32178]_ ;
  assign \new_[32180]_  = \new_[32179]_  & \new_[32174]_ ;
  assign \new_[32184]_  = A167 & A169;
  assign \new_[32185]_  = ~A170 & \new_[32184]_ ;
  assign \new_[32189]_  = ~A200 & ~A199;
  assign \new_[32190]_  = A166 & \new_[32189]_ ;
  assign \new_[32191]_  = \new_[32190]_  & \new_[32185]_ ;
  assign \new_[32195]_  = A265 & A233;
  assign \new_[32196]_  = A232 & \new_[32195]_ ;
  assign \new_[32200]_  = A299 & A298;
  assign \new_[32201]_  = ~A267 & \new_[32200]_ ;
  assign \new_[32202]_  = \new_[32201]_  & \new_[32196]_ ;
  assign \new_[32206]_  = A167 & A169;
  assign \new_[32207]_  = ~A170 & \new_[32206]_ ;
  assign \new_[32211]_  = ~A200 & ~A199;
  assign \new_[32212]_  = A166 & \new_[32211]_ ;
  assign \new_[32213]_  = \new_[32212]_  & \new_[32207]_ ;
  assign \new_[32217]_  = A265 & A233;
  assign \new_[32218]_  = A232 & \new_[32217]_ ;
  assign \new_[32222]_  = ~A299 & ~A298;
  assign \new_[32223]_  = ~A267 & \new_[32222]_ ;
  assign \new_[32224]_  = \new_[32223]_  & \new_[32218]_ ;
  assign \new_[32228]_  = A167 & A169;
  assign \new_[32229]_  = ~A170 & \new_[32228]_ ;
  assign \new_[32233]_  = ~A200 & ~A199;
  assign \new_[32234]_  = A166 & \new_[32233]_ ;
  assign \new_[32235]_  = \new_[32234]_  & \new_[32229]_ ;
  assign \new_[32239]_  = A265 & A233;
  assign \new_[32240]_  = A232 & \new_[32239]_ ;
  assign \new_[32244]_  = ~A300 & ~A299;
  assign \new_[32245]_  = A266 & \new_[32244]_ ;
  assign \new_[32246]_  = \new_[32245]_  & \new_[32240]_ ;
  assign \new_[32250]_  = A167 & A169;
  assign \new_[32251]_  = ~A170 & \new_[32250]_ ;
  assign \new_[32255]_  = ~A200 & ~A199;
  assign \new_[32256]_  = A166 & \new_[32255]_ ;
  assign \new_[32257]_  = \new_[32256]_  & \new_[32251]_ ;
  assign \new_[32261]_  = A265 & A233;
  assign \new_[32262]_  = A232 & \new_[32261]_ ;
  assign \new_[32266]_  = A299 & A298;
  assign \new_[32267]_  = A266 & \new_[32266]_ ;
  assign \new_[32268]_  = \new_[32267]_  & \new_[32262]_ ;
  assign \new_[32272]_  = A167 & A169;
  assign \new_[32273]_  = ~A170 & \new_[32272]_ ;
  assign \new_[32277]_  = ~A200 & ~A199;
  assign \new_[32278]_  = A166 & \new_[32277]_ ;
  assign \new_[32279]_  = \new_[32278]_  & \new_[32273]_ ;
  assign \new_[32283]_  = A265 & A233;
  assign \new_[32284]_  = A232 & \new_[32283]_ ;
  assign \new_[32288]_  = ~A299 & ~A298;
  assign \new_[32289]_  = A266 & \new_[32288]_ ;
  assign \new_[32290]_  = \new_[32289]_  & \new_[32284]_ ;
  assign \new_[32294]_  = A167 & A169;
  assign \new_[32295]_  = ~A170 & \new_[32294]_ ;
  assign \new_[32299]_  = ~A200 & ~A199;
  assign \new_[32300]_  = A166 & \new_[32299]_ ;
  assign \new_[32301]_  = \new_[32300]_  & \new_[32295]_ ;
  assign \new_[32305]_  = ~A265 & A233;
  assign \new_[32306]_  = A232 & \new_[32305]_ ;
  assign \new_[32310]_  = ~A300 & ~A299;
  assign \new_[32311]_  = ~A266 & \new_[32310]_ ;
  assign \new_[32312]_  = \new_[32311]_  & \new_[32306]_ ;
  assign \new_[32316]_  = A167 & A169;
  assign \new_[32317]_  = ~A170 & \new_[32316]_ ;
  assign \new_[32321]_  = ~A200 & ~A199;
  assign \new_[32322]_  = A166 & \new_[32321]_ ;
  assign \new_[32323]_  = \new_[32322]_  & \new_[32317]_ ;
  assign \new_[32327]_  = ~A265 & A233;
  assign \new_[32328]_  = A232 & \new_[32327]_ ;
  assign \new_[32332]_  = A299 & A298;
  assign \new_[32333]_  = ~A266 & \new_[32332]_ ;
  assign \new_[32334]_  = \new_[32333]_  & \new_[32328]_ ;
  assign \new_[32338]_  = A167 & A169;
  assign \new_[32339]_  = ~A170 & \new_[32338]_ ;
  assign \new_[32343]_  = ~A200 & ~A199;
  assign \new_[32344]_  = A166 & \new_[32343]_ ;
  assign \new_[32345]_  = \new_[32344]_  & \new_[32339]_ ;
  assign \new_[32349]_  = ~A265 & A233;
  assign \new_[32350]_  = A232 & \new_[32349]_ ;
  assign \new_[32354]_  = ~A299 & ~A298;
  assign \new_[32355]_  = ~A266 & \new_[32354]_ ;
  assign \new_[32356]_  = \new_[32355]_  & \new_[32350]_ ;
  assign \new_[32360]_  = A167 & A169;
  assign \new_[32361]_  = ~A170 & \new_[32360]_ ;
  assign \new_[32365]_  = ~A200 & ~A199;
  assign \new_[32366]_  = A166 & \new_[32365]_ ;
  assign \new_[32367]_  = \new_[32366]_  & \new_[32361]_ ;
  assign \new_[32371]_  = A298 & A233;
  assign \new_[32372]_  = ~A232 & \new_[32371]_ ;
  assign \new_[32376]_  = A301 & A300;
  assign \new_[32377]_  = ~A299 & \new_[32376]_ ;
  assign \new_[32378]_  = \new_[32377]_  & \new_[32372]_ ;
  assign \new_[32382]_  = A167 & A169;
  assign \new_[32383]_  = ~A170 & \new_[32382]_ ;
  assign \new_[32387]_  = ~A200 & ~A199;
  assign \new_[32388]_  = A166 & \new_[32387]_ ;
  assign \new_[32389]_  = \new_[32388]_  & \new_[32383]_ ;
  assign \new_[32393]_  = A298 & A233;
  assign \new_[32394]_  = ~A232 & \new_[32393]_ ;
  assign \new_[32398]_  = A302 & A300;
  assign \new_[32399]_  = ~A299 & \new_[32398]_ ;
  assign \new_[32400]_  = \new_[32399]_  & \new_[32394]_ ;
  assign \new_[32404]_  = A167 & A169;
  assign \new_[32405]_  = ~A170 & \new_[32404]_ ;
  assign \new_[32409]_  = ~A200 & ~A199;
  assign \new_[32410]_  = A166 & \new_[32409]_ ;
  assign \new_[32411]_  = \new_[32410]_  & \new_[32405]_ ;
  assign \new_[32415]_  = A265 & A233;
  assign \new_[32416]_  = ~A232 & \new_[32415]_ ;
  assign \new_[32420]_  = A268 & A267;
  assign \new_[32421]_  = ~A266 & \new_[32420]_ ;
  assign \new_[32422]_  = \new_[32421]_  & \new_[32416]_ ;
  assign \new_[32426]_  = A167 & A169;
  assign \new_[32427]_  = ~A170 & \new_[32426]_ ;
  assign \new_[32431]_  = ~A200 & ~A199;
  assign \new_[32432]_  = A166 & \new_[32431]_ ;
  assign \new_[32433]_  = \new_[32432]_  & \new_[32427]_ ;
  assign \new_[32437]_  = A265 & A233;
  assign \new_[32438]_  = ~A232 & \new_[32437]_ ;
  assign \new_[32442]_  = A269 & A267;
  assign \new_[32443]_  = ~A266 & \new_[32442]_ ;
  assign \new_[32444]_  = \new_[32443]_  & \new_[32438]_ ;
  assign \new_[32448]_  = A167 & A169;
  assign \new_[32449]_  = ~A170 & \new_[32448]_ ;
  assign \new_[32453]_  = ~A200 & ~A199;
  assign \new_[32454]_  = A166 & \new_[32453]_ ;
  assign \new_[32455]_  = \new_[32454]_  & \new_[32449]_ ;
  assign \new_[32459]_  = A265 & ~A234;
  assign \new_[32460]_  = ~A233 & \new_[32459]_ ;
  assign \new_[32464]_  = ~A300 & A298;
  assign \new_[32465]_  = A266 & \new_[32464]_ ;
  assign \new_[32466]_  = \new_[32465]_  & \new_[32460]_ ;
  assign \new_[32470]_  = A167 & A169;
  assign \new_[32471]_  = ~A170 & \new_[32470]_ ;
  assign \new_[32475]_  = ~A200 & ~A199;
  assign \new_[32476]_  = A166 & \new_[32475]_ ;
  assign \new_[32477]_  = \new_[32476]_  & \new_[32471]_ ;
  assign \new_[32481]_  = A265 & ~A234;
  assign \new_[32482]_  = ~A233 & \new_[32481]_ ;
  assign \new_[32486]_  = A299 & A298;
  assign \new_[32487]_  = A266 & \new_[32486]_ ;
  assign \new_[32488]_  = \new_[32487]_  & \new_[32482]_ ;
  assign \new_[32492]_  = A167 & A169;
  assign \new_[32493]_  = ~A170 & \new_[32492]_ ;
  assign \new_[32497]_  = ~A200 & ~A199;
  assign \new_[32498]_  = A166 & \new_[32497]_ ;
  assign \new_[32499]_  = \new_[32498]_  & \new_[32493]_ ;
  assign \new_[32503]_  = A265 & ~A234;
  assign \new_[32504]_  = ~A233 & \new_[32503]_ ;
  assign \new_[32508]_  = ~A299 & ~A298;
  assign \new_[32509]_  = A266 & \new_[32508]_ ;
  assign \new_[32510]_  = \new_[32509]_  & \new_[32504]_ ;
  assign \new_[32514]_  = A167 & A169;
  assign \new_[32515]_  = ~A170 & \new_[32514]_ ;
  assign \new_[32519]_  = ~A200 & ~A199;
  assign \new_[32520]_  = A166 & \new_[32519]_ ;
  assign \new_[32521]_  = \new_[32520]_  & \new_[32515]_ ;
  assign \new_[32525]_  = ~A266 & ~A234;
  assign \new_[32526]_  = ~A233 & \new_[32525]_ ;
  assign \new_[32530]_  = ~A300 & A298;
  assign \new_[32531]_  = ~A267 & \new_[32530]_ ;
  assign \new_[32532]_  = \new_[32531]_  & \new_[32526]_ ;
  assign \new_[32536]_  = A167 & A169;
  assign \new_[32537]_  = ~A170 & \new_[32536]_ ;
  assign \new_[32541]_  = ~A200 & ~A199;
  assign \new_[32542]_  = A166 & \new_[32541]_ ;
  assign \new_[32543]_  = \new_[32542]_  & \new_[32537]_ ;
  assign \new_[32547]_  = ~A266 & ~A234;
  assign \new_[32548]_  = ~A233 & \new_[32547]_ ;
  assign \new_[32552]_  = A299 & A298;
  assign \new_[32553]_  = ~A267 & \new_[32552]_ ;
  assign \new_[32554]_  = \new_[32553]_  & \new_[32548]_ ;
  assign \new_[32558]_  = A167 & A169;
  assign \new_[32559]_  = ~A170 & \new_[32558]_ ;
  assign \new_[32563]_  = ~A200 & ~A199;
  assign \new_[32564]_  = A166 & \new_[32563]_ ;
  assign \new_[32565]_  = \new_[32564]_  & \new_[32559]_ ;
  assign \new_[32569]_  = ~A266 & ~A234;
  assign \new_[32570]_  = ~A233 & \new_[32569]_ ;
  assign \new_[32574]_  = ~A299 & ~A298;
  assign \new_[32575]_  = ~A267 & \new_[32574]_ ;
  assign \new_[32576]_  = \new_[32575]_  & \new_[32570]_ ;
  assign \new_[32580]_  = A167 & A169;
  assign \new_[32581]_  = ~A170 & \new_[32580]_ ;
  assign \new_[32585]_  = ~A200 & ~A199;
  assign \new_[32586]_  = A166 & \new_[32585]_ ;
  assign \new_[32587]_  = \new_[32586]_  & \new_[32581]_ ;
  assign \new_[32591]_  = ~A265 & ~A234;
  assign \new_[32592]_  = ~A233 & \new_[32591]_ ;
  assign \new_[32596]_  = ~A300 & A298;
  assign \new_[32597]_  = ~A266 & \new_[32596]_ ;
  assign \new_[32598]_  = \new_[32597]_  & \new_[32592]_ ;
  assign \new_[32602]_  = A167 & A169;
  assign \new_[32603]_  = ~A170 & \new_[32602]_ ;
  assign \new_[32607]_  = ~A200 & ~A199;
  assign \new_[32608]_  = A166 & \new_[32607]_ ;
  assign \new_[32609]_  = \new_[32608]_  & \new_[32603]_ ;
  assign \new_[32613]_  = ~A265 & ~A234;
  assign \new_[32614]_  = ~A233 & \new_[32613]_ ;
  assign \new_[32618]_  = A299 & A298;
  assign \new_[32619]_  = ~A266 & \new_[32618]_ ;
  assign \new_[32620]_  = \new_[32619]_  & \new_[32614]_ ;
  assign \new_[32624]_  = A167 & A169;
  assign \new_[32625]_  = ~A170 & \new_[32624]_ ;
  assign \new_[32629]_  = ~A200 & ~A199;
  assign \new_[32630]_  = A166 & \new_[32629]_ ;
  assign \new_[32631]_  = \new_[32630]_  & \new_[32625]_ ;
  assign \new_[32635]_  = ~A265 & ~A234;
  assign \new_[32636]_  = ~A233 & \new_[32635]_ ;
  assign \new_[32640]_  = ~A299 & ~A298;
  assign \new_[32641]_  = ~A266 & \new_[32640]_ ;
  assign \new_[32642]_  = \new_[32641]_  & \new_[32636]_ ;
  assign \new_[32646]_  = A167 & A169;
  assign \new_[32647]_  = ~A170 & \new_[32646]_ ;
  assign \new_[32651]_  = ~A200 & ~A199;
  assign \new_[32652]_  = A166 & \new_[32651]_ ;
  assign \new_[32653]_  = \new_[32652]_  & \new_[32647]_ ;
  assign \new_[32657]_  = A234 & ~A233;
  assign \new_[32658]_  = A232 & \new_[32657]_ ;
  assign \new_[32662]_  = A299 & ~A298;
  assign \new_[32663]_  = A235 & \new_[32662]_ ;
  assign \new_[32664]_  = \new_[32663]_  & \new_[32658]_ ;
  assign \new_[32668]_  = A167 & A169;
  assign \new_[32669]_  = ~A170 & \new_[32668]_ ;
  assign \new_[32673]_  = ~A200 & ~A199;
  assign \new_[32674]_  = A166 & \new_[32673]_ ;
  assign \new_[32675]_  = \new_[32674]_  & \new_[32669]_ ;
  assign \new_[32679]_  = A234 & ~A233;
  assign \new_[32680]_  = A232 & \new_[32679]_ ;
  assign \new_[32684]_  = A266 & ~A265;
  assign \new_[32685]_  = A235 & \new_[32684]_ ;
  assign \new_[32686]_  = \new_[32685]_  & \new_[32680]_ ;
  assign \new_[32690]_  = A167 & A169;
  assign \new_[32691]_  = ~A170 & \new_[32690]_ ;
  assign \new_[32695]_  = ~A200 & ~A199;
  assign \new_[32696]_  = A166 & \new_[32695]_ ;
  assign \new_[32697]_  = \new_[32696]_  & \new_[32691]_ ;
  assign \new_[32701]_  = A234 & ~A233;
  assign \new_[32702]_  = A232 & \new_[32701]_ ;
  assign \new_[32706]_  = A299 & ~A298;
  assign \new_[32707]_  = A236 & \new_[32706]_ ;
  assign \new_[32708]_  = \new_[32707]_  & \new_[32702]_ ;
  assign \new_[32712]_  = A167 & A169;
  assign \new_[32713]_  = ~A170 & \new_[32712]_ ;
  assign \new_[32717]_  = ~A200 & ~A199;
  assign \new_[32718]_  = A166 & \new_[32717]_ ;
  assign \new_[32719]_  = \new_[32718]_  & \new_[32713]_ ;
  assign \new_[32723]_  = A234 & ~A233;
  assign \new_[32724]_  = A232 & \new_[32723]_ ;
  assign \new_[32728]_  = A266 & ~A265;
  assign \new_[32729]_  = A236 & \new_[32728]_ ;
  assign \new_[32730]_  = \new_[32729]_  & \new_[32724]_ ;
  assign \new_[32734]_  = A167 & A169;
  assign \new_[32735]_  = ~A170 & \new_[32734]_ ;
  assign \new_[32739]_  = ~A200 & ~A199;
  assign \new_[32740]_  = A166 & \new_[32739]_ ;
  assign \new_[32741]_  = \new_[32740]_  & \new_[32735]_ ;
  assign \new_[32745]_  = A265 & ~A233;
  assign \new_[32746]_  = ~A232 & \new_[32745]_ ;
  assign \new_[32750]_  = ~A300 & A298;
  assign \new_[32751]_  = A266 & \new_[32750]_ ;
  assign \new_[32752]_  = \new_[32751]_  & \new_[32746]_ ;
  assign \new_[32756]_  = A167 & A169;
  assign \new_[32757]_  = ~A170 & \new_[32756]_ ;
  assign \new_[32761]_  = ~A200 & ~A199;
  assign \new_[32762]_  = A166 & \new_[32761]_ ;
  assign \new_[32763]_  = \new_[32762]_  & \new_[32757]_ ;
  assign \new_[32767]_  = A265 & ~A233;
  assign \new_[32768]_  = ~A232 & \new_[32767]_ ;
  assign \new_[32772]_  = A299 & A298;
  assign \new_[32773]_  = A266 & \new_[32772]_ ;
  assign \new_[32774]_  = \new_[32773]_  & \new_[32768]_ ;
  assign \new_[32778]_  = A167 & A169;
  assign \new_[32779]_  = ~A170 & \new_[32778]_ ;
  assign \new_[32783]_  = ~A200 & ~A199;
  assign \new_[32784]_  = A166 & \new_[32783]_ ;
  assign \new_[32785]_  = \new_[32784]_  & \new_[32779]_ ;
  assign \new_[32789]_  = A265 & ~A233;
  assign \new_[32790]_  = ~A232 & \new_[32789]_ ;
  assign \new_[32794]_  = ~A299 & ~A298;
  assign \new_[32795]_  = A266 & \new_[32794]_ ;
  assign \new_[32796]_  = \new_[32795]_  & \new_[32790]_ ;
  assign \new_[32800]_  = A167 & A169;
  assign \new_[32801]_  = ~A170 & \new_[32800]_ ;
  assign \new_[32805]_  = ~A200 & ~A199;
  assign \new_[32806]_  = A166 & \new_[32805]_ ;
  assign \new_[32807]_  = \new_[32806]_  & \new_[32801]_ ;
  assign \new_[32811]_  = ~A266 & ~A233;
  assign \new_[32812]_  = ~A232 & \new_[32811]_ ;
  assign \new_[32816]_  = ~A300 & A298;
  assign \new_[32817]_  = ~A267 & \new_[32816]_ ;
  assign \new_[32818]_  = \new_[32817]_  & \new_[32812]_ ;
  assign \new_[32822]_  = A167 & A169;
  assign \new_[32823]_  = ~A170 & \new_[32822]_ ;
  assign \new_[32827]_  = ~A200 & ~A199;
  assign \new_[32828]_  = A166 & \new_[32827]_ ;
  assign \new_[32829]_  = \new_[32828]_  & \new_[32823]_ ;
  assign \new_[32833]_  = ~A266 & ~A233;
  assign \new_[32834]_  = ~A232 & \new_[32833]_ ;
  assign \new_[32838]_  = A299 & A298;
  assign \new_[32839]_  = ~A267 & \new_[32838]_ ;
  assign \new_[32840]_  = \new_[32839]_  & \new_[32834]_ ;
  assign \new_[32844]_  = A167 & A169;
  assign \new_[32845]_  = ~A170 & \new_[32844]_ ;
  assign \new_[32849]_  = ~A200 & ~A199;
  assign \new_[32850]_  = A166 & \new_[32849]_ ;
  assign \new_[32851]_  = \new_[32850]_  & \new_[32845]_ ;
  assign \new_[32855]_  = ~A266 & ~A233;
  assign \new_[32856]_  = ~A232 & \new_[32855]_ ;
  assign \new_[32860]_  = ~A299 & ~A298;
  assign \new_[32861]_  = ~A267 & \new_[32860]_ ;
  assign \new_[32862]_  = \new_[32861]_  & \new_[32856]_ ;
  assign \new_[32866]_  = A167 & A169;
  assign \new_[32867]_  = ~A170 & \new_[32866]_ ;
  assign \new_[32871]_  = ~A200 & ~A199;
  assign \new_[32872]_  = A166 & \new_[32871]_ ;
  assign \new_[32873]_  = \new_[32872]_  & \new_[32867]_ ;
  assign \new_[32877]_  = ~A265 & ~A233;
  assign \new_[32878]_  = ~A232 & \new_[32877]_ ;
  assign \new_[32882]_  = ~A300 & A298;
  assign \new_[32883]_  = ~A266 & \new_[32882]_ ;
  assign \new_[32884]_  = \new_[32883]_  & \new_[32878]_ ;
  assign \new_[32888]_  = A167 & A169;
  assign \new_[32889]_  = ~A170 & \new_[32888]_ ;
  assign \new_[32893]_  = ~A200 & ~A199;
  assign \new_[32894]_  = A166 & \new_[32893]_ ;
  assign \new_[32895]_  = \new_[32894]_  & \new_[32889]_ ;
  assign \new_[32899]_  = ~A265 & ~A233;
  assign \new_[32900]_  = ~A232 & \new_[32899]_ ;
  assign \new_[32904]_  = A299 & A298;
  assign \new_[32905]_  = ~A266 & \new_[32904]_ ;
  assign \new_[32906]_  = \new_[32905]_  & \new_[32900]_ ;
  assign \new_[32910]_  = A167 & A169;
  assign \new_[32911]_  = ~A170 & \new_[32910]_ ;
  assign \new_[32915]_  = ~A200 & ~A199;
  assign \new_[32916]_  = A166 & \new_[32915]_ ;
  assign \new_[32917]_  = \new_[32916]_  & \new_[32911]_ ;
  assign \new_[32921]_  = ~A265 & ~A233;
  assign \new_[32922]_  = ~A232 & \new_[32921]_ ;
  assign \new_[32926]_  = ~A299 & ~A298;
  assign \new_[32927]_  = ~A266 & \new_[32926]_ ;
  assign \new_[32928]_  = \new_[32927]_  & \new_[32922]_ ;
  assign \new_[32932]_  = ~A167 & A169;
  assign \new_[32933]_  = ~A170 & \new_[32932]_ ;
  assign \new_[32937]_  = A200 & A199;
  assign \new_[32938]_  = ~A166 & \new_[32937]_ ;
  assign \new_[32939]_  = \new_[32938]_  & \new_[32933]_ ;
  assign \new_[32943]_  = A265 & A233;
  assign \new_[32944]_  = A232 & \new_[32943]_ ;
  assign \new_[32948]_  = ~A300 & ~A299;
  assign \new_[32949]_  = ~A267 & \new_[32948]_ ;
  assign \new_[32950]_  = \new_[32949]_  & \new_[32944]_ ;
  assign \new_[32954]_  = ~A167 & A169;
  assign \new_[32955]_  = ~A170 & \new_[32954]_ ;
  assign \new_[32959]_  = A200 & A199;
  assign \new_[32960]_  = ~A166 & \new_[32959]_ ;
  assign \new_[32961]_  = \new_[32960]_  & \new_[32955]_ ;
  assign \new_[32965]_  = A265 & A233;
  assign \new_[32966]_  = A232 & \new_[32965]_ ;
  assign \new_[32970]_  = A299 & A298;
  assign \new_[32971]_  = ~A267 & \new_[32970]_ ;
  assign \new_[32972]_  = \new_[32971]_  & \new_[32966]_ ;
  assign \new_[32976]_  = ~A167 & A169;
  assign \new_[32977]_  = ~A170 & \new_[32976]_ ;
  assign \new_[32981]_  = A200 & A199;
  assign \new_[32982]_  = ~A166 & \new_[32981]_ ;
  assign \new_[32983]_  = \new_[32982]_  & \new_[32977]_ ;
  assign \new_[32987]_  = A265 & A233;
  assign \new_[32988]_  = A232 & \new_[32987]_ ;
  assign \new_[32992]_  = ~A299 & ~A298;
  assign \new_[32993]_  = ~A267 & \new_[32992]_ ;
  assign \new_[32994]_  = \new_[32993]_  & \new_[32988]_ ;
  assign \new_[32998]_  = ~A167 & A169;
  assign \new_[32999]_  = ~A170 & \new_[32998]_ ;
  assign \new_[33003]_  = A200 & A199;
  assign \new_[33004]_  = ~A166 & \new_[33003]_ ;
  assign \new_[33005]_  = \new_[33004]_  & \new_[32999]_ ;
  assign \new_[33009]_  = A265 & A233;
  assign \new_[33010]_  = A232 & \new_[33009]_ ;
  assign \new_[33014]_  = ~A300 & ~A299;
  assign \new_[33015]_  = A266 & \new_[33014]_ ;
  assign \new_[33016]_  = \new_[33015]_  & \new_[33010]_ ;
  assign \new_[33020]_  = ~A167 & A169;
  assign \new_[33021]_  = ~A170 & \new_[33020]_ ;
  assign \new_[33025]_  = A200 & A199;
  assign \new_[33026]_  = ~A166 & \new_[33025]_ ;
  assign \new_[33027]_  = \new_[33026]_  & \new_[33021]_ ;
  assign \new_[33031]_  = A265 & A233;
  assign \new_[33032]_  = A232 & \new_[33031]_ ;
  assign \new_[33036]_  = A299 & A298;
  assign \new_[33037]_  = A266 & \new_[33036]_ ;
  assign \new_[33038]_  = \new_[33037]_  & \new_[33032]_ ;
  assign \new_[33042]_  = ~A167 & A169;
  assign \new_[33043]_  = ~A170 & \new_[33042]_ ;
  assign \new_[33047]_  = A200 & A199;
  assign \new_[33048]_  = ~A166 & \new_[33047]_ ;
  assign \new_[33049]_  = \new_[33048]_  & \new_[33043]_ ;
  assign \new_[33053]_  = A265 & A233;
  assign \new_[33054]_  = A232 & \new_[33053]_ ;
  assign \new_[33058]_  = ~A299 & ~A298;
  assign \new_[33059]_  = A266 & \new_[33058]_ ;
  assign \new_[33060]_  = \new_[33059]_  & \new_[33054]_ ;
  assign \new_[33064]_  = ~A167 & A169;
  assign \new_[33065]_  = ~A170 & \new_[33064]_ ;
  assign \new_[33069]_  = A200 & A199;
  assign \new_[33070]_  = ~A166 & \new_[33069]_ ;
  assign \new_[33071]_  = \new_[33070]_  & \new_[33065]_ ;
  assign \new_[33075]_  = ~A265 & A233;
  assign \new_[33076]_  = A232 & \new_[33075]_ ;
  assign \new_[33080]_  = ~A300 & ~A299;
  assign \new_[33081]_  = ~A266 & \new_[33080]_ ;
  assign \new_[33082]_  = \new_[33081]_  & \new_[33076]_ ;
  assign \new_[33086]_  = ~A167 & A169;
  assign \new_[33087]_  = ~A170 & \new_[33086]_ ;
  assign \new_[33091]_  = A200 & A199;
  assign \new_[33092]_  = ~A166 & \new_[33091]_ ;
  assign \new_[33093]_  = \new_[33092]_  & \new_[33087]_ ;
  assign \new_[33097]_  = ~A265 & A233;
  assign \new_[33098]_  = A232 & \new_[33097]_ ;
  assign \new_[33102]_  = A299 & A298;
  assign \new_[33103]_  = ~A266 & \new_[33102]_ ;
  assign \new_[33104]_  = \new_[33103]_  & \new_[33098]_ ;
  assign \new_[33108]_  = ~A167 & A169;
  assign \new_[33109]_  = ~A170 & \new_[33108]_ ;
  assign \new_[33113]_  = A200 & A199;
  assign \new_[33114]_  = ~A166 & \new_[33113]_ ;
  assign \new_[33115]_  = \new_[33114]_  & \new_[33109]_ ;
  assign \new_[33119]_  = ~A265 & A233;
  assign \new_[33120]_  = A232 & \new_[33119]_ ;
  assign \new_[33124]_  = ~A299 & ~A298;
  assign \new_[33125]_  = ~A266 & \new_[33124]_ ;
  assign \new_[33126]_  = \new_[33125]_  & \new_[33120]_ ;
  assign \new_[33130]_  = ~A167 & A169;
  assign \new_[33131]_  = ~A170 & \new_[33130]_ ;
  assign \new_[33135]_  = A200 & A199;
  assign \new_[33136]_  = ~A166 & \new_[33135]_ ;
  assign \new_[33137]_  = \new_[33136]_  & \new_[33131]_ ;
  assign \new_[33141]_  = A298 & A233;
  assign \new_[33142]_  = ~A232 & \new_[33141]_ ;
  assign \new_[33146]_  = A301 & A300;
  assign \new_[33147]_  = ~A299 & \new_[33146]_ ;
  assign \new_[33148]_  = \new_[33147]_  & \new_[33142]_ ;
  assign \new_[33152]_  = ~A167 & A169;
  assign \new_[33153]_  = ~A170 & \new_[33152]_ ;
  assign \new_[33157]_  = A200 & A199;
  assign \new_[33158]_  = ~A166 & \new_[33157]_ ;
  assign \new_[33159]_  = \new_[33158]_  & \new_[33153]_ ;
  assign \new_[33163]_  = A298 & A233;
  assign \new_[33164]_  = ~A232 & \new_[33163]_ ;
  assign \new_[33168]_  = A302 & A300;
  assign \new_[33169]_  = ~A299 & \new_[33168]_ ;
  assign \new_[33170]_  = \new_[33169]_  & \new_[33164]_ ;
  assign \new_[33174]_  = ~A167 & A169;
  assign \new_[33175]_  = ~A170 & \new_[33174]_ ;
  assign \new_[33179]_  = A200 & A199;
  assign \new_[33180]_  = ~A166 & \new_[33179]_ ;
  assign \new_[33181]_  = \new_[33180]_  & \new_[33175]_ ;
  assign \new_[33185]_  = A265 & A233;
  assign \new_[33186]_  = ~A232 & \new_[33185]_ ;
  assign \new_[33190]_  = A268 & A267;
  assign \new_[33191]_  = ~A266 & \new_[33190]_ ;
  assign \new_[33192]_  = \new_[33191]_  & \new_[33186]_ ;
  assign \new_[33196]_  = ~A167 & A169;
  assign \new_[33197]_  = ~A170 & \new_[33196]_ ;
  assign \new_[33201]_  = A200 & A199;
  assign \new_[33202]_  = ~A166 & \new_[33201]_ ;
  assign \new_[33203]_  = \new_[33202]_  & \new_[33197]_ ;
  assign \new_[33207]_  = A265 & A233;
  assign \new_[33208]_  = ~A232 & \new_[33207]_ ;
  assign \new_[33212]_  = A269 & A267;
  assign \new_[33213]_  = ~A266 & \new_[33212]_ ;
  assign \new_[33214]_  = \new_[33213]_  & \new_[33208]_ ;
  assign \new_[33218]_  = ~A167 & A169;
  assign \new_[33219]_  = ~A170 & \new_[33218]_ ;
  assign \new_[33223]_  = A200 & A199;
  assign \new_[33224]_  = ~A166 & \new_[33223]_ ;
  assign \new_[33225]_  = \new_[33224]_  & \new_[33219]_ ;
  assign \new_[33229]_  = A265 & ~A234;
  assign \new_[33230]_  = ~A233 & \new_[33229]_ ;
  assign \new_[33234]_  = ~A300 & A298;
  assign \new_[33235]_  = A266 & \new_[33234]_ ;
  assign \new_[33236]_  = \new_[33235]_  & \new_[33230]_ ;
  assign \new_[33240]_  = ~A167 & A169;
  assign \new_[33241]_  = ~A170 & \new_[33240]_ ;
  assign \new_[33245]_  = A200 & A199;
  assign \new_[33246]_  = ~A166 & \new_[33245]_ ;
  assign \new_[33247]_  = \new_[33246]_  & \new_[33241]_ ;
  assign \new_[33251]_  = A265 & ~A234;
  assign \new_[33252]_  = ~A233 & \new_[33251]_ ;
  assign \new_[33256]_  = A299 & A298;
  assign \new_[33257]_  = A266 & \new_[33256]_ ;
  assign \new_[33258]_  = \new_[33257]_  & \new_[33252]_ ;
  assign \new_[33262]_  = ~A167 & A169;
  assign \new_[33263]_  = ~A170 & \new_[33262]_ ;
  assign \new_[33267]_  = A200 & A199;
  assign \new_[33268]_  = ~A166 & \new_[33267]_ ;
  assign \new_[33269]_  = \new_[33268]_  & \new_[33263]_ ;
  assign \new_[33273]_  = A265 & ~A234;
  assign \new_[33274]_  = ~A233 & \new_[33273]_ ;
  assign \new_[33278]_  = ~A299 & ~A298;
  assign \new_[33279]_  = A266 & \new_[33278]_ ;
  assign \new_[33280]_  = \new_[33279]_  & \new_[33274]_ ;
  assign \new_[33284]_  = ~A167 & A169;
  assign \new_[33285]_  = ~A170 & \new_[33284]_ ;
  assign \new_[33289]_  = A200 & A199;
  assign \new_[33290]_  = ~A166 & \new_[33289]_ ;
  assign \new_[33291]_  = \new_[33290]_  & \new_[33285]_ ;
  assign \new_[33295]_  = ~A266 & ~A234;
  assign \new_[33296]_  = ~A233 & \new_[33295]_ ;
  assign \new_[33300]_  = ~A300 & A298;
  assign \new_[33301]_  = ~A267 & \new_[33300]_ ;
  assign \new_[33302]_  = \new_[33301]_  & \new_[33296]_ ;
  assign \new_[33306]_  = ~A167 & A169;
  assign \new_[33307]_  = ~A170 & \new_[33306]_ ;
  assign \new_[33311]_  = A200 & A199;
  assign \new_[33312]_  = ~A166 & \new_[33311]_ ;
  assign \new_[33313]_  = \new_[33312]_  & \new_[33307]_ ;
  assign \new_[33317]_  = ~A266 & ~A234;
  assign \new_[33318]_  = ~A233 & \new_[33317]_ ;
  assign \new_[33322]_  = A299 & A298;
  assign \new_[33323]_  = ~A267 & \new_[33322]_ ;
  assign \new_[33324]_  = \new_[33323]_  & \new_[33318]_ ;
  assign \new_[33328]_  = ~A167 & A169;
  assign \new_[33329]_  = ~A170 & \new_[33328]_ ;
  assign \new_[33333]_  = A200 & A199;
  assign \new_[33334]_  = ~A166 & \new_[33333]_ ;
  assign \new_[33335]_  = \new_[33334]_  & \new_[33329]_ ;
  assign \new_[33339]_  = ~A266 & ~A234;
  assign \new_[33340]_  = ~A233 & \new_[33339]_ ;
  assign \new_[33344]_  = ~A299 & ~A298;
  assign \new_[33345]_  = ~A267 & \new_[33344]_ ;
  assign \new_[33346]_  = \new_[33345]_  & \new_[33340]_ ;
  assign \new_[33350]_  = ~A167 & A169;
  assign \new_[33351]_  = ~A170 & \new_[33350]_ ;
  assign \new_[33355]_  = A200 & A199;
  assign \new_[33356]_  = ~A166 & \new_[33355]_ ;
  assign \new_[33357]_  = \new_[33356]_  & \new_[33351]_ ;
  assign \new_[33361]_  = ~A265 & ~A234;
  assign \new_[33362]_  = ~A233 & \new_[33361]_ ;
  assign \new_[33366]_  = ~A300 & A298;
  assign \new_[33367]_  = ~A266 & \new_[33366]_ ;
  assign \new_[33368]_  = \new_[33367]_  & \new_[33362]_ ;
  assign \new_[33372]_  = ~A167 & A169;
  assign \new_[33373]_  = ~A170 & \new_[33372]_ ;
  assign \new_[33377]_  = A200 & A199;
  assign \new_[33378]_  = ~A166 & \new_[33377]_ ;
  assign \new_[33379]_  = \new_[33378]_  & \new_[33373]_ ;
  assign \new_[33383]_  = ~A265 & ~A234;
  assign \new_[33384]_  = ~A233 & \new_[33383]_ ;
  assign \new_[33388]_  = A299 & A298;
  assign \new_[33389]_  = ~A266 & \new_[33388]_ ;
  assign \new_[33390]_  = \new_[33389]_  & \new_[33384]_ ;
  assign \new_[33394]_  = ~A167 & A169;
  assign \new_[33395]_  = ~A170 & \new_[33394]_ ;
  assign \new_[33399]_  = A200 & A199;
  assign \new_[33400]_  = ~A166 & \new_[33399]_ ;
  assign \new_[33401]_  = \new_[33400]_  & \new_[33395]_ ;
  assign \new_[33405]_  = ~A265 & ~A234;
  assign \new_[33406]_  = ~A233 & \new_[33405]_ ;
  assign \new_[33410]_  = ~A299 & ~A298;
  assign \new_[33411]_  = ~A266 & \new_[33410]_ ;
  assign \new_[33412]_  = \new_[33411]_  & \new_[33406]_ ;
  assign \new_[33416]_  = ~A167 & A169;
  assign \new_[33417]_  = ~A170 & \new_[33416]_ ;
  assign \new_[33421]_  = A200 & A199;
  assign \new_[33422]_  = ~A166 & \new_[33421]_ ;
  assign \new_[33423]_  = \new_[33422]_  & \new_[33417]_ ;
  assign \new_[33427]_  = A234 & ~A233;
  assign \new_[33428]_  = A232 & \new_[33427]_ ;
  assign \new_[33432]_  = A299 & ~A298;
  assign \new_[33433]_  = A235 & \new_[33432]_ ;
  assign \new_[33434]_  = \new_[33433]_  & \new_[33428]_ ;
  assign \new_[33438]_  = ~A167 & A169;
  assign \new_[33439]_  = ~A170 & \new_[33438]_ ;
  assign \new_[33443]_  = A200 & A199;
  assign \new_[33444]_  = ~A166 & \new_[33443]_ ;
  assign \new_[33445]_  = \new_[33444]_  & \new_[33439]_ ;
  assign \new_[33449]_  = A234 & ~A233;
  assign \new_[33450]_  = A232 & \new_[33449]_ ;
  assign \new_[33454]_  = A266 & ~A265;
  assign \new_[33455]_  = A235 & \new_[33454]_ ;
  assign \new_[33456]_  = \new_[33455]_  & \new_[33450]_ ;
  assign \new_[33460]_  = ~A167 & A169;
  assign \new_[33461]_  = ~A170 & \new_[33460]_ ;
  assign \new_[33465]_  = A200 & A199;
  assign \new_[33466]_  = ~A166 & \new_[33465]_ ;
  assign \new_[33467]_  = \new_[33466]_  & \new_[33461]_ ;
  assign \new_[33471]_  = A234 & ~A233;
  assign \new_[33472]_  = A232 & \new_[33471]_ ;
  assign \new_[33476]_  = A299 & ~A298;
  assign \new_[33477]_  = A236 & \new_[33476]_ ;
  assign \new_[33478]_  = \new_[33477]_  & \new_[33472]_ ;
  assign \new_[33482]_  = ~A167 & A169;
  assign \new_[33483]_  = ~A170 & \new_[33482]_ ;
  assign \new_[33487]_  = A200 & A199;
  assign \new_[33488]_  = ~A166 & \new_[33487]_ ;
  assign \new_[33489]_  = \new_[33488]_  & \new_[33483]_ ;
  assign \new_[33493]_  = A234 & ~A233;
  assign \new_[33494]_  = A232 & \new_[33493]_ ;
  assign \new_[33498]_  = A266 & ~A265;
  assign \new_[33499]_  = A236 & \new_[33498]_ ;
  assign \new_[33500]_  = \new_[33499]_  & \new_[33494]_ ;
  assign \new_[33504]_  = ~A167 & A169;
  assign \new_[33505]_  = ~A170 & \new_[33504]_ ;
  assign \new_[33509]_  = A200 & A199;
  assign \new_[33510]_  = ~A166 & \new_[33509]_ ;
  assign \new_[33511]_  = \new_[33510]_  & \new_[33505]_ ;
  assign \new_[33515]_  = A265 & ~A233;
  assign \new_[33516]_  = ~A232 & \new_[33515]_ ;
  assign \new_[33520]_  = ~A300 & A298;
  assign \new_[33521]_  = A266 & \new_[33520]_ ;
  assign \new_[33522]_  = \new_[33521]_  & \new_[33516]_ ;
  assign \new_[33526]_  = ~A167 & A169;
  assign \new_[33527]_  = ~A170 & \new_[33526]_ ;
  assign \new_[33531]_  = A200 & A199;
  assign \new_[33532]_  = ~A166 & \new_[33531]_ ;
  assign \new_[33533]_  = \new_[33532]_  & \new_[33527]_ ;
  assign \new_[33537]_  = A265 & ~A233;
  assign \new_[33538]_  = ~A232 & \new_[33537]_ ;
  assign \new_[33542]_  = A299 & A298;
  assign \new_[33543]_  = A266 & \new_[33542]_ ;
  assign \new_[33544]_  = \new_[33543]_  & \new_[33538]_ ;
  assign \new_[33548]_  = ~A167 & A169;
  assign \new_[33549]_  = ~A170 & \new_[33548]_ ;
  assign \new_[33553]_  = A200 & A199;
  assign \new_[33554]_  = ~A166 & \new_[33553]_ ;
  assign \new_[33555]_  = \new_[33554]_  & \new_[33549]_ ;
  assign \new_[33559]_  = A265 & ~A233;
  assign \new_[33560]_  = ~A232 & \new_[33559]_ ;
  assign \new_[33564]_  = ~A299 & ~A298;
  assign \new_[33565]_  = A266 & \new_[33564]_ ;
  assign \new_[33566]_  = \new_[33565]_  & \new_[33560]_ ;
  assign \new_[33570]_  = ~A167 & A169;
  assign \new_[33571]_  = ~A170 & \new_[33570]_ ;
  assign \new_[33575]_  = A200 & A199;
  assign \new_[33576]_  = ~A166 & \new_[33575]_ ;
  assign \new_[33577]_  = \new_[33576]_  & \new_[33571]_ ;
  assign \new_[33581]_  = ~A266 & ~A233;
  assign \new_[33582]_  = ~A232 & \new_[33581]_ ;
  assign \new_[33586]_  = ~A300 & A298;
  assign \new_[33587]_  = ~A267 & \new_[33586]_ ;
  assign \new_[33588]_  = \new_[33587]_  & \new_[33582]_ ;
  assign \new_[33592]_  = ~A167 & A169;
  assign \new_[33593]_  = ~A170 & \new_[33592]_ ;
  assign \new_[33597]_  = A200 & A199;
  assign \new_[33598]_  = ~A166 & \new_[33597]_ ;
  assign \new_[33599]_  = \new_[33598]_  & \new_[33593]_ ;
  assign \new_[33603]_  = ~A266 & ~A233;
  assign \new_[33604]_  = ~A232 & \new_[33603]_ ;
  assign \new_[33608]_  = A299 & A298;
  assign \new_[33609]_  = ~A267 & \new_[33608]_ ;
  assign \new_[33610]_  = \new_[33609]_  & \new_[33604]_ ;
  assign \new_[33614]_  = ~A167 & A169;
  assign \new_[33615]_  = ~A170 & \new_[33614]_ ;
  assign \new_[33619]_  = A200 & A199;
  assign \new_[33620]_  = ~A166 & \new_[33619]_ ;
  assign \new_[33621]_  = \new_[33620]_  & \new_[33615]_ ;
  assign \new_[33625]_  = ~A266 & ~A233;
  assign \new_[33626]_  = ~A232 & \new_[33625]_ ;
  assign \new_[33630]_  = ~A299 & ~A298;
  assign \new_[33631]_  = ~A267 & \new_[33630]_ ;
  assign \new_[33632]_  = \new_[33631]_  & \new_[33626]_ ;
  assign \new_[33636]_  = ~A167 & A169;
  assign \new_[33637]_  = ~A170 & \new_[33636]_ ;
  assign \new_[33641]_  = A200 & A199;
  assign \new_[33642]_  = ~A166 & \new_[33641]_ ;
  assign \new_[33643]_  = \new_[33642]_  & \new_[33637]_ ;
  assign \new_[33647]_  = ~A265 & ~A233;
  assign \new_[33648]_  = ~A232 & \new_[33647]_ ;
  assign \new_[33652]_  = ~A300 & A298;
  assign \new_[33653]_  = ~A266 & \new_[33652]_ ;
  assign \new_[33654]_  = \new_[33653]_  & \new_[33648]_ ;
  assign \new_[33658]_  = ~A167 & A169;
  assign \new_[33659]_  = ~A170 & \new_[33658]_ ;
  assign \new_[33663]_  = A200 & A199;
  assign \new_[33664]_  = ~A166 & \new_[33663]_ ;
  assign \new_[33665]_  = \new_[33664]_  & \new_[33659]_ ;
  assign \new_[33669]_  = ~A265 & ~A233;
  assign \new_[33670]_  = ~A232 & \new_[33669]_ ;
  assign \new_[33674]_  = A299 & A298;
  assign \new_[33675]_  = ~A266 & \new_[33674]_ ;
  assign \new_[33676]_  = \new_[33675]_  & \new_[33670]_ ;
  assign \new_[33680]_  = ~A167 & A169;
  assign \new_[33681]_  = ~A170 & \new_[33680]_ ;
  assign \new_[33685]_  = A200 & A199;
  assign \new_[33686]_  = ~A166 & \new_[33685]_ ;
  assign \new_[33687]_  = \new_[33686]_  & \new_[33681]_ ;
  assign \new_[33691]_  = ~A265 & ~A233;
  assign \new_[33692]_  = ~A232 & \new_[33691]_ ;
  assign \new_[33696]_  = ~A299 & ~A298;
  assign \new_[33697]_  = ~A266 & \new_[33696]_ ;
  assign \new_[33698]_  = \new_[33697]_  & \new_[33692]_ ;
  assign \new_[33702]_  = ~A167 & A169;
  assign \new_[33703]_  = ~A170 & \new_[33702]_ ;
  assign \new_[33707]_  = ~A201 & ~A200;
  assign \new_[33708]_  = ~A166 & \new_[33707]_ ;
  assign \new_[33709]_  = \new_[33708]_  & \new_[33703]_ ;
  assign \new_[33713]_  = A265 & A233;
  assign \new_[33714]_  = A232 & \new_[33713]_ ;
  assign \new_[33718]_  = ~A300 & ~A299;
  assign \new_[33719]_  = ~A267 & \new_[33718]_ ;
  assign \new_[33720]_  = \new_[33719]_  & \new_[33714]_ ;
  assign \new_[33724]_  = ~A167 & A169;
  assign \new_[33725]_  = ~A170 & \new_[33724]_ ;
  assign \new_[33729]_  = ~A201 & ~A200;
  assign \new_[33730]_  = ~A166 & \new_[33729]_ ;
  assign \new_[33731]_  = \new_[33730]_  & \new_[33725]_ ;
  assign \new_[33735]_  = A265 & A233;
  assign \new_[33736]_  = A232 & \new_[33735]_ ;
  assign \new_[33740]_  = A299 & A298;
  assign \new_[33741]_  = ~A267 & \new_[33740]_ ;
  assign \new_[33742]_  = \new_[33741]_  & \new_[33736]_ ;
  assign \new_[33746]_  = ~A167 & A169;
  assign \new_[33747]_  = ~A170 & \new_[33746]_ ;
  assign \new_[33751]_  = ~A201 & ~A200;
  assign \new_[33752]_  = ~A166 & \new_[33751]_ ;
  assign \new_[33753]_  = \new_[33752]_  & \new_[33747]_ ;
  assign \new_[33757]_  = A265 & A233;
  assign \new_[33758]_  = A232 & \new_[33757]_ ;
  assign \new_[33762]_  = ~A299 & ~A298;
  assign \new_[33763]_  = ~A267 & \new_[33762]_ ;
  assign \new_[33764]_  = \new_[33763]_  & \new_[33758]_ ;
  assign \new_[33768]_  = ~A167 & A169;
  assign \new_[33769]_  = ~A170 & \new_[33768]_ ;
  assign \new_[33773]_  = ~A201 & ~A200;
  assign \new_[33774]_  = ~A166 & \new_[33773]_ ;
  assign \new_[33775]_  = \new_[33774]_  & \new_[33769]_ ;
  assign \new_[33779]_  = A265 & A233;
  assign \new_[33780]_  = A232 & \new_[33779]_ ;
  assign \new_[33784]_  = ~A300 & ~A299;
  assign \new_[33785]_  = A266 & \new_[33784]_ ;
  assign \new_[33786]_  = \new_[33785]_  & \new_[33780]_ ;
  assign \new_[33790]_  = ~A167 & A169;
  assign \new_[33791]_  = ~A170 & \new_[33790]_ ;
  assign \new_[33795]_  = ~A201 & ~A200;
  assign \new_[33796]_  = ~A166 & \new_[33795]_ ;
  assign \new_[33797]_  = \new_[33796]_  & \new_[33791]_ ;
  assign \new_[33801]_  = A265 & A233;
  assign \new_[33802]_  = A232 & \new_[33801]_ ;
  assign \new_[33806]_  = A299 & A298;
  assign \new_[33807]_  = A266 & \new_[33806]_ ;
  assign \new_[33808]_  = \new_[33807]_  & \new_[33802]_ ;
  assign \new_[33812]_  = ~A167 & A169;
  assign \new_[33813]_  = ~A170 & \new_[33812]_ ;
  assign \new_[33817]_  = ~A201 & ~A200;
  assign \new_[33818]_  = ~A166 & \new_[33817]_ ;
  assign \new_[33819]_  = \new_[33818]_  & \new_[33813]_ ;
  assign \new_[33823]_  = A265 & A233;
  assign \new_[33824]_  = A232 & \new_[33823]_ ;
  assign \new_[33828]_  = ~A299 & ~A298;
  assign \new_[33829]_  = A266 & \new_[33828]_ ;
  assign \new_[33830]_  = \new_[33829]_  & \new_[33824]_ ;
  assign \new_[33834]_  = ~A167 & A169;
  assign \new_[33835]_  = ~A170 & \new_[33834]_ ;
  assign \new_[33839]_  = ~A201 & ~A200;
  assign \new_[33840]_  = ~A166 & \new_[33839]_ ;
  assign \new_[33841]_  = \new_[33840]_  & \new_[33835]_ ;
  assign \new_[33845]_  = ~A265 & A233;
  assign \new_[33846]_  = A232 & \new_[33845]_ ;
  assign \new_[33850]_  = ~A300 & ~A299;
  assign \new_[33851]_  = ~A266 & \new_[33850]_ ;
  assign \new_[33852]_  = \new_[33851]_  & \new_[33846]_ ;
  assign \new_[33856]_  = ~A167 & A169;
  assign \new_[33857]_  = ~A170 & \new_[33856]_ ;
  assign \new_[33861]_  = ~A201 & ~A200;
  assign \new_[33862]_  = ~A166 & \new_[33861]_ ;
  assign \new_[33863]_  = \new_[33862]_  & \new_[33857]_ ;
  assign \new_[33867]_  = ~A265 & A233;
  assign \new_[33868]_  = A232 & \new_[33867]_ ;
  assign \new_[33872]_  = A299 & A298;
  assign \new_[33873]_  = ~A266 & \new_[33872]_ ;
  assign \new_[33874]_  = \new_[33873]_  & \new_[33868]_ ;
  assign \new_[33878]_  = ~A167 & A169;
  assign \new_[33879]_  = ~A170 & \new_[33878]_ ;
  assign \new_[33883]_  = ~A201 & ~A200;
  assign \new_[33884]_  = ~A166 & \new_[33883]_ ;
  assign \new_[33885]_  = \new_[33884]_  & \new_[33879]_ ;
  assign \new_[33889]_  = ~A265 & A233;
  assign \new_[33890]_  = A232 & \new_[33889]_ ;
  assign \new_[33894]_  = ~A299 & ~A298;
  assign \new_[33895]_  = ~A266 & \new_[33894]_ ;
  assign \new_[33896]_  = \new_[33895]_  & \new_[33890]_ ;
  assign \new_[33900]_  = ~A167 & A169;
  assign \new_[33901]_  = ~A170 & \new_[33900]_ ;
  assign \new_[33905]_  = ~A201 & ~A200;
  assign \new_[33906]_  = ~A166 & \new_[33905]_ ;
  assign \new_[33907]_  = \new_[33906]_  & \new_[33901]_ ;
  assign \new_[33911]_  = A298 & A233;
  assign \new_[33912]_  = ~A232 & \new_[33911]_ ;
  assign \new_[33916]_  = A301 & A300;
  assign \new_[33917]_  = ~A299 & \new_[33916]_ ;
  assign \new_[33918]_  = \new_[33917]_  & \new_[33912]_ ;
  assign \new_[33922]_  = ~A167 & A169;
  assign \new_[33923]_  = ~A170 & \new_[33922]_ ;
  assign \new_[33927]_  = ~A201 & ~A200;
  assign \new_[33928]_  = ~A166 & \new_[33927]_ ;
  assign \new_[33929]_  = \new_[33928]_  & \new_[33923]_ ;
  assign \new_[33933]_  = A298 & A233;
  assign \new_[33934]_  = ~A232 & \new_[33933]_ ;
  assign \new_[33938]_  = A302 & A300;
  assign \new_[33939]_  = ~A299 & \new_[33938]_ ;
  assign \new_[33940]_  = \new_[33939]_  & \new_[33934]_ ;
  assign \new_[33944]_  = ~A167 & A169;
  assign \new_[33945]_  = ~A170 & \new_[33944]_ ;
  assign \new_[33949]_  = ~A201 & ~A200;
  assign \new_[33950]_  = ~A166 & \new_[33949]_ ;
  assign \new_[33951]_  = \new_[33950]_  & \new_[33945]_ ;
  assign \new_[33955]_  = A265 & A233;
  assign \new_[33956]_  = ~A232 & \new_[33955]_ ;
  assign \new_[33960]_  = A268 & A267;
  assign \new_[33961]_  = ~A266 & \new_[33960]_ ;
  assign \new_[33962]_  = \new_[33961]_  & \new_[33956]_ ;
  assign \new_[33966]_  = ~A167 & A169;
  assign \new_[33967]_  = ~A170 & \new_[33966]_ ;
  assign \new_[33971]_  = ~A201 & ~A200;
  assign \new_[33972]_  = ~A166 & \new_[33971]_ ;
  assign \new_[33973]_  = \new_[33972]_  & \new_[33967]_ ;
  assign \new_[33977]_  = A265 & A233;
  assign \new_[33978]_  = ~A232 & \new_[33977]_ ;
  assign \new_[33982]_  = A269 & A267;
  assign \new_[33983]_  = ~A266 & \new_[33982]_ ;
  assign \new_[33984]_  = \new_[33983]_  & \new_[33978]_ ;
  assign \new_[33988]_  = ~A167 & A169;
  assign \new_[33989]_  = ~A170 & \new_[33988]_ ;
  assign \new_[33993]_  = ~A201 & ~A200;
  assign \new_[33994]_  = ~A166 & \new_[33993]_ ;
  assign \new_[33995]_  = \new_[33994]_  & \new_[33989]_ ;
  assign \new_[33999]_  = A265 & ~A234;
  assign \new_[34000]_  = ~A233 & \new_[33999]_ ;
  assign \new_[34004]_  = ~A300 & A298;
  assign \new_[34005]_  = A266 & \new_[34004]_ ;
  assign \new_[34006]_  = \new_[34005]_  & \new_[34000]_ ;
  assign \new_[34010]_  = ~A167 & A169;
  assign \new_[34011]_  = ~A170 & \new_[34010]_ ;
  assign \new_[34015]_  = ~A201 & ~A200;
  assign \new_[34016]_  = ~A166 & \new_[34015]_ ;
  assign \new_[34017]_  = \new_[34016]_  & \new_[34011]_ ;
  assign \new_[34021]_  = A265 & ~A234;
  assign \new_[34022]_  = ~A233 & \new_[34021]_ ;
  assign \new_[34026]_  = A299 & A298;
  assign \new_[34027]_  = A266 & \new_[34026]_ ;
  assign \new_[34028]_  = \new_[34027]_  & \new_[34022]_ ;
  assign \new_[34032]_  = ~A167 & A169;
  assign \new_[34033]_  = ~A170 & \new_[34032]_ ;
  assign \new_[34037]_  = ~A201 & ~A200;
  assign \new_[34038]_  = ~A166 & \new_[34037]_ ;
  assign \new_[34039]_  = \new_[34038]_  & \new_[34033]_ ;
  assign \new_[34043]_  = A265 & ~A234;
  assign \new_[34044]_  = ~A233 & \new_[34043]_ ;
  assign \new_[34048]_  = ~A299 & ~A298;
  assign \new_[34049]_  = A266 & \new_[34048]_ ;
  assign \new_[34050]_  = \new_[34049]_  & \new_[34044]_ ;
  assign \new_[34054]_  = ~A167 & A169;
  assign \new_[34055]_  = ~A170 & \new_[34054]_ ;
  assign \new_[34059]_  = ~A201 & ~A200;
  assign \new_[34060]_  = ~A166 & \new_[34059]_ ;
  assign \new_[34061]_  = \new_[34060]_  & \new_[34055]_ ;
  assign \new_[34065]_  = ~A266 & ~A234;
  assign \new_[34066]_  = ~A233 & \new_[34065]_ ;
  assign \new_[34070]_  = ~A300 & A298;
  assign \new_[34071]_  = ~A267 & \new_[34070]_ ;
  assign \new_[34072]_  = \new_[34071]_  & \new_[34066]_ ;
  assign \new_[34076]_  = ~A167 & A169;
  assign \new_[34077]_  = ~A170 & \new_[34076]_ ;
  assign \new_[34081]_  = ~A201 & ~A200;
  assign \new_[34082]_  = ~A166 & \new_[34081]_ ;
  assign \new_[34083]_  = \new_[34082]_  & \new_[34077]_ ;
  assign \new_[34087]_  = ~A266 & ~A234;
  assign \new_[34088]_  = ~A233 & \new_[34087]_ ;
  assign \new_[34092]_  = A299 & A298;
  assign \new_[34093]_  = ~A267 & \new_[34092]_ ;
  assign \new_[34094]_  = \new_[34093]_  & \new_[34088]_ ;
  assign \new_[34098]_  = ~A167 & A169;
  assign \new_[34099]_  = ~A170 & \new_[34098]_ ;
  assign \new_[34103]_  = ~A201 & ~A200;
  assign \new_[34104]_  = ~A166 & \new_[34103]_ ;
  assign \new_[34105]_  = \new_[34104]_  & \new_[34099]_ ;
  assign \new_[34109]_  = ~A266 & ~A234;
  assign \new_[34110]_  = ~A233 & \new_[34109]_ ;
  assign \new_[34114]_  = ~A299 & ~A298;
  assign \new_[34115]_  = ~A267 & \new_[34114]_ ;
  assign \new_[34116]_  = \new_[34115]_  & \new_[34110]_ ;
  assign \new_[34120]_  = ~A167 & A169;
  assign \new_[34121]_  = ~A170 & \new_[34120]_ ;
  assign \new_[34125]_  = ~A201 & ~A200;
  assign \new_[34126]_  = ~A166 & \new_[34125]_ ;
  assign \new_[34127]_  = \new_[34126]_  & \new_[34121]_ ;
  assign \new_[34131]_  = ~A265 & ~A234;
  assign \new_[34132]_  = ~A233 & \new_[34131]_ ;
  assign \new_[34136]_  = ~A300 & A298;
  assign \new_[34137]_  = ~A266 & \new_[34136]_ ;
  assign \new_[34138]_  = \new_[34137]_  & \new_[34132]_ ;
  assign \new_[34142]_  = ~A167 & A169;
  assign \new_[34143]_  = ~A170 & \new_[34142]_ ;
  assign \new_[34147]_  = ~A201 & ~A200;
  assign \new_[34148]_  = ~A166 & \new_[34147]_ ;
  assign \new_[34149]_  = \new_[34148]_  & \new_[34143]_ ;
  assign \new_[34153]_  = ~A265 & ~A234;
  assign \new_[34154]_  = ~A233 & \new_[34153]_ ;
  assign \new_[34158]_  = A299 & A298;
  assign \new_[34159]_  = ~A266 & \new_[34158]_ ;
  assign \new_[34160]_  = \new_[34159]_  & \new_[34154]_ ;
  assign \new_[34164]_  = ~A167 & A169;
  assign \new_[34165]_  = ~A170 & \new_[34164]_ ;
  assign \new_[34169]_  = ~A201 & ~A200;
  assign \new_[34170]_  = ~A166 & \new_[34169]_ ;
  assign \new_[34171]_  = \new_[34170]_  & \new_[34165]_ ;
  assign \new_[34175]_  = ~A265 & ~A234;
  assign \new_[34176]_  = ~A233 & \new_[34175]_ ;
  assign \new_[34180]_  = ~A299 & ~A298;
  assign \new_[34181]_  = ~A266 & \new_[34180]_ ;
  assign \new_[34182]_  = \new_[34181]_  & \new_[34176]_ ;
  assign \new_[34186]_  = ~A167 & A169;
  assign \new_[34187]_  = ~A170 & \new_[34186]_ ;
  assign \new_[34191]_  = ~A201 & ~A200;
  assign \new_[34192]_  = ~A166 & \new_[34191]_ ;
  assign \new_[34193]_  = \new_[34192]_  & \new_[34187]_ ;
  assign \new_[34197]_  = A234 & ~A233;
  assign \new_[34198]_  = A232 & \new_[34197]_ ;
  assign \new_[34202]_  = A299 & ~A298;
  assign \new_[34203]_  = A235 & \new_[34202]_ ;
  assign \new_[34204]_  = \new_[34203]_  & \new_[34198]_ ;
  assign \new_[34208]_  = ~A167 & A169;
  assign \new_[34209]_  = ~A170 & \new_[34208]_ ;
  assign \new_[34213]_  = ~A201 & ~A200;
  assign \new_[34214]_  = ~A166 & \new_[34213]_ ;
  assign \new_[34215]_  = \new_[34214]_  & \new_[34209]_ ;
  assign \new_[34219]_  = A234 & ~A233;
  assign \new_[34220]_  = A232 & \new_[34219]_ ;
  assign \new_[34224]_  = A266 & ~A265;
  assign \new_[34225]_  = A235 & \new_[34224]_ ;
  assign \new_[34226]_  = \new_[34225]_  & \new_[34220]_ ;
  assign \new_[34230]_  = ~A167 & A169;
  assign \new_[34231]_  = ~A170 & \new_[34230]_ ;
  assign \new_[34235]_  = ~A201 & ~A200;
  assign \new_[34236]_  = ~A166 & \new_[34235]_ ;
  assign \new_[34237]_  = \new_[34236]_  & \new_[34231]_ ;
  assign \new_[34241]_  = A234 & ~A233;
  assign \new_[34242]_  = A232 & \new_[34241]_ ;
  assign \new_[34246]_  = A299 & ~A298;
  assign \new_[34247]_  = A236 & \new_[34246]_ ;
  assign \new_[34248]_  = \new_[34247]_  & \new_[34242]_ ;
  assign \new_[34252]_  = ~A167 & A169;
  assign \new_[34253]_  = ~A170 & \new_[34252]_ ;
  assign \new_[34257]_  = ~A201 & ~A200;
  assign \new_[34258]_  = ~A166 & \new_[34257]_ ;
  assign \new_[34259]_  = \new_[34258]_  & \new_[34253]_ ;
  assign \new_[34263]_  = A234 & ~A233;
  assign \new_[34264]_  = A232 & \new_[34263]_ ;
  assign \new_[34268]_  = A266 & ~A265;
  assign \new_[34269]_  = A236 & \new_[34268]_ ;
  assign \new_[34270]_  = \new_[34269]_  & \new_[34264]_ ;
  assign \new_[34274]_  = ~A167 & A169;
  assign \new_[34275]_  = ~A170 & \new_[34274]_ ;
  assign \new_[34279]_  = ~A201 & ~A200;
  assign \new_[34280]_  = ~A166 & \new_[34279]_ ;
  assign \new_[34281]_  = \new_[34280]_  & \new_[34275]_ ;
  assign \new_[34285]_  = A265 & ~A233;
  assign \new_[34286]_  = ~A232 & \new_[34285]_ ;
  assign \new_[34290]_  = ~A300 & A298;
  assign \new_[34291]_  = A266 & \new_[34290]_ ;
  assign \new_[34292]_  = \new_[34291]_  & \new_[34286]_ ;
  assign \new_[34296]_  = ~A167 & A169;
  assign \new_[34297]_  = ~A170 & \new_[34296]_ ;
  assign \new_[34301]_  = ~A201 & ~A200;
  assign \new_[34302]_  = ~A166 & \new_[34301]_ ;
  assign \new_[34303]_  = \new_[34302]_  & \new_[34297]_ ;
  assign \new_[34307]_  = A265 & ~A233;
  assign \new_[34308]_  = ~A232 & \new_[34307]_ ;
  assign \new_[34312]_  = A299 & A298;
  assign \new_[34313]_  = A266 & \new_[34312]_ ;
  assign \new_[34314]_  = \new_[34313]_  & \new_[34308]_ ;
  assign \new_[34318]_  = ~A167 & A169;
  assign \new_[34319]_  = ~A170 & \new_[34318]_ ;
  assign \new_[34323]_  = ~A201 & ~A200;
  assign \new_[34324]_  = ~A166 & \new_[34323]_ ;
  assign \new_[34325]_  = \new_[34324]_  & \new_[34319]_ ;
  assign \new_[34329]_  = A265 & ~A233;
  assign \new_[34330]_  = ~A232 & \new_[34329]_ ;
  assign \new_[34334]_  = ~A299 & ~A298;
  assign \new_[34335]_  = A266 & \new_[34334]_ ;
  assign \new_[34336]_  = \new_[34335]_  & \new_[34330]_ ;
  assign \new_[34340]_  = ~A167 & A169;
  assign \new_[34341]_  = ~A170 & \new_[34340]_ ;
  assign \new_[34345]_  = ~A201 & ~A200;
  assign \new_[34346]_  = ~A166 & \new_[34345]_ ;
  assign \new_[34347]_  = \new_[34346]_  & \new_[34341]_ ;
  assign \new_[34351]_  = ~A266 & ~A233;
  assign \new_[34352]_  = ~A232 & \new_[34351]_ ;
  assign \new_[34356]_  = ~A300 & A298;
  assign \new_[34357]_  = ~A267 & \new_[34356]_ ;
  assign \new_[34358]_  = \new_[34357]_  & \new_[34352]_ ;
  assign \new_[34362]_  = ~A167 & A169;
  assign \new_[34363]_  = ~A170 & \new_[34362]_ ;
  assign \new_[34367]_  = ~A201 & ~A200;
  assign \new_[34368]_  = ~A166 & \new_[34367]_ ;
  assign \new_[34369]_  = \new_[34368]_  & \new_[34363]_ ;
  assign \new_[34373]_  = ~A266 & ~A233;
  assign \new_[34374]_  = ~A232 & \new_[34373]_ ;
  assign \new_[34378]_  = A299 & A298;
  assign \new_[34379]_  = ~A267 & \new_[34378]_ ;
  assign \new_[34380]_  = \new_[34379]_  & \new_[34374]_ ;
  assign \new_[34384]_  = ~A167 & A169;
  assign \new_[34385]_  = ~A170 & \new_[34384]_ ;
  assign \new_[34389]_  = ~A201 & ~A200;
  assign \new_[34390]_  = ~A166 & \new_[34389]_ ;
  assign \new_[34391]_  = \new_[34390]_  & \new_[34385]_ ;
  assign \new_[34395]_  = ~A266 & ~A233;
  assign \new_[34396]_  = ~A232 & \new_[34395]_ ;
  assign \new_[34400]_  = ~A299 & ~A298;
  assign \new_[34401]_  = ~A267 & \new_[34400]_ ;
  assign \new_[34402]_  = \new_[34401]_  & \new_[34396]_ ;
  assign \new_[34406]_  = ~A167 & A169;
  assign \new_[34407]_  = ~A170 & \new_[34406]_ ;
  assign \new_[34411]_  = ~A201 & ~A200;
  assign \new_[34412]_  = ~A166 & \new_[34411]_ ;
  assign \new_[34413]_  = \new_[34412]_  & \new_[34407]_ ;
  assign \new_[34417]_  = ~A265 & ~A233;
  assign \new_[34418]_  = ~A232 & \new_[34417]_ ;
  assign \new_[34422]_  = ~A300 & A298;
  assign \new_[34423]_  = ~A266 & \new_[34422]_ ;
  assign \new_[34424]_  = \new_[34423]_  & \new_[34418]_ ;
  assign \new_[34428]_  = ~A167 & A169;
  assign \new_[34429]_  = ~A170 & \new_[34428]_ ;
  assign \new_[34433]_  = ~A201 & ~A200;
  assign \new_[34434]_  = ~A166 & \new_[34433]_ ;
  assign \new_[34435]_  = \new_[34434]_  & \new_[34429]_ ;
  assign \new_[34439]_  = ~A265 & ~A233;
  assign \new_[34440]_  = ~A232 & \new_[34439]_ ;
  assign \new_[34444]_  = A299 & A298;
  assign \new_[34445]_  = ~A266 & \new_[34444]_ ;
  assign \new_[34446]_  = \new_[34445]_  & \new_[34440]_ ;
  assign \new_[34450]_  = ~A167 & A169;
  assign \new_[34451]_  = ~A170 & \new_[34450]_ ;
  assign \new_[34455]_  = ~A201 & ~A200;
  assign \new_[34456]_  = ~A166 & \new_[34455]_ ;
  assign \new_[34457]_  = \new_[34456]_  & \new_[34451]_ ;
  assign \new_[34461]_  = ~A265 & ~A233;
  assign \new_[34462]_  = ~A232 & \new_[34461]_ ;
  assign \new_[34466]_  = ~A299 & ~A298;
  assign \new_[34467]_  = ~A266 & \new_[34466]_ ;
  assign \new_[34468]_  = \new_[34467]_  & \new_[34462]_ ;
  assign \new_[34472]_  = ~A167 & A169;
  assign \new_[34473]_  = ~A170 & \new_[34472]_ ;
  assign \new_[34477]_  = ~A200 & ~A199;
  assign \new_[34478]_  = ~A166 & \new_[34477]_ ;
  assign \new_[34479]_  = \new_[34478]_  & \new_[34473]_ ;
  assign \new_[34483]_  = A265 & A233;
  assign \new_[34484]_  = A232 & \new_[34483]_ ;
  assign \new_[34488]_  = ~A300 & ~A299;
  assign \new_[34489]_  = ~A267 & \new_[34488]_ ;
  assign \new_[34490]_  = \new_[34489]_  & \new_[34484]_ ;
  assign \new_[34494]_  = ~A167 & A169;
  assign \new_[34495]_  = ~A170 & \new_[34494]_ ;
  assign \new_[34499]_  = ~A200 & ~A199;
  assign \new_[34500]_  = ~A166 & \new_[34499]_ ;
  assign \new_[34501]_  = \new_[34500]_  & \new_[34495]_ ;
  assign \new_[34505]_  = A265 & A233;
  assign \new_[34506]_  = A232 & \new_[34505]_ ;
  assign \new_[34510]_  = A299 & A298;
  assign \new_[34511]_  = ~A267 & \new_[34510]_ ;
  assign \new_[34512]_  = \new_[34511]_  & \new_[34506]_ ;
  assign \new_[34516]_  = ~A167 & A169;
  assign \new_[34517]_  = ~A170 & \new_[34516]_ ;
  assign \new_[34521]_  = ~A200 & ~A199;
  assign \new_[34522]_  = ~A166 & \new_[34521]_ ;
  assign \new_[34523]_  = \new_[34522]_  & \new_[34517]_ ;
  assign \new_[34527]_  = A265 & A233;
  assign \new_[34528]_  = A232 & \new_[34527]_ ;
  assign \new_[34532]_  = ~A299 & ~A298;
  assign \new_[34533]_  = ~A267 & \new_[34532]_ ;
  assign \new_[34534]_  = \new_[34533]_  & \new_[34528]_ ;
  assign \new_[34538]_  = ~A167 & A169;
  assign \new_[34539]_  = ~A170 & \new_[34538]_ ;
  assign \new_[34543]_  = ~A200 & ~A199;
  assign \new_[34544]_  = ~A166 & \new_[34543]_ ;
  assign \new_[34545]_  = \new_[34544]_  & \new_[34539]_ ;
  assign \new_[34549]_  = A265 & A233;
  assign \new_[34550]_  = A232 & \new_[34549]_ ;
  assign \new_[34554]_  = ~A300 & ~A299;
  assign \new_[34555]_  = A266 & \new_[34554]_ ;
  assign \new_[34556]_  = \new_[34555]_  & \new_[34550]_ ;
  assign \new_[34560]_  = ~A167 & A169;
  assign \new_[34561]_  = ~A170 & \new_[34560]_ ;
  assign \new_[34565]_  = ~A200 & ~A199;
  assign \new_[34566]_  = ~A166 & \new_[34565]_ ;
  assign \new_[34567]_  = \new_[34566]_  & \new_[34561]_ ;
  assign \new_[34571]_  = A265 & A233;
  assign \new_[34572]_  = A232 & \new_[34571]_ ;
  assign \new_[34576]_  = A299 & A298;
  assign \new_[34577]_  = A266 & \new_[34576]_ ;
  assign \new_[34578]_  = \new_[34577]_  & \new_[34572]_ ;
  assign \new_[34582]_  = ~A167 & A169;
  assign \new_[34583]_  = ~A170 & \new_[34582]_ ;
  assign \new_[34587]_  = ~A200 & ~A199;
  assign \new_[34588]_  = ~A166 & \new_[34587]_ ;
  assign \new_[34589]_  = \new_[34588]_  & \new_[34583]_ ;
  assign \new_[34593]_  = A265 & A233;
  assign \new_[34594]_  = A232 & \new_[34593]_ ;
  assign \new_[34598]_  = ~A299 & ~A298;
  assign \new_[34599]_  = A266 & \new_[34598]_ ;
  assign \new_[34600]_  = \new_[34599]_  & \new_[34594]_ ;
  assign \new_[34604]_  = ~A167 & A169;
  assign \new_[34605]_  = ~A170 & \new_[34604]_ ;
  assign \new_[34609]_  = ~A200 & ~A199;
  assign \new_[34610]_  = ~A166 & \new_[34609]_ ;
  assign \new_[34611]_  = \new_[34610]_  & \new_[34605]_ ;
  assign \new_[34615]_  = ~A265 & A233;
  assign \new_[34616]_  = A232 & \new_[34615]_ ;
  assign \new_[34620]_  = ~A300 & ~A299;
  assign \new_[34621]_  = ~A266 & \new_[34620]_ ;
  assign \new_[34622]_  = \new_[34621]_  & \new_[34616]_ ;
  assign \new_[34626]_  = ~A167 & A169;
  assign \new_[34627]_  = ~A170 & \new_[34626]_ ;
  assign \new_[34631]_  = ~A200 & ~A199;
  assign \new_[34632]_  = ~A166 & \new_[34631]_ ;
  assign \new_[34633]_  = \new_[34632]_  & \new_[34627]_ ;
  assign \new_[34637]_  = ~A265 & A233;
  assign \new_[34638]_  = A232 & \new_[34637]_ ;
  assign \new_[34642]_  = A299 & A298;
  assign \new_[34643]_  = ~A266 & \new_[34642]_ ;
  assign \new_[34644]_  = \new_[34643]_  & \new_[34638]_ ;
  assign \new_[34648]_  = ~A167 & A169;
  assign \new_[34649]_  = ~A170 & \new_[34648]_ ;
  assign \new_[34653]_  = ~A200 & ~A199;
  assign \new_[34654]_  = ~A166 & \new_[34653]_ ;
  assign \new_[34655]_  = \new_[34654]_  & \new_[34649]_ ;
  assign \new_[34659]_  = ~A265 & A233;
  assign \new_[34660]_  = A232 & \new_[34659]_ ;
  assign \new_[34664]_  = ~A299 & ~A298;
  assign \new_[34665]_  = ~A266 & \new_[34664]_ ;
  assign \new_[34666]_  = \new_[34665]_  & \new_[34660]_ ;
  assign \new_[34670]_  = ~A167 & A169;
  assign \new_[34671]_  = ~A170 & \new_[34670]_ ;
  assign \new_[34675]_  = ~A200 & ~A199;
  assign \new_[34676]_  = ~A166 & \new_[34675]_ ;
  assign \new_[34677]_  = \new_[34676]_  & \new_[34671]_ ;
  assign \new_[34681]_  = A298 & A233;
  assign \new_[34682]_  = ~A232 & \new_[34681]_ ;
  assign \new_[34686]_  = A301 & A300;
  assign \new_[34687]_  = ~A299 & \new_[34686]_ ;
  assign \new_[34688]_  = \new_[34687]_  & \new_[34682]_ ;
  assign \new_[34692]_  = ~A167 & A169;
  assign \new_[34693]_  = ~A170 & \new_[34692]_ ;
  assign \new_[34697]_  = ~A200 & ~A199;
  assign \new_[34698]_  = ~A166 & \new_[34697]_ ;
  assign \new_[34699]_  = \new_[34698]_  & \new_[34693]_ ;
  assign \new_[34703]_  = A298 & A233;
  assign \new_[34704]_  = ~A232 & \new_[34703]_ ;
  assign \new_[34708]_  = A302 & A300;
  assign \new_[34709]_  = ~A299 & \new_[34708]_ ;
  assign \new_[34710]_  = \new_[34709]_  & \new_[34704]_ ;
  assign \new_[34714]_  = ~A167 & A169;
  assign \new_[34715]_  = ~A170 & \new_[34714]_ ;
  assign \new_[34719]_  = ~A200 & ~A199;
  assign \new_[34720]_  = ~A166 & \new_[34719]_ ;
  assign \new_[34721]_  = \new_[34720]_  & \new_[34715]_ ;
  assign \new_[34725]_  = A265 & A233;
  assign \new_[34726]_  = ~A232 & \new_[34725]_ ;
  assign \new_[34730]_  = A268 & A267;
  assign \new_[34731]_  = ~A266 & \new_[34730]_ ;
  assign \new_[34732]_  = \new_[34731]_  & \new_[34726]_ ;
  assign \new_[34736]_  = ~A167 & A169;
  assign \new_[34737]_  = ~A170 & \new_[34736]_ ;
  assign \new_[34741]_  = ~A200 & ~A199;
  assign \new_[34742]_  = ~A166 & \new_[34741]_ ;
  assign \new_[34743]_  = \new_[34742]_  & \new_[34737]_ ;
  assign \new_[34747]_  = A265 & A233;
  assign \new_[34748]_  = ~A232 & \new_[34747]_ ;
  assign \new_[34752]_  = A269 & A267;
  assign \new_[34753]_  = ~A266 & \new_[34752]_ ;
  assign \new_[34754]_  = \new_[34753]_  & \new_[34748]_ ;
  assign \new_[34758]_  = ~A167 & A169;
  assign \new_[34759]_  = ~A170 & \new_[34758]_ ;
  assign \new_[34763]_  = ~A200 & ~A199;
  assign \new_[34764]_  = ~A166 & \new_[34763]_ ;
  assign \new_[34765]_  = \new_[34764]_  & \new_[34759]_ ;
  assign \new_[34769]_  = A265 & ~A234;
  assign \new_[34770]_  = ~A233 & \new_[34769]_ ;
  assign \new_[34774]_  = ~A300 & A298;
  assign \new_[34775]_  = A266 & \new_[34774]_ ;
  assign \new_[34776]_  = \new_[34775]_  & \new_[34770]_ ;
  assign \new_[34780]_  = ~A167 & A169;
  assign \new_[34781]_  = ~A170 & \new_[34780]_ ;
  assign \new_[34785]_  = ~A200 & ~A199;
  assign \new_[34786]_  = ~A166 & \new_[34785]_ ;
  assign \new_[34787]_  = \new_[34786]_  & \new_[34781]_ ;
  assign \new_[34791]_  = A265 & ~A234;
  assign \new_[34792]_  = ~A233 & \new_[34791]_ ;
  assign \new_[34796]_  = A299 & A298;
  assign \new_[34797]_  = A266 & \new_[34796]_ ;
  assign \new_[34798]_  = \new_[34797]_  & \new_[34792]_ ;
  assign \new_[34802]_  = ~A167 & A169;
  assign \new_[34803]_  = ~A170 & \new_[34802]_ ;
  assign \new_[34807]_  = ~A200 & ~A199;
  assign \new_[34808]_  = ~A166 & \new_[34807]_ ;
  assign \new_[34809]_  = \new_[34808]_  & \new_[34803]_ ;
  assign \new_[34813]_  = A265 & ~A234;
  assign \new_[34814]_  = ~A233 & \new_[34813]_ ;
  assign \new_[34818]_  = ~A299 & ~A298;
  assign \new_[34819]_  = A266 & \new_[34818]_ ;
  assign \new_[34820]_  = \new_[34819]_  & \new_[34814]_ ;
  assign \new_[34824]_  = ~A167 & A169;
  assign \new_[34825]_  = ~A170 & \new_[34824]_ ;
  assign \new_[34829]_  = ~A200 & ~A199;
  assign \new_[34830]_  = ~A166 & \new_[34829]_ ;
  assign \new_[34831]_  = \new_[34830]_  & \new_[34825]_ ;
  assign \new_[34835]_  = ~A266 & ~A234;
  assign \new_[34836]_  = ~A233 & \new_[34835]_ ;
  assign \new_[34840]_  = ~A300 & A298;
  assign \new_[34841]_  = ~A267 & \new_[34840]_ ;
  assign \new_[34842]_  = \new_[34841]_  & \new_[34836]_ ;
  assign \new_[34846]_  = ~A167 & A169;
  assign \new_[34847]_  = ~A170 & \new_[34846]_ ;
  assign \new_[34851]_  = ~A200 & ~A199;
  assign \new_[34852]_  = ~A166 & \new_[34851]_ ;
  assign \new_[34853]_  = \new_[34852]_  & \new_[34847]_ ;
  assign \new_[34857]_  = ~A266 & ~A234;
  assign \new_[34858]_  = ~A233 & \new_[34857]_ ;
  assign \new_[34862]_  = A299 & A298;
  assign \new_[34863]_  = ~A267 & \new_[34862]_ ;
  assign \new_[34864]_  = \new_[34863]_  & \new_[34858]_ ;
  assign \new_[34868]_  = ~A167 & A169;
  assign \new_[34869]_  = ~A170 & \new_[34868]_ ;
  assign \new_[34873]_  = ~A200 & ~A199;
  assign \new_[34874]_  = ~A166 & \new_[34873]_ ;
  assign \new_[34875]_  = \new_[34874]_  & \new_[34869]_ ;
  assign \new_[34879]_  = ~A266 & ~A234;
  assign \new_[34880]_  = ~A233 & \new_[34879]_ ;
  assign \new_[34884]_  = ~A299 & ~A298;
  assign \new_[34885]_  = ~A267 & \new_[34884]_ ;
  assign \new_[34886]_  = \new_[34885]_  & \new_[34880]_ ;
  assign \new_[34890]_  = ~A167 & A169;
  assign \new_[34891]_  = ~A170 & \new_[34890]_ ;
  assign \new_[34895]_  = ~A200 & ~A199;
  assign \new_[34896]_  = ~A166 & \new_[34895]_ ;
  assign \new_[34897]_  = \new_[34896]_  & \new_[34891]_ ;
  assign \new_[34901]_  = ~A265 & ~A234;
  assign \new_[34902]_  = ~A233 & \new_[34901]_ ;
  assign \new_[34906]_  = ~A300 & A298;
  assign \new_[34907]_  = ~A266 & \new_[34906]_ ;
  assign \new_[34908]_  = \new_[34907]_  & \new_[34902]_ ;
  assign \new_[34912]_  = ~A167 & A169;
  assign \new_[34913]_  = ~A170 & \new_[34912]_ ;
  assign \new_[34917]_  = ~A200 & ~A199;
  assign \new_[34918]_  = ~A166 & \new_[34917]_ ;
  assign \new_[34919]_  = \new_[34918]_  & \new_[34913]_ ;
  assign \new_[34923]_  = ~A265 & ~A234;
  assign \new_[34924]_  = ~A233 & \new_[34923]_ ;
  assign \new_[34928]_  = A299 & A298;
  assign \new_[34929]_  = ~A266 & \new_[34928]_ ;
  assign \new_[34930]_  = \new_[34929]_  & \new_[34924]_ ;
  assign \new_[34934]_  = ~A167 & A169;
  assign \new_[34935]_  = ~A170 & \new_[34934]_ ;
  assign \new_[34939]_  = ~A200 & ~A199;
  assign \new_[34940]_  = ~A166 & \new_[34939]_ ;
  assign \new_[34941]_  = \new_[34940]_  & \new_[34935]_ ;
  assign \new_[34945]_  = ~A265 & ~A234;
  assign \new_[34946]_  = ~A233 & \new_[34945]_ ;
  assign \new_[34950]_  = ~A299 & ~A298;
  assign \new_[34951]_  = ~A266 & \new_[34950]_ ;
  assign \new_[34952]_  = \new_[34951]_  & \new_[34946]_ ;
  assign \new_[34956]_  = ~A167 & A169;
  assign \new_[34957]_  = ~A170 & \new_[34956]_ ;
  assign \new_[34961]_  = ~A200 & ~A199;
  assign \new_[34962]_  = ~A166 & \new_[34961]_ ;
  assign \new_[34963]_  = \new_[34962]_  & \new_[34957]_ ;
  assign \new_[34967]_  = A234 & ~A233;
  assign \new_[34968]_  = A232 & \new_[34967]_ ;
  assign \new_[34972]_  = A299 & ~A298;
  assign \new_[34973]_  = A235 & \new_[34972]_ ;
  assign \new_[34974]_  = \new_[34973]_  & \new_[34968]_ ;
  assign \new_[34978]_  = ~A167 & A169;
  assign \new_[34979]_  = ~A170 & \new_[34978]_ ;
  assign \new_[34983]_  = ~A200 & ~A199;
  assign \new_[34984]_  = ~A166 & \new_[34983]_ ;
  assign \new_[34985]_  = \new_[34984]_  & \new_[34979]_ ;
  assign \new_[34989]_  = A234 & ~A233;
  assign \new_[34990]_  = A232 & \new_[34989]_ ;
  assign \new_[34994]_  = A266 & ~A265;
  assign \new_[34995]_  = A235 & \new_[34994]_ ;
  assign \new_[34996]_  = \new_[34995]_  & \new_[34990]_ ;
  assign \new_[35000]_  = ~A167 & A169;
  assign \new_[35001]_  = ~A170 & \new_[35000]_ ;
  assign \new_[35005]_  = ~A200 & ~A199;
  assign \new_[35006]_  = ~A166 & \new_[35005]_ ;
  assign \new_[35007]_  = \new_[35006]_  & \new_[35001]_ ;
  assign \new_[35011]_  = A234 & ~A233;
  assign \new_[35012]_  = A232 & \new_[35011]_ ;
  assign \new_[35016]_  = A299 & ~A298;
  assign \new_[35017]_  = A236 & \new_[35016]_ ;
  assign \new_[35018]_  = \new_[35017]_  & \new_[35012]_ ;
  assign \new_[35022]_  = ~A167 & A169;
  assign \new_[35023]_  = ~A170 & \new_[35022]_ ;
  assign \new_[35027]_  = ~A200 & ~A199;
  assign \new_[35028]_  = ~A166 & \new_[35027]_ ;
  assign \new_[35029]_  = \new_[35028]_  & \new_[35023]_ ;
  assign \new_[35033]_  = A234 & ~A233;
  assign \new_[35034]_  = A232 & \new_[35033]_ ;
  assign \new_[35038]_  = A266 & ~A265;
  assign \new_[35039]_  = A236 & \new_[35038]_ ;
  assign \new_[35040]_  = \new_[35039]_  & \new_[35034]_ ;
  assign \new_[35044]_  = ~A167 & A169;
  assign \new_[35045]_  = ~A170 & \new_[35044]_ ;
  assign \new_[35049]_  = ~A200 & ~A199;
  assign \new_[35050]_  = ~A166 & \new_[35049]_ ;
  assign \new_[35051]_  = \new_[35050]_  & \new_[35045]_ ;
  assign \new_[35055]_  = A265 & ~A233;
  assign \new_[35056]_  = ~A232 & \new_[35055]_ ;
  assign \new_[35060]_  = ~A300 & A298;
  assign \new_[35061]_  = A266 & \new_[35060]_ ;
  assign \new_[35062]_  = \new_[35061]_  & \new_[35056]_ ;
  assign \new_[35066]_  = ~A167 & A169;
  assign \new_[35067]_  = ~A170 & \new_[35066]_ ;
  assign \new_[35071]_  = ~A200 & ~A199;
  assign \new_[35072]_  = ~A166 & \new_[35071]_ ;
  assign \new_[35073]_  = \new_[35072]_  & \new_[35067]_ ;
  assign \new_[35077]_  = A265 & ~A233;
  assign \new_[35078]_  = ~A232 & \new_[35077]_ ;
  assign \new_[35082]_  = A299 & A298;
  assign \new_[35083]_  = A266 & \new_[35082]_ ;
  assign \new_[35084]_  = \new_[35083]_  & \new_[35078]_ ;
  assign \new_[35088]_  = ~A167 & A169;
  assign \new_[35089]_  = ~A170 & \new_[35088]_ ;
  assign \new_[35093]_  = ~A200 & ~A199;
  assign \new_[35094]_  = ~A166 & \new_[35093]_ ;
  assign \new_[35095]_  = \new_[35094]_  & \new_[35089]_ ;
  assign \new_[35099]_  = A265 & ~A233;
  assign \new_[35100]_  = ~A232 & \new_[35099]_ ;
  assign \new_[35104]_  = ~A299 & ~A298;
  assign \new_[35105]_  = A266 & \new_[35104]_ ;
  assign \new_[35106]_  = \new_[35105]_  & \new_[35100]_ ;
  assign \new_[35110]_  = ~A167 & A169;
  assign \new_[35111]_  = ~A170 & \new_[35110]_ ;
  assign \new_[35115]_  = ~A200 & ~A199;
  assign \new_[35116]_  = ~A166 & \new_[35115]_ ;
  assign \new_[35117]_  = \new_[35116]_  & \new_[35111]_ ;
  assign \new_[35121]_  = ~A266 & ~A233;
  assign \new_[35122]_  = ~A232 & \new_[35121]_ ;
  assign \new_[35126]_  = ~A300 & A298;
  assign \new_[35127]_  = ~A267 & \new_[35126]_ ;
  assign \new_[35128]_  = \new_[35127]_  & \new_[35122]_ ;
  assign \new_[35132]_  = ~A167 & A169;
  assign \new_[35133]_  = ~A170 & \new_[35132]_ ;
  assign \new_[35137]_  = ~A200 & ~A199;
  assign \new_[35138]_  = ~A166 & \new_[35137]_ ;
  assign \new_[35139]_  = \new_[35138]_  & \new_[35133]_ ;
  assign \new_[35143]_  = ~A266 & ~A233;
  assign \new_[35144]_  = ~A232 & \new_[35143]_ ;
  assign \new_[35148]_  = A299 & A298;
  assign \new_[35149]_  = ~A267 & \new_[35148]_ ;
  assign \new_[35150]_  = \new_[35149]_  & \new_[35144]_ ;
  assign \new_[35154]_  = ~A167 & A169;
  assign \new_[35155]_  = ~A170 & \new_[35154]_ ;
  assign \new_[35159]_  = ~A200 & ~A199;
  assign \new_[35160]_  = ~A166 & \new_[35159]_ ;
  assign \new_[35161]_  = \new_[35160]_  & \new_[35155]_ ;
  assign \new_[35165]_  = ~A266 & ~A233;
  assign \new_[35166]_  = ~A232 & \new_[35165]_ ;
  assign \new_[35170]_  = ~A299 & ~A298;
  assign \new_[35171]_  = ~A267 & \new_[35170]_ ;
  assign \new_[35172]_  = \new_[35171]_  & \new_[35166]_ ;
  assign \new_[35176]_  = ~A167 & A169;
  assign \new_[35177]_  = ~A170 & \new_[35176]_ ;
  assign \new_[35181]_  = ~A200 & ~A199;
  assign \new_[35182]_  = ~A166 & \new_[35181]_ ;
  assign \new_[35183]_  = \new_[35182]_  & \new_[35177]_ ;
  assign \new_[35187]_  = ~A265 & ~A233;
  assign \new_[35188]_  = ~A232 & \new_[35187]_ ;
  assign \new_[35192]_  = ~A300 & A298;
  assign \new_[35193]_  = ~A266 & \new_[35192]_ ;
  assign \new_[35194]_  = \new_[35193]_  & \new_[35188]_ ;
  assign \new_[35198]_  = ~A167 & A169;
  assign \new_[35199]_  = ~A170 & \new_[35198]_ ;
  assign \new_[35203]_  = ~A200 & ~A199;
  assign \new_[35204]_  = ~A166 & \new_[35203]_ ;
  assign \new_[35205]_  = \new_[35204]_  & \new_[35199]_ ;
  assign \new_[35209]_  = ~A265 & ~A233;
  assign \new_[35210]_  = ~A232 & \new_[35209]_ ;
  assign \new_[35214]_  = A299 & A298;
  assign \new_[35215]_  = ~A266 & \new_[35214]_ ;
  assign \new_[35216]_  = \new_[35215]_  & \new_[35210]_ ;
  assign \new_[35220]_  = ~A167 & A169;
  assign \new_[35221]_  = ~A170 & \new_[35220]_ ;
  assign \new_[35225]_  = ~A200 & ~A199;
  assign \new_[35226]_  = ~A166 & \new_[35225]_ ;
  assign \new_[35227]_  = \new_[35226]_  & \new_[35221]_ ;
  assign \new_[35231]_  = ~A265 & ~A233;
  assign \new_[35232]_  = ~A232 & \new_[35231]_ ;
  assign \new_[35236]_  = ~A299 & ~A298;
  assign \new_[35237]_  = ~A266 & \new_[35236]_ ;
  assign \new_[35238]_  = \new_[35237]_  & \new_[35232]_ ;
  assign \new_[35242]_  = ~A166 & ~A167;
  assign \new_[35243]_  = ~A169 & \new_[35242]_ ;
  assign \new_[35247]_  = A232 & A200;
  assign \new_[35248]_  = ~A199 & \new_[35247]_ ;
  assign \new_[35249]_  = \new_[35248]_  & \new_[35243]_ ;
  assign \new_[35253]_  = ~A268 & A265;
  assign \new_[35254]_  = A233 & \new_[35253]_ ;
  assign \new_[35258]_  = ~A300 & ~A299;
  assign \new_[35259]_  = ~A269 & \new_[35258]_ ;
  assign \new_[35260]_  = \new_[35259]_  & \new_[35254]_ ;
  assign \new_[35264]_  = ~A166 & ~A167;
  assign \new_[35265]_  = ~A169 & \new_[35264]_ ;
  assign \new_[35269]_  = A232 & A200;
  assign \new_[35270]_  = ~A199 & \new_[35269]_ ;
  assign \new_[35271]_  = \new_[35270]_  & \new_[35265]_ ;
  assign \new_[35275]_  = ~A268 & A265;
  assign \new_[35276]_  = A233 & \new_[35275]_ ;
  assign \new_[35280]_  = A299 & A298;
  assign \new_[35281]_  = ~A269 & \new_[35280]_ ;
  assign \new_[35282]_  = \new_[35281]_  & \new_[35276]_ ;
  assign \new_[35286]_  = ~A166 & ~A167;
  assign \new_[35287]_  = ~A169 & \new_[35286]_ ;
  assign \new_[35291]_  = A232 & A200;
  assign \new_[35292]_  = ~A199 & \new_[35291]_ ;
  assign \new_[35293]_  = \new_[35292]_  & \new_[35287]_ ;
  assign \new_[35297]_  = ~A268 & A265;
  assign \new_[35298]_  = A233 & \new_[35297]_ ;
  assign \new_[35302]_  = ~A299 & ~A298;
  assign \new_[35303]_  = ~A269 & \new_[35302]_ ;
  assign \new_[35304]_  = \new_[35303]_  & \new_[35298]_ ;
  assign \new_[35308]_  = ~A166 & ~A167;
  assign \new_[35309]_  = ~A169 & \new_[35308]_ ;
  assign \new_[35313]_  = A232 & A200;
  assign \new_[35314]_  = ~A199 & \new_[35313]_ ;
  assign \new_[35315]_  = \new_[35314]_  & \new_[35309]_ ;
  assign \new_[35319]_  = ~A267 & A265;
  assign \new_[35320]_  = A233 & \new_[35319]_ ;
  assign \new_[35324]_  = ~A302 & ~A301;
  assign \new_[35325]_  = ~A299 & \new_[35324]_ ;
  assign \new_[35326]_  = \new_[35325]_  & \new_[35320]_ ;
  assign \new_[35330]_  = ~A166 & ~A167;
  assign \new_[35331]_  = ~A169 & \new_[35330]_ ;
  assign \new_[35335]_  = A232 & A200;
  assign \new_[35336]_  = ~A199 & \new_[35335]_ ;
  assign \new_[35337]_  = \new_[35336]_  & \new_[35331]_ ;
  assign \new_[35341]_  = A266 & A265;
  assign \new_[35342]_  = A233 & \new_[35341]_ ;
  assign \new_[35346]_  = ~A302 & ~A301;
  assign \new_[35347]_  = ~A299 & \new_[35346]_ ;
  assign \new_[35348]_  = \new_[35347]_  & \new_[35342]_ ;
  assign \new_[35352]_  = ~A166 & ~A167;
  assign \new_[35353]_  = ~A169 & \new_[35352]_ ;
  assign \new_[35357]_  = A232 & A200;
  assign \new_[35358]_  = ~A199 & \new_[35357]_ ;
  assign \new_[35359]_  = \new_[35358]_  & \new_[35353]_ ;
  assign \new_[35363]_  = ~A266 & ~A265;
  assign \new_[35364]_  = A233 & \new_[35363]_ ;
  assign \new_[35368]_  = ~A302 & ~A301;
  assign \new_[35369]_  = ~A299 & \new_[35368]_ ;
  assign \new_[35370]_  = \new_[35369]_  & \new_[35364]_ ;
  assign \new_[35374]_  = ~A166 & ~A167;
  assign \new_[35375]_  = ~A169 & \new_[35374]_ ;
  assign \new_[35379]_  = ~A233 & A200;
  assign \new_[35380]_  = ~A199 & \new_[35379]_ ;
  assign \new_[35381]_  = \new_[35380]_  & \new_[35375]_ ;
  assign \new_[35385]_  = A265 & ~A236;
  assign \new_[35386]_  = ~A235 & \new_[35385]_ ;
  assign \new_[35390]_  = ~A300 & A298;
  assign \new_[35391]_  = A266 & \new_[35390]_ ;
  assign \new_[35392]_  = \new_[35391]_  & \new_[35386]_ ;
  assign \new_[35396]_  = ~A166 & ~A167;
  assign \new_[35397]_  = ~A169 & \new_[35396]_ ;
  assign \new_[35401]_  = ~A233 & A200;
  assign \new_[35402]_  = ~A199 & \new_[35401]_ ;
  assign \new_[35403]_  = \new_[35402]_  & \new_[35397]_ ;
  assign \new_[35407]_  = A265 & ~A236;
  assign \new_[35408]_  = ~A235 & \new_[35407]_ ;
  assign \new_[35412]_  = A299 & A298;
  assign \new_[35413]_  = A266 & \new_[35412]_ ;
  assign \new_[35414]_  = \new_[35413]_  & \new_[35408]_ ;
  assign \new_[35418]_  = ~A166 & ~A167;
  assign \new_[35419]_  = ~A169 & \new_[35418]_ ;
  assign \new_[35423]_  = ~A233 & A200;
  assign \new_[35424]_  = ~A199 & \new_[35423]_ ;
  assign \new_[35425]_  = \new_[35424]_  & \new_[35419]_ ;
  assign \new_[35429]_  = A265 & ~A236;
  assign \new_[35430]_  = ~A235 & \new_[35429]_ ;
  assign \new_[35434]_  = ~A299 & ~A298;
  assign \new_[35435]_  = A266 & \new_[35434]_ ;
  assign \new_[35436]_  = \new_[35435]_  & \new_[35430]_ ;
  assign \new_[35440]_  = ~A166 & ~A167;
  assign \new_[35441]_  = ~A169 & \new_[35440]_ ;
  assign \new_[35445]_  = ~A233 & A200;
  assign \new_[35446]_  = ~A199 & \new_[35445]_ ;
  assign \new_[35447]_  = \new_[35446]_  & \new_[35441]_ ;
  assign \new_[35451]_  = ~A266 & ~A236;
  assign \new_[35452]_  = ~A235 & \new_[35451]_ ;
  assign \new_[35456]_  = ~A300 & A298;
  assign \new_[35457]_  = ~A267 & \new_[35456]_ ;
  assign \new_[35458]_  = \new_[35457]_  & \new_[35452]_ ;
  assign \new_[35462]_  = ~A166 & ~A167;
  assign \new_[35463]_  = ~A169 & \new_[35462]_ ;
  assign \new_[35467]_  = ~A233 & A200;
  assign \new_[35468]_  = ~A199 & \new_[35467]_ ;
  assign \new_[35469]_  = \new_[35468]_  & \new_[35463]_ ;
  assign \new_[35473]_  = ~A266 & ~A236;
  assign \new_[35474]_  = ~A235 & \new_[35473]_ ;
  assign \new_[35478]_  = A299 & A298;
  assign \new_[35479]_  = ~A267 & \new_[35478]_ ;
  assign \new_[35480]_  = \new_[35479]_  & \new_[35474]_ ;
  assign \new_[35484]_  = ~A166 & ~A167;
  assign \new_[35485]_  = ~A169 & \new_[35484]_ ;
  assign \new_[35489]_  = ~A233 & A200;
  assign \new_[35490]_  = ~A199 & \new_[35489]_ ;
  assign \new_[35491]_  = \new_[35490]_  & \new_[35485]_ ;
  assign \new_[35495]_  = ~A266 & ~A236;
  assign \new_[35496]_  = ~A235 & \new_[35495]_ ;
  assign \new_[35500]_  = ~A299 & ~A298;
  assign \new_[35501]_  = ~A267 & \new_[35500]_ ;
  assign \new_[35502]_  = \new_[35501]_  & \new_[35496]_ ;
  assign \new_[35506]_  = ~A166 & ~A167;
  assign \new_[35507]_  = ~A169 & \new_[35506]_ ;
  assign \new_[35511]_  = ~A233 & A200;
  assign \new_[35512]_  = ~A199 & \new_[35511]_ ;
  assign \new_[35513]_  = \new_[35512]_  & \new_[35507]_ ;
  assign \new_[35517]_  = ~A265 & ~A236;
  assign \new_[35518]_  = ~A235 & \new_[35517]_ ;
  assign \new_[35522]_  = ~A300 & A298;
  assign \new_[35523]_  = ~A266 & \new_[35522]_ ;
  assign \new_[35524]_  = \new_[35523]_  & \new_[35518]_ ;
  assign \new_[35528]_  = ~A166 & ~A167;
  assign \new_[35529]_  = ~A169 & \new_[35528]_ ;
  assign \new_[35533]_  = ~A233 & A200;
  assign \new_[35534]_  = ~A199 & \new_[35533]_ ;
  assign \new_[35535]_  = \new_[35534]_  & \new_[35529]_ ;
  assign \new_[35539]_  = ~A265 & ~A236;
  assign \new_[35540]_  = ~A235 & \new_[35539]_ ;
  assign \new_[35544]_  = A299 & A298;
  assign \new_[35545]_  = ~A266 & \new_[35544]_ ;
  assign \new_[35546]_  = \new_[35545]_  & \new_[35540]_ ;
  assign \new_[35550]_  = ~A166 & ~A167;
  assign \new_[35551]_  = ~A169 & \new_[35550]_ ;
  assign \new_[35555]_  = ~A233 & A200;
  assign \new_[35556]_  = ~A199 & \new_[35555]_ ;
  assign \new_[35557]_  = \new_[35556]_  & \new_[35551]_ ;
  assign \new_[35561]_  = ~A265 & ~A236;
  assign \new_[35562]_  = ~A235 & \new_[35561]_ ;
  assign \new_[35566]_  = ~A299 & ~A298;
  assign \new_[35567]_  = ~A266 & \new_[35566]_ ;
  assign \new_[35568]_  = \new_[35567]_  & \new_[35562]_ ;
  assign \new_[35572]_  = ~A166 & ~A167;
  assign \new_[35573]_  = ~A169 & \new_[35572]_ ;
  assign \new_[35577]_  = ~A233 & A200;
  assign \new_[35578]_  = ~A199 & \new_[35577]_ ;
  assign \new_[35579]_  = \new_[35578]_  & \new_[35573]_ ;
  assign \new_[35583]_  = A266 & A265;
  assign \new_[35584]_  = ~A234 & \new_[35583]_ ;
  assign \new_[35588]_  = ~A302 & ~A301;
  assign \new_[35589]_  = A298 & \new_[35588]_ ;
  assign \new_[35590]_  = \new_[35589]_  & \new_[35584]_ ;
  assign \new_[35594]_  = ~A166 & ~A167;
  assign \new_[35595]_  = ~A169 & \new_[35594]_ ;
  assign \new_[35599]_  = ~A233 & A200;
  assign \new_[35600]_  = ~A199 & \new_[35599]_ ;
  assign \new_[35601]_  = \new_[35600]_  & \new_[35595]_ ;
  assign \new_[35605]_  = ~A268 & ~A266;
  assign \new_[35606]_  = ~A234 & \new_[35605]_ ;
  assign \new_[35610]_  = ~A300 & A298;
  assign \new_[35611]_  = ~A269 & \new_[35610]_ ;
  assign \new_[35612]_  = \new_[35611]_  & \new_[35606]_ ;
  assign \new_[35616]_  = ~A166 & ~A167;
  assign \new_[35617]_  = ~A169 & \new_[35616]_ ;
  assign \new_[35621]_  = ~A233 & A200;
  assign \new_[35622]_  = ~A199 & \new_[35621]_ ;
  assign \new_[35623]_  = \new_[35622]_  & \new_[35617]_ ;
  assign \new_[35627]_  = ~A268 & ~A266;
  assign \new_[35628]_  = ~A234 & \new_[35627]_ ;
  assign \new_[35632]_  = A299 & A298;
  assign \new_[35633]_  = ~A269 & \new_[35632]_ ;
  assign \new_[35634]_  = \new_[35633]_  & \new_[35628]_ ;
  assign \new_[35638]_  = ~A166 & ~A167;
  assign \new_[35639]_  = ~A169 & \new_[35638]_ ;
  assign \new_[35643]_  = ~A233 & A200;
  assign \new_[35644]_  = ~A199 & \new_[35643]_ ;
  assign \new_[35645]_  = \new_[35644]_  & \new_[35639]_ ;
  assign \new_[35649]_  = ~A268 & ~A266;
  assign \new_[35650]_  = ~A234 & \new_[35649]_ ;
  assign \new_[35654]_  = ~A299 & ~A298;
  assign \new_[35655]_  = ~A269 & \new_[35654]_ ;
  assign \new_[35656]_  = \new_[35655]_  & \new_[35650]_ ;
  assign \new_[35660]_  = ~A166 & ~A167;
  assign \new_[35661]_  = ~A169 & \new_[35660]_ ;
  assign \new_[35665]_  = ~A233 & A200;
  assign \new_[35666]_  = ~A199 & \new_[35665]_ ;
  assign \new_[35667]_  = \new_[35666]_  & \new_[35661]_ ;
  assign \new_[35671]_  = ~A267 & ~A266;
  assign \new_[35672]_  = ~A234 & \new_[35671]_ ;
  assign \new_[35676]_  = ~A302 & ~A301;
  assign \new_[35677]_  = A298 & \new_[35676]_ ;
  assign \new_[35678]_  = \new_[35677]_  & \new_[35672]_ ;
  assign \new_[35682]_  = ~A166 & ~A167;
  assign \new_[35683]_  = ~A169 & \new_[35682]_ ;
  assign \new_[35687]_  = ~A233 & A200;
  assign \new_[35688]_  = ~A199 & \new_[35687]_ ;
  assign \new_[35689]_  = \new_[35688]_  & \new_[35683]_ ;
  assign \new_[35693]_  = ~A266 & ~A265;
  assign \new_[35694]_  = ~A234 & \new_[35693]_ ;
  assign \new_[35698]_  = ~A302 & ~A301;
  assign \new_[35699]_  = A298 & \new_[35698]_ ;
  assign \new_[35700]_  = \new_[35699]_  & \new_[35694]_ ;
  assign \new_[35704]_  = ~A166 & ~A167;
  assign \new_[35705]_  = ~A169 & \new_[35704]_ ;
  assign \new_[35709]_  = ~A232 & A200;
  assign \new_[35710]_  = ~A199 & \new_[35709]_ ;
  assign \new_[35711]_  = \new_[35710]_  & \new_[35705]_ ;
  assign \new_[35715]_  = A266 & A265;
  assign \new_[35716]_  = ~A233 & \new_[35715]_ ;
  assign \new_[35720]_  = ~A302 & ~A301;
  assign \new_[35721]_  = A298 & \new_[35720]_ ;
  assign \new_[35722]_  = \new_[35721]_  & \new_[35716]_ ;
  assign \new_[35726]_  = ~A166 & ~A167;
  assign \new_[35727]_  = ~A169 & \new_[35726]_ ;
  assign \new_[35731]_  = ~A232 & A200;
  assign \new_[35732]_  = ~A199 & \new_[35731]_ ;
  assign \new_[35733]_  = \new_[35732]_  & \new_[35727]_ ;
  assign \new_[35737]_  = ~A268 & ~A266;
  assign \new_[35738]_  = ~A233 & \new_[35737]_ ;
  assign \new_[35742]_  = ~A300 & A298;
  assign \new_[35743]_  = ~A269 & \new_[35742]_ ;
  assign \new_[35744]_  = \new_[35743]_  & \new_[35738]_ ;
  assign \new_[35748]_  = ~A166 & ~A167;
  assign \new_[35749]_  = ~A169 & \new_[35748]_ ;
  assign \new_[35753]_  = ~A232 & A200;
  assign \new_[35754]_  = ~A199 & \new_[35753]_ ;
  assign \new_[35755]_  = \new_[35754]_  & \new_[35749]_ ;
  assign \new_[35759]_  = ~A268 & ~A266;
  assign \new_[35760]_  = ~A233 & \new_[35759]_ ;
  assign \new_[35764]_  = A299 & A298;
  assign \new_[35765]_  = ~A269 & \new_[35764]_ ;
  assign \new_[35766]_  = \new_[35765]_  & \new_[35760]_ ;
  assign \new_[35770]_  = ~A166 & ~A167;
  assign \new_[35771]_  = ~A169 & \new_[35770]_ ;
  assign \new_[35775]_  = ~A232 & A200;
  assign \new_[35776]_  = ~A199 & \new_[35775]_ ;
  assign \new_[35777]_  = \new_[35776]_  & \new_[35771]_ ;
  assign \new_[35781]_  = ~A268 & ~A266;
  assign \new_[35782]_  = ~A233 & \new_[35781]_ ;
  assign \new_[35786]_  = ~A299 & ~A298;
  assign \new_[35787]_  = ~A269 & \new_[35786]_ ;
  assign \new_[35788]_  = \new_[35787]_  & \new_[35782]_ ;
  assign \new_[35792]_  = ~A166 & ~A167;
  assign \new_[35793]_  = ~A169 & \new_[35792]_ ;
  assign \new_[35797]_  = ~A232 & A200;
  assign \new_[35798]_  = ~A199 & \new_[35797]_ ;
  assign \new_[35799]_  = \new_[35798]_  & \new_[35793]_ ;
  assign \new_[35803]_  = ~A267 & ~A266;
  assign \new_[35804]_  = ~A233 & \new_[35803]_ ;
  assign \new_[35808]_  = ~A302 & ~A301;
  assign \new_[35809]_  = A298 & \new_[35808]_ ;
  assign \new_[35810]_  = \new_[35809]_  & \new_[35804]_ ;
  assign \new_[35814]_  = ~A166 & ~A167;
  assign \new_[35815]_  = ~A169 & \new_[35814]_ ;
  assign \new_[35819]_  = ~A232 & A200;
  assign \new_[35820]_  = ~A199 & \new_[35819]_ ;
  assign \new_[35821]_  = \new_[35820]_  & \new_[35815]_ ;
  assign \new_[35825]_  = ~A266 & ~A265;
  assign \new_[35826]_  = ~A233 & \new_[35825]_ ;
  assign \new_[35830]_  = ~A302 & ~A301;
  assign \new_[35831]_  = A298 & \new_[35830]_ ;
  assign \new_[35832]_  = \new_[35831]_  & \new_[35826]_ ;
  assign \new_[35836]_  = A167 & ~A168;
  assign \new_[35837]_  = ~A169 & \new_[35836]_ ;
  assign \new_[35841]_  = A200 & ~A199;
  assign \new_[35842]_  = A166 & \new_[35841]_ ;
  assign \new_[35843]_  = \new_[35842]_  & \new_[35837]_ ;
  assign \new_[35847]_  = A265 & A233;
  assign \new_[35848]_  = A232 & \new_[35847]_ ;
  assign \new_[35852]_  = ~A300 & ~A299;
  assign \new_[35853]_  = ~A267 & \new_[35852]_ ;
  assign \new_[35854]_  = \new_[35853]_  & \new_[35848]_ ;
  assign \new_[35858]_  = A167 & ~A168;
  assign \new_[35859]_  = ~A169 & \new_[35858]_ ;
  assign \new_[35863]_  = A200 & ~A199;
  assign \new_[35864]_  = A166 & \new_[35863]_ ;
  assign \new_[35865]_  = \new_[35864]_  & \new_[35859]_ ;
  assign \new_[35869]_  = A265 & A233;
  assign \new_[35870]_  = A232 & \new_[35869]_ ;
  assign \new_[35874]_  = A299 & A298;
  assign \new_[35875]_  = ~A267 & \new_[35874]_ ;
  assign \new_[35876]_  = \new_[35875]_  & \new_[35870]_ ;
  assign \new_[35880]_  = A167 & ~A168;
  assign \new_[35881]_  = ~A169 & \new_[35880]_ ;
  assign \new_[35885]_  = A200 & ~A199;
  assign \new_[35886]_  = A166 & \new_[35885]_ ;
  assign \new_[35887]_  = \new_[35886]_  & \new_[35881]_ ;
  assign \new_[35891]_  = A265 & A233;
  assign \new_[35892]_  = A232 & \new_[35891]_ ;
  assign \new_[35896]_  = ~A299 & ~A298;
  assign \new_[35897]_  = ~A267 & \new_[35896]_ ;
  assign \new_[35898]_  = \new_[35897]_  & \new_[35892]_ ;
  assign \new_[35902]_  = A167 & ~A168;
  assign \new_[35903]_  = ~A169 & \new_[35902]_ ;
  assign \new_[35907]_  = A200 & ~A199;
  assign \new_[35908]_  = A166 & \new_[35907]_ ;
  assign \new_[35909]_  = \new_[35908]_  & \new_[35903]_ ;
  assign \new_[35913]_  = A265 & A233;
  assign \new_[35914]_  = A232 & \new_[35913]_ ;
  assign \new_[35918]_  = ~A300 & ~A299;
  assign \new_[35919]_  = A266 & \new_[35918]_ ;
  assign \new_[35920]_  = \new_[35919]_  & \new_[35914]_ ;
  assign \new_[35924]_  = A167 & ~A168;
  assign \new_[35925]_  = ~A169 & \new_[35924]_ ;
  assign \new_[35929]_  = A200 & ~A199;
  assign \new_[35930]_  = A166 & \new_[35929]_ ;
  assign \new_[35931]_  = \new_[35930]_  & \new_[35925]_ ;
  assign \new_[35935]_  = A265 & A233;
  assign \new_[35936]_  = A232 & \new_[35935]_ ;
  assign \new_[35940]_  = A299 & A298;
  assign \new_[35941]_  = A266 & \new_[35940]_ ;
  assign \new_[35942]_  = \new_[35941]_  & \new_[35936]_ ;
  assign \new_[35946]_  = A167 & ~A168;
  assign \new_[35947]_  = ~A169 & \new_[35946]_ ;
  assign \new_[35951]_  = A200 & ~A199;
  assign \new_[35952]_  = A166 & \new_[35951]_ ;
  assign \new_[35953]_  = \new_[35952]_  & \new_[35947]_ ;
  assign \new_[35957]_  = A265 & A233;
  assign \new_[35958]_  = A232 & \new_[35957]_ ;
  assign \new_[35962]_  = ~A299 & ~A298;
  assign \new_[35963]_  = A266 & \new_[35962]_ ;
  assign \new_[35964]_  = \new_[35963]_  & \new_[35958]_ ;
  assign \new_[35968]_  = A167 & ~A168;
  assign \new_[35969]_  = ~A169 & \new_[35968]_ ;
  assign \new_[35973]_  = A200 & ~A199;
  assign \new_[35974]_  = A166 & \new_[35973]_ ;
  assign \new_[35975]_  = \new_[35974]_  & \new_[35969]_ ;
  assign \new_[35979]_  = ~A265 & A233;
  assign \new_[35980]_  = A232 & \new_[35979]_ ;
  assign \new_[35984]_  = ~A300 & ~A299;
  assign \new_[35985]_  = ~A266 & \new_[35984]_ ;
  assign \new_[35986]_  = \new_[35985]_  & \new_[35980]_ ;
  assign \new_[35990]_  = A167 & ~A168;
  assign \new_[35991]_  = ~A169 & \new_[35990]_ ;
  assign \new_[35995]_  = A200 & ~A199;
  assign \new_[35996]_  = A166 & \new_[35995]_ ;
  assign \new_[35997]_  = \new_[35996]_  & \new_[35991]_ ;
  assign \new_[36001]_  = ~A265 & A233;
  assign \new_[36002]_  = A232 & \new_[36001]_ ;
  assign \new_[36006]_  = A299 & A298;
  assign \new_[36007]_  = ~A266 & \new_[36006]_ ;
  assign \new_[36008]_  = \new_[36007]_  & \new_[36002]_ ;
  assign \new_[36012]_  = A167 & ~A168;
  assign \new_[36013]_  = ~A169 & \new_[36012]_ ;
  assign \new_[36017]_  = A200 & ~A199;
  assign \new_[36018]_  = A166 & \new_[36017]_ ;
  assign \new_[36019]_  = \new_[36018]_  & \new_[36013]_ ;
  assign \new_[36023]_  = ~A265 & A233;
  assign \new_[36024]_  = A232 & \new_[36023]_ ;
  assign \new_[36028]_  = ~A299 & ~A298;
  assign \new_[36029]_  = ~A266 & \new_[36028]_ ;
  assign \new_[36030]_  = \new_[36029]_  & \new_[36024]_ ;
  assign \new_[36034]_  = A167 & ~A168;
  assign \new_[36035]_  = ~A169 & \new_[36034]_ ;
  assign \new_[36039]_  = A200 & ~A199;
  assign \new_[36040]_  = A166 & \new_[36039]_ ;
  assign \new_[36041]_  = \new_[36040]_  & \new_[36035]_ ;
  assign \new_[36045]_  = A298 & A233;
  assign \new_[36046]_  = ~A232 & \new_[36045]_ ;
  assign \new_[36050]_  = A301 & A300;
  assign \new_[36051]_  = ~A299 & \new_[36050]_ ;
  assign \new_[36052]_  = \new_[36051]_  & \new_[36046]_ ;
  assign \new_[36056]_  = A167 & ~A168;
  assign \new_[36057]_  = ~A169 & \new_[36056]_ ;
  assign \new_[36061]_  = A200 & ~A199;
  assign \new_[36062]_  = A166 & \new_[36061]_ ;
  assign \new_[36063]_  = \new_[36062]_  & \new_[36057]_ ;
  assign \new_[36067]_  = A298 & A233;
  assign \new_[36068]_  = ~A232 & \new_[36067]_ ;
  assign \new_[36072]_  = A302 & A300;
  assign \new_[36073]_  = ~A299 & \new_[36072]_ ;
  assign \new_[36074]_  = \new_[36073]_  & \new_[36068]_ ;
  assign \new_[36078]_  = A167 & ~A168;
  assign \new_[36079]_  = ~A169 & \new_[36078]_ ;
  assign \new_[36083]_  = A200 & ~A199;
  assign \new_[36084]_  = A166 & \new_[36083]_ ;
  assign \new_[36085]_  = \new_[36084]_  & \new_[36079]_ ;
  assign \new_[36089]_  = A265 & A233;
  assign \new_[36090]_  = ~A232 & \new_[36089]_ ;
  assign \new_[36094]_  = A268 & A267;
  assign \new_[36095]_  = ~A266 & \new_[36094]_ ;
  assign \new_[36096]_  = \new_[36095]_  & \new_[36090]_ ;
  assign \new_[36100]_  = A167 & ~A168;
  assign \new_[36101]_  = ~A169 & \new_[36100]_ ;
  assign \new_[36105]_  = A200 & ~A199;
  assign \new_[36106]_  = A166 & \new_[36105]_ ;
  assign \new_[36107]_  = \new_[36106]_  & \new_[36101]_ ;
  assign \new_[36111]_  = A265 & A233;
  assign \new_[36112]_  = ~A232 & \new_[36111]_ ;
  assign \new_[36116]_  = A269 & A267;
  assign \new_[36117]_  = ~A266 & \new_[36116]_ ;
  assign \new_[36118]_  = \new_[36117]_  & \new_[36112]_ ;
  assign \new_[36122]_  = A167 & ~A168;
  assign \new_[36123]_  = ~A169 & \new_[36122]_ ;
  assign \new_[36127]_  = A200 & ~A199;
  assign \new_[36128]_  = A166 & \new_[36127]_ ;
  assign \new_[36129]_  = \new_[36128]_  & \new_[36123]_ ;
  assign \new_[36133]_  = A265 & ~A234;
  assign \new_[36134]_  = ~A233 & \new_[36133]_ ;
  assign \new_[36138]_  = ~A300 & A298;
  assign \new_[36139]_  = A266 & \new_[36138]_ ;
  assign \new_[36140]_  = \new_[36139]_  & \new_[36134]_ ;
  assign \new_[36144]_  = A167 & ~A168;
  assign \new_[36145]_  = ~A169 & \new_[36144]_ ;
  assign \new_[36149]_  = A200 & ~A199;
  assign \new_[36150]_  = A166 & \new_[36149]_ ;
  assign \new_[36151]_  = \new_[36150]_  & \new_[36145]_ ;
  assign \new_[36155]_  = A265 & ~A234;
  assign \new_[36156]_  = ~A233 & \new_[36155]_ ;
  assign \new_[36160]_  = A299 & A298;
  assign \new_[36161]_  = A266 & \new_[36160]_ ;
  assign \new_[36162]_  = \new_[36161]_  & \new_[36156]_ ;
  assign \new_[36166]_  = A167 & ~A168;
  assign \new_[36167]_  = ~A169 & \new_[36166]_ ;
  assign \new_[36171]_  = A200 & ~A199;
  assign \new_[36172]_  = A166 & \new_[36171]_ ;
  assign \new_[36173]_  = \new_[36172]_  & \new_[36167]_ ;
  assign \new_[36177]_  = A265 & ~A234;
  assign \new_[36178]_  = ~A233 & \new_[36177]_ ;
  assign \new_[36182]_  = ~A299 & ~A298;
  assign \new_[36183]_  = A266 & \new_[36182]_ ;
  assign \new_[36184]_  = \new_[36183]_  & \new_[36178]_ ;
  assign \new_[36188]_  = A167 & ~A168;
  assign \new_[36189]_  = ~A169 & \new_[36188]_ ;
  assign \new_[36193]_  = A200 & ~A199;
  assign \new_[36194]_  = A166 & \new_[36193]_ ;
  assign \new_[36195]_  = \new_[36194]_  & \new_[36189]_ ;
  assign \new_[36199]_  = ~A266 & ~A234;
  assign \new_[36200]_  = ~A233 & \new_[36199]_ ;
  assign \new_[36204]_  = ~A300 & A298;
  assign \new_[36205]_  = ~A267 & \new_[36204]_ ;
  assign \new_[36206]_  = \new_[36205]_  & \new_[36200]_ ;
  assign \new_[36210]_  = A167 & ~A168;
  assign \new_[36211]_  = ~A169 & \new_[36210]_ ;
  assign \new_[36215]_  = A200 & ~A199;
  assign \new_[36216]_  = A166 & \new_[36215]_ ;
  assign \new_[36217]_  = \new_[36216]_  & \new_[36211]_ ;
  assign \new_[36221]_  = ~A266 & ~A234;
  assign \new_[36222]_  = ~A233 & \new_[36221]_ ;
  assign \new_[36226]_  = A299 & A298;
  assign \new_[36227]_  = ~A267 & \new_[36226]_ ;
  assign \new_[36228]_  = \new_[36227]_  & \new_[36222]_ ;
  assign \new_[36232]_  = A167 & ~A168;
  assign \new_[36233]_  = ~A169 & \new_[36232]_ ;
  assign \new_[36237]_  = A200 & ~A199;
  assign \new_[36238]_  = A166 & \new_[36237]_ ;
  assign \new_[36239]_  = \new_[36238]_  & \new_[36233]_ ;
  assign \new_[36243]_  = ~A266 & ~A234;
  assign \new_[36244]_  = ~A233 & \new_[36243]_ ;
  assign \new_[36248]_  = ~A299 & ~A298;
  assign \new_[36249]_  = ~A267 & \new_[36248]_ ;
  assign \new_[36250]_  = \new_[36249]_  & \new_[36244]_ ;
  assign \new_[36254]_  = A167 & ~A168;
  assign \new_[36255]_  = ~A169 & \new_[36254]_ ;
  assign \new_[36259]_  = A200 & ~A199;
  assign \new_[36260]_  = A166 & \new_[36259]_ ;
  assign \new_[36261]_  = \new_[36260]_  & \new_[36255]_ ;
  assign \new_[36265]_  = ~A265 & ~A234;
  assign \new_[36266]_  = ~A233 & \new_[36265]_ ;
  assign \new_[36270]_  = ~A300 & A298;
  assign \new_[36271]_  = ~A266 & \new_[36270]_ ;
  assign \new_[36272]_  = \new_[36271]_  & \new_[36266]_ ;
  assign \new_[36276]_  = A167 & ~A168;
  assign \new_[36277]_  = ~A169 & \new_[36276]_ ;
  assign \new_[36281]_  = A200 & ~A199;
  assign \new_[36282]_  = A166 & \new_[36281]_ ;
  assign \new_[36283]_  = \new_[36282]_  & \new_[36277]_ ;
  assign \new_[36287]_  = ~A265 & ~A234;
  assign \new_[36288]_  = ~A233 & \new_[36287]_ ;
  assign \new_[36292]_  = A299 & A298;
  assign \new_[36293]_  = ~A266 & \new_[36292]_ ;
  assign \new_[36294]_  = \new_[36293]_  & \new_[36288]_ ;
  assign \new_[36298]_  = A167 & ~A168;
  assign \new_[36299]_  = ~A169 & \new_[36298]_ ;
  assign \new_[36303]_  = A200 & ~A199;
  assign \new_[36304]_  = A166 & \new_[36303]_ ;
  assign \new_[36305]_  = \new_[36304]_  & \new_[36299]_ ;
  assign \new_[36309]_  = ~A265 & ~A234;
  assign \new_[36310]_  = ~A233 & \new_[36309]_ ;
  assign \new_[36314]_  = ~A299 & ~A298;
  assign \new_[36315]_  = ~A266 & \new_[36314]_ ;
  assign \new_[36316]_  = \new_[36315]_  & \new_[36310]_ ;
  assign \new_[36320]_  = A167 & ~A168;
  assign \new_[36321]_  = ~A169 & \new_[36320]_ ;
  assign \new_[36325]_  = A200 & ~A199;
  assign \new_[36326]_  = A166 & \new_[36325]_ ;
  assign \new_[36327]_  = \new_[36326]_  & \new_[36321]_ ;
  assign \new_[36331]_  = A234 & ~A233;
  assign \new_[36332]_  = A232 & \new_[36331]_ ;
  assign \new_[36336]_  = A299 & ~A298;
  assign \new_[36337]_  = A235 & \new_[36336]_ ;
  assign \new_[36338]_  = \new_[36337]_  & \new_[36332]_ ;
  assign \new_[36342]_  = A167 & ~A168;
  assign \new_[36343]_  = ~A169 & \new_[36342]_ ;
  assign \new_[36347]_  = A200 & ~A199;
  assign \new_[36348]_  = A166 & \new_[36347]_ ;
  assign \new_[36349]_  = \new_[36348]_  & \new_[36343]_ ;
  assign \new_[36353]_  = A234 & ~A233;
  assign \new_[36354]_  = A232 & \new_[36353]_ ;
  assign \new_[36358]_  = A266 & ~A265;
  assign \new_[36359]_  = A235 & \new_[36358]_ ;
  assign \new_[36360]_  = \new_[36359]_  & \new_[36354]_ ;
  assign \new_[36364]_  = A167 & ~A168;
  assign \new_[36365]_  = ~A169 & \new_[36364]_ ;
  assign \new_[36369]_  = A200 & ~A199;
  assign \new_[36370]_  = A166 & \new_[36369]_ ;
  assign \new_[36371]_  = \new_[36370]_  & \new_[36365]_ ;
  assign \new_[36375]_  = A234 & ~A233;
  assign \new_[36376]_  = A232 & \new_[36375]_ ;
  assign \new_[36380]_  = A299 & ~A298;
  assign \new_[36381]_  = A236 & \new_[36380]_ ;
  assign \new_[36382]_  = \new_[36381]_  & \new_[36376]_ ;
  assign \new_[36386]_  = A167 & ~A168;
  assign \new_[36387]_  = ~A169 & \new_[36386]_ ;
  assign \new_[36391]_  = A200 & ~A199;
  assign \new_[36392]_  = A166 & \new_[36391]_ ;
  assign \new_[36393]_  = \new_[36392]_  & \new_[36387]_ ;
  assign \new_[36397]_  = A234 & ~A233;
  assign \new_[36398]_  = A232 & \new_[36397]_ ;
  assign \new_[36402]_  = A266 & ~A265;
  assign \new_[36403]_  = A236 & \new_[36402]_ ;
  assign \new_[36404]_  = \new_[36403]_  & \new_[36398]_ ;
  assign \new_[36408]_  = A167 & ~A168;
  assign \new_[36409]_  = ~A169 & \new_[36408]_ ;
  assign \new_[36413]_  = A200 & ~A199;
  assign \new_[36414]_  = A166 & \new_[36413]_ ;
  assign \new_[36415]_  = \new_[36414]_  & \new_[36409]_ ;
  assign \new_[36419]_  = A265 & ~A233;
  assign \new_[36420]_  = ~A232 & \new_[36419]_ ;
  assign \new_[36424]_  = ~A300 & A298;
  assign \new_[36425]_  = A266 & \new_[36424]_ ;
  assign \new_[36426]_  = \new_[36425]_  & \new_[36420]_ ;
  assign \new_[36430]_  = A167 & ~A168;
  assign \new_[36431]_  = ~A169 & \new_[36430]_ ;
  assign \new_[36435]_  = A200 & ~A199;
  assign \new_[36436]_  = A166 & \new_[36435]_ ;
  assign \new_[36437]_  = \new_[36436]_  & \new_[36431]_ ;
  assign \new_[36441]_  = A265 & ~A233;
  assign \new_[36442]_  = ~A232 & \new_[36441]_ ;
  assign \new_[36446]_  = A299 & A298;
  assign \new_[36447]_  = A266 & \new_[36446]_ ;
  assign \new_[36448]_  = \new_[36447]_  & \new_[36442]_ ;
  assign \new_[36452]_  = A167 & ~A168;
  assign \new_[36453]_  = ~A169 & \new_[36452]_ ;
  assign \new_[36457]_  = A200 & ~A199;
  assign \new_[36458]_  = A166 & \new_[36457]_ ;
  assign \new_[36459]_  = \new_[36458]_  & \new_[36453]_ ;
  assign \new_[36463]_  = A265 & ~A233;
  assign \new_[36464]_  = ~A232 & \new_[36463]_ ;
  assign \new_[36468]_  = ~A299 & ~A298;
  assign \new_[36469]_  = A266 & \new_[36468]_ ;
  assign \new_[36470]_  = \new_[36469]_  & \new_[36464]_ ;
  assign \new_[36474]_  = A167 & ~A168;
  assign \new_[36475]_  = ~A169 & \new_[36474]_ ;
  assign \new_[36479]_  = A200 & ~A199;
  assign \new_[36480]_  = A166 & \new_[36479]_ ;
  assign \new_[36481]_  = \new_[36480]_  & \new_[36475]_ ;
  assign \new_[36485]_  = ~A266 & ~A233;
  assign \new_[36486]_  = ~A232 & \new_[36485]_ ;
  assign \new_[36490]_  = ~A300 & A298;
  assign \new_[36491]_  = ~A267 & \new_[36490]_ ;
  assign \new_[36492]_  = \new_[36491]_  & \new_[36486]_ ;
  assign \new_[36496]_  = A167 & ~A168;
  assign \new_[36497]_  = ~A169 & \new_[36496]_ ;
  assign \new_[36501]_  = A200 & ~A199;
  assign \new_[36502]_  = A166 & \new_[36501]_ ;
  assign \new_[36503]_  = \new_[36502]_  & \new_[36497]_ ;
  assign \new_[36507]_  = ~A266 & ~A233;
  assign \new_[36508]_  = ~A232 & \new_[36507]_ ;
  assign \new_[36512]_  = A299 & A298;
  assign \new_[36513]_  = ~A267 & \new_[36512]_ ;
  assign \new_[36514]_  = \new_[36513]_  & \new_[36508]_ ;
  assign \new_[36518]_  = A167 & ~A168;
  assign \new_[36519]_  = ~A169 & \new_[36518]_ ;
  assign \new_[36523]_  = A200 & ~A199;
  assign \new_[36524]_  = A166 & \new_[36523]_ ;
  assign \new_[36525]_  = \new_[36524]_  & \new_[36519]_ ;
  assign \new_[36529]_  = ~A266 & ~A233;
  assign \new_[36530]_  = ~A232 & \new_[36529]_ ;
  assign \new_[36534]_  = ~A299 & ~A298;
  assign \new_[36535]_  = ~A267 & \new_[36534]_ ;
  assign \new_[36536]_  = \new_[36535]_  & \new_[36530]_ ;
  assign \new_[36540]_  = A167 & ~A168;
  assign \new_[36541]_  = ~A169 & \new_[36540]_ ;
  assign \new_[36545]_  = A200 & ~A199;
  assign \new_[36546]_  = A166 & \new_[36545]_ ;
  assign \new_[36547]_  = \new_[36546]_  & \new_[36541]_ ;
  assign \new_[36551]_  = ~A265 & ~A233;
  assign \new_[36552]_  = ~A232 & \new_[36551]_ ;
  assign \new_[36556]_  = ~A300 & A298;
  assign \new_[36557]_  = ~A266 & \new_[36556]_ ;
  assign \new_[36558]_  = \new_[36557]_  & \new_[36552]_ ;
  assign \new_[36562]_  = A167 & ~A168;
  assign \new_[36563]_  = ~A169 & \new_[36562]_ ;
  assign \new_[36567]_  = A200 & ~A199;
  assign \new_[36568]_  = A166 & \new_[36567]_ ;
  assign \new_[36569]_  = \new_[36568]_  & \new_[36563]_ ;
  assign \new_[36573]_  = ~A265 & ~A233;
  assign \new_[36574]_  = ~A232 & \new_[36573]_ ;
  assign \new_[36578]_  = A299 & A298;
  assign \new_[36579]_  = ~A266 & \new_[36578]_ ;
  assign \new_[36580]_  = \new_[36579]_  & \new_[36574]_ ;
  assign \new_[36584]_  = A167 & ~A168;
  assign \new_[36585]_  = ~A169 & \new_[36584]_ ;
  assign \new_[36589]_  = A200 & ~A199;
  assign \new_[36590]_  = A166 & \new_[36589]_ ;
  assign \new_[36591]_  = \new_[36590]_  & \new_[36585]_ ;
  assign \new_[36595]_  = ~A265 & ~A233;
  assign \new_[36596]_  = ~A232 & \new_[36595]_ ;
  assign \new_[36600]_  = ~A299 & ~A298;
  assign \new_[36601]_  = ~A266 & \new_[36600]_ ;
  assign \new_[36602]_  = \new_[36601]_  & \new_[36596]_ ;
  assign \new_[36606]_  = A167 & ~A168;
  assign \new_[36607]_  = ~A169 & \new_[36606]_ ;
  assign \new_[36611]_  = ~A200 & A199;
  assign \new_[36612]_  = A166 & \new_[36611]_ ;
  assign \new_[36613]_  = \new_[36612]_  & \new_[36607]_ ;
  assign \new_[36617]_  = ~A232 & A202;
  assign \new_[36618]_  = A201 & \new_[36617]_ ;
  assign \new_[36622]_  = A299 & ~A298;
  assign \new_[36623]_  = A233 & \new_[36622]_ ;
  assign \new_[36624]_  = \new_[36623]_  & \new_[36618]_ ;
  assign \new_[36628]_  = A167 & ~A168;
  assign \new_[36629]_  = ~A169 & \new_[36628]_ ;
  assign \new_[36633]_  = ~A200 & A199;
  assign \new_[36634]_  = A166 & \new_[36633]_ ;
  assign \new_[36635]_  = \new_[36634]_  & \new_[36629]_ ;
  assign \new_[36639]_  = ~A232 & A202;
  assign \new_[36640]_  = A201 & \new_[36639]_ ;
  assign \new_[36644]_  = A266 & ~A265;
  assign \new_[36645]_  = A233 & \new_[36644]_ ;
  assign \new_[36646]_  = \new_[36645]_  & \new_[36640]_ ;
  assign \new_[36650]_  = A167 & ~A168;
  assign \new_[36651]_  = ~A169 & \new_[36650]_ ;
  assign \new_[36655]_  = ~A200 & A199;
  assign \new_[36656]_  = A166 & \new_[36655]_ ;
  assign \new_[36657]_  = \new_[36656]_  & \new_[36651]_ ;
  assign \new_[36661]_  = ~A232 & A203;
  assign \new_[36662]_  = A201 & \new_[36661]_ ;
  assign \new_[36666]_  = A299 & ~A298;
  assign \new_[36667]_  = A233 & \new_[36666]_ ;
  assign \new_[36668]_  = \new_[36667]_  & \new_[36662]_ ;
  assign \new_[36672]_  = A167 & ~A168;
  assign \new_[36673]_  = ~A169 & \new_[36672]_ ;
  assign \new_[36677]_  = ~A200 & A199;
  assign \new_[36678]_  = A166 & \new_[36677]_ ;
  assign \new_[36679]_  = \new_[36678]_  & \new_[36673]_ ;
  assign \new_[36683]_  = ~A232 & A203;
  assign \new_[36684]_  = A201 & \new_[36683]_ ;
  assign \new_[36688]_  = A266 & ~A265;
  assign \new_[36689]_  = A233 & \new_[36688]_ ;
  assign \new_[36690]_  = \new_[36689]_  & \new_[36684]_ ;
  assign \new_[36694]_  = A167 & ~A169;
  assign \new_[36695]_  = A170 & \new_[36694]_ ;
  assign \new_[36699]_  = A200 & A199;
  assign \new_[36700]_  = ~A166 & \new_[36699]_ ;
  assign \new_[36701]_  = \new_[36700]_  & \new_[36695]_ ;
  assign \new_[36705]_  = A265 & A233;
  assign \new_[36706]_  = A232 & \new_[36705]_ ;
  assign \new_[36710]_  = ~A300 & ~A299;
  assign \new_[36711]_  = ~A267 & \new_[36710]_ ;
  assign \new_[36712]_  = \new_[36711]_  & \new_[36706]_ ;
  assign \new_[36716]_  = A167 & ~A169;
  assign \new_[36717]_  = A170 & \new_[36716]_ ;
  assign \new_[36721]_  = A200 & A199;
  assign \new_[36722]_  = ~A166 & \new_[36721]_ ;
  assign \new_[36723]_  = \new_[36722]_  & \new_[36717]_ ;
  assign \new_[36727]_  = A265 & A233;
  assign \new_[36728]_  = A232 & \new_[36727]_ ;
  assign \new_[36732]_  = A299 & A298;
  assign \new_[36733]_  = ~A267 & \new_[36732]_ ;
  assign \new_[36734]_  = \new_[36733]_  & \new_[36728]_ ;
  assign \new_[36738]_  = A167 & ~A169;
  assign \new_[36739]_  = A170 & \new_[36738]_ ;
  assign \new_[36743]_  = A200 & A199;
  assign \new_[36744]_  = ~A166 & \new_[36743]_ ;
  assign \new_[36745]_  = \new_[36744]_  & \new_[36739]_ ;
  assign \new_[36749]_  = A265 & A233;
  assign \new_[36750]_  = A232 & \new_[36749]_ ;
  assign \new_[36754]_  = ~A299 & ~A298;
  assign \new_[36755]_  = ~A267 & \new_[36754]_ ;
  assign \new_[36756]_  = \new_[36755]_  & \new_[36750]_ ;
  assign \new_[36760]_  = A167 & ~A169;
  assign \new_[36761]_  = A170 & \new_[36760]_ ;
  assign \new_[36765]_  = A200 & A199;
  assign \new_[36766]_  = ~A166 & \new_[36765]_ ;
  assign \new_[36767]_  = \new_[36766]_  & \new_[36761]_ ;
  assign \new_[36771]_  = A265 & A233;
  assign \new_[36772]_  = A232 & \new_[36771]_ ;
  assign \new_[36776]_  = ~A300 & ~A299;
  assign \new_[36777]_  = A266 & \new_[36776]_ ;
  assign \new_[36778]_  = \new_[36777]_  & \new_[36772]_ ;
  assign \new_[36782]_  = A167 & ~A169;
  assign \new_[36783]_  = A170 & \new_[36782]_ ;
  assign \new_[36787]_  = A200 & A199;
  assign \new_[36788]_  = ~A166 & \new_[36787]_ ;
  assign \new_[36789]_  = \new_[36788]_  & \new_[36783]_ ;
  assign \new_[36793]_  = A265 & A233;
  assign \new_[36794]_  = A232 & \new_[36793]_ ;
  assign \new_[36798]_  = A299 & A298;
  assign \new_[36799]_  = A266 & \new_[36798]_ ;
  assign \new_[36800]_  = \new_[36799]_  & \new_[36794]_ ;
  assign \new_[36804]_  = A167 & ~A169;
  assign \new_[36805]_  = A170 & \new_[36804]_ ;
  assign \new_[36809]_  = A200 & A199;
  assign \new_[36810]_  = ~A166 & \new_[36809]_ ;
  assign \new_[36811]_  = \new_[36810]_  & \new_[36805]_ ;
  assign \new_[36815]_  = A265 & A233;
  assign \new_[36816]_  = A232 & \new_[36815]_ ;
  assign \new_[36820]_  = ~A299 & ~A298;
  assign \new_[36821]_  = A266 & \new_[36820]_ ;
  assign \new_[36822]_  = \new_[36821]_  & \new_[36816]_ ;
  assign \new_[36826]_  = A167 & ~A169;
  assign \new_[36827]_  = A170 & \new_[36826]_ ;
  assign \new_[36831]_  = A200 & A199;
  assign \new_[36832]_  = ~A166 & \new_[36831]_ ;
  assign \new_[36833]_  = \new_[36832]_  & \new_[36827]_ ;
  assign \new_[36837]_  = ~A265 & A233;
  assign \new_[36838]_  = A232 & \new_[36837]_ ;
  assign \new_[36842]_  = ~A300 & ~A299;
  assign \new_[36843]_  = ~A266 & \new_[36842]_ ;
  assign \new_[36844]_  = \new_[36843]_  & \new_[36838]_ ;
  assign \new_[36848]_  = A167 & ~A169;
  assign \new_[36849]_  = A170 & \new_[36848]_ ;
  assign \new_[36853]_  = A200 & A199;
  assign \new_[36854]_  = ~A166 & \new_[36853]_ ;
  assign \new_[36855]_  = \new_[36854]_  & \new_[36849]_ ;
  assign \new_[36859]_  = ~A265 & A233;
  assign \new_[36860]_  = A232 & \new_[36859]_ ;
  assign \new_[36864]_  = A299 & A298;
  assign \new_[36865]_  = ~A266 & \new_[36864]_ ;
  assign \new_[36866]_  = \new_[36865]_  & \new_[36860]_ ;
  assign \new_[36870]_  = A167 & ~A169;
  assign \new_[36871]_  = A170 & \new_[36870]_ ;
  assign \new_[36875]_  = A200 & A199;
  assign \new_[36876]_  = ~A166 & \new_[36875]_ ;
  assign \new_[36877]_  = \new_[36876]_  & \new_[36871]_ ;
  assign \new_[36881]_  = ~A265 & A233;
  assign \new_[36882]_  = A232 & \new_[36881]_ ;
  assign \new_[36886]_  = ~A299 & ~A298;
  assign \new_[36887]_  = ~A266 & \new_[36886]_ ;
  assign \new_[36888]_  = \new_[36887]_  & \new_[36882]_ ;
  assign \new_[36892]_  = A167 & ~A169;
  assign \new_[36893]_  = A170 & \new_[36892]_ ;
  assign \new_[36897]_  = A200 & A199;
  assign \new_[36898]_  = ~A166 & \new_[36897]_ ;
  assign \new_[36899]_  = \new_[36898]_  & \new_[36893]_ ;
  assign \new_[36903]_  = A298 & A233;
  assign \new_[36904]_  = ~A232 & \new_[36903]_ ;
  assign \new_[36908]_  = A301 & A300;
  assign \new_[36909]_  = ~A299 & \new_[36908]_ ;
  assign \new_[36910]_  = \new_[36909]_  & \new_[36904]_ ;
  assign \new_[36914]_  = A167 & ~A169;
  assign \new_[36915]_  = A170 & \new_[36914]_ ;
  assign \new_[36919]_  = A200 & A199;
  assign \new_[36920]_  = ~A166 & \new_[36919]_ ;
  assign \new_[36921]_  = \new_[36920]_  & \new_[36915]_ ;
  assign \new_[36925]_  = A298 & A233;
  assign \new_[36926]_  = ~A232 & \new_[36925]_ ;
  assign \new_[36930]_  = A302 & A300;
  assign \new_[36931]_  = ~A299 & \new_[36930]_ ;
  assign \new_[36932]_  = \new_[36931]_  & \new_[36926]_ ;
  assign \new_[36936]_  = A167 & ~A169;
  assign \new_[36937]_  = A170 & \new_[36936]_ ;
  assign \new_[36941]_  = A200 & A199;
  assign \new_[36942]_  = ~A166 & \new_[36941]_ ;
  assign \new_[36943]_  = \new_[36942]_  & \new_[36937]_ ;
  assign \new_[36947]_  = A265 & A233;
  assign \new_[36948]_  = ~A232 & \new_[36947]_ ;
  assign \new_[36952]_  = A268 & A267;
  assign \new_[36953]_  = ~A266 & \new_[36952]_ ;
  assign \new_[36954]_  = \new_[36953]_  & \new_[36948]_ ;
  assign \new_[36958]_  = A167 & ~A169;
  assign \new_[36959]_  = A170 & \new_[36958]_ ;
  assign \new_[36963]_  = A200 & A199;
  assign \new_[36964]_  = ~A166 & \new_[36963]_ ;
  assign \new_[36965]_  = \new_[36964]_  & \new_[36959]_ ;
  assign \new_[36969]_  = A265 & A233;
  assign \new_[36970]_  = ~A232 & \new_[36969]_ ;
  assign \new_[36974]_  = A269 & A267;
  assign \new_[36975]_  = ~A266 & \new_[36974]_ ;
  assign \new_[36976]_  = \new_[36975]_  & \new_[36970]_ ;
  assign \new_[36980]_  = A167 & ~A169;
  assign \new_[36981]_  = A170 & \new_[36980]_ ;
  assign \new_[36985]_  = A200 & A199;
  assign \new_[36986]_  = ~A166 & \new_[36985]_ ;
  assign \new_[36987]_  = \new_[36986]_  & \new_[36981]_ ;
  assign \new_[36991]_  = A265 & ~A234;
  assign \new_[36992]_  = ~A233 & \new_[36991]_ ;
  assign \new_[36996]_  = ~A300 & A298;
  assign \new_[36997]_  = A266 & \new_[36996]_ ;
  assign \new_[36998]_  = \new_[36997]_  & \new_[36992]_ ;
  assign \new_[37002]_  = A167 & ~A169;
  assign \new_[37003]_  = A170 & \new_[37002]_ ;
  assign \new_[37007]_  = A200 & A199;
  assign \new_[37008]_  = ~A166 & \new_[37007]_ ;
  assign \new_[37009]_  = \new_[37008]_  & \new_[37003]_ ;
  assign \new_[37013]_  = A265 & ~A234;
  assign \new_[37014]_  = ~A233 & \new_[37013]_ ;
  assign \new_[37018]_  = A299 & A298;
  assign \new_[37019]_  = A266 & \new_[37018]_ ;
  assign \new_[37020]_  = \new_[37019]_  & \new_[37014]_ ;
  assign \new_[37024]_  = A167 & ~A169;
  assign \new_[37025]_  = A170 & \new_[37024]_ ;
  assign \new_[37029]_  = A200 & A199;
  assign \new_[37030]_  = ~A166 & \new_[37029]_ ;
  assign \new_[37031]_  = \new_[37030]_  & \new_[37025]_ ;
  assign \new_[37035]_  = A265 & ~A234;
  assign \new_[37036]_  = ~A233 & \new_[37035]_ ;
  assign \new_[37040]_  = ~A299 & ~A298;
  assign \new_[37041]_  = A266 & \new_[37040]_ ;
  assign \new_[37042]_  = \new_[37041]_  & \new_[37036]_ ;
  assign \new_[37046]_  = A167 & ~A169;
  assign \new_[37047]_  = A170 & \new_[37046]_ ;
  assign \new_[37051]_  = A200 & A199;
  assign \new_[37052]_  = ~A166 & \new_[37051]_ ;
  assign \new_[37053]_  = \new_[37052]_  & \new_[37047]_ ;
  assign \new_[37057]_  = ~A266 & ~A234;
  assign \new_[37058]_  = ~A233 & \new_[37057]_ ;
  assign \new_[37062]_  = ~A300 & A298;
  assign \new_[37063]_  = ~A267 & \new_[37062]_ ;
  assign \new_[37064]_  = \new_[37063]_  & \new_[37058]_ ;
  assign \new_[37068]_  = A167 & ~A169;
  assign \new_[37069]_  = A170 & \new_[37068]_ ;
  assign \new_[37073]_  = A200 & A199;
  assign \new_[37074]_  = ~A166 & \new_[37073]_ ;
  assign \new_[37075]_  = \new_[37074]_  & \new_[37069]_ ;
  assign \new_[37079]_  = ~A266 & ~A234;
  assign \new_[37080]_  = ~A233 & \new_[37079]_ ;
  assign \new_[37084]_  = A299 & A298;
  assign \new_[37085]_  = ~A267 & \new_[37084]_ ;
  assign \new_[37086]_  = \new_[37085]_  & \new_[37080]_ ;
  assign \new_[37090]_  = A167 & ~A169;
  assign \new_[37091]_  = A170 & \new_[37090]_ ;
  assign \new_[37095]_  = A200 & A199;
  assign \new_[37096]_  = ~A166 & \new_[37095]_ ;
  assign \new_[37097]_  = \new_[37096]_  & \new_[37091]_ ;
  assign \new_[37101]_  = ~A266 & ~A234;
  assign \new_[37102]_  = ~A233 & \new_[37101]_ ;
  assign \new_[37106]_  = ~A299 & ~A298;
  assign \new_[37107]_  = ~A267 & \new_[37106]_ ;
  assign \new_[37108]_  = \new_[37107]_  & \new_[37102]_ ;
  assign \new_[37112]_  = A167 & ~A169;
  assign \new_[37113]_  = A170 & \new_[37112]_ ;
  assign \new_[37117]_  = A200 & A199;
  assign \new_[37118]_  = ~A166 & \new_[37117]_ ;
  assign \new_[37119]_  = \new_[37118]_  & \new_[37113]_ ;
  assign \new_[37123]_  = ~A265 & ~A234;
  assign \new_[37124]_  = ~A233 & \new_[37123]_ ;
  assign \new_[37128]_  = ~A300 & A298;
  assign \new_[37129]_  = ~A266 & \new_[37128]_ ;
  assign \new_[37130]_  = \new_[37129]_  & \new_[37124]_ ;
  assign \new_[37134]_  = A167 & ~A169;
  assign \new_[37135]_  = A170 & \new_[37134]_ ;
  assign \new_[37139]_  = A200 & A199;
  assign \new_[37140]_  = ~A166 & \new_[37139]_ ;
  assign \new_[37141]_  = \new_[37140]_  & \new_[37135]_ ;
  assign \new_[37145]_  = ~A265 & ~A234;
  assign \new_[37146]_  = ~A233 & \new_[37145]_ ;
  assign \new_[37150]_  = A299 & A298;
  assign \new_[37151]_  = ~A266 & \new_[37150]_ ;
  assign \new_[37152]_  = \new_[37151]_  & \new_[37146]_ ;
  assign \new_[37156]_  = A167 & ~A169;
  assign \new_[37157]_  = A170 & \new_[37156]_ ;
  assign \new_[37161]_  = A200 & A199;
  assign \new_[37162]_  = ~A166 & \new_[37161]_ ;
  assign \new_[37163]_  = \new_[37162]_  & \new_[37157]_ ;
  assign \new_[37167]_  = ~A265 & ~A234;
  assign \new_[37168]_  = ~A233 & \new_[37167]_ ;
  assign \new_[37172]_  = ~A299 & ~A298;
  assign \new_[37173]_  = ~A266 & \new_[37172]_ ;
  assign \new_[37174]_  = \new_[37173]_  & \new_[37168]_ ;
  assign \new_[37178]_  = A167 & ~A169;
  assign \new_[37179]_  = A170 & \new_[37178]_ ;
  assign \new_[37183]_  = A200 & A199;
  assign \new_[37184]_  = ~A166 & \new_[37183]_ ;
  assign \new_[37185]_  = \new_[37184]_  & \new_[37179]_ ;
  assign \new_[37189]_  = A234 & ~A233;
  assign \new_[37190]_  = A232 & \new_[37189]_ ;
  assign \new_[37194]_  = A299 & ~A298;
  assign \new_[37195]_  = A235 & \new_[37194]_ ;
  assign \new_[37196]_  = \new_[37195]_  & \new_[37190]_ ;
  assign \new_[37200]_  = A167 & ~A169;
  assign \new_[37201]_  = A170 & \new_[37200]_ ;
  assign \new_[37205]_  = A200 & A199;
  assign \new_[37206]_  = ~A166 & \new_[37205]_ ;
  assign \new_[37207]_  = \new_[37206]_  & \new_[37201]_ ;
  assign \new_[37211]_  = A234 & ~A233;
  assign \new_[37212]_  = A232 & \new_[37211]_ ;
  assign \new_[37216]_  = A266 & ~A265;
  assign \new_[37217]_  = A235 & \new_[37216]_ ;
  assign \new_[37218]_  = \new_[37217]_  & \new_[37212]_ ;
  assign \new_[37222]_  = A167 & ~A169;
  assign \new_[37223]_  = A170 & \new_[37222]_ ;
  assign \new_[37227]_  = A200 & A199;
  assign \new_[37228]_  = ~A166 & \new_[37227]_ ;
  assign \new_[37229]_  = \new_[37228]_  & \new_[37223]_ ;
  assign \new_[37233]_  = A234 & ~A233;
  assign \new_[37234]_  = A232 & \new_[37233]_ ;
  assign \new_[37238]_  = A299 & ~A298;
  assign \new_[37239]_  = A236 & \new_[37238]_ ;
  assign \new_[37240]_  = \new_[37239]_  & \new_[37234]_ ;
  assign \new_[37244]_  = A167 & ~A169;
  assign \new_[37245]_  = A170 & \new_[37244]_ ;
  assign \new_[37249]_  = A200 & A199;
  assign \new_[37250]_  = ~A166 & \new_[37249]_ ;
  assign \new_[37251]_  = \new_[37250]_  & \new_[37245]_ ;
  assign \new_[37255]_  = A234 & ~A233;
  assign \new_[37256]_  = A232 & \new_[37255]_ ;
  assign \new_[37260]_  = A266 & ~A265;
  assign \new_[37261]_  = A236 & \new_[37260]_ ;
  assign \new_[37262]_  = \new_[37261]_  & \new_[37256]_ ;
  assign \new_[37266]_  = A167 & ~A169;
  assign \new_[37267]_  = A170 & \new_[37266]_ ;
  assign \new_[37271]_  = A200 & A199;
  assign \new_[37272]_  = ~A166 & \new_[37271]_ ;
  assign \new_[37273]_  = \new_[37272]_  & \new_[37267]_ ;
  assign \new_[37277]_  = A265 & ~A233;
  assign \new_[37278]_  = ~A232 & \new_[37277]_ ;
  assign \new_[37282]_  = ~A300 & A298;
  assign \new_[37283]_  = A266 & \new_[37282]_ ;
  assign \new_[37284]_  = \new_[37283]_  & \new_[37278]_ ;
  assign \new_[37288]_  = A167 & ~A169;
  assign \new_[37289]_  = A170 & \new_[37288]_ ;
  assign \new_[37293]_  = A200 & A199;
  assign \new_[37294]_  = ~A166 & \new_[37293]_ ;
  assign \new_[37295]_  = \new_[37294]_  & \new_[37289]_ ;
  assign \new_[37299]_  = A265 & ~A233;
  assign \new_[37300]_  = ~A232 & \new_[37299]_ ;
  assign \new_[37304]_  = A299 & A298;
  assign \new_[37305]_  = A266 & \new_[37304]_ ;
  assign \new_[37306]_  = \new_[37305]_  & \new_[37300]_ ;
  assign \new_[37310]_  = A167 & ~A169;
  assign \new_[37311]_  = A170 & \new_[37310]_ ;
  assign \new_[37315]_  = A200 & A199;
  assign \new_[37316]_  = ~A166 & \new_[37315]_ ;
  assign \new_[37317]_  = \new_[37316]_  & \new_[37311]_ ;
  assign \new_[37321]_  = A265 & ~A233;
  assign \new_[37322]_  = ~A232 & \new_[37321]_ ;
  assign \new_[37326]_  = ~A299 & ~A298;
  assign \new_[37327]_  = A266 & \new_[37326]_ ;
  assign \new_[37328]_  = \new_[37327]_  & \new_[37322]_ ;
  assign \new_[37332]_  = A167 & ~A169;
  assign \new_[37333]_  = A170 & \new_[37332]_ ;
  assign \new_[37337]_  = A200 & A199;
  assign \new_[37338]_  = ~A166 & \new_[37337]_ ;
  assign \new_[37339]_  = \new_[37338]_  & \new_[37333]_ ;
  assign \new_[37343]_  = ~A266 & ~A233;
  assign \new_[37344]_  = ~A232 & \new_[37343]_ ;
  assign \new_[37348]_  = ~A300 & A298;
  assign \new_[37349]_  = ~A267 & \new_[37348]_ ;
  assign \new_[37350]_  = \new_[37349]_  & \new_[37344]_ ;
  assign \new_[37354]_  = A167 & ~A169;
  assign \new_[37355]_  = A170 & \new_[37354]_ ;
  assign \new_[37359]_  = A200 & A199;
  assign \new_[37360]_  = ~A166 & \new_[37359]_ ;
  assign \new_[37361]_  = \new_[37360]_  & \new_[37355]_ ;
  assign \new_[37365]_  = ~A266 & ~A233;
  assign \new_[37366]_  = ~A232 & \new_[37365]_ ;
  assign \new_[37370]_  = A299 & A298;
  assign \new_[37371]_  = ~A267 & \new_[37370]_ ;
  assign \new_[37372]_  = \new_[37371]_  & \new_[37366]_ ;
  assign \new_[37376]_  = A167 & ~A169;
  assign \new_[37377]_  = A170 & \new_[37376]_ ;
  assign \new_[37381]_  = A200 & A199;
  assign \new_[37382]_  = ~A166 & \new_[37381]_ ;
  assign \new_[37383]_  = \new_[37382]_  & \new_[37377]_ ;
  assign \new_[37387]_  = ~A266 & ~A233;
  assign \new_[37388]_  = ~A232 & \new_[37387]_ ;
  assign \new_[37392]_  = ~A299 & ~A298;
  assign \new_[37393]_  = ~A267 & \new_[37392]_ ;
  assign \new_[37394]_  = \new_[37393]_  & \new_[37388]_ ;
  assign \new_[37398]_  = A167 & ~A169;
  assign \new_[37399]_  = A170 & \new_[37398]_ ;
  assign \new_[37403]_  = A200 & A199;
  assign \new_[37404]_  = ~A166 & \new_[37403]_ ;
  assign \new_[37405]_  = \new_[37404]_  & \new_[37399]_ ;
  assign \new_[37409]_  = ~A265 & ~A233;
  assign \new_[37410]_  = ~A232 & \new_[37409]_ ;
  assign \new_[37414]_  = ~A300 & A298;
  assign \new_[37415]_  = ~A266 & \new_[37414]_ ;
  assign \new_[37416]_  = \new_[37415]_  & \new_[37410]_ ;
  assign \new_[37420]_  = A167 & ~A169;
  assign \new_[37421]_  = A170 & \new_[37420]_ ;
  assign \new_[37425]_  = A200 & A199;
  assign \new_[37426]_  = ~A166 & \new_[37425]_ ;
  assign \new_[37427]_  = \new_[37426]_  & \new_[37421]_ ;
  assign \new_[37431]_  = ~A265 & ~A233;
  assign \new_[37432]_  = ~A232 & \new_[37431]_ ;
  assign \new_[37436]_  = A299 & A298;
  assign \new_[37437]_  = ~A266 & \new_[37436]_ ;
  assign \new_[37438]_  = \new_[37437]_  & \new_[37432]_ ;
  assign \new_[37442]_  = A167 & ~A169;
  assign \new_[37443]_  = A170 & \new_[37442]_ ;
  assign \new_[37447]_  = A200 & A199;
  assign \new_[37448]_  = ~A166 & \new_[37447]_ ;
  assign \new_[37449]_  = \new_[37448]_  & \new_[37443]_ ;
  assign \new_[37453]_  = ~A265 & ~A233;
  assign \new_[37454]_  = ~A232 & \new_[37453]_ ;
  assign \new_[37458]_  = ~A299 & ~A298;
  assign \new_[37459]_  = ~A266 & \new_[37458]_ ;
  assign \new_[37460]_  = \new_[37459]_  & \new_[37454]_ ;
  assign \new_[37464]_  = A167 & ~A169;
  assign \new_[37465]_  = A170 & \new_[37464]_ ;
  assign \new_[37469]_  = ~A201 & ~A200;
  assign \new_[37470]_  = ~A166 & \new_[37469]_ ;
  assign \new_[37471]_  = \new_[37470]_  & \new_[37465]_ ;
  assign \new_[37475]_  = A265 & A233;
  assign \new_[37476]_  = A232 & \new_[37475]_ ;
  assign \new_[37480]_  = ~A300 & ~A299;
  assign \new_[37481]_  = ~A267 & \new_[37480]_ ;
  assign \new_[37482]_  = \new_[37481]_  & \new_[37476]_ ;
  assign \new_[37486]_  = A167 & ~A169;
  assign \new_[37487]_  = A170 & \new_[37486]_ ;
  assign \new_[37491]_  = ~A201 & ~A200;
  assign \new_[37492]_  = ~A166 & \new_[37491]_ ;
  assign \new_[37493]_  = \new_[37492]_  & \new_[37487]_ ;
  assign \new_[37497]_  = A265 & A233;
  assign \new_[37498]_  = A232 & \new_[37497]_ ;
  assign \new_[37502]_  = A299 & A298;
  assign \new_[37503]_  = ~A267 & \new_[37502]_ ;
  assign \new_[37504]_  = \new_[37503]_  & \new_[37498]_ ;
  assign \new_[37508]_  = A167 & ~A169;
  assign \new_[37509]_  = A170 & \new_[37508]_ ;
  assign \new_[37513]_  = ~A201 & ~A200;
  assign \new_[37514]_  = ~A166 & \new_[37513]_ ;
  assign \new_[37515]_  = \new_[37514]_  & \new_[37509]_ ;
  assign \new_[37519]_  = A265 & A233;
  assign \new_[37520]_  = A232 & \new_[37519]_ ;
  assign \new_[37524]_  = ~A299 & ~A298;
  assign \new_[37525]_  = ~A267 & \new_[37524]_ ;
  assign \new_[37526]_  = \new_[37525]_  & \new_[37520]_ ;
  assign \new_[37530]_  = A167 & ~A169;
  assign \new_[37531]_  = A170 & \new_[37530]_ ;
  assign \new_[37535]_  = ~A201 & ~A200;
  assign \new_[37536]_  = ~A166 & \new_[37535]_ ;
  assign \new_[37537]_  = \new_[37536]_  & \new_[37531]_ ;
  assign \new_[37541]_  = A265 & A233;
  assign \new_[37542]_  = A232 & \new_[37541]_ ;
  assign \new_[37546]_  = ~A300 & ~A299;
  assign \new_[37547]_  = A266 & \new_[37546]_ ;
  assign \new_[37548]_  = \new_[37547]_  & \new_[37542]_ ;
  assign \new_[37552]_  = A167 & ~A169;
  assign \new_[37553]_  = A170 & \new_[37552]_ ;
  assign \new_[37557]_  = ~A201 & ~A200;
  assign \new_[37558]_  = ~A166 & \new_[37557]_ ;
  assign \new_[37559]_  = \new_[37558]_  & \new_[37553]_ ;
  assign \new_[37563]_  = A265 & A233;
  assign \new_[37564]_  = A232 & \new_[37563]_ ;
  assign \new_[37568]_  = A299 & A298;
  assign \new_[37569]_  = A266 & \new_[37568]_ ;
  assign \new_[37570]_  = \new_[37569]_  & \new_[37564]_ ;
  assign \new_[37574]_  = A167 & ~A169;
  assign \new_[37575]_  = A170 & \new_[37574]_ ;
  assign \new_[37579]_  = ~A201 & ~A200;
  assign \new_[37580]_  = ~A166 & \new_[37579]_ ;
  assign \new_[37581]_  = \new_[37580]_  & \new_[37575]_ ;
  assign \new_[37585]_  = A265 & A233;
  assign \new_[37586]_  = A232 & \new_[37585]_ ;
  assign \new_[37590]_  = ~A299 & ~A298;
  assign \new_[37591]_  = A266 & \new_[37590]_ ;
  assign \new_[37592]_  = \new_[37591]_  & \new_[37586]_ ;
  assign \new_[37596]_  = A167 & ~A169;
  assign \new_[37597]_  = A170 & \new_[37596]_ ;
  assign \new_[37601]_  = ~A201 & ~A200;
  assign \new_[37602]_  = ~A166 & \new_[37601]_ ;
  assign \new_[37603]_  = \new_[37602]_  & \new_[37597]_ ;
  assign \new_[37607]_  = ~A265 & A233;
  assign \new_[37608]_  = A232 & \new_[37607]_ ;
  assign \new_[37612]_  = ~A300 & ~A299;
  assign \new_[37613]_  = ~A266 & \new_[37612]_ ;
  assign \new_[37614]_  = \new_[37613]_  & \new_[37608]_ ;
  assign \new_[37618]_  = A167 & ~A169;
  assign \new_[37619]_  = A170 & \new_[37618]_ ;
  assign \new_[37623]_  = ~A201 & ~A200;
  assign \new_[37624]_  = ~A166 & \new_[37623]_ ;
  assign \new_[37625]_  = \new_[37624]_  & \new_[37619]_ ;
  assign \new_[37629]_  = ~A265 & A233;
  assign \new_[37630]_  = A232 & \new_[37629]_ ;
  assign \new_[37634]_  = A299 & A298;
  assign \new_[37635]_  = ~A266 & \new_[37634]_ ;
  assign \new_[37636]_  = \new_[37635]_  & \new_[37630]_ ;
  assign \new_[37640]_  = A167 & ~A169;
  assign \new_[37641]_  = A170 & \new_[37640]_ ;
  assign \new_[37645]_  = ~A201 & ~A200;
  assign \new_[37646]_  = ~A166 & \new_[37645]_ ;
  assign \new_[37647]_  = \new_[37646]_  & \new_[37641]_ ;
  assign \new_[37651]_  = ~A265 & A233;
  assign \new_[37652]_  = A232 & \new_[37651]_ ;
  assign \new_[37656]_  = ~A299 & ~A298;
  assign \new_[37657]_  = ~A266 & \new_[37656]_ ;
  assign \new_[37658]_  = \new_[37657]_  & \new_[37652]_ ;
  assign \new_[37662]_  = A167 & ~A169;
  assign \new_[37663]_  = A170 & \new_[37662]_ ;
  assign \new_[37667]_  = ~A201 & ~A200;
  assign \new_[37668]_  = ~A166 & \new_[37667]_ ;
  assign \new_[37669]_  = \new_[37668]_  & \new_[37663]_ ;
  assign \new_[37673]_  = A298 & A233;
  assign \new_[37674]_  = ~A232 & \new_[37673]_ ;
  assign \new_[37678]_  = A301 & A300;
  assign \new_[37679]_  = ~A299 & \new_[37678]_ ;
  assign \new_[37680]_  = \new_[37679]_  & \new_[37674]_ ;
  assign \new_[37684]_  = A167 & ~A169;
  assign \new_[37685]_  = A170 & \new_[37684]_ ;
  assign \new_[37689]_  = ~A201 & ~A200;
  assign \new_[37690]_  = ~A166 & \new_[37689]_ ;
  assign \new_[37691]_  = \new_[37690]_  & \new_[37685]_ ;
  assign \new_[37695]_  = A298 & A233;
  assign \new_[37696]_  = ~A232 & \new_[37695]_ ;
  assign \new_[37700]_  = A302 & A300;
  assign \new_[37701]_  = ~A299 & \new_[37700]_ ;
  assign \new_[37702]_  = \new_[37701]_  & \new_[37696]_ ;
  assign \new_[37706]_  = A167 & ~A169;
  assign \new_[37707]_  = A170 & \new_[37706]_ ;
  assign \new_[37711]_  = ~A201 & ~A200;
  assign \new_[37712]_  = ~A166 & \new_[37711]_ ;
  assign \new_[37713]_  = \new_[37712]_  & \new_[37707]_ ;
  assign \new_[37717]_  = A265 & A233;
  assign \new_[37718]_  = ~A232 & \new_[37717]_ ;
  assign \new_[37722]_  = A268 & A267;
  assign \new_[37723]_  = ~A266 & \new_[37722]_ ;
  assign \new_[37724]_  = \new_[37723]_  & \new_[37718]_ ;
  assign \new_[37728]_  = A167 & ~A169;
  assign \new_[37729]_  = A170 & \new_[37728]_ ;
  assign \new_[37733]_  = ~A201 & ~A200;
  assign \new_[37734]_  = ~A166 & \new_[37733]_ ;
  assign \new_[37735]_  = \new_[37734]_  & \new_[37729]_ ;
  assign \new_[37739]_  = A265 & A233;
  assign \new_[37740]_  = ~A232 & \new_[37739]_ ;
  assign \new_[37744]_  = A269 & A267;
  assign \new_[37745]_  = ~A266 & \new_[37744]_ ;
  assign \new_[37746]_  = \new_[37745]_  & \new_[37740]_ ;
  assign \new_[37750]_  = A167 & ~A169;
  assign \new_[37751]_  = A170 & \new_[37750]_ ;
  assign \new_[37755]_  = ~A201 & ~A200;
  assign \new_[37756]_  = ~A166 & \new_[37755]_ ;
  assign \new_[37757]_  = \new_[37756]_  & \new_[37751]_ ;
  assign \new_[37761]_  = A265 & ~A234;
  assign \new_[37762]_  = ~A233 & \new_[37761]_ ;
  assign \new_[37766]_  = ~A300 & A298;
  assign \new_[37767]_  = A266 & \new_[37766]_ ;
  assign \new_[37768]_  = \new_[37767]_  & \new_[37762]_ ;
  assign \new_[37772]_  = A167 & ~A169;
  assign \new_[37773]_  = A170 & \new_[37772]_ ;
  assign \new_[37777]_  = ~A201 & ~A200;
  assign \new_[37778]_  = ~A166 & \new_[37777]_ ;
  assign \new_[37779]_  = \new_[37778]_  & \new_[37773]_ ;
  assign \new_[37783]_  = A265 & ~A234;
  assign \new_[37784]_  = ~A233 & \new_[37783]_ ;
  assign \new_[37788]_  = A299 & A298;
  assign \new_[37789]_  = A266 & \new_[37788]_ ;
  assign \new_[37790]_  = \new_[37789]_  & \new_[37784]_ ;
  assign \new_[37794]_  = A167 & ~A169;
  assign \new_[37795]_  = A170 & \new_[37794]_ ;
  assign \new_[37799]_  = ~A201 & ~A200;
  assign \new_[37800]_  = ~A166 & \new_[37799]_ ;
  assign \new_[37801]_  = \new_[37800]_  & \new_[37795]_ ;
  assign \new_[37805]_  = A265 & ~A234;
  assign \new_[37806]_  = ~A233 & \new_[37805]_ ;
  assign \new_[37810]_  = ~A299 & ~A298;
  assign \new_[37811]_  = A266 & \new_[37810]_ ;
  assign \new_[37812]_  = \new_[37811]_  & \new_[37806]_ ;
  assign \new_[37816]_  = A167 & ~A169;
  assign \new_[37817]_  = A170 & \new_[37816]_ ;
  assign \new_[37821]_  = ~A201 & ~A200;
  assign \new_[37822]_  = ~A166 & \new_[37821]_ ;
  assign \new_[37823]_  = \new_[37822]_  & \new_[37817]_ ;
  assign \new_[37827]_  = ~A266 & ~A234;
  assign \new_[37828]_  = ~A233 & \new_[37827]_ ;
  assign \new_[37832]_  = ~A300 & A298;
  assign \new_[37833]_  = ~A267 & \new_[37832]_ ;
  assign \new_[37834]_  = \new_[37833]_  & \new_[37828]_ ;
  assign \new_[37838]_  = A167 & ~A169;
  assign \new_[37839]_  = A170 & \new_[37838]_ ;
  assign \new_[37843]_  = ~A201 & ~A200;
  assign \new_[37844]_  = ~A166 & \new_[37843]_ ;
  assign \new_[37845]_  = \new_[37844]_  & \new_[37839]_ ;
  assign \new_[37849]_  = ~A266 & ~A234;
  assign \new_[37850]_  = ~A233 & \new_[37849]_ ;
  assign \new_[37854]_  = A299 & A298;
  assign \new_[37855]_  = ~A267 & \new_[37854]_ ;
  assign \new_[37856]_  = \new_[37855]_  & \new_[37850]_ ;
  assign \new_[37860]_  = A167 & ~A169;
  assign \new_[37861]_  = A170 & \new_[37860]_ ;
  assign \new_[37865]_  = ~A201 & ~A200;
  assign \new_[37866]_  = ~A166 & \new_[37865]_ ;
  assign \new_[37867]_  = \new_[37866]_  & \new_[37861]_ ;
  assign \new_[37871]_  = ~A266 & ~A234;
  assign \new_[37872]_  = ~A233 & \new_[37871]_ ;
  assign \new_[37876]_  = ~A299 & ~A298;
  assign \new_[37877]_  = ~A267 & \new_[37876]_ ;
  assign \new_[37878]_  = \new_[37877]_  & \new_[37872]_ ;
  assign \new_[37882]_  = A167 & ~A169;
  assign \new_[37883]_  = A170 & \new_[37882]_ ;
  assign \new_[37887]_  = ~A201 & ~A200;
  assign \new_[37888]_  = ~A166 & \new_[37887]_ ;
  assign \new_[37889]_  = \new_[37888]_  & \new_[37883]_ ;
  assign \new_[37893]_  = ~A265 & ~A234;
  assign \new_[37894]_  = ~A233 & \new_[37893]_ ;
  assign \new_[37898]_  = ~A300 & A298;
  assign \new_[37899]_  = ~A266 & \new_[37898]_ ;
  assign \new_[37900]_  = \new_[37899]_  & \new_[37894]_ ;
  assign \new_[37904]_  = A167 & ~A169;
  assign \new_[37905]_  = A170 & \new_[37904]_ ;
  assign \new_[37909]_  = ~A201 & ~A200;
  assign \new_[37910]_  = ~A166 & \new_[37909]_ ;
  assign \new_[37911]_  = \new_[37910]_  & \new_[37905]_ ;
  assign \new_[37915]_  = ~A265 & ~A234;
  assign \new_[37916]_  = ~A233 & \new_[37915]_ ;
  assign \new_[37920]_  = A299 & A298;
  assign \new_[37921]_  = ~A266 & \new_[37920]_ ;
  assign \new_[37922]_  = \new_[37921]_  & \new_[37916]_ ;
  assign \new_[37926]_  = A167 & ~A169;
  assign \new_[37927]_  = A170 & \new_[37926]_ ;
  assign \new_[37931]_  = ~A201 & ~A200;
  assign \new_[37932]_  = ~A166 & \new_[37931]_ ;
  assign \new_[37933]_  = \new_[37932]_  & \new_[37927]_ ;
  assign \new_[37937]_  = ~A265 & ~A234;
  assign \new_[37938]_  = ~A233 & \new_[37937]_ ;
  assign \new_[37942]_  = ~A299 & ~A298;
  assign \new_[37943]_  = ~A266 & \new_[37942]_ ;
  assign \new_[37944]_  = \new_[37943]_  & \new_[37938]_ ;
  assign \new_[37948]_  = A167 & ~A169;
  assign \new_[37949]_  = A170 & \new_[37948]_ ;
  assign \new_[37953]_  = ~A201 & ~A200;
  assign \new_[37954]_  = ~A166 & \new_[37953]_ ;
  assign \new_[37955]_  = \new_[37954]_  & \new_[37949]_ ;
  assign \new_[37959]_  = A234 & ~A233;
  assign \new_[37960]_  = A232 & \new_[37959]_ ;
  assign \new_[37964]_  = A299 & ~A298;
  assign \new_[37965]_  = A235 & \new_[37964]_ ;
  assign \new_[37966]_  = \new_[37965]_  & \new_[37960]_ ;
  assign \new_[37970]_  = A167 & ~A169;
  assign \new_[37971]_  = A170 & \new_[37970]_ ;
  assign \new_[37975]_  = ~A201 & ~A200;
  assign \new_[37976]_  = ~A166 & \new_[37975]_ ;
  assign \new_[37977]_  = \new_[37976]_  & \new_[37971]_ ;
  assign \new_[37981]_  = A234 & ~A233;
  assign \new_[37982]_  = A232 & \new_[37981]_ ;
  assign \new_[37986]_  = A266 & ~A265;
  assign \new_[37987]_  = A235 & \new_[37986]_ ;
  assign \new_[37988]_  = \new_[37987]_  & \new_[37982]_ ;
  assign \new_[37992]_  = A167 & ~A169;
  assign \new_[37993]_  = A170 & \new_[37992]_ ;
  assign \new_[37997]_  = ~A201 & ~A200;
  assign \new_[37998]_  = ~A166 & \new_[37997]_ ;
  assign \new_[37999]_  = \new_[37998]_  & \new_[37993]_ ;
  assign \new_[38003]_  = A234 & ~A233;
  assign \new_[38004]_  = A232 & \new_[38003]_ ;
  assign \new_[38008]_  = A299 & ~A298;
  assign \new_[38009]_  = A236 & \new_[38008]_ ;
  assign \new_[38010]_  = \new_[38009]_  & \new_[38004]_ ;
  assign \new_[38014]_  = A167 & ~A169;
  assign \new_[38015]_  = A170 & \new_[38014]_ ;
  assign \new_[38019]_  = ~A201 & ~A200;
  assign \new_[38020]_  = ~A166 & \new_[38019]_ ;
  assign \new_[38021]_  = \new_[38020]_  & \new_[38015]_ ;
  assign \new_[38025]_  = A234 & ~A233;
  assign \new_[38026]_  = A232 & \new_[38025]_ ;
  assign \new_[38030]_  = A266 & ~A265;
  assign \new_[38031]_  = A236 & \new_[38030]_ ;
  assign \new_[38032]_  = \new_[38031]_  & \new_[38026]_ ;
  assign \new_[38036]_  = A167 & ~A169;
  assign \new_[38037]_  = A170 & \new_[38036]_ ;
  assign \new_[38041]_  = ~A201 & ~A200;
  assign \new_[38042]_  = ~A166 & \new_[38041]_ ;
  assign \new_[38043]_  = \new_[38042]_  & \new_[38037]_ ;
  assign \new_[38047]_  = A265 & ~A233;
  assign \new_[38048]_  = ~A232 & \new_[38047]_ ;
  assign \new_[38052]_  = ~A300 & A298;
  assign \new_[38053]_  = A266 & \new_[38052]_ ;
  assign \new_[38054]_  = \new_[38053]_  & \new_[38048]_ ;
  assign \new_[38058]_  = A167 & ~A169;
  assign \new_[38059]_  = A170 & \new_[38058]_ ;
  assign \new_[38063]_  = ~A201 & ~A200;
  assign \new_[38064]_  = ~A166 & \new_[38063]_ ;
  assign \new_[38065]_  = \new_[38064]_  & \new_[38059]_ ;
  assign \new_[38069]_  = A265 & ~A233;
  assign \new_[38070]_  = ~A232 & \new_[38069]_ ;
  assign \new_[38074]_  = A299 & A298;
  assign \new_[38075]_  = A266 & \new_[38074]_ ;
  assign \new_[38076]_  = \new_[38075]_  & \new_[38070]_ ;
  assign \new_[38080]_  = A167 & ~A169;
  assign \new_[38081]_  = A170 & \new_[38080]_ ;
  assign \new_[38085]_  = ~A201 & ~A200;
  assign \new_[38086]_  = ~A166 & \new_[38085]_ ;
  assign \new_[38087]_  = \new_[38086]_  & \new_[38081]_ ;
  assign \new_[38091]_  = A265 & ~A233;
  assign \new_[38092]_  = ~A232 & \new_[38091]_ ;
  assign \new_[38096]_  = ~A299 & ~A298;
  assign \new_[38097]_  = A266 & \new_[38096]_ ;
  assign \new_[38098]_  = \new_[38097]_  & \new_[38092]_ ;
  assign \new_[38102]_  = A167 & ~A169;
  assign \new_[38103]_  = A170 & \new_[38102]_ ;
  assign \new_[38107]_  = ~A201 & ~A200;
  assign \new_[38108]_  = ~A166 & \new_[38107]_ ;
  assign \new_[38109]_  = \new_[38108]_  & \new_[38103]_ ;
  assign \new_[38113]_  = ~A266 & ~A233;
  assign \new_[38114]_  = ~A232 & \new_[38113]_ ;
  assign \new_[38118]_  = ~A300 & A298;
  assign \new_[38119]_  = ~A267 & \new_[38118]_ ;
  assign \new_[38120]_  = \new_[38119]_  & \new_[38114]_ ;
  assign \new_[38124]_  = A167 & ~A169;
  assign \new_[38125]_  = A170 & \new_[38124]_ ;
  assign \new_[38129]_  = ~A201 & ~A200;
  assign \new_[38130]_  = ~A166 & \new_[38129]_ ;
  assign \new_[38131]_  = \new_[38130]_  & \new_[38125]_ ;
  assign \new_[38135]_  = ~A266 & ~A233;
  assign \new_[38136]_  = ~A232 & \new_[38135]_ ;
  assign \new_[38140]_  = A299 & A298;
  assign \new_[38141]_  = ~A267 & \new_[38140]_ ;
  assign \new_[38142]_  = \new_[38141]_  & \new_[38136]_ ;
  assign \new_[38146]_  = A167 & ~A169;
  assign \new_[38147]_  = A170 & \new_[38146]_ ;
  assign \new_[38151]_  = ~A201 & ~A200;
  assign \new_[38152]_  = ~A166 & \new_[38151]_ ;
  assign \new_[38153]_  = \new_[38152]_  & \new_[38147]_ ;
  assign \new_[38157]_  = ~A266 & ~A233;
  assign \new_[38158]_  = ~A232 & \new_[38157]_ ;
  assign \new_[38162]_  = ~A299 & ~A298;
  assign \new_[38163]_  = ~A267 & \new_[38162]_ ;
  assign \new_[38164]_  = \new_[38163]_  & \new_[38158]_ ;
  assign \new_[38168]_  = A167 & ~A169;
  assign \new_[38169]_  = A170 & \new_[38168]_ ;
  assign \new_[38173]_  = ~A201 & ~A200;
  assign \new_[38174]_  = ~A166 & \new_[38173]_ ;
  assign \new_[38175]_  = \new_[38174]_  & \new_[38169]_ ;
  assign \new_[38179]_  = ~A265 & ~A233;
  assign \new_[38180]_  = ~A232 & \new_[38179]_ ;
  assign \new_[38184]_  = ~A300 & A298;
  assign \new_[38185]_  = ~A266 & \new_[38184]_ ;
  assign \new_[38186]_  = \new_[38185]_  & \new_[38180]_ ;
  assign \new_[38190]_  = A167 & ~A169;
  assign \new_[38191]_  = A170 & \new_[38190]_ ;
  assign \new_[38195]_  = ~A201 & ~A200;
  assign \new_[38196]_  = ~A166 & \new_[38195]_ ;
  assign \new_[38197]_  = \new_[38196]_  & \new_[38191]_ ;
  assign \new_[38201]_  = ~A265 & ~A233;
  assign \new_[38202]_  = ~A232 & \new_[38201]_ ;
  assign \new_[38206]_  = A299 & A298;
  assign \new_[38207]_  = ~A266 & \new_[38206]_ ;
  assign \new_[38208]_  = \new_[38207]_  & \new_[38202]_ ;
  assign \new_[38212]_  = A167 & ~A169;
  assign \new_[38213]_  = A170 & \new_[38212]_ ;
  assign \new_[38217]_  = ~A201 & ~A200;
  assign \new_[38218]_  = ~A166 & \new_[38217]_ ;
  assign \new_[38219]_  = \new_[38218]_  & \new_[38213]_ ;
  assign \new_[38223]_  = ~A265 & ~A233;
  assign \new_[38224]_  = ~A232 & \new_[38223]_ ;
  assign \new_[38228]_  = ~A299 & ~A298;
  assign \new_[38229]_  = ~A266 & \new_[38228]_ ;
  assign \new_[38230]_  = \new_[38229]_  & \new_[38224]_ ;
  assign \new_[38234]_  = A167 & ~A169;
  assign \new_[38235]_  = A170 & \new_[38234]_ ;
  assign \new_[38239]_  = ~A200 & ~A199;
  assign \new_[38240]_  = ~A166 & \new_[38239]_ ;
  assign \new_[38241]_  = \new_[38240]_  & \new_[38235]_ ;
  assign \new_[38245]_  = A265 & A233;
  assign \new_[38246]_  = A232 & \new_[38245]_ ;
  assign \new_[38250]_  = ~A300 & ~A299;
  assign \new_[38251]_  = ~A267 & \new_[38250]_ ;
  assign \new_[38252]_  = \new_[38251]_  & \new_[38246]_ ;
  assign \new_[38256]_  = A167 & ~A169;
  assign \new_[38257]_  = A170 & \new_[38256]_ ;
  assign \new_[38261]_  = ~A200 & ~A199;
  assign \new_[38262]_  = ~A166 & \new_[38261]_ ;
  assign \new_[38263]_  = \new_[38262]_  & \new_[38257]_ ;
  assign \new_[38267]_  = A265 & A233;
  assign \new_[38268]_  = A232 & \new_[38267]_ ;
  assign \new_[38272]_  = A299 & A298;
  assign \new_[38273]_  = ~A267 & \new_[38272]_ ;
  assign \new_[38274]_  = \new_[38273]_  & \new_[38268]_ ;
  assign \new_[38278]_  = A167 & ~A169;
  assign \new_[38279]_  = A170 & \new_[38278]_ ;
  assign \new_[38283]_  = ~A200 & ~A199;
  assign \new_[38284]_  = ~A166 & \new_[38283]_ ;
  assign \new_[38285]_  = \new_[38284]_  & \new_[38279]_ ;
  assign \new_[38289]_  = A265 & A233;
  assign \new_[38290]_  = A232 & \new_[38289]_ ;
  assign \new_[38294]_  = ~A299 & ~A298;
  assign \new_[38295]_  = ~A267 & \new_[38294]_ ;
  assign \new_[38296]_  = \new_[38295]_  & \new_[38290]_ ;
  assign \new_[38300]_  = A167 & ~A169;
  assign \new_[38301]_  = A170 & \new_[38300]_ ;
  assign \new_[38305]_  = ~A200 & ~A199;
  assign \new_[38306]_  = ~A166 & \new_[38305]_ ;
  assign \new_[38307]_  = \new_[38306]_  & \new_[38301]_ ;
  assign \new_[38311]_  = A265 & A233;
  assign \new_[38312]_  = A232 & \new_[38311]_ ;
  assign \new_[38316]_  = ~A300 & ~A299;
  assign \new_[38317]_  = A266 & \new_[38316]_ ;
  assign \new_[38318]_  = \new_[38317]_  & \new_[38312]_ ;
  assign \new_[38322]_  = A167 & ~A169;
  assign \new_[38323]_  = A170 & \new_[38322]_ ;
  assign \new_[38327]_  = ~A200 & ~A199;
  assign \new_[38328]_  = ~A166 & \new_[38327]_ ;
  assign \new_[38329]_  = \new_[38328]_  & \new_[38323]_ ;
  assign \new_[38333]_  = A265 & A233;
  assign \new_[38334]_  = A232 & \new_[38333]_ ;
  assign \new_[38338]_  = A299 & A298;
  assign \new_[38339]_  = A266 & \new_[38338]_ ;
  assign \new_[38340]_  = \new_[38339]_  & \new_[38334]_ ;
  assign \new_[38344]_  = A167 & ~A169;
  assign \new_[38345]_  = A170 & \new_[38344]_ ;
  assign \new_[38349]_  = ~A200 & ~A199;
  assign \new_[38350]_  = ~A166 & \new_[38349]_ ;
  assign \new_[38351]_  = \new_[38350]_  & \new_[38345]_ ;
  assign \new_[38355]_  = A265 & A233;
  assign \new_[38356]_  = A232 & \new_[38355]_ ;
  assign \new_[38360]_  = ~A299 & ~A298;
  assign \new_[38361]_  = A266 & \new_[38360]_ ;
  assign \new_[38362]_  = \new_[38361]_  & \new_[38356]_ ;
  assign \new_[38366]_  = A167 & ~A169;
  assign \new_[38367]_  = A170 & \new_[38366]_ ;
  assign \new_[38371]_  = ~A200 & ~A199;
  assign \new_[38372]_  = ~A166 & \new_[38371]_ ;
  assign \new_[38373]_  = \new_[38372]_  & \new_[38367]_ ;
  assign \new_[38377]_  = ~A265 & A233;
  assign \new_[38378]_  = A232 & \new_[38377]_ ;
  assign \new_[38382]_  = ~A300 & ~A299;
  assign \new_[38383]_  = ~A266 & \new_[38382]_ ;
  assign \new_[38384]_  = \new_[38383]_  & \new_[38378]_ ;
  assign \new_[38388]_  = A167 & ~A169;
  assign \new_[38389]_  = A170 & \new_[38388]_ ;
  assign \new_[38393]_  = ~A200 & ~A199;
  assign \new_[38394]_  = ~A166 & \new_[38393]_ ;
  assign \new_[38395]_  = \new_[38394]_  & \new_[38389]_ ;
  assign \new_[38399]_  = ~A265 & A233;
  assign \new_[38400]_  = A232 & \new_[38399]_ ;
  assign \new_[38404]_  = A299 & A298;
  assign \new_[38405]_  = ~A266 & \new_[38404]_ ;
  assign \new_[38406]_  = \new_[38405]_  & \new_[38400]_ ;
  assign \new_[38410]_  = A167 & ~A169;
  assign \new_[38411]_  = A170 & \new_[38410]_ ;
  assign \new_[38415]_  = ~A200 & ~A199;
  assign \new_[38416]_  = ~A166 & \new_[38415]_ ;
  assign \new_[38417]_  = \new_[38416]_  & \new_[38411]_ ;
  assign \new_[38421]_  = ~A265 & A233;
  assign \new_[38422]_  = A232 & \new_[38421]_ ;
  assign \new_[38426]_  = ~A299 & ~A298;
  assign \new_[38427]_  = ~A266 & \new_[38426]_ ;
  assign \new_[38428]_  = \new_[38427]_  & \new_[38422]_ ;
  assign \new_[38432]_  = A167 & ~A169;
  assign \new_[38433]_  = A170 & \new_[38432]_ ;
  assign \new_[38437]_  = ~A200 & ~A199;
  assign \new_[38438]_  = ~A166 & \new_[38437]_ ;
  assign \new_[38439]_  = \new_[38438]_  & \new_[38433]_ ;
  assign \new_[38443]_  = A298 & A233;
  assign \new_[38444]_  = ~A232 & \new_[38443]_ ;
  assign \new_[38448]_  = A301 & A300;
  assign \new_[38449]_  = ~A299 & \new_[38448]_ ;
  assign \new_[38450]_  = \new_[38449]_  & \new_[38444]_ ;
  assign \new_[38454]_  = A167 & ~A169;
  assign \new_[38455]_  = A170 & \new_[38454]_ ;
  assign \new_[38459]_  = ~A200 & ~A199;
  assign \new_[38460]_  = ~A166 & \new_[38459]_ ;
  assign \new_[38461]_  = \new_[38460]_  & \new_[38455]_ ;
  assign \new_[38465]_  = A298 & A233;
  assign \new_[38466]_  = ~A232 & \new_[38465]_ ;
  assign \new_[38470]_  = A302 & A300;
  assign \new_[38471]_  = ~A299 & \new_[38470]_ ;
  assign \new_[38472]_  = \new_[38471]_  & \new_[38466]_ ;
  assign \new_[38476]_  = A167 & ~A169;
  assign \new_[38477]_  = A170 & \new_[38476]_ ;
  assign \new_[38481]_  = ~A200 & ~A199;
  assign \new_[38482]_  = ~A166 & \new_[38481]_ ;
  assign \new_[38483]_  = \new_[38482]_  & \new_[38477]_ ;
  assign \new_[38487]_  = A265 & A233;
  assign \new_[38488]_  = ~A232 & \new_[38487]_ ;
  assign \new_[38492]_  = A268 & A267;
  assign \new_[38493]_  = ~A266 & \new_[38492]_ ;
  assign \new_[38494]_  = \new_[38493]_  & \new_[38488]_ ;
  assign \new_[38498]_  = A167 & ~A169;
  assign \new_[38499]_  = A170 & \new_[38498]_ ;
  assign \new_[38503]_  = ~A200 & ~A199;
  assign \new_[38504]_  = ~A166 & \new_[38503]_ ;
  assign \new_[38505]_  = \new_[38504]_  & \new_[38499]_ ;
  assign \new_[38509]_  = A265 & A233;
  assign \new_[38510]_  = ~A232 & \new_[38509]_ ;
  assign \new_[38514]_  = A269 & A267;
  assign \new_[38515]_  = ~A266 & \new_[38514]_ ;
  assign \new_[38516]_  = \new_[38515]_  & \new_[38510]_ ;
  assign \new_[38520]_  = A167 & ~A169;
  assign \new_[38521]_  = A170 & \new_[38520]_ ;
  assign \new_[38525]_  = ~A200 & ~A199;
  assign \new_[38526]_  = ~A166 & \new_[38525]_ ;
  assign \new_[38527]_  = \new_[38526]_  & \new_[38521]_ ;
  assign \new_[38531]_  = A265 & ~A234;
  assign \new_[38532]_  = ~A233 & \new_[38531]_ ;
  assign \new_[38536]_  = ~A300 & A298;
  assign \new_[38537]_  = A266 & \new_[38536]_ ;
  assign \new_[38538]_  = \new_[38537]_  & \new_[38532]_ ;
  assign \new_[38542]_  = A167 & ~A169;
  assign \new_[38543]_  = A170 & \new_[38542]_ ;
  assign \new_[38547]_  = ~A200 & ~A199;
  assign \new_[38548]_  = ~A166 & \new_[38547]_ ;
  assign \new_[38549]_  = \new_[38548]_  & \new_[38543]_ ;
  assign \new_[38553]_  = A265 & ~A234;
  assign \new_[38554]_  = ~A233 & \new_[38553]_ ;
  assign \new_[38558]_  = A299 & A298;
  assign \new_[38559]_  = A266 & \new_[38558]_ ;
  assign \new_[38560]_  = \new_[38559]_  & \new_[38554]_ ;
  assign \new_[38564]_  = A167 & ~A169;
  assign \new_[38565]_  = A170 & \new_[38564]_ ;
  assign \new_[38569]_  = ~A200 & ~A199;
  assign \new_[38570]_  = ~A166 & \new_[38569]_ ;
  assign \new_[38571]_  = \new_[38570]_  & \new_[38565]_ ;
  assign \new_[38575]_  = A265 & ~A234;
  assign \new_[38576]_  = ~A233 & \new_[38575]_ ;
  assign \new_[38580]_  = ~A299 & ~A298;
  assign \new_[38581]_  = A266 & \new_[38580]_ ;
  assign \new_[38582]_  = \new_[38581]_  & \new_[38576]_ ;
  assign \new_[38586]_  = A167 & ~A169;
  assign \new_[38587]_  = A170 & \new_[38586]_ ;
  assign \new_[38591]_  = ~A200 & ~A199;
  assign \new_[38592]_  = ~A166 & \new_[38591]_ ;
  assign \new_[38593]_  = \new_[38592]_  & \new_[38587]_ ;
  assign \new_[38597]_  = ~A266 & ~A234;
  assign \new_[38598]_  = ~A233 & \new_[38597]_ ;
  assign \new_[38602]_  = ~A300 & A298;
  assign \new_[38603]_  = ~A267 & \new_[38602]_ ;
  assign \new_[38604]_  = \new_[38603]_  & \new_[38598]_ ;
  assign \new_[38608]_  = A167 & ~A169;
  assign \new_[38609]_  = A170 & \new_[38608]_ ;
  assign \new_[38613]_  = ~A200 & ~A199;
  assign \new_[38614]_  = ~A166 & \new_[38613]_ ;
  assign \new_[38615]_  = \new_[38614]_  & \new_[38609]_ ;
  assign \new_[38619]_  = ~A266 & ~A234;
  assign \new_[38620]_  = ~A233 & \new_[38619]_ ;
  assign \new_[38624]_  = A299 & A298;
  assign \new_[38625]_  = ~A267 & \new_[38624]_ ;
  assign \new_[38626]_  = \new_[38625]_  & \new_[38620]_ ;
  assign \new_[38630]_  = A167 & ~A169;
  assign \new_[38631]_  = A170 & \new_[38630]_ ;
  assign \new_[38635]_  = ~A200 & ~A199;
  assign \new_[38636]_  = ~A166 & \new_[38635]_ ;
  assign \new_[38637]_  = \new_[38636]_  & \new_[38631]_ ;
  assign \new_[38641]_  = ~A266 & ~A234;
  assign \new_[38642]_  = ~A233 & \new_[38641]_ ;
  assign \new_[38646]_  = ~A299 & ~A298;
  assign \new_[38647]_  = ~A267 & \new_[38646]_ ;
  assign \new_[38648]_  = \new_[38647]_  & \new_[38642]_ ;
  assign \new_[38652]_  = A167 & ~A169;
  assign \new_[38653]_  = A170 & \new_[38652]_ ;
  assign \new_[38657]_  = ~A200 & ~A199;
  assign \new_[38658]_  = ~A166 & \new_[38657]_ ;
  assign \new_[38659]_  = \new_[38658]_  & \new_[38653]_ ;
  assign \new_[38663]_  = ~A265 & ~A234;
  assign \new_[38664]_  = ~A233 & \new_[38663]_ ;
  assign \new_[38668]_  = ~A300 & A298;
  assign \new_[38669]_  = ~A266 & \new_[38668]_ ;
  assign \new_[38670]_  = \new_[38669]_  & \new_[38664]_ ;
  assign \new_[38674]_  = A167 & ~A169;
  assign \new_[38675]_  = A170 & \new_[38674]_ ;
  assign \new_[38679]_  = ~A200 & ~A199;
  assign \new_[38680]_  = ~A166 & \new_[38679]_ ;
  assign \new_[38681]_  = \new_[38680]_  & \new_[38675]_ ;
  assign \new_[38685]_  = ~A265 & ~A234;
  assign \new_[38686]_  = ~A233 & \new_[38685]_ ;
  assign \new_[38690]_  = A299 & A298;
  assign \new_[38691]_  = ~A266 & \new_[38690]_ ;
  assign \new_[38692]_  = \new_[38691]_  & \new_[38686]_ ;
  assign \new_[38696]_  = A167 & ~A169;
  assign \new_[38697]_  = A170 & \new_[38696]_ ;
  assign \new_[38701]_  = ~A200 & ~A199;
  assign \new_[38702]_  = ~A166 & \new_[38701]_ ;
  assign \new_[38703]_  = \new_[38702]_  & \new_[38697]_ ;
  assign \new_[38707]_  = ~A265 & ~A234;
  assign \new_[38708]_  = ~A233 & \new_[38707]_ ;
  assign \new_[38712]_  = ~A299 & ~A298;
  assign \new_[38713]_  = ~A266 & \new_[38712]_ ;
  assign \new_[38714]_  = \new_[38713]_  & \new_[38708]_ ;
  assign \new_[38718]_  = A167 & ~A169;
  assign \new_[38719]_  = A170 & \new_[38718]_ ;
  assign \new_[38723]_  = ~A200 & ~A199;
  assign \new_[38724]_  = ~A166 & \new_[38723]_ ;
  assign \new_[38725]_  = \new_[38724]_  & \new_[38719]_ ;
  assign \new_[38729]_  = A234 & ~A233;
  assign \new_[38730]_  = A232 & \new_[38729]_ ;
  assign \new_[38734]_  = A299 & ~A298;
  assign \new_[38735]_  = A235 & \new_[38734]_ ;
  assign \new_[38736]_  = \new_[38735]_  & \new_[38730]_ ;
  assign \new_[38740]_  = A167 & ~A169;
  assign \new_[38741]_  = A170 & \new_[38740]_ ;
  assign \new_[38745]_  = ~A200 & ~A199;
  assign \new_[38746]_  = ~A166 & \new_[38745]_ ;
  assign \new_[38747]_  = \new_[38746]_  & \new_[38741]_ ;
  assign \new_[38751]_  = A234 & ~A233;
  assign \new_[38752]_  = A232 & \new_[38751]_ ;
  assign \new_[38756]_  = A266 & ~A265;
  assign \new_[38757]_  = A235 & \new_[38756]_ ;
  assign \new_[38758]_  = \new_[38757]_  & \new_[38752]_ ;
  assign \new_[38762]_  = A167 & ~A169;
  assign \new_[38763]_  = A170 & \new_[38762]_ ;
  assign \new_[38767]_  = ~A200 & ~A199;
  assign \new_[38768]_  = ~A166 & \new_[38767]_ ;
  assign \new_[38769]_  = \new_[38768]_  & \new_[38763]_ ;
  assign \new_[38773]_  = A234 & ~A233;
  assign \new_[38774]_  = A232 & \new_[38773]_ ;
  assign \new_[38778]_  = A299 & ~A298;
  assign \new_[38779]_  = A236 & \new_[38778]_ ;
  assign \new_[38780]_  = \new_[38779]_  & \new_[38774]_ ;
  assign \new_[38784]_  = A167 & ~A169;
  assign \new_[38785]_  = A170 & \new_[38784]_ ;
  assign \new_[38789]_  = ~A200 & ~A199;
  assign \new_[38790]_  = ~A166 & \new_[38789]_ ;
  assign \new_[38791]_  = \new_[38790]_  & \new_[38785]_ ;
  assign \new_[38795]_  = A234 & ~A233;
  assign \new_[38796]_  = A232 & \new_[38795]_ ;
  assign \new_[38800]_  = A266 & ~A265;
  assign \new_[38801]_  = A236 & \new_[38800]_ ;
  assign \new_[38802]_  = \new_[38801]_  & \new_[38796]_ ;
  assign \new_[38806]_  = A167 & ~A169;
  assign \new_[38807]_  = A170 & \new_[38806]_ ;
  assign \new_[38811]_  = ~A200 & ~A199;
  assign \new_[38812]_  = ~A166 & \new_[38811]_ ;
  assign \new_[38813]_  = \new_[38812]_  & \new_[38807]_ ;
  assign \new_[38817]_  = A265 & ~A233;
  assign \new_[38818]_  = ~A232 & \new_[38817]_ ;
  assign \new_[38822]_  = ~A300 & A298;
  assign \new_[38823]_  = A266 & \new_[38822]_ ;
  assign \new_[38824]_  = \new_[38823]_  & \new_[38818]_ ;
  assign \new_[38828]_  = A167 & ~A169;
  assign \new_[38829]_  = A170 & \new_[38828]_ ;
  assign \new_[38833]_  = ~A200 & ~A199;
  assign \new_[38834]_  = ~A166 & \new_[38833]_ ;
  assign \new_[38835]_  = \new_[38834]_  & \new_[38829]_ ;
  assign \new_[38839]_  = A265 & ~A233;
  assign \new_[38840]_  = ~A232 & \new_[38839]_ ;
  assign \new_[38844]_  = A299 & A298;
  assign \new_[38845]_  = A266 & \new_[38844]_ ;
  assign \new_[38846]_  = \new_[38845]_  & \new_[38840]_ ;
  assign \new_[38850]_  = A167 & ~A169;
  assign \new_[38851]_  = A170 & \new_[38850]_ ;
  assign \new_[38855]_  = ~A200 & ~A199;
  assign \new_[38856]_  = ~A166 & \new_[38855]_ ;
  assign \new_[38857]_  = \new_[38856]_  & \new_[38851]_ ;
  assign \new_[38861]_  = A265 & ~A233;
  assign \new_[38862]_  = ~A232 & \new_[38861]_ ;
  assign \new_[38866]_  = ~A299 & ~A298;
  assign \new_[38867]_  = A266 & \new_[38866]_ ;
  assign \new_[38868]_  = \new_[38867]_  & \new_[38862]_ ;
  assign \new_[38872]_  = A167 & ~A169;
  assign \new_[38873]_  = A170 & \new_[38872]_ ;
  assign \new_[38877]_  = ~A200 & ~A199;
  assign \new_[38878]_  = ~A166 & \new_[38877]_ ;
  assign \new_[38879]_  = \new_[38878]_  & \new_[38873]_ ;
  assign \new_[38883]_  = ~A266 & ~A233;
  assign \new_[38884]_  = ~A232 & \new_[38883]_ ;
  assign \new_[38888]_  = ~A300 & A298;
  assign \new_[38889]_  = ~A267 & \new_[38888]_ ;
  assign \new_[38890]_  = \new_[38889]_  & \new_[38884]_ ;
  assign \new_[38894]_  = A167 & ~A169;
  assign \new_[38895]_  = A170 & \new_[38894]_ ;
  assign \new_[38899]_  = ~A200 & ~A199;
  assign \new_[38900]_  = ~A166 & \new_[38899]_ ;
  assign \new_[38901]_  = \new_[38900]_  & \new_[38895]_ ;
  assign \new_[38905]_  = ~A266 & ~A233;
  assign \new_[38906]_  = ~A232 & \new_[38905]_ ;
  assign \new_[38910]_  = A299 & A298;
  assign \new_[38911]_  = ~A267 & \new_[38910]_ ;
  assign \new_[38912]_  = \new_[38911]_  & \new_[38906]_ ;
  assign \new_[38916]_  = A167 & ~A169;
  assign \new_[38917]_  = A170 & \new_[38916]_ ;
  assign \new_[38921]_  = ~A200 & ~A199;
  assign \new_[38922]_  = ~A166 & \new_[38921]_ ;
  assign \new_[38923]_  = \new_[38922]_  & \new_[38917]_ ;
  assign \new_[38927]_  = ~A266 & ~A233;
  assign \new_[38928]_  = ~A232 & \new_[38927]_ ;
  assign \new_[38932]_  = ~A299 & ~A298;
  assign \new_[38933]_  = ~A267 & \new_[38932]_ ;
  assign \new_[38934]_  = \new_[38933]_  & \new_[38928]_ ;
  assign \new_[38938]_  = A167 & ~A169;
  assign \new_[38939]_  = A170 & \new_[38938]_ ;
  assign \new_[38943]_  = ~A200 & ~A199;
  assign \new_[38944]_  = ~A166 & \new_[38943]_ ;
  assign \new_[38945]_  = \new_[38944]_  & \new_[38939]_ ;
  assign \new_[38949]_  = ~A265 & ~A233;
  assign \new_[38950]_  = ~A232 & \new_[38949]_ ;
  assign \new_[38954]_  = ~A300 & A298;
  assign \new_[38955]_  = ~A266 & \new_[38954]_ ;
  assign \new_[38956]_  = \new_[38955]_  & \new_[38950]_ ;
  assign \new_[38960]_  = A167 & ~A169;
  assign \new_[38961]_  = A170 & \new_[38960]_ ;
  assign \new_[38965]_  = ~A200 & ~A199;
  assign \new_[38966]_  = ~A166 & \new_[38965]_ ;
  assign \new_[38967]_  = \new_[38966]_  & \new_[38961]_ ;
  assign \new_[38971]_  = ~A265 & ~A233;
  assign \new_[38972]_  = ~A232 & \new_[38971]_ ;
  assign \new_[38976]_  = A299 & A298;
  assign \new_[38977]_  = ~A266 & \new_[38976]_ ;
  assign \new_[38978]_  = \new_[38977]_  & \new_[38972]_ ;
  assign \new_[38982]_  = A167 & ~A169;
  assign \new_[38983]_  = A170 & \new_[38982]_ ;
  assign \new_[38987]_  = ~A200 & ~A199;
  assign \new_[38988]_  = ~A166 & \new_[38987]_ ;
  assign \new_[38989]_  = \new_[38988]_  & \new_[38983]_ ;
  assign \new_[38993]_  = ~A265 & ~A233;
  assign \new_[38994]_  = ~A232 & \new_[38993]_ ;
  assign \new_[38998]_  = ~A299 & ~A298;
  assign \new_[38999]_  = ~A266 & \new_[38998]_ ;
  assign \new_[39000]_  = \new_[38999]_  & \new_[38994]_ ;
  assign \new_[39004]_  = ~A167 & ~A169;
  assign \new_[39005]_  = A170 & \new_[39004]_ ;
  assign \new_[39009]_  = A200 & A199;
  assign \new_[39010]_  = A166 & \new_[39009]_ ;
  assign \new_[39011]_  = \new_[39010]_  & \new_[39005]_ ;
  assign \new_[39015]_  = A265 & A233;
  assign \new_[39016]_  = A232 & \new_[39015]_ ;
  assign \new_[39020]_  = ~A300 & ~A299;
  assign \new_[39021]_  = ~A267 & \new_[39020]_ ;
  assign \new_[39022]_  = \new_[39021]_  & \new_[39016]_ ;
  assign \new_[39026]_  = ~A167 & ~A169;
  assign \new_[39027]_  = A170 & \new_[39026]_ ;
  assign \new_[39031]_  = A200 & A199;
  assign \new_[39032]_  = A166 & \new_[39031]_ ;
  assign \new_[39033]_  = \new_[39032]_  & \new_[39027]_ ;
  assign \new_[39037]_  = A265 & A233;
  assign \new_[39038]_  = A232 & \new_[39037]_ ;
  assign \new_[39042]_  = A299 & A298;
  assign \new_[39043]_  = ~A267 & \new_[39042]_ ;
  assign \new_[39044]_  = \new_[39043]_  & \new_[39038]_ ;
  assign \new_[39048]_  = ~A167 & ~A169;
  assign \new_[39049]_  = A170 & \new_[39048]_ ;
  assign \new_[39053]_  = A200 & A199;
  assign \new_[39054]_  = A166 & \new_[39053]_ ;
  assign \new_[39055]_  = \new_[39054]_  & \new_[39049]_ ;
  assign \new_[39059]_  = A265 & A233;
  assign \new_[39060]_  = A232 & \new_[39059]_ ;
  assign \new_[39064]_  = ~A299 & ~A298;
  assign \new_[39065]_  = ~A267 & \new_[39064]_ ;
  assign \new_[39066]_  = \new_[39065]_  & \new_[39060]_ ;
  assign \new_[39070]_  = ~A167 & ~A169;
  assign \new_[39071]_  = A170 & \new_[39070]_ ;
  assign \new_[39075]_  = A200 & A199;
  assign \new_[39076]_  = A166 & \new_[39075]_ ;
  assign \new_[39077]_  = \new_[39076]_  & \new_[39071]_ ;
  assign \new_[39081]_  = A265 & A233;
  assign \new_[39082]_  = A232 & \new_[39081]_ ;
  assign \new_[39086]_  = ~A300 & ~A299;
  assign \new_[39087]_  = A266 & \new_[39086]_ ;
  assign \new_[39088]_  = \new_[39087]_  & \new_[39082]_ ;
  assign \new_[39092]_  = ~A167 & ~A169;
  assign \new_[39093]_  = A170 & \new_[39092]_ ;
  assign \new_[39097]_  = A200 & A199;
  assign \new_[39098]_  = A166 & \new_[39097]_ ;
  assign \new_[39099]_  = \new_[39098]_  & \new_[39093]_ ;
  assign \new_[39103]_  = A265 & A233;
  assign \new_[39104]_  = A232 & \new_[39103]_ ;
  assign \new_[39108]_  = A299 & A298;
  assign \new_[39109]_  = A266 & \new_[39108]_ ;
  assign \new_[39110]_  = \new_[39109]_  & \new_[39104]_ ;
  assign \new_[39114]_  = ~A167 & ~A169;
  assign \new_[39115]_  = A170 & \new_[39114]_ ;
  assign \new_[39119]_  = A200 & A199;
  assign \new_[39120]_  = A166 & \new_[39119]_ ;
  assign \new_[39121]_  = \new_[39120]_  & \new_[39115]_ ;
  assign \new_[39125]_  = A265 & A233;
  assign \new_[39126]_  = A232 & \new_[39125]_ ;
  assign \new_[39130]_  = ~A299 & ~A298;
  assign \new_[39131]_  = A266 & \new_[39130]_ ;
  assign \new_[39132]_  = \new_[39131]_  & \new_[39126]_ ;
  assign \new_[39136]_  = ~A167 & ~A169;
  assign \new_[39137]_  = A170 & \new_[39136]_ ;
  assign \new_[39141]_  = A200 & A199;
  assign \new_[39142]_  = A166 & \new_[39141]_ ;
  assign \new_[39143]_  = \new_[39142]_  & \new_[39137]_ ;
  assign \new_[39147]_  = ~A265 & A233;
  assign \new_[39148]_  = A232 & \new_[39147]_ ;
  assign \new_[39152]_  = ~A300 & ~A299;
  assign \new_[39153]_  = ~A266 & \new_[39152]_ ;
  assign \new_[39154]_  = \new_[39153]_  & \new_[39148]_ ;
  assign \new_[39158]_  = ~A167 & ~A169;
  assign \new_[39159]_  = A170 & \new_[39158]_ ;
  assign \new_[39163]_  = A200 & A199;
  assign \new_[39164]_  = A166 & \new_[39163]_ ;
  assign \new_[39165]_  = \new_[39164]_  & \new_[39159]_ ;
  assign \new_[39169]_  = ~A265 & A233;
  assign \new_[39170]_  = A232 & \new_[39169]_ ;
  assign \new_[39174]_  = A299 & A298;
  assign \new_[39175]_  = ~A266 & \new_[39174]_ ;
  assign \new_[39176]_  = \new_[39175]_  & \new_[39170]_ ;
  assign \new_[39180]_  = ~A167 & ~A169;
  assign \new_[39181]_  = A170 & \new_[39180]_ ;
  assign \new_[39185]_  = A200 & A199;
  assign \new_[39186]_  = A166 & \new_[39185]_ ;
  assign \new_[39187]_  = \new_[39186]_  & \new_[39181]_ ;
  assign \new_[39191]_  = ~A265 & A233;
  assign \new_[39192]_  = A232 & \new_[39191]_ ;
  assign \new_[39196]_  = ~A299 & ~A298;
  assign \new_[39197]_  = ~A266 & \new_[39196]_ ;
  assign \new_[39198]_  = \new_[39197]_  & \new_[39192]_ ;
  assign \new_[39202]_  = ~A167 & ~A169;
  assign \new_[39203]_  = A170 & \new_[39202]_ ;
  assign \new_[39207]_  = A200 & A199;
  assign \new_[39208]_  = A166 & \new_[39207]_ ;
  assign \new_[39209]_  = \new_[39208]_  & \new_[39203]_ ;
  assign \new_[39213]_  = A298 & A233;
  assign \new_[39214]_  = ~A232 & \new_[39213]_ ;
  assign \new_[39218]_  = A301 & A300;
  assign \new_[39219]_  = ~A299 & \new_[39218]_ ;
  assign \new_[39220]_  = \new_[39219]_  & \new_[39214]_ ;
  assign \new_[39224]_  = ~A167 & ~A169;
  assign \new_[39225]_  = A170 & \new_[39224]_ ;
  assign \new_[39229]_  = A200 & A199;
  assign \new_[39230]_  = A166 & \new_[39229]_ ;
  assign \new_[39231]_  = \new_[39230]_  & \new_[39225]_ ;
  assign \new_[39235]_  = A298 & A233;
  assign \new_[39236]_  = ~A232 & \new_[39235]_ ;
  assign \new_[39240]_  = A302 & A300;
  assign \new_[39241]_  = ~A299 & \new_[39240]_ ;
  assign \new_[39242]_  = \new_[39241]_  & \new_[39236]_ ;
  assign \new_[39246]_  = ~A167 & ~A169;
  assign \new_[39247]_  = A170 & \new_[39246]_ ;
  assign \new_[39251]_  = A200 & A199;
  assign \new_[39252]_  = A166 & \new_[39251]_ ;
  assign \new_[39253]_  = \new_[39252]_  & \new_[39247]_ ;
  assign \new_[39257]_  = A265 & A233;
  assign \new_[39258]_  = ~A232 & \new_[39257]_ ;
  assign \new_[39262]_  = A268 & A267;
  assign \new_[39263]_  = ~A266 & \new_[39262]_ ;
  assign \new_[39264]_  = \new_[39263]_  & \new_[39258]_ ;
  assign \new_[39268]_  = ~A167 & ~A169;
  assign \new_[39269]_  = A170 & \new_[39268]_ ;
  assign \new_[39273]_  = A200 & A199;
  assign \new_[39274]_  = A166 & \new_[39273]_ ;
  assign \new_[39275]_  = \new_[39274]_  & \new_[39269]_ ;
  assign \new_[39279]_  = A265 & A233;
  assign \new_[39280]_  = ~A232 & \new_[39279]_ ;
  assign \new_[39284]_  = A269 & A267;
  assign \new_[39285]_  = ~A266 & \new_[39284]_ ;
  assign \new_[39286]_  = \new_[39285]_  & \new_[39280]_ ;
  assign \new_[39290]_  = ~A167 & ~A169;
  assign \new_[39291]_  = A170 & \new_[39290]_ ;
  assign \new_[39295]_  = A200 & A199;
  assign \new_[39296]_  = A166 & \new_[39295]_ ;
  assign \new_[39297]_  = \new_[39296]_  & \new_[39291]_ ;
  assign \new_[39301]_  = A265 & ~A234;
  assign \new_[39302]_  = ~A233 & \new_[39301]_ ;
  assign \new_[39306]_  = ~A300 & A298;
  assign \new_[39307]_  = A266 & \new_[39306]_ ;
  assign \new_[39308]_  = \new_[39307]_  & \new_[39302]_ ;
  assign \new_[39312]_  = ~A167 & ~A169;
  assign \new_[39313]_  = A170 & \new_[39312]_ ;
  assign \new_[39317]_  = A200 & A199;
  assign \new_[39318]_  = A166 & \new_[39317]_ ;
  assign \new_[39319]_  = \new_[39318]_  & \new_[39313]_ ;
  assign \new_[39323]_  = A265 & ~A234;
  assign \new_[39324]_  = ~A233 & \new_[39323]_ ;
  assign \new_[39328]_  = A299 & A298;
  assign \new_[39329]_  = A266 & \new_[39328]_ ;
  assign \new_[39330]_  = \new_[39329]_  & \new_[39324]_ ;
  assign \new_[39334]_  = ~A167 & ~A169;
  assign \new_[39335]_  = A170 & \new_[39334]_ ;
  assign \new_[39339]_  = A200 & A199;
  assign \new_[39340]_  = A166 & \new_[39339]_ ;
  assign \new_[39341]_  = \new_[39340]_  & \new_[39335]_ ;
  assign \new_[39345]_  = A265 & ~A234;
  assign \new_[39346]_  = ~A233 & \new_[39345]_ ;
  assign \new_[39350]_  = ~A299 & ~A298;
  assign \new_[39351]_  = A266 & \new_[39350]_ ;
  assign \new_[39352]_  = \new_[39351]_  & \new_[39346]_ ;
  assign \new_[39356]_  = ~A167 & ~A169;
  assign \new_[39357]_  = A170 & \new_[39356]_ ;
  assign \new_[39361]_  = A200 & A199;
  assign \new_[39362]_  = A166 & \new_[39361]_ ;
  assign \new_[39363]_  = \new_[39362]_  & \new_[39357]_ ;
  assign \new_[39367]_  = ~A266 & ~A234;
  assign \new_[39368]_  = ~A233 & \new_[39367]_ ;
  assign \new_[39372]_  = ~A300 & A298;
  assign \new_[39373]_  = ~A267 & \new_[39372]_ ;
  assign \new_[39374]_  = \new_[39373]_  & \new_[39368]_ ;
  assign \new_[39378]_  = ~A167 & ~A169;
  assign \new_[39379]_  = A170 & \new_[39378]_ ;
  assign \new_[39383]_  = A200 & A199;
  assign \new_[39384]_  = A166 & \new_[39383]_ ;
  assign \new_[39385]_  = \new_[39384]_  & \new_[39379]_ ;
  assign \new_[39389]_  = ~A266 & ~A234;
  assign \new_[39390]_  = ~A233 & \new_[39389]_ ;
  assign \new_[39394]_  = A299 & A298;
  assign \new_[39395]_  = ~A267 & \new_[39394]_ ;
  assign \new_[39396]_  = \new_[39395]_  & \new_[39390]_ ;
  assign \new_[39400]_  = ~A167 & ~A169;
  assign \new_[39401]_  = A170 & \new_[39400]_ ;
  assign \new_[39405]_  = A200 & A199;
  assign \new_[39406]_  = A166 & \new_[39405]_ ;
  assign \new_[39407]_  = \new_[39406]_  & \new_[39401]_ ;
  assign \new_[39411]_  = ~A266 & ~A234;
  assign \new_[39412]_  = ~A233 & \new_[39411]_ ;
  assign \new_[39416]_  = ~A299 & ~A298;
  assign \new_[39417]_  = ~A267 & \new_[39416]_ ;
  assign \new_[39418]_  = \new_[39417]_  & \new_[39412]_ ;
  assign \new_[39422]_  = ~A167 & ~A169;
  assign \new_[39423]_  = A170 & \new_[39422]_ ;
  assign \new_[39427]_  = A200 & A199;
  assign \new_[39428]_  = A166 & \new_[39427]_ ;
  assign \new_[39429]_  = \new_[39428]_  & \new_[39423]_ ;
  assign \new_[39433]_  = ~A265 & ~A234;
  assign \new_[39434]_  = ~A233 & \new_[39433]_ ;
  assign \new_[39438]_  = ~A300 & A298;
  assign \new_[39439]_  = ~A266 & \new_[39438]_ ;
  assign \new_[39440]_  = \new_[39439]_  & \new_[39434]_ ;
  assign \new_[39444]_  = ~A167 & ~A169;
  assign \new_[39445]_  = A170 & \new_[39444]_ ;
  assign \new_[39449]_  = A200 & A199;
  assign \new_[39450]_  = A166 & \new_[39449]_ ;
  assign \new_[39451]_  = \new_[39450]_  & \new_[39445]_ ;
  assign \new_[39455]_  = ~A265 & ~A234;
  assign \new_[39456]_  = ~A233 & \new_[39455]_ ;
  assign \new_[39460]_  = A299 & A298;
  assign \new_[39461]_  = ~A266 & \new_[39460]_ ;
  assign \new_[39462]_  = \new_[39461]_  & \new_[39456]_ ;
  assign \new_[39466]_  = ~A167 & ~A169;
  assign \new_[39467]_  = A170 & \new_[39466]_ ;
  assign \new_[39471]_  = A200 & A199;
  assign \new_[39472]_  = A166 & \new_[39471]_ ;
  assign \new_[39473]_  = \new_[39472]_  & \new_[39467]_ ;
  assign \new_[39477]_  = ~A265 & ~A234;
  assign \new_[39478]_  = ~A233 & \new_[39477]_ ;
  assign \new_[39482]_  = ~A299 & ~A298;
  assign \new_[39483]_  = ~A266 & \new_[39482]_ ;
  assign \new_[39484]_  = \new_[39483]_  & \new_[39478]_ ;
  assign \new_[39488]_  = ~A167 & ~A169;
  assign \new_[39489]_  = A170 & \new_[39488]_ ;
  assign \new_[39493]_  = A200 & A199;
  assign \new_[39494]_  = A166 & \new_[39493]_ ;
  assign \new_[39495]_  = \new_[39494]_  & \new_[39489]_ ;
  assign \new_[39499]_  = A234 & ~A233;
  assign \new_[39500]_  = A232 & \new_[39499]_ ;
  assign \new_[39504]_  = A299 & ~A298;
  assign \new_[39505]_  = A235 & \new_[39504]_ ;
  assign \new_[39506]_  = \new_[39505]_  & \new_[39500]_ ;
  assign \new_[39510]_  = ~A167 & ~A169;
  assign \new_[39511]_  = A170 & \new_[39510]_ ;
  assign \new_[39515]_  = A200 & A199;
  assign \new_[39516]_  = A166 & \new_[39515]_ ;
  assign \new_[39517]_  = \new_[39516]_  & \new_[39511]_ ;
  assign \new_[39521]_  = A234 & ~A233;
  assign \new_[39522]_  = A232 & \new_[39521]_ ;
  assign \new_[39526]_  = A266 & ~A265;
  assign \new_[39527]_  = A235 & \new_[39526]_ ;
  assign \new_[39528]_  = \new_[39527]_  & \new_[39522]_ ;
  assign \new_[39532]_  = ~A167 & ~A169;
  assign \new_[39533]_  = A170 & \new_[39532]_ ;
  assign \new_[39537]_  = A200 & A199;
  assign \new_[39538]_  = A166 & \new_[39537]_ ;
  assign \new_[39539]_  = \new_[39538]_  & \new_[39533]_ ;
  assign \new_[39543]_  = A234 & ~A233;
  assign \new_[39544]_  = A232 & \new_[39543]_ ;
  assign \new_[39548]_  = A299 & ~A298;
  assign \new_[39549]_  = A236 & \new_[39548]_ ;
  assign \new_[39550]_  = \new_[39549]_  & \new_[39544]_ ;
  assign \new_[39554]_  = ~A167 & ~A169;
  assign \new_[39555]_  = A170 & \new_[39554]_ ;
  assign \new_[39559]_  = A200 & A199;
  assign \new_[39560]_  = A166 & \new_[39559]_ ;
  assign \new_[39561]_  = \new_[39560]_  & \new_[39555]_ ;
  assign \new_[39565]_  = A234 & ~A233;
  assign \new_[39566]_  = A232 & \new_[39565]_ ;
  assign \new_[39570]_  = A266 & ~A265;
  assign \new_[39571]_  = A236 & \new_[39570]_ ;
  assign \new_[39572]_  = \new_[39571]_  & \new_[39566]_ ;
  assign \new_[39576]_  = ~A167 & ~A169;
  assign \new_[39577]_  = A170 & \new_[39576]_ ;
  assign \new_[39581]_  = A200 & A199;
  assign \new_[39582]_  = A166 & \new_[39581]_ ;
  assign \new_[39583]_  = \new_[39582]_  & \new_[39577]_ ;
  assign \new_[39587]_  = A265 & ~A233;
  assign \new_[39588]_  = ~A232 & \new_[39587]_ ;
  assign \new_[39592]_  = ~A300 & A298;
  assign \new_[39593]_  = A266 & \new_[39592]_ ;
  assign \new_[39594]_  = \new_[39593]_  & \new_[39588]_ ;
  assign \new_[39598]_  = ~A167 & ~A169;
  assign \new_[39599]_  = A170 & \new_[39598]_ ;
  assign \new_[39603]_  = A200 & A199;
  assign \new_[39604]_  = A166 & \new_[39603]_ ;
  assign \new_[39605]_  = \new_[39604]_  & \new_[39599]_ ;
  assign \new_[39609]_  = A265 & ~A233;
  assign \new_[39610]_  = ~A232 & \new_[39609]_ ;
  assign \new_[39614]_  = A299 & A298;
  assign \new_[39615]_  = A266 & \new_[39614]_ ;
  assign \new_[39616]_  = \new_[39615]_  & \new_[39610]_ ;
  assign \new_[39620]_  = ~A167 & ~A169;
  assign \new_[39621]_  = A170 & \new_[39620]_ ;
  assign \new_[39625]_  = A200 & A199;
  assign \new_[39626]_  = A166 & \new_[39625]_ ;
  assign \new_[39627]_  = \new_[39626]_  & \new_[39621]_ ;
  assign \new_[39631]_  = A265 & ~A233;
  assign \new_[39632]_  = ~A232 & \new_[39631]_ ;
  assign \new_[39636]_  = ~A299 & ~A298;
  assign \new_[39637]_  = A266 & \new_[39636]_ ;
  assign \new_[39638]_  = \new_[39637]_  & \new_[39632]_ ;
  assign \new_[39642]_  = ~A167 & ~A169;
  assign \new_[39643]_  = A170 & \new_[39642]_ ;
  assign \new_[39647]_  = A200 & A199;
  assign \new_[39648]_  = A166 & \new_[39647]_ ;
  assign \new_[39649]_  = \new_[39648]_  & \new_[39643]_ ;
  assign \new_[39653]_  = ~A266 & ~A233;
  assign \new_[39654]_  = ~A232 & \new_[39653]_ ;
  assign \new_[39658]_  = ~A300 & A298;
  assign \new_[39659]_  = ~A267 & \new_[39658]_ ;
  assign \new_[39660]_  = \new_[39659]_  & \new_[39654]_ ;
  assign \new_[39664]_  = ~A167 & ~A169;
  assign \new_[39665]_  = A170 & \new_[39664]_ ;
  assign \new_[39669]_  = A200 & A199;
  assign \new_[39670]_  = A166 & \new_[39669]_ ;
  assign \new_[39671]_  = \new_[39670]_  & \new_[39665]_ ;
  assign \new_[39675]_  = ~A266 & ~A233;
  assign \new_[39676]_  = ~A232 & \new_[39675]_ ;
  assign \new_[39680]_  = A299 & A298;
  assign \new_[39681]_  = ~A267 & \new_[39680]_ ;
  assign \new_[39682]_  = \new_[39681]_  & \new_[39676]_ ;
  assign \new_[39686]_  = ~A167 & ~A169;
  assign \new_[39687]_  = A170 & \new_[39686]_ ;
  assign \new_[39691]_  = A200 & A199;
  assign \new_[39692]_  = A166 & \new_[39691]_ ;
  assign \new_[39693]_  = \new_[39692]_  & \new_[39687]_ ;
  assign \new_[39697]_  = ~A266 & ~A233;
  assign \new_[39698]_  = ~A232 & \new_[39697]_ ;
  assign \new_[39702]_  = ~A299 & ~A298;
  assign \new_[39703]_  = ~A267 & \new_[39702]_ ;
  assign \new_[39704]_  = \new_[39703]_  & \new_[39698]_ ;
  assign \new_[39708]_  = ~A167 & ~A169;
  assign \new_[39709]_  = A170 & \new_[39708]_ ;
  assign \new_[39713]_  = A200 & A199;
  assign \new_[39714]_  = A166 & \new_[39713]_ ;
  assign \new_[39715]_  = \new_[39714]_  & \new_[39709]_ ;
  assign \new_[39719]_  = ~A265 & ~A233;
  assign \new_[39720]_  = ~A232 & \new_[39719]_ ;
  assign \new_[39724]_  = ~A300 & A298;
  assign \new_[39725]_  = ~A266 & \new_[39724]_ ;
  assign \new_[39726]_  = \new_[39725]_  & \new_[39720]_ ;
  assign \new_[39730]_  = ~A167 & ~A169;
  assign \new_[39731]_  = A170 & \new_[39730]_ ;
  assign \new_[39735]_  = A200 & A199;
  assign \new_[39736]_  = A166 & \new_[39735]_ ;
  assign \new_[39737]_  = \new_[39736]_  & \new_[39731]_ ;
  assign \new_[39741]_  = ~A265 & ~A233;
  assign \new_[39742]_  = ~A232 & \new_[39741]_ ;
  assign \new_[39746]_  = A299 & A298;
  assign \new_[39747]_  = ~A266 & \new_[39746]_ ;
  assign \new_[39748]_  = \new_[39747]_  & \new_[39742]_ ;
  assign \new_[39752]_  = ~A167 & ~A169;
  assign \new_[39753]_  = A170 & \new_[39752]_ ;
  assign \new_[39757]_  = A200 & A199;
  assign \new_[39758]_  = A166 & \new_[39757]_ ;
  assign \new_[39759]_  = \new_[39758]_  & \new_[39753]_ ;
  assign \new_[39763]_  = ~A265 & ~A233;
  assign \new_[39764]_  = ~A232 & \new_[39763]_ ;
  assign \new_[39768]_  = ~A299 & ~A298;
  assign \new_[39769]_  = ~A266 & \new_[39768]_ ;
  assign \new_[39770]_  = \new_[39769]_  & \new_[39764]_ ;
  assign \new_[39774]_  = ~A167 & ~A169;
  assign \new_[39775]_  = A170 & \new_[39774]_ ;
  assign \new_[39779]_  = ~A201 & ~A200;
  assign \new_[39780]_  = A166 & \new_[39779]_ ;
  assign \new_[39781]_  = \new_[39780]_  & \new_[39775]_ ;
  assign \new_[39785]_  = A265 & A233;
  assign \new_[39786]_  = A232 & \new_[39785]_ ;
  assign \new_[39790]_  = ~A300 & ~A299;
  assign \new_[39791]_  = ~A267 & \new_[39790]_ ;
  assign \new_[39792]_  = \new_[39791]_  & \new_[39786]_ ;
  assign \new_[39796]_  = ~A167 & ~A169;
  assign \new_[39797]_  = A170 & \new_[39796]_ ;
  assign \new_[39801]_  = ~A201 & ~A200;
  assign \new_[39802]_  = A166 & \new_[39801]_ ;
  assign \new_[39803]_  = \new_[39802]_  & \new_[39797]_ ;
  assign \new_[39807]_  = A265 & A233;
  assign \new_[39808]_  = A232 & \new_[39807]_ ;
  assign \new_[39812]_  = A299 & A298;
  assign \new_[39813]_  = ~A267 & \new_[39812]_ ;
  assign \new_[39814]_  = \new_[39813]_  & \new_[39808]_ ;
  assign \new_[39818]_  = ~A167 & ~A169;
  assign \new_[39819]_  = A170 & \new_[39818]_ ;
  assign \new_[39823]_  = ~A201 & ~A200;
  assign \new_[39824]_  = A166 & \new_[39823]_ ;
  assign \new_[39825]_  = \new_[39824]_  & \new_[39819]_ ;
  assign \new_[39829]_  = A265 & A233;
  assign \new_[39830]_  = A232 & \new_[39829]_ ;
  assign \new_[39834]_  = ~A299 & ~A298;
  assign \new_[39835]_  = ~A267 & \new_[39834]_ ;
  assign \new_[39836]_  = \new_[39835]_  & \new_[39830]_ ;
  assign \new_[39840]_  = ~A167 & ~A169;
  assign \new_[39841]_  = A170 & \new_[39840]_ ;
  assign \new_[39845]_  = ~A201 & ~A200;
  assign \new_[39846]_  = A166 & \new_[39845]_ ;
  assign \new_[39847]_  = \new_[39846]_  & \new_[39841]_ ;
  assign \new_[39851]_  = A265 & A233;
  assign \new_[39852]_  = A232 & \new_[39851]_ ;
  assign \new_[39856]_  = ~A300 & ~A299;
  assign \new_[39857]_  = A266 & \new_[39856]_ ;
  assign \new_[39858]_  = \new_[39857]_  & \new_[39852]_ ;
  assign \new_[39862]_  = ~A167 & ~A169;
  assign \new_[39863]_  = A170 & \new_[39862]_ ;
  assign \new_[39867]_  = ~A201 & ~A200;
  assign \new_[39868]_  = A166 & \new_[39867]_ ;
  assign \new_[39869]_  = \new_[39868]_  & \new_[39863]_ ;
  assign \new_[39873]_  = A265 & A233;
  assign \new_[39874]_  = A232 & \new_[39873]_ ;
  assign \new_[39878]_  = A299 & A298;
  assign \new_[39879]_  = A266 & \new_[39878]_ ;
  assign \new_[39880]_  = \new_[39879]_  & \new_[39874]_ ;
  assign \new_[39884]_  = ~A167 & ~A169;
  assign \new_[39885]_  = A170 & \new_[39884]_ ;
  assign \new_[39889]_  = ~A201 & ~A200;
  assign \new_[39890]_  = A166 & \new_[39889]_ ;
  assign \new_[39891]_  = \new_[39890]_  & \new_[39885]_ ;
  assign \new_[39895]_  = A265 & A233;
  assign \new_[39896]_  = A232 & \new_[39895]_ ;
  assign \new_[39900]_  = ~A299 & ~A298;
  assign \new_[39901]_  = A266 & \new_[39900]_ ;
  assign \new_[39902]_  = \new_[39901]_  & \new_[39896]_ ;
  assign \new_[39906]_  = ~A167 & ~A169;
  assign \new_[39907]_  = A170 & \new_[39906]_ ;
  assign \new_[39911]_  = ~A201 & ~A200;
  assign \new_[39912]_  = A166 & \new_[39911]_ ;
  assign \new_[39913]_  = \new_[39912]_  & \new_[39907]_ ;
  assign \new_[39917]_  = ~A265 & A233;
  assign \new_[39918]_  = A232 & \new_[39917]_ ;
  assign \new_[39922]_  = ~A300 & ~A299;
  assign \new_[39923]_  = ~A266 & \new_[39922]_ ;
  assign \new_[39924]_  = \new_[39923]_  & \new_[39918]_ ;
  assign \new_[39928]_  = ~A167 & ~A169;
  assign \new_[39929]_  = A170 & \new_[39928]_ ;
  assign \new_[39933]_  = ~A201 & ~A200;
  assign \new_[39934]_  = A166 & \new_[39933]_ ;
  assign \new_[39935]_  = \new_[39934]_  & \new_[39929]_ ;
  assign \new_[39939]_  = ~A265 & A233;
  assign \new_[39940]_  = A232 & \new_[39939]_ ;
  assign \new_[39944]_  = A299 & A298;
  assign \new_[39945]_  = ~A266 & \new_[39944]_ ;
  assign \new_[39946]_  = \new_[39945]_  & \new_[39940]_ ;
  assign \new_[39950]_  = ~A167 & ~A169;
  assign \new_[39951]_  = A170 & \new_[39950]_ ;
  assign \new_[39955]_  = ~A201 & ~A200;
  assign \new_[39956]_  = A166 & \new_[39955]_ ;
  assign \new_[39957]_  = \new_[39956]_  & \new_[39951]_ ;
  assign \new_[39961]_  = ~A265 & A233;
  assign \new_[39962]_  = A232 & \new_[39961]_ ;
  assign \new_[39966]_  = ~A299 & ~A298;
  assign \new_[39967]_  = ~A266 & \new_[39966]_ ;
  assign \new_[39968]_  = \new_[39967]_  & \new_[39962]_ ;
  assign \new_[39972]_  = ~A167 & ~A169;
  assign \new_[39973]_  = A170 & \new_[39972]_ ;
  assign \new_[39977]_  = ~A201 & ~A200;
  assign \new_[39978]_  = A166 & \new_[39977]_ ;
  assign \new_[39979]_  = \new_[39978]_  & \new_[39973]_ ;
  assign \new_[39983]_  = A298 & A233;
  assign \new_[39984]_  = ~A232 & \new_[39983]_ ;
  assign \new_[39988]_  = A301 & A300;
  assign \new_[39989]_  = ~A299 & \new_[39988]_ ;
  assign \new_[39990]_  = \new_[39989]_  & \new_[39984]_ ;
  assign \new_[39994]_  = ~A167 & ~A169;
  assign \new_[39995]_  = A170 & \new_[39994]_ ;
  assign \new_[39999]_  = ~A201 & ~A200;
  assign \new_[40000]_  = A166 & \new_[39999]_ ;
  assign \new_[40001]_  = \new_[40000]_  & \new_[39995]_ ;
  assign \new_[40005]_  = A298 & A233;
  assign \new_[40006]_  = ~A232 & \new_[40005]_ ;
  assign \new_[40010]_  = A302 & A300;
  assign \new_[40011]_  = ~A299 & \new_[40010]_ ;
  assign \new_[40012]_  = \new_[40011]_  & \new_[40006]_ ;
  assign \new_[40016]_  = ~A167 & ~A169;
  assign \new_[40017]_  = A170 & \new_[40016]_ ;
  assign \new_[40021]_  = ~A201 & ~A200;
  assign \new_[40022]_  = A166 & \new_[40021]_ ;
  assign \new_[40023]_  = \new_[40022]_  & \new_[40017]_ ;
  assign \new_[40027]_  = A265 & A233;
  assign \new_[40028]_  = ~A232 & \new_[40027]_ ;
  assign \new_[40032]_  = A268 & A267;
  assign \new_[40033]_  = ~A266 & \new_[40032]_ ;
  assign \new_[40034]_  = \new_[40033]_  & \new_[40028]_ ;
  assign \new_[40038]_  = ~A167 & ~A169;
  assign \new_[40039]_  = A170 & \new_[40038]_ ;
  assign \new_[40043]_  = ~A201 & ~A200;
  assign \new_[40044]_  = A166 & \new_[40043]_ ;
  assign \new_[40045]_  = \new_[40044]_  & \new_[40039]_ ;
  assign \new_[40049]_  = A265 & A233;
  assign \new_[40050]_  = ~A232 & \new_[40049]_ ;
  assign \new_[40054]_  = A269 & A267;
  assign \new_[40055]_  = ~A266 & \new_[40054]_ ;
  assign \new_[40056]_  = \new_[40055]_  & \new_[40050]_ ;
  assign \new_[40060]_  = ~A167 & ~A169;
  assign \new_[40061]_  = A170 & \new_[40060]_ ;
  assign \new_[40065]_  = ~A201 & ~A200;
  assign \new_[40066]_  = A166 & \new_[40065]_ ;
  assign \new_[40067]_  = \new_[40066]_  & \new_[40061]_ ;
  assign \new_[40071]_  = A265 & ~A234;
  assign \new_[40072]_  = ~A233 & \new_[40071]_ ;
  assign \new_[40076]_  = ~A300 & A298;
  assign \new_[40077]_  = A266 & \new_[40076]_ ;
  assign \new_[40078]_  = \new_[40077]_  & \new_[40072]_ ;
  assign \new_[40082]_  = ~A167 & ~A169;
  assign \new_[40083]_  = A170 & \new_[40082]_ ;
  assign \new_[40087]_  = ~A201 & ~A200;
  assign \new_[40088]_  = A166 & \new_[40087]_ ;
  assign \new_[40089]_  = \new_[40088]_  & \new_[40083]_ ;
  assign \new_[40093]_  = A265 & ~A234;
  assign \new_[40094]_  = ~A233 & \new_[40093]_ ;
  assign \new_[40098]_  = A299 & A298;
  assign \new_[40099]_  = A266 & \new_[40098]_ ;
  assign \new_[40100]_  = \new_[40099]_  & \new_[40094]_ ;
  assign \new_[40104]_  = ~A167 & ~A169;
  assign \new_[40105]_  = A170 & \new_[40104]_ ;
  assign \new_[40109]_  = ~A201 & ~A200;
  assign \new_[40110]_  = A166 & \new_[40109]_ ;
  assign \new_[40111]_  = \new_[40110]_  & \new_[40105]_ ;
  assign \new_[40115]_  = A265 & ~A234;
  assign \new_[40116]_  = ~A233 & \new_[40115]_ ;
  assign \new_[40120]_  = ~A299 & ~A298;
  assign \new_[40121]_  = A266 & \new_[40120]_ ;
  assign \new_[40122]_  = \new_[40121]_  & \new_[40116]_ ;
  assign \new_[40126]_  = ~A167 & ~A169;
  assign \new_[40127]_  = A170 & \new_[40126]_ ;
  assign \new_[40131]_  = ~A201 & ~A200;
  assign \new_[40132]_  = A166 & \new_[40131]_ ;
  assign \new_[40133]_  = \new_[40132]_  & \new_[40127]_ ;
  assign \new_[40137]_  = ~A266 & ~A234;
  assign \new_[40138]_  = ~A233 & \new_[40137]_ ;
  assign \new_[40142]_  = ~A300 & A298;
  assign \new_[40143]_  = ~A267 & \new_[40142]_ ;
  assign \new_[40144]_  = \new_[40143]_  & \new_[40138]_ ;
  assign \new_[40148]_  = ~A167 & ~A169;
  assign \new_[40149]_  = A170 & \new_[40148]_ ;
  assign \new_[40153]_  = ~A201 & ~A200;
  assign \new_[40154]_  = A166 & \new_[40153]_ ;
  assign \new_[40155]_  = \new_[40154]_  & \new_[40149]_ ;
  assign \new_[40159]_  = ~A266 & ~A234;
  assign \new_[40160]_  = ~A233 & \new_[40159]_ ;
  assign \new_[40164]_  = A299 & A298;
  assign \new_[40165]_  = ~A267 & \new_[40164]_ ;
  assign \new_[40166]_  = \new_[40165]_  & \new_[40160]_ ;
  assign \new_[40170]_  = ~A167 & ~A169;
  assign \new_[40171]_  = A170 & \new_[40170]_ ;
  assign \new_[40175]_  = ~A201 & ~A200;
  assign \new_[40176]_  = A166 & \new_[40175]_ ;
  assign \new_[40177]_  = \new_[40176]_  & \new_[40171]_ ;
  assign \new_[40181]_  = ~A266 & ~A234;
  assign \new_[40182]_  = ~A233 & \new_[40181]_ ;
  assign \new_[40186]_  = ~A299 & ~A298;
  assign \new_[40187]_  = ~A267 & \new_[40186]_ ;
  assign \new_[40188]_  = \new_[40187]_  & \new_[40182]_ ;
  assign \new_[40192]_  = ~A167 & ~A169;
  assign \new_[40193]_  = A170 & \new_[40192]_ ;
  assign \new_[40197]_  = ~A201 & ~A200;
  assign \new_[40198]_  = A166 & \new_[40197]_ ;
  assign \new_[40199]_  = \new_[40198]_  & \new_[40193]_ ;
  assign \new_[40203]_  = ~A265 & ~A234;
  assign \new_[40204]_  = ~A233 & \new_[40203]_ ;
  assign \new_[40208]_  = ~A300 & A298;
  assign \new_[40209]_  = ~A266 & \new_[40208]_ ;
  assign \new_[40210]_  = \new_[40209]_  & \new_[40204]_ ;
  assign \new_[40214]_  = ~A167 & ~A169;
  assign \new_[40215]_  = A170 & \new_[40214]_ ;
  assign \new_[40219]_  = ~A201 & ~A200;
  assign \new_[40220]_  = A166 & \new_[40219]_ ;
  assign \new_[40221]_  = \new_[40220]_  & \new_[40215]_ ;
  assign \new_[40225]_  = ~A265 & ~A234;
  assign \new_[40226]_  = ~A233 & \new_[40225]_ ;
  assign \new_[40230]_  = A299 & A298;
  assign \new_[40231]_  = ~A266 & \new_[40230]_ ;
  assign \new_[40232]_  = \new_[40231]_  & \new_[40226]_ ;
  assign \new_[40236]_  = ~A167 & ~A169;
  assign \new_[40237]_  = A170 & \new_[40236]_ ;
  assign \new_[40241]_  = ~A201 & ~A200;
  assign \new_[40242]_  = A166 & \new_[40241]_ ;
  assign \new_[40243]_  = \new_[40242]_  & \new_[40237]_ ;
  assign \new_[40247]_  = ~A265 & ~A234;
  assign \new_[40248]_  = ~A233 & \new_[40247]_ ;
  assign \new_[40252]_  = ~A299 & ~A298;
  assign \new_[40253]_  = ~A266 & \new_[40252]_ ;
  assign \new_[40254]_  = \new_[40253]_  & \new_[40248]_ ;
  assign \new_[40258]_  = ~A167 & ~A169;
  assign \new_[40259]_  = A170 & \new_[40258]_ ;
  assign \new_[40263]_  = ~A201 & ~A200;
  assign \new_[40264]_  = A166 & \new_[40263]_ ;
  assign \new_[40265]_  = \new_[40264]_  & \new_[40259]_ ;
  assign \new_[40269]_  = A234 & ~A233;
  assign \new_[40270]_  = A232 & \new_[40269]_ ;
  assign \new_[40274]_  = A299 & ~A298;
  assign \new_[40275]_  = A235 & \new_[40274]_ ;
  assign \new_[40276]_  = \new_[40275]_  & \new_[40270]_ ;
  assign \new_[40280]_  = ~A167 & ~A169;
  assign \new_[40281]_  = A170 & \new_[40280]_ ;
  assign \new_[40285]_  = ~A201 & ~A200;
  assign \new_[40286]_  = A166 & \new_[40285]_ ;
  assign \new_[40287]_  = \new_[40286]_  & \new_[40281]_ ;
  assign \new_[40291]_  = A234 & ~A233;
  assign \new_[40292]_  = A232 & \new_[40291]_ ;
  assign \new_[40296]_  = A266 & ~A265;
  assign \new_[40297]_  = A235 & \new_[40296]_ ;
  assign \new_[40298]_  = \new_[40297]_  & \new_[40292]_ ;
  assign \new_[40302]_  = ~A167 & ~A169;
  assign \new_[40303]_  = A170 & \new_[40302]_ ;
  assign \new_[40307]_  = ~A201 & ~A200;
  assign \new_[40308]_  = A166 & \new_[40307]_ ;
  assign \new_[40309]_  = \new_[40308]_  & \new_[40303]_ ;
  assign \new_[40313]_  = A234 & ~A233;
  assign \new_[40314]_  = A232 & \new_[40313]_ ;
  assign \new_[40318]_  = A299 & ~A298;
  assign \new_[40319]_  = A236 & \new_[40318]_ ;
  assign \new_[40320]_  = \new_[40319]_  & \new_[40314]_ ;
  assign \new_[40324]_  = ~A167 & ~A169;
  assign \new_[40325]_  = A170 & \new_[40324]_ ;
  assign \new_[40329]_  = ~A201 & ~A200;
  assign \new_[40330]_  = A166 & \new_[40329]_ ;
  assign \new_[40331]_  = \new_[40330]_  & \new_[40325]_ ;
  assign \new_[40335]_  = A234 & ~A233;
  assign \new_[40336]_  = A232 & \new_[40335]_ ;
  assign \new_[40340]_  = A266 & ~A265;
  assign \new_[40341]_  = A236 & \new_[40340]_ ;
  assign \new_[40342]_  = \new_[40341]_  & \new_[40336]_ ;
  assign \new_[40346]_  = ~A167 & ~A169;
  assign \new_[40347]_  = A170 & \new_[40346]_ ;
  assign \new_[40351]_  = ~A201 & ~A200;
  assign \new_[40352]_  = A166 & \new_[40351]_ ;
  assign \new_[40353]_  = \new_[40352]_  & \new_[40347]_ ;
  assign \new_[40357]_  = A265 & ~A233;
  assign \new_[40358]_  = ~A232 & \new_[40357]_ ;
  assign \new_[40362]_  = ~A300 & A298;
  assign \new_[40363]_  = A266 & \new_[40362]_ ;
  assign \new_[40364]_  = \new_[40363]_  & \new_[40358]_ ;
  assign \new_[40368]_  = ~A167 & ~A169;
  assign \new_[40369]_  = A170 & \new_[40368]_ ;
  assign \new_[40373]_  = ~A201 & ~A200;
  assign \new_[40374]_  = A166 & \new_[40373]_ ;
  assign \new_[40375]_  = \new_[40374]_  & \new_[40369]_ ;
  assign \new_[40379]_  = A265 & ~A233;
  assign \new_[40380]_  = ~A232 & \new_[40379]_ ;
  assign \new_[40384]_  = A299 & A298;
  assign \new_[40385]_  = A266 & \new_[40384]_ ;
  assign \new_[40386]_  = \new_[40385]_  & \new_[40380]_ ;
  assign \new_[40390]_  = ~A167 & ~A169;
  assign \new_[40391]_  = A170 & \new_[40390]_ ;
  assign \new_[40395]_  = ~A201 & ~A200;
  assign \new_[40396]_  = A166 & \new_[40395]_ ;
  assign \new_[40397]_  = \new_[40396]_  & \new_[40391]_ ;
  assign \new_[40401]_  = A265 & ~A233;
  assign \new_[40402]_  = ~A232 & \new_[40401]_ ;
  assign \new_[40406]_  = ~A299 & ~A298;
  assign \new_[40407]_  = A266 & \new_[40406]_ ;
  assign \new_[40408]_  = \new_[40407]_  & \new_[40402]_ ;
  assign \new_[40412]_  = ~A167 & ~A169;
  assign \new_[40413]_  = A170 & \new_[40412]_ ;
  assign \new_[40417]_  = ~A201 & ~A200;
  assign \new_[40418]_  = A166 & \new_[40417]_ ;
  assign \new_[40419]_  = \new_[40418]_  & \new_[40413]_ ;
  assign \new_[40423]_  = ~A266 & ~A233;
  assign \new_[40424]_  = ~A232 & \new_[40423]_ ;
  assign \new_[40428]_  = ~A300 & A298;
  assign \new_[40429]_  = ~A267 & \new_[40428]_ ;
  assign \new_[40430]_  = \new_[40429]_  & \new_[40424]_ ;
  assign \new_[40434]_  = ~A167 & ~A169;
  assign \new_[40435]_  = A170 & \new_[40434]_ ;
  assign \new_[40439]_  = ~A201 & ~A200;
  assign \new_[40440]_  = A166 & \new_[40439]_ ;
  assign \new_[40441]_  = \new_[40440]_  & \new_[40435]_ ;
  assign \new_[40445]_  = ~A266 & ~A233;
  assign \new_[40446]_  = ~A232 & \new_[40445]_ ;
  assign \new_[40450]_  = A299 & A298;
  assign \new_[40451]_  = ~A267 & \new_[40450]_ ;
  assign \new_[40452]_  = \new_[40451]_  & \new_[40446]_ ;
  assign \new_[40456]_  = ~A167 & ~A169;
  assign \new_[40457]_  = A170 & \new_[40456]_ ;
  assign \new_[40461]_  = ~A201 & ~A200;
  assign \new_[40462]_  = A166 & \new_[40461]_ ;
  assign \new_[40463]_  = \new_[40462]_  & \new_[40457]_ ;
  assign \new_[40467]_  = ~A266 & ~A233;
  assign \new_[40468]_  = ~A232 & \new_[40467]_ ;
  assign \new_[40472]_  = ~A299 & ~A298;
  assign \new_[40473]_  = ~A267 & \new_[40472]_ ;
  assign \new_[40474]_  = \new_[40473]_  & \new_[40468]_ ;
  assign \new_[40478]_  = ~A167 & ~A169;
  assign \new_[40479]_  = A170 & \new_[40478]_ ;
  assign \new_[40483]_  = ~A201 & ~A200;
  assign \new_[40484]_  = A166 & \new_[40483]_ ;
  assign \new_[40485]_  = \new_[40484]_  & \new_[40479]_ ;
  assign \new_[40489]_  = ~A265 & ~A233;
  assign \new_[40490]_  = ~A232 & \new_[40489]_ ;
  assign \new_[40494]_  = ~A300 & A298;
  assign \new_[40495]_  = ~A266 & \new_[40494]_ ;
  assign \new_[40496]_  = \new_[40495]_  & \new_[40490]_ ;
  assign \new_[40500]_  = ~A167 & ~A169;
  assign \new_[40501]_  = A170 & \new_[40500]_ ;
  assign \new_[40505]_  = ~A201 & ~A200;
  assign \new_[40506]_  = A166 & \new_[40505]_ ;
  assign \new_[40507]_  = \new_[40506]_  & \new_[40501]_ ;
  assign \new_[40511]_  = ~A265 & ~A233;
  assign \new_[40512]_  = ~A232 & \new_[40511]_ ;
  assign \new_[40516]_  = A299 & A298;
  assign \new_[40517]_  = ~A266 & \new_[40516]_ ;
  assign \new_[40518]_  = \new_[40517]_  & \new_[40512]_ ;
  assign \new_[40522]_  = ~A167 & ~A169;
  assign \new_[40523]_  = A170 & \new_[40522]_ ;
  assign \new_[40527]_  = ~A201 & ~A200;
  assign \new_[40528]_  = A166 & \new_[40527]_ ;
  assign \new_[40529]_  = \new_[40528]_  & \new_[40523]_ ;
  assign \new_[40533]_  = ~A265 & ~A233;
  assign \new_[40534]_  = ~A232 & \new_[40533]_ ;
  assign \new_[40538]_  = ~A299 & ~A298;
  assign \new_[40539]_  = ~A266 & \new_[40538]_ ;
  assign \new_[40540]_  = \new_[40539]_  & \new_[40534]_ ;
  assign \new_[40544]_  = ~A167 & ~A169;
  assign \new_[40545]_  = A170 & \new_[40544]_ ;
  assign \new_[40549]_  = ~A200 & ~A199;
  assign \new_[40550]_  = A166 & \new_[40549]_ ;
  assign \new_[40551]_  = \new_[40550]_  & \new_[40545]_ ;
  assign \new_[40555]_  = A265 & A233;
  assign \new_[40556]_  = A232 & \new_[40555]_ ;
  assign \new_[40560]_  = ~A300 & ~A299;
  assign \new_[40561]_  = ~A267 & \new_[40560]_ ;
  assign \new_[40562]_  = \new_[40561]_  & \new_[40556]_ ;
  assign \new_[40566]_  = ~A167 & ~A169;
  assign \new_[40567]_  = A170 & \new_[40566]_ ;
  assign \new_[40571]_  = ~A200 & ~A199;
  assign \new_[40572]_  = A166 & \new_[40571]_ ;
  assign \new_[40573]_  = \new_[40572]_  & \new_[40567]_ ;
  assign \new_[40577]_  = A265 & A233;
  assign \new_[40578]_  = A232 & \new_[40577]_ ;
  assign \new_[40582]_  = A299 & A298;
  assign \new_[40583]_  = ~A267 & \new_[40582]_ ;
  assign \new_[40584]_  = \new_[40583]_  & \new_[40578]_ ;
  assign \new_[40588]_  = ~A167 & ~A169;
  assign \new_[40589]_  = A170 & \new_[40588]_ ;
  assign \new_[40593]_  = ~A200 & ~A199;
  assign \new_[40594]_  = A166 & \new_[40593]_ ;
  assign \new_[40595]_  = \new_[40594]_  & \new_[40589]_ ;
  assign \new_[40599]_  = A265 & A233;
  assign \new_[40600]_  = A232 & \new_[40599]_ ;
  assign \new_[40604]_  = ~A299 & ~A298;
  assign \new_[40605]_  = ~A267 & \new_[40604]_ ;
  assign \new_[40606]_  = \new_[40605]_  & \new_[40600]_ ;
  assign \new_[40610]_  = ~A167 & ~A169;
  assign \new_[40611]_  = A170 & \new_[40610]_ ;
  assign \new_[40615]_  = ~A200 & ~A199;
  assign \new_[40616]_  = A166 & \new_[40615]_ ;
  assign \new_[40617]_  = \new_[40616]_  & \new_[40611]_ ;
  assign \new_[40621]_  = A265 & A233;
  assign \new_[40622]_  = A232 & \new_[40621]_ ;
  assign \new_[40626]_  = ~A300 & ~A299;
  assign \new_[40627]_  = A266 & \new_[40626]_ ;
  assign \new_[40628]_  = \new_[40627]_  & \new_[40622]_ ;
  assign \new_[40632]_  = ~A167 & ~A169;
  assign \new_[40633]_  = A170 & \new_[40632]_ ;
  assign \new_[40637]_  = ~A200 & ~A199;
  assign \new_[40638]_  = A166 & \new_[40637]_ ;
  assign \new_[40639]_  = \new_[40638]_  & \new_[40633]_ ;
  assign \new_[40643]_  = A265 & A233;
  assign \new_[40644]_  = A232 & \new_[40643]_ ;
  assign \new_[40648]_  = A299 & A298;
  assign \new_[40649]_  = A266 & \new_[40648]_ ;
  assign \new_[40650]_  = \new_[40649]_  & \new_[40644]_ ;
  assign \new_[40654]_  = ~A167 & ~A169;
  assign \new_[40655]_  = A170 & \new_[40654]_ ;
  assign \new_[40659]_  = ~A200 & ~A199;
  assign \new_[40660]_  = A166 & \new_[40659]_ ;
  assign \new_[40661]_  = \new_[40660]_  & \new_[40655]_ ;
  assign \new_[40665]_  = A265 & A233;
  assign \new_[40666]_  = A232 & \new_[40665]_ ;
  assign \new_[40670]_  = ~A299 & ~A298;
  assign \new_[40671]_  = A266 & \new_[40670]_ ;
  assign \new_[40672]_  = \new_[40671]_  & \new_[40666]_ ;
  assign \new_[40676]_  = ~A167 & ~A169;
  assign \new_[40677]_  = A170 & \new_[40676]_ ;
  assign \new_[40681]_  = ~A200 & ~A199;
  assign \new_[40682]_  = A166 & \new_[40681]_ ;
  assign \new_[40683]_  = \new_[40682]_  & \new_[40677]_ ;
  assign \new_[40687]_  = ~A265 & A233;
  assign \new_[40688]_  = A232 & \new_[40687]_ ;
  assign \new_[40692]_  = ~A300 & ~A299;
  assign \new_[40693]_  = ~A266 & \new_[40692]_ ;
  assign \new_[40694]_  = \new_[40693]_  & \new_[40688]_ ;
  assign \new_[40698]_  = ~A167 & ~A169;
  assign \new_[40699]_  = A170 & \new_[40698]_ ;
  assign \new_[40703]_  = ~A200 & ~A199;
  assign \new_[40704]_  = A166 & \new_[40703]_ ;
  assign \new_[40705]_  = \new_[40704]_  & \new_[40699]_ ;
  assign \new_[40709]_  = ~A265 & A233;
  assign \new_[40710]_  = A232 & \new_[40709]_ ;
  assign \new_[40714]_  = A299 & A298;
  assign \new_[40715]_  = ~A266 & \new_[40714]_ ;
  assign \new_[40716]_  = \new_[40715]_  & \new_[40710]_ ;
  assign \new_[40720]_  = ~A167 & ~A169;
  assign \new_[40721]_  = A170 & \new_[40720]_ ;
  assign \new_[40725]_  = ~A200 & ~A199;
  assign \new_[40726]_  = A166 & \new_[40725]_ ;
  assign \new_[40727]_  = \new_[40726]_  & \new_[40721]_ ;
  assign \new_[40731]_  = ~A265 & A233;
  assign \new_[40732]_  = A232 & \new_[40731]_ ;
  assign \new_[40736]_  = ~A299 & ~A298;
  assign \new_[40737]_  = ~A266 & \new_[40736]_ ;
  assign \new_[40738]_  = \new_[40737]_  & \new_[40732]_ ;
  assign \new_[40742]_  = ~A167 & ~A169;
  assign \new_[40743]_  = A170 & \new_[40742]_ ;
  assign \new_[40747]_  = ~A200 & ~A199;
  assign \new_[40748]_  = A166 & \new_[40747]_ ;
  assign \new_[40749]_  = \new_[40748]_  & \new_[40743]_ ;
  assign \new_[40753]_  = A298 & A233;
  assign \new_[40754]_  = ~A232 & \new_[40753]_ ;
  assign \new_[40758]_  = A301 & A300;
  assign \new_[40759]_  = ~A299 & \new_[40758]_ ;
  assign \new_[40760]_  = \new_[40759]_  & \new_[40754]_ ;
  assign \new_[40764]_  = ~A167 & ~A169;
  assign \new_[40765]_  = A170 & \new_[40764]_ ;
  assign \new_[40769]_  = ~A200 & ~A199;
  assign \new_[40770]_  = A166 & \new_[40769]_ ;
  assign \new_[40771]_  = \new_[40770]_  & \new_[40765]_ ;
  assign \new_[40775]_  = A298 & A233;
  assign \new_[40776]_  = ~A232 & \new_[40775]_ ;
  assign \new_[40780]_  = A302 & A300;
  assign \new_[40781]_  = ~A299 & \new_[40780]_ ;
  assign \new_[40782]_  = \new_[40781]_  & \new_[40776]_ ;
  assign \new_[40786]_  = ~A167 & ~A169;
  assign \new_[40787]_  = A170 & \new_[40786]_ ;
  assign \new_[40791]_  = ~A200 & ~A199;
  assign \new_[40792]_  = A166 & \new_[40791]_ ;
  assign \new_[40793]_  = \new_[40792]_  & \new_[40787]_ ;
  assign \new_[40797]_  = A265 & A233;
  assign \new_[40798]_  = ~A232 & \new_[40797]_ ;
  assign \new_[40802]_  = A268 & A267;
  assign \new_[40803]_  = ~A266 & \new_[40802]_ ;
  assign \new_[40804]_  = \new_[40803]_  & \new_[40798]_ ;
  assign \new_[40808]_  = ~A167 & ~A169;
  assign \new_[40809]_  = A170 & \new_[40808]_ ;
  assign \new_[40813]_  = ~A200 & ~A199;
  assign \new_[40814]_  = A166 & \new_[40813]_ ;
  assign \new_[40815]_  = \new_[40814]_  & \new_[40809]_ ;
  assign \new_[40819]_  = A265 & A233;
  assign \new_[40820]_  = ~A232 & \new_[40819]_ ;
  assign \new_[40824]_  = A269 & A267;
  assign \new_[40825]_  = ~A266 & \new_[40824]_ ;
  assign \new_[40826]_  = \new_[40825]_  & \new_[40820]_ ;
  assign \new_[40830]_  = ~A167 & ~A169;
  assign \new_[40831]_  = A170 & \new_[40830]_ ;
  assign \new_[40835]_  = ~A200 & ~A199;
  assign \new_[40836]_  = A166 & \new_[40835]_ ;
  assign \new_[40837]_  = \new_[40836]_  & \new_[40831]_ ;
  assign \new_[40841]_  = A265 & ~A234;
  assign \new_[40842]_  = ~A233 & \new_[40841]_ ;
  assign \new_[40846]_  = ~A300 & A298;
  assign \new_[40847]_  = A266 & \new_[40846]_ ;
  assign \new_[40848]_  = \new_[40847]_  & \new_[40842]_ ;
  assign \new_[40852]_  = ~A167 & ~A169;
  assign \new_[40853]_  = A170 & \new_[40852]_ ;
  assign \new_[40857]_  = ~A200 & ~A199;
  assign \new_[40858]_  = A166 & \new_[40857]_ ;
  assign \new_[40859]_  = \new_[40858]_  & \new_[40853]_ ;
  assign \new_[40863]_  = A265 & ~A234;
  assign \new_[40864]_  = ~A233 & \new_[40863]_ ;
  assign \new_[40868]_  = A299 & A298;
  assign \new_[40869]_  = A266 & \new_[40868]_ ;
  assign \new_[40870]_  = \new_[40869]_  & \new_[40864]_ ;
  assign \new_[40874]_  = ~A167 & ~A169;
  assign \new_[40875]_  = A170 & \new_[40874]_ ;
  assign \new_[40879]_  = ~A200 & ~A199;
  assign \new_[40880]_  = A166 & \new_[40879]_ ;
  assign \new_[40881]_  = \new_[40880]_  & \new_[40875]_ ;
  assign \new_[40885]_  = A265 & ~A234;
  assign \new_[40886]_  = ~A233 & \new_[40885]_ ;
  assign \new_[40890]_  = ~A299 & ~A298;
  assign \new_[40891]_  = A266 & \new_[40890]_ ;
  assign \new_[40892]_  = \new_[40891]_  & \new_[40886]_ ;
  assign \new_[40896]_  = ~A167 & ~A169;
  assign \new_[40897]_  = A170 & \new_[40896]_ ;
  assign \new_[40901]_  = ~A200 & ~A199;
  assign \new_[40902]_  = A166 & \new_[40901]_ ;
  assign \new_[40903]_  = \new_[40902]_  & \new_[40897]_ ;
  assign \new_[40907]_  = ~A266 & ~A234;
  assign \new_[40908]_  = ~A233 & \new_[40907]_ ;
  assign \new_[40912]_  = ~A300 & A298;
  assign \new_[40913]_  = ~A267 & \new_[40912]_ ;
  assign \new_[40914]_  = \new_[40913]_  & \new_[40908]_ ;
  assign \new_[40918]_  = ~A167 & ~A169;
  assign \new_[40919]_  = A170 & \new_[40918]_ ;
  assign \new_[40923]_  = ~A200 & ~A199;
  assign \new_[40924]_  = A166 & \new_[40923]_ ;
  assign \new_[40925]_  = \new_[40924]_  & \new_[40919]_ ;
  assign \new_[40929]_  = ~A266 & ~A234;
  assign \new_[40930]_  = ~A233 & \new_[40929]_ ;
  assign \new_[40934]_  = A299 & A298;
  assign \new_[40935]_  = ~A267 & \new_[40934]_ ;
  assign \new_[40936]_  = \new_[40935]_  & \new_[40930]_ ;
  assign \new_[40940]_  = ~A167 & ~A169;
  assign \new_[40941]_  = A170 & \new_[40940]_ ;
  assign \new_[40945]_  = ~A200 & ~A199;
  assign \new_[40946]_  = A166 & \new_[40945]_ ;
  assign \new_[40947]_  = \new_[40946]_  & \new_[40941]_ ;
  assign \new_[40951]_  = ~A266 & ~A234;
  assign \new_[40952]_  = ~A233 & \new_[40951]_ ;
  assign \new_[40956]_  = ~A299 & ~A298;
  assign \new_[40957]_  = ~A267 & \new_[40956]_ ;
  assign \new_[40958]_  = \new_[40957]_  & \new_[40952]_ ;
  assign \new_[40962]_  = ~A167 & ~A169;
  assign \new_[40963]_  = A170 & \new_[40962]_ ;
  assign \new_[40967]_  = ~A200 & ~A199;
  assign \new_[40968]_  = A166 & \new_[40967]_ ;
  assign \new_[40969]_  = \new_[40968]_  & \new_[40963]_ ;
  assign \new_[40973]_  = ~A265 & ~A234;
  assign \new_[40974]_  = ~A233 & \new_[40973]_ ;
  assign \new_[40978]_  = ~A300 & A298;
  assign \new_[40979]_  = ~A266 & \new_[40978]_ ;
  assign \new_[40980]_  = \new_[40979]_  & \new_[40974]_ ;
  assign \new_[40984]_  = ~A167 & ~A169;
  assign \new_[40985]_  = A170 & \new_[40984]_ ;
  assign \new_[40989]_  = ~A200 & ~A199;
  assign \new_[40990]_  = A166 & \new_[40989]_ ;
  assign \new_[40991]_  = \new_[40990]_  & \new_[40985]_ ;
  assign \new_[40995]_  = ~A265 & ~A234;
  assign \new_[40996]_  = ~A233 & \new_[40995]_ ;
  assign \new_[41000]_  = A299 & A298;
  assign \new_[41001]_  = ~A266 & \new_[41000]_ ;
  assign \new_[41002]_  = \new_[41001]_  & \new_[40996]_ ;
  assign \new_[41006]_  = ~A167 & ~A169;
  assign \new_[41007]_  = A170 & \new_[41006]_ ;
  assign \new_[41011]_  = ~A200 & ~A199;
  assign \new_[41012]_  = A166 & \new_[41011]_ ;
  assign \new_[41013]_  = \new_[41012]_  & \new_[41007]_ ;
  assign \new_[41017]_  = ~A265 & ~A234;
  assign \new_[41018]_  = ~A233 & \new_[41017]_ ;
  assign \new_[41022]_  = ~A299 & ~A298;
  assign \new_[41023]_  = ~A266 & \new_[41022]_ ;
  assign \new_[41024]_  = \new_[41023]_  & \new_[41018]_ ;
  assign \new_[41028]_  = ~A167 & ~A169;
  assign \new_[41029]_  = A170 & \new_[41028]_ ;
  assign \new_[41033]_  = ~A200 & ~A199;
  assign \new_[41034]_  = A166 & \new_[41033]_ ;
  assign \new_[41035]_  = \new_[41034]_  & \new_[41029]_ ;
  assign \new_[41039]_  = A234 & ~A233;
  assign \new_[41040]_  = A232 & \new_[41039]_ ;
  assign \new_[41044]_  = A299 & ~A298;
  assign \new_[41045]_  = A235 & \new_[41044]_ ;
  assign \new_[41046]_  = \new_[41045]_  & \new_[41040]_ ;
  assign \new_[41050]_  = ~A167 & ~A169;
  assign \new_[41051]_  = A170 & \new_[41050]_ ;
  assign \new_[41055]_  = ~A200 & ~A199;
  assign \new_[41056]_  = A166 & \new_[41055]_ ;
  assign \new_[41057]_  = \new_[41056]_  & \new_[41051]_ ;
  assign \new_[41061]_  = A234 & ~A233;
  assign \new_[41062]_  = A232 & \new_[41061]_ ;
  assign \new_[41066]_  = A266 & ~A265;
  assign \new_[41067]_  = A235 & \new_[41066]_ ;
  assign \new_[41068]_  = \new_[41067]_  & \new_[41062]_ ;
  assign \new_[41072]_  = ~A167 & ~A169;
  assign \new_[41073]_  = A170 & \new_[41072]_ ;
  assign \new_[41077]_  = ~A200 & ~A199;
  assign \new_[41078]_  = A166 & \new_[41077]_ ;
  assign \new_[41079]_  = \new_[41078]_  & \new_[41073]_ ;
  assign \new_[41083]_  = A234 & ~A233;
  assign \new_[41084]_  = A232 & \new_[41083]_ ;
  assign \new_[41088]_  = A299 & ~A298;
  assign \new_[41089]_  = A236 & \new_[41088]_ ;
  assign \new_[41090]_  = \new_[41089]_  & \new_[41084]_ ;
  assign \new_[41094]_  = ~A167 & ~A169;
  assign \new_[41095]_  = A170 & \new_[41094]_ ;
  assign \new_[41099]_  = ~A200 & ~A199;
  assign \new_[41100]_  = A166 & \new_[41099]_ ;
  assign \new_[41101]_  = \new_[41100]_  & \new_[41095]_ ;
  assign \new_[41105]_  = A234 & ~A233;
  assign \new_[41106]_  = A232 & \new_[41105]_ ;
  assign \new_[41110]_  = A266 & ~A265;
  assign \new_[41111]_  = A236 & \new_[41110]_ ;
  assign \new_[41112]_  = \new_[41111]_  & \new_[41106]_ ;
  assign \new_[41116]_  = ~A167 & ~A169;
  assign \new_[41117]_  = A170 & \new_[41116]_ ;
  assign \new_[41121]_  = ~A200 & ~A199;
  assign \new_[41122]_  = A166 & \new_[41121]_ ;
  assign \new_[41123]_  = \new_[41122]_  & \new_[41117]_ ;
  assign \new_[41127]_  = A265 & ~A233;
  assign \new_[41128]_  = ~A232 & \new_[41127]_ ;
  assign \new_[41132]_  = ~A300 & A298;
  assign \new_[41133]_  = A266 & \new_[41132]_ ;
  assign \new_[41134]_  = \new_[41133]_  & \new_[41128]_ ;
  assign \new_[41138]_  = ~A167 & ~A169;
  assign \new_[41139]_  = A170 & \new_[41138]_ ;
  assign \new_[41143]_  = ~A200 & ~A199;
  assign \new_[41144]_  = A166 & \new_[41143]_ ;
  assign \new_[41145]_  = \new_[41144]_  & \new_[41139]_ ;
  assign \new_[41149]_  = A265 & ~A233;
  assign \new_[41150]_  = ~A232 & \new_[41149]_ ;
  assign \new_[41154]_  = A299 & A298;
  assign \new_[41155]_  = A266 & \new_[41154]_ ;
  assign \new_[41156]_  = \new_[41155]_  & \new_[41150]_ ;
  assign \new_[41160]_  = ~A167 & ~A169;
  assign \new_[41161]_  = A170 & \new_[41160]_ ;
  assign \new_[41165]_  = ~A200 & ~A199;
  assign \new_[41166]_  = A166 & \new_[41165]_ ;
  assign \new_[41167]_  = \new_[41166]_  & \new_[41161]_ ;
  assign \new_[41171]_  = A265 & ~A233;
  assign \new_[41172]_  = ~A232 & \new_[41171]_ ;
  assign \new_[41176]_  = ~A299 & ~A298;
  assign \new_[41177]_  = A266 & \new_[41176]_ ;
  assign \new_[41178]_  = \new_[41177]_  & \new_[41172]_ ;
  assign \new_[41182]_  = ~A167 & ~A169;
  assign \new_[41183]_  = A170 & \new_[41182]_ ;
  assign \new_[41187]_  = ~A200 & ~A199;
  assign \new_[41188]_  = A166 & \new_[41187]_ ;
  assign \new_[41189]_  = \new_[41188]_  & \new_[41183]_ ;
  assign \new_[41193]_  = ~A266 & ~A233;
  assign \new_[41194]_  = ~A232 & \new_[41193]_ ;
  assign \new_[41198]_  = ~A300 & A298;
  assign \new_[41199]_  = ~A267 & \new_[41198]_ ;
  assign \new_[41200]_  = \new_[41199]_  & \new_[41194]_ ;
  assign \new_[41204]_  = ~A167 & ~A169;
  assign \new_[41205]_  = A170 & \new_[41204]_ ;
  assign \new_[41209]_  = ~A200 & ~A199;
  assign \new_[41210]_  = A166 & \new_[41209]_ ;
  assign \new_[41211]_  = \new_[41210]_  & \new_[41205]_ ;
  assign \new_[41215]_  = ~A266 & ~A233;
  assign \new_[41216]_  = ~A232 & \new_[41215]_ ;
  assign \new_[41220]_  = A299 & A298;
  assign \new_[41221]_  = ~A267 & \new_[41220]_ ;
  assign \new_[41222]_  = \new_[41221]_  & \new_[41216]_ ;
  assign \new_[41226]_  = ~A167 & ~A169;
  assign \new_[41227]_  = A170 & \new_[41226]_ ;
  assign \new_[41231]_  = ~A200 & ~A199;
  assign \new_[41232]_  = A166 & \new_[41231]_ ;
  assign \new_[41233]_  = \new_[41232]_  & \new_[41227]_ ;
  assign \new_[41237]_  = ~A266 & ~A233;
  assign \new_[41238]_  = ~A232 & \new_[41237]_ ;
  assign \new_[41242]_  = ~A299 & ~A298;
  assign \new_[41243]_  = ~A267 & \new_[41242]_ ;
  assign \new_[41244]_  = \new_[41243]_  & \new_[41238]_ ;
  assign \new_[41248]_  = ~A167 & ~A169;
  assign \new_[41249]_  = A170 & \new_[41248]_ ;
  assign \new_[41253]_  = ~A200 & ~A199;
  assign \new_[41254]_  = A166 & \new_[41253]_ ;
  assign \new_[41255]_  = \new_[41254]_  & \new_[41249]_ ;
  assign \new_[41259]_  = ~A265 & ~A233;
  assign \new_[41260]_  = ~A232 & \new_[41259]_ ;
  assign \new_[41264]_  = ~A300 & A298;
  assign \new_[41265]_  = ~A266 & \new_[41264]_ ;
  assign \new_[41266]_  = \new_[41265]_  & \new_[41260]_ ;
  assign \new_[41270]_  = ~A167 & ~A169;
  assign \new_[41271]_  = A170 & \new_[41270]_ ;
  assign \new_[41275]_  = ~A200 & ~A199;
  assign \new_[41276]_  = A166 & \new_[41275]_ ;
  assign \new_[41277]_  = \new_[41276]_  & \new_[41271]_ ;
  assign \new_[41281]_  = ~A265 & ~A233;
  assign \new_[41282]_  = ~A232 & \new_[41281]_ ;
  assign \new_[41286]_  = A299 & A298;
  assign \new_[41287]_  = ~A266 & \new_[41286]_ ;
  assign \new_[41288]_  = \new_[41287]_  & \new_[41282]_ ;
  assign \new_[41292]_  = ~A167 & ~A169;
  assign \new_[41293]_  = A170 & \new_[41292]_ ;
  assign \new_[41297]_  = ~A200 & ~A199;
  assign \new_[41298]_  = A166 & \new_[41297]_ ;
  assign \new_[41299]_  = \new_[41298]_  & \new_[41293]_ ;
  assign \new_[41303]_  = ~A265 & ~A233;
  assign \new_[41304]_  = ~A232 & \new_[41303]_ ;
  assign \new_[41308]_  = ~A299 & ~A298;
  assign \new_[41309]_  = ~A266 & \new_[41308]_ ;
  assign \new_[41310]_  = \new_[41309]_  & \new_[41304]_ ;
  assign \new_[41314]_  = A199 & A166;
  assign \new_[41315]_  = A168 & \new_[41314]_ ;
  assign \new_[41319]_  = ~A235 & ~A233;
  assign \new_[41320]_  = A200 & \new_[41319]_ ;
  assign \new_[41321]_  = \new_[41320]_  & \new_[41315]_ ;
  assign \new_[41325]_  = ~A268 & ~A266;
  assign \new_[41326]_  = ~A236 & \new_[41325]_ ;
  assign \new_[41329]_  = A298 & ~A269;
  assign \new_[41332]_  = ~A302 & ~A301;
  assign \new_[41333]_  = \new_[41332]_  & \new_[41329]_ ;
  assign \new_[41334]_  = \new_[41333]_  & \new_[41326]_ ;
  assign \new_[41338]_  = ~A200 & A166;
  assign \new_[41339]_  = A168 & \new_[41338]_ ;
  assign \new_[41343]_  = A232 & ~A203;
  assign \new_[41344]_  = ~A202 & \new_[41343]_ ;
  assign \new_[41345]_  = \new_[41344]_  & \new_[41339]_ ;
  assign \new_[41349]_  = ~A268 & A265;
  assign \new_[41350]_  = A233 & \new_[41349]_ ;
  assign \new_[41353]_  = ~A299 & ~A269;
  assign \new_[41356]_  = ~A302 & ~A301;
  assign \new_[41357]_  = \new_[41356]_  & \new_[41353]_ ;
  assign \new_[41358]_  = \new_[41357]_  & \new_[41350]_ ;
  assign \new_[41362]_  = ~A200 & A166;
  assign \new_[41363]_  = A168 & \new_[41362]_ ;
  assign \new_[41367]_  = ~A233 & ~A203;
  assign \new_[41368]_  = ~A202 & \new_[41367]_ ;
  assign \new_[41369]_  = \new_[41368]_  & \new_[41363]_ ;
  assign \new_[41373]_  = A265 & ~A236;
  assign \new_[41374]_  = ~A235 & \new_[41373]_ ;
  assign \new_[41377]_  = A298 & A266;
  assign \new_[41380]_  = ~A302 & ~A301;
  assign \new_[41381]_  = \new_[41380]_  & \new_[41377]_ ;
  assign \new_[41382]_  = \new_[41381]_  & \new_[41374]_ ;
  assign \new_[41386]_  = ~A200 & A166;
  assign \new_[41387]_  = A168 & \new_[41386]_ ;
  assign \new_[41391]_  = ~A233 & ~A203;
  assign \new_[41392]_  = ~A202 & \new_[41391]_ ;
  assign \new_[41393]_  = \new_[41392]_  & \new_[41387]_ ;
  assign \new_[41397]_  = ~A266 & ~A236;
  assign \new_[41398]_  = ~A235 & \new_[41397]_ ;
  assign \new_[41401]_  = ~A269 & ~A268;
  assign \new_[41404]_  = ~A300 & A298;
  assign \new_[41405]_  = \new_[41404]_  & \new_[41401]_ ;
  assign \new_[41406]_  = \new_[41405]_  & \new_[41398]_ ;
  assign \new_[41410]_  = ~A200 & A166;
  assign \new_[41411]_  = A168 & \new_[41410]_ ;
  assign \new_[41415]_  = ~A233 & ~A203;
  assign \new_[41416]_  = ~A202 & \new_[41415]_ ;
  assign \new_[41417]_  = \new_[41416]_  & \new_[41411]_ ;
  assign \new_[41421]_  = ~A266 & ~A236;
  assign \new_[41422]_  = ~A235 & \new_[41421]_ ;
  assign \new_[41425]_  = ~A269 & ~A268;
  assign \new_[41428]_  = A299 & A298;
  assign \new_[41429]_  = \new_[41428]_  & \new_[41425]_ ;
  assign \new_[41430]_  = \new_[41429]_  & \new_[41422]_ ;
  assign \new_[41434]_  = ~A200 & A166;
  assign \new_[41435]_  = A168 & \new_[41434]_ ;
  assign \new_[41439]_  = ~A233 & ~A203;
  assign \new_[41440]_  = ~A202 & \new_[41439]_ ;
  assign \new_[41441]_  = \new_[41440]_  & \new_[41435]_ ;
  assign \new_[41445]_  = ~A266 & ~A236;
  assign \new_[41446]_  = ~A235 & \new_[41445]_ ;
  assign \new_[41449]_  = ~A269 & ~A268;
  assign \new_[41452]_  = ~A299 & ~A298;
  assign \new_[41453]_  = \new_[41452]_  & \new_[41449]_ ;
  assign \new_[41454]_  = \new_[41453]_  & \new_[41446]_ ;
  assign \new_[41458]_  = ~A200 & A166;
  assign \new_[41459]_  = A168 & \new_[41458]_ ;
  assign \new_[41463]_  = ~A233 & ~A203;
  assign \new_[41464]_  = ~A202 & \new_[41463]_ ;
  assign \new_[41465]_  = \new_[41464]_  & \new_[41459]_ ;
  assign \new_[41469]_  = ~A266 & ~A236;
  assign \new_[41470]_  = ~A235 & \new_[41469]_ ;
  assign \new_[41473]_  = A298 & ~A267;
  assign \new_[41476]_  = ~A302 & ~A301;
  assign \new_[41477]_  = \new_[41476]_  & \new_[41473]_ ;
  assign \new_[41478]_  = \new_[41477]_  & \new_[41470]_ ;
  assign \new_[41482]_  = ~A200 & A166;
  assign \new_[41483]_  = A168 & \new_[41482]_ ;
  assign \new_[41487]_  = ~A233 & ~A203;
  assign \new_[41488]_  = ~A202 & \new_[41487]_ ;
  assign \new_[41489]_  = \new_[41488]_  & \new_[41483]_ ;
  assign \new_[41493]_  = ~A265 & ~A236;
  assign \new_[41494]_  = ~A235 & \new_[41493]_ ;
  assign \new_[41497]_  = A298 & ~A266;
  assign \new_[41500]_  = ~A302 & ~A301;
  assign \new_[41501]_  = \new_[41500]_  & \new_[41497]_ ;
  assign \new_[41502]_  = \new_[41501]_  & \new_[41494]_ ;
  assign \new_[41506]_  = ~A200 & A166;
  assign \new_[41507]_  = A168 & \new_[41506]_ ;
  assign \new_[41511]_  = ~A233 & ~A203;
  assign \new_[41512]_  = ~A202 & \new_[41511]_ ;
  assign \new_[41513]_  = \new_[41512]_  & \new_[41507]_ ;
  assign \new_[41517]_  = ~A268 & ~A266;
  assign \new_[41518]_  = ~A234 & \new_[41517]_ ;
  assign \new_[41521]_  = A298 & ~A269;
  assign \new_[41524]_  = ~A302 & ~A301;
  assign \new_[41525]_  = \new_[41524]_  & \new_[41521]_ ;
  assign \new_[41526]_  = \new_[41525]_  & \new_[41518]_ ;
  assign \new_[41530]_  = ~A200 & A166;
  assign \new_[41531]_  = A168 & \new_[41530]_ ;
  assign \new_[41535]_  = A232 & ~A203;
  assign \new_[41536]_  = ~A202 & \new_[41535]_ ;
  assign \new_[41537]_  = \new_[41536]_  & \new_[41531]_ ;
  assign \new_[41541]_  = A235 & A234;
  assign \new_[41542]_  = ~A233 & \new_[41541]_ ;
  assign \new_[41545]_  = ~A299 & A298;
  assign \new_[41548]_  = A301 & A300;
  assign \new_[41549]_  = \new_[41548]_  & \new_[41545]_ ;
  assign \new_[41550]_  = \new_[41549]_  & \new_[41542]_ ;
  assign \new_[41554]_  = ~A200 & A166;
  assign \new_[41555]_  = A168 & \new_[41554]_ ;
  assign \new_[41559]_  = A232 & ~A203;
  assign \new_[41560]_  = ~A202 & \new_[41559]_ ;
  assign \new_[41561]_  = \new_[41560]_  & \new_[41555]_ ;
  assign \new_[41565]_  = A235 & A234;
  assign \new_[41566]_  = ~A233 & \new_[41565]_ ;
  assign \new_[41569]_  = ~A299 & A298;
  assign \new_[41572]_  = A302 & A300;
  assign \new_[41573]_  = \new_[41572]_  & \new_[41569]_ ;
  assign \new_[41574]_  = \new_[41573]_  & \new_[41566]_ ;
  assign \new_[41578]_  = ~A200 & A166;
  assign \new_[41579]_  = A168 & \new_[41578]_ ;
  assign \new_[41583]_  = A232 & ~A203;
  assign \new_[41584]_  = ~A202 & \new_[41583]_ ;
  assign \new_[41585]_  = \new_[41584]_  & \new_[41579]_ ;
  assign \new_[41589]_  = A235 & A234;
  assign \new_[41590]_  = ~A233 & \new_[41589]_ ;
  assign \new_[41593]_  = ~A266 & A265;
  assign \new_[41596]_  = A268 & A267;
  assign \new_[41597]_  = \new_[41596]_  & \new_[41593]_ ;
  assign \new_[41598]_  = \new_[41597]_  & \new_[41590]_ ;
  assign \new_[41602]_  = ~A200 & A166;
  assign \new_[41603]_  = A168 & \new_[41602]_ ;
  assign \new_[41607]_  = A232 & ~A203;
  assign \new_[41608]_  = ~A202 & \new_[41607]_ ;
  assign \new_[41609]_  = \new_[41608]_  & \new_[41603]_ ;
  assign \new_[41613]_  = A235 & A234;
  assign \new_[41614]_  = ~A233 & \new_[41613]_ ;
  assign \new_[41617]_  = ~A266 & A265;
  assign \new_[41620]_  = A269 & A267;
  assign \new_[41621]_  = \new_[41620]_  & \new_[41617]_ ;
  assign \new_[41622]_  = \new_[41621]_  & \new_[41614]_ ;
  assign \new_[41626]_  = ~A200 & A166;
  assign \new_[41627]_  = A168 & \new_[41626]_ ;
  assign \new_[41631]_  = A232 & ~A203;
  assign \new_[41632]_  = ~A202 & \new_[41631]_ ;
  assign \new_[41633]_  = \new_[41632]_  & \new_[41627]_ ;
  assign \new_[41637]_  = A236 & A234;
  assign \new_[41638]_  = ~A233 & \new_[41637]_ ;
  assign \new_[41641]_  = ~A299 & A298;
  assign \new_[41644]_  = A301 & A300;
  assign \new_[41645]_  = \new_[41644]_  & \new_[41641]_ ;
  assign \new_[41646]_  = \new_[41645]_  & \new_[41638]_ ;
  assign \new_[41650]_  = ~A200 & A166;
  assign \new_[41651]_  = A168 & \new_[41650]_ ;
  assign \new_[41655]_  = A232 & ~A203;
  assign \new_[41656]_  = ~A202 & \new_[41655]_ ;
  assign \new_[41657]_  = \new_[41656]_  & \new_[41651]_ ;
  assign \new_[41661]_  = A236 & A234;
  assign \new_[41662]_  = ~A233 & \new_[41661]_ ;
  assign \new_[41665]_  = ~A299 & A298;
  assign \new_[41668]_  = A302 & A300;
  assign \new_[41669]_  = \new_[41668]_  & \new_[41665]_ ;
  assign \new_[41670]_  = \new_[41669]_  & \new_[41662]_ ;
  assign \new_[41674]_  = ~A200 & A166;
  assign \new_[41675]_  = A168 & \new_[41674]_ ;
  assign \new_[41679]_  = A232 & ~A203;
  assign \new_[41680]_  = ~A202 & \new_[41679]_ ;
  assign \new_[41681]_  = \new_[41680]_  & \new_[41675]_ ;
  assign \new_[41685]_  = A236 & A234;
  assign \new_[41686]_  = ~A233 & \new_[41685]_ ;
  assign \new_[41689]_  = ~A266 & A265;
  assign \new_[41692]_  = A268 & A267;
  assign \new_[41693]_  = \new_[41692]_  & \new_[41689]_ ;
  assign \new_[41694]_  = \new_[41693]_  & \new_[41686]_ ;
  assign \new_[41698]_  = ~A200 & A166;
  assign \new_[41699]_  = A168 & \new_[41698]_ ;
  assign \new_[41703]_  = A232 & ~A203;
  assign \new_[41704]_  = ~A202 & \new_[41703]_ ;
  assign \new_[41705]_  = \new_[41704]_  & \new_[41699]_ ;
  assign \new_[41709]_  = A236 & A234;
  assign \new_[41710]_  = ~A233 & \new_[41709]_ ;
  assign \new_[41713]_  = ~A266 & A265;
  assign \new_[41716]_  = A269 & A267;
  assign \new_[41717]_  = \new_[41716]_  & \new_[41713]_ ;
  assign \new_[41718]_  = \new_[41717]_  & \new_[41710]_ ;
  assign \new_[41722]_  = ~A200 & A166;
  assign \new_[41723]_  = A168 & \new_[41722]_ ;
  assign \new_[41727]_  = ~A232 & ~A203;
  assign \new_[41728]_  = ~A202 & \new_[41727]_ ;
  assign \new_[41729]_  = \new_[41728]_  & \new_[41723]_ ;
  assign \new_[41733]_  = ~A268 & ~A266;
  assign \new_[41734]_  = ~A233 & \new_[41733]_ ;
  assign \new_[41737]_  = A298 & ~A269;
  assign \new_[41740]_  = ~A302 & ~A301;
  assign \new_[41741]_  = \new_[41740]_  & \new_[41737]_ ;
  assign \new_[41742]_  = \new_[41741]_  & \new_[41734]_ ;
  assign \new_[41746]_  = ~A200 & A166;
  assign \new_[41747]_  = A168 & \new_[41746]_ ;
  assign \new_[41751]_  = ~A235 & ~A233;
  assign \new_[41752]_  = ~A201 & \new_[41751]_ ;
  assign \new_[41753]_  = \new_[41752]_  & \new_[41747]_ ;
  assign \new_[41757]_  = ~A268 & ~A266;
  assign \new_[41758]_  = ~A236 & \new_[41757]_ ;
  assign \new_[41761]_  = A298 & ~A269;
  assign \new_[41764]_  = ~A302 & ~A301;
  assign \new_[41765]_  = \new_[41764]_  & \new_[41761]_ ;
  assign \new_[41766]_  = \new_[41765]_  & \new_[41758]_ ;
  assign \new_[41770]_  = ~A199 & A166;
  assign \new_[41771]_  = A168 & \new_[41770]_ ;
  assign \new_[41775]_  = ~A235 & ~A233;
  assign \new_[41776]_  = ~A200 & \new_[41775]_ ;
  assign \new_[41777]_  = \new_[41776]_  & \new_[41771]_ ;
  assign \new_[41781]_  = ~A268 & ~A266;
  assign \new_[41782]_  = ~A236 & \new_[41781]_ ;
  assign \new_[41785]_  = A298 & ~A269;
  assign \new_[41788]_  = ~A302 & ~A301;
  assign \new_[41789]_  = \new_[41788]_  & \new_[41785]_ ;
  assign \new_[41790]_  = \new_[41789]_  & \new_[41782]_ ;
  assign \new_[41794]_  = A199 & A167;
  assign \new_[41795]_  = A168 & \new_[41794]_ ;
  assign \new_[41799]_  = ~A235 & ~A233;
  assign \new_[41800]_  = A200 & \new_[41799]_ ;
  assign \new_[41801]_  = \new_[41800]_  & \new_[41795]_ ;
  assign \new_[41805]_  = ~A268 & ~A266;
  assign \new_[41806]_  = ~A236 & \new_[41805]_ ;
  assign \new_[41809]_  = A298 & ~A269;
  assign \new_[41812]_  = ~A302 & ~A301;
  assign \new_[41813]_  = \new_[41812]_  & \new_[41809]_ ;
  assign \new_[41814]_  = \new_[41813]_  & \new_[41806]_ ;
  assign \new_[41818]_  = ~A200 & A167;
  assign \new_[41819]_  = A168 & \new_[41818]_ ;
  assign \new_[41823]_  = A232 & ~A203;
  assign \new_[41824]_  = ~A202 & \new_[41823]_ ;
  assign \new_[41825]_  = \new_[41824]_  & \new_[41819]_ ;
  assign \new_[41829]_  = ~A268 & A265;
  assign \new_[41830]_  = A233 & \new_[41829]_ ;
  assign \new_[41833]_  = ~A299 & ~A269;
  assign \new_[41836]_  = ~A302 & ~A301;
  assign \new_[41837]_  = \new_[41836]_  & \new_[41833]_ ;
  assign \new_[41838]_  = \new_[41837]_  & \new_[41830]_ ;
  assign \new_[41842]_  = ~A200 & A167;
  assign \new_[41843]_  = A168 & \new_[41842]_ ;
  assign \new_[41847]_  = ~A233 & ~A203;
  assign \new_[41848]_  = ~A202 & \new_[41847]_ ;
  assign \new_[41849]_  = \new_[41848]_  & \new_[41843]_ ;
  assign \new_[41853]_  = A265 & ~A236;
  assign \new_[41854]_  = ~A235 & \new_[41853]_ ;
  assign \new_[41857]_  = A298 & A266;
  assign \new_[41860]_  = ~A302 & ~A301;
  assign \new_[41861]_  = \new_[41860]_  & \new_[41857]_ ;
  assign \new_[41862]_  = \new_[41861]_  & \new_[41854]_ ;
  assign \new_[41866]_  = ~A200 & A167;
  assign \new_[41867]_  = A168 & \new_[41866]_ ;
  assign \new_[41871]_  = ~A233 & ~A203;
  assign \new_[41872]_  = ~A202 & \new_[41871]_ ;
  assign \new_[41873]_  = \new_[41872]_  & \new_[41867]_ ;
  assign \new_[41877]_  = ~A266 & ~A236;
  assign \new_[41878]_  = ~A235 & \new_[41877]_ ;
  assign \new_[41881]_  = ~A269 & ~A268;
  assign \new_[41884]_  = ~A300 & A298;
  assign \new_[41885]_  = \new_[41884]_  & \new_[41881]_ ;
  assign \new_[41886]_  = \new_[41885]_  & \new_[41878]_ ;
  assign \new_[41890]_  = ~A200 & A167;
  assign \new_[41891]_  = A168 & \new_[41890]_ ;
  assign \new_[41895]_  = ~A233 & ~A203;
  assign \new_[41896]_  = ~A202 & \new_[41895]_ ;
  assign \new_[41897]_  = \new_[41896]_  & \new_[41891]_ ;
  assign \new_[41901]_  = ~A266 & ~A236;
  assign \new_[41902]_  = ~A235 & \new_[41901]_ ;
  assign \new_[41905]_  = ~A269 & ~A268;
  assign \new_[41908]_  = A299 & A298;
  assign \new_[41909]_  = \new_[41908]_  & \new_[41905]_ ;
  assign \new_[41910]_  = \new_[41909]_  & \new_[41902]_ ;
  assign \new_[41914]_  = ~A200 & A167;
  assign \new_[41915]_  = A168 & \new_[41914]_ ;
  assign \new_[41919]_  = ~A233 & ~A203;
  assign \new_[41920]_  = ~A202 & \new_[41919]_ ;
  assign \new_[41921]_  = \new_[41920]_  & \new_[41915]_ ;
  assign \new_[41925]_  = ~A266 & ~A236;
  assign \new_[41926]_  = ~A235 & \new_[41925]_ ;
  assign \new_[41929]_  = ~A269 & ~A268;
  assign \new_[41932]_  = ~A299 & ~A298;
  assign \new_[41933]_  = \new_[41932]_  & \new_[41929]_ ;
  assign \new_[41934]_  = \new_[41933]_  & \new_[41926]_ ;
  assign \new_[41938]_  = ~A200 & A167;
  assign \new_[41939]_  = A168 & \new_[41938]_ ;
  assign \new_[41943]_  = ~A233 & ~A203;
  assign \new_[41944]_  = ~A202 & \new_[41943]_ ;
  assign \new_[41945]_  = \new_[41944]_  & \new_[41939]_ ;
  assign \new_[41949]_  = ~A266 & ~A236;
  assign \new_[41950]_  = ~A235 & \new_[41949]_ ;
  assign \new_[41953]_  = A298 & ~A267;
  assign \new_[41956]_  = ~A302 & ~A301;
  assign \new_[41957]_  = \new_[41956]_  & \new_[41953]_ ;
  assign \new_[41958]_  = \new_[41957]_  & \new_[41950]_ ;
  assign \new_[41962]_  = ~A200 & A167;
  assign \new_[41963]_  = A168 & \new_[41962]_ ;
  assign \new_[41967]_  = ~A233 & ~A203;
  assign \new_[41968]_  = ~A202 & \new_[41967]_ ;
  assign \new_[41969]_  = \new_[41968]_  & \new_[41963]_ ;
  assign \new_[41973]_  = ~A265 & ~A236;
  assign \new_[41974]_  = ~A235 & \new_[41973]_ ;
  assign \new_[41977]_  = A298 & ~A266;
  assign \new_[41980]_  = ~A302 & ~A301;
  assign \new_[41981]_  = \new_[41980]_  & \new_[41977]_ ;
  assign \new_[41982]_  = \new_[41981]_  & \new_[41974]_ ;
  assign \new_[41986]_  = ~A200 & A167;
  assign \new_[41987]_  = A168 & \new_[41986]_ ;
  assign \new_[41991]_  = ~A233 & ~A203;
  assign \new_[41992]_  = ~A202 & \new_[41991]_ ;
  assign \new_[41993]_  = \new_[41992]_  & \new_[41987]_ ;
  assign \new_[41997]_  = ~A268 & ~A266;
  assign \new_[41998]_  = ~A234 & \new_[41997]_ ;
  assign \new_[42001]_  = A298 & ~A269;
  assign \new_[42004]_  = ~A302 & ~A301;
  assign \new_[42005]_  = \new_[42004]_  & \new_[42001]_ ;
  assign \new_[42006]_  = \new_[42005]_  & \new_[41998]_ ;
  assign \new_[42010]_  = ~A200 & A167;
  assign \new_[42011]_  = A168 & \new_[42010]_ ;
  assign \new_[42015]_  = A232 & ~A203;
  assign \new_[42016]_  = ~A202 & \new_[42015]_ ;
  assign \new_[42017]_  = \new_[42016]_  & \new_[42011]_ ;
  assign \new_[42021]_  = A235 & A234;
  assign \new_[42022]_  = ~A233 & \new_[42021]_ ;
  assign \new_[42025]_  = ~A299 & A298;
  assign \new_[42028]_  = A301 & A300;
  assign \new_[42029]_  = \new_[42028]_  & \new_[42025]_ ;
  assign \new_[42030]_  = \new_[42029]_  & \new_[42022]_ ;
  assign \new_[42034]_  = ~A200 & A167;
  assign \new_[42035]_  = A168 & \new_[42034]_ ;
  assign \new_[42039]_  = A232 & ~A203;
  assign \new_[42040]_  = ~A202 & \new_[42039]_ ;
  assign \new_[42041]_  = \new_[42040]_  & \new_[42035]_ ;
  assign \new_[42045]_  = A235 & A234;
  assign \new_[42046]_  = ~A233 & \new_[42045]_ ;
  assign \new_[42049]_  = ~A299 & A298;
  assign \new_[42052]_  = A302 & A300;
  assign \new_[42053]_  = \new_[42052]_  & \new_[42049]_ ;
  assign \new_[42054]_  = \new_[42053]_  & \new_[42046]_ ;
  assign \new_[42058]_  = ~A200 & A167;
  assign \new_[42059]_  = A168 & \new_[42058]_ ;
  assign \new_[42063]_  = A232 & ~A203;
  assign \new_[42064]_  = ~A202 & \new_[42063]_ ;
  assign \new_[42065]_  = \new_[42064]_  & \new_[42059]_ ;
  assign \new_[42069]_  = A235 & A234;
  assign \new_[42070]_  = ~A233 & \new_[42069]_ ;
  assign \new_[42073]_  = ~A266 & A265;
  assign \new_[42076]_  = A268 & A267;
  assign \new_[42077]_  = \new_[42076]_  & \new_[42073]_ ;
  assign \new_[42078]_  = \new_[42077]_  & \new_[42070]_ ;
  assign \new_[42082]_  = ~A200 & A167;
  assign \new_[42083]_  = A168 & \new_[42082]_ ;
  assign \new_[42087]_  = A232 & ~A203;
  assign \new_[42088]_  = ~A202 & \new_[42087]_ ;
  assign \new_[42089]_  = \new_[42088]_  & \new_[42083]_ ;
  assign \new_[42093]_  = A235 & A234;
  assign \new_[42094]_  = ~A233 & \new_[42093]_ ;
  assign \new_[42097]_  = ~A266 & A265;
  assign \new_[42100]_  = A269 & A267;
  assign \new_[42101]_  = \new_[42100]_  & \new_[42097]_ ;
  assign \new_[42102]_  = \new_[42101]_  & \new_[42094]_ ;
  assign \new_[42106]_  = ~A200 & A167;
  assign \new_[42107]_  = A168 & \new_[42106]_ ;
  assign \new_[42111]_  = A232 & ~A203;
  assign \new_[42112]_  = ~A202 & \new_[42111]_ ;
  assign \new_[42113]_  = \new_[42112]_  & \new_[42107]_ ;
  assign \new_[42117]_  = A236 & A234;
  assign \new_[42118]_  = ~A233 & \new_[42117]_ ;
  assign \new_[42121]_  = ~A299 & A298;
  assign \new_[42124]_  = A301 & A300;
  assign \new_[42125]_  = \new_[42124]_  & \new_[42121]_ ;
  assign \new_[42126]_  = \new_[42125]_  & \new_[42118]_ ;
  assign \new_[42130]_  = ~A200 & A167;
  assign \new_[42131]_  = A168 & \new_[42130]_ ;
  assign \new_[42135]_  = A232 & ~A203;
  assign \new_[42136]_  = ~A202 & \new_[42135]_ ;
  assign \new_[42137]_  = \new_[42136]_  & \new_[42131]_ ;
  assign \new_[42141]_  = A236 & A234;
  assign \new_[42142]_  = ~A233 & \new_[42141]_ ;
  assign \new_[42145]_  = ~A299 & A298;
  assign \new_[42148]_  = A302 & A300;
  assign \new_[42149]_  = \new_[42148]_  & \new_[42145]_ ;
  assign \new_[42150]_  = \new_[42149]_  & \new_[42142]_ ;
  assign \new_[42154]_  = ~A200 & A167;
  assign \new_[42155]_  = A168 & \new_[42154]_ ;
  assign \new_[42159]_  = A232 & ~A203;
  assign \new_[42160]_  = ~A202 & \new_[42159]_ ;
  assign \new_[42161]_  = \new_[42160]_  & \new_[42155]_ ;
  assign \new_[42165]_  = A236 & A234;
  assign \new_[42166]_  = ~A233 & \new_[42165]_ ;
  assign \new_[42169]_  = ~A266 & A265;
  assign \new_[42172]_  = A268 & A267;
  assign \new_[42173]_  = \new_[42172]_  & \new_[42169]_ ;
  assign \new_[42174]_  = \new_[42173]_  & \new_[42166]_ ;
  assign \new_[42178]_  = ~A200 & A167;
  assign \new_[42179]_  = A168 & \new_[42178]_ ;
  assign \new_[42183]_  = A232 & ~A203;
  assign \new_[42184]_  = ~A202 & \new_[42183]_ ;
  assign \new_[42185]_  = \new_[42184]_  & \new_[42179]_ ;
  assign \new_[42189]_  = A236 & A234;
  assign \new_[42190]_  = ~A233 & \new_[42189]_ ;
  assign \new_[42193]_  = ~A266 & A265;
  assign \new_[42196]_  = A269 & A267;
  assign \new_[42197]_  = \new_[42196]_  & \new_[42193]_ ;
  assign \new_[42198]_  = \new_[42197]_  & \new_[42190]_ ;
  assign \new_[42202]_  = ~A200 & A167;
  assign \new_[42203]_  = A168 & \new_[42202]_ ;
  assign \new_[42207]_  = ~A232 & ~A203;
  assign \new_[42208]_  = ~A202 & \new_[42207]_ ;
  assign \new_[42209]_  = \new_[42208]_  & \new_[42203]_ ;
  assign \new_[42213]_  = ~A268 & ~A266;
  assign \new_[42214]_  = ~A233 & \new_[42213]_ ;
  assign \new_[42217]_  = A298 & ~A269;
  assign \new_[42220]_  = ~A302 & ~A301;
  assign \new_[42221]_  = \new_[42220]_  & \new_[42217]_ ;
  assign \new_[42222]_  = \new_[42221]_  & \new_[42214]_ ;
  assign \new_[42226]_  = ~A200 & A167;
  assign \new_[42227]_  = A168 & \new_[42226]_ ;
  assign \new_[42231]_  = ~A235 & ~A233;
  assign \new_[42232]_  = ~A201 & \new_[42231]_ ;
  assign \new_[42233]_  = \new_[42232]_  & \new_[42227]_ ;
  assign \new_[42237]_  = ~A268 & ~A266;
  assign \new_[42238]_  = ~A236 & \new_[42237]_ ;
  assign \new_[42241]_  = A298 & ~A269;
  assign \new_[42244]_  = ~A302 & ~A301;
  assign \new_[42245]_  = \new_[42244]_  & \new_[42241]_ ;
  assign \new_[42246]_  = \new_[42245]_  & \new_[42238]_ ;
  assign \new_[42250]_  = ~A199 & A167;
  assign \new_[42251]_  = A168 & \new_[42250]_ ;
  assign \new_[42255]_  = ~A235 & ~A233;
  assign \new_[42256]_  = ~A200 & \new_[42255]_ ;
  assign \new_[42257]_  = \new_[42256]_  & \new_[42251]_ ;
  assign \new_[42261]_  = ~A268 & ~A266;
  assign \new_[42262]_  = ~A236 & \new_[42261]_ ;
  assign \new_[42265]_  = A298 & ~A269;
  assign \new_[42268]_  = ~A302 & ~A301;
  assign \new_[42269]_  = \new_[42268]_  & \new_[42265]_ ;
  assign \new_[42270]_  = \new_[42269]_  & \new_[42262]_ ;
  assign \new_[42274]_  = ~A166 & ~A167;
  assign \new_[42275]_  = A170 & \new_[42274]_ ;
  assign \new_[42279]_  = A232 & A200;
  assign \new_[42280]_  = ~A199 & \new_[42279]_ ;
  assign \new_[42281]_  = \new_[42280]_  & \new_[42275]_ ;
  assign \new_[42285]_  = ~A268 & A265;
  assign \new_[42286]_  = A233 & \new_[42285]_ ;
  assign \new_[42289]_  = ~A299 & ~A269;
  assign \new_[42292]_  = ~A302 & ~A301;
  assign \new_[42293]_  = \new_[42292]_  & \new_[42289]_ ;
  assign \new_[42294]_  = \new_[42293]_  & \new_[42286]_ ;
  assign \new_[42298]_  = ~A166 & ~A167;
  assign \new_[42299]_  = A170 & \new_[42298]_ ;
  assign \new_[42303]_  = ~A233 & A200;
  assign \new_[42304]_  = ~A199 & \new_[42303]_ ;
  assign \new_[42305]_  = \new_[42304]_  & \new_[42299]_ ;
  assign \new_[42309]_  = A265 & ~A236;
  assign \new_[42310]_  = ~A235 & \new_[42309]_ ;
  assign \new_[42313]_  = A298 & A266;
  assign \new_[42316]_  = ~A302 & ~A301;
  assign \new_[42317]_  = \new_[42316]_  & \new_[42313]_ ;
  assign \new_[42318]_  = \new_[42317]_  & \new_[42310]_ ;
  assign \new_[42322]_  = ~A166 & ~A167;
  assign \new_[42323]_  = A170 & \new_[42322]_ ;
  assign \new_[42327]_  = ~A233 & A200;
  assign \new_[42328]_  = ~A199 & \new_[42327]_ ;
  assign \new_[42329]_  = \new_[42328]_  & \new_[42323]_ ;
  assign \new_[42333]_  = ~A266 & ~A236;
  assign \new_[42334]_  = ~A235 & \new_[42333]_ ;
  assign \new_[42337]_  = ~A269 & ~A268;
  assign \new_[42340]_  = ~A300 & A298;
  assign \new_[42341]_  = \new_[42340]_  & \new_[42337]_ ;
  assign \new_[42342]_  = \new_[42341]_  & \new_[42334]_ ;
  assign \new_[42346]_  = ~A166 & ~A167;
  assign \new_[42347]_  = A170 & \new_[42346]_ ;
  assign \new_[42351]_  = ~A233 & A200;
  assign \new_[42352]_  = ~A199 & \new_[42351]_ ;
  assign \new_[42353]_  = \new_[42352]_  & \new_[42347]_ ;
  assign \new_[42357]_  = ~A266 & ~A236;
  assign \new_[42358]_  = ~A235 & \new_[42357]_ ;
  assign \new_[42361]_  = ~A269 & ~A268;
  assign \new_[42364]_  = A299 & A298;
  assign \new_[42365]_  = \new_[42364]_  & \new_[42361]_ ;
  assign \new_[42366]_  = \new_[42365]_  & \new_[42358]_ ;
  assign \new_[42370]_  = ~A166 & ~A167;
  assign \new_[42371]_  = A170 & \new_[42370]_ ;
  assign \new_[42375]_  = ~A233 & A200;
  assign \new_[42376]_  = ~A199 & \new_[42375]_ ;
  assign \new_[42377]_  = \new_[42376]_  & \new_[42371]_ ;
  assign \new_[42381]_  = ~A266 & ~A236;
  assign \new_[42382]_  = ~A235 & \new_[42381]_ ;
  assign \new_[42385]_  = ~A269 & ~A268;
  assign \new_[42388]_  = ~A299 & ~A298;
  assign \new_[42389]_  = \new_[42388]_  & \new_[42385]_ ;
  assign \new_[42390]_  = \new_[42389]_  & \new_[42382]_ ;
  assign \new_[42394]_  = ~A166 & ~A167;
  assign \new_[42395]_  = A170 & \new_[42394]_ ;
  assign \new_[42399]_  = ~A233 & A200;
  assign \new_[42400]_  = ~A199 & \new_[42399]_ ;
  assign \new_[42401]_  = \new_[42400]_  & \new_[42395]_ ;
  assign \new_[42405]_  = ~A266 & ~A236;
  assign \new_[42406]_  = ~A235 & \new_[42405]_ ;
  assign \new_[42409]_  = A298 & ~A267;
  assign \new_[42412]_  = ~A302 & ~A301;
  assign \new_[42413]_  = \new_[42412]_  & \new_[42409]_ ;
  assign \new_[42414]_  = \new_[42413]_  & \new_[42406]_ ;
  assign \new_[42418]_  = ~A166 & ~A167;
  assign \new_[42419]_  = A170 & \new_[42418]_ ;
  assign \new_[42423]_  = ~A233 & A200;
  assign \new_[42424]_  = ~A199 & \new_[42423]_ ;
  assign \new_[42425]_  = \new_[42424]_  & \new_[42419]_ ;
  assign \new_[42429]_  = ~A265 & ~A236;
  assign \new_[42430]_  = ~A235 & \new_[42429]_ ;
  assign \new_[42433]_  = A298 & ~A266;
  assign \new_[42436]_  = ~A302 & ~A301;
  assign \new_[42437]_  = \new_[42436]_  & \new_[42433]_ ;
  assign \new_[42438]_  = \new_[42437]_  & \new_[42430]_ ;
  assign \new_[42442]_  = ~A166 & ~A167;
  assign \new_[42443]_  = A170 & \new_[42442]_ ;
  assign \new_[42447]_  = ~A233 & A200;
  assign \new_[42448]_  = ~A199 & \new_[42447]_ ;
  assign \new_[42449]_  = \new_[42448]_  & \new_[42443]_ ;
  assign \new_[42453]_  = ~A268 & ~A266;
  assign \new_[42454]_  = ~A234 & \new_[42453]_ ;
  assign \new_[42457]_  = A298 & ~A269;
  assign \new_[42460]_  = ~A302 & ~A301;
  assign \new_[42461]_  = \new_[42460]_  & \new_[42457]_ ;
  assign \new_[42462]_  = \new_[42461]_  & \new_[42454]_ ;
  assign \new_[42466]_  = ~A166 & ~A167;
  assign \new_[42467]_  = A170 & \new_[42466]_ ;
  assign \new_[42471]_  = A232 & A200;
  assign \new_[42472]_  = ~A199 & \new_[42471]_ ;
  assign \new_[42473]_  = \new_[42472]_  & \new_[42467]_ ;
  assign \new_[42477]_  = A235 & A234;
  assign \new_[42478]_  = ~A233 & \new_[42477]_ ;
  assign \new_[42481]_  = ~A299 & A298;
  assign \new_[42484]_  = A301 & A300;
  assign \new_[42485]_  = \new_[42484]_  & \new_[42481]_ ;
  assign \new_[42486]_  = \new_[42485]_  & \new_[42478]_ ;
  assign \new_[42490]_  = ~A166 & ~A167;
  assign \new_[42491]_  = A170 & \new_[42490]_ ;
  assign \new_[42495]_  = A232 & A200;
  assign \new_[42496]_  = ~A199 & \new_[42495]_ ;
  assign \new_[42497]_  = \new_[42496]_  & \new_[42491]_ ;
  assign \new_[42501]_  = A235 & A234;
  assign \new_[42502]_  = ~A233 & \new_[42501]_ ;
  assign \new_[42505]_  = ~A299 & A298;
  assign \new_[42508]_  = A302 & A300;
  assign \new_[42509]_  = \new_[42508]_  & \new_[42505]_ ;
  assign \new_[42510]_  = \new_[42509]_  & \new_[42502]_ ;
  assign \new_[42514]_  = ~A166 & ~A167;
  assign \new_[42515]_  = A170 & \new_[42514]_ ;
  assign \new_[42519]_  = A232 & A200;
  assign \new_[42520]_  = ~A199 & \new_[42519]_ ;
  assign \new_[42521]_  = \new_[42520]_  & \new_[42515]_ ;
  assign \new_[42525]_  = A235 & A234;
  assign \new_[42526]_  = ~A233 & \new_[42525]_ ;
  assign \new_[42529]_  = ~A266 & A265;
  assign \new_[42532]_  = A268 & A267;
  assign \new_[42533]_  = \new_[42532]_  & \new_[42529]_ ;
  assign \new_[42534]_  = \new_[42533]_  & \new_[42526]_ ;
  assign \new_[42538]_  = ~A166 & ~A167;
  assign \new_[42539]_  = A170 & \new_[42538]_ ;
  assign \new_[42543]_  = A232 & A200;
  assign \new_[42544]_  = ~A199 & \new_[42543]_ ;
  assign \new_[42545]_  = \new_[42544]_  & \new_[42539]_ ;
  assign \new_[42549]_  = A235 & A234;
  assign \new_[42550]_  = ~A233 & \new_[42549]_ ;
  assign \new_[42553]_  = ~A266 & A265;
  assign \new_[42556]_  = A269 & A267;
  assign \new_[42557]_  = \new_[42556]_  & \new_[42553]_ ;
  assign \new_[42558]_  = \new_[42557]_  & \new_[42550]_ ;
  assign \new_[42562]_  = ~A166 & ~A167;
  assign \new_[42563]_  = A170 & \new_[42562]_ ;
  assign \new_[42567]_  = A232 & A200;
  assign \new_[42568]_  = ~A199 & \new_[42567]_ ;
  assign \new_[42569]_  = \new_[42568]_  & \new_[42563]_ ;
  assign \new_[42573]_  = A236 & A234;
  assign \new_[42574]_  = ~A233 & \new_[42573]_ ;
  assign \new_[42577]_  = ~A299 & A298;
  assign \new_[42580]_  = A301 & A300;
  assign \new_[42581]_  = \new_[42580]_  & \new_[42577]_ ;
  assign \new_[42582]_  = \new_[42581]_  & \new_[42574]_ ;
  assign \new_[42586]_  = ~A166 & ~A167;
  assign \new_[42587]_  = A170 & \new_[42586]_ ;
  assign \new_[42591]_  = A232 & A200;
  assign \new_[42592]_  = ~A199 & \new_[42591]_ ;
  assign \new_[42593]_  = \new_[42592]_  & \new_[42587]_ ;
  assign \new_[42597]_  = A236 & A234;
  assign \new_[42598]_  = ~A233 & \new_[42597]_ ;
  assign \new_[42601]_  = ~A299 & A298;
  assign \new_[42604]_  = A302 & A300;
  assign \new_[42605]_  = \new_[42604]_  & \new_[42601]_ ;
  assign \new_[42606]_  = \new_[42605]_  & \new_[42598]_ ;
  assign \new_[42610]_  = ~A166 & ~A167;
  assign \new_[42611]_  = A170 & \new_[42610]_ ;
  assign \new_[42615]_  = A232 & A200;
  assign \new_[42616]_  = ~A199 & \new_[42615]_ ;
  assign \new_[42617]_  = \new_[42616]_  & \new_[42611]_ ;
  assign \new_[42621]_  = A236 & A234;
  assign \new_[42622]_  = ~A233 & \new_[42621]_ ;
  assign \new_[42625]_  = ~A266 & A265;
  assign \new_[42628]_  = A268 & A267;
  assign \new_[42629]_  = \new_[42628]_  & \new_[42625]_ ;
  assign \new_[42630]_  = \new_[42629]_  & \new_[42622]_ ;
  assign \new_[42634]_  = ~A166 & ~A167;
  assign \new_[42635]_  = A170 & \new_[42634]_ ;
  assign \new_[42639]_  = A232 & A200;
  assign \new_[42640]_  = ~A199 & \new_[42639]_ ;
  assign \new_[42641]_  = \new_[42640]_  & \new_[42635]_ ;
  assign \new_[42645]_  = A236 & A234;
  assign \new_[42646]_  = ~A233 & \new_[42645]_ ;
  assign \new_[42649]_  = ~A266 & A265;
  assign \new_[42652]_  = A269 & A267;
  assign \new_[42653]_  = \new_[42652]_  & \new_[42649]_ ;
  assign \new_[42654]_  = \new_[42653]_  & \new_[42646]_ ;
  assign \new_[42658]_  = ~A166 & ~A167;
  assign \new_[42659]_  = A170 & \new_[42658]_ ;
  assign \new_[42663]_  = ~A232 & A200;
  assign \new_[42664]_  = ~A199 & \new_[42663]_ ;
  assign \new_[42665]_  = \new_[42664]_  & \new_[42659]_ ;
  assign \new_[42669]_  = ~A268 & ~A266;
  assign \new_[42670]_  = ~A233 & \new_[42669]_ ;
  assign \new_[42673]_  = A298 & ~A269;
  assign \new_[42676]_  = ~A302 & ~A301;
  assign \new_[42677]_  = \new_[42676]_  & \new_[42673]_ ;
  assign \new_[42678]_  = \new_[42677]_  & \new_[42670]_ ;
  assign \new_[42682]_  = ~A166 & ~A167;
  assign \new_[42683]_  = A170 & \new_[42682]_ ;
  assign \new_[42687]_  = A201 & ~A200;
  assign \new_[42688]_  = A199 & \new_[42687]_ ;
  assign \new_[42689]_  = \new_[42688]_  & \new_[42683]_ ;
  assign \new_[42693]_  = A233 & A232;
  assign \new_[42694]_  = A202 & \new_[42693]_ ;
  assign \new_[42697]_  = ~A267 & A265;
  assign \new_[42700]_  = ~A300 & ~A299;
  assign \new_[42701]_  = \new_[42700]_  & \new_[42697]_ ;
  assign \new_[42702]_  = \new_[42701]_  & \new_[42694]_ ;
  assign \new_[42706]_  = ~A166 & ~A167;
  assign \new_[42707]_  = A170 & \new_[42706]_ ;
  assign \new_[42711]_  = A201 & ~A200;
  assign \new_[42712]_  = A199 & \new_[42711]_ ;
  assign \new_[42713]_  = \new_[42712]_  & \new_[42707]_ ;
  assign \new_[42717]_  = A233 & A232;
  assign \new_[42718]_  = A202 & \new_[42717]_ ;
  assign \new_[42721]_  = ~A267 & A265;
  assign \new_[42724]_  = A299 & A298;
  assign \new_[42725]_  = \new_[42724]_  & \new_[42721]_ ;
  assign \new_[42726]_  = \new_[42725]_  & \new_[42718]_ ;
  assign \new_[42730]_  = ~A166 & ~A167;
  assign \new_[42731]_  = A170 & \new_[42730]_ ;
  assign \new_[42735]_  = A201 & ~A200;
  assign \new_[42736]_  = A199 & \new_[42735]_ ;
  assign \new_[42737]_  = \new_[42736]_  & \new_[42731]_ ;
  assign \new_[42741]_  = A233 & A232;
  assign \new_[42742]_  = A202 & \new_[42741]_ ;
  assign \new_[42745]_  = ~A267 & A265;
  assign \new_[42748]_  = ~A299 & ~A298;
  assign \new_[42749]_  = \new_[42748]_  & \new_[42745]_ ;
  assign \new_[42750]_  = \new_[42749]_  & \new_[42742]_ ;
  assign \new_[42754]_  = ~A166 & ~A167;
  assign \new_[42755]_  = A170 & \new_[42754]_ ;
  assign \new_[42759]_  = A201 & ~A200;
  assign \new_[42760]_  = A199 & \new_[42759]_ ;
  assign \new_[42761]_  = \new_[42760]_  & \new_[42755]_ ;
  assign \new_[42765]_  = A233 & A232;
  assign \new_[42766]_  = A202 & \new_[42765]_ ;
  assign \new_[42769]_  = A266 & A265;
  assign \new_[42772]_  = ~A300 & ~A299;
  assign \new_[42773]_  = \new_[42772]_  & \new_[42769]_ ;
  assign \new_[42774]_  = \new_[42773]_  & \new_[42766]_ ;
  assign \new_[42778]_  = ~A166 & ~A167;
  assign \new_[42779]_  = A170 & \new_[42778]_ ;
  assign \new_[42783]_  = A201 & ~A200;
  assign \new_[42784]_  = A199 & \new_[42783]_ ;
  assign \new_[42785]_  = \new_[42784]_  & \new_[42779]_ ;
  assign \new_[42789]_  = A233 & A232;
  assign \new_[42790]_  = A202 & \new_[42789]_ ;
  assign \new_[42793]_  = A266 & A265;
  assign \new_[42796]_  = A299 & A298;
  assign \new_[42797]_  = \new_[42796]_  & \new_[42793]_ ;
  assign \new_[42798]_  = \new_[42797]_  & \new_[42790]_ ;
  assign \new_[42802]_  = ~A166 & ~A167;
  assign \new_[42803]_  = A170 & \new_[42802]_ ;
  assign \new_[42807]_  = A201 & ~A200;
  assign \new_[42808]_  = A199 & \new_[42807]_ ;
  assign \new_[42809]_  = \new_[42808]_  & \new_[42803]_ ;
  assign \new_[42813]_  = A233 & A232;
  assign \new_[42814]_  = A202 & \new_[42813]_ ;
  assign \new_[42817]_  = A266 & A265;
  assign \new_[42820]_  = ~A299 & ~A298;
  assign \new_[42821]_  = \new_[42820]_  & \new_[42817]_ ;
  assign \new_[42822]_  = \new_[42821]_  & \new_[42814]_ ;
  assign \new_[42826]_  = ~A166 & ~A167;
  assign \new_[42827]_  = A170 & \new_[42826]_ ;
  assign \new_[42831]_  = A201 & ~A200;
  assign \new_[42832]_  = A199 & \new_[42831]_ ;
  assign \new_[42833]_  = \new_[42832]_  & \new_[42827]_ ;
  assign \new_[42837]_  = A233 & A232;
  assign \new_[42838]_  = A202 & \new_[42837]_ ;
  assign \new_[42841]_  = ~A266 & ~A265;
  assign \new_[42844]_  = ~A300 & ~A299;
  assign \new_[42845]_  = \new_[42844]_  & \new_[42841]_ ;
  assign \new_[42846]_  = \new_[42845]_  & \new_[42838]_ ;
  assign \new_[42850]_  = ~A166 & ~A167;
  assign \new_[42851]_  = A170 & \new_[42850]_ ;
  assign \new_[42855]_  = A201 & ~A200;
  assign \new_[42856]_  = A199 & \new_[42855]_ ;
  assign \new_[42857]_  = \new_[42856]_  & \new_[42851]_ ;
  assign \new_[42861]_  = A233 & A232;
  assign \new_[42862]_  = A202 & \new_[42861]_ ;
  assign \new_[42865]_  = ~A266 & ~A265;
  assign \new_[42868]_  = A299 & A298;
  assign \new_[42869]_  = \new_[42868]_  & \new_[42865]_ ;
  assign \new_[42870]_  = \new_[42869]_  & \new_[42862]_ ;
  assign \new_[42874]_  = ~A166 & ~A167;
  assign \new_[42875]_  = A170 & \new_[42874]_ ;
  assign \new_[42879]_  = A201 & ~A200;
  assign \new_[42880]_  = A199 & \new_[42879]_ ;
  assign \new_[42881]_  = \new_[42880]_  & \new_[42875]_ ;
  assign \new_[42885]_  = A233 & A232;
  assign \new_[42886]_  = A202 & \new_[42885]_ ;
  assign \new_[42889]_  = ~A266 & ~A265;
  assign \new_[42892]_  = ~A299 & ~A298;
  assign \new_[42893]_  = \new_[42892]_  & \new_[42889]_ ;
  assign \new_[42894]_  = \new_[42893]_  & \new_[42886]_ ;
  assign \new_[42898]_  = ~A166 & ~A167;
  assign \new_[42899]_  = A170 & \new_[42898]_ ;
  assign \new_[42903]_  = A201 & ~A200;
  assign \new_[42904]_  = A199 & \new_[42903]_ ;
  assign \new_[42905]_  = \new_[42904]_  & \new_[42899]_ ;
  assign \new_[42909]_  = A233 & ~A232;
  assign \new_[42910]_  = A202 & \new_[42909]_ ;
  assign \new_[42913]_  = ~A299 & A298;
  assign \new_[42916]_  = A301 & A300;
  assign \new_[42917]_  = \new_[42916]_  & \new_[42913]_ ;
  assign \new_[42918]_  = \new_[42917]_  & \new_[42910]_ ;
  assign \new_[42922]_  = ~A166 & ~A167;
  assign \new_[42923]_  = A170 & \new_[42922]_ ;
  assign \new_[42927]_  = A201 & ~A200;
  assign \new_[42928]_  = A199 & \new_[42927]_ ;
  assign \new_[42929]_  = \new_[42928]_  & \new_[42923]_ ;
  assign \new_[42933]_  = A233 & ~A232;
  assign \new_[42934]_  = A202 & \new_[42933]_ ;
  assign \new_[42937]_  = ~A299 & A298;
  assign \new_[42940]_  = A302 & A300;
  assign \new_[42941]_  = \new_[42940]_  & \new_[42937]_ ;
  assign \new_[42942]_  = \new_[42941]_  & \new_[42934]_ ;
  assign \new_[42946]_  = ~A166 & ~A167;
  assign \new_[42947]_  = A170 & \new_[42946]_ ;
  assign \new_[42951]_  = A201 & ~A200;
  assign \new_[42952]_  = A199 & \new_[42951]_ ;
  assign \new_[42953]_  = \new_[42952]_  & \new_[42947]_ ;
  assign \new_[42957]_  = A233 & ~A232;
  assign \new_[42958]_  = A202 & \new_[42957]_ ;
  assign \new_[42961]_  = ~A266 & A265;
  assign \new_[42964]_  = A268 & A267;
  assign \new_[42965]_  = \new_[42964]_  & \new_[42961]_ ;
  assign \new_[42966]_  = \new_[42965]_  & \new_[42958]_ ;
  assign \new_[42970]_  = ~A166 & ~A167;
  assign \new_[42971]_  = A170 & \new_[42970]_ ;
  assign \new_[42975]_  = A201 & ~A200;
  assign \new_[42976]_  = A199 & \new_[42975]_ ;
  assign \new_[42977]_  = \new_[42976]_  & \new_[42971]_ ;
  assign \new_[42981]_  = A233 & ~A232;
  assign \new_[42982]_  = A202 & \new_[42981]_ ;
  assign \new_[42985]_  = ~A266 & A265;
  assign \new_[42988]_  = A269 & A267;
  assign \new_[42989]_  = \new_[42988]_  & \new_[42985]_ ;
  assign \new_[42990]_  = \new_[42989]_  & \new_[42982]_ ;
  assign \new_[42994]_  = ~A166 & ~A167;
  assign \new_[42995]_  = A170 & \new_[42994]_ ;
  assign \new_[42999]_  = A201 & ~A200;
  assign \new_[43000]_  = A199 & \new_[42999]_ ;
  assign \new_[43001]_  = \new_[43000]_  & \new_[42995]_ ;
  assign \new_[43005]_  = ~A234 & ~A233;
  assign \new_[43006]_  = A202 & \new_[43005]_ ;
  assign \new_[43009]_  = A266 & A265;
  assign \new_[43012]_  = ~A300 & A298;
  assign \new_[43013]_  = \new_[43012]_  & \new_[43009]_ ;
  assign \new_[43014]_  = \new_[43013]_  & \new_[43006]_ ;
  assign \new_[43018]_  = ~A166 & ~A167;
  assign \new_[43019]_  = A170 & \new_[43018]_ ;
  assign \new_[43023]_  = A201 & ~A200;
  assign \new_[43024]_  = A199 & \new_[43023]_ ;
  assign \new_[43025]_  = \new_[43024]_  & \new_[43019]_ ;
  assign \new_[43029]_  = ~A234 & ~A233;
  assign \new_[43030]_  = A202 & \new_[43029]_ ;
  assign \new_[43033]_  = A266 & A265;
  assign \new_[43036]_  = A299 & A298;
  assign \new_[43037]_  = \new_[43036]_  & \new_[43033]_ ;
  assign \new_[43038]_  = \new_[43037]_  & \new_[43030]_ ;
  assign \new_[43042]_  = ~A166 & ~A167;
  assign \new_[43043]_  = A170 & \new_[43042]_ ;
  assign \new_[43047]_  = A201 & ~A200;
  assign \new_[43048]_  = A199 & \new_[43047]_ ;
  assign \new_[43049]_  = \new_[43048]_  & \new_[43043]_ ;
  assign \new_[43053]_  = ~A234 & ~A233;
  assign \new_[43054]_  = A202 & \new_[43053]_ ;
  assign \new_[43057]_  = A266 & A265;
  assign \new_[43060]_  = ~A299 & ~A298;
  assign \new_[43061]_  = \new_[43060]_  & \new_[43057]_ ;
  assign \new_[43062]_  = \new_[43061]_  & \new_[43054]_ ;
  assign \new_[43066]_  = ~A166 & ~A167;
  assign \new_[43067]_  = A170 & \new_[43066]_ ;
  assign \new_[43071]_  = A201 & ~A200;
  assign \new_[43072]_  = A199 & \new_[43071]_ ;
  assign \new_[43073]_  = \new_[43072]_  & \new_[43067]_ ;
  assign \new_[43077]_  = ~A234 & ~A233;
  assign \new_[43078]_  = A202 & \new_[43077]_ ;
  assign \new_[43081]_  = ~A267 & ~A266;
  assign \new_[43084]_  = ~A300 & A298;
  assign \new_[43085]_  = \new_[43084]_  & \new_[43081]_ ;
  assign \new_[43086]_  = \new_[43085]_  & \new_[43078]_ ;
  assign \new_[43090]_  = ~A166 & ~A167;
  assign \new_[43091]_  = A170 & \new_[43090]_ ;
  assign \new_[43095]_  = A201 & ~A200;
  assign \new_[43096]_  = A199 & \new_[43095]_ ;
  assign \new_[43097]_  = \new_[43096]_  & \new_[43091]_ ;
  assign \new_[43101]_  = ~A234 & ~A233;
  assign \new_[43102]_  = A202 & \new_[43101]_ ;
  assign \new_[43105]_  = ~A267 & ~A266;
  assign \new_[43108]_  = A299 & A298;
  assign \new_[43109]_  = \new_[43108]_  & \new_[43105]_ ;
  assign \new_[43110]_  = \new_[43109]_  & \new_[43102]_ ;
  assign \new_[43114]_  = ~A166 & ~A167;
  assign \new_[43115]_  = A170 & \new_[43114]_ ;
  assign \new_[43119]_  = A201 & ~A200;
  assign \new_[43120]_  = A199 & \new_[43119]_ ;
  assign \new_[43121]_  = \new_[43120]_  & \new_[43115]_ ;
  assign \new_[43125]_  = ~A234 & ~A233;
  assign \new_[43126]_  = A202 & \new_[43125]_ ;
  assign \new_[43129]_  = ~A267 & ~A266;
  assign \new_[43132]_  = ~A299 & ~A298;
  assign \new_[43133]_  = \new_[43132]_  & \new_[43129]_ ;
  assign \new_[43134]_  = \new_[43133]_  & \new_[43126]_ ;
  assign \new_[43138]_  = ~A166 & ~A167;
  assign \new_[43139]_  = A170 & \new_[43138]_ ;
  assign \new_[43143]_  = A201 & ~A200;
  assign \new_[43144]_  = A199 & \new_[43143]_ ;
  assign \new_[43145]_  = \new_[43144]_  & \new_[43139]_ ;
  assign \new_[43149]_  = ~A234 & ~A233;
  assign \new_[43150]_  = A202 & \new_[43149]_ ;
  assign \new_[43153]_  = ~A266 & ~A265;
  assign \new_[43156]_  = ~A300 & A298;
  assign \new_[43157]_  = \new_[43156]_  & \new_[43153]_ ;
  assign \new_[43158]_  = \new_[43157]_  & \new_[43150]_ ;
  assign \new_[43162]_  = ~A166 & ~A167;
  assign \new_[43163]_  = A170 & \new_[43162]_ ;
  assign \new_[43167]_  = A201 & ~A200;
  assign \new_[43168]_  = A199 & \new_[43167]_ ;
  assign \new_[43169]_  = \new_[43168]_  & \new_[43163]_ ;
  assign \new_[43173]_  = ~A234 & ~A233;
  assign \new_[43174]_  = A202 & \new_[43173]_ ;
  assign \new_[43177]_  = ~A266 & ~A265;
  assign \new_[43180]_  = A299 & A298;
  assign \new_[43181]_  = \new_[43180]_  & \new_[43177]_ ;
  assign \new_[43182]_  = \new_[43181]_  & \new_[43174]_ ;
  assign \new_[43186]_  = ~A166 & ~A167;
  assign \new_[43187]_  = A170 & \new_[43186]_ ;
  assign \new_[43191]_  = A201 & ~A200;
  assign \new_[43192]_  = A199 & \new_[43191]_ ;
  assign \new_[43193]_  = \new_[43192]_  & \new_[43187]_ ;
  assign \new_[43197]_  = ~A234 & ~A233;
  assign \new_[43198]_  = A202 & \new_[43197]_ ;
  assign \new_[43201]_  = ~A266 & ~A265;
  assign \new_[43204]_  = ~A299 & ~A298;
  assign \new_[43205]_  = \new_[43204]_  & \new_[43201]_ ;
  assign \new_[43206]_  = \new_[43205]_  & \new_[43198]_ ;
  assign \new_[43210]_  = ~A166 & ~A167;
  assign \new_[43211]_  = A170 & \new_[43210]_ ;
  assign \new_[43215]_  = A201 & ~A200;
  assign \new_[43216]_  = A199 & \new_[43215]_ ;
  assign \new_[43217]_  = \new_[43216]_  & \new_[43211]_ ;
  assign \new_[43221]_  = ~A233 & A232;
  assign \new_[43222]_  = A202 & \new_[43221]_ ;
  assign \new_[43225]_  = A235 & A234;
  assign \new_[43228]_  = A299 & ~A298;
  assign \new_[43229]_  = \new_[43228]_  & \new_[43225]_ ;
  assign \new_[43230]_  = \new_[43229]_  & \new_[43222]_ ;
  assign \new_[43234]_  = ~A166 & ~A167;
  assign \new_[43235]_  = A170 & \new_[43234]_ ;
  assign \new_[43239]_  = A201 & ~A200;
  assign \new_[43240]_  = A199 & \new_[43239]_ ;
  assign \new_[43241]_  = \new_[43240]_  & \new_[43235]_ ;
  assign \new_[43245]_  = ~A233 & A232;
  assign \new_[43246]_  = A202 & \new_[43245]_ ;
  assign \new_[43249]_  = A235 & A234;
  assign \new_[43252]_  = A266 & ~A265;
  assign \new_[43253]_  = \new_[43252]_  & \new_[43249]_ ;
  assign \new_[43254]_  = \new_[43253]_  & \new_[43246]_ ;
  assign \new_[43258]_  = ~A166 & ~A167;
  assign \new_[43259]_  = A170 & \new_[43258]_ ;
  assign \new_[43263]_  = A201 & ~A200;
  assign \new_[43264]_  = A199 & \new_[43263]_ ;
  assign \new_[43265]_  = \new_[43264]_  & \new_[43259]_ ;
  assign \new_[43269]_  = ~A233 & A232;
  assign \new_[43270]_  = A202 & \new_[43269]_ ;
  assign \new_[43273]_  = A236 & A234;
  assign \new_[43276]_  = A299 & ~A298;
  assign \new_[43277]_  = \new_[43276]_  & \new_[43273]_ ;
  assign \new_[43278]_  = \new_[43277]_  & \new_[43270]_ ;
  assign \new_[43282]_  = ~A166 & ~A167;
  assign \new_[43283]_  = A170 & \new_[43282]_ ;
  assign \new_[43287]_  = A201 & ~A200;
  assign \new_[43288]_  = A199 & \new_[43287]_ ;
  assign \new_[43289]_  = \new_[43288]_  & \new_[43283]_ ;
  assign \new_[43293]_  = ~A233 & A232;
  assign \new_[43294]_  = A202 & \new_[43293]_ ;
  assign \new_[43297]_  = A236 & A234;
  assign \new_[43300]_  = A266 & ~A265;
  assign \new_[43301]_  = \new_[43300]_  & \new_[43297]_ ;
  assign \new_[43302]_  = \new_[43301]_  & \new_[43294]_ ;
  assign \new_[43306]_  = ~A166 & ~A167;
  assign \new_[43307]_  = A170 & \new_[43306]_ ;
  assign \new_[43311]_  = A201 & ~A200;
  assign \new_[43312]_  = A199 & \new_[43311]_ ;
  assign \new_[43313]_  = \new_[43312]_  & \new_[43307]_ ;
  assign \new_[43317]_  = ~A233 & ~A232;
  assign \new_[43318]_  = A202 & \new_[43317]_ ;
  assign \new_[43321]_  = A266 & A265;
  assign \new_[43324]_  = ~A300 & A298;
  assign \new_[43325]_  = \new_[43324]_  & \new_[43321]_ ;
  assign \new_[43326]_  = \new_[43325]_  & \new_[43318]_ ;
  assign \new_[43330]_  = ~A166 & ~A167;
  assign \new_[43331]_  = A170 & \new_[43330]_ ;
  assign \new_[43335]_  = A201 & ~A200;
  assign \new_[43336]_  = A199 & \new_[43335]_ ;
  assign \new_[43337]_  = \new_[43336]_  & \new_[43331]_ ;
  assign \new_[43341]_  = ~A233 & ~A232;
  assign \new_[43342]_  = A202 & \new_[43341]_ ;
  assign \new_[43345]_  = A266 & A265;
  assign \new_[43348]_  = A299 & A298;
  assign \new_[43349]_  = \new_[43348]_  & \new_[43345]_ ;
  assign \new_[43350]_  = \new_[43349]_  & \new_[43342]_ ;
  assign \new_[43354]_  = ~A166 & ~A167;
  assign \new_[43355]_  = A170 & \new_[43354]_ ;
  assign \new_[43359]_  = A201 & ~A200;
  assign \new_[43360]_  = A199 & \new_[43359]_ ;
  assign \new_[43361]_  = \new_[43360]_  & \new_[43355]_ ;
  assign \new_[43365]_  = ~A233 & ~A232;
  assign \new_[43366]_  = A202 & \new_[43365]_ ;
  assign \new_[43369]_  = A266 & A265;
  assign \new_[43372]_  = ~A299 & ~A298;
  assign \new_[43373]_  = \new_[43372]_  & \new_[43369]_ ;
  assign \new_[43374]_  = \new_[43373]_  & \new_[43366]_ ;
  assign \new_[43378]_  = ~A166 & ~A167;
  assign \new_[43379]_  = A170 & \new_[43378]_ ;
  assign \new_[43383]_  = A201 & ~A200;
  assign \new_[43384]_  = A199 & \new_[43383]_ ;
  assign \new_[43385]_  = \new_[43384]_  & \new_[43379]_ ;
  assign \new_[43389]_  = ~A233 & ~A232;
  assign \new_[43390]_  = A202 & \new_[43389]_ ;
  assign \new_[43393]_  = ~A267 & ~A266;
  assign \new_[43396]_  = ~A300 & A298;
  assign \new_[43397]_  = \new_[43396]_  & \new_[43393]_ ;
  assign \new_[43398]_  = \new_[43397]_  & \new_[43390]_ ;
  assign \new_[43402]_  = ~A166 & ~A167;
  assign \new_[43403]_  = A170 & \new_[43402]_ ;
  assign \new_[43407]_  = A201 & ~A200;
  assign \new_[43408]_  = A199 & \new_[43407]_ ;
  assign \new_[43409]_  = \new_[43408]_  & \new_[43403]_ ;
  assign \new_[43413]_  = ~A233 & ~A232;
  assign \new_[43414]_  = A202 & \new_[43413]_ ;
  assign \new_[43417]_  = ~A267 & ~A266;
  assign \new_[43420]_  = A299 & A298;
  assign \new_[43421]_  = \new_[43420]_  & \new_[43417]_ ;
  assign \new_[43422]_  = \new_[43421]_  & \new_[43414]_ ;
  assign \new_[43426]_  = ~A166 & ~A167;
  assign \new_[43427]_  = A170 & \new_[43426]_ ;
  assign \new_[43431]_  = A201 & ~A200;
  assign \new_[43432]_  = A199 & \new_[43431]_ ;
  assign \new_[43433]_  = \new_[43432]_  & \new_[43427]_ ;
  assign \new_[43437]_  = ~A233 & ~A232;
  assign \new_[43438]_  = A202 & \new_[43437]_ ;
  assign \new_[43441]_  = ~A267 & ~A266;
  assign \new_[43444]_  = ~A299 & ~A298;
  assign \new_[43445]_  = \new_[43444]_  & \new_[43441]_ ;
  assign \new_[43446]_  = \new_[43445]_  & \new_[43438]_ ;
  assign \new_[43450]_  = ~A166 & ~A167;
  assign \new_[43451]_  = A170 & \new_[43450]_ ;
  assign \new_[43455]_  = A201 & ~A200;
  assign \new_[43456]_  = A199 & \new_[43455]_ ;
  assign \new_[43457]_  = \new_[43456]_  & \new_[43451]_ ;
  assign \new_[43461]_  = ~A233 & ~A232;
  assign \new_[43462]_  = A202 & \new_[43461]_ ;
  assign \new_[43465]_  = ~A266 & ~A265;
  assign \new_[43468]_  = ~A300 & A298;
  assign \new_[43469]_  = \new_[43468]_  & \new_[43465]_ ;
  assign \new_[43470]_  = \new_[43469]_  & \new_[43462]_ ;
  assign \new_[43474]_  = ~A166 & ~A167;
  assign \new_[43475]_  = A170 & \new_[43474]_ ;
  assign \new_[43479]_  = A201 & ~A200;
  assign \new_[43480]_  = A199 & \new_[43479]_ ;
  assign \new_[43481]_  = \new_[43480]_  & \new_[43475]_ ;
  assign \new_[43485]_  = ~A233 & ~A232;
  assign \new_[43486]_  = A202 & \new_[43485]_ ;
  assign \new_[43489]_  = ~A266 & ~A265;
  assign \new_[43492]_  = A299 & A298;
  assign \new_[43493]_  = \new_[43492]_  & \new_[43489]_ ;
  assign \new_[43494]_  = \new_[43493]_  & \new_[43486]_ ;
  assign \new_[43498]_  = ~A166 & ~A167;
  assign \new_[43499]_  = A170 & \new_[43498]_ ;
  assign \new_[43503]_  = A201 & ~A200;
  assign \new_[43504]_  = A199 & \new_[43503]_ ;
  assign \new_[43505]_  = \new_[43504]_  & \new_[43499]_ ;
  assign \new_[43509]_  = ~A233 & ~A232;
  assign \new_[43510]_  = A202 & \new_[43509]_ ;
  assign \new_[43513]_  = ~A266 & ~A265;
  assign \new_[43516]_  = ~A299 & ~A298;
  assign \new_[43517]_  = \new_[43516]_  & \new_[43513]_ ;
  assign \new_[43518]_  = \new_[43517]_  & \new_[43510]_ ;
  assign \new_[43522]_  = ~A166 & ~A167;
  assign \new_[43523]_  = A170 & \new_[43522]_ ;
  assign \new_[43527]_  = A201 & ~A200;
  assign \new_[43528]_  = A199 & \new_[43527]_ ;
  assign \new_[43529]_  = \new_[43528]_  & \new_[43523]_ ;
  assign \new_[43533]_  = A233 & A232;
  assign \new_[43534]_  = A203 & \new_[43533]_ ;
  assign \new_[43537]_  = ~A267 & A265;
  assign \new_[43540]_  = ~A300 & ~A299;
  assign \new_[43541]_  = \new_[43540]_  & \new_[43537]_ ;
  assign \new_[43542]_  = \new_[43541]_  & \new_[43534]_ ;
  assign \new_[43546]_  = ~A166 & ~A167;
  assign \new_[43547]_  = A170 & \new_[43546]_ ;
  assign \new_[43551]_  = A201 & ~A200;
  assign \new_[43552]_  = A199 & \new_[43551]_ ;
  assign \new_[43553]_  = \new_[43552]_  & \new_[43547]_ ;
  assign \new_[43557]_  = A233 & A232;
  assign \new_[43558]_  = A203 & \new_[43557]_ ;
  assign \new_[43561]_  = ~A267 & A265;
  assign \new_[43564]_  = A299 & A298;
  assign \new_[43565]_  = \new_[43564]_  & \new_[43561]_ ;
  assign \new_[43566]_  = \new_[43565]_  & \new_[43558]_ ;
  assign \new_[43570]_  = ~A166 & ~A167;
  assign \new_[43571]_  = A170 & \new_[43570]_ ;
  assign \new_[43575]_  = A201 & ~A200;
  assign \new_[43576]_  = A199 & \new_[43575]_ ;
  assign \new_[43577]_  = \new_[43576]_  & \new_[43571]_ ;
  assign \new_[43581]_  = A233 & A232;
  assign \new_[43582]_  = A203 & \new_[43581]_ ;
  assign \new_[43585]_  = ~A267 & A265;
  assign \new_[43588]_  = ~A299 & ~A298;
  assign \new_[43589]_  = \new_[43588]_  & \new_[43585]_ ;
  assign \new_[43590]_  = \new_[43589]_  & \new_[43582]_ ;
  assign \new_[43594]_  = ~A166 & ~A167;
  assign \new_[43595]_  = A170 & \new_[43594]_ ;
  assign \new_[43599]_  = A201 & ~A200;
  assign \new_[43600]_  = A199 & \new_[43599]_ ;
  assign \new_[43601]_  = \new_[43600]_  & \new_[43595]_ ;
  assign \new_[43605]_  = A233 & A232;
  assign \new_[43606]_  = A203 & \new_[43605]_ ;
  assign \new_[43609]_  = A266 & A265;
  assign \new_[43612]_  = ~A300 & ~A299;
  assign \new_[43613]_  = \new_[43612]_  & \new_[43609]_ ;
  assign \new_[43614]_  = \new_[43613]_  & \new_[43606]_ ;
  assign \new_[43618]_  = ~A166 & ~A167;
  assign \new_[43619]_  = A170 & \new_[43618]_ ;
  assign \new_[43623]_  = A201 & ~A200;
  assign \new_[43624]_  = A199 & \new_[43623]_ ;
  assign \new_[43625]_  = \new_[43624]_  & \new_[43619]_ ;
  assign \new_[43629]_  = A233 & A232;
  assign \new_[43630]_  = A203 & \new_[43629]_ ;
  assign \new_[43633]_  = A266 & A265;
  assign \new_[43636]_  = A299 & A298;
  assign \new_[43637]_  = \new_[43636]_  & \new_[43633]_ ;
  assign \new_[43638]_  = \new_[43637]_  & \new_[43630]_ ;
  assign \new_[43642]_  = ~A166 & ~A167;
  assign \new_[43643]_  = A170 & \new_[43642]_ ;
  assign \new_[43647]_  = A201 & ~A200;
  assign \new_[43648]_  = A199 & \new_[43647]_ ;
  assign \new_[43649]_  = \new_[43648]_  & \new_[43643]_ ;
  assign \new_[43653]_  = A233 & A232;
  assign \new_[43654]_  = A203 & \new_[43653]_ ;
  assign \new_[43657]_  = A266 & A265;
  assign \new_[43660]_  = ~A299 & ~A298;
  assign \new_[43661]_  = \new_[43660]_  & \new_[43657]_ ;
  assign \new_[43662]_  = \new_[43661]_  & \new_[43654]_ ;
  assign \new_[43666]_  = ~A166 & ~A167;
  assign \new_[43667]_  = A170 & \new_[43666]_ ;
  assign \new_[43671]_  = A201 & ~A200;
  assign \new_[43672]_  = A199 & \new_[43671]_ ;
  assign \new_[43673]_  = \new_[43672]_  & \new_[43667]_ ;
  assign \new_[43677]_  = A233 & A232;
  assign \new_[43678]_  = A203 & \new_[43677]_ ;
  assign \new_[43681]_  = ~A266 & ~A265;
  assign \new_[43684]_  = ~A300 & ~A299;
  assign \new_[43685]_  = \new_[43684]_  & \new_[43681]_ ;
  assign \new_[43686]_  = \new_[43685]_  & \new_[43678]_ ;
  assign \new_[43690]_  = ~A166 & ~A167;
  assign \new_[43691]_  = A170 & \new_[43690]_ ;
  assign \new_[43695]_  = A201 & ~A200;
  assign \new_[43696]_  = A199 & \new_[43695]_ ;
  assign \new_[43697]_  = \new_[43696]_  & \new_[43691]_ ;
  assign \new_[43701]_  = A233 & A232;
  assign \new_[43702]_  = A203 & \new_[43701]_ ;
  assign \new_[43705]_  = ~A266 & ~A265;
  assign \new_[43708]_  = A299 & A298;
  assign \new_[43709]_  = \new_[43708]_  & \new_[43705]_ ;
  assign \new_[43710]_  = \new_[43709]_  & \new_[43702]_ ;
  assign \new_[43714]_  = ~A166 & ~A167;
  assign \new_[43715]_  = A170 & \new_[43714]_ ;
  assign \new_[43719]_  = A201 & ~A200;
  assign \new_[43720]_  = A199 & \new_[43719]_ ;
  assign \new_[43721]_  = \new_[43720]_  & \new_[43715]_ ;
  assign \new_[43725]_  = A233 & A232;
  assign \new_[43726]_  = A203 & \new_[43725]_ ;
  assign \new_[43729]_  = ~A266 & ~A265;
  assign \new_[43732]_  = ~A299 & ~A298;
  assign \new_[43733]_  = \new_[43732]_  & \new_[43729]_ ;
  assign \new_[43734]_  = \new_[43733]_  & \new_[43726]_ ;
  assign \new_[43738]_  = ~A166 & ~A167;
  assign \new_[43739]_  = A170 & \new_[43738]_ ;
  assign \new_[43743]_  = A201 & ~A200;
  assign \new_[43744]_  = A199 & \new_[43743]_ ;
  assign \new_[43745]_  = \new_[43744]_  & \new_[43739]_ ;
  assign \new_[43749]_  = A233 & ~A232;
  assign \new_[43750]_  = A203 & \new_[43749]_ ;
  assign \new_[43753]_  = ~A299 & A298;
  assign \new_[43756]_  = A301 & A300;
  assign \new_[43757]_  = \new_[43756]_  & \new_[43753]_ ;
  assign \new_[43758]_  = \new_[43757]_  & \new_[43750]_ ;
  assign \new_[43762]_  = ~A166 & ~A167;
  assign \new_[43763]_  = A170 & \new_[43762]_ ;
  assign \new_[43767]_  = A201 & ~A200;
  assign \new_[43768]_  = A199 & \new_[43767]_ ;
  assign \new_[43769]_  = \new_[43768]_  & \new_[43763]_ ;
  assign \new_[43773]_  = A233 & ~A232;
  assign \new_[43774]_  = A203 & \new_[43773]_ ;
  assign \new_[43777]_  = ~A299 & A298;
  assign \new_[43780]_  = A302 & A300;
  assign \new_[43781]_  = \new_[43780]_  & \new_[43777]_ ;
  assign \new_[43782]_  = \new_[43781]_  & \new_[43774]_ ;
  assign \new_[43786]_  = ~A166 & ~A167;
  assign \new_[43787]_  = A170 & \new_[43786]_ ;
  assign \new_[43791]_  = A201 & ~A200;
  assign \new_[43792]_  = A199 & \new_[43791]_ ;
  assign \new_[43793]_  = \new_[43792]_  & \new_[43787]_ ;
  assign \new_[43797]_  = A233 & ~A232;
  assign \new_[43798]_  = A203 & \new_[43797]_ ;
  assign \new_[43801]_  = ~A266 & A265;
  assign \new_[43804]_  = A268 & A267;
  assign \new_[43805]_  = \new_[43804]_  & \new_[43801]_ ;
  assign \new_[43806]_  = \new_[43805]_  & \new_[43798]_ ;
  assign \new_[43810]_  = ~A166 & ~A167;
  assign \new_[43811]_  = A170 & \new_[43810]_ ;
  assign \new_[43815]_  = A201 & ~A200;
  assign \new_[43816]_  = A199 & \new_[43815]_ ;
  assign \new_[43817]_  = \new_[43816]_  & \new_[43811]_ ;
  assign \new_[43821]_  = A233 & ~A232;
  assign \new_[43822]_  = A203 & \new_[43821]_ ;
  assign \new_[43825]_  = ~A266 & A265;
  assign \new_[43828]_  = A269 & A267;
  assign \new_[43829]_  = \new_[43828]_  & \new_[43825]_ ;
  assign \new_[43830]_  = \new_[43829]_  & \new_[43822]_ ;
  assign \new_[43834]_  = ~A166 & ~A167;
  assign \new_[43835]_  = A170 & \new_[43834]_ ;
  assign \new_[43839]_  = A201 & ~A200;
  assign \new_[43840]_  = A199 & \new_[43839]_ ;
  assign \new_[43841]_  = \new_[43840]_  & \new_[43835]_ ;
  assign \new_[43845]_  = ~A234 & ~A233;
  assign \new_[43846]_  = A203 & \new_[43845]_ ;
  assign \new_[43849]_  = A266 & A265;
  assign \new_[43852]_  = ~A300 & A298;
  assign \new_[43853]_  = \new_[43852]_  & \new_[43849]_ ;
  assign \new_[43854]_  = \new_[43853]_  & \new_[43846]_ ;
  assign \new_[43858]_  = ~A166 & ~A167;
  assign \new_[43859]_  = A170 & \new_[43858]_ ;
  assign \new_[43863]_  = A201 & ~A200;
  assign \new_[43864]_  = A199 & \new_[43863]_ ;
  assign \new_[43865]_  = \new_[43864]_  & \new_[43859]_ ;
  assign \new_[43869]_  = ~A234 & ~A233;
  assign \new_[43870]_  = A203 & \new_[43869]_ ;
  assign \new_[43873]_  = A266 & A265;
  assign \new_[43876]_  = A299 & A298;
  assign \new_[43877]_  = \new_[43876]_  & \new_[43873]_ ;
  assign \new_[43878]_  = \new_[43877]_  & \new_[43870]_ ;
  assign \new_[43882]_  = ~A166 & ~A167;
  assign \new_[43883]_  = A170 & \new_[43882]_ ;
  assign \new_[43887]_  = A201 & ~A200;
  assign \new_[43888]_  = A199 & \new_[43887]_ ;
  assign \new_[43889]_  = \new_[43888]_  & \new_[43883]_ ;
  assign \new_[43893]_  = ~A234 & ~A233;
  assign \new_[43894]_  = A203 & \new_[43893]_ ;
  assign \new_[43897]_  = A266 & A265;
  assign \new_[43900]_  = ~A299 & ~A298;
  assign \new_[43901]_  = \new_[43900]_  & \new_[43897]_ ;
  assign \new_[43902]_  = \new_[43901]_  & \new_[43894]_ ;
  assign \new_[43906]_  = ~A166 & ~A167;
  assign \new_[43907]_  = A170 & \new_[43906]_ ;
  assign \new_[43911]_  = A201 & ~A200;
  assign \new_[43912]_  = A199 & \new_[43911]_ ;
  assign \new_[43913]_  = \new_[43912]_  & \new_[43907]_ ;
  assign \new_[43917]_  = ~A234 & ~A233;
  assign \new_[43918]_  = A203 & \new_[43917]_ ;
  assign \new_[43921]_  = ~A267 & ~A266;
  assign \new_[43924]_  = ~A300 & A298;
  assign \new_[43925]_  = \new_[43924]_  & \new_[43921]_ ;
  assign \new_[43926]_  = \new_[43925]_  & \new_[43918]_ ;
  assign \new_[43930]_  = ~A166 & ~A167;
  assign \new_[43931]_  = A170 & \new_[43930]_ ;
  assign \new_[43935]_  = A201 & ~A200;
  assign \new_[43936]_  = A199 & \new_[43935]_ ;
  assign \new_[43937]_  = \new_[43936]_  & \new_[43931]_ ;
  assign \new_[43941]_  = ~A234 & ~A233;
  assign \new_[43942]_  = A203 & \new_[43941]_ ;
  assign \new_[43945]_  = ~A267 & ~A266;
  assign \new_[43948]_  = A299 & A298;
  assign \new_[43949]_  = \new_[43948]_  & \new_[43945]_ ;
  assign \new_[43950]_  = \new_[43949]_  & \new_[43942]_ ;
  assign \new_[43954]_  = ~A166 & ~A167;
  assign \new_[43955]_  = A170 & \new_[43954]_ ;
  assign \new_[43959]_  = A201 & ~A200;
  assign \new_[43960]_  = A199 & \new_[43959]_ ;
  assign \new_[43961]_  = \new_[43960]_  & \new_[43955]_ ;
  assign \new_[43965]_  = ~A234 & ~A233;
  assign \new_[43966]_  = A203 & \new_[43965]_ ;
  assign \new_[43969]_  = ~A267 & ~A266;
  assign \new_[43972]_  = ~A299 & ~A298;
  assign \new_[43973]_  = \new_[43972]_  & \new_[43969]_ ;
  assign \new_[43974]_  = \new_[43973]_  & \new_[43966]_ ;
  assign \new_[43978]_  = ~A166 & ~A167;
  assign \new_[43979]_  = A170 & \new_[43978]_ ;
  assign \new_[43983]_  = A201 & ~A200;
  assign \new_[43984]_  = A199 & \new_[43983]_ ;
  assign \new_[43985]_  = \new_[43984]_  & \new_[43979]_ ;
  assign \new_[43989]_  = ~A234 & ~A233;
  assign \new_[43990]_  = A203 & \new_[43989]_ ;
  assign \new_[43993]_  = ~A266 & ~A265;
  assign \new_[43996]_  = ~A300 & A298;
  assign \new_[43997]_  = \new_[43996]_  & \new_[43993]_ ;
  assign \new_[43998]_  = \new_[43997]_  & \new_[43990]_ ;
  assign \new_[44002]_  = ~A166 & ~A167;
  assign \new_[44003]_  = A170 & \new_[44002]_ ;
  assign \new_[44007]_  = A201 & ~A200;
  assign \new_[44008]_  = A199 & \new_[44007]_ ;
  assign \new_[44009]_  = \new_[44008]_  & \new_[44003]_ ;
  assign \new_[44013]_  = ~A234 & ~A233;
  assign \new_[44014]_  = A203 & \new_[44013]_ ;
  assign \new_[44017]_  = ~A266 & ~A265;
  assign \new_[44020]_  = A299 & A298;
  assign \new_[44021]_  = \new_[44020]_  & \new_[44017]_ ;
  assign \new_[44022]_  = \new_[44021]_  & \new_[44014]_ ;
  assign \new_[44026]_  = ~A166 & ~A167;
  assign \new_[44027]_  = A170 & \new_[44026]_ ;
  assign \new_[44031]_  = A201 & ~A200;
  assign \new_[44032]_  = A199 & \new_[44031]_ ;
  assign \new_[44033]_  = \new_[44032]_  & \new_[44027]_ ;
  assign \new_[44037]_  = ~A234 & ~A233;
  assign \new_[44038]_  = A203 & \new_[44037]_ ;
  assign \new_[44041]_  = ~A266 & ~A265;
  assign \new_[44044]_  = ~A299 & ~A298;
  assign \new_[44045]_  = \new_[44044]_  & \new_[44041]_ ;
  assign \new_[44046]_  = \new_[44045]_  & \new_[44038]_ ;
  assign \new_[44050]_  = ~A166 & ~A167;
  assign \new_[44051]_  = A170 & \new_[44050]_ ;
  assign \new_[44055]_  = A201 & ~A200;
  assign \new_[44056]_  = A199 & \new_[44055]_ ;
  assign \new_[44057]_  = \new_[44056]_  & \new_[44051]_ ;
  assign \new_[44061]_  = ~A233 & A232;
  assign \new_[44062]_  = A203 & \new_[44061]_ ;
  assign \new_[44065]_  = A235 & A234;
  assign \new_[44068]_  = A299 & ~A298;
  assign \new_[44069]_  = \new_[44068]_  & \new_[44065]_ ;
  assign \new_[44070]_  = \new_[44069]_  & \new_[44062]_ ;
  assign \new_[44074]_  = ~A166 & ~A167;
  assign \new_[44075]_  = A170 & \new_[44074]_ ;
  assign \new_[44079]_  = A201 & ~A200;
  assign \new_[44080]_  = A199 & \new_[44079]_ ;
  assign \new_[44081]_  = \new_[44080]_  & \new_[44075]_ ;
  assign \new_[44085]_  = ~A233 & A232;
  assign \new_[44086]_  = A203 & \new_[44085]_ ;
  assign \new_[44089]_  = A235 & A234;
  assign \new_[44092]_  = A266 & ~A265;
  assign \new_[44093]_  = \new_[44092]_  & \new_[44089]_ ;
  assign \new_[44094]_  = \new_[44093]_  & \new_[44086]_ ;
  assign \new_[44098]_  = ~A166 & ~A167;
  assign \new_[44099]_  = A170 & \new_[44098]_ ;
  assign \new_[44103]_  = A201 & ~A200;
  assign \new_[44104]_  = A199 & \new_[44103]_ ;
  assign \new_[44105]_  = \new_[44104]_  & \new_[44099]_ ;
  assign \new_[44109]_  = ~A233 & A232;
  assign \new_[44110]_  = A203 & \new_[44109]_ ;
  assign \new_[44113]_  = A236 & A234;
  assign \new_[44116]_  = A299 & ~A298;
  assign \new_[44117]_  = \new_[44116]_  & \new_[44113]_ ;
  assign \new_[44118]_  = \new_[44117]_  & \new_[44110]_ ;
  assign \new_[44122]_  = ~A166 & ~A167;
  assign \new_[44123]_  = A170 & \new_[44122]_ ;
  assign \new_[44127]_  = A201 & ~A200;
  assign \new_[44128]_  = A199 & \new_[44127]_ ;
  assign \new_[44129]_  = \new_[44128]_  & \new_[44123]_ ;
  assign \new_[44133]_  = ~A233 & A232;
  assign \new_[44134]_  = A203 & \new_[44133]_ ;
  assign \new_[44137]_  = A236 & A234;
  assign \new_[44140]_  = A266 & ~A265;
  assign \new_[44141]_  = \new_[44140]_  & \new_[44137]_ ;
  assign \new_[44142]_  = \new_[44141]_  & \new_[44134]_ ;
  assign \new_[44146]_  = ~A166 & ~A167;
  assign \new_[44147]_  = A170 & \new_[44146]_ ;
  assign \new_[44151]_  = A201 & ~A200;
  assign \new_[44152]_  = A199 & \new_[44151]_ ;
  assign \new_[44153]_  = \new_[44152]_  & \new_[44147]_ ;
  assign \new_[44157]_  = ~A233 & ~A232;
  assign \new_[44158]_  = A203 & \new_[44157]_ ;
  assign \new_[44161]_  = A266 & A265;
  assign \new_[44164]_  = ~A300 & A298;
  assign \new_[44165]_  = \new_[44164]_  & \new_[44161]_ ;
  assign \new_[44166]_  = \new_[44165]_  & \new_[44158]_ ;
  assign \new_[44170]_  = ~A166 & ~A167;
  assign \new_[44171]_  = A170 & \new_[44170]_ ;
  assign \new_[44175]_  = A201 & ~A200;
  assign \new_[44176]_  = A199 & \new_[44175]_ ;
  assign \new_[44177]_  = \new_[44176]_  & \new_[44171]_ ;
  assign \new_[44181]_  = ~A233 & ~A232;
  assign \new_[44182]_  = A203 & \new_[44181]_ ;
  assign \new_[44185]_  = A266 & A265;
  assign \new_[44188]_  = A299 & A298;
  assign \new_[44189]_  = \new_[44188]_  & \new_[44185]_ ;
  assign \new_[44190]_  = \new_[44189]_  & \new_[44182]_ ;
  assign \new_[44194]_  = ~A166 & ~A167;
  assign \new_[44195]_  = A170 & \new_[44194]_ ;
  assign \new_[44199]_  = A201 & ~A200;
  assign \new_[44200]_  = A199 & \new_[44199]_ ;
  assign \new_[44201]_  = \new_[44200]_  & \new_[44195]_ ;
  assign \new_[44205]_  = ~A233 & ~A232;
  assign \new_[44206]_  = A203 & \new_[44205]_ ;
  assign \new_[44209]_  = A266 & A265;
  assign \new_[44212]_  = ~A299 & ~A298;
  assign \new_[44213]_  = \new_[44212]_  & \new_[44209]_ ;
  assign \new_[44214]_  = \new_[44213]_  & \new_[44206]_ ;
  assign \new_[44218]_  = ~A166 & ~A167;
  assign \new_[44219]_  = A170 & \new_[44218]_ ;
  assign \new_[44223]_  = A201 & ~A200;
  assign \new_[44224]_  = A199 & \new_[44223]_ ;
  assign \new_[44225]_  = \new_[44224]_  & \new_[44219]_ ;
  assign \new_[44229]_  = ~A233 & ~A232;
  assign \new_[44230]_  = A203 & \new_[44229]_ ;
  assign \new_[44233]_  = ~A267 & ~A266;
  assign \new_[44236]_  = ~A300 & A298;
  assign \new_[44237]_  = \new_[44236]_  & \new_[44233]_ ;
  assign \new_[44238]_  = \new_[44237]_  & \new_[44230]_ ;
  assign \new_[44242]_  = ~A166 & ~A167;
  assign \new_[44243]_  = A170 & \new_[44242]_ ;
  assign \new_[44247]_  = A201 & ~A200;
  assign \new_[44248]_  = A199 & \new_[44247]_ ;
  assign \new_[44249]_  = \new_[44248]_  & \new_[44243]_ ;
  assign \new_[44253]_  = ~A233 & ~A232;
  assign \new_[44254]_  = A203 & \new_[44253]_ ;
  assign \new_[44257]_  = ~A267 & ~A266;
  assign \new_[44260]_  = A299 & A298;
  assign \new_[44261]_  = \new_[44260]_  & \new_[44257]_ ;
  assign \new_[44262]_  = \new_[44261]_  & \new_[44254]_ ;
  assign \new_[44266]_  = ~A166 & ~A167;
  assign \new_[44267]_  = A170 & \new_[44266]_ ;
  assign \new_[44271]_  = A201 & ~A200;
  assign \new_[44272]_  = A199 & \new_[44271]_ ;
  assign \new_[44273]_  = \new_[44272]_  & \new_[44267]_ ;
  assign \new_[44277]_  = ~A233 & ~A232;
  assign \new_[44278]_  = A203 & \new_[44277]_ ;
  assign \new_[44281]_  = ~A267 & ~A266;
  assign \new_[44284]_  = ~A299 & ~A298;
  assign \new_[44285]_  = \new_[44284]_  & \new_[44281]_ ;
  assign \new_[44286]_  = \new_[44285]_  & \new_[44278]_ ;
  assign \new_[44290]_  = ~A166 & ~A167;
  assign \new_[44291]_  = A170 & \new_[44290]_ ;
  assign \new_[44295]_  = A201 & ~A200;
  assign \new_[44296]_  = A199 & \new_[44295]_ ;
  assign \new_[44297]_  = \new_[44296]_  & \new_[44291]_ ;
  assign \new_[44301]_  = ~A233 & ~A232;
  assign \new_[44302]_  = A203 & \new_[44301]_ ;
  assign \new_[44305]_  = ~A266 & ~A265;
  assign \new_[44308]_  = ~A300 & A298;
  assign \new_[44309]_  = \new_[44308]_  & \new_[44305]_ ;
  assign \new_[44310]_  = \new_[44309]_  & \new_[44302]_ ;
  assign \new_[44314]_  = ~A166 & ~A167;
  assign \new_[44315]_  = A170 & \new_[44314]_ ;
  assign \new_[44319]_  = A201 & ~A200;
  assign \new_[44320]_  = A199 & \new_[44319]_ ;
  assign \new_[44321]_  = \new_[44320]_  & \new_[44315]_ ;
  assign \new_[44325]_  = ~A233 & ~A232;
  assign \new_[44326]_  = A203 & \new_[44325]_ ;
  assign \new_[44329]_  = ~A266 & ~A265;
  assign \new_[44332]_  = A299 & A298;
  assign \new_[44333]_  = \new_[44332]_  & \new_[44329]_ ;
  assign \new_[44334]_  = \new_[44333]_  & \new_[44326]_ ;
  assign \new_[44338]_  = ~A166 & ~A167;
  assign \new_[44339]_  = A170 & \new_[44338]_ ;
  assign \new_[44343]_  = A201 & ~A200;
  assign \new_[44344]_  = A199 & \new_[44343]_ ;
  assign \new_[44345]_  = \new_[44344]_  & \new_[44339]_ ;
  assign \new_[44349]_  = ~A233 & ~A232;
  assign \new_[44350]_  = A203 & \new_[44349]_ ;
  assign \new_[44353]_  = ~A266 & ~A265;
  assign \new_[44356]_  = ~A299 & ~A298;
  assign \new_[44357]_  = \new_[44356]_  & \new_[44353]_ ;
  assign \new_[44358]_  = \new_[44357]_  & \new_[44350]_ ;
  assign \new_[44362]_  = A167 & ~A168;
  assign \new_[44363]_  = A170 & \new_[44362]_ ;
  assign \new_[44367]_  = A200 & ~A199;
  assign \new_[44368]_  = A166 & \new_[44367]_ ;
  assign \new_[44369]_  = \new_[44368]_  & \new_[44363]_ ;
  assign \new_[44373]_  = A265 & A233;
  assign \new_[44374]_  = A232 & \new_[44373]_ ;
  assign \new_[44377]_  = ~A269 & ~A268;
  assign \new_[44380]_  = ~A300 & ~A299;
  assign \new_[44381]_  = \new_[44380]_  & \new_[44377]_ ;
  assign \new_[44382]_  = \new_[44381]_  & \new_[44374]_ ;
  assign \new_[44386]_  = A167 & ~A168;
  assign \new_[44387]_  = A170 & \new_[44386]_ ;
  assign \new_[44391]_  = A200 & ~A199;
  assign \new_[44392]_  = A166 & \new_[44391]_ ;
  assign \new_[44393]_  = \new_[44392]_  & \new_[44387]_ ;
  assign \new_[44397]_  = A265 & A233;
  assign \new_[44398]_  = A232 & \new_[44397]_ ;
  assign \new_[44401]_  = ~A269 & ~A268;
  assign \new_[44404]_  = A299 & A298;
  assign \new_[44405]_  = \new_[44404]_  & \new_[44401]_ ;
  assign \new_[44406]_  = \new_[44405]_  & \new_[44398]_ ;
  assign \new_[44410]_  = A167 & ~A168;
  assign \new_[44411]_  = A170 & \new_[44410]_ ;
  assign \new_[44415]_  = A200 & ~A199;
  assign \new_[44416]_  = A166 & \new_[44415]_ ;
  assign \new_[44417]_  = \new_[44416]_  & \new_[44411]_ ;
  assign \new_[44421]_  = A265 & A233;
  assign \new_[44422]_  = A232 & \new_[44421]_ ;
  assign \new_[44425]_  = ~A269 & ~A268;
  assign \new_[44428]_  = ~A299 & ~A298;
  assign \new_[44429]_  = \new_[44428]_  & \new_[44425]_ ;
  assign \new_[44430]_  = \new_[44429]_  & \new_[44422]_ ;
  assign \new_[44434]_  = A167 & ~A168;
  assign \new_[44435]_  = A170 & \new_[44434]_ ;
  assign \new_[44439]_  = A200 & ~A199;
  assign \new_[44440]_  = A166 & \new_[44439]_ ;
  assign \new_[44441]_  = \new_[44440]_  & \new_[44435]_ ;
  assign \new_[44445]_  = A265 & A233;
  assign \new_[44446]_  = A232 & \new_[44445]_ ;
  assign \new_[44449]_  = ~A299 & ~A267;
  assign \new_[44452]_  = ~A302 & ~A301;
  assign \new_[44453]_  = \new_[44452]_  & \new_[44449]_ ;
  assign \new_[44454]_  = \new_[44453]_  & \new_[44446]_ ;
  assign \new_[44458]_  = A167 & ~A168;
  assign \new_[44459]_  = A170 & \new_[44458]_ ;
  assign \new_[44463]_  = A200 & ~A199;
  assign \new_[44464]_  = A166 & \new_[44463]_ ;
  assign \new_[44465]_  = \new_[44464]_  & \new_[44459]_ ;
  assign \new_[44469]_  = A265 & A233;
  assign \new_[44470]_  = A232 & \new_[44469]_ ;
  assign \new_[44473]_  = ~A299 & A266;
  assign \new_[44476]_  = ~A302 & ~A301;
  assign \new_[44477]_  = \new_[44476]_  & \new_[44473]_ ;
  assign \new_[44478]_  = \new_[44477]_  & \new_[44470]_ ;
  assign \new_[44482]_  = A167 & ~A168;
  assign \new_[44483]_  = A170 & \new_[44482]_ ;
  assign \new_[44487]_  = A200 & ~A199;
  assign \new_[44488]_  = A166 & \new_[44487]_ ;
  assign \new_[44489]_  = \new_[44488]_  & \new_[44483]_ ;
  assign \new_[44493]_  = ~A265 & A233;
  assign \new_[44494]_  = A232 & \new_[44493]_ ;
  assign \new_[44497]_  = ~A299 & ~A266;
  assign \new_[44500]_  = ~A302 & ~A301;
  assign \new_[44501]_  = \new_[44500]_  & \new_[44497]_ ;
  assign \new_[44502]_  = \new_[44501]_  & \new_[44494]_ ;
  assign \new_[44506]_  = A167 & ~A168;
  assign \new_[44507]_  = A170 & \new_[44506]_ ;
  assign \new_[44511]_  = A200 & ~A199;
  assign \new_[44512]_  = A166 & \new_[44511]_ ;
  assign \new_[44513]_  = \new_[44512]_  & \new_[44507]_ ;
  assign \new_[44517]_  = ~A236 & ~A235;
  assign \new_[44518]_  = ~A233 & \new_[44517]_ ;
  assign \new_[44521]_  = A266 & A265;
  assign \new_[44524]_  = ~A300 & A298;
  assign \new_[44525]_  = \new_[44524]_  & \new_[44521]_ ;
  assign \new_[44526]_  = \new_[44525]_  & \new_[44518]_ ;
  assign \new_[44530]_  = A167 & ~A168;
  assign \new_[44531]_  = A170 & \new_[44530]_ ;
  assign \new_[44535]_  = A200 & ~A199;
  assign \new_[44536]_  = A166 & \new_[44535]_ ;
  assign \new_[44537]_  = \new_[44536]_  & \new_[44531]_ ;
  assign \new_[44541]_  = ~A236 & ~A235;
  assign \new_[44542]_  = ~A233 & \new_[44541]_ ;
  assign \new_[44545]_  = A266 & A265;
  assign \new_[44548]_  = A299 & A298;
  assign \new_[44549]_  = \new_[44548]_  & \new_[44545]_ ;
  assign \new_[44550]_  = \new_[44549]_  & \new_[44542]_ ;
  assign \new_[44554]_  = A167 & ~A168;
  assign \new_[44555]_  = A170 & \new_[44554]_ ;
  assign \new_[44559]_  = A200 & ~A199;
  assign \new_[44560]_  = A166 & \new_[44559]_ ;
  assign \new_[44561]_  = \new_[44560]_  & \new_[44555]_ ;
  assign \new_[44565]_  = ~A236 & ~A235;
  assign \new_[44566]_  = ~A233 & \new_[44565]_ ;
  assign \new_[44569]_  = A266 & A265;
  assign \new_[44572]_  = ~A299 & ~A298;
  assign \new_[44573]_  = \new_[44572]_  & \new_[44569]_ ;
  assign \new_[44574]_  = \new_[44573]_  & \new_[44566]_ ;
  assign \new_[44578]_  = A167 & ~A168;
  assign \new_[44579]_  = A170 & \new_[44578]_ ;
  assign \new_[44583]_  = A200 & ~A199;
  assign \new_[44584]_  = A166 & \new_[44583]_ ;
  assign \new_[44585]_  = \new_[44584]_  & \new_[44579]_ ;
  assign \new_[44589]_  = ~A236 & ~A235;
  assign \new_[44590]_  = ~A233 & \new_[44589]_ ;
  assign \new_[44593]_  = ~A267 & ~A266;
  assign \new_[44596]_  = ~A300 & A298;
  assign \new_[44597]_  = \new_[44596]_  & \new_[44593]_ ;
  assign \new_[44598]_  = \new_[44597]_  & \new_[44590]_ ;
  assign \new_[44602]_  = A167 & ~A168;
  assign \new_[44603]_  = A170 & \new_[44602]_ ;
  assign \new_[44607]_  = A200 & ~A199;
  assign \new_[44608]_  = A166 & \new_[44607]_ ;
  assign \new_[44609]_  = \new_[44608]_  & \new_[44603]_ ;
  assign \new_[44613]_  = ~A236 & ~A235;
  assign \new_[44614]_  = ~A233 & \new_[44613]_ ;
  assign \new_[44617]_  = ~A267 & ~A266;
  assign \new_[44620]_  = A299 & A298;
  assign \new_[44621]_  = \new_[44620]_  & \new_[44617]_ ;
  assign \new_[44622]_  = \new_[44621]_  & \new_[44614]_ ;
  assign \new_[44626]_  = A167 & ~A168;
  assign \new_[44627]_  = A170 & \new_[44626]_ ;
  assign \new_[44631]_  = A200 & ~A199;
  assign \new_[44632]_  = A166 & \new_[44631]_ ;
  assign \new_[44633]_  = \new_[44632]_  & \new_[44627]_ ;
  assign \new_[44637]_  = ~A236 & ~A235;
  assign \new_[44638]_  = ~A233 & \new_[44637]_ ;
  assign \new_[44641]_  = ~A267 & ~A266;
  assign \new_[44644]_  = ~A299 & ~A298;
  assign \new_[44645]_  = \new_[44644]_  & \new_[44641]_ ;
  assign \new_[44646]_  = \new_[44645]_  & \new_[44638]_ ;
  assign \new_[44650]_  = A167 & ~A168;
  assign \new_[44651]_  = A170 & \new_[44650]_ ;
  assign \new_[44655]_  = A200 & ~A199;
  assign \new_[44656]_  = A166 & \new_[44655]_ ;
  assign \new_[44657]_  = \new_[44656]_  & \new_[44651]_ ;
  assign \new_[44661]_  = ~A236 & ~A235;
  assign \new_[44662]_  = ~A233 & \new_[44661]_ ;
  assign \new_[44665]_  = ~A266 & ~A265;
  assign \new_[44668]_  = ~A300 & A298;
  assign \new_[44669]_  = \new_[44668]_  & \new_[44665]_ ;
  assign \new_[44670]_  = \new_[44669]_  & \new_[44662]_ ;
  assign \new_[44674]_  = A167 & ~A168;
  assign \new_[44675]_  = A170 & \new_[44674]_ ;
  assign \new_[44679]_  = A200 & ~A199;
  assign \new_[44680]_  = A166 & \new_[44679]_ ;
  assign \new_[44681]_  = \new_[44680]_  & \new_[44675]_ ;
  assign \new_[44685]_  = ~A236 & ~A235;
  assign \new_[44686]_  = ~A233 & \new_[44685]_ ;
  assign \new_[44689]_  = ~A266 & ~A265;
  assign \new_[44692]_  = A299 & A298;
  assign \new_[44693]_  = \new_[44692]_  & \new_[44689]_ ;
  assign \new_[44694]_  = \new_[44693]_  & \new_[44686]_ ;
  assign \new_[44698]_  = A167 & ~A168;
  assign \new_[44699]_  = A170 & \new_[44698]_ ;
  assign \new_[44703]_  = A200 & ~A199;
  assign \new_[44704]_  = A166 & \new_[44703]_ ;
  assign \new_[44705]_  = \new_[44704]_  & \new_[44699]_ ;
  assign \new_[44709]_  = ~A236 & ~A235;
  assign \new_[44710]_  = ~A233 & \new_[44709]_ ;
  assign \new_[44713]_  = ~A266 & ~A265;
  assign \new_[44716]_  = ~A299 & ~A298;
  assign \new_[44717]_  = \new_[44716]_  & \new_[44713]_ ;
  assign \new_[44718]_  = \new_[44717]_  & \new_[44710]_ ;
  assign \new_[44722]_  = A167 & ~A168;
  assign \new_[44723]_  = A170 & \new_[44722]_ ;
  assign \new_[44727]_  = A200 & ~A199;
  assign \new_[44728]_  = A166 & \new_[44727]_ ;
  assign \new_[44729]_  = \new_[44728]_  & \new_[44723]_ ;
  assign \new_[44733]_  = A265 & ~A234;
  assign \new_[44734]_  = ~A233 & \new_[44733]_ ;
  assign \new_[44737]_  = A298 & A266;
  assign \new_[44740]_  = ~A302 & ~A301;
  assign \new_[44741]_  = \new_[44740]_  & \new_[44737]_ ;
  assign \new_[44742]_  = \new_[44741]_  & \new_[44734]_ ;
  assign \new_[44746]_  = A167 & ~A168;
  assign \new_[44747]_  = A170 & \new_[44746]_ ;
  assign \new_[44751]_  = A200 & ~A199;
  assign \new_[44752]_  = A166 & \new_[44751]_ ;
  assign \new_[44753]_  = \new_[44752]_  & \new_[44747]_ ;
  assign \new_[44757]_  = ~A266 & ~A234;
  assign \new_[44758]_  = ~A233 & \new_[44757]_ ;
  assign \new_[44761]_  = ~A269 & ~A268;
  assign \new_[44764]_  = ~A300 & A298;
  assign \new_[44765]_  = \new_[44764]_  & \new_[44761]_ ;
  assign \new_[44766]_  = \new_[44765]_  & \new_[44758]_ ;
  assign \new_[44770]_  = A167 & ~A168;
  assign \new_[44771]_  = A170 & \new_[44770]_ ;
  assign \new_[44775]_  = A200 & ~A199;
  assign \new_[44776]_  = A166 & \new_[44775]_ ;
  assign \new_[44777]_  = \new_[44776]_  & \new_[44771]_ ;
  assign \new_[44781]_  = ~A266 & ~A234;
  assign \new_[44782]_  = ~A233 & \new_[44781]_ ;
  assign \new_[44785]_  = ~A269 & ~A268;
  assign \new_[44788]_  = A299 & A298;
  assign \new_[44789]_  = \new_[44788]_  & \new_[44785]_ ;
  assign \new_[44790]_  = \new_[44789]_  & \new_[44782]_ ;
  assign \new_[44794]_  = A167 & ~A168;
  assign \new_[44795]_  = A170 & \new_[44794]_ ;
  assign \new_[44799]_  = A200 & ~A199;
  assign \new_[44800]_  = A166 & \new_[44799]_ ;
  assign \new_[44801]_  = \new_[44800]_  & \new_[44795]_ ;
  assign \new_[44805]_  = ~A266 & ~A234;
  assign \new_[44806]_  = ~A233 & \new_[44805]_ ;
  assign \new_[44809]_  = ~A269 & ~A268;
  assign \new_[44812]_  = ~A299 & ~A298;
  assign \new_[44813]_  = \new_[44812]_  & \new_[44809]_ ;
  assign \new_[44814]_  = \new_[44813]_  & \new_[44806]_ ;
  assign \new_[44818]_  = A167 & ~A168;
  assign \new_[44819]_  = A170 & \new_[44818]_ ;
  assign \new_[44823]_  = A200 & ~A199;
  assign \new_[44824]_  = A166 & \new_[44823]_ ;
  assign \new_[44825]_  = \new_[44824]_  & \new_[44819]_ ;
  assign \new_[44829]_  = ~A266 & ~A234;
  assign \new_[44830]_  = ~A233 & \new_[44829]_ ;
  assign \new_[44833]_  = A298 & ~A267;
  assign \new_[44836]_  = ~A302 & ~A301;
  assign \new_[44837]_  = \new_[44836]_  & \new_[44833]_ ;
  assign \new_[44838]_  = \new_[44837]_  & \new_[44830]_ ;
  assign \new_[44842]_  = A167 & ~A168;
  assign \new_[44843]_  = A170 & \new_[44842]_ ;
  assign \new_[44847]_  = A200 & ~A199;
  assign \new_[44848]_  = A166 & \new_[44847]_ ;
  assign \new_[44849]_  = \new_[44848]_  & \new_[44843]_ ;
  assign \new_[44853]_  = ~A265 & ~A234;
  assign \new_[44854]_  = ~A233 & \new_[44853]_ ;
  assign \new_[44857]_  = A298 & ~A266;
  assign \new_[44860]_  = ~A302 & ~A301;
  assign \new_[44861]_  = \new_[44860]_  & \new_[44857]_ ;
  assign \new_[44862]_  = \new_[44861]_  & \new_[44854]_ ;
  assign \new_[44866]_  = A167 & ~A168;
  assign \new_[44867]_  = A170 & \new_[44866]_ ;
  assign \new_[44871]_  = A200 & ~A199;
  assign \new_[44872]_  = A166 & \new_[44871]_ ;
  assign \new_[44873]_  = \new_[44872]_  & \new_[44867]_ ;
  assign \new_[44877]_  = A265 & ~A233;
  assign \new_[44878]_  = ~A232 & \new_[44877]_ ;
  assign \new_[44881]_  = A298 & A266;
  assign \new_[44884]_  = ~A302 & ~A301;
  assign \new_[44885]_  = \new_[44884]_  & \new_[44881]_ ;
  assign \new_[44886]_  = \new_[44885]_  & \new_[44878]_ ;
  assign \new_[44890]_  = A167 & ~A168;
  assign \new_[44891]_  = A170 & \new_[44890]_ ;
  assign \new_[44895]_  = A200 & ~A199;
  assign \new_[44896]_  = A166 & \new_[44895]_ ;
  assign \new_[44897]_  = \new_[44896]_  & \new_[44891]_ ;
  assign \new_[44901]_  = ~A266 & ~A233;
  assign \new_[44902]_  = ~A232 & \new_[44901]_ ;
  assign \new_[44905]_  = ~A269 & ~A268;
  assign \new_[44908]_  = ~A300 & A298;
  assign \new_[44909]_  = \new_[44908]_  & \new_[44905]_ ;
  assign \new_[44910]_  = \new_[44909]_  & \new_[44902]_ ;
  assign \new_[44914]_  = A167 & ~A168;
  assign \new_[44915]_  = A170 & \new_[44914]_ ;
  assign \new_[44919]_  = A200 & ~A199;
  assign \new_[44920]_  = A166 & \new_[44919]_ ;
  assign \new_[44921]_  = \new_[44920]_  & \new_[44915]_ ;
  assign \new_[44925]_  = ~A266 & ~A233;
  assign \new_[44926]_  = ~A232 & \new_[44925]_ ;
  assign \new_[44929]_  = ~A269 & ~A268;
  assign \new_[44932]_  = A299 & A298;
  assign \new_[44933]_  = \new_[44932]_  & \new_[44929]_ ;
  assign \new_[44934]_  = \new_[44933]_  & \new_[44926]_ ;
  assign \new_[44938]_  = A167 & ~A168;
  assign \new_[44939]_  = A170 & \new_[44938]_ ;
  assign \new_[44943]_  = A200 & ~A199;
  assign \new_[44944]_  = A166 & \new_[44943]_ ;
  assign \new_[44945]_  = \new_[44944]_  & \new_[44939]_ ;
  assign \new_[44949]_  = ~A266 & ~A233;
  assign \new_[44950]_  = ~A232 & \new_[44949]_ ;
  assign \new_[44953]_  = ~A269 & ~A268;
  assign \new_[44956]_  = ~A299 & ~A298;
  assign \new_[44957]_  = \new_[44956]_  & \new_[44953]_ ;
  assign \new_[44958]_  = \new_[44957]_  & \new_[44950]_ ;
  assign \new_[44962]_  = A167 & ~A168;
  assign \new_[44963]_  = A170 & \new_[44962]_ ;
  assign \new_[44967]_  = A200 & ~A199;
  assign \new_[44968]_  = A166 & \new_[44967]_ ;
  assign \new_[44969]_  = \new_[44968]_  & \new_[44963]_ ;
  assign \new_[44973]_  = ~A266 & ~A233;
  assign \new_[44974]_  = ~A232 & \new_[44973]_ ;
  assign \new_[44977]_  = A298 & ~A267;
  assign \new_[44980]_  = ~A302 & ~A301;
  assign \new_[44981]_  = \new_[44980]_  & \new_[44977]_ ;
  assign \new_[44982]_  = \new_[44981]_  & \new_[44974]_ ;
  assign \new_[44986]_  = A167 & ~A168;
  assign \new_[44987]_  = A170 & \new_[44986]_ ;
  assign \new_[44991]_  = A200 & ~A199;
  assign \new_[44992]_  = A166 & \new_[44991]_ ;
  assign \new_[44993]_  = \new_[44992]_  & \new_[44987]_ ;
  assign \new_[44997]_  = ~A265 & ~A233;
  assign \new_[44998]_  = ~A232 & \new_[44997]_ ;
  assign \new_[45001]_  = A298 & ~A266;
  assign \new_[45004]_  = ~A302 & ~A301;
  assign \new_[45005]_  = \new_[45004]_  & \new_[45001]_ ;
  assign \new_[45006]_  = \new_[45005]_  & \new_[44998]_ ;
  assign \new_[45010]_  = A167 & ~A168;
  assign \new_[45011]_  = ~A170 & \new_[45010]_ ;
  assign \new_[45015]_  = A200 & ~A199;
  assign \new_[45016]_  = ~A166 & \new_[45015]_ ;
  assign \new_[45017]_  = \new_[45016]_  & \new_[45011]_ ;
  assign \new_[45021]_  = A265 & A233;
  assign \new_[45022]_  = A232 & \new_[45021]_ ;
  assign \new_[45025]_  = ~A269 & ~A268;
  assign \new_[45028]_  = ~A300 & ~A299;
  assign \new_[45029]_  = \new_[45028]_  & \new_[45025]_ ;
  assign \new_[45030]_  = \new_[45029]_  & \new_[45022]_ ;
  assign \new_[45034]_  = A167 & ~A168;
  assign \new_[45035]_  = ~A170 & \new_[45034]_ ;
  assign \new_[45039]_  = A200 & ~A199;
  assign \new_[45040]_  = ~A166 & \new_[45039]_ ;
  assign \new_[45041]_  = \new_[45040]_  & \new_[45035]_ ;
  assign \new_[45045]_  = A265 & A233;
  assign \new_[45046]_  = A232 & \new_[45045]_ ;
  assign \new_[45049]_  = ~A269 & ~A268;
  assign \new_[45052]_  = A299 & A298;
  assign \new_[45053]_  = \new_[45052]_  & \new_[45049]_ ;
  assign \new_[45054]_  = \new_[45053]_  & \new_[45046]_ ;
  assign \new_[45058]_  = A167 & ~A168;
  assign \new_[45059]_  = ~A170 & \new_[45058]_ ;
  assign \new_[45063]_  = A200 & ~A199;
  assign \new_[45064]_  = ~A166 & \new_[45063]_ ;
  assign \new_[45065]_  = \new_[45064]_  & \new_[45059]_ ;
  assign \new_[45069]_  = A265 & A233;
  assign \new_[45070]_  = A232 & \new_[45069]_ ;
  assign \new_[45073]_  = ~A269 & ~A268;
  assign \new_[45076]_  = ~A299 & ~A298;
  assign \new_[45077]_  = \new_[45076]_  & \new_[45073]_ ;
  assign \new_[45078]_  = \new_[45077]_  & \new_[45070]_ ;
  assign \new_[45082]_  = A167 & ~A168;
  assign \new_[45083]_  = ~A170 & \new_[45082]_ ;
  assign \new_[45087]_  = A200 & ~A199;
  assign \new_[45088]_  = ~A166 & \new_[45087]_ ;
  assign \new_[45089]_  = \new_[45088]_  & \new_[45083]_ ;
  assign \new_[45093]_  = A265 & A233;
  assign \new_[45094]_  = A232 & \new_[45093]_ ;
  assign \new_[45097]_  = ~A299 & ~A267;
  assign \new_[45100]_  = ~A302 & ~A301;
  assign \new_[45101]_  = \new_[45100]_  & \new_[45097]_ ;
  assign \new_[45102]_  = \new_[45101]_  & \new_[45094]_ ;
  assign \new_[45106]_  = A167 & ~A168;
  assign \new_[45107]_  = ~A170 & \new_[45106]_ ;
  assign \new_[45111]_  = A200 & ~A199;
  assign \new_[45112]_  = ~A166 & \new_[45111]_ ;
  assign \new_[45113]_  = \new_[45112]_  & \new_[45107]_ ;
  assign \new_[45117]_  = A265 & A233;
  assign \new_[45118]_  = A232 & \new_[45117]_ ;
  assign \new_[45121]_  = ~A299 & A266;
  assign \new_[45124]_  = ~A302 & ~A301;
  assign \new_[45125]_  = \new_[45124]_  & \new_[45121]_ ;
  assign \new_[45126]_  = \new_[45125]_  & \new_[45118]_ ;
  assign \new_[45130]_  = A167 & ~A168;
  assign \new_[45131]_  = ~A170 & \new_[45130]_ ;
  assign \new_[45135]_  = A200 & ~A199;
  assign \new_[45136]_  = ~A166 & \new_[45135]_ ;
  assign \new_[45137]_  = \new_[45136]_  & \new_[45131]_ ;
  assign \new_[45141]_  = ~A265 & A233;
  assign \new_[45142]_  = A232 & \new_[45141]_ ;
  assign \new_[45145]_  = ~A299 & ~A266;
  assign \new_[45148]_  = ~A302 & ~A301;
  assign \new_[45149]_  = \new_[45148]_  & \new_[45145]_ ;
  assign \new_[45150]_  = \new_[45149]_  & \new_[45142]_ ;
  assign \new_[45154]_  = A167 & ~A168;
  assign \new_[45155]_  = ~A170 & \new_[45154]_ ;
  assign \new_[45159]_  = A200 & ~A199;
  assign \new_[45160]_  = ~A166 & \new_[45159]_ ;
  assign \new_[45161]_  = \new_[45160]_  & \new_[45155]_ ;
  assign \new_[45165]_  = ~A236 & ~A235;
  assign \new_[45166]_  = ~A233 & \new_[45165]_ ;
  assign \new_[45169]_  = A266 & A265;
  assign \new_[45172]_  = ~A300 & A298;
  assign \new_[45173]_  = \new_[45172]_  & \new_[45169]_ ;
  assign \new_[45174]_  = \new_[45173]_  & \new_[45166]_ ;
  assign \new_[45178]_  = A167 & ~A168;
  assign \new_[45179]_  = ~A170 & \new_[45178]_ ;
  assign \new_[45183]_  = A200 & ~A199;
  assign \new_[45184]_  = ~A166 & \new_[45183]_ ;
  assign \new_[45185]_  = \new_[45184]_  & \new_[45179]_ ;
  assign \new_[45189]_  = ~A236 & ~A235;
  assign \new_[45190]_  = ~A233 & \new_[45189]_ ;
  assign \new_[45193]_  = A266 & A265;
  assign \new_[45196]_  = A299 & A298;
  assign \new_[45197]_  = \new_[45196]_  & \new_[45193]_ ;
  assign \new_[45198]_  = \new_[45197]_  & \new_[45190]_ ;
  assign \new_[45202]_  = A167 & ~A168;
  assign \new_[45203]_  = ~A170 & \new_[45202]_ ;
  assign \new_[45207]_  = A200 & ~A199;
  assign \new_[45208]_  = ~A166 & \new_[45207]_ ;
  assign \new_[45209]_  = \new_[45208]_  & \new_[45203]_ ;
  assign \new_[45213]_  = ~A236 & ~A235;
  assign \new_[45214]_  = ~A233 & \new_[45213]_ ;
  assign \new_[45217]_  = A266 & A265;
  assign \new_[45220]_  = ~A299 & ~A298;
  assign \new_[45221]_  = \new_[45220]_  & \new_[45217]_ ;
  assign \new_[45222]_  = \new_[45221]_  & \new_[45214]_ ;
  assign \new_[45226]_  = A167 & ~A168;
  assign \new_[45227]_  = ~A170 & \new_[45226]_ ;
  assign \new_[45231]_  = A200 & ~A199;
  assign \new_[45232]_  = ~A166 & \new_[45231]_ ;
  assign \new_[45233]_  = \new_[45232]_  & \new_[45227]_ ;
  assign \new_[45237]_  = ~A236 & ~A235;
  assign \new_[45238]_  = ~A233 & \new_[45237]_ ;
  assign \new_[45241]_  = ~A267 & ~A266;
  assign \new_[45244]_  = ~A300 & A298;
  assign \new_[45245]_  = \new_[45244]_  & \new_[45241]_ ;
  assign \new_[45246]_  = \new_[45245]_  & \new_[45238]_ ;
  assign \new_[45250]_  = A167 & ~A168;
  assign \new_[45251]_  = ~A170 & \new_[45250]_ ;
  assign \new_[45255]_  = A200 & ~A199;
  assign \new_[45256]_  = ~A166 & \new_[45255]_ ;
  assign \new_[45257]_  = \new_[45256]_  & \new_[45251]_ ;
  assign \new_[45261]_  = ~A236 & ~A235;
  assign \new_[45262]_  = ~A233 & \new_[45261]_ ;
  assign \new_[45265]_  = ~A267 & ~A266;
  assign \new_[45268]_  = A299 & A298;
  assign \new_[45269]_  = \new_[45268]_  & \new_[45265]_ ;
  assign \new_[45270]_  = \new_[45269]_  & \new_[45262]_ ;
  assign \new_[45274]_  = A167 & ~A168;
  assign \new_[45275]_  = ~A170 & \new_[45274]_ ;
  assign \new_[45279]_  = A200 & ~A199;
  assign \new_[45280]_  = ~A166 & \new_[45279]_ ;
  assign \new_[45281]_  = \new_[45280]_  & \new_[45275]_ ;
  assign \new_[45285]_  = ~A236 & ~A235;
  assign \new_[45286]_  = ~A233 & \new_[45285]_ ;
  assign \new_[45289]_  = ~A267 & ~A266;
  assign \new_[45292]_  = ~A299 & ~A298;
  assign \new_[45293]_  = \new_[45292]_  & \new_[45289]_ ;
  assign \new_[45294]_  = \new_[45293]_  & \new_[45286]_ ;
  assign \new_[45298]_  = A167 & ~A168;
  assign \new_[45299]_  = ~A170 & \new_[45298]_ ;
  assign \new_[45303]_  = A200 & ~A199;
  assign \new_[45304]_  = ~A166 & \new_[45303]_ ;
  assign \new_[45305]_  = \new_[45304]_  & \new_[45299]_ ;
  assign \new_[45309]_  = ~A236 & ~A235;
  assign \new_[45310]_  = ~A233 & \new_[45309]_ ;
  assign \new_[45313]_  = ~A266 & ~A265;
  assign \new_[45316]_  = ~A300 & A298;
  assign \new_[45317]_  = \new_[45316]_  & \new_[45313]_ ;
  assign \new_[45318]_  = \new_[45317]_  & \new_[45310]_ ;
  assign \new_[45322]_  = A167 & ~A168;
  assign \new_[45323]_  = ~A170 & \new_[45322]_ ;
  assign \new_[45327]_  = A200 & ~A199;
  assign \new_[45328]_  = ~A166 & \new_[45327]_ ;
  assign \new_[45329]_  = \new_[45328]_  & \new_[45323]_ ;
  assign \new_[45333]_  = ~A236 & ~A235;
  assign \new_[45334]_  = ~A233 & \new_[45333]_ ;
  assign \new_[45337]_  = ~A266 & ~A265;
  assign \new_[45340]_  = A299 & A298;
  assign \new_[45341]_  = \new_[45340]_  & \new_[45337]_ ;
  assign \new_[45342]_  = \new_[45341]_  & \new_[45334]_ ;
  assign \new_[45346]_  = A167 & ~A168;
  assign \new_[45347]_  = ~A170 & \new_[45346]_ ;
  assign \new_[45351]_  = A200 & ~A199;
  assign \new_[45352]_  = ~A166 & \new_[45351]_ ;
  assign \new_[45353]_  = \new_[45352]_  & \new_[45347]_ ;
  assign \new_[45357]_  = ~A236 & ~A235;
  assign \new_[45358]_  = ~A233 & \new_[45357]_ ;
  assign \new_[45361]_  = ~A266 & ~A265;
  assign \new_[45364]_  = ~A299 & ~A298;
  assign \new_[45365]_  = \new_[45364]_  & \new_[45361]_ ;
  assign \new_[45366]_  = \new_[45365]_  & \new_[45358]_ ;
  assign \new_[45370]_  = A167 & ~A168;
  assign \new_[45371]_  = ~A170 & \new_[45370]_ ;
  assign \new_[45375]_  = A200 & ~A199;
  assign \new_[45376]_  = ~A166 & \new_[45375]_ ;
  assign \new_[45377]_  = \new_[45376]_  & \new_[45371]_ ;
  assign \new_[45381]_  = A265 & ~A234;
  assign \new_[45382]_  = ~A233 & \new_[45381]_ ;
  assign \new_[45385]_  = A298 & A266;
  assign \new_[45388]_  = ~A302 & ~A301;
  assign \new_[45389]_  = \new_[45388]_  & \new_[45385]_ ;
  assign \new_[45390]_  = \new_[45389]_  & \new_[45382]_ ;
  assign \new_[45394]_  = A167 & ~A168;
  assign \new_[45395]_  = ~A170 & \new_[45394]_ ;
  assign \new_[45399]_  = A200 & ~A199;
  assign \new_[45400]_  = ~A166 & \new_[45399]_ ;
  assign \new_[45401]_  = \new_[45400]_  & \new_[45395]_ ;
  assign \new_[45405]_  = ~A266 & ~A234;
  assign \new_[45406]_  = ~A233 & \new_[45405]_ ;
  assign \new_[45409]_  = ~A269 & ~A268;
  assign \new_[45412]_  = ~A300 & A298;
  assign \new_[45413]_  = \new_[45412]_  & \new_[45409]_ ;
  assign \new_[45414]_  = \new_[45413]_  & \new_[45406]_ ;
  assign \new_[45418]_  = A167 & ~A168;
  assign \new_[45419]_  = ~A170 & \new_[45418]_ ;
  assign \new_[45423]_  = A200 & ~A199;
  assign \new_[45424]_  = ~A166 & \new_[45423]_ ;
  assign \new_[45425]_  = \new_[45424]_  & \new_[45419]_ ;
  assign \new_[45429]_  = ~A266 & ~A234;
  assign \new_[45430]_  = ~A233 & \new_[45429]_ ;
  assign \new_[45433]_  = ~A269 & ~A268;
  assign \new_[45436]_  = A299 & A298;
  assign \new_[45437]_  = \new_[45436]_  & \new_[45433]_ ;
  assign \new_[45438]_  = \new_[45437]_  & \new_[45430]_ ;
  assign \new_[45442]_  = A167 & ~A168;
  assign \new_[45443]_  = ~A170 & \new_[45442]_ ;
  assign \new_[45447]_  = A200 & ~A199;
  assign \new_[45448]_  = ~A166 & \new_[45447]_ ;
  assign \new_[45449]_  = \new_[45448]_  & \new_[45443]_ ;
  assign \new_[45453]_  = ~A266 & ~A234;
  assign \new_[45454]_  = ~A233 & \new_[45453]_ ;
  assign \new_[45457]_  = ~A269 & ~A268;
  assign \new_[45460]_  = ~A299 & ~A298;
  assign \new_[45461]_  = \new_[45460]_  & \new_[45457]_ ;
  assign \new_[45462]_  = \new_[45461]_  & \new_[45454]_ ;
  assign \new_[45466]_  = A167 & ~A168;
  assign \new_[45467]_  = ~A170 & \new_[45466]_ ;
  assign \new_[45471]_  = A200 & ~A199;
  assign \new_[45472]_  = ~A166 & \new_[45471]_ ;
  assign \new_[45473]_  = \new_[45472]_  & \new_[45467]_ ;
  assign \new_[45477]_  = ~A266 & ~A234;
  assign \new_[45478]_  = ~A233 & \new_[45477]_ ;
  assign \new_[45481]_  = A298 & ~A267;
  assign \new_[45484]_  = ~A302 & ~A301;
  assign \new_[45485]_  = \new_[45484]_  & \new_[45481]_ ;
  assign \new_[45486]_  = \new_[45485]_  & \new_[45478]_ ;
  assign \new_[45490]_  = A167 & ~A168;
  assign \new_[45491]_  = ~A170 & \new_[45490]_ ;
  assign \new_[45495]_  = A200 & ~A199;
  assign \new_[45496]_  = ~A166 & \new_[45495]_ ;
  assign \new_[45497]_  = \new_[45496]_  & \new_[45491]_ ;
  assign \new_[45501]_  = ~A265 & ~A234;
  assign \new_[45502]_  = ~A233 & \new_[45501]_ ;
  assign \new_[45505]_  = A298 & ~A266;
  assign \new_[45508]_  = ~A302 & ~A301;
  assign \new_[45509]_  = \new_[45508]_  & \new_[45505]_ ;
  assign \new_[45510]_  = \new_[45509]_  & \new_[45502]_ ;
  assign \new_[45514]_  = A167 & ~A168;
  assign \new_[45515]_  = ~A170 & \new_[45514]_ ;
  assign \new_[45519]_  = A200 & ~A199;
  assign \new_[45520]_  = ~A166 & \new_[45519]_ ;
  assign \new_[45521]_  = \new_[45520]_  & \new_[45515]_ ;
  assign \new_[45525]_  = A265 & ~A233;
  assign \new_[45526]_  = ~A232 & \new_[45525]_ ;
  assign \new_[45529]_  = A298 & A266;
  assign \new_[45532]_  = ~A302 & ~A301;
  assign \new_[45533]_  = \new_[45532]_  & \new_[45529]_ ;
  assign \new_[45534]_  = \new_[45533]_  & \new_[45526]_ ;
  assign \new_[45538]_  = A167 & ~A168;
  assign \new_[45539]_  = ~A170 & \new_[45538]_ ;
  assign \new_[45543]_  = A200 & ~A199;
  assign \new_[45544]_  = ~A166 & \new_[45543]_ ;
  assign \new_[45545]_  = \new_[45544]_  & \new_[45539]_ ;
  assign \new_[45549]_  = ~A266 & ~A233;
  assign \new_[45550]_  = ~A232 & \new_[45549]_ ;
  assign \new_[45553]_  = ~A269 & ~A268;
  assign \new_[45556]_  = ~A300 & A298;
  assign \new_[45557]_  = \new_[45556]_  & \new_[45553]_ ;
  assign \new_[45558]_  = \new_[45557]_  & \new_[45550]_ ;
  assign \new_[45562]_  = A167 & ~A168;
  assign \new_[45563]_  = ~A170 & \new_[45562]_ ;
  assign \new_[45567]_  = A200 & ~A199;
  assign \new_[45568]_  = ~A166 & \new_[45567]_ ;
  assign \new_[45569]_  = \new_[45568]_  & \new_[45563]_ ;
  assign \new_[45573]_  = ~A266 & ~A233;
  assign \new_[45574]_  = ~A232 & \new_[45573]_ ;
  assign \new_[45577]_  = ~A269 & ~A268;
  assign \new_[45580]_  = A299 & A298;
  assign \new_[45581]_  = \new_[45580]_  & \new_[45577]_ ;
  assign \new_[45582]_  = \new_[45581]_  & \new_[45574]_ ;
  assign \new_[45586]_  = A167 & ~A168;
  assign \new_[45587]_  = ~A170 & \new_[45586]_ ;
  assign \new_[45591]_  = A200 & ~A199;
  assign \new_[45592]_  = ~A166 & \new_[45591]_ ;
  assign \new_[45593]_  = \new_[45592]_  & \new_[45587]_ ;
  assign \new_[45597]_  = ~A266 & ~A233;
  assign \new_[45598]_  = ~A232 & \new_[45597]_ ;
  assign \new_[45601]_  = ~A269 & ~A268;
  assign \new_[45604]_  = ~A299 & ~A298;
  assign \new_[45605]_  = \new_[45604]_  & \new_[45601]_ ;
  assign \new_[45606]_  = \new_[45605]_  & \new_[45598]_ ;
  assign \new_[45610]_  = A167 & ~A168;
  assign \new_[45611]_  = ~A170 & \new_[45610]_ ;
  assign \new_[45615]_  = A200 & ~A199;
  assign \new_[45616]_  = ~A166 & \new_[45615]_ ;
  assign \new_[45617]_  = \new_[45616]_  & \new_[45611]_ ;
  assign \new_[45621]_  = ~A266 & ~A233;
  assign \new_[45622]_  = ~A232 & \new_[45621]_ ;
  assign \new_[45625]_  = A298 & ~A267;
  assign \new_[45628]_  = ~A302 & ~A301;
  assign \new_[45629]_  = \new_[45628]_  & \new_[45625]_ ;
  assign \new_[45630]_  = \new_[45629]_  & \new_[45622]_ ;
  assign \new_[45634]_  = A167 & ~A168;
  assign \new_[45635]_  = ~A170 & \new_[45634]_ ;
  assign \new_[45639]_  = A200 & ~A199;
  assign \new_[45640]_  = ~A166 & \new_[45639]_ ;
  assign \new_[45641]_  = \new_[45640]_  & \new_[45635]_ ;
  assign \new_[45645]_  = ~A265 & ~A233;
  assign \new_[45646]_  = ~A232 & \new_[45645]_ ;
  assign \new_[45649]_  = A298 & ~A266;
  assign \new_[45652]_  = ~A302 & ~A301;
  assign \new_[45653]_  = \new_[45652]_  & \new_[45649]_ ;
  assign \new_[45654]_  = \new_[45653]_  & \new_[45646]_ ;
  assign \new_[45658]_  = ~A167 & ~A168;
  assign \new_[45659]_  = ~A170 & \new_[45658]_ ;
  assign \new_[45663]_  = A200 & ~A199;
  assign \new_[45664]_  = A166 & \new_[45663]_ ;
  assign \new_[45665]_  = \new_[45664]_  & \new_[45659]_ ;
  assign \new_[45669]_  = A265 & A233;
  assign \new_[45670]_  = A232 & \new_[45669]_ ;
  assign \new_[45673]_  = ~A269 & ~A268;
  assign \new_[45676]_  = ~A300 & ~A299;
  assign \new_[45677]_  = \new_[45676]_  & \new_[45673]_ ;
  assign \new_[45678]_  = \new_[45677]_  & \new_[45670]_ ;
  assign \new_[45682]_  = ~A167 & ~A168;
  assign \new_[45683]_  = ~A170 & \new_[45682]_ ;
  assign \new_[45687]_  = A200 & ~A199;
  assign \new_[45688]_  = A166 & \new_[45687]_ ;
  assign \new_[45689]_  = \new_[45688]_  & \new_[45683]_ ;
  assign \new_[45693]_  = A265 & A233;
  assign \new_[45694]_  = A232 & \new_[45693]_ ;
  assign \new_[45697]_  = ~A269 & ~A268;
  assign \new_[45700]_  = A299 & A298;
  assign \new_[45701]_  = \new_[45700]_  & \new_[45697]_ ;
  assign \new_[45702]_  = \new_[45701]_  & \new_[45694]_ ;
  assign \new_[45706]_  = ~A167 & ~A168;
  assign \new_[45707]_  = ~A170 & \new_[45706]_ ;
  assign \new_[45711]_  = A200 & ~A199;
  assign \new_[45712]_  = A166 & \new_[45711]_ ;
  assign \new_[45713]_  = \new_[45712]_  & \new_[45707]_ ;
  assign \new_[45717]_  = A265 & A233;
  assign \new_[45718]_  = A232 & \new_[45717]_ ;
  assign \new_[45721]_  = ~A269 & ~A268;
  assign \new_[45724]_  = ~A299 & ~A298;
  assign \new_[45725]_  = \new_[45724]_  & \new_[45721]_ ;
  assign \new_[45726]_  = \new_[45725]_  & \new_[45718]_ ;
  assign \new_[45730]_  = ~A167 & ~A168;
  assign \new_[45731]_  = ~A170 & \new_[45730]_ ;
  assign \new_[45735]_  = A200 & ~A199;
  assign \new_[45736]_  = A166 & \new_[45735]_ ;
  assign \new_[45737]_  = \new_[45736]_  & \new_[45731]_ ;
  assign \new_[45741]_  = A265 & A233;
  assign \new_[45742]_  = A232 & \new_[45741]_ ;
  assign \new_[45745]_  = ~A299 & ~A267;
  assign \new_[45748]_  = ~A302 & ~A301;
  assign \new_[45749]_  = \new_[45748]_  & \new_[45745]_ ;
  assign \new_[45750]_  = \new_[45749]_  & \new_[45742]_ ;
  assign \new_[45754]_  = ~A167 & ~A168;
  assign \new_[45755]_  = ~A170 & \new_[45754]_ ;
  assign \new_[45759]_  = A200 & ~A199;
  assign \new_[45760]_  = A166 & \new_[45759]_ ;
  assign \new_[45761]_  = \new_[45760]_  & \new_[45755]_ ;
  assign \new_[45765]_  = A265 & A233;
  assign \new_[45766]_  = A232 & \new_[45765]_ ;
  assign \new_[45769]_  = ~A299 & A266;
  assign \new_[45772]_  = ~A302 & ~A301;
  assign \new_[45773]_  = \new_[45772]_  & \new_[45769]_ ;
  assign \new_[45774]_  = \new_[45773]_  & \new_[45766]_ ;
  assign \new_[45778]_  = ~A167 & ~A168;
  assign \new_[45779]_  = ~A170 & \new_[45778]_ ;
  assign \new_[45783]_  = A200 & ~A199;
  assign \new_[45784]_  = A166 & \new_[45783]_ ;
  assign \new_[45785]_  = \new_[45784]_  & \new_[45779]_ ;
  assign \new_[45789]_  = ~A265 & A233;
  assign \new_[45790]_  = A232 & \new_[45789]_ ;
  assign \new_[45793]_  = ~A299 & ~A266;
  assign \new_[45796]_  = ~A302 & ~A301;
  assign \new_[45797]_  = \new_[45796]_  & \new_[45793]_ ;
  assign \new_[45798]_  = \new_[45797]_  & \new_[45790]_ ;
  assign \new_[45802]_  = ~A167 & ~A168;
  assign \new_[45803]_  = ~A170 & \new_[45802]_ ;
  assign \new_[45807]_  = A200 & ~A199;
  assign \new_[45808]_  = A166 & \new_[45807]_ ;
  assign \new_[45809]_  = \new_[45808]_  & \new_[45803]_ ;
  assign \new_[45813]_  = ~A236 & ~A235;
  assign \new_[45814]_  = ~A233 & \new_[45813]_ ;
  assign \new_[45817]_  = A266 & A265;
  assign \new_[45820]_  = ~A300 & A298;
  assign \new_[45821]_  = \new_[45820]_  & \new_[45817]_ ;
  assign \new_[45822]_  = \new_[45821]_  & \new_[45814]_ ;
  assign \new_[45826]_  = ~A167 & ~A168;
  assign \new_[45827]_  = ~A170 & \new_[45826]_ ;
  assign \new_[45831]_  = A200 & ~A199;
  assign \new_[45832]_  = A166 & \new_[45831]_ ;
  assign \new_[45833]_  = \new_[45832]_  & \new_[45827]_ ;
  assign \new_[45837]_  = ~A236 & ~A235;
  assign \new_[45838]_  = ~A233 & \new_[45837]_ ;
  assign \new_[45841]_  = A266 & A265;
  assign \new_[45844]_  = A299 & A298;
  assign \new_[45845]_  = \new_[45844]_  & \new_[45841]_ ;
  assign \new_[45846]_  = \new_[45845]_  & \new_[45838]_ ;
  assign \new_[45850]_  = ~A167 & ~A168;
  assign \new_[45851]_  = ~A170 & \new_[45850]_ ;
  assign \new_[45855]_  = A200 & ~A199;
  assign \new_[45856]_  = A166 & \new_[45855]_ ;
  assign \new_[45857]_  = \new_[45856]_  & \new_[45851]_ ;
  assign \new_[45861]_  = ~A236 & ~A235;
  assign \new_[45862]_  = ~A233 & \new_[45861]_ ;
  assign \new_[45865]_  = A266 & A265;
  assign \new_[45868]_  = ~A299 & ~A298;
  assign \new_[45869]_  = \new_[45868]_  & \new_[45865]_ ;
  assign \new_[45870]_  = \new_[45869]_  & \new_[45862]_ ;
  assign \new_[45874]_  = ~A167 & ~A168;
  assign \new_[45875]_  = ~A170 & \new_[45874]_ ;
  assign \new_[45879]_  = A200 & ~A199;
  assign \new_[45880]_  = A166 & \new_[45879]_ ;
  assign \new_[45881]_  = \new_[45880]_  & \new_[45875]_ ;
  assign \new_[45885]_  = ~A236 & ~A235;
  assign \new_[45886]_  = ~A233 & \new_[45885]_ ;
  assign \new_[45889]_  = ~A267 & ~A266;
  assign \new_[45892]_  = ~A300 & A298;
  assign \new_[45893]_  = \new_[45892]_  & \new_[45889]_ ;
  assign \new_[45894]_  = \new_[45893]_  & \new_[45886]_ ;
  assign \new_[45898]_  = ~A167 & ~A168;
  assign \new_[45899]_  = ~A170 & \new_[45898]_ ;
  assign \new_[45903]_  = A200 & ~A199;
  assign \new_[45904]_  = A166 & \new_[45903]_ ;
  assign \new_[45905]_  = \new_[45904]_  & \new_[45899]_ ;
  assign \new_[45909]_  = ~A236 & ~A235;
  assign \new_[45910]_  = ~A233 & \new_[45909]_ ;
  assign \new_[45913]_  = ~A267 & ~A266;
  assign \new_[45916]_  = A299 & A298;
  assign \new_[45917]_  = \new_[45916]_  & \new_[45913]_ ;
  assign \new_[45918]_  = \new_[45917]_  & \new_[45910]_ ;
  assign \new_[45922]_  = ~A167 & ~A168;
  assign \new_[45923]_  = ~A170 & \new_[45922]_ ;
  assign \new_[45927]_  = A200 & ~A199;
  assign \new_[45928]_  = A166 & \new_[45927]_ ;
  assign \new_[45929]_  = \new_[45928]_  & \new_[45923]_ ;
  assign \new_[45933]_  = ~A236 & ~A235;
  assign \new_[45934]_  = ~A233 & \new_[45933]_ ;
  assign \new_[45937]_  = ~A267 & ~A266;
  assign \new_[45940]_  = ~A299 & ~A298;
  assign \new_[45941]_  = \new_[45940]_  & \new_[45937]_ ;
  assign \new_[45942]_  = \new_[45941]_  & \new_[45934]_ ;
  assign \new_[45946]_  = ~A167 & ~A168;
  assign \new_[45947]_  = ~A170 & \new_[45946]_ ;
  assign \new_[45951]_  = A200 & ~A199;
  assign \new_[45952]_  = A166 & \new_[45951]_ ;
  assign \new_[45953]_  = \new_[45952]_  & \new_[45947]_ ;
  assign \new_[45957]_  = ~A236 & ~A235;
  assign \new_[45958]_  = ~A233 & \new_[45957]_ ;
  assign \new_[45961]_  = ~A266 & ~A265;
  assign \new_[45964]_  = ~A300 & A298;
  assign \new_[45965]_  = \new_[45964]_  & \new_[45961]_ ;
  assign \new_[45966]_  = \new_[45965]_  & \new_[45958]_ ;
  assign \new_[45970]_  = ~A167 & ~A168;
  assign \new_[45971]_  = ~A170 & \new_[45970]_ ;
  assign \new_[45975]_  = A200 & ~A199;
  assign \new_[45976]_  = A166 & \new_[45975]_ ;
  assign \new_[45977]_  = \new_[45976]_  & \new_[45971]_ ;
  assign \new_[45981]_  = ~A236 & ~A235;
  assign \new_[45982]_  = ~A233 & \new_[45981]_ ;
  assign \new_[45985]_  = ~A266 & ~A265;
  assign \new_[45988]_  = A299 & A298;
  assign \new_[45989]_  = \new_[45988]_  & \new_[45985]_ ;
  assign \new_[45990]_  = \new_[45989]_  & \new_[45982]_ ;
  assign \new_[45994]_  = ~A167 & ~A168;
  assign \new_[45995]_  = ~A170 & \new_[45994]_ ;
  assign \new_[45999]_  = A200 & ~A199;
  assign \new_[46000]_  = A166 & \new_[45999]_ ;
  assign \new_[46001]_  = \new_[46000]_  & \new_[45995]_ ;
  assign \new_[46005]_  = ~A236 & ~A235;
  assign \new_[46006]_  = ~A233 & \new_[46005]_ ;
  assign \new_[46009]_  = ~A266 & ~A265;
  assign \new_[46012]_  = ~A299 & ~A298;
  assign \new_[46013]_  = \new_[46012]_  & \new_[46009]_ ;
  assign \new_[46014]_  = \new_[46013]_  & \new_[46006]_ ;
  assign \new_[46018]_  = ~A167 & ~A168;
  assign \new_[46019]_  = ~A170 & \new_[46018]_ ;
  assign \new_[46023]_  = A200 & ~A199;
  assign \new_[46024]_  = A166 & \new_[46023]_ ;
  assign \new_[46025]_  = \new_[46024]_  & \new_[46019]_ ;
  assign \new_[46029]_  = A265 & ~A234;
  assign \new_[46030]_  = ~A233 & \new_[46029]_ ;
  assign \new_[46033]_  = A298 & A266;
  assign \new_[46036]_  = ~A302 & ~A301;
  assign \new_[46037]_  = \new_[46036]_  & \new_[46033]_ ;
  assign \new_[46038]_  = \new_[46037]_  & \new_[46030]_ ;
  assign \new_[46042]_  = ~A167 & ~A168;
  assign \new_[46043]_  = ~A170 & \new_[46042]_ ;
  assign \new_[46047]_  = A200 & ~A199;
  assign \new_[46048]_  = A166 & \new_[46047]_ ;
  assign \new_[46049]_  = \new_[46048]_  & \new_[46043]_ ;
  assign \new_[46053]_  = ~A266 & ~A234;
  assign \new_[46054]_  = ~A233 & \new_[46053]_ ;
  assign \new_[46057]_  = ~A269 & ~A268;
  assign \new_[46060]_  = ~A300 & A298;
  assign \new_[46061]_  = \new_[46060]_  & \new_[46057]_ ;
  assign \new_[46062]_  = \new_[46061]_  & \new_[46054]_ ;
  assign \new_[46066]_  = ~A167 & ~A168;
  assign \new_[46067]_  = ~A170 & \new_[46066]_ ;
  assign \new_[46071]_  = A200 & ~A199;
  assign \new_[46072]_  = A166 & \new_[46071]_ ;
  assign \new_[46073]_  = \new_[46072]_  & \new_[46067]_ ;
  assign \new_[46077]_  = ~A266 & ~A234;
  assign \new_[46078]_  = ~A233 & \new_[46077]_ ;
  assign \new_[46081]_  = ~A269 & ~A268;
  assign \new_[46084]_  = A299 & A298;
  assign \new_[46085]_  = \new_[46084]_  & \new_[46081]_ ;
  assign \new_[46086]_  = \new_[46085]_  & \new_[46078]_ ;
  assign \new_[46090]_  = ~A167 & ~A168;
  assign \new_[46091]_  = ~A170 & \new_[46090]_ ;
  assign \new_[46095]_  = A200 & ~A199;
  assign \new_[46096]_  = A166 & \new_[46095]_ ;
  assign \new_[46097]_  = \new_[46096]_  & \new_[46091]_ ;
  assign \new_[46101]_  = ~A266 & ~A234;
  assign \new_[46102]_  = ~A233 & \new_[46101]_ ;
  assign \new_[46105]_  = ~A269 & ~A268;
  assign \new_[46108]_  = ~A299 & ~A298;
  assign \new_[46109]_  = \new_[46108]_  & \new_[46105]_ ;
  assign \new_[46110]_  = \new_[46109]_  & \new_[46102]_ ;
  assign \new_[46114]_  = ~A167 & ~A168;
  assign \new_[46115]_  = ~A170 & \new_[46114]_ ;
  assign \new_[46119]_  = A200 & ~A199;
  assign \new_[46120]_  = A166 & \new_[46119]_ ;
  assign \new_[46121]_  = \new_[46120]_  & \new_[46115]_ ;
  assign \new_[46125]_  = ~A266 & ~A234;
  assign \new_[46126]_  = ~A233 & \new_[46125]_ ;
  assign \new_[46129]_  = A298 & ~A267;
  assign \new_[46132]_  = ~A302 & ~A301;
  assign \new_[46133]_  = \new_[46132]_  & \new_[46129]_ ;
  assign \new_[46134]_  = \new_[46133]_  & \new_[46126]_ ;
  assign \new_[46138]_  = ~A167 & ~A168;
  assign \new_[46139]_  = ~A170 & \new_[46138]_ ;
  assign \new_[46143]_  = A200 & ~A199;
  assign \new_[46144]_  = A166 & \new_[46143]_ ;
  assign \new_[46145]_  = \new_[46144]_  & \new_[46139]_ ;
  assign \new_[46149]_  = ~A265 & ~A234;
  assign \new_[46150]_  = ~A233 & \new_[46149]_ ;
  assign \new_[46153]_  = A298 & ~A266;
  assign \new_[46156]_  = ~A302 & ~A301;
  assign \new_[46157]_  = \new_[46156]_  & \new_[46153]_ ;
  assign \new_[46158]_  = \new_[46157]_  & \new_[46150]_ ;
  assign \new_[46162]_  = ~A167 & ~A168;
  assign \new_[46163]_  = ~A170 & \new_[46162]_ ;
  assign \new_[46167]_  = A200 & ~A199;
  assign \new_[46168]_  = A166 & \new_[46167]_ ;
  assign \new_[46169]_  = \new_[46168]_  & \new_[46163]_ ;
  assign \new_[46173]_  = A265 & ~A233;
  assign \new_[46174]_  = ~A232 & \new_[46173]_ ;
  assign \new_[46177]_  = A298 & A266;
  assign \new_[46180]_  = ~A302 & ~A301;
  assign \new_[46181]_  = \new_[46180]_  & \new_[46177]_ ;
  assign \new_[46182]_  = \new_[46181]_  & \new_[46174]_ ;
  assign \new_[46186]_  = ~A167 & ~A168;
  assign \new_[46187]_  = ~A170 & \new_[46186]_ ;
  assign \new_[46191]_  = A200 & ~A199;
  assign \new_[46192]_  = A166 & \new_[46191]_ ;
  assign \new_[46193]_  = \new_[46192]_  & \new_[46187]_ ;
  assign \new_[46197]_  = ~A266 & ~A233;
  assign \new_[46198]_  = ~A232 & \new_[46197]_ ;
  assign \new_[46201]_  = ~A269 & ~A268;
  assign \new_[46204]_  = ~A300 & A298;
  assign \new_[46205]_  = \new_[46204]_  & \new_[46201]_ ;
  assign \new_[46206]_  = \new_[46205]_  & \new_[46198]_ ;
  assign \new_[46210]_  = ~A167 & ~A168;
  assign \new_[46211]_  = ~A170 & \new_[46210]_ ;
  assign \new_[46215]_  = A200 & ~A199;
  assign \new_[46216]_  = A166 & \new_[46215]_ ;
  assign \new_[46217]_  = \new_[46216]_  & \new_[46211]_ ;
  assign \new_[46221]_  = ~A266 & ~A233;
  assign \new_[46222]_  = ~A232 & \new_[46221]_ ;
  assign \new_[46225]_  = ~A269 & ~A268;
  assign \new_[46228]_  = A299 & A298;
  assign \new_[46229]_  = \new_[46228]_  & \new_[46225]_ ;
  assign \new_[46230]_  = \new_[46229]_  & \new_[46222]_ ;
  assign \new_[46234]_  = ~A167 & ~A168;
  assign \new_[46235]_  = ~A170 & \new_[46234]_ ;
  assign \new_[46239]_  = A200 & ~A199;
  assign \new_[46240]_  = A166 & \new_[46239]_ ;
  assign \new_[46241]_  = \new_[46240]_  & \new_[46235]_ ;
  assign \new_[46245]_  = ~A266 & ~A233;
  assign \new_[46246]_  = ~A232 & \new_[46245]_ ;
  assign \new_[46249]_  = ~A269 & ~A268;
  assign \new_[46252]_  = ~A299 & ~A298;
  assign \new_[46253]_  = \new_[46252]_  & \new_[46249]_ ;
  assign \new_[46254]_  = \new_[46253]_  & \new_[46246]_ ;
  assign \new_[46258]_  = ~A167 & ~A168;
  assign \new_[46259]_  = ~A170 & \new_[46258]_ ;
  assign \new_[46263]_  = A200 & ~A199;
  assign \new_[46264]_  = A166 & \new_[46263]_ ;
  assign \new_[46265]_  = \new_[46264]_  & \new_[46259]_ ;
  assign \new_[46269]_  = ~A266 & ~A233;
  assign \new_[46270]_  = ~A232 & \new_[46269]_ ;
  assign \new_[46273]_  = A298 & ~A267;
  assign \new_[46276]_  = ~A302 & ~A301;
  assign \new_[46277]_  = \new_[46276]_  & \new_[46273]_ ;
  assign \new_[46278]_  = \new_[46277]_  & \new_[46270]_ ;
  assign \new_[46282]_  = ~A167 & ~A168;
  assign \new_[46283]_  = ~A170 & \new_[46282]_ ;
  assign \new_[46287]_  = A200 & ~A199;
  assign \new_[46288]_  = A166 & \new_[46287]_ ;
  assign \new_[46289]_  = \new_[46288]_  & \new_[46283]_ ;
  assign \new_[46293]_  = ~A265 & ~A233;
  assign \new_[46294]_  = ~A232 & \new_[46293]_ ;
  assign \new_[46297]_  = A298 & ~A266;
  assign \new_[46300]_  = ~A302 & ~A301;
  assign \new_[46301]_  = \new_[46300]_  & \new_[46297]_ ;
  assign \new_[46302]_  = \new_[46301]_  & \new_[46294]_ ;
  assign \new_[46306]_  = A167 & ~A168;
  assign \new_[46307]_  = A169 & \new_[46306]_ ;
  assign \new_[46311]_  = A200 & ~A199;
  assign \new_[46312]_  = ~A166 & \new_[46311]_ ;
  assign \new_[46313]_  = \new_[46312]_  & \new_[46307]_ ;
  assign \new_[46317]_  = A265 & A233;
  assign \new_[46318]_  = A232 & \new_[46317]_ ;
  assign \new_[46321]_  = ~A269 & ~A268;
  assign \new_[46324]_  = ~A300 & ~A299;
  assign \new_[46325]_  = \new_[46324]_  & \new_[46321]_ ;
  assign \new_[46326]_  = \new_[46325]_  & \new_[46318]_ ;
  assign \new_[46330]_  = A167 & ~A168;
  assign \new_[46331]_  = A169 & \new_[46330]_ ;
  assign \new_[46335]_  = A200 & ~A199;
  assign \new_[46336]_  = ~A166 & \new_[46335]_ ;
  assign \new_[46337]_  = \new_[46336]_  & \new_[46331]_ ;
  assign \new_[46341]_  = A265 & A233;
  assign \new_[46342]_  = A232 & \new_[46341]_ ;
  assign \new_[46345]_  = ~A269 & ~A268;
  assign \new_[46348]_  = A299 & A298;
  assign \new_[46349]_  = \new_[46348]_  & \new_[46345]_ ;
  assign \new_[46350]_  = \new_[46349]_  & \new_[46342]_ ;
  assign \new_[46354]_  = A167 & ~A168;
  assign \new_[46355]_  = A169 & \new_[46354]_ ;
  assign \new_[46359]_  = A200 & ~A199;
  assign \new_[46360]_  = ~A166 & \new_[46359]_ ;
  assign \new_[46361]_  = \new_[46360]_  & \new_[46355]_ ;
  assign \new_[46365]_  = A265 & A233;
  assign \new_[46366]_  = A232 & \new_[46365]_ ;
  assign \new_[46369]_  = ~A269 & ~A268;
  assign \new_[46372]_  = ~A299 & ~A298;
  assign \new_[46373]_  = \new_[46372]_  & \new_[46369]_ ;
  assign \new_[46374]_  = \new_[46373]_  & \new_[46366]_ ;
  assign \new_[46378]_  = A167 & ~A168;
  assign \new_[46379]_  = A169 & \new_[46378]_ ;
  assign \new_[46383]_  = A200 & ~A199;
  assign \new_[46384]_  = ~A166 & \new_[46383]_ ;
  assign \new_[46385]_  = \new_[46384]_  & \new_[46379]_ ;
  assign \new_[46389]_  = A265 & A233;
  assign \new_[46390]_  = A232 & \new_[46389]_ ;
  assign \new_[46393]_  = ~A299 & ~A267;
  assign \new_[46396]_  = ~A302 & ~A301;
  assign \new_[46397]_  = \new_[46396]_  & \new_[46393]_ ;
  assign \new_[46398]_  = \new_[46397]_  & \new_[46390]_ ;
  assign \new_[46402]_  = A167 & ~A168;
  assign \new_[46403]_  = A169 & \new_[46402]_ ;
  assign \new_[46407]_  = A200 & ~A199;
  assign \new_[46408]_  = ~A166 & \new_[46407]_ ;
  assign \new_[46409]_  = \new_[46408]_  & \new_[46403]_ ;
  assign \new_[46413]_  = A265 & A233;
  assign \new_[46414]_  = A232 & \new_[46413]_ ;
  assign \new_[46417]_  = ~A299 & A266;
  assign \new_[46420]_  = ~A302 & ~A301;
  assign \new_[46421]_  = \new_[46420]_  & \new_[46417]_ ;
  assign \new_[46422]_  = \new_[46421]_  & \new_[46414]_ ;
  assign \new_[46426]_  = A167 & ~A168;
  assign \new_[46427]_  = A169 & \new_[46426]_ ;
  assign \new_[46431]_  = A200 & ~A199;
  assign \new_[46432]_  = ~A166 & \new_[46431]_ ;
  assign \new_[46433]_  = \new_[46432]_  & \new_[46427]_ ;
  assign \new_[46437]_  = ~A265 & A233;
  assign \new_[46438]_  = A232 & \new_[46437]_ ;
  assign \new_[46441]_  = ~A299 & ~A266;
  assign \new_[46444]_  = ~A302 & ~A301;
  assign \new_[46445]_  = \new_[46444]_  & \new_[46441]_ ;
  assign \new_[46446]_  = \new_[46445]_  & \new_[46438]_ ;
  assign \new_[46450]_  = A167 & ~A168;
  assign \new_[46451]_  = A169 & \new_[46450]_ ;
  assign \new_[46455]_  = A200 & ~A199;
  assign \new_[46456]_  = ~A166 & \new_[46455]_ ;
  assign \new_[46457]_  = \new_[46456]_  & \new_[46451]_ ;
  assign \new_[46461]_  = ~A236 & ~A235;
  assign \new_[46462]_  = ~A233 & \new_[46461]_ ;
  assign \new_[46465]_  = A266 & A265;
  assign \new_[46468]_  = ~A300 & A298;
  assign \new_[46469]_  = \new_[46468]_  & \new_[46465]_ ;
  assign \new_[46470]_  = \new_[46469]_  & \new_[46462]_ ;
  assign \new_[46474]_  = A167 & ~A168;
  assign \new_[46475]_  = A169 & \new_[46474]_ ;
  assign \new_[46479]_  = A200 & ~A199;
  assign \new_[46480]_  = ~A166 & \new_[46479]_ ;
  assign \new_[46481]_  = \new_[46480]_  & \new_[46475]_ ;
  assign \new_[46485]_  = ~A236 & ~A235;
  assign \new_[46486]_  = ~A233 & \new_[46485]_ ;
  assign \new_[46489]_  = A266 & A265;
  assign \new_[46492]_  = A299 & A298;
  assign \new_[46493]_  = \new_[46492]_  & \new_[46489]_ ;
  assign \new_[46494]_  = \new_[46493]_  & \new_[46486]_ ;
  assign \new_[46498]_  = A167 & ~A168;
  assign \new_[46499]_  = A169 & \new_[46498]_ ;
  assign \new_[46503]_  = A200 & ~A199;
  assign \new_[46504]_  = ~A166 & \new_[46503]_ ;
  assign \new_[46505]_  = \new_[46504]_  & \new_[46499]_ ;
  assign \new_[46509]_  = ~A236 & ~A235;
  assign \new_[46510]_  = ~A233 & \new_[46509]_ ;
  assign \new_[46513]_  = A266 & A265;
  assign \new_[46516]_  = ~A299 & ~A298;
  assign \new_[46517]_  = \new_[46516]_  & \new_[46513]_ ;
  assign \new_[46518]_  = \new_[46517]_  & \new_[46510]_ ;
  assign \new_[46522]_  = A167 & ~A168;
  assign \new_[46523]_  = A169 & \new_[46522]_ ;
  assign \new_[46527]_  = A200 & ~A199;
  assign \new_[46528]_  = ~A166 & \new_[46527]_ ;
  assign \new_[46529]_  = \new_[46528]_  & \new_[46523]_ ;
  assign \new_[46533]_  = ~A236 & ~A235;
  assign \new_[46534]_  = ~A233 & \new_[46533]_ ;
  assign \new_[46537]_  = ~A267 & ~A266;
  assign \new_[46540]_  = ~A300 & A298;
  assign \new_[46541]_  = \new_[46540]_  & \new_[46537]_ ;
  assign \new_[46542]_  = \new_[46541]_  & \new_[46534]_ ;
  assign \new_[46546]_  = A167 & ~A168;
  assign \new_[46547]_  = A169 & \new_[46546]_ ;
  assign \new_[46551]_  = A200 & ~A199;
  assign \new_[46552]_  = ~A166 & \new_[46551]_ ;
  assign \new_[46553]_  = \new_[46552]_  & \new_[46547]_ ;
  assign \new_[46557]_  = ~A236 & ~A235;
  assign \new_[46558]_  = ~A233 & \new_[46557]_ ;
  assign \new_[46561]_  = ~A267 & ~A266;
  assign \new_[46564]_  = A299 & A298;
  assign \new_[46565]_  = \new_[46564]_  & \new_[46561]_ ;
  assign \new_[46566]_  = \new_[46565]_  & \new_[46558]_ ;
  assign \new_[46570]_  = A167 & ~A168;
  assign \new_[46571]_  = A169 & \new_[46570]_ ;
  assign \new_[46575]_  = A200 & ~A199;
  assign \new_[46576]_  = ~A166 & \new_[46575]_ ;
  assign \new_[46577]_  = \new_[46576]_  & \new_[46571]_ ;
  assign \new_[46581]_  = ~A236 & ~A235;
  assign \new_[46582]_  = ~A233 & \new_[46581]_ ;
  assign \new_[46585]_  = ~A267 & ~A266;
  assign \new_[46588]_  = ~A299 & ~A298;
  assign \new_[46589]_  = \new_[46588]_  & \new_[46585]_ ;
  assign \new_[46590]_  = \new_[46589]_  & \new_[46582]_ ;
  assign \new_[46594]_  = A167 & ~A168;
  assign \new_[46595]_  = A169 & \new_[46594]_ ;
  assign \new_[46599]_  = A200 & ~A199;
  assign \new_[46600]_  = ~A166 & \new_[46599]_ ;
  assign \new_[46601]_  = \new_[46600]_  & \new_[46595]_ ;
  assign \new_[46605]_  = ~A236 & ~A235;
  assign \new_[46606]_  = ~A233 & \new_[46605]_ ;
  assign \new_[46609]_  = ~A266 & ~A265;
  assign \new_[46612]_  = ~A300 & A298;
  assign \new_[46613]_  = \new_[46612]_  & \new_[46609]_ ;
  assign \new_[46614]_  = \new_[46613]_  & \new_[46606]_ ;
  assign \new_[46618]_  = A167 & ~A168;
  assign \new_[46619]_  = A169 & \new_[46618]_ ;
  assign \new_[46623]_  = A200 & ~A199;
  assign \new_[46624]_  = ~A166 & \new_[46623]_ ;
  assign \new_[46625]_  = \new_[46624]_  & \new_[46619]_ ;
  assign \new_[46629]_  = ~A236 & ~A235;
  assign \new_[46630]_  = ~A233 & \new_[46629]_ ;
  assign \new_[46633]_  = ~A266 & ~A265;
  assign \new_[46636]_  = A299 & A298;
  assign \new_[46637]_  = \new_[46636]_  & \new_[46633]_ ;
  assign \new_[46638]_  = \new_[46637]_  & \new_[46630]_ ;
  assign \new_[46642]_  = A167 & ~A168;
  assign \new_[46643]_  = A169 & \new_[46642]_ ;
  assign \new_[46647]_  = A200 & ~A199;
  assign \new_[46648]_  = ~A166 & \new_[46647]_ ;
  assign \new_[46649]_  = \new_[46648]_  & \new_[46643]_ ;
  assign \new_[46653]_  = ~A236 & ~A235;
  assign \new_[46654]_  = ~A233 & \new_[46653]_ ;
  assign \new_[46657]_  = ~A266 & ~A265;
  assign \new_[46660]_  = ~A299 & ~A298;
  assign \new_[46661]_  = \new_[46660]_  & \new_[46657]_ ;
  assign \new_[46662]_  = \new_[46661]_  & \new_[46654]_ ;
  assign \new_[46666]_  = A167 & ~A168;
  assign \new_[46667]_  = A169 & \new_[46666]_ ;
  assign \new_[46671]_  = A200 & ~A199;
  assign \new_[46672]_  = ~A166 & \new_[46671]_ ;
  assign \new_[46673]_  = \new_[46672]_  & \new_[46667]_ ;
  assign \new_[46677]_  = A265 & ~A234;
  assign \new_[46678]_  = ~A233 & \new_[46677]_ ;
  assign \new_[46681]_  = A298 & A266;
  assign \new_[46684]_  = ~A302 & ~A301;
  assign \new_[46685]_  = \new_[46684]_  & \new_[46681]_ ;
  assign \new_[46686]_  = \new_[46685]_  & \new_[46678]_ ;
  assign \new_[46690]_  = A167 & ~A168;
  assign \new_[46691]_  = A169 & \new_[46690]_ ;
  assign \new_[46695]_  = A200 & ~A199;
  assign \new_[46696]_  = ~A166 & \new_[46695]_ ;
  assign \new_[46697]_  = \new_[46696]_  & \new_[46691]_ ;
  assign \new_[46701]_  = ~A266 & ~A234;
  assign \new_[46702]_  = ~A233 & \new_[46701]_ ;
  assign \new_[46705]_  = ~A269 & ~A268;
  assign \new_[46708]_  = ~A300 & A298;
  assign \new_[46709]_  = \new_[46708]_  & \new_[46705]_ ;
  assign \new_[46710]_  = \new_[46709]_  & \new_[46702]_ ;
  assign \new_[46714]_  = A167 & ~A168;
  assign \new_[46715]_  = A169 & \new_[46714]_ ;
  assign \new_[46719]_  = A200 & ~A199;
  assign \new_[46720]_  = ~A166 & \new_[46719]_ ;
  assign \new_[46721]_  = \new_[46720]_  & \new_[46715]_ ;
  assign \new_[46725]_  = ~A266 & ~A234;
  assign \new_[46726]_  = ~A233 & \new_[46725]_ ;
  assign \new_[46729]_  = ~A269 & ~A268;
  assign \new_[46732]_  = A299 & A298;
  assign \new_[46733]_  = \new_[46732]_  & \new_[46729]_ ;
  assign \new_[46734]_  = \new_[46733]_  & \new_[46726]_ ;
  assign \new_[46738]_  = A167 & ~A168;
  assign \new_[46739]_  = A169 & \new_[46738]_ ;
  assign \new_[46743]_  = A200 & ~A199;
  assign \new_[46744]_  = ~A166 & \new_[46743]_ ;
  assign \new_[46745]_  = \new_[46744]_  & \new_[46739]_ ;
  assign \new_[46749]_  = ~A266 & ~A234;
  assign \new_[46750]_  = ~A233 & \new_[46749]_ ;
  assign \new_[46753]_  = ~A269 & ~A268;
  assign \new_[46756]_  = ~A299 & ~A298;
  assign \new_[46757]_  = \new_[46756]_  & \new_[46753]_ ;
  assign \new_[46758]_  = \new_[46757]_  & \new_[46750]_ ;
  assign \new_[46762]_  = A167 & ~A168;
  assign \new_[46763]_  = A169 & \new_[46762]_ ;
  assign \new_[46767]_  = A200 & ~A199;
  assign \new_[46768]_  = ~A166 & \new_[46767]_ ;
  assign \new_[46769]_  = \new_[46768]_  & \new_[46763]_ ;
  assign \new_[46773]_  = ~A266 & ~A234;
  assign \new_[46774]_  = ~A233 & \new_[46773]_ ;
  assign \new_[46777]_  = A298 & ~A267;
  assign \new_[46780]_  = ~A302 & ~A301;
  assign \new_[46781]_  = \new_[46780]_  & \new_[46777]_ ;
  assign \new_[46782]_  = \new_[46781]_  & \new_[46774]_ ;
  assign \new_[46786]_  = A167 & ~A168;
  assign \new_[46787]_  = A169 & \new_[46786]_ ;
  assign \new_[46791]_  = A200 & ~A199;
  assign \new_[46792]_  = ~A166 & \new_[46791]_ ;
  assign \new_[46793]_  = \new_[46792]_  & \new_[46787]_ ;
  assign \new_[46797]_  = ~A265 & ~A234;
  assign \new_[46798]_  = ~A233 & \new_[46797]_ ;
  assign \new_[46801]_  = A298 & ~A266;
  assign \new_[46804]_  = ~A302 & ~A301;
  assign \new_[46805]_  = \new_[46804]_  & \new_[46801]_ ;
  assign \new_[46806]_  = \new_[46805]_  & \new_[46798]_ ;
  assign \new_[46810]_  = A167 & ~A168;
  assign \new_[46811]_  = A169 & \new_[46810]_ ;
  assign \new_[46815]_  = A200 & ~A199;
  assign \new_[46816]_  = ~A166 & \new_[46815]_ ;
  assign \new_[46817]_  = \new_[46816]_  & \new_[46811]_ ;
  assign \new_[46821]_  = A265 & ~A233;
  assign \new_[46822]_  = ~A232 & \new_[46821]_ ;
  assign \new_[46825]_  = A298 & A266;
  assign \new_[46828]_  = ~A302 & ~A301;
  assign \new_[46829]_  = \new_[46828]_  & \new_[46825]_ ;
  assign \new_[46830]_  = \new_[46829]_  & \new_[46822]_ ;
  assign \new_[46834]_  = A167 & ~A168;
  assign \new_[46835]_  = A169 & \new_[46834]_ ;
  assign \new_[46839]_  = A200 & ~A199;
  assign \new_[46840]_  = ~A166 & \new_[46839]_ ;
  assign \new_[46841]_  = \new_[46840]_  & \new_[46835]_ ;
  assign \new_[46845]_  = ~A266 & ~A233;
  assign \new_[46846]_  = ~A232 & \new_[46845]_ ;
  assign \new_[46849]_  = ~A269 & ~A268;
  assign \new_[46852]_  = ~A300 & A298;
  assign \new_[46853]_  = \new_[46852]_  & \new_[46849]_ ;
  assign \new_[46854]_  = \new_[46853]_  & \new_[46846]_ ;
  assign \new_[46858]_  = A167 & ~A168;
  assign \new_[46859]_  = A169 & \new_[46858]_ ;
  assign \new_[46863]_  = A200 & ~A199;
  assign \new_[46864]_  = ~A166 & \new_[46863]_ ;
  assign \new_[46865]_  = \new_[46864]_  & \new_[46859]_ ;
  assign \new_[46869]_  = ~A266 & ~A233;
  assign \new_[46870]_  = ~A232 & \new_[46869]_ ;
  assign \new_[46873]_  = ~A269 & ~A268;
  assign \new_[46876]_  = A299 & A298;
  assign \new_[46877]_  = \new_[46876]_  & \new_[46873]_ ;
  assign \new_[46878]_  = \new_[46877]_  & \new_[46870]_ ;
  assign \new_[46882]_  = A167 & ~A168;
  assign \new_[46883]_  = A169 & \new_[46882]_ ;
  assign \new_[46887]_  = A200 & ~A199;
  assign \new_[46888]_  = ~A166 & \new_[46887]_ ;
  assign \new_[46889]_  = \new_[46888]_  & \new_[46883]_ ;
  assign \new_[46893]_  = ~A266 & ~A233;
  assign \new_[46894]_  = ~A232 & \new_[46893]_ ;
  assign \new_[46897]_  = ~A269 & ~A268;
  assign \new_[46900]_  = ~A299 & ~A298;
  assign \new_[46901]_  = \new_[46900]_  & \new_[46897]_ ;
  assign \new_[46902]_  = \new_[46901]_  & \new_[46894]_ ;
  assign \new_[46906]_  = A167 & ~A168;
  assign \new_[46907]_  = A169 & \new_[46906]_ ;
  assign \new_[46911]_  = A200 & ~A199;
  assign \new_[46912]_  = ~A166 & \new_[46911]_ ;
  assign \new_[46913]_  = \new_[46912]_  & \new_[46907]_ ;
  assign \new_[46917]_  = ~A266 & ~A233;
  assign \new_[46918]_  = ~A232 & \new_[46917]_ ;
  assign \new_[46921]_  = A298 & ~A267;
  assign \new_[46924]_  = ~A302 & ~A301;
  assign \new_[46925]_  = \new_[46924]_  & \new_[46921]_ ;
  assign \new_[46926]_  = \new_[46925]_  & \new_[46918]_ ;
  assign \new_[46930]_  = A167 & ~A168;
  assign \new_[46931]_  = A169 & \new_[46930]_ ;
  assign \new_[46935]_  = A200 & ~A199;
  assign \new_[46936]_  = ~A166 & \new_[46935]_ ;
  assign \new_[46937]_  = \new_[46936]_  & \new_[46931]_ ;
  assign \new_[46941]_  = ~A265 & ~A233;
  assign \new_[46942]_  = ~A232 & \new_[46941]_ ;
  assign \new_[46945]_  = A298 & ~A266;
  assign \new_[46948]_  = ~A302 & ~A301;
  assign \new_[46949]_  = \new_[46948]_  & \new_[46945]_ ;
  assign \new_[46950]_  = \new_[46949]_  & \new_[46942]_ ;
  assign \new_[46954]_  = ~A167 & ~A168;
  assign \new_[46955]_  = A169 & \new_[46954]_ ;
  assign \new_[46959]_  = A200 & ~A199;
  assign \new_[46960]_  = A166 & \new_[46959]_ ;
  assign \new_[46961]_  = \new_[46960]_  & \new_[46955]_ ;
  assign \new_[46965]_  = A265 & A233;
  assign \new_[46966]_  = A232 & \new_[46965]_ ;
  assign \new_[46969]_  = ~A269 & ~A268;
  assign \new_[46972]_  = ~A300 & ~A299;
  assign \new_[46973]_  = \new_[46972]_  & \new_[46969]_ ;
  assign \new_[46974]_  = \new_[46973]_  & \new_[46966]_ ;
  assign \new_[46978]_  = ~A167 & ~A168;
  assign \new_[46979]_  = A169 & \new_[46978]_ ;
  assign \new_[46983]_  = A200 & ~A199;
  assign \new_[46984]_  = A166 & \new_[46983]_ ;
  assign \new_[46985]_  = \new_[46984]_  & \new_[46979]_ ;
  assign \new_[46989]_  = A265 & A233;
  assign \new_[46990]_  = A232 & \new_[46989]_ ;
  assign \new_[46993]_  = ~A269 & ~A268;
  assign \new_[46996]_  = A299 & A298;
  assign \new_[46997]_  = \new_[46996]_  & \new_[46993]_ ;
  assign \new_[46998]_  = \new_[46997]_  & \new_[46990]_ ;
  assign \new_[47002]_  = ~A167 & ~A168;
  assign \new_[47003]_  = A169 & \new_[47002]_ ;
  assign \new_[47007]_  = A200 & ~A199;
  assign \new_[47008]_  = A166 & \new_[47007]_ ;
  assign \new_[47009]_  = \new_[47008]_  & \new_[47003]_ ;
  assign \new_[47013]_  = A265 & A233;
  assign \new_[47014]_  = A232 & \new_[47013]_ ;
  assign \new_[47017]_  = ~A269 & ~A268;
  assign \new_[47020]_  = ~A299 & ~A298;
  assign \new_[47021]_  = \new_[47020]_  & \new_[47017]_ ;
  assign \new_[47022]_  = \new_[47021]_  & \new_[47014]_ ;
  assign \new_[47026]_  = ~A167 & ~A168;
  assign \new_[47027]_  = A169 & \new_[47026]_ ;
  assign \new_[47031]_  = A200 & ~A199;
  assign \new_[47032]_  = A166 & \new_[47031]_ ;
  assign \new_[47033]_  = \new_[47032]_  & \new_[47027]_ ;
  assign \new_[47037]_  = A265 & A233;
  assign \new_[47038]_  = A232 & \new_[47037]_ ;
  assign \new_[47041]_  = ~A299 & ~A267;
  assign \new_[47044]_  = ~A302 & ~A301;
  assign \new_[47045]_  = \new_[47044]_  & \new_[47041]_ ;
  assign \new_[47046]_  = \new_[47045]_  & \new_[47038]_ ;
  assign \new_[47050]_  = ~A167 & ~A168;
  assign \new_[47051]_  = A169 & \new_[47050]_ ;
  assign \new_[47055]_  = A200 & ~A199;
  assign \new_[47056]_  = A166 & \new_[47055]_ ;
  assign \new_[47057]_  = \new_[47056]_  & \new_[47051]_ ;
  assign \new_[47061]_  = A265 & A233;
  assign \new_[47062]_  = A232 & \new_[47061]_ ;
  assign \new_[47065]_  = ~A299 & A266;
  assign \new_[47068]_  = ~A302 & ~A301;
  assign \new_[47069]_  = \new_[47068]_  & \new_[47065]_ ;
  assign \new_[47070]_  = \new_[47069]_  & \new_[47062]_ ;
  assign \new_[47074]_  = ~A167 & ~A168;
  assign \new_[47075]_  = A169 & \new_[47074]_ ;
  assign \new_[47079]_  = A200 & ~A199;
  assign \new_[47080]_  = A166 & \new_[47079]_ ;
  assign \new_[47081]_  = \new_[47080]_  & \new_[47075]_ ;
  assign \new_[47085]_  = ~A265 & A233;
  assign \new_[47086]_  = A232 & \new_[47085]_ ;
  assign \new_[47089]_  = ~A299 & ~A266;
  assign \new_[47092]_  = ~A302 & ~A301;
  assign \new_[47093]_  = \new_[47092]_  & \new_[47089]_ ;
  assign \new_[47094]_  = \new_[47093]_  & \new_[47086]_ ;
  assign \new_[47098]_  = ~A167 & ~A168;
  assign \new_[47099]_  = A169 & \new_[47098]_ ;
  assign \new_[47103]_  = A200 & ~A199;
  assign \new_[47104]_  = A166 & \new_[47103]_ ;
  assign \new_[47105]_  = \new_[47104]_  & \new_[47099]_ ;
  assign \new_[47109]_  = ~A236 & ~A235;
  assign \new_[47110]_  = ~A233 & \new_[47109]_ ;
  assign \new_[47113]_  = A266 & A265;
  assign \new_[47116]_  = ~A300 & A298;
  assign \new_[47117]_  = \new_[47116]_  & \new_[47113]_ ;
  assign \new_[47118]_  = \new_[47117]_  & \new_[47110]_ ;
  assign \new_[47122]_  = ~A167 & ~A168;
  assign \new_[47123]_  = A169 & \new_[47122]_ ;
  assign \new_[47127]_  = A200 & ~A199;
  assign \new_[47128]_  = A166 & \new_[47127]_ ;
  assign \new_[47129]_  = \new_[47128]_  & \new_[47123]_ ;
  assign \new_[47133]_  = ~A236 & ~A235;
  assign \new_[47134]_  = ~A233 & \new_[47133]_ ;
  assign \new_[47137]_  = A266 & A265;
  assign \new_[47140]_  = A299 & A298;
  assign \new_[47141]_  = \new_[47140]_  & \new_[47137]_ ;
  assign \new_[47142]_  = \new_[47141]_  & \new_[47134]_ ;
  assign \new_[47146]_  = ~A167 & ~A168;
  assign \new_[47147]_  = A169 & \new_[47146]_ ;
  assign \new_[47151]_  = A200 & ~A199;
  assign \new_[47152]_  = A166 & \new_[47151]_ ;
  assign \new_[47153]_  = \new_[47152]_  & \new_[47147]_ ;
  assign \new_[47157]_  = ~A236 & ~A235;
  assign \new_[47158]_  = ~A233 & \new_[47157]_ ;
  assign \new_[47161]_  = A266 & A265;
  assign \new_[47164]_  = ~A299 & ~A298;
  assign \new_[47165]_  = \new_[47164]_  & \new_[47161]_ ;
  assign \new_[47166]_  = \new_[47165]_  & \new_[47158]_ ;
  assign \new_[47170]_  = ~A167 & ~A168;
  assign \new_[47171]_  = A169 & \new_[47170]_ ;
  assign \new_[47175]_  = A200 & ~A199;
  assign \new_[47176]_  = A166 & \new_[47175]_ ;
  assign \new_[47177]_  = \new_[47176]_  & \new_[47171]_ ;
  assign \new_[47181]_  = ~A236 & ~A235;
  assign \new_[47182]_  = ~A233 & \new_[47181]_ ;
  assign \new_[47185]_  = ~A267 & ~A266;
  assign \new_[47188]_  = ~A300 & A298;
  assign \new_[47189]_  = \new_[47188]_  & \new_[47185]_ ;
  assign \new_[47190]_  = \new_[47189]_  & \new_[47182]_ ;
  assign \new_[47194]_  = ~A167 & ~A168;
  assign \new_[47195]_  = A169 & \new_[47194]_ ;
  assign \new_[47199]_  = A200 & ~A199;
  assign \new_[47200]_  = A166 & \new_[47199]_ ;
  assign \new_[47201]_  = \new_[47200]_  & \new_[47195]_ ;
  assign \new_[47205]_  = ~A236 & ~A235;
  assign \new_[47206]_  = ~A233 & \new_[47205]_ ;
  assign \new_[47209]_  = ~A267 & ~A266;
  assign \new_[47212]_  = A299 & A298;
  assign \new_[47213]_  = \new_[47212]_  & \new_[47209]_ ;
  assign \new_[47214]_  = \new_[47213]_  & \new_[47206]_ ;
  assign \new_[47218]_  = ~A167 & ~A168;
  assign \new_[47219]_  = A169 & \new_[47218]_ ;
  assign \new_[47223]_  = A200 & ~A199;
  assign \new_[47224]_  = A166 & \new_[47223]_ ;
  assign \new_[47225]_  = \new_[47224]_  & \new_[47219]_ ;
  assign \new_[47229]_  = ~A236 & ~A235;
  assign \new_[47230]_  = ~A233 & \new_[47229]_ ;
  assign \new_[47233]_  = ~A267 & ~A266;
  assign \new_[47236]_  = ~A299 & ~A298;
  assign \new_[47237]_  = \new_[47236]_  & \new_[47233]_ ;
  assign \new_[47238]_  = \new_[47237]_  & \new_[47230]_ ;
  assign \new_[47242]_  = ~A167 & ~A168;
  assign \new_[47243]_  = A169 & \new_[47242]_ ;
  assign \new_[47247]_  = A200 & ~A199;
  assign \new_[47248]_  = A166 & \new_[47247]_ ;
  assign \new_[47249]_  = \new_[47248]_  & \new_[47243]_ ;
  assign \new_[47253]_  = ~A236 & ~A235;
  assign \new_[47254]_  = ~A233 & \new_[47253]_ ;
  assign \new_[47257]_  = ~A266 & ~A265;
  assign \new_[47260]_  = ~A300 & A298;
  assign \new_[47261]_  = \new_[47260]_  & \new_[47257]_ ;
  assign \new_[47262]_  = \new_[47261]_  & \new_[47254]_ ;
  assign \new_[47266]_  = ~A167 & ~A168;
  assign \new_[47267]_  = A169 & \new_[47266]_ ;
  assign \new_[47271]_  = A200 & ~A199;
  assign \new_[47272]_  = A166 & \new_[47271]_ ;
  assign \new_[47273]_  = \new_[47272]_  & \new_[47267]_ ;
  assign \new_[47277]_  = ~A236 & ~A235;
  assign \new_[47278]_  = ~A233 & \new_[47277]_ ;
  assign \new_[47281]_  = ~A266 & ~A265;
  assign \new_[47284]_  = A299 & A298;
  assign \new_[47285]_  = \new_[47284]_  & \new_[47281]_ ;
  assign \new_[47286]_  = \new_[47285]_  & \new_[47278]_ ;
  assign \new_[47290]_  = ~A167 & ~A168;
  assign \new_[47291]_  = A169 & \new_[47290]_ ;
  assign \new_[47295]_  = A200 & ~A199;
  assign \new_[47296]_  = A166 & \new_[47295]_ ;
  assign \new_[47297]_  = \new_[47296]_  & \new_[47291]_ ;
  assign \new_[47301]_  = ~A236 & ~A235;
  assign \new_[47302]_  = ~A233 & \new_[47301]_ ;
  assign \new_[47305]_  = ~A266 & ~A265;
  assign \new_[47308]_  = ~A299 & ~A298;
  assign \new_[47309]_  = \new_[47308]_  & \new_[47305]_ ;
  assign \new_[47310]_  = \new_[47309]_  & \new_[47302]_ ;
  assign \new_[47314]_  = ~A167 & ~A168;
  assign \new_[47315]_  = A169 & \new_[47314]_ ;
  assign \new_[47319]_  = A200 & ~A199;
  assign \new_[47320]_  = A166 & \new_[47319]_ ;
  assign \new_[47321]_  = \new_[47320]_  & \new_[47315]_ ;
  assign \new_[47325]_  = A265 & ~A234;
  assign \new_[47326]_  = ~A233 & \new_[47325]_ ;
  assign \new_[47329]_  = A298 & A266;
  assign \new_[47332]_  = ~A302 & ~A301;
  assign \new_[47333]_  = \new_[47332]_  & \new_[47329]_ ;
  assign \new_[47334]_  = \new_[47333]_  & \new_[47326]_ ;
  assign \new_[47338]_  = ~A167 & ~A168;
  assign \new_[47339]_  = A169 & \new_[47338]_ ;
  assign \new_[47343]_  = A200 & ~A199;
  assign \new_[47344]_  = A166 & \new_[47343]_ ;
  assign \new_[47345]_  = \new_[47344]_  & \new_[47339]_ ;
  assign \new_[47349]_  = ~A266 & ~A234;
  assign \new_[47350]_  = ~A233 & \new_[47349]_ ;
  assign \new_[47353]_  = ~A269 & ~A268;
  assign \new_[47356]_  = ~A300 & A298;
  assign \new_[47357]_  = \new_[47356]_  & \new_[47353]_ ;
  assign \new_[47358]_  = \new_[47357]_  & \new_[47350]_ ;
  assign \new_[47362]_  = ~A167 & ~A168;
  assign \new_[47363]_  = A169 & \new_[47362]_ ;
  assign \new_[47367]_  = A200 & ~A199;
  assign \new_[47368]_  = A166 & \new_[47367]_ ;
  assign \new_[47369]_  = \new_[47368]_  & \new_[47363]_ ;
  assign \new_[47373]_  = ~A266 & ~A234;
  assign \new_[47374]_  = ~A233 & \new_[47373]_ ;
  assign \new_[47377]_  = ~A269 & ~A268;
  assign \new_[47380]_  = A299 & A298;
  assign \new_[47381]_  = \new_[47380]_  & \new_[47377]_ ;
  assign \new_[47382]_  = \new_[47381]_  & \new_[47374]_ ;
  assign \new_[47386]_  = ~A167 & ~A168;
  assign \new_[47387]_  = A169 & \new_[47386]_ ;
  assign \new_[47391]_  = A200 & ~A199;
  assign \new_[47392]_  = A166 & \new_[47391]_ ;
  assign \new_[47393]_  = \new_[47392]_  & \new_[47387]_ ;
  assign \new_[47397]_  = ~A266 & ~A234;
  assign \new_[47398]_  = ~A233 & \new_[47397]_ ;
  assign \new_[47401]_  = ~A269 & ~A268;
  assign \new_[47404]_  = ~A299 & ~A298;
  assign \new_[47405]_  = \new_[47404]_  & \new_[47401]_ ;
  assign \new_[47406]_  = \new_[47405]_  & \new_[47398]_ ;
  assign \new_[47410]_  = ~A167 & ~A168;
  assign \new_[47411]_  = A169 & \new_[47410]_ ;
  assign \new_[47415]_  = A200 & ~A199;
  assign \new_[47416]_  = A166 & \new_[47415]_ ;
  assign \new_[47417]_  = \new_[47416]_  & \new_[47411]_ ;
  assign \new_[47421]_  = ~A266 & ~A234;
  assign \new_[47422]_  = ~A233 & \new_[47421]_ ;
  assign \new_[47425]_  = A298 & ~A267;
  assign \new_[47428]_  = ~A302 & ~A301;
  assign \new_[47429]_  = \new_[47428]_  & \new_[47425]_ ;
  assign \new_[47430]_  = \new_[47429]_  & \new_[47422]_ ;
  assign \new_[47434]_  = ~A167 & ~A168;
  assign \new_[47435]_  = A169 & \new_[47434]_ ;
  assign \new_[47439]_  = A200 & ~A199;
  assign \new_[47440]_  = A166 & \new_[47439]_ ;
  assign \new_[47441]_  = \new_[47440]_  & \new_[47435]_ ;
  assign \new_[47445]_  = ~A265 & ~A234;
  assign \new_[47446]_  = ~A233 & \new_[47445]_ ;
  assign \new_[47449]_  = A298 & ~A266;
  assign \new_[47452]_  = ~A302 & ~A301;
  assign \new_[47453]_  = \new_[47452]_  & \new_[47449]_ ;
  assign \new_[47454]_  = \new_[47453]_  & \new_[47446]_ ;
  assign \new_[47458]_  = ~A167 & ~A168;
  assign \new_[47459]_  = A169 & \new_[47458]_ ;
  assign \new_[47463]_  = A200 & ~A199;
  assign \new_[47464]_  = A166 & \new_[47463]_ ;
  assign \new_[47465]_  = \new_[47464]_  & \new_[47459]_ ;
  assign \new_[47469]_  = A265 & ~A233;
  assign \new_[47470]_  = ~A232 & \new_[47469]_ ;
  assign \new_[47473]_  = A298 & A266;
  assign \new_[47476]_  = ~A302 & ~A301;
  assign \new_[47477]_  = \new_[47476]_  & \new_[47473]_ ;
  assign \new_[47478]_  = \new_[47477]_  & \new_[47470]_ ;
  assign \new_[47482]_  = ~A167 & ~A168;
  assign \new_[47483]_  = A169 & \new_[47482]_ ;
  assign \new_[47487]_  = A200 & ~A199;
  assign \new_[47488]_  = A166 & \new_[47487]_ ;
  assign \new_[47489]_  = \new_[47488]_  & \new_[47483]_ ;
  assign \new_[47493]_  = ~A266 & ~A233;
  assign \new_[47494]_  = ~A232 & \new_[47493]_ ;
  assign \new_[47497]_  = ~A269 & ~A268;
  assign \new_[47500]_  = ~A300 & A298;
  assign \new_[47501]_  = \new_[47500]_  & \new_[47497]_ ;
  assign \new_[47502]_  = \new_[47501]_  & \new_[47494]_ ;
  assign \new_[47506]_  = ~A167 & ~A168;
  assign \new_[47507]_  = A169 & \new_[47506]_ ;
  assign \new_[47511]_  = A200 & ~A199;
  assign \new_[47512]_  = A166 & \new_[47511]_ ;
  assign \new_[47513]_  = \new_[47512]_  & \new_[47507]_ ;
  assign \new_[47517]_  = ~A266 & ~A233;
  assign \new_[47518]_  = ~A232 & \new_[47517]_ ;
  assign \new_[47521]_  = ~A269 & ~A268;
  assign \new_[47524]_  = A299 & A298;
  assign \new_[47525]_  = \new_[47524]_  & \new_[47521]_ ;
  assign \new_[47526]_  = \new_[47525]_  & \new_[47518]_ ;
  assign \new_[47530]_  = ~A167 & ~A168;
  assign \new_[47531]_  = A169 & \new_[47530]_ ;
  assign \new_[47535]_  = A200 & ~A199;
  assign \new_[47536]_  = A166 & \new_[47535]_ ;
  assign \new_[47537]_  = \new_[47536]_  & \new_[47531]_ ;
  assign \new_[47541]_  = ~A266 & ~A233;
  assign \new_[47542]_  = ~A232 & \new_[47541]_ ;
  assign \new_[47545]_  = ~A269 & ~A268;
  assign \new_[47548]_  = ~A299 & ~A298;
  assign \new_[47549]_  = \new_[47548]_  & \new_[47545]_ ;
  assign \new_[47550]_  = \new_[47549]_  & \new_[47542]_ ;
  assign \new_[47554]_  = ~A167 & ~A168;
  assign \new_[47555]_  = A169 & \new_[47554]_ ;
  assign \new_[47559]_  = A200 & ~A199;
  assign \new_[47560]_  = A166 & \new_[47559]_ ;
  assign \new_[47561]_  = \new_[47560]_  & \new_[47555]_ ;
  assign \new_[47565]_  = ~A266 & ~A233;
  assign \new_[47566]_  = ~A232 & \new_[47565]_ ;
  assign \new_[47569]_  = A298 & ~A267;
  assign \new_[47572]_  = ~A302 & ~A301;
  assign \new_[47573]_  = \new_[47572]_  & \new_[47569]_ ;
  assign \new_[47574]_  = \new_[47573]_  & \new_[47566]_ ;
  assign \new_[47578]_  = ~A167 & ~A168;
  assign \new_[47579]_  = A169 & \new_[47578]_ ;
  assign \new_[47583]_  = A200 & ~A199;
  assign \new_[47584]_  = A166 & \new_[47583]_ ;
  assign \new_[47585]_  = \new_[47584]_  & \new_[47579]_ ;
  assign \new_[47589]_  = ~A265 & ~A233;
  assign \new_[47590]_  = ~A232 & \new_[47589]_ ;
  assign \new_[47593]_  = A298 & ~A266;
  assign \new_[47596]_  = ~A302 & ~A301;
  assign \new_[47597]_  = \new_[47596]_  & \new_[47593]_ ;
  assign \new_[47598]_  = \new_[47597]_  & \new_[47590]_ ;
  assign \new_[47602]_  = ~A168 & A169;
  assign \new_[47603]_  = A170 & \new_[47602]_ ;
  assign \new_[47607]_  = A201 & ~A200;
  assign \new_[47608]_  = A199 & \new_[47607]_ ;
  assign \new_[47609]_  = \new_[47608]_  & \new_[47603]_ ;
  assign \new_[47613]_  = A233 & A232;
  assign \new_[47614]_  = A202 & \new_[47613]_ ;
  assign \new_[47617]_  = ~A267 & A265;
  assign \new_[47620]_  = ~A300 & ~A299;
  assign \new_[47621]_  = \new_[47620]_  & \new_[47617]_ ;
  assign \new_[47622]_  = \new_[47621]_  & \new_[47614]_ ;
  assign \new_[47626]_  = ~A168 & A169;
  assign \new_[47627]_  = A170 & \new_[47626]_ ;
  assign \new_[47631]_  = A201 & ~A200;
  assign \new_[47632]_  = A199 & \new_[47631]_ ;
  assign \new_[47633]_  = \new_[47632]_  & \new_[47627]_ ;
  assign \new_[47637]_  = A233 & A232;
  assign \new_[47638]_  = A202 & \new_[47637]_ ;
  assign \new_[47641]_  = ~A267 & A265;
  assign \new_[47644]_  = A299 & A298;
  assign \new_[47645]_  = \new_[47644]_  & \new_[47641]_ ;
  assign \new_[47646]_  = \new_[47645]_  & \new_[47638]_ ;
  assign \new_[47650]_  = ~A168 & A169;
  assign \new_[47651]_  = A170 & \new_[47650]_ ;
  assign \new_[47655]_  = A201 & ~A200;
  assign \new_[47656]_  = A199 & \new_[47655]_ ;
  assign \new_[47657]_  = \new_[47656]_  & \new_[47651]_ ;
  assign \new_[47661]_  = A233 & A232;
  assign \new_[47662]_  = A202 & \new_[47661]_ ;
  assign \new_[47665]_  = ~A267 & A265;
  assign \new_[47668]_  = ~A299 & ~A298;
  assign \new_[47669]_  = \new_[47668]_  & \new_[47665]_ ;
  assign \new_[47670]_  = \new_[47669]_  & \new_[47662]_ ;
  assign \new_[47674]_  = ~A168 & A169;
  assign \new_[47675]_  = A170 & \new_[47674]_ ;
  assign \new_[47679]_  = A201 & ~A200;
  assign \new_[47680]_  = A199 & \new_[47679]_ ;
  assign \new_[47681]_  = \new_[47680]_  & \new_[47675]_ ;
  assign \new_[47685]_  = A233 & A232;
  assign \new_[47686]_  = A202 & \new_[47685]_ ;
  assign \new_[47689]_  = A266 & A265;
  assign \new_[47692]_  = ~A300 & ~A299;
  assign \new_[47693]_  = \new_[47692]_  & \new_[47689]_ ;
  assign \new_[47694]_  = \new_[47693]_  & \new_[47686]_ ;
  assign \new_[47698]_  = ~A168 & A169;
  assign \new_[47699]_  = A170 & \new_[47698]_ ;
  assign \new_[47703]_  = A201 & ~A200;
  assign \new_[47704]_  = A199 & \new_[47703]_ ;
  assign \new_[47705]_  = \new_[47704]_  & \new_[47699]_ ;
  assign \new_[47709]_  = A233 & A232;
  assign \new_[47710]_  = A202 & \new_[47709]_ ;
  assign \new_[47713]_  = A266 & A265;
  assign \new_[47716]_  = A299 & A298;
  assign \new_[47717]_  = \new_[47716]_  & \new_[47713]_ ;
  assign \new_[47718]_  = \new_[47717]_  & \new_[47710]_ ;
  assign \new_[47722]_  = ~A168 & A169;
  assign \new_[47723]_  = A170 & \new_[47722]_ ;
  assign \new_[47727]_  = A201 & ~A200;
  assign \new_[47728]_  = A199 & \new_[47727]_ ;
  assign \new_[47729]_  = \new_[47728]_  & \new_[47723]_ ;
  assign \new_[47733]_  = A233 & A232;
  assign \new_[47734]_  = A202 & \new_[47733]_ ;
  assign \new_[47737]_  = A266 & A265;
  assign \new_[47740]_  = ~A299 & ~A298;
  assign \new_[47741]_  = \new_[47740]_  & \new_[47737]_ ;
  assign \new_[47742]_  = \new_[47741]_  & \new_[47734]_ ;
  assign \new_[47746]_  = ~A168 & A169;
  assign \new_[47747]_  = A170 & \new_[47746]_ ;
  assign \new_[47751]_  = A201 & ~A200;
  assign \new_[47752]_  = A199 & \new_[47751]_ ;
  assign \new_[47753]_  = \new_[47752]_  & \new_[47747]_ ;
  assign \new_[47757]_  = A233 & A232;
  assign \new_[47758]_  = A202 & \new_[47757]_ ;
  assign \new_[47761]_  = ~A266 & ~A265;
  assign \new_[47764]_  = ~A300 & ~A299;
  assign \new_[47765]_  = \new_[47764]_  & \new_[47761]_ ;
  assign \new_[47766]_  = \new_[47765]_  & \new_[47758]_ ;
  assign \new_[47770]_  = ~A168 & A169;
  assign \new_[47771]_  = A170 & \new_[47770]_ ;
  assign \new_[47775]_  = A201 & ~A200;
  assign \new_[47776]_  = A199 & \new_[47775]_ ;
  assign \new_[47777]_  = \new_[47776]_  & \new_[47771]_ ;
  assign \new_[47781]_  = A233 & A232;
  assign \new_[47782]_  = A202 & \new_[47781]_ ;
  assign \new_[47785]_  = ~A266 & ~A265;
  assign \new_[47788]_  = A299 & A298;
  assign \new_[47789]_  = \new_[47788]_  & \new_[47785]_ ;
  assign \new_[47790]_  = \new_[47789]_  & \new_[47782]_ ;
  assign \new_[47794]_  = ~A168 & A169;
  assign \new_[47795]_  = A170 & \new_[47794]_ ;
  assign \new_[47799]_  = A201 & ~A200;
  assign \new_[47800]_  = A199 & \new_[47799]_ ;
  assign \new_[47801]_  = \new_[47800]_  & \new_[47795]_ ;
  assign \new_[47805]_  = A233 & A232;
  assign \new_[47806]_  = A202 & \new_[47805]_ ;
  assign \new_[47809]_  = ~A266 & ~A265;
  assign \new_[47812]_  = ~A299 & ~A298;
  assign \new_[47813]_  = \new_[47812]_  & \new_[47809]_ ;
  assign \new_[47814]_  = \new_[47813]_  & \new_[47806]_ ;
  assign \new_[47818]_  = ~A168 & A169;
  assign \new_[47819]_  = A170 & \new_[47818]_ ;
  assign \new_[47823]_  = A201 & ~A200;
  assign \new_[47824]_  = A199 & \new_[47823]_ ;
  assign \new_[47825]_  = \new_[47824]_  & \new_[47819]_ ;
  assign \new_[47829]_  = ~A234 & ~A233;
  assign \new_[47830]_  = A202 & \new_[47829]_ ;
  assign \new_[47833]_  = A266 & A265;
  assign \new_[47836]_  = ~A300 & A298;
  assign \new_[47837]_  = \new_[47836]_  & \new_[47833]_ ;
  assign \new_[47838]_  = \new_[47837]_  & \new_[47830]_ ;
  assign \new_[47842]_  = ~A168 & A169;
  assign \new_[47843]_  = A170 & \new_[47842]_ ;
  assign \new_[47847]_  = A201 & ~A200;
  assign \new_[47848]_  = A199 & \new_[47847]_ ;
  assign \new_[47849]_  = \new_[47848]_  & \new_[47843]_ ;
  assign \new_[47853]_  = ~A234 & ~A233;
  assign \new_[47854]_  = A202 & \new_[47853]_ ;
  assign \new_[47857]_  = A266 & A265;
  assign \new_[47860]_  = A299 & A298;
  assign \new_[47861]_  = \new_[47860]_  & \new_[47857]_ ;
  assign \new_[47862]_  = \new_[47861]_  & \new_[47854]_ ;
  assign \new_[47866]_  = ~A168 & A169;
  assign \new_[47867]_  = A170 & \new_[47866]_ ;
  assign \new_[47871]_  = A201 & ~A200;
  assign \new_[47872]_  = A199 & \new_[47871]_ ;
  assign \new_[47873]_  = \new_[47872]_  & \new_[47867]_ ;
  assign \new_[47877]_  = ~A234 & ~A233;
  assign \new_[47878]_  = A202 & \new_[47877]_ ;
  assign \new_[47881]_  = A266 & A265;
  assign \new_[47884]_  = ~A299 & ~A298;
  assign \new_[47885]_  = \new_[47884]_  & \new_[47881]_ ;
  assign \new_[47886]_  = \new_[47885]_  & \new_[47878]_ ;
  assign \new_[47890]_  = ~A168 & A169;
  assign \new_[47891]_  = A170 & \new_[47890]_ ;
  assign \new_[47895]_  = A201 & ~A200;
  assign \new_[47896]_  = A199 & \new_[47895]_ ;
  assign \new_[47897]_  = \new_[47896]_  & \new_[47891]_ ;
  assign \new_[47901]_  = ~A234 & ~A233;
  assign \new_[47902]_  = A202 & \new_[47901]_ ;
  assign \new_[47905]_  = ~A267 & ~A266;
  assign \new_[47908]_  = ~A300 & A298;
  assign \new_[47909]_  = \new_[47908]_  & \new_[47905]_ ;
  assign \new_[47910]_  = \new_[47909]_  & \new_[47902]_ ;
  assign \new_[47914]_  = ~A168 & A169;
  assign \new_[47915]_  = A170 & \new_[47914]_ ;
  assign \new_[47919]_  = A201 & ~A200;
  assign \new_[47920]_  = A199 & \new_[47919]_ ;
  assign \new_[47921]_  = \new_[47920]_  & \new_[47915]_ ;
  assign \new_[47925]_  = ~A234 & ~A233;
  assign \new_[47926]_  = A202 & \new_[47925]_ ;
  assign \new_[47929]_  = ~A267 & ~A266;
  assign \new_[47932]_  = A299 & A298;
  assign \new_[47933]_  = \new_[47932]_  & \new_[47929]_ ;
  assign \new_[47934]_  = \new_[47933]_  & \new_[47926]_ ;
  assign \new_[47938]_  = ~A168 & A169;
  assign \new_[47939]_  = A170 & \new_[47938]_ ;
  assign \new_[47943]_  = A201 & ~A200;
  assign \new_[47944]_  = A199 & \new_[47943]_ ;
  assign \new_[47945]_  = \new_[47944]_  & \new_[47939]_ ;
  assign \new_[47949]_  = ~A234 & ~A233;
  assign \new_[47950]_  = A202 & \new_[47949]_ ;
  assign \new_[47953]_  = ~A267 & ~A266;
  assign \new_[47956]_  = ~A299 & ~A298;
  assign \new_[47957]_  = \new_[47956]_  & \new_[47953]_ ;
  assign \new_[47958]_  = \new_[47957]_  & \new_[47950]_ ;
  assign \new_[47962]_  = ~A168 & A169;
  assign \new_[47963]_  = A170 & \new_[47962]_ ;
  assign \new_[47967]_  = A201 & ~A200;
  assign \new_[47968]_  = A199 & \new_[47967]_ ;
  assign \new_[47969]_  = \new_[47968]_  & \new_[47963]_ ;
  assign \new_[47973]_  = ~A234 & ~A233;
  assign \new_[47974]_  = A202 & \new_[47973]_ ;
  assign \new_[47977]_  = ~A266 & ~A265;
  assign \new_[47980]_  = ~A300 & A298;
  assign \new_[47981]_  = \new_[47980]_  & \new_[47977]_ ;
  assign \new_[47982]_  = \new_[47981]_  & \new_[47974]_ ;
  assign \new_[47986]_  = ~A168 & A169;
  assign \new_[47987]_  = A170 & \new_[47986]_ ;
  assign \new_[47991]_  = A201 & ~A200;
  assign \new_[47992]_  = A199 & \new_[47991]_ ;
  assign \new_[47993]_  = \new_[47992]_  & \new_[47987]_ ;
  assign \new_[47997]_  = ~A234 & ~A233;
  assign \new_[47998]_  = A202 & \new_[47997]_ ;
  assign \new_[48001]_  = ~A266 & ~A265;
  assign \new_[48004]_  = A299 & A298;
  assign \new_[48005]_  = \new_[48004]_  & \new_[48001]_ ;
  assign \new_[48006]_  = \new_[48005]_  & \new_[47998]_ ;
  assign \new_[48010]_  = ~A168 & A169;
  assign \new_[48011]_  = A170 & \new_[48010]_ ;
  assign \new_[48015]_  = A201 & ~A200;
  assign \new_[48016]_  = A199 & \new_[48015]_ ;
  assign \new_[48017]_  = \new_[48016]_  & \new_[48011]_ ;
  assign \new_[48021]_  = ~A234 & ~A233;
  assign \new_[48022]_  = A202 & \new_[48021]_ ;
  assign \new_[48025]_  = ~A266 & ~A265;
  assign \new_[48028]_  = ~A299 & ~A298;
  assign \new_[48029]_  = \new_[48028]_  & \new_[48025]_ ;
  assign \new_[48030]_  = \new_[48029]_  & \new_[48022]_ ;
  assign \new_[48034]_  = ~A168 & A169;
  assign \new_[48035]_  = A170 & \new_[48034]_ ;
  assign \new_[48039]_  = A201 & ~A200;
  assign \new_[48040]_  = A199 & \new_[48039]_ ;
  assign \new_[48041]_  = \new_[48040]_  & \new_[48035]_ ;
  assign \new_[48045]_  = ~A233 & A232;
  assign \new_[48046]_  = A202 & \new_[48045]_ ;
  assign \new_[48049]_  = A235 & A234;
  assign \new_[48052]_  = A299 & ~A298;
  assign \new_[48053]_  = \new_[48052]_  & \new_[48049]_ ;
  assign \new_[48054]_  = \new_[48053]_  & \new_[48046]_ ;
  assign \new_[48058]_  = ~A168 & A169;
  assign \new_[48059]_  = A170 & \new_[48058]_ ;
  assign \new_[48063]_  = A201 & ~A200;
  assign \new_[48064]_  = A199 & \new_[48063]_ ;
  assign \new_[48065]_  = \new_[48064]_  & \new_[48059]_ ;
  assign \new_[48069]_  = ~A233 & A232;
  assign \new_[48070]_  = A202 & \new_[48069]_ ;
  assign \new_[48073]_  = A235 & A234;
  assign \new_[48076]_  = A266 & ~A265;
  assign \new_[48077]_  = \new_[48076]_  & \new_[48073]_ ;
  assign \new_[48078]_  = \new_[48077]_  & \new_[48070]_ ;
  assign \new_[48082]_  = ~A168 & A169;
  assign \new_[48083]_  = A170 & \new_[48082]_ ;
  assign \new_[48087]_  = A201 & ~A200;
  assign \new_[48088]_  = A199 & \new_[48087]_ ;
  assign \new_[48089]_  = \new_[48088]_  & \new_[48083]_ ;
  assign \new_[48093]_  = ~A233 & A232;
  assign \new_[48094]_  = A202 & \new_[48093]_ ;
  assign \new_[48097]_  = A236 & A234;
  assign \new_[48100]_  = A299 & ~A298;
  assign \new_[48101]_  = \new_[48100]_  & \new_[48097]_ ;
  assign \new_[48102]_  = \new_[48101]_  & \new_[48094]_ ;
  assign \new_[48106]_  = ~A168 & A169;
  assign \new_[48107]_  = A170 & \new_[48106]_ ;
  assign \new_[48111]_  = A201 & ~A200;
  assign \new_[48112]_  = A199 & \new_[48111]_ ;
  assign \new_[48113]_  = \new_[48112]_  & \new_[48107]_ ;
  assign \new_[48117]_  = ~A233 & A232;
  assign \new_[48118]_  = A202 & \new_[48117]_ ;
  assign \new_[48121]_  = A236 & A234;
  assign \new_[48124]_  = A266 & ~A265;
  assign \new_[48125]_  = \new_[48124]_  & \new_[48121]_ ;
  assign \new_[48126]_  = \new_[48125]_  & \new_[48118]_ ;
  assign \new_[48130]_  = ~A168 & A169;
  assign \new_[48131]_  = A170 & \new_[48130]_ ;
  assign \new_[48135]_  = A201 & ~A200;
  assign \new_[48136]_  = A199 & \new_[48135]_ ;
  assign \new_[48137]_  = \new_[48136]_  & \new_[48131]_ ;
  assign \new_[48141]_  = ~A233 & ~A232;
  assign \new_[48142]_  = A202 & \new_[48141]_ ;
  assign \new_[48145]_  = A266 & A265;
  assign \new_[48148]_  = ~A300 & A298;
  assign \new_[48149]_  = \new_[48148]_  & \new_[48145]_ ;
  assign \new_[48150]_  = \new_[48149]_  & \new_[48142]_ ;
  assign \new_[48154]_  = ~A168 & A169;
  assign \new_[48155]_  = A170 & \new_[48154]_ ;
  assign \new_[48159]_  = A201 & ~A200;
  assign \new_[48160]_  = A199 & \new_[48159]_ ;
  assign \new_[48161]_  = \new_[48160]_  & \new_[48155]_ ;
  assign \new_[48165]_  = ~A233 & ~A232;
  assign \new_[48166]_  = A202 & \new_[48165]_ ;
  assign \new_[48169]_  = A266 & A265;
  assign \new_[48172]_  = A299 & A298;
  assign \new_[48173]_  = \new_[48172]_  & \new_[48169]_ ;
  assign \new_[48174]_  = \new_[48173]_  & \new_[48166]_ ;
  assign \new_[48178]_  = ~A168 & A169;
  assign \new_[48179]_  = A170 & \new_[48178]_ ;
  assign \new_[48183]_  = A201 & ~A200;
  assign \new_[48184]_  = A199 & \new_[48183]_ ;
  assign \new_[48185]_  = \new_[48184]_  & \new_[48179]_ ;
  assign \new_[48189]_  = ~A233 & ~A232;
  assign \new_[48190]_  = A202 & \new_[48189]_ ;
  assign \new_[48193]_  = A266 & A265;
  assign \new_[48196]_  = ~A299 & ~A298;
  assign \new_[48197]_  = \new_[48196]_  & \new_[48193]_ ;
  assign \new_[48198]_  = \new_[48197]_  & \new_[48190]_ ;
  assign \new_[48202]_  = ~A168 & A169;
  assign \new_[48203]_  = A170 & \new_[48202]_ ;
  assign \new_[48207]_  = A201 & ~A200;
  assign \new_[48208]_  = A199 & \new_[48207]_ ;
  assign \new_[48209]_  = \new_[48208]_  & \new_[48203]_ ;
  assign \new_[48213]_  = ~A233 & ~A232;
  assign \new_[48214]_  = A202 & \new_[48213]_ ;
  assign \new_[48217]_  = ~A267 & ~A266;
  assign \new_[48220]_  = ~A300 & A298;
  assign \new_[48221]_  = \new_[48220]_  & \new_[48217]_ ;
  assign \new_[48222]_  = \new_[48221]_  & \new_[48214]_ ;
  assign \new_[48226]_  = ~A168 & A169;
  assign \new_[48227]_  = A170 & \new_[48226]_ ;
  assign \new_[48231]_  = A201 & ~A200;
  assign \new_[48232]_  = A199 & \new_[48231]_ ;
  assign \new_[48233]_  = \new_[48232]_  & \new_[48227]_ ;
  assign \new_[48237]_  = ~A233 & ~A232;
  assign \new_[48238]_  = A202 & \new_[48237]_ ;
  assign \new_[48241]_  = ~A267 & ~A266;
  assign \new_[48244]_  = A299 & A298;
  assign \new_[48245]_  = \new_[48244]_  & \new_[48241]_ ;
  assign \new_[48246]_  = \new_[48245]_  & \new_[48238]_ ;
  assign \new_[48250]_  = ~A168 & A169;
  assign \new_[48251]_  = A170 & \new_[48250]_ ;
  assign \new_[48255]_  = A201 & ~A200;
  assign \new_[48256]_  = A199 & \new_[48255]_ ;
  assign \new_[48257]_  = \new_[48256]_  & \new_[48251]_ ;
  assign \new_[48261]_  = ~A233 & ~A232;
  assign \new_[48262]_  = A202 & \new_[48261]_ ;
  assign \new_[48265]_  = ~A267 & ~A266;
  assign \new_[48268]_  = ~A299 & ~A298;
  assign \new_[48269]_  = \new_[48268]_  & \new_[48265]_ ;
  assign \new_[48270]_  = \new_[48269]_  & \new_[48262]_ ;
  assign \new_[48274]_  = ~A168 & A169;
  assign \new_[48275]_  = A170 & \new_[48274]_ ;
  assign \new_[48279]_  = A201 & ~A200;
  assign \new_[48280]_  = A199 & \new_[48279]_ ;
  assign \new_[48281]_  = \new_[48280]_  & \new_[48275]_ ;
  assign \new_[48285]_  = ~A233 & ~A232;
  assign \new_[48286]_  = A202 & \new_[48285]_ ;
  assign \new_[48289]_  = ~A266 & ~A265;
  assign \new_[48292]_  = ~A300 & A298;
  assign \new_[48293]_  = \new_[48292]_  & \new_[48289]_ ;
  assign \new_[48294]_  = \new_[48293]_  & \new_[48286]_ ;
  assign \new_[48298]_  = ~A168 & A169;
  assign \new_[48299]_  = A170 & \new_[48298]_ ;
  assign \new_[48303]_  = A201 & ~A200;
  assign \new_[48304]_  = A199 & \new_[48303]_ ;
  assign \new_[48305]_  = \new_[48304]_  & \new_[48299]_ ;
  assign \new_[48309]_  = ~A233 & ~A232;
  assign \new_[48310]_  = A202 & \new_[48309]_ ;
  assign \new_[48313]_  = ~A266 & ~A265;
  assign \new_[48316]_  = A299 & A298;
  assign \new_[48317]_  = \new_[48316]_  & \new_[48313]_ ;
  assign \new_[48318]_  = \new_[48317]_  & \new_[48310]_ ;
  assign \new_[48322]_  = ~A168 & A169;
  assign \new_[48323]_  = A170 & \new_[48322]_ ;
  assign \new_[48327]_  = A201 & ~A200;
  assign \new_[48328]_  = A199 & \new_[48327]_ ;
  assign \new_[48329]_  = \new_[48328]_  & \new_[48323]_ ;
  assign \new_[48333]_  = ~A233 & ~A232;
  assign \new_[48334]_  = A202 & \new_[48333]_ ;
  assign \new_[48337]_  = ~A266 & ~A265;
  assign \new_[48340]_  = ~A299 & ~A298;
  assign \new_[48341]_  = \new_[48340]_  & \new_[48337]_ ;
  assign \new_[48342]_  = \new_[48341]_  & \new_[48334]_ ;
  assign \new_[48346]_  = ~A168 & A169;
  assign \new_[48347]_  = A170 & \new_[48346]_ ;
  assign \new_[48351]_  = A201 & ~A200;
  assign \new_[48352]_  = A199 & \new_[48351]_ ;
  assign \new_[48353]_  = \new_[48352]_  & \new_[48347]_ ;
  assign \new_[48357]_  = A233 & A232;
  assign \new_[48358]_  = A203 & \new_[48357]_ ;
  assign \new_[48361]_  = ~A267 & A265;
  assign \new_[48364]_  = ~A300 & ~A299;
  assign \new_[48365]_  = \new_[48364]_  & \new_[48361]_ ;
  assign \new_[48366]_  = \new_[48365]_  & \new_[48358]_ ;
  assign \new_[48370]_  = ~A168 & A169;
  assign \new_[48371]_  = A170 & \new_[48370]_ ;
  assign \new_[48375]_  = A201 & ~A200;
  assign \new_[48376]_  = A199 & \new_[48375]_ ;
  assign \new_[48377]_  = \new_[48376]_  & \new_[48371]_ ;
  assign \new_[48381]_  = A233 & A232;
  assign \new_[48382]_  = A203 & \new_[48381]_ ;
  assign \new_[48385]_  = ~A267 & A265;
  assign \new_[48388]_  = A299 & A298;
  assign \new_[48389]_  = \new_[48388]_  & \new_[48385]_ ;
  assign \new_[48390]_  = \new_[48389]_  & \new_[48382]_ ;
  assign \new_[48394]_  = ~A168 & A169;
  assign \new_[48395]_  = A170 & \new_[48394]_ ;
  assign \new_[48399]_  = A201 & ~A200;
  assign \new_[48400]_  = A199 & \new_[48399]_ ;
  assign \new_[48401]_  = \new_[48400]_  & \new_[48395]_ ;
  assign \new_[48405]_  = A233 & A232;
  assign \new_[48406]_  = A203 & \new_[48405]_ ;
  assign \new_[48409]_  = ~A267 & A265;
  assign \new_[48412]_  = ~A299 & ~A298;
  assign \new_[48413]_  = \new_[48412]_  & \new_[48409]_ ;
  assign \new_[48414]_  = \new_[48413]_  & \new_[48406]_ ;
  assign \new_[48418]_  = ~A168 & A169;
  assign \new_[48419]_  = A170 & \new_[48418]_ ;
  assign \new_[48423]_  = A201 & ~A200;
  assign \new_[48424]_  = A199 & \new_[48423]_ ;
  assign \new_[48425]_  = \new_[48424]_  & \new_[48419]_ ;
  assign \new_[48429]_  = A233 & A232;
  assign \new_[48430]_  = A203 & \new_[48429]_ ;
  assign \new_[48433]_  = A266 & A265;
  assign \new_[48436]_  = ~A300 & ~A299;
  assign \new_[48437]_  = \new_[48436]_  & \new_[48433]_ ;
  assign \new_[48438]_  = \new_[48437]_  & \new_[48430]_ ;
  assign \new_[48442]_  = ~A168 & A169;
  assign \new_[48443]_  = A170 & \new_[48442]_ ;
  assign \new_[48447]_  = A201 & ~A200;
  assign \new_[48448]_  = A199 & \new_[48447]_ ;
  assign \new_[48449]_  = \new_[48448]_  & \new_[48443]_ ;
  assign \new_[48453]_  = A233 & A232;
  assign \new_[48454]_  = A203 & \new_[48453]_ ;
  assign \new_[48457]_  = A266 & A265;
  assign \new_[48460]_  = A299 & A298;
  assign \new_[48461]_  = \new_[48460]_  & \new_[48457]_ ;
  assign \new_[48462]_  = \new_[48461]_  & \new_[48454]_ ;
  assign \new_[48466]_  = ~A168 & A169;
  assign \new_[48467]_  = A170 & \new_[48466]_ ;
  assign \new_[48471]_  = A201 & ~A200;
  assign \new_[48472]_  = A199 & \new_[48471]_ ;
  assign \new_[48473]_  = \new_[48472]_  & \new_[48467]_ ;
  assign \new_[48477]_  = A233 & A232;
  assign \new_[48478]_  = A203 & \new_[48477]_ ;
  assign \new_[48481]_  = A266 & A265;
  assign \new_[48484]_  = ~A299 & ~A298;
  assign \new_[48485]_  = \new_[48484]_  & \new_[48481]_ ;
  assign \new_[48486]_  = \new_[48485]_  & \new_[48478]_ ;
  assign \new_[48490]_  = ~A168 & A169;
  assign \new_[48491]_  = A170 & \new_[48490]_ ;
  assign \new_[48495]_  = A201 & ~A200;
  assign \new_[48496]_  = A199 & \new_[48495]_ ;
  assign \new_[48497]_  = \new_[48496]_  & \new_[48491]_ ;
  assign \new_[48501]_  = A233 & A232;
  assign \new_[48502]_  = A203 & \new_[48501]_ ;
  assign \new_[48505]_  = ~A266 & ~A265;
  assign \new_[48508]_  = ~A300 & ~A299;
  assign \new_[48509]_  = \new_[48508]_  & \new_[48505]_ ;
  assign \new_[48510]_  = \new_[48509]_  & \new_[48502]_ ;
  assign \new_[48514]_  = ~A168 & A169;
  assign \new_[48515]_  = A170 & \new_[48514]_ ;
  assign \new_[48519]_  = A201 & ~A200;
  assign \new_[48520]_  = A199 & \new_[48519]_ ;
  assign \new_[48521]_  = \new_[48520]_  & \new_[48515]_ ;
  assign \new_[48525]_  = A233 & A232;
  assign \new_[48526]_  = A203 & \new_[48525]_ ;
  assign \new_[48529]_  = ~A266 & ~A265;
  assign \new_[48532]_  = A299 & A298;
  assign \new_[48533]_  = \new_[48532]_  & \new_[48529]_ ;
  assign \new_[48534]_  = \new_[48533]_  & \new_[48526]_ ;
  assign \new_[48538]_  = ~A168 & A169;
  assign \new_[48539]_  = A170 & \new_[48538]_ ;
  assign \new_[48543]_  = A201 & ~A200;
  assign \new_[48544]_  = A199 & \new_[48543]_ ;
  assign \new_[48545]_  = \new_[48544]_  & \new_[48539]_ ;
  assign \new_[48549]_  = A233 & A232;
  assign \new_[48550]_  = A203 & \new_[48549]_ ;
  assign \new_[48553]_  = ~A266 & ~A265;
  assign \new_[48556]_  = ~A299 & ~A298;
  assign \new_[48557]_  = \new_[48556]_  & \new_[48553]_ ;
  assign \new_[48558]_  = \new_[48557]_  & \new_[48550]_ ;
  assign \new_[48562]_  = ~A168 & A169;
  assign \new_[48563]_  = A170 & \new_[48562]_ ;
  assign \new_[48567]_  = A201 & ~A200;
  assign \new_[48568]_  = A199 & \new_[48567]_ ;
  assign \new_[48569]_  = \new_[48568]_  & \new_[48563]_ ;
  assign \new_[48573]_  = ~A234 & ~A233;
  assign \new_[48574]_  = A203 & \new_[48573]_ ;
  assign \new_[48577]_  = A266 & A265;
  assign \new_[48580]_  = ~A300 & A298;
  assign \new_[48581]_  = \new_[48580]_  & \new_[48577]_ ;
  assign \new_[48582]_  = \new_[48581]_  & \new_[48574]_ ;
  assign \new_[48586]_  = ~A168 & A169;
  assign \new_[48587]_  = A170 & \new_[48586]_ ;
  assign \new_[48591]_  = A201 & ~A200;
  assign \new_[48592]_  = A199 & \new_[48591]_ ;
  assign \new_[48593]_  = \new_[48592]_  & \new_[48587]_ ;
  assign \new_[48597]_  = ~A234 & ~A233;
  assign \new_[48598]_  = A203 & \new_[48597]_ ;
  assign \new_[48601]_  = A266 & A265;
  assign \new_[48604]_  = A299 & A298;
  assign \new_[48605]_  = \new_[48604]_  & \new_[48601]_ ;
  assign \new_[48606]_  = \new_[48605]_  & \new_[48598]_ ;
  assign \new_[48610]_  = ~A168 & A169;
  assign \new_[48611]_  = A170 & \new_[48610]_ ;
  assign \new_[48615]_  = A201 & ~A200;
  assign \new_[48616]_  = A199 & \new_[48615]_ ;
  assign \new_[48617]_  = \new_[48616]_  & \new_[48611]_ ;
  assign \new_[48621]_  = ~A234 & ~A233;
  assign \new_[48622]_  = A203 & \new_[48621]_ ;
  assign \new_[48625]_  = A266 & A265;
  assign \new_[48628]_  = ~A299 & ~A298;
  assign \new_[48629]_  = \new_[48628]_  & \new_[48625]_ ;
  assign \new_[48630]_  = \new_[48629]_  & \new_[48622]_ ;
  assign \new_[48634]_  = ~A168 & A169;
  assign \new_[48635]_  = A170 & \new_[48634]_ ;
  assign \new_[48639]_  = A201 & ~A200;
  assign \new_[48640]_  = A199 & \new_[48639]_ ;
  assign \new_[48641]_  = \new_[48640]_  & \new_[48635]_ ;
  assign \new_[48645]_  = ~A234 & ~A233;
  assign \new_[48646]_  = A203 & \new_[48645]_ ;
  assign \new_[48649]_  = ~A267 & ~A266;
  assign \new_[48652]_  = ~A300 & A298;
  assign \new_[48653]_  = \new_[48652]_  & \new_[48649]_ ;
  assign \new_[48654]_  = \new_[48653]_  & \new_[48646]_ ;
  assign \new_[48658]_  = ~A168 & A169;
  assign \new_[48659]_  = A170 & \new_[48658]_ ;
  assign \new_[48663]_  = A201 & ~A200;
  assign \new_[48664]_  = A199 & \new_[48663]_ ;
  assign \new_[48665]_  = \new_[48664]_  & \new_[48659]_ ;
  assign \new_[48669]_  = ~A234 & ~A233;
  assign \new_[48670]_  = A203 & \new_[48669]_ ;
  assign \new_[48673]_  = ~A267 & ~A266;
  assign \new_[48676]_  = A299 & A298;
  assign \new_[48677]_  = \new_[48676]_  & \new_[48673]_ ;
  assign \new_[48678]_  = \new_[48677]_  & \new_[48670]_ ;
  assign \new_[48682]_  = ~A168 & A169;
  assign \new_[48683]_  = A170 & \new_[48682]_ ;
  assign \new_[48687]_  = A201 & ~A200;
  assign \new_[48688]_  = A199 & \new_[48687]_ ;
  assign \new_[48689]_  = \new_[48688]_  & \new_[48683]_ ;
  assign \new_[48693]_  = ~A234 & ~A233;
  assign \new_[48694]_  = A203 & \new_[48693]_ ;
  assign \new_[48697]_  = ~A267 & ~A266;
  assign \new_[48700]_  = ~A299 & ~A298;
  assign \new_[48701]_  = \new_[48700]_  & \new_[48697]_ ;
  assign \new_[48702]_  = \new_[48701]_  & \new_[48694]_ ;
  assign \new_[48706]_  = ~A168 & A169;
  assign \new_[48707]_  = A170 & \new_[48706]_ ;
  assign \new_[48711]_  = A201 & ~A200;
  assign \new_[48712]_  = A199 & \new_[48711]_ ;
  assign \new_[48713]_  = \new_[48712]_  & \new_[48707]_ ;
  assign \new_[48717]_  = ~A234 & ~A233;
  assign \new_[48718]_  = A203 & \new_[48717]_ ;
  assign \new_[48721]_  = ~A266 & ~A265;
  assign \new_[48724]_  = ~A300 & A298;
  assign \new_[48725]_  = \new_[48724]_  & \new_[48721]_ ;
  assign \new_[48726]_  = \new_[48725]_  & \new_[48718]_ ;
  assign \new_[48730]_  = ~A168 & A169;
  assign \new_[48731]_  = A170 & \new_[48730]_ ;
  assign \new_[48735]_  = A201 & ~A200;
  assign \new_[48736]_  = A199 & \new_[48735]_ ;
  assign \new_[48737]_  = \new_[48736]_  & \new_[48731]_ ;
  assign \new_[48741]_  = ~A234 & ~A233;
  assign \new_[48742]_  = A203 & \new_[48741]_ ;
  assign \new_[48745]_  = ~A266 & ~A265;
  assign \new_[48748]_  = A299 & A298;
  assign \new_[48749]_  = \new_[48748]_  & \new_[48745]_ ;
  assign \new_[48750]_  = \new_[48749]_  & \new_[48742]_ ;
  assign \new_[48754]_  = ~A168 & A169;
  assign \new_[48755]_  = A170 & \new_[48754]_ ;
  assign \new_[48759]_  = A201 & ~A200;
  assign \new_[48760]_  = A199 & \new_[48759]_ ;
  assign \new_[48761]_  = \new_[48760]_  & \new_[48755]_ ;
  assign \new_[48765]_  = ~A234 & ~A233;
  assign \new_[48766]_  = A203 & \new_[48765]_ ;
  assign \new_[48769]_  = ~A266 & ~A265;
  assign \new_[48772]_  = ~A299 & ~A298;
  assign \new_[48773]_  = \new_[48772]_  & \new_[48769]_ ;
  assign \new_[48774]_  = \new_[48773]_  & \new_[48766]_ ;
  assign \new_[48778]_  = ~A168 & A169;
  assign \new_[48779]_  = A170 & \new_[48778]_ ;
  assign \new_[48783]_  = A201 & ~A200;
  assign \new_[48784]_  = A199 & \new_[48783]_ ;
  assign \new_[48785]_  = \new_[48784]_  & \new_[48779]_ ;
  assign \new_[48789]_  = ~A233 & A232;
  assign \new_[48790]_  = A203 & \new_[48789]_ ;
  assign \new_[48793]_  = A235 & A234;
  assign \new_[48796]_  = A299 & ~A298;
  assign \new_[48797]_  = \new_[48796]_  & \new_[48793]_ ;
  assign \new_[48798]_  = \new_[48797]_  & \new_[48790]_ ;
  assign \new_[48802]_  = ~A168 & A169;
  assign \new_[48803]_  = A170 & \new_[48802]_ ;
  assign \new_[48807]_  = A201 & ~A200;
  assign \new_[48808]_  = A199 & \new_[48807]_ ;
  assign \new_[48809]_  = \new_[48808]_  & \new_[48803]_ ;
  assign \new_[48813]_  = ~A233 & A232;
  assign \new_[48814]_  = A203 & \new_[48813]_ ;
  assign \new_[48817]_  = A235 & A234;
  assign \new_[48820]_  = A266 & ~A265;
  assign \new_[48821]_  = \new_[48820]_  & \new_[48817]_ ;
  assign \new_[48822]_  = \new_[48821]_  & \new_[48814]_ ;
  assign \new_[48826]_  = ~A168 & A169;
  assign \new_[48827]_  = A170 & \new_[48826]_ ;
  assign \new_[48831]_  = A201 & ~A200;
  assign \new_[48832]_  = A199 & \new_[48831]_ ;
  assign \new_[48833]_  = \new_[48832]_  & \new_[48827]_ ;
  assign \new_[48837]_  = ~A233 & A232;
  assign \new_[48838]_  = A203 & \new_[48837]_ ;
  assign \new_[48841]_  = A236 & A234;
  assign \new_[48844]_  = A299 & ~A298;
  assign \new_[48845]_  = \new_[48844]_  & \new_[48841]_ ;
  assign \new_[48846]_  = \new_[48845]_  & \new_[48838]_ ;
  assign \new_[48850]_  = ~A168 & A169;
  assign \new_[48851]_  = A170 & \new_[48850]_ ;
  assign \new_[48855]_  = A201 & ~A200;
  assign \new_[48856]_  = A199 & \new_[48855]_ ;
  assign \new_[48857]_  = \new_[48856]_  & \new_[48851]_ ;
  assign \new_[48861]_  = ~A233 & A232;
  assign \new_[48862]_  = A203 & \new_[48861]_ ;
  assign \new_[48865]_  = A236 & A234;
  assign \new_[48868]_  = A266 & ~A265;
  assign \new_[48869]_  = \new_[48868]_  & \new_[48865]_ ;
  assign \new_[48870]_  = \new_[48869]_  & \new_[48862]_ ;
  assign \new_[48874]_  = ~A168 & A169;
  assign \new_[48875]_  = A170 & \new_[48874]_ ;
  assign \new_[48879]_  = A201 & ~A200;
  assign \new_[48880]_  = A199 & \new_[48879]_ ;
  assign \new_[48881]_  = \new_[48880]_  & \new_[48875]_ ;
  assign \new_[48885]_  = ~A233 & ~A232;
  assign \new_[48886]_  = A203 & \new_[48885]_ ;
  assign \new_[48889]_  = A266 & A265;
  assign \new_[48892]_  = ~A300 & A298;
  assign \new_[48893]_  = \new_[48892]_  & \new_[48889]_ ;
  assign \new_[48894]_  = \new_[48893]_  & \new_[48886]_ ;
  assign \new_[48898]_  = ~A168 & A169;
  assign \new_[48899]_  = A170 & \new_[48898]_ ;
  assign \new_[48903]_  = A201 & ~A200;
  assign \new_[48904]_  = A199 & \new_[48903]_ ;
  assign \new_[48905]_  = \new_[48904]_  & \new_[48899]_ ;
  assign \new_[48909]_  = ~A233 & ~A232;
  assign \new_[48910]_  = A203 & \new_[48909]_ ;
  assign \new_[48913]_  = A266 & A265;
  assign \new_[48916]_  = A299 & A298;
  assign \new_[48917]_  = \new_[48916]_  & \new_[48913]_ ;
  assign \new_[48918]_  = \new_[48917]_  & \new_[48910]_ ;
  assign \new_[48922]_  = ~A168 & A169;
  assign \new_[48923]_  = A170 & \new_[48922]_ ;
  assign \new_[48927]_  = A201 & ~A200;
  assign \new_[48928]_  = A199 & \new_[48927]_ ;
  assign \new_[48929]_  = \new_[48928]_  & \new_[48923]_ ;
  assign \new_[48933]_  = ~A233 & ~A232;
  assign \new_[48934]_  = A203 & \new_[48933]_ ;
  assign \new_[48937]_  = A266 & A265;
  assign \new_[48940]_  = ~A299 & ~A298;
  assign \new_[48941]_  = \new_[48940]_  & \new_[48937]_ ;
  assign \new_[48942]_  = \new_[48941]_  & \new_[48934]_ ;
  assign \new_[48946]_  = ~A168 & A169;
  assign \new_[48947]_  = A170 & \new_[48946]_ ;
  assign \new_[48951]_  = A201 & ~A200;
  assign \new_[48952]_  = A199 & \new_[48951]_ ;
  assign \new_[48953]_  = \new_[48952]_  & \new_[48947]_ ;
  assign \new_[48957]_  = ~A233 & ~A232;
  assign \new_[48958]_  = A203 & \new_[48957]_ ;
  assign \new_[48961]_  = ~A267 & ~A266;
  assign \new_[48964]_  = ~A300 & A298;
  assign \new_[48965]_  = \new_[48964]_  & \new_[48961]_ ;
  assign \new_[48966]_  = \new_[48965]_  & \new_[48958]_ ;
  assign \new_[48970]_  = ~A168 & A169;
  assign \new_[48971]_  = A170 & \new_[48970]_ ;
  assign \new_[48975]_  = A201 & ~A200;
  assign \new_[48976]_  = A199 & \new_[48975]_ ;
  assign \new_[48977]_  = \new_[48976]_  & \new_[48971]_ ;
  assign \new_[48981]_  = ~A233 & ~A232;
  assign \new_[48982]_  = A203 & \new_[48981]_ ;
  assign \new_[48985]_  = ~A267 & ~A266;
  assign \new_[48988]_  = A299 & A298;
  assign \new_[48989]_  = \new_[48988]_  & \new_[48985]_ ;
  assign \new_[48990]_  = \new_[48989]_  & \new_[48982]_ ;
  assign \new_[48994]_  = ~A168 & A169;
  assign \new_[48995]_  = A170 & \new_[48994]_ ;
  assign \new_[48999]_  = A201 & ~A200;
  assign \new_[49000]_  = A199 & \new_[48999]_ ;
  assign \new_[49001]_  = \new_[49000]_  & \new_[48995]_ ;
  assign \new_[49005]_  = ~A233 & ~A232;
  assign \new_[49006]_  = A203 & \new_[49005]_ ;
  assign \new_[49009]_  = ~A267 & ~A266;
  assign \new_[49012]_  = ~A299 & ~A298;
  assign \new_[49013]_  = \new_[49012]_  & \new_[49009]_ ;
  assign \new_[49014]_  = \new_[49013]_  & \new_[49006]_ ;
  assign \new_[49018]_  = ~A168 & A169;
  assign \new_[49019]_  = A170 & \new_[49018]_ ;
  assign \new_[49023]_  = A201 & ~A200;
  assign \new_[49024]_  = A199 & \new_[49023]_ ;
  assign \new_[49025]_  = \new_[49024]_  & \new_[49019]_ ;
  assign \new_[49029]_  = ~A233 & ~A232;
  assign \new_[49030]_  = A203 & \new_[49029]_ ;
  assign \new_[49033]_  = ~A266 & ~A265;
  assign \new_[49036]_  = ~A300 & A298;
  assign \new_[49037]_  = \new_[49036]_  & \new_[49033]_ ;
  assign \new_[49038]_  = \new_[49037]_  & \new_[49030]_ ;
  assign \new_[49042]_  = ~A168 & A169;
  assign \new_[49043]_  = A170 & \new_[49042]_ ;
  assign \new_[49047]_  = A201 & ~A200;
  assign \new_[49048]_  = A199 & \new_[49047]_ ;
  assign \new_[49049]_  = \new_[49048]_  & \new_[49043]_ ;
  assign \new_[49053]_  = ~A233 & ~A232;
  assign \new_[49054]_  = A203 & \new_[49053]_ ;
  assign \new_[49057]_  = ~A266 & ~A265;
  assign \new_[49060]_  = A299 & A298;
  assign \new_[49061]_  = \new_[49060]_  & \new_[49057]_ ;
  assign \new_[49062]_  = \new_[49061]_  & \new_[49054]_ ;
  assign \new_[49066]_  = ~A168 & A169;
  assign \new_[49067]_  = A170 & \new_[49066]_ ;
  assign \new_[49071]_  = A201 & ~A200;
  assign \new_[49072]_  = A199 & \new_[49071]_ ;
  assign \new_[49073]_  = \new_[49072]_  & \new_[49067]_ ;
  assign \new_[49077]_  = ~A233 & ~A232;
  assign \new_[49078]_  = A203 & \new_[49077]_ ;
  assign \new_[49081]_  = ~A266 & ~A265;
  assign \new_[49084]_  = ~A299 & ~A298;
  assign \new_[49085]_  = \new_[49084]_  & \new_[49081]_ ;
  assign \new_[49086]_  = \new_[49085]_  & \new_[49078]_ ;
  assign \new_[49090]_  = A167 & A169;
  assign \new_[49091]_  = ~A170 & \new_[49090]_ ;
  assign \new_[49095]_  = A200 & A199;
  assign \new_[49096]_  = A166 & \new_[49095]_ ;
  assign \new_[49097]_  = \new_[49096]_  & \new_[49091]_ ;
  assign \new_[49101]_  = A265 & A233;
  assign \new_[49102]_  = A232 & \new_[49101]_ ;
  assign \new_[49105]_  = ~A269 & ~A268;
  assign \new_[49108]_  = ~A300 & ~A299;
  assign \new_[49109]_  = \new_[49108]_  & \new_[49105]_ ;
  assign \new_[49110]_  = \new_[49109]_  & \new_[49102]_ ;
  assign \new_[49114]_  = A167 & A169;
  assign \new_[49115]_  = ~A170 & \new_[49114]_ ;
  assign \new_[49119]_  = A200 & A199;
  assign \new_[49120]_  = A166 & \new_[49119]_ ;
  assign \new_[49121]_  = \new_[49120]_  & \new_[49115]_ ;
  assign \new_[49125]_  = A265 & A233;
  assign \new_[49126]_  = A232 & \new_[49125]_ ;
  assign \new_[49129]_  = ~A269 & ~A268;
  assign \new_[49132]_  = A299 & A298;
  assign \new_[49133]_  = \new_[49132]_  & \new_[49129]_ ;
  assign \new_[49134]_  = \new_[49133]_  & \new_[49126]_ ;
  assign \new_[49138]_  = A167 & A169;
  assign \new_[49139]_  = ~A170 & \new_[49138]_ ;
  assign \new_[49143]_  = A200 & A199;
  assign \new_[49144]_  = A166 & \new_[49143]_ ;
  assign \new_[49145]_  = \new_[49144]_  & \new_[49139]_ ;
  assign \new_[49149]_  = A265 & A233;
  assign \new_[49150]_  = A232 & \new_[49149]_ ;
  assign \new_[49153]_  = ~A269 & ~A268;
  assign \new_[49156]_  = ~A299 & ~A298;
  assign \new_[49157]_  = \new_[49156]_  & \new_[49153]_ ;
  assign \new_[49158]_  = \new_[49157]_  & \new_[49150]_ ;
  assign \new_[49162]_  = A167 & A169;
  assign \new_[49163]_  = ~A170 & \new_[49162]_ ;
  assign \new_[49167]_  = A200 & A199;
  assign \new_[49168]_  = A166 & \new_[49167]_ ;
  assign \new_[49169]_  = \new_[49168]_  & \new_[49163]_ ;
  assign \new_[49173]_  = A265 & A233;
  assign \new_[49174]_  = A232 & \new_[49173]_ ;
  assign \new_[49177]_  = ~A299 & ~A267;
  assign \new_[49180]_  = ~A302 & ~A301;
  assign \new_[49181]_  = \new_[49180]_  & \new_[49177]_ ;
  assign \new_[49182]_  = \new_[49181]_  & \new_[49174]_ ;
  assign \new_[49186]_  = A167 & A169;
  assign \new_[49187]_  = ~A170 & \new_[49186]_ ;
  assign \new_[49191]_  = A200 & A199;
  assign \new_[49192]_  = A166 & \new_[49191]_ ;
  assign \new_[49193]_  = \new_[49192]_  & \new_[49187]_ ;
  assign \new_[49197]_  = A265 & A233;
  assign \new_[49198]_  = A232 & \new_[49197]_ ;
  assign \new_[49201]_  = ~A299 & A266;
  assign \new_[49204]_  = ~A302 & ~A301;
  assign \new_[49205]_  = \new_[49204]_  & \new_[49201]_ ;
  assign \new_[49206]_  = \new_[49205]_  & \new_[49198]_ ;
  assign \new_[49210]_  = A167 & A169;
  assign \new_[49211]_  = ~A170 & \new_[49210]_ ;
  assign \new_[49215]_  = A200 & A199;
  assign \new_[49216]_  = A166 & \new_[49215]_ ;
  assign \new_[49217]_  = \new_[49216]_  & \new_[49211]_ ;
  assign \new_[49221]_  = ~A265 & A233;
  assign \new_[49222]_  = A232 & \new_[49221]_ ;
  assign \new_[49225]_  = ~A299 & ~A266;
  assign \new_[49228]_  = ~A302 & ~A301;
  assign \new_[49229]_  = \new_[49228]_  & \new_[49225]_ ;
  assign \new_[49230]_  = \new_[49229]_  & \new_[49222]_ ;
  assign \new_[49234]_  = A167 & A169;
  assign \new_[49235]_  = ~A170 & \new_[49234]_ ;
  assign \new_[49239]_  = A200 & A199;
  assign \new_[49240]_  = A166 & \new_[49239]_ ;
  assign \new_[49241]_  = \new_[49240]_  & \new_[49235]_ ;
  assign \new_[49245]_  = ~A236 & ~A235;
  assign \new_[49246]_  = ~A233 & \new_[49245]_ ;
  assign \new_[49249]_  = A266 & A265;
  assign \new_[49252]_  = ~A300 & A298;
  assign \new_[49253]_  = \new_[49252]_  & \new_[49249]_ ;
  assign \new_[49254]_  = \new_[49253]_  & \new_[49246]_ ;
  assign \new_[49258]_  = A167 & A169;
  assign \new_[49259]_  = ~A170 & \new_[49258]_ ;
  assign \new_[49263]_  = A200 & A199;
  assign \new_[49264]_  = A166 & \new_[49263]_ ;
  assign \new_[49265]_  = \new_[49264]_  & \new_[49259]_ ;
  assign \new_[49269]_  = ~A236 & ~A235;
  assign \new_[49270]_  = ~A233 & \new_[49269]_ ;
  assign \new_[49273]_  = A266 & A265;
  assign \new_[49276]_  = A299 & A298;
  assign \new_[49277]_  = \new_[49276]_  & \new_[49273]_ ;
  assign \new_[49278]_  = \new_[49277]_  & \new_[49270]_ ;
  assign \new_[49282]_  = A167 & A169;
  assign \new_[49283]_  = ~A170 & \new_[49282]_ ;
  assign \new_[49287]_  = A200 & A199;
  assign \new_[49288]_  = A166 & \new_[49287]_ ;
  assign \new_[49289]_  = \new_[49288]_  & \new_[49283]_ ;
  assign \new_[49293]_  = ~A236 & ~A235;
  assign \new_[49294]_  = ~A233 & \new_[49293]_ ;
  assign \new_[49297]_  = A266 & A265;
  assign \new_[49300]_  = ~A299 & ~A298;
  assign \new_[49301]_  = \new_[49300]_  & \new_[49297]_ ;
  assign \new_[49302]_  = \new_[49301]_  & \new_[49294]_ ;
  assign \new_[49306]_  = A167 & A169;
  assign \new_[49307]_  = ~A170 & \new_[49306]_ ;
  assign \new_[49311]_  = A200 & A199;
  assign \new_[49312]_  = A166 & \new_[49311]_ ;
  assign \new_[49313]_  = \new_[49312]_  & \new_[49307]_ ;
  assign \new_[49317]_  = ~A236 & ~A235;
  assign \new_[49318]_  = ~A233 & \new_[49317]_ ;
  assign \new_[49321]_  = ~A267 & ~A266;
  assign \new_[49324]_  = ~A300 & A298;
  assign \new_[49325]_  = \new_[49324]_  & \new_[49321]_ ;
  assign \new_[49326]_  = \new_[49325]_  & \new_[49318]_ ;
  assign \new_[49330]_  = A167 & A169;
  assign \new_[49331]_  = ~A170 & \new_[49330]_ ;
  assign \new_[49335]_  = A200 & A199;
  assign \new_[49336]_  = A166 & \new_[49335]_ ;
  assign \new_[49337]_  = \new_[49336]_  & \new_[49331]_ ;
  assign \new_[49341]_  = ~A236 & ~A235;
  assign \new_[49342]_  = ~A233 & \new_[49341]_ ;
  assign \new_[49345]_  = ~A267 & ~A266;
  assign \new_[49348]_  = A299 & A298;
  assign \new_[49349]_  = \new_[49348]_  & \new_[49345]_ ;
  assign \new_[49350]_  = \new_[49349]_  & \new_[49342]_ ;
  assign \new_[49354]_  = A167 & A169;
  assign \new_[49355]_  = ~A170 & \new_[49354]_ ;
  assign \new_[49359]_  = A200 & A199;
  assign \new_[49360]_  = A166 & \new_[49359]_ ;
  assign \new_[49361]_  = \new_[49360]_  & \new_[49355]_ ;
  assign \new_[49365]_  = ~A236 & ~A235;
  assign \new_[49366]_  = ~A233 & \new_[49365]_ ;
  assign \new_[49369]_  = ~A267 & ~A266;
  assign \new_[49372]_  = ~A299 & ~A298;
  assign \new_[49373]_  = \new_[49372]_  & \new_[49369]_ ;
  assign \new_[49374]_  = \new_[49373]_  & \new_[49366]_ ;
  assign \new_[49378]_  = A167 & A169;
  assign \new_[49379]_  = ~A170 & \new_[49378]_ ;
  assign \new_[49383]_  = A200 & A199;
  assign \new_[49384]_  = A166 & \new_[49383]_ ;
  assign \new_[49385]_  = \new_[49384]_  & \new_[49379]_ ;
  assign \new_[49389]_  = ~A236 & ~A235;
  assign \new_[49390]_  = ~A233 & \new_[49389]_ ;
  assign \new_[49393]_  = ~A266 & ~A265;
  assign \new_[49396]_  = ~A300 & A298;
  assign \new_[49397]_  = \new_[49396]_  & \new_[49393]_ ;
  assign \new_[49398]_  = \new_[49397]_  & \new_[49390]_ ;
  assign \new_[49402]_  = A167 & A169;
  assign \new_[49403]_  = ~A170 & \new_[49402]_ ;
  assign \new_[49407]_  = A200 & A199;
  assign \new_[49408]_  = A166 & \new_[49407]_ ;
  assign \new_[49409]_  = \new_[49408]_  & \new_[49403]_ ;
  assign \new_[49413]_  = ~A236 & ~A235;
  assign \new_[49414]_  = ~A233 & \new_[49413]_ ;
  assign \new_[49417]_  = ~A266 & ~A265;
  assign \new_[49420]_  = A299 & A298;
  assign \new_[49421]_  = \new_[49420]_  & \new_[49417]_ ;
  assign \new_[49422]_  = \new_[49421]_  & \new_[49414]_ ;
  assign \new_[49426]_  = A167 & A169;
  assign \new_[49427]_  = ~A170 & \new_[49426]_ ;
  assign \new_[49431]_  = A200 & A199;
  assign \new_[49432]_  = A166 & \new_[49431]_ ;
  assign \new_[49433]_  = \new_[49432]_  & \new_[49427]_ ;
  assign \new_[49437]_  = ~A236 & ~A235;
  assign \new_[49438]_  = ~A233 & \new_[49437]_ ;
  assign \new_[49441]_  = ~A266 & ~A265;
  assign \new_[49444]_  = ~A299 & ~A298;
  assign \new_[49445]_  = \new_[49444]_  & \new_[49441]_ ;
  assign \new_[49446]_  = \new_[49445]_  & \new_[49438]_ ;
  assign \new_[49450]_  = A167 & A169;
  assign \new_[49451]_  = ~A170 & \new_[49450]_ ;
  assign \new_[49455]_  = A200 & A199;
  assign \new_[49456]_  = A166 & \new_[49455]_ ;
  assign \new_[49457]_  = \new_[49456]_  & \new_[49451]_ ;
  assign \new_[49461]_  = A265 & ~A234;
  assign \new_[49462]_  = ~A233 & \new_[49461]_ ;
  assign \new_[49465]_  = A298 & A266;
  assign \new_[49468]_  = ~A302 & ~A301;
  assign \new_[49469]_  = \new_[49468]_  & \new_[49465]_ ;
  assign \new_[49470]_  = \new_[49469]_  & \new_[49462]_ ;
  assign \new_[49474]_  = A167 & A169;
  assign \new_[49475]_  = ~A170 & \new_[49474]_ ;
  assign \new_[49479]_  = A200 & A199;
  assign \new_[49480]_  = A166 & \new_[49479]_ ;
  assign \new_[49481]_  = \new_[49480]_  & \new_[49475]_ ;
  assign \new_[49485]_  = ~A266 & ~A234;
  assign \new_[49486]_  = ~A233 & \new_[49485]_ ;
  assign \new_[49489]_  = ~A269 & ~A268;
  assign \new_[49492]_  = ~A300 & A298;
  assign \new_[49493]_  = \new_[49492]_  & \new_[49489]_ ;
  assign \new_[49494]_  = \new_[49493]_  & \new_[49486]_ ;
  assign \new_[49498]_  = A167 & A169;
  assign \new_[49499]_  = ~A170 & \new_[49498]_ ;
  assign \new_[49503]_  = A200 & A199;
  assign \new_[49504]_  = A166 & \new_[49503]_ ;
  assign \new_[49505]_  = \new_[49504]_  & \new_[49499]_ ;
  assign \new_[49509]_  = ~A266 & ~A234;
  assign \new_[49510]_  = ~A233 & \new_[49509]_ ;
  assign \new_[49513]_  = ~A269 & ~A268;
  assign \new_[49516]_  = A299 & A298;
  assign \new_[49517]_  = \new_[49516]_  & \new_[49513]_ ;
  assign \new_[49518]_  = \new_[49517]_  & \new_[49510]_ ;
  assign \new_[49522]_  = A167 & A169;
  assign \new_[49523]_  = ~A170 & \new_[49522]_ ;
  assign \new_[49527]_  = A200 & A199;
  assign \new_[49528]_  = A166 & \new_[49527]_ ;
  assign \new_[49529]_  = \new_[49528]_  & \new_[49523]_ ;
  assign \new_[49533]_  = ~A266 & ~A234;
  assign \new_[49534]_  = ~A233 & \new_[49533]_ ;
  assign \new_[49537]_  = ~A269 & ~A268;
  assign \new_[49540]_  = ~A299 & ~A298;
  assign \new_[49541]_  = \new_[49540]_  & \new_[49537]_ ;
  assign \new_[49542]_  = \new_[49541]_  & \new_[49534]_ ;
  assign \new_[49546]_  = A167 & A169;
  assign \new_[49547]_  = ~A170 & \new_[49546]_ ;
  assign \new_[49551]_  = A200 & A199;
  assign \new_[49552]_  = A166 & \new_[49551]_ ;
  assign \new_[49553]_  = \new_[49552]_  & \new_[49547]_ ;
  assign \new_[49557]_  = ~A266 & ~A234;
  assign \new_[49558]_  = ~A233 & \new_[49557]_ ;
  assign \new_[49561]_  = A298 & ~A267;
  assign \new_[49564]_  = ~A302 & ~A301;
  assign \new_[49565]_  = \new_[49564]_  & \new_[49561]_ ;
  assign \new_[49566]_  = \new_[49565]_  & \new_[49558]_ ;
  assign \new_[49570]_  = A167 & A169;
  assign \new_[49571]_  = ~A170 & \new_[49570]_ ;
  assign \new_[49575]_  = A200 & A199;
  assign \new_[49576]_  = A166 & \new_[49575]_ ;
  assign \new_[49577]_  = \new_[49576]_  & \new_[49571]_ ;
  assign \new_[49581]_  = ~A265 & ~A234;
  assign \new_[49582]_  = ~A233 & \new_[49581]_ ;
  assign \new_[49585]_  = A298 & ~A266;
  assign \new_[49588]_  = ~A302 & ~A301;
  assign \new_[49589]_  = \new_[49588]_  & \new_[49585]_ ;
  assign \new_[49590]_  = \new_[49589]_  & \new_[49582]_ ;
  assign \new_[49594]_  = A167 & A169;
  assign \new_[49595]_  = ~A170 & \new_[49594]_ ;
  assign \new_[49599]_  = A200 & A199;
  assign \new_[49600]_  = A166 & \new_[49599]_ ;
  assign \new_[49601]_  = \new_[49600]_  & \new_[49595]_ ;
  assign \new_[49605]_  = A265 & ~A233;
  assign \new_[49606]_  = ~A232 & \new_[49605]_ ;
  assign \new_[49609]_  = A298 & A266;
  assign \new_[49612]_  = ~A302 & ~A301;
  assign \new_[49613]_  = \new_[49612]_  & \new_[49609]_ ;
  assign \new_[49614]_  = \new_[49613]_  & \new_[49606]_ ;
  assign \new_[49618]_  = A167 & A169;
  assign \new_[49619]_  = ~A170 & \new_[49618]_ ;
  assign \new_[49623]_  = A200 & A199;
  assign \new_[49624]_  = A166 & \new_[49623]_ ;
  assign \new_[49625]_  = \new_[49624]_  & \new_[49619]_ ;
  assign \new_[49629]_  = ~A266 & ~A233;
  assign \new_[49630]_  = ~A232 & \new_[49629]_ ;
  assign \new_[49633]_  = ~A269 & ~A268;
  assign \new_[49636]_  = ~A300 & A298;
  assign \new_[49637]_  = \new_[49636]_  & \new_[49633]_ ;
  assign \new_[49638]_  = \new_[49637]_  & \new_[49630]_ ;
  assign \new_[49642]_  = A167 & A169;
  assign \new_[49643]_  = ~A170 & \new_[49642]_ ;
  assign \new_[49647]_  = A200 & A199;
  assign \new_[49648]_  = A166 & \new_[49647]_ ;
  assign \new_[49649]_  = \new_[49648]_  & \new_[49643]_ ;
  assign \new_[49653]_  = ~A266 & ~A233;
  assign \new_[49654]_  = ~A232 & \new_[49653]_ ;
  assign \new_[49657]_  = ~A269 & ~A268;
  assign \new_[49660]_  = A299 & A298;
  assign \new_[49661]_  = \new_[49660]_  & \new_[49657]_ ;
  assign \new_[49662]_  = \new_[49661]_  & \new_[49654]_ ;
  assign \new_[49666]_  = A167 & A169;
  assign \new_[49667]_  = ~A170 & \new_[49666]_ ;
  assign \new_[49671]_  = A200 & A199;
  assign \new_[49672]_  = A166 & \new_[49671]_ ;
  assign \new_[49673]_  = \new_[49672]_  & \new_[49667]_ ;
  assign \new_[49677]_  = ~A266 & ~A233;
  assign \new_[49678]_  = ~A232 & \new_[49677]_ ;
  assign \new_[49681]_  = ~A269 & ~A268;
  assign \new_[49684]_  = ~A299 & ~A298;
  assign \new_[49685]_  = \new_[49684]_  & \new_[49681]_ ;
  assign \new_[49686]_  = \new_[49685]_  & \new_[49678]_ ;
  assign \new_[49690]_  = A167 & A169;
  assign \new_[49691]_  = ~A170 & \new_[49690]_ ;
  assign \new_[49695]_  = A200 & A199;
  assign \new_[49696]_  = A166 & \new_[49695]_ ;
  assign \new_[49697]_  = \new_[49696]_  & \new_[49691]_ ;
  assign \new_[49701]_  = ~A266 & ~A233;
  assign \new_[49702]_  = ~A232 & \new_[49701]_ ;
  assign \new_[49705]_  = A298 & ~A267;
  assign \new_[49708]_  = ~A302 & ~A301;
  assign \new_[49709]_  = \new_[49708]_  & \new_[49705]_ ;
  assign \new_[49710]_  = \new_[49709]_  & \new_[49702]_ ;
  assign \new_[49714]_  = A167 & A169;
  assign \new_[49715]_  = ~A170 & \new_[49714]_ ;
  assign \new_[49719]_  = A200 & A199;
  assign \new_[49720]_  = A166 & \new_[49719]_ ;
  assign \new_[49721]_  = \new_[49720]_  & \new_[49715]_ ;
  assign \new_[49725]_  = ~A265 & ~A233;
  assign \new_[49726]_  = ~A232 & \new_[49725]_ ;
  assign \new_[49729]_  = A298 & ~A266;
  assign \new_[49732]_  = ~A302 & ~A301;
  assign \new_[49733]_  = \new_[49732]_  & \new_[49729]_ ;
  assign \new_[49734]_  = \new_[49733]_  & \new_[49726]_ ;
  assign \new_[49738]_  = A167 & A169;
  assign \new_[49739]_  = ~A170 & \new_[49738]_ ;
  assign \new_[49743]_  = ~A202 & ~A200;
  assign \new_[49744]_  = A166 & \new_[49743]_ ;
  assign \new_[49745]_  = \new_[49744]_  & \new_[49739]_ ;
  assign \new_[49749]_  = A233 & A232;
  assign \new_[49750]_  = ~A203 & \new_[49749]_ ;
  assign \new_[49753]_  = ~A267 & A265;
  assign \new_[49756]_  = ~A300 & ~A299;
  assign \new_[49757]_  = \new_[49756]_  & \new_[49753]_ ;
  assign \new_[49758]_  = \new_[49757]_  & \new_[49750]_ ;
  assign \new_[49762]_  = A167 & A169;
  assign \new_[49763]_  = ~A170 & \new_[49762]_ ;
  assign \new_[49767]_  = ~A202 & ~A200;
  assign \new_[49768]_  = A166 & \new_[49767]_ ;
  assign \new_[49769]_  = \new_[49768]_  & \new_[49763]_ ;
  assign \new_[49773]_  = A233 & A232;
  assign \new_[49774]_  = ~A203 & \new_[49773]_ ;
  assign \new_[49777]_  = ~A267 & A265;
  assign \new_[49780]_  = A299 & A298;
  assign \new_[49781]_  = \new_[49780]_  & \new_[49777]_ ;
  assign \new_[49782]_  = \new_[49781]_  & \new_[49774]_ ;
  assign \new_[49786]_  = A167 & A169;
  assign \new_[49787]_  = ~A170 & \new_[49786]_ ;
  assign \new_[49791]_  = ~A202 & ~A200;
  assign \new_[49792]_  = A166 & \new_[49791]_ ;
  assign \new_[49793]_  = \new_[49792]_  & \new_[49787]_ ;
  assign \new_[49797]_  = A233 & A232;
  assign \new_[49798]_  = ~A203 & \new_[49797]_ ;
  assign \new_[49801]_  = ~A267 & A265;
  assign \new_[49804]_  = ~A299 & ~A298;
  assign \new_[49805]_  = \new_[49804]_  & \new_[49801]_ ;
  assign \new_[49806]_  = \new_[49805]_  & \new_[49798]_ ;
  assign \new_[49810]_  = A167 & A169;
  assign \new_[49811]_  = ~A170 & \new_[49810]_ ;
  assign \new_[49815]_  = ~A202 & ~A200;
  assign \new_[49816]_  = A166 & \new_[49815]_ ;
  assign \new_[49817]_  = \new_[49816]_  & \new_[49811]_ ;
  assign \new_[49821]_  = A233 & A232;
  assign \new_[49822]_  = ~A203 & \new_[49821]_ ;
  assign \new_[49825]_  = A266 & A265;
  assign \new_[49828]_  = ~A300 & ~A299;
  assign \new_[49829]_  = \new_[49828]_  & \new_[49825]_ ;
  assign \new_[49830]_  = \new_[49829]_  & \new_[49822]_ ;
  assign \new_[49834]_  = A167 & A169;
  assign \new_[49835]_  = ~A170 & \new_[49834]_ ;
  assign \new_[49839]_  = ~A202 & ~A200;
  assign \new_[49840]_  = A166 & \new_[49839]_ ;
  assign \new_[49841]_  = \new_[49840]_  & \new_[49835]_ ;
  assign \new_[49845]_  = A233 & A232;
  assign \new_[49846]_  = ~A203 & \new_[49845]_ ;
  assign \new_[49849]_  = A266 & A265;
  assign \new_[49852]_  = A299 & A298;
  assign \new_[49853]_  = \new_[49852]_  & \new_[49849]_ ;
  assign \new_[49854]_  = \new_[49853]_  & \new_[49846]_ ;
  assign \new_[49858]_  = A167 & A169;
  assign \new_[49859]_  = ~A170 & \new_[49858]_ ;
  assign \new_[49863]_  = ~A202 & ~A200;
  assign \new_[49864]_  = A166 & \new_[49863]_ ;
  assign \new_[49865]_  = \new_[49864]_  & \new_[49859]_ ;
  assign \new_[49869]_  = A233 & A232;
  assign \new_[49870]_  = ~A203 & \new_[49869]_ ;
  assign \new_[49873]_  = A266 & A265;
  assign \new_[49876]_  = ~A299 & ~A298;
  assign \new_[49877]_  = \new_[49876]_  & \new_[49873]_ ;
  assign \new_[49878]_  = \new_[49877]_  & \new_[49870]_ ;
  assign \new_[49882]_  = A167 & A169;
  assign \new_[49883]_  = ~A170 & \new_[49882]_ ;
  assign \new_[49887]_  = ~A202 & ~A200;
  assign \new_[49888]_  = A166 & \new_[49887]_ ;
  assign \new_[49889]_  = \new_[49888]_  & \new_[49883]_ ;
  assign \new_[49893]_  = A233 & A232;
  assign \new_[49894]_  = ~A203 & \new_[49893]_ ;
  assign \new_[49897]_  = ~A266 & ~A265;
  assign \new_[49900]_  = ~A300 & ~A299;
  assign \new_[49901]_  = \new_[49900]_  & \new_[49897]_ ;
  assign \new_[49902]_  = \new_[49901]_  & \new_[49894]_ ;
  assign \new_[49906]_  = A167 & A169;
  assign \new_[49907]_  = ~A170 & \new_[49906]_ ;
  assign \new_[49911]_  = ~A202 & ~A200;
  assign \new_[49912]_  = A166 & \new_[49911]_ ;
  assign \new_[49913]_  = \new_[49912]_  & \new_[49907]_ ;
  assign \new_[49917]_  = A233 & A232;
  assign \new_[49918]_  = ~A203 & \new_[49917]_ ;
  assign \new_[49921]_  = ~A266 & ~A265;
  assign \new_[49924]_  = A299 & A298;
  assign \new_[49925]_  = \new_[49924]_  & \new_[49921]_ ;
  assign \new_[49926]_  = \new_[49925]_  & \new_[49918]_ ;
  assign \new_[49930]_  = A167 & A169;
  assign \new_[49931]_  = ~A170 & \new_[49930]_ ;
  assign \new_[49935]_  = ~A202 & ~A200;
  assign \new_[49936]_  = A166 & \new_[49935]_ ;
  assign \new_[49937]_  = \new_[49936]_  & \new_[49931]_ ;
  assign \new_[49941]_  = A233 & A232;
  assign \new_[49942]_  = ~A203 & \new_[49941]_ ;
  assign \new_[49945]_  = ~A266 & ~A265;
  assign \new_[49948]_  = ~A299 & ~A298;
  assign \new_[49949]_  = \new_[49948]_  & \new_[49945]_ ;
  assign \new_[49950]_  = \new_[49949]_  & \new_[49942]_ ;
  assign \new_[49954]_  = A167 & A169;
  assign \new_[49955]_  = ~A170 & \new_[49954]_ ;
  assign \new_[49959]_  = ~A202 & ~A200;
  assign \new_[49960]_  = A166 & \new_[49959]_ ;
  assign \new_[49961]_  = \new_[49960]_  & \new_[49955]_ ;
  assign \new_[49965]_  = A233 & ~A232;
  assign \new_[49966]_  = ~A203 & \new_[49965]_ ;
  assign \new_[49969]_  = ~A299 & A298;
  assign \new_[49972]_  = A301 & A300;
  assign \new_[49973]_  = \new_[49972]_  & \new_[49969]_ ;
  assign \new_[49974]_  = \new_[49973]_  & \new_[49966]_ ;
  assign \new_[49978]_  = A167 & A169;
  assign \new_[49979]_  = ~A170 & \new_[49978]_ ;
  assign \new_[49983]_  = ~A202 & ~A200;
  assign \new_[49984]_  = A166 & \new_[49983]_ ;
  assign \new_[49985]_  = \new_[49984]_  & \new_[49979]_ ;
  assign \new_[49989]_  = A233 & ~A232;
  assign \new_[49990]_  = ~A203 & \new_[49989]_ ;
  assign \new_[49993]_  = ~A299 & A298;
  assign \new_[49996]_  = A302 & A300;
  assign \new_[49997]_  = \new_[49996]_  & \new_[49993]_ ;
  assign \new_[49998]_  = \new_[49997]_  & \new_[49990]_ ;
  assign \new_[50002]_  = A167 & A169;
  assign \new_[50003]_  = ~A170 & \new_[50002]_ ;
  assign \new_[50007]_  = ~A202 & ~A200;
  assign \new_[50008]_  = A166 & \new_[50007]_ ;
  assign \new_[50009]_  = \new_[50008]_  & \new_[50003]_ ;
  assign \new_[50013]_  = A233 & ~A232;
  assign \new_[50014]_  = ~A203 & \new_[50013]_ ;
  assign \new_[50017]_  = ~A266 & A265;
  assign \new_[50020]_  = A268 & A267;
  assign \new_[50021]_  = \new_[50020]_  & \new_[50017]_ ;
  assign \new_[50022]_  = \new_[50021]_  & \new_[50014]_ ;
  assign \new_[50026]_  = A167 & A169;
  assign \new_[50027]_  = ~A170 & \new_[50026]_ ;
  assign \new_[50031]_  = ~A202 & ~A200;
  assign \new_[50032]_  = A166 & \new_[50031]_ ;
  assign \new_[50033]_  = \new_[50032]_  & \new_[50027]_ ;
  assign \new_[50037]_  = A233 & ~A232;
  assign \new_[50038]_  = ~A203 & \new_[50037]_ ;
  assign \new_[50041]_  = ~A266 & A265;
  assign \new_[50044]_  = A269 & A267;
  assign \new_[50045]_  = \new_[50044]_  & \new_[50041]_ ;
  assign \new_[50046]_  = \new_[50045]_  & \new_[50038]_ ;
  assign \new_[50050]_  = A167 & A169;
  assign \new_[50051]_  = ~A170 & \new_[50050]_ ;
  assign \new_[50055]_  = ~A202 & ~A200;
  assign \new_[50056]_  = A166 & \new_[50055]_ ;
  assign \new_[50057]_  = \new_[50056]_  & \new_[50051]_ ;
  assign \new_[50061]_  = ~A234 & ~A233;
  assign \new_[50062]_  = ~A203 & \new_[50061]_ ;
  assign \new_[50065]_  = A266 & A265;
  assign \new_[50068]_  = ~A300 & A298;
  assign \new_[50069]_  = \new_[50068]_  & \new_[50065]_ ;
  assign \new_[50070]_  = \new_[50069]_  & \new_[50062]_ ;
  assign \new_[50074]_  = A167 & A169;
  assign \new_[50075]_  = ~A170 & \new_[50074]_ ;
  assign \new_[50079]_  = ~A202 & ~A200;
  assign \new_[50080]_  = A166 & \new_[50079]_ ;
  assign \new_[50081]_  = \new_[50080]_  & \new_[50075]_ ;
  assign \new_[50085]_  = ~A234 & ~A233;
  assign \new_[50086]_  = ~A203 & \new_[50085]_ ;
  assign \new_[50089]_  = A266 & A265;
  assign \new_[50092]_  = A299 & A298;
  assign \new_[50093]_  = \new_[50092]_  & \new_[50089]_ ;
  assign \new_[50094]_  = \new_[50093]_  & \new_[50086]_ ;
  assign \new_[50098]_  = A167 & A169;
  assign \new_[50099]_  = ~A170 & \new_[50098]_ ;
  assign \new_[50103]_  = ~A202 & ~A200;
  assign \new_[50104]_  = A166 & \new_[50103]_ ;
  assign \new_[50105]_  = \new_[50104]_  & \new_[50099]_ ;
  assign \new_[50109]_  = ~A234 & ~A233;
  assign \new_[50110]_  = ~A203 & \new_[50109]_ ;
  assign \new_[50113]_  = A266 & A265;
  assign \new_[50116]_  = ~A299 & ~A298;
  assign \new_[50117]_  = \new_[50116]_  & \new_[50113]_ ;
  assign \new_[50118]_  = \new_[50117]_  & \new_[50110]_ ;
  assign \new_[50122]_  = A167 & A169;
  assign \new_[50123]_  = ~A170 & \new_[50122]_ ;
  assign \new_[50127]_  = ~A202 & ~A200;
  assign \new_[50128]_  = A166 & \new_[50127]_ ;
  assign \new_[50129]_  = \new_[50128]_  & \new_[50123]_ ;
  assign \new_[50133]_  = ~A234 & ~A233;
  assign \new_[50134]_  = ~A203 & \new_[50133]_ ;
  assign \new_[50137]_  = ~A267 & ~A266;
  assign \new_[50140]_  = ~A300 & A298;
  assign \new_[50141]_  = \new_[50140]_  & \new_[50137]_ ;
  assign \new_[50142]_  = \new_[50141]_  & \new_[50134]_ ;
  assign \new_[50146]_  = A167 & A169;
  assign \new_[50147]_  = ~A170 & \new_[50146]_ ;
  assign \new_[50151]_  = ~A202 & ~A200;
  assign \new_[50152]_  = A166 & \new_[50151]_ ;
  assign \new_[50153]_  = \new_[50152]_  & \new_[50147]_ ;
  assign \new_[50157]_  = ~A234 & ~A233;
  assign \new_[50158]_  = ~A203 & \new_[50157]_ ;
  assign \new_[50161]_  = ~A267 & ~A266;
  assign \new_[50164]_  = A299 & A298;
  assign \new_[50165]_  = \new_[50164]_  & \new_[50161]_ ;
  assign \new_[50166]_  = \new_[50165]_  & \new_[50158]_ ;
  assign \new_[50170]_  = A167 & A169;
  assign \new_[50171]_  = ~A170 & \new_[50170]_ ;
  assign \new_[50175]_  = ~A202 & ~A200;
  assign \new_[50176]_  = A166 & \new_[50175]_ ;
  assign \new_[50177]_  = \new_[50176]_  & \new_[50171]_ ;
  assign \new_[50181]_  = ~A234 & ~A233;
  assign \new_[50182]_  = ~A203 & \new_[50181]_ ;
  assign \new_[50185]_  = ~A267 & ~A266;
  assign \new_[50188]_  = ~A299 & ~A298;
  assign \new_[50189]_  = \new_[50188]_  & \new_[50185]_ ;
  assign \new_[50190]_  = \new_[50189]_  & \new_[50182]_ ;
  assign \new_[50194]_  = A167 & A169;
  assign \new_[50195]_  = ~A170 & \new_[50194]_ ;
  assign \new_[50199]_  = ~A202 & ~A200;
  assign \new_[50200]_  = A166 & \new_[50199]_ ;
  assign \new_[50201]_  = \new_[50200]_  & \new_[50195]_ ;
  assign \new_[50205]_  = ~A234 & ~A233;
  assign \new_[50206]_  = ~A203 & \new_[50205]_ ;
  assign \new_[50209]_  = ~A266 & ~A265;
  assign \new_[50212]_  = ~A300 & A298;
  assign \new_[50213]_  = \new_[50212]_  & \new_[50209]_ ;
  assign \new_[50214]_  = \new_[50213]_  & \new_[50206]_ ;
  assign \new_[50218]_  = A167 & A169;
  assign \new_[50219]_  = ~A170 & \new_[50218]_ ;
  assign \new_[50223]_  = ~A202 & ~A200;
  assign \new_[50224]_  = A166 & \new_[50223]_ ;
  assign \new_[50225]_  = \new_[50224]_  & \new_[50219]_ ;
  assign \new_[50229]_  = ~A234 & ~A233;
  assign \new_[50230]_  = ~A203 & \new_[50229]_ ;
  assign \new_[50233]_  = ~A266 & ~A265;
  assign \new_[50236]_  = A299 & A298;
  assign \new_[50237]_  = \new_[50236]_  & \new_[50233]_ ;
  assign \new_[50238]_  = \new_[50237]_  & \new_[50230]_ ;
  assign \new_[50242]_  = A167 & A169;
  assign \new_[50243]_  = ~A170 & \new_[50242]_ ;
  assign \new_[50247]_  = ~A202 & ~A200;
  assign \new_[50248]_  = A166 & \new_[50247]_ ;
  assign \new_[50249]_  = \new_[50248]_  & \new_[50243]_ ;
  assign \new_[50253]_  = ~A234 & ~A233;
  assign \new_[50254]_  = ~A203 & \new_[50253]_ ;
  assign \new_[50257]_  = ~A266 & ~A265;
  assign \new_[50260]_  = ~A299 & ~A298;
  assign \new_[50261]_  = \new_[50260]_  & \new_[50257]_ ;
  assign \new_[50262]_  = \new_[50261]_  & \new_[50254]_ ;
  assign \new_[50266]_  = A167 & A169;
  assign \new_[50267]_  = ~A170 & \new_[50266]_ ;
  assign \new_[50271]_  = ~A202 & ~A200;
  assign \new_[50272]_  = A166 & \new_[50271]_ ;
  assign \new_[50273]_  = \new_[50272]_  & \new_[50267]_ ;
  assign \new_[50277]_  = ~A233 & A232;
  assign \new_[50278]_  = ~A203 & \new_[50277]_ ;
  assign \new_[50281]_  = A235 & A234;
  assign \new_[50284]_  = A299 & ~A298;
  assign \new_[50285]_  = \new_[50284]_  & \new_[50281]_ ;
  assign \new_[50286]_  = \new_[50285]_  & \new_[50278]_ ;
  assign \new_[50290]_  = A167 & A169;
  assign \new_[50291]_  = ~A170 & \new_[50290]_ ;
  assign \new_[50295]_  = ~A202 & ~A200;
  assign \new_[50296]_  = A166 & \new_[50295]_ ;
  assign \new_[50297]_  = \new_[50296]_  & \new_[50291]_ ;
  assign \new_[50301]_  = ~A233 & A232;
  assign \new_[50302]_  = ~A203 & \new_[50301]_ ;
  assign \new_[50305]_  = A235 & A234;
  assign \new_[50308]_  = A266 & ~A265;
  assign \new_[50309]_  = \new_[50308]_  & \new_[50305]_ ;
  assign \new_[50310]_  = \new_[50309]_  & \new_[50302]_ ;
  assign \new_[50314]_  = A167 & A169;
  assign \new_[50315]_  = ~A170 & \new_[50314]_ ;
  assign \new_[50319]_  = ~A202 & ~A200;
  assign \new_[50320]_  = A166 & \new_[50319]_ ;
  assign \new_[50321]_  = \new_[50320]_  & \new_[50315]_ ;
  assign \new_[50325]_  = ~A233 & A232;
  assign \new_[50326]_  = ~A203 & \new_[50325]_ ;
  assign \new_[50329]_  = A236 & A234;
  assign \new_[50332]_  = A299 & ~A298;
  assign \new_[50333]_  = \new_[50332]_  & \new_[50329]_ ;
  assign \new_[50334]_  = \new_[50333]_  & \new_[50326]_ ;
  assign \new_[50338]_  = A167 & A169;
  assign \new_[50339]_  = ~A170 & \new_[50338]_ ;
  assign \new_[50343]_  = ~A202 & ~A200;
  assign \new_[50344]_  = A166 & \new_[50343]_ ;
  assign \new_[50345]_  = \new_[50344]_  & \new_[50339]_ ;
  assign \new_[50349]_  = ~A233 & A232;
  assign \new_[50350]_  = ~A203 & \new_[50349]_ ;
  assign \new_[50353]_  = A236 & A234;
  assign \new_[50356]_  = A266 & ~A265;
  assign \new_[50357]_  = \new_[50356]_  & \new_[50353]_ ;
  assign \new_[50358]_  = \new_[50357]_  & \new_[50350]_ ;
  assign \new_[50362]_  = A167 & A169;
  assign \new_[50363]_  = ~A170 & \new_[50362]_ ;
  assign \new_[50367]_  = ~A202 & ~A200;
  assign \new_[50368]_  = A166 & \new_[50367]_ ;
  assign \new_[50369]_  = \new_[50368]_  & \new_[50363]_ ;
  assign \new_[50373]_  = ~A233 & ~A232;
  assign \new_[50374]_  = ~A203 & \new_[50373]_ ;
  assign \new_[50377]_  = A266 & A265;
  assign \new_[50380]_  = ~A300 & A298;
  assign \new_[50381]_  = \new_[50380]_  & \new_[50377]_ ;
  assign \new_[50382]_  = \new_[50381]_  & \new_[50374]_ ;
  assign \new_[50386]_  = A167 & A169;
  assign \new_[50387]_  = ~A170 & \new_[50386]_ ;
  assign \new_[50391]_  = ~A202 & ~A200;
  assign \new_[50392]_  = A166 & \new_[50391]_ ;
  assign \new_[50393]_  = \new_[50392]_  & \new_[50387]_ ;
  assign \new_[50397]_  = ~A233 & ~A232;
  assign \new_[50398]_  = ~A203 & \new_[50397]_ ;
  assign \new_[50401]_  = A266 & A265;
  assign \new_[50404]_  = A299 & A298;
  assign \new_[50405]_  = \new_[50404]_  & \new_[50401]_ ;
  assign \new_[50406]_  = \new_[50405]_  & \new_[50398]_ ;
  assign \new_[50410]_  = A167 & A169;
  assign \new_[50411]_  = ~A170 & \new_[50410]_ ;
  assign \new_[50415]_  = ~A202 & ~A200;
  assign \new_[50416]_  = A166 & \new_[50415]_ ;
  assign \new_[50417]_  = \new_[50416]_  & \new_[50411]_ ;
  assign \new_[50421]_  = ~A233 & ~A232;
  assign \new_[50422]_  = ~A203 & \new_[50421]_ ;
  assign \new_[50425]_  = A266 & A265;
  assign \new_[50428]_  = ~A299 & ~A298;
  assign \new_[50429]_  = \new_[50428]_  & \new_[50425]_ ;
  assign \new_[50430]_  = \new_[50429]_  & \new_[50422]_ ;
  assign \new_[50434]_  = A167 & A169;
  assign \new_[50435]_  = ~A170 & \new_[50434]_ ;
  assign \new_[50439]_  = ~A202 & ~A200;
  assign \new_[50440]_  = A166 & \new_[50439]_ ;
  assign \new_[50441]_  = \new_[50440]_  & \new_[50435]_ ;
  assign \new_[50445]_  = ~A233 & ~A232;
  assign \new_[50446]_  = ~A203 & \new_[50445]_ ;
  assign \new_[50449]_  = ~A267 & ~A266;
  assign \new_[50452]_  = ~A300 & A298;
  assign \new_[50453]_  = \new_[50452]_  & \new_[50449]_ ;
  assign \new_[50454]_  = \new_[50453]_  & \new_[50446]_ ;
  assign \new_[50458]_  = A167 & A169;
  assign \new_[50459]_  = ~A170 & \new_[50458]_ ;
  assign \new_[50463]_  = ~A202 & ~A200;
  assign \new_[50464]_  = A166 & \new_[50463]_ ;
  assign \new_[50465]_  = \new_[50464]_  & \new_[50459]_ ;
  assign \new_[50469]_  = ~A233 & ~A232;
  assign \new_[50470]_  = ~A203 & \new_[50469]_ ;
  assign \new_[50473]_  = ~A267 & ~A266;
  assign \new_[50476]_  = A299 & A298;
  assign \new_[50477]_  = \new_[50476]_  & \new_[50473]_ ;
  assign \new_[50478]_  = \new_[50477]_  & \new_[50470]_ ;
  assign \new_[50482]_  = A167 & A169;
  assign \new_[50483]_  = ~A170 & \new_[50482]_ ;
  assign \new_[50487]_  = ~A202 & ~A200;
  assign \new_[50488]_  = A166 & \new_[50487]_ ;
  assign \new_[50489]_  = \new_[50488]_  & \new_[50483]_ ;
  assign \new_[50493]_  = ~A233 & ~A232;
  assign \new_[50494]_  = ~A203 & \new_[50493]_ ;
  assign \new_[50497]_  = ~A267 & ~A266;
  assign \new_[50500]_  = ~A299 & ~A298;
  assign \new_[50501]_  = \new_[50500]_  & \new_[50497]_ ;
  assign \new_[50502]_  = \new_[50501]_  & \new_[50494]_ ;
  assign \new_[50506]_  = A167 & A169;
  assign \new_[50507]_  = ~A170 & \new_[50506]_ ;
  assign \new_[50511]_  = ~A202 & ~A200;
  assign \new_[50512]_  = A166 & \new_[50511]_ ;
  assign \new_[50513]_  = \new_[50512]_  & \new_[50507]_ ;
  assign \new_[50517]_  = ~A233 & ~A232;
  assign \new_[50518]_  = ~A203 & \new_[50517]_ ;
  assign \new_[50521]_  = ~A266 & ~A265;
  assign \new_[50524]_  = ~A300 & A298;
  assign \new_[50525]_  = \new_[50524]_  & \new_[50521]_ ;
  assign \new_[50526]_  = \new_[50525]_  & \new_[50518]_ ;
  assign \new_[50530]_  = A167 & A169;
  assign \new_[50531]_  = ~A170 & \new_[50530]_ ;
  assign \new_[50535]_  = ~A202 & ~A200;
  assign \new_[50536]_  = A166 & \new_[50535]_ ;
  assign \new_[50537]_  = \new_[50536]_  & \new_[50531]_ ;
  assign \new_[50541]_  = ~A233 & ~A232;
  assign \new_[50542]_  = ~A203 & \new_[50541]_ ;
  assign \new_[50545]_  = ~A266 & ~A265;
  assign \new_[50548]_  = A299 & A298;
  assign \new_[50549]_  = \new_[50548]_  & \new_[50545]_ ;
  assign \new_[50550]_  = \new_[50549]_  & \new_[50542]_ ;
  assign \new_[50554]_  = A167 & A169;
  assign \new_[50555]_  = ~A170 & \new_[50554]_ ;
  assign \new_[50559]_  = ~A202 & ~A200;
  assign \new_[50560]_  = A166 & \new_[50559]_ ;
  assign \new_[50561]_  = \new_[50560]_  & \new_[50555]_ ;
  assign \new_[50565]_  = ~A233 & ~A232;
  assign \new_[50566]_  = ~A203 & \new_[50565]_ ;
  assign \new_[50569]_  = ~A266 & ~A265;
  assign \new_[50572]_  = ~A299 & ~A298;
  assign \new_[50573]_  = \new_[50572]_  & \new_[50569]_ ;
  assign \new_[50574]_  = \new_[50573]_  & \new_[50566]_ ;
  assign \new_[50578]_  = A167 & A169;
  assign \new_[50579]_  = ~A170 & \new_[50578]_ ;
  assign \new_[50583]_  = ~A201 & ~A200;
  assign \new_[50584]_  = A166 & \new_[50583]_ ;
  assign \new_[50585]_  = \new_[50584]_  & \new_[50579]_ ;
  assign \new_[50589]_  = A265 & A233;
  assign \new_[50590]_  = A232 & \new_[50589]_ ;
  assign \new_[50593]_  = ~A269 & ~A268;
  assign \new_[50596]_  = ~A300 & ~A299;
  assign \new_[50597]_  = \new_[50596]_  & \new_[50593]_ ;
  assign \new_[50598]_  = \new_[50597]_  & \new_[50590]_ ;
  assign \new_[50602]_  = A167 & A169;
  assign \new_[50603]_  = ~A170 & \new_[50602]_ ;
  assign \new_[50607]_  = ~A201 & ~A200;
  assign \new_[50608]_  = A166 & \new_[50607]_ ;
  assign \new_[50609]_  = \new_[50608]_  & \new_[50603]_ ;
  assign \new_[50613]_  = A265 & A233;
  assign \new_[50614]_  = A232 & \new_[50613]_ ;
  assign \new_[50617]_  = ~A269 & ~A268;
  assign \new_[50620]_  = A299 & A298;
  assign \new_[50621]_  = \new_[50620]_  & \new_[50617]_ ;
  assign \new_[50622]_  = \new_[50621]_  & \new_[50614]_ ;
  assign \new_[50626]_  = A167 & A169;
  assign \new_[50627]_  = ~A170 & \new_[50626]_ ;
  assign \new_[50631]_  = ~A201 & ~A200;
  assign \new_[50632]_  = A166 & \new_[50631]_ ;
  assign \new_[50633]_  = \new_[50632]_  & \new_[50627]_ ;
  assign \new_[50637]_  = A265 & A233;
  assign \new_[50638]_  = A232 & \new_[50637]_ ;
  assign \new_[50641]_  = ~A269 & ~A268;
  assign \new_[50644]_  = ~A299 & ~A298;
  assign \new_[50645]_  = \new_[50644]_  & \new_[50641]_ ;
  assign \new_[50646]_  = \new_[50645]_  & \new_[50638]_ ;
  assign \new_[50650]_  = A167 & A169;
  assign \new_[50651]_  = ~A170 & \new_[50650]_ ;
  assign \new_[50655]_  = ~A201 & ~A200;
  assign \new_[50656]_  = A166 & \new_[50655]_ ;
  assign \new_[50657]_  = \new_[50656]_  & \new_[50651]_ ;
  assign \new_[50661]_  = A265 & A233;
  assign \new_[50662]_  = A232 & \new_[50661]_ ;
  assign \new_[50665]_  = ~A299 & ~A267;
  assign \new_[50668]_  = ~A302 & ~A301;
  assign \new_[50669]_  = \new_[50668]_  & \new_[50665]_ ;
  assign \new_[50670]_  = \new_[50669]_  & \new_[50662]_ ;
  assign \new_[50674]_  = A167 & A169;
  assign \new_[50675]_  = ~A170 & \new_[50674]_ ;
  assign \new_[50679]_  = ~A201 & ~A200;
  assign \new_[50680]_  = A166 & \new_[50679]_ ;
  assign \new_[50681]_  = \new_[50680]_  & \new_[50675]_ ;
  assign \new_[50685]_  = A265 & A233;
  assign \new_[50686]_  = A232 & \new_[50685]_ ;
  assign \new_[50689]_  = ~A299 & A266;
  assign \new_[50692]_  = ~A302 & ~A301;
  assign \new_[50693]_  = \new_[50692]_  & \new_[50689]_ ;
  assign \new_[50694]_  = \new_[50693]_  & \new_[50686]_ ;
  assign \new_[50698]_  = A167 & A169;
  assign \new_[50699]_  = ~A170 & \new_[50698]_ ;
  assign \new_[50703]_  = ~A201 & ~A200;
  assign \new_[50704]_  = A166 & \new_[50703]_ ;
  assign \new_[50705]_  = \new_[50704]_  & \new_[50699]_ ;
  assign \new_[50709]_  = ~A265 & A233;
  assign \new_[50710]_  = A232 & \new_[50709]_ ;
  assign \new_[50713]_  = ~A299 & ~A266;
  assign \new_[50716]_  = ~A302 & ~A301;
  assign \new_[50717]_  = \new_[50716]_  & \new_[50713]_ ;
  assign \new_[50718]_  = \new_[50717]_  & \new_[50710]_ ;
  assign \new_[50722]_  = A167 & A169;
  assign \new_[50723]_  = ~A170 & \new_[50722]_ ;
  assign \new_[50727]_  = ~A201 & ~A200;
  assign \new_[50728]_  = A166 & \new_[50727]_ ;
  assign \new_[50729]_  = \new_[50728]_  & \new_[50723]_ ;
  assign \new_[50733]_  = ~A236 & ~A235;
  assign \new_[50734]_  = ~A233 & \new_[50733]_ ;
  assign \new_[50737]_  = A266 & A265;
  assign \new_[50740]_  = ~A300 & A298;
  assign \new_[50741]_  = \new_[50740]_  & \new_[50737]_ ;
  assign \new_[50742]_  = \new_[50741]_  & \new_[50734]_ ;
  assign \new_[50746]_  = A167 & A169;
  assign \new_[50747]_  = ~A170 & \new_[50746]_ ;
  assign \new_[50751]_  = ~A201 & ~A200;
  assign \new_[50752]_  = A166 & \new_[50751]_ ;
  assign \new_[50753]_  = \new_[50752]_  & \new_[50747]_ ;
  assign \new_[50757]_  = ~A236 & ~A235;
  assign \new_[50758]_  = ~A233 & \new_[50757]_ ;
  assign \new_[50761]_  = A266 & A265;
  assign \new_[50764]_  = A299 & A298;
  assign \new_[50765]_  = \new_[50764]_  & \new_[50761]_ ;
  assign \new_[50766]_  = \new_[50765]_  & \new_[50758]_ ;
  assign \new_[50770]_  = A167 & A169;
  assign \new_[50771]_  = ~A170 & \new_[50770]_ ;
  assign \new_[50775]_  = ~A201 & ~A200;
  assign \new_[50776]_  = A166 & \new_[50775]_ ;
  assign \new_[50777]_  = \new_[50776]_  & \new_[50771]_ ;
  assign \new_[50781]_  = ~A236 & ~A235;
  assign \new_[50782]_  = ~A233 & \new_[50781]_ ;
  assign \new_[50785]_  = A266 & A265;
  assign \new_[50788]_  = ~A299 & ~A298;
  assign \new_[50789]_  = \new_[50788]_  & \new_[50785]_ ;
  assign \new_[50790]_  = \new_[50789]_  & \new_[50782]_ ;
  assign \new_[50794]_  = A167 & A169;
  assign \new_[50795]_  = ~A170 & \new_[50794]_ ;
  assign \new_[50799]_  = ~A201 & ~A200;
  assign \new_[50800]_  = A166 & \new_[50799]_ ;
  assign \new_[50801]_  = \new_[50800]_  & \new_[50795]_ ;
  assign \new_[50805]_  = ~A236 & ~A235;
  assign \new_[50806]_  = ~A233 & \new_[50805]_ ;
  assign \new_[50809]_  = ~A267 & ~A266;
  assign \new_[50812]_  = ~A300 & A298;
  assign \new_[50813]_  = \new_[50812]_  & \new_[50809]_ ;
  assign \new_[50814]_  = \new_[50813]_  & \new_[50806]_ ;
  assign \new_[50818]_  = A167 & A169;
  assign \new_[50819]_  = ~A170 & \new_[50818]_ ;
  assign \new_[50823]_  = ~A201 & ~A200;
  assign \new_[50824]_  = A166 & \new_[50823]_ ;
  assign \new_[50825]_  = \new_[50824]_  & \new_[50819]_ ;
  assign \new_[50829]_  = ~A236 & ~A235;
  assign \new_[50830]_  = ~A233 & \new_[50829]_ ;
  assign \new_[50833]_  = ~A267 & ~A266;
  assign \new_[50836]_  = A299 & A298;
  assign \new_[50837]_  = \new_[50836]_  & \new_[50833]_ ;
  assign \new_[50838]_  = \new_[50837]_  & \new_[50830]_ ;
  assign \new_[50842]_  = A167 & A169;
  assign \new_[50843]_  = ~A170 & \new_[50842]_ ;
  assign \new_[50847]_  = ~A201 & ~A200;
  assign \new_[50848]_  = A166 & \new_[50847]_ ;
  assign \new_[50849]_  = \new_[50848]_  & \new_[50843]_ ;
  assign \new_[50853]_  = ~A236 & ~A235;
  assign \new_[50854]_  = ~A233 & \new_[50853]_ ;
  assign \new_[50857]_  = ~A267 & ~A266;
  assign \new_[50860]_  = ~A299 & ~A298;
  assign \new_[50861]_  = \new_[50860]_  & \new_[50857]_ ;
  assign \new_[50862]_  = \new_[50861]_  & \new_[50854]_ ;
  assign \new_[50866]_  = A167 & A169;
  assign \new_[50867]_  = ~A170 & \new_[50866]_ ;
  assign \new_[50871]_  = ~A201 & ~A200;
  assign \new_[50872]_  = A166 & \new_[50871]_ ;
  assign \new_[50873]_  = \new_[50872]_  & \new_[50867]_ ;
  assign \new_[50877]_  = ~A236 & ~A235;
  assign \new_[50878]_  = ~A233 & \new_[50877]_ ;
  assign \new_[50881]_  = ~A266 & ~A265;
  assign \new_[50884]_  = ~A300 & A298;
  assign \new_[50885]_  = \new_[50884]_  & \new_[50881]_ ;
  assign \new_[50886]_  = \new_[50885]_  & \new_[50878]_ ;
  assign \new_[50890]_  = A167 & A169;
  assign \new_[50891]_  = ~A170 & \new_[50890]_ ;
  assign \new_[50895]_  = ~A201 & ~A200;
  assign \new_[50896]_  = A166 & \new_[50895]_ ;
  assign \new_[50897]_  = \new_[50896]_  & \new_[50891]_ ;
  assign \new_[50901]_  = ~A236 & ~A235;
  assign \new_[50902]_  = ~A233 & \new_[50901]_ ;
  assign \new_[50905]_  = ~A266 & ~A265;
  assign \new_[50908]_  = A299 & A298;
  assign \new_[50909]_  = \new_[50908]_  & \new_[50905]_ ;
  assign \new_[50910]_  = \new_[50909]_  & \new_[50902]_ ;
  assign \new_[50914]_  = A167 & A169;
  assign \new_[50915]_  = ~A170 & \new_[50914]_ ;
  assign \new_[50919]_  = ~A201 & ~A200;
  assign \new_[50920]_  = A166 & \new_[50919]_ ;
  assign \new_[50921]_  = \new_[50920]_  & \new_[50915]_ ;
  assign \new_[50925]_  = ~A236 & ~A235;
  assign \new_[50926]_  = ~A233 & \new_[50925]_ ;
  assign \new_[50929]_  = ~A266 & ~A265;
  assign \new_[50932]_  = ~A299 & ~A298;
  assign \new_[50933]_  = \new_[50932]_  & \new_[50929]_ ;
  assign \new_[50934]_  = \new_[50933]_  & \new_[50926]_ ;
  assign \new_[50938]_  = A167 & A169;
  assign \new_[50939]_  = ~A170 & \new_[50938]_ ;
  assign \new_[50943]_  = ~A201 & ~A200;
  assign \new_[50944]_  = A166 & \new_[50943]_ ;
  assign \new_[50945]_  = \new_[50944]_  & \new_[50939]_ ;
  assign \new_[50949]_  = A265 & ~A234;
  assign \new_[50950]_  = ~A233 & \new_[50949]_ ;
  assign \new_[50953]_  = A298 & A266;
  assign \new_[50956]_  = ~A302 & ~A301;
  assign \new_[50957]_  = \new_[50956]_  & \new_[50953]_ ;
  assign \new_[50958]_  = \new_[50957]_  & \new_[50950]_ ;
  assign \new_[50962]_  = A167 & A169;
  assign \new_[50963]_  = ~A170 & \new_[50962]_ ;
  assign \new_[50967]_  = ~A201 & ~A200;
  assign \new_[50968]_  = A166 & \new_[50967]_ ;
  assign \new_[50969]_  = \new_[50968]_  & \new_[50963]_ ;
  assign \new_[50973]_  = ~A266 & ~A234;
  assign \new_[50974]_  = ~A233 & \new_[50973]_ ;
  assign \new_[50977]_  = ~A269 & ~A268;
  assign \new_[50980]_  = ~A300 & A298;
  assign \new_[50981]_  = \new_[50980]_  & \new_[50977]_ ;
  assign \new_[50982]_  = \new_[50981]_  & \new_[50974]_ ;
  assign \new_[50986]_  = A167 & A169;
  assign \new_[50987]_  = ~A170 & \new_[50986]_ ;
  assign \new_[50991]_  = ~A201 & ~A200;
  assign \new_[50992]_  = A166 & \new_[50991]_ ;
  assign \new_[50993]_  = \new_[50992]_  & \new_[50987]_ ;
  assign \new_[50997]_  = ~A266 & ~A234;
  assign \new_[50998]_  = ~A233 & \new_[50997]_ ;
  assign \new_[51001]_  = ~A269 & ~A268;
  assign \new_[51004]_  = A299 & A298;
  assign \new_[51005]_  = \new_[51004]_  & \new_[51001]_ ;
  assign \new_[51006]_  = \new_[51005]_  & \new_[50998]_ ;
  assign \new_[51010]_  = A167 & A169;
  assign \new_[51011]_  = ~A170 & \new_[51010]_ ;
  assign \new_[51015]_  = ~A201 & ~A200;
  assign \new_[51016]_  = A166 & \new_[51015]_ ;
  assign \new_[51017]_  = \new_[51016]_  & \new_[51011]_ ;
  assign \new_[51021]_  = ~A266 & ~A234;
  assign \new_[51022]_  = ~A233 & \new_[51021]_ ;
  assign \new_[51025]_  = ~A269 & ~A268;
  assign \new_[51028]_  = ~A299 & ~A298;
  assign \new_[51029]_  = \new_[51028]_  & \new_[51025]_ ;
  assign \new_[51030]_  = \new_[51029]_  & \new_[51022]_ ;
  assign \new_[51034]_  = A167 & A169;
  assign \new_[51035]_  = ~A170 & \new_[51034]_ ;
  assign \new_[51039]_  = ~A201 & ~A200;
  assign \new_[51040]_  = A166 & \new_[51039]_ ;
  assign \new_[51041]_  = \new_[51040]_  & \new_[51035]_ ;
  assign \new_[51045]_  = ~A266 & ~A234;
  assign \new_[51046]_  = ~A233 & \new_[51045]_ ;
  assign \new_[51049]_  = A298 & ~A267;
  assign \new_[51052]_  = ~A302 & ~A301;
  assign \new_[51053]_  = \new_[51052]_  & \new_[51049]_ ;
  assign \new_[51054]_  = \new_[51053]_  & \new_[51046]_ ;
  assign \new_[51058]_  = A167 & A169;
  assign \new_[51059]_  = ~A170 & \new_[51058]_ ;
  assign \new_[51063]_  = ~A201 & ~A200;
  assign \new_[51064]_  = A166 & \new_[51063]_ ;
  assign \new_[51065]_  = \new_[51064]_  & \new_[51059]_ ;
  assign \new_[51069]_  = ~A265 & ~A234;
  assign \new_[51070]_  = ~A233 & \new_[51069]_ ;
  assign \new_[51073]_  = A298 & ~A266;
  assign \new_[51076]_  = ~A302 & ~A301;
  assign \new_[51077]_  = \new_[51076]_  & \new_[51073]_ ;
  assign \new_[51078]_  = \new_[51077]_  & \new_[51070]_ ;
  assign \new_[51082]_  = A167 & A169;
  assign \new_[51083]_  = ~A170 & \new_[51082]_ ;
  assign \new_[51087]_  = ~A201 & ~A200;
  assign \new_[51088]_  = A166 & \new_[51087]_ ;
  assign \new_[51089]_  = \new_[51088]_  & \new_[51083]_ ;
  assign \new_[51093]_  = A265 & ~A233;
  assign \new_[51094]_  = ~A232 & \new_[51093]_ ;
  assign \new_[51097]_  = A298 & A266;
  assign \new_[51100]_  = ~A302 & ~A301;
  assign \new_[51101]_  = \new_[51100]_  & \new_[51097]_ ;
  assign \new_[51102]_  = \new_[51101]_  & \new_[51094]_ ;
  assign \new_[51106]_  = A167 & A169;
  assign \new_[51107]_  = ~A170 & \new_[51106]_ ;
  assign \new_[51111]_  = ~A201 & ~A200;
  assign \new_[51112]_  = A166 & \new_[51111]_ ;
  assign \new_[51113]_  = \new_[51112]_  & \new_[51107]_ ;
  assign \new_[51117]_  = ~A266 & ~A233;
  assign \new_[51118]_  = ~A232 & \new_[51117]_ ;
  assign \new_[51121]_  = ~A269 & ~A268;
  assign \new_[51124]_  = ~A300 & A298;
  assign \new_[51125]_  = \new_[51124]_  & \new_[51121]_ ;
  assign \new_[51126]_  = \new_[51125]_  & \new_[51118]_ ;
  assign \new_[51130]_  = A167 & A169;
  assign \new_[51131]_  = ~A170 & \new_[51130]_ ;
  assign \new_[51135]_  = ~A201 & ~A200;
  assign \new_[51136]_  = A166 & \new_[51135]_ ;
  assign \new_[51137]_  = \new_[51136]_  & \new_[51131]_ ;
  assign \new_[51141]_  = ~A266 & ~A233;
  assign \new_[51142]_  = ~A232 & \new_[51141]_ ;
  assign \new_[51145]_  = ~A269 & ~A268;
  assign \new_[51148]_  = A299 & A298;
  assign \new_[51149]_  = \new_[51148]_  & \new_[51145]_ ;
  assign \new_[51150]_  = \new_[51149]_  & \new_[51142]_ ;
  assign \new_[51154]_  = A167 & A169;
  assign \new_[51155]_  = ~A170 & \new_[51154]_ ;
  assign \new_[51159]_  = ~A201 & ~A200;
  assign \new_[51160]_  = A166 & \new_[51159]_ ;
  assign \new_[51161]_  = \new_[51160]_  & \new_[51155]_ ;
  assign \new_[51165]_  = ~A266 & ~A233;
  assign \new_[51166]_  = ~A232 & \new_[51165]_ ;
  assign \new_[51169]_  = ~A269 & ~A268;
  assign \new_[51172]_  = ~A299 & ~A298;
  assign \new_[51173]_  = \new_[51172]_  & \new_[51169]_ ;
  assign \new_[51174]_  = \new_[51173]_  & \new_[51166]_ ;
  assign \new_[51178]_  = A167 & A169;
  assign \new_[51179]_  = ~A170 & \new_[51178]_ ;
  assign \new_[51183]_  = ~A201 & ~A200;
  assign \new_[51184]_  = A166 & \new_[51183]_ ;
  assign \new_[51185]_  = \new_[51184]_  & \new_[51179]_ ;
  assign \new_[51189]_  = ~A266 & ~A233;
  assign \new_[51190]_  = ~A232 & \new_[51189]_ ;
  assign \new_[51193]_  = A298 & ~A267;
  assign \new_[51196]_  = ~A302 & ~A301;
  assign \new_[51197]_  = \new_[51196]_  & \new_[51193]_ ;
  assign \new_[51198]_  = \new_[51197]_  & \new_[51190]_ ;
  assign \new_[51202]_  = A167 & A169;
  assign \new_[51203]_  = ~A170 & \new_[51202]_ ;
  assign \new_[51207]_  = ~A201 & ~A200;
  assign \new_[51208]_  = A166 & \new_[51207]_ ;
  assign \new_[51209]_  = \new_[51208]_  & \new_[51203]_ ;
  assign \new_[51213]_  = ~A265 & ~A233;
  assign \new_[51214]_  = ~A232 & \new_[51213]_ ;
  assign \new_[51217]_  = A298 & ~A266;
  assign \new_[51220]_  = ~A302 & ~A301;
  assign \new_[51221]_  = \new_[51220]_  & \new_[51217]_ ;
  assign \new_[51222]_  = \new_[51221]_  & \new_[51214]_ ;
  assign \new_[51226]_  = A167 & A169;
  assign \new_[51227]_  = ~A170 & \new_[51226]_ ;
  assign \new_[51231]_  = ~A200 & ~A199;
  assign \new_[51232]_  = A166 & \new_[51231]_ ;
  assign \new_[51233]_  = \new_[51232]_  & \new_[51227]_ ;
  assign \new_[51237]_  = A265 & A233;
  assign \new_[51238]_  = A232 & \new_[51237]_ ;
  assign \new_[51241]_  = ~A269 & ~A268;
  assign \new_[51244]_  = ~A300 & ~A299;
  assign \new_[51245]_  = \new_[51244]_  & \new_[51241]_ ;
  assign \new_[51246]_  = \new_[51245]_  & \new_[51238]_ ;
  assign \new_[51250]_  = A167 & A169;
  assign \new_[51251]_  = ~A170 & \new_[51250]_ ;
  assign \new_[51255]_  = ~A200 & ~A199;
  assign \new_[51256]_  = A166 & \new_[51255]_ ;
  assign \new_[51257]_  = \new_[51256]_  & \new_[51251]_ ;
  assign \new_[51261]_  = A265 & A233;
  assign \new_[51262]_  = A232 & \new_[51261]_ ;
  assign \new_[51265]_  = ~A269 & ~A268;
  assign \new_[51268]_  = A299 & A298;
  assign \new_[51269]_  = \new_[51268]_  & \new_[51265]_ ;
  assign \new_[51270]_  = \new_[51269]_  & \new_[51262]_ ;
  assign \new_[51274]_  = A167 & A169;
  assign \new_[51275]_  = ~A170 & \new_[51274]_ ;
  assign \new_[51279]_  = ~A200 & ~A199;
  assign \new_[51280]_  = A166 & \new_[51279]_ ;
  assign \new_[51281]_  = \new_[51280]_  & \new_[51275]_ ;
  assign \new_[51285]_  = A265 & A233;
  assign \new_[51286]_  = A232 & \new_[51285]_ ;
  assign \new_[51289]_  = ~A269 & ~A268;
  assign \new_[51292]_  = ~A299 & ~A298;
  assign \new_[51293]_  = \new_[51292]_  & \new_[51289]_ ;
  assign \new_[51294]_  = \new_[51293]_  & \new_[51286]_ ;
  assign \new_[51298]_  = A167 & A169;
  assign \new_[51299]_  = ~A170 & \new_[51298]_ ;
  assign \new_[51303]_  = ~A200 & ~A199;
  assign \new_[51304]_  = A166 & \new_[51303]_ ;
  assign \new_[51305]_  = \new_[51304]_  & \new_[51299]_ ;
  assign \new_[51309]_  = A265 & A233;
  assign \new_[51310]_  = A232 & \new_[51309]_ ;
  assign \new_[51313]_  = ~A299 & ~A267;
  assign \new_[51316]_  = ~A302 & ~A301;
  assign \new_[51317]_  = \new_[51316]_  & \new_[51313]_ ;
  assign \new_[51318]_  = \new_[51317]_  & \new_[51310]_ ;
  assign \new_[51322]_  = A167 & A169;
  assign \new_[51323]_  = ~A170 & \new_[51322]_ ;
  assign \new_[51327]_  = ~A200 & ~A199;
  assign \new_[51328]_  = A166 & \new_[51327]_ ;
  assign \new_[51329]_  = \new_[51328]_  & \new_[51323]_ ;
  assign \new_[51333]_  = A265 & A233;
  assign \new_[51334]_  = A232 & \new_[51333]_ ;
  assign \new_[51337]_  = ~A299 & A266;
  assign \new_[51340]_  = ~A302 & ~A301;
  assign \new_[51341]_  = \new_[51340]_  & \new_[51337]_ ;
  assign \new_[51342]_  = \new_[51341]_  & \new_[51334]_ ;
  assign \new_[51346]_  = A167 & A169;
  assign \new_[51347]_  = ~A170 & \new_[51346]_ ;
  assign \new_[51351]_  = ~A200 & ~A199;
  assign \new_[51352]_  = A166 & \new_[51351]_ ;
  assign \new_[51353]_  = \new_[51352]_  & \new_[51347]_ ;
  assign \new_[51357]_  = ~A265 & A233;
  assign \new_[51358]_  = A232 & \new_[51357]_ ;
  assign \new_[51361]_  = ~A299 & ~A266;
  assign \new_[51364]_  = ~A302 & ~A301;
  assign \new_[51365]_  = \new_[51364]_  & \new_[51361]_ ;
  assign \new_[51366]_  = \new_[51365]_  & \new_[51358]_ ;
  assign \new_[51370]_  = A167 & A169;
  assign \new_[51371]_  = ~A170 & \new_[51370]_ ;
  assign \new_[51375]_  = ~A200 & ~A199;
  assign \new_[51376]_  = A166 & \new_[51375]_ ;
  assign \new_[51377]_  = \new_[51376]_  & \new_[51371]_ ;
  assign \new_[51381]_  = ~A236 & ~A235;
  assign \new_[51382]_  = ~A233 & \new_[51381]_ ;
  assign \new_[51385]_  = A266 & A265;
  assign \new_[51388]_  = ~A300 & A298;
  assign \new_[51389]_  = \new_[51388]_  & \new_[51385]_ ;
  assign \new_[51390]_  = \new_[51389]_  & \new_[51382]_ ;
  assign \new_[51394]_  = A167 & A169;
  assign \new_[51395]_  = ~A170 & \new_[51394]_ ;
  assign \new_[51399]_  = ~A200 & ~A199;
  assign \new_[51400]_  = A166 & \new_[51399]_ ;
  assign \new_[51401]_  = \new_[51400]_  & \new_[51395]_ ;
  assign \new_[51405]_  = ~A236 & ~A235;
  assign \new_[51406]_  = ~A233 & \new_[51405]_ ;
  assign \new_[51409]_  = A266 & A265;
  assign \new_[51412]_  = A299 & A298;
  assign \new_[51413]_  = \new_[51412]_  & \new_[51409]_ ;
  assign \new_[51414]_  = \new_[51413]_  & \new_[51406]_ ;
  assign \new_[51418]_  = A167 & A169;
  assign \new_[51419]_  = ~A170 & \new_[51418]_ ;
  assign \new_[51423]_  = ~A200 & ~A199;
  assign \new_[51424]_  = A166 & \new_[51423]_ ;
  assign \new_[51425]_  = \new_[51424]_  & \new_[51419]_ ;
  assign \new_[51429]_  = ~A236 & ~A235;
  assign \new_[51430]_  = ~A233 & \new_[51429]_ ;
  assign \new_[51433]_  = A266 & A265;
  assign \new_[51436]_  = ~A299 & ~A298;
  assign \new_[51437]_  = \new_[51436]_  & \new_[51433]_ ;
  assign \new_[51438]_  = \new_[51437]_  & \new_[51430]_ ;
  assign \new_[51442]_  = A167 & A169;
  assign \new_[51443]_  = ~A170 & \new_[51442]_ ;
  assign \new_[51447]_  = ~A200 & ~A199;
  assign \new_[51448]_  = A166 & \new_[51447]_ ;
  assign \new_[51449]_  = \new_[51448]_  & \new_[51443]_ ;
  assign \new_[51453]_  = ~A236 & ~A235;
  assign \new_[51454]_  = ~A233 & \new_[51453]_ ;
  assign \new_[51457]_  = ~A267 & ~A266;
  assign \new_[51460]_  = ~A300 & A298;
  assign \new_[51461]_  = \new_[51460]_  & \new_[51457]_ ;
  assign \new_[51462]_  = \new_[51461]_  & \new_[51454]_ ;
  assign \new_[51466]_  = A167 & A169;
  assign \new_[51467]_  = ~A170 & \new_[51466]_ ;
  assign \new_[51471]_  = ~A200 & ~A199;
  assign \new_[51472]_  = A166 & \new_[51471]_ ;
  assign \new_[51473]_  = \new_[51472]_  & \new_[51467]_ ;
  assign \new_[51477]_  = ~A236 & ~A235;
  assign \new_[51478]_  = ~A233 & \new_[51477]_ ;
  assign \new_[51481]_  = ~A267 & ~A266;
  assign \new_[51484]_  = A299 & A298;
  assign \new_[51485]_  = \new_[51484]_  & \new_[51481]_ ;
  assign \new_[51486]_  = \new_[51485]_  & \new_[51478]_ ;
  assign \new_[51490]_  = A167 & A169;
  assign \new_[51491]_  = ~A170 & \new_[51490]_ ;
  assign \new_[51495]_  = ~A200 & ~A199;
  assign \new_[51496]_  = A166 & \new_[51495]_ ;
  assign \new_[51497]_  = \new_[51496]_  & \new_[51491]_ ;
  assign \new_[51501]_  = ~A236 & ~A235;
  assign \new_[51502]_  = ~A233 & \new_[51501]_ ;
  assign \new_[51505]_  = ~A267 & ~A266;
  assign \new_[51508]_  = ~A299 & ~A298;
  assign \new_[51509]_  = \new_[51508]_  & \new_[51505]_ ;
  assign \new_[51510]_  = \new_[51509]_  & \new_[51502]_ ;
  assign \new_[51514]_  = A167 & A169;
  assign \new_[51515]_  = ~A170 & \new_[51514]_ ;
  assign \new_[51519]_  = ~A200 & ~A199;
  assign \new_[51520]_  = A166 & \new_[51519]_ ;
  assign \new_[51521]_  = \new_[51520]_  & \new_[51515]_ ;
  assign \new_[51525]_  = ~A236 & ~A235;
  assign \new_[51526]_  = ~A233 & \new_[51525]_ ;
  assign \new_[51529]_  = ~A266 & ~A265;
  assign \new_[51532]_  = ~A300 & A298;
  assign \new_[51533]_  = \new_[51532]_  & \new_[51529]_ ;
  assign \new_[51534]_  = \new_[51533]_  & \new_[51526]_ ;
  assign \new_[51538]_  = A167 & A169;
  assign \new_[51539]_  = ~A170 & \new_[51538]_ ;
  assign \new_[51543]_  = ~A200 & ~A199;
  assign \new_[51544]_  = A166 & \new_[51543]_ ;
  assign \new_[51545]_  = \new_[51544]_  & \new_[51539]_ ;
  assign \new_[51549]_  = ~A236 & ~A235;
  assign \new_[51550]_  = ~A233 & \new_[51549]_ ;
  assign \new_[51553]_  = ~A266 & ~A265;
  assign \new_[51556]_  = A299 & A298;
  assign \new_[51557]_  = \new_[51556]_  & \new_[51553]_ ;
  assign \new_[51558]_  = \new_[51557]_  & \new_[51550]_ ;
  assign \new_[51562]_  = A167 & A169;
  assign \new_[51563]_  = ~A170 & \new_[51562]_ ;
  assign \new_[51567]_  = ~A200 & ~A199;
  assign \new_[51568]_  = A166 & \new_[51567]_ ;
  assign \new_[51569]_  = \new_[51568]_  & \new_[51563]_ ;
  assign \new_[51573]_  = ~A236 & ~A235;
  assign \new_[51574]_  = ~A233 & \new_[51573]_ ;
  assign \new_[51577]_  = ~A266 & ~A265;
  assign \new_[51580]_  = ~A299 & ~A298;
  assign \new_[51581]_  = \new_[51580]_  & \new_[51577]_ ;
  assign \new_[51582]_  = \new_[51581]_  & \new_[51574]_ ;
  assign \new_[51586]_  = A167 & A169;
  assign \new_[51587]_  = ~A170 & \new_[51586]_ ;
  assign \new_[51591]_  = ~A200 & ~A199;
  assign \new_[51592]_  = A166 & \new_[51591]_ ;
  assign \new_[51593]_  = \new_[51592]_  & \new_[51587]_ ;
  assign \new_[51597]_  = A265 & ~A234;
  assign \new_[51598]_  = ~A233 & \new_[51597]_ ;
  assign \new_[51601]_  = A298 & A266;
  assign \new_[51604]_  = ~A302 & ~A301;
  assign \new_[51605]_  = \new_[51604]_  & \new_[51601]_ ;
  assign \new_[51606]_  = \new_[51605]_  & \new_[51598]_ ;
  assign \new_[51610]_  = A167 & A169;
  assign \new_[51611]_  = ~A170 & \new_[51610]_ ;
  assign \new_[51615]_  = ~A200 & ~A199;
  assign \new_[51616]_  = A166 & \new_[51615]_ ;
  assign \new_[51617]_  = \new_[51616]_  & \new_[51611]_ ;
  assign \new_[51621]_  = ~A266 & ~A234;
  assign \new_[51622]_  = ~A233 & \new_[51621]_ ;
  assign \new_[51625]_  = ~A269 & ~A268;
  assign \new_[51628]_  = ~A300 & A298;
  assign \new_[51629]_  = \new_[51628]_  & \new_[51625]_ ;
  assign \new_[51630]_  = \new_[51629]_  & \new_[51622]_ ;
  assign \new_[51634]_  = A167 & A169;
  assign \new_[51635]_  = ~A170 & \new_[51634]_ ;
  assign \new_[51639]_  = ~A200 & ~A199;
  assign \new_[51640]_  = A166 & \new_[51639]_ ;
  assign \new_[51641]_  = \new_[51640]_  & \new_[51635]_ ;
  assign \new_[51645]_  = ~A266 & ~A234;
  assign \new_[51646]_  = ~A233 & \new_[51645]_ ;
  assign \new_[51649]_  = ~A269 & ~A268;
  assign \new_[51652]_  = A299 & A298;
  assign \new_[51653]_  = \new_[51652]_  & \new_[51649]_ ;
  assign \new_[51654]_  = \new_[51653]_  & \new_[51646]_ ;
  assign \new_[51658]_  = A167 & A169;
  assign \new_[51659]_  = ~A170 & \new_[51658]_ ;
  assign \new_[51663]_  = ~A200 & ~A199;
  assign \new_[51664]_  = A166 & \new_[51663]_ ;
  assign \new_[51665]_  = \new_[51664]_  & \new_[51659]_ ;
  assign \new_[51669]_  = ~A266 & ~A234;
  assign \new_[51670]_  = ~A233 & \new_[51669]_ ;
  assign \new_[51673]_  = ~A269 & ~A268;
  assign \new_[51676]_  = ~A299 & ~A298;
  assign \new_[51677]_  = \new_[51676]_  & \new_[51673]_ ;
  assign \new_[51678]_  = \new_[51677]_  & \new_[51670]_ ;
  assign \new_[51682]_  = A167 & A169;
  assign \new_[51683]_  = ~A170 & \new_[51682]_ ;
  assign \new_[51687]_  = ~A200 & ~A199;
  assign \new_[51688]_  = A166 & \new_[51687]_ ;
  assign \new_[51689]_  = \new_[51688]_  & \new_[51683]_ ;
  assign \new_[51693]_  = ~A266 & ~A234;
  assign \new_[51694]_  = ~A233 & \new_[51693]_ ;
  assign \new_[51697]_  = A298 & ~A267;
  assign \new_[51700]_  = ~A302 & ~A301;
  assign \new_[51701]_  = \new_[51700]_  & \new_[51697]_ ;
  assign \new_[51702]_  = \new_[51701]_  & \new_[51694]_ ;
  assign \new_[51706]_  = A167 & A169;
  assign \new_[51707]_  = ~A170 & \new_[51706]_ ;
  assign \new_[51711]_  = ~A200 & ~A199;
  assign \new_[51712]_  = A166 & \new_[51711]_ ;
  assign \new_[51713]_  = \new_[51712]_  & \new_[51707]_ ;
  assign \new_[51717]_  = ~A265 & ~A234;
  assign \new_[51718]_  = ~A233 & \new_[51717]_ ;
  assign \new_[51721]_  = A298 & ~A266;
  assign \new_[51724]_  = ~A302 & ~A301;
  assign \new_[51725]_  = \new_[51724]_  & \new_[51721]_ ;
  assign \new_[51726]_  = \new_[51725]_  & \new_[51718]_ ;
  assign \new_[51730]_  = A167 & A169;
  assign \new_[51731]_  = ~A170 & \new_[51730]_ ;
  assign \new_[51735]_  = ~A200 & ~A199;
  assign \new_[51736]_  = A166 & \new_[51735]_ ;
  assign \new_[51737]_  = \new_[51736]_  & \new_[51731]_ ;
  assign \new_[51741]_  = A265 & ~A233;
  assign \new_[51742]_  = ~A232 & \new_[51741]_ ;
  assign \new_[51745]_  = A298 & A266;
  assign \new_[51748]_  = ~A302 & ~A301;
  assign \new_[51749]_  = \new_[51748]_  & \new_[51745]_ ;
  assign \new_[51750]_  = \new_[51749]_  & \new_[51742]_ ;
  assign \new_[51754]_  = A167 & A169;
  assign \new_[51755]_  = ~A170 & \new_[51754]_ ;
  assign \new_[51759]_  = ~A200 & ~A199;
  assign \new_[51760]_  = A166 & \new_[51759]_ ;
  assign \new_[51761]_  = \new_[51760]_  & \new_[51755]_ ;
  assign \new_[51765]_  = ~A266 & ~A233;
  assign \new_[51766]_  = ~A232 & \new_[51765]_ ;
  assign \new_[51769]_  = ~A269 & ~A268;
  assign \new_[51772]_  = ~A300 & A298;
  assign \new_[51773]_  = \new_[51772]_  & \new_[51769]_ ;
  assign \new_[51774]_  = \new_[51773]_  & \new_[51766]_ ;
  assign \new_[51778]_  = A167 & A169;
  assign \new_[51779]_  = ~A170 & \new_[51778]_ ;
  assign \new_[51783]_  = ~A200 & ~A199;
  assign \new_[51784]_  = A166 & \new_[51783]_ ;
  assign \new_[51785]_  = \new_[51784]_  & \new_[51779]_ ;
  assign \new_[51789]_  = ~A266 & ~A233;
  assign \new_[51790]_  = ~A232 & \new_[51789]_ ;
  assign \new_[51793]_  = ~A269 & ~A268;
  assign \new_[51796]_  = A299 & A298;
  assign \new_[51797]_  = \new_[51796]_  & \new_[51793]_ ;
  assign \new_[51798]_  = \new_[51797]_  & \new_[51790]_ ;
  assign \new_[51802]_  = A167 & A169;
  assign \new_[51803]_  = ~A170 & \new_[51802]_ ;
  assign \new_[51807]_  = ~A200 & ~A199;
  assign \new_[51808]_  = A166 & \new_[51807]_ ;
  assign \new_[51809]_  = \new_[51808]_  & \new_[51803]_ ;
  assign \new_[51813]_  = ~A266 & ~A233;
  assign \new_[51814]_  = ~A232 & \new_[51813]_ ;
  assign \new_[51817]_  = ~A269 & ~A268;
  assign \new_[51820]_  = ~A299 & ~A298;
  assign \new_[51821]_  = \new_[51820]_  & \new_[51817]_ ;
  assign \new_[51822]_  = \new_[51821]_  & \new_[51814]_ ;
  assign \new_[51826]_  = A167 & A169;
  assign \new_[51827]_  = ~A170 & \new_[51826]_ ;
  assign \new_[51831]_  = ~A200 & ~A199;
  assign \new_[51832]_  = A166 & \new_[51831]_ ;
  assign \new_[51833]_  = \new_[51832]_  & \new_[51827]_ ;
  assign \new_[51837]_  = ~A266 & ~A233;
  assign \new_[51838]_  = ~A232 & \new_[51837]_ ;
  assign \new_[51841]_  = A298 & ~A267;
  assign \new_[51844]_  = ~A302 & ~A301;
  assign \new_[51845]_  = \new_[51844]_  & \new_[51841]_ ;
  assign \new_[51846]_  = \new_[51845]_  & \new_[51838]_ ;
  assign \new_[51850]_  = A167 & A169;
  assign \new_[51851]_  = ~A170 & \new_[51850]_ ;
  assign \new_[51855]_  = ~A200 & ~A199;
  assign \new_[51856]_  = A166 & \new_[51855]_ ;
  assign \new_[51857]_  = \new_[51856]_  & \new_[51851]_ ;
  assign \new_[51861]_  = ~A265 & ~A233;
  assign \new_[51862]_  = ~A232 & \new_[51861]_ ;
  assign \new_[51865]_  = A298 & ~A266;
  assign \new_[51868]_  = ~A302 & ~A301;
  assign \new_[51869]_  = \new_[51868]_  & \new_[51865]_ ;
  assign \new_[51870]_  = \new_[51869]_  & \new_[51862]_ ;
  assign \new_[51874]_  = ~A167 & A169;
  assign \new_[51875]_  = ~A170 & \new_[51874]_ ;
  assign \new_[51879]_  = A200 & A199;
  assign \new_[51880]_  = ~A166 & \new_[51879]_ ;
  assign \new_[51881]_  = \new_[51880]_  & \new_[51875]_ ;
  assign \new_[51885]_  = A265 & A233;
  assign \new_[51886]_  = A232 & \new_[51885]_ ;
  assign \new_[51889]_  = ~A269 & ~A268;
  assign \new_[51892]_  = ~A300 & ~A299;
  assign \new_[51893]_  = \new_[51892]_  & \new_[51889]_ ;
  assign \new_[51894]_  = \new_[51893]_  & \new_[51886]_ ;
  assign \new_[51898]_  = ~A167 & A169;
  assign \new_[51899]_  = ~A170 & \new_[51898]_ ;
  assign \new_[51903]_  = A200 & A199;
  assign \new_[51904]_  = ~A166 & \new_[51903]_ ;
  assign \new_[51905]_  = \new_[51904]_  & \new_[51899]_ ;
  assign \new_[51909]_  = A265 & A233;
  assign \new_[51910]_  = A232 & \new_[51909]_ ;
  assign \new_[51913]_  = ~A269 & ~A268;
  assign \new_[51916]_  = A299 & A298;
  assign \new_[51917]_  = \new_[51916]_  & \new_[51913]_ ;
  assign \new_[51918]_  = \new_[51917]_  & \new_[51910]_ ;
  assign \new_[51922]_  = ~A167 & A169;
  assign \new_[51923]_  = ~A170 & \new_[51922]_ ;
  assign \new_[51927]_  = A200 & A199;
  assign \new_[51928]_  = ~A166 & \new_[51927]_ ;
  assign \new_[51929]_  = \new_[51928]_  & \new_[51923]_ ;
  assign \new_[51933]_  = A265 & A233;
  assign \new_[51934]_  = A232 & \new_[51933]_ ;
  assign \new_[51937]_  = ~A269 & ~A268;
  assign \new_[51940]_  = ~A299 & ~A298;
  assign \new_[51941]_  = \new_[51940]_  & \new_[51937]_ ;
  assign \new_[51942]_  = \new_[51941]_  & \new_[51934]_ ;
  assign \new_[51946]_  = ~A167 & A169;
  assign \new_[51947]_  = ~A170 & \new_[51946]_ ;
  assign \new_[51951]_  = A200 & A199;
  assign \new_[51952]_  = ~A166 & \new_[51951]_ ;
  assign \new_[51953]_  = \new_[51952]_  & \new_[51947]_ ;
  assign \new_[51957]_  = A265 & A233;
  assign \new_[51958]_  = A232 & \new_[51957]_ ;
  assign \new_[51961]_  = ~A299 & ~A267;
  assign \new_[51964]_  = ~A302 & ~A301;
  assign \new_[51965]_  = \new_[51964]_  & \new_[51961]_ ;
  assign \new_[51966]_  = \new_[51965]_  & \new_[51958]_ ;
  assign \new_[51970]_  = ~A167 & A169;
  assign \new_[51971]_  = ~A170 & \new_[51970]_ ;
  assign \new_[51975]_  = A200 & A199;
  assign \new_[51976]_  = ~A166 & \new_[51975]_ ;
  assign \new_[51977]_  = \new_[51976]_  & \new_[51971]_ ;
  assign \new_[51981]_  = A265 & A233;
  assign \new_[51982]_  = A232 & \new_[51981]_ ;
  assign \new_[51985]_  = ~A299 & A266;
  assign \new_[51988]_  = ~A302 & ~A301;
  assign \new_[51989]_  = \new_[51988]_  & \new_[51985]_ ;
  assign \new_[51990]_  = \new_[51989]_  & \new_[51982]_ ;
  assign \new_[51994]_  = ~A167 & A169;
  assign \new_[51995]_  = ~A170 & \new_[51994]_ ;
  assign \new_[51999]_  = A200 & A199;
  assign \new_[52000]_  = ~A166 & \new_[51999]_ ;
  assign \new_[52001]_  = \new_[52000]_  & \new_[51995]_ ;
  assign \new_[52005]_  = ~A265 & A233;
  assign \new_[52006]_  = A232 & \new_[52005]_ ;
  assign \new_[52009]_  = ~A299 & ~A266;
  assign \new_[52012]_  = ~A302 & ~A301;
  assign \new_[52013]_  = \new_[52012]_  & \new_[52009]_ ;
  assign \new_[52014]_  = \new_[52013]_  & \new_[52006]_ ;
  assign \new_[52018]_  = ~A167 & A169;
  assign \new_[52019]_  = ~A170 & \new_[52018]_ ;
  assign \new_[52023]_  = A200 & A199;
  assign \new_[52024]_  = ~A166 & \new_[52023]_ ;
  assign \new_[52025]_  = \new_[52024]_  & \new_[52019]_ ;
  assign \new_[52029]_  = ~A236 & ~A235;
  assign \new_[52030]_  = ~A233 & \new_[52029]_ ;
  assign \new_[52033]_  = A266 & A265;
  assign \new_[52036]_  = ~A300 & A298;
  assign \new_[52037]_  = \new_[52036]_  & \new_[52033]_ ;
  assign \new_[52038]_  = \new_[52037]_  & \new_[52030]_ ;
  assign \new_[52042]_  = ~A167 & A169;
  assign \new_[52043]_  = ~A170 & \new_[52042]_ ;
  assign \new_[52047]_  = A200 & A199;
  assign \new_[52048]_  = ~A166 & \new_[52047]_ ;
  assign \new_[52049]_  = \new_[52048]_  & \new_[52043]_ ;
  assign \new_[52053]_  = ~A236 & ~A235;
  assign \new_[52054]_  = ~A233 & \new_[52053]_ ;
  assign \new_[52057]_  = A266 & A265;
  assign \new_[52060]_  = A299 & A298;
  assign \new_[52061]_  = \new_[52060]_  & \new_[52057]_ ;
  assign \new_[52062]_  = \new_[52061]_  & \new_[52054]_ ;
  assign \new_[52066]_  = ~A167 & A169;
  assign \new_[52067]_  = ~A170 & \new_[52066]_ ;
  assign \new_[52071]_  = A200 & A199;
  assign \new_[52072]_  = ~A166 & \new_[52071]_ ;
  assign \new_[52073]_  = \new_[52072]_  & \new_[52067]_ ;
  assign \new_[52077]_  = ~A236 & ~A235;
  assign \new_[52078]_  = ~A233 & \new_[52077]_ ;
  assign \new_[52081]_  = A266 & A265;
  assign \new_[52084]_  = ~A299 & ~A298;
  assign \new_[52085]_  = \new_[52084]_  & \new_[52081]_ ;
  assign \new_[52086]_  = \new_[52085]_  & \new_[52078]_ ;
  assign \new_[52090]_  = ~A167 & A169;
  assign \new_[52091]_  = ~A170 & \new_[52090]_ ;
  assign \new_[52095]_  = A200 & A199;
  assign \new_[52096]_  = ~A166 & \new_[52095]_ ;
  assign \new_[52097]_  = \new_[52096]_  & \new_[52091]_ ;
  assign \new_[52101]_  = ~A236 & ~A235;
  assign \new_[52102]_  = ~A233 & \new_[52101]_ ;
  assign \new_[52105]_  = ~A267 & ~A266;
  assign \new_[52108]_  = ~A300 & A298;
  assign \new_[52109]_  = \new_[52108]_  & \new_[52105]_ ;
  assign \new_[52110]_  = \new_[52109]_  & \new_[52102]_ ;
  assign \new_[52114]_  = ~A167 & A169;
  assign \new_[52115]_  = ~A170 & \new_[52114]_ ;
  assign \new_[52119]_  = A200 & A199;
  assign \new_[52120]_  = ~A166 & \new_[52119]_ ;
  assign \new_[52121]_  = \new_[52120]_  & \new_[52115]_ ;
  assign \new_[52125]_  = ~A236 & ~A235;
  assign \new_[52126]_  = ~A233 & \new_[52125]_ ;
  assign \new_[52129]_  = ~A267 & ~A266;
  assign \new_[52132]_  = A299 & A298;
  assign \new_[52133]_  = \new_[52132]_  & \new_[52129]_ ;
  assign \new_[52134]_  = \new_[52133]_  & \new_[52126]_ ;
  assign \new_[52138]_  = ~A167 & A169;
  assign \new_[52139]_  = ~A170 & \new_[52138]_ ;
  assign \new_[52143]_  = A200 & A199;
  assign \new_[52144]_  = ~A166 & \new_[52143]_ ;
  assign \new_[52145]_  = \new_[52144]_  & \new_[52139]_ ;
  assign \new_[52149]_  = ~A236 & ~A235;
  assign \new_[52150]_  = ~A233 & \new_[52149]_ ;
  assign \new_[52153]_  = ~A267 & ~A266;
  assign \new_[52156]_  = ~A299 & ~A298;
  assign \new_[52157]_  = \new_[52156]_  & \new_[52153]_ ;
  assign \new_[52158]_  = \new_[52157]_  & \new_[52150]_ ;
  assign \new_[52162]_  = ~A167 & A169;
  assign \new_[52163]_  = ~A170 & \new_[52162]_ ;
  assign \new_[52167]_  = A200 & A199;
  assign \new_[52168]_  = ~A166 & \new_[52167]_ ;
  assign \new_[52169]_  = \new_[52168]_  & \new_[52163]_ ;
  assign \new_[52173]_  = ~A236 & ~A235;
  assign \new_[52174]_  = ~A233 & \new_[52173]_ ;
  assign \new_[52177]_  = ~A266 & ~A265;
  assign \new_[52180]_  = ~A300 & A298;
  assign \new_[52181]_  = \new_[52180]_  & \new_[52177]_ ;
  assign \new_[52182]_  = \new_[52181]_  & \new_[52174]_ ;
  assign \new_[52186]_  = ~A167 & A169;
  assign \new_[52187]_  = ~A170 & \new_[52186]_ ;
  assign \new_[52191]_  = A200 & A199;
  assign \new_[52192]_  = ~A166 & \new_[52191]_ ;
  assign \new_[52193]_  = \new_[52192]_  & \new_[52187]_ ;
  assign \new_[52197]_  = ~A236 & ~A235;
  assign \new_[52198]_  = ~A233 & \new_[52197]_ ;
  assign \new_[52201]_  = ~A266 & ~A265;
  assign \new_[52204]_  = A299 & A298;
  assign \new_[52205]_  = \new_[52204]_  & \new_[52201]_ ;
  assign \new_[52206]_  = \new_[52205]_  & \new_[52198]_ ;
  assign \new_[52210]_  = ~A167 & A169;
  assign \new_[52211]_  = ~A170 & \new_[52210]_ ;
  assign \new_[52215]_  = A200 & A199;
  assign \new_[52216]_  = ~A166 & \new_[52215]_ ;
  assign \new_[52217]_  = \new_[52216]_  & \new_[52211]_ ;
  assign \new_[52221]_  = ~A236 & ~A235;
  assign \new_[52222]_  = ~A233 & \new_[52221]_ ;
  assign \new_[52225]_  = ~A266 & ~A265;
  assign \new_[52228]_  = ~A299 & ~A298;
  assign \new_[52229]_  = \new_[52228]_  & \new_[52225]_ ;
  assign \new_[52230]_  = \new_[52229]_  & \new_[52222]_ ;
  assign \new_[52234]_  = ~A167 & A169;
  assign \new_[52235]_  = ~A170 & \new_[52234]_ ;
  assign \new_[52239]_  = A200 & A199;
  assign \new_[52240]_  = ~A166 & \new_[52239]_ ;
  assign \new_[52241]_  = \new_[52240]_  & \new_[52235]_ ;
  assign \new_[52245]_  = A265 & ~A234;
  assign \new_[52246]_  = ~A233 & \new_[52245]_ ;
  assign \new_[52249]_  = A298 & A266;
  assign \new_[52252]_  = ~A302 & ~A301;
  assign \new_[52253]_  = \new_[52252]_  & \new_[52249]_ ;
  assign \new_[52254]_  = \new_[52253]_  & \new_[52246]_ ;
  assign \new_[52258]_  = ~A167 & A169;
  assign \new_[52259]_  = ~A170 & \new_[52258]_ ;
  assign \new_[52263]_  = A200 & A199;
  assign \new_[52264]_  = ~A166 & \new_[52263]_ ;
  assign \new_[52265]_  = \new_[52264]_  & \new_[52259]_ ;
  assign \new_[52269]_  = ~A266 & ~A234;
  assign \new_[52270]_  = ~A233 & \new_[52269]_ ;
  assign \new_[52273]_  = ~A269 & ~A268;
  assign \new_[52276]_  = ~A300 & A298;
  assign \new_[52277]_  = \new_[52276]_  & \new_[52273]_ ;
  assign \new_[52278]_  = \new_[52277]_  & \new_[52270]_ ;
  assign \new_[52282]_  = ~A167 & A169;
  assign \new_[52283]_  = ~A170 & \new_[52282]_ ;
  assign \new_[52287]_  = A200 & A199;
  assign \new_[52288]_  = ~A166 & \new_[52287]_ ;
  assign \new_[52289]_  = \new_[52288]_  & \new_[52283]_ ;
  assign \new_[52293]_  = ~A266 & ~A234;
  assign \new_[52294]_  = ~A233 & \new_[52293]_ ;
  assign \new_[52297]_  = ~A269 & ~A268;
  assign \new_[52300]_  = A299 & A298;
  assign \new_[52301]_  = \new_[52300]_  & \new_[52297]_ ;
  assign \new_[52302]_  = \new_[52301]_  & \new_[52294]_ ;
  assign \new_[52306]_  = ~A167 & A169;
  assign \new_[52307]_  = ~A170 & \new_[52306]_ ;
  assign \new_[52311]_  = A200 & A199;
  assign \new_[52312]_  = ~A166 & \new_[52311]_ ;
  assign \new_[52313]_  = \new_[52312]_  & \new_[52307]_ ;
  assign \new_[52317]_  = ~A266 & ~A234;
  assign \new_[52318]_  = ~A233 & \new_[52317]_ ;
  assign \new_[52321]_  = ~A269 & ~A268;
  assign \new_[52324]_  = ~A299 & ~A298;
  assign \new_[52325]_  = \new_[52324]_  & \new_[52321]_ ;
  assign \new_[52326]_  = \new_[52325]_  & \new_[52318]_ ;
  assign \new_[52330]_  = ~A167 & A169;
  assign \new_[52331]_  = ~A170 & \new_[52330]_ ;
  assign \new_[52335]_  = A200 & A199;
  assign \new_[52336]_  = ~A166 & \new_[52335]_ ;
  assign \new_[52337]_  = \new_[52336]_  & \new_[52331]_ ;
  assign \new_[52341]_  = ~A266 & ~A234;
  assign \new_[52342]_  = ~A233 & \new_[52341]_ ;
  assign \new_[52345]_  = A298 & ~A267;
  assign \new_[52348]_  = ~A302 & ~A301;
  assign \new_[52349]_  = \new_[52348]_  & \new_[52345]_ ;
  assign \new_[52350]_  = \new_[52349]_  & \new_[52342]_ ;
  assign \new_[52354]_  = ~A167 & A169;
  assign \new_[52355]_  = ~A170 & \new_[52354]_ ;
  assign \new_[52359]_  = A200 & A199;
  assign \new_[52360]_  = ~A166 & \new_[52359]_ ;
  assign \new_[52361]_  = \new_[52360]_  & \new_[52355]_ ;
  assign \new_[52365]_  = ~A265 & ~A234;
  assign \new_[52366]_  = ~A233 & \new_[52365]_ ;
  assign \new_[52369]_  = A298 & ~A266;
  assign \new_[52372]_  = ~A302 & ~A301;
  assign \new_[52373]_  = \new_[52372]_  & \new_[52369]_ ;
  assign \new_[52374]_  = \new_[52373]_  & \new_[52366]_ ;
  assign \new_[52378]_  = ~A167 & A169;
  assign \new_[52379]_  = ~A170 & \new_[52378]_ ;
  assign \new_[52383]_  = A200 & A199;
  assign \new_[52384]_  = ~A166 & \new_[52383]_ ;
  assign \new_[52385]_  = \new_[52384]_  & \new_[52379]_ ;
  assign \new_[52389]_  = A265 & ~A233;
  assign \new_[52390]_  = ~A232 & \new_[52389]_ ;
  assign \new_[52393]_  = A298 & A266;
  assign \new_[52396]_  = ~A302 & ~A301;
  assign \new_[52397]_  = \new_[52396]_  & \new_[52393]_ ;
  assign \new_[52398]_  = \new_[52397]_  & \new_[52390]_ ;
  assign \new_[52402]_  = ~A167 & A169;
  assign \new_[52403]_  = ~A170 & \new_[52402]_ ;
  assign \new_[52407]_  = A200 & A199;
  assign \new_[52408]_  = ~A166 & \new_[52407]_ ;
  assign \new_[52409]_  = \new_[52408]_  & \new_[52403]_ ;
  assign \new_[52413]_  = ~A266 & ~A233;
  assign \new_[52414]_  = ~A232 & \new_[52413]_ ;
  assign \new_[52417]_  = ~A269 & ~A268;
  assign \new_[52420]_  = ~A300 & A298;
  assign \new_[52421]_  = \new_[52420]_  & \new_[52417]_ ;
  assign \new_[52422]_  = \new_[52421]_  & \new_[52414]_ ;
  assign \new_[52426]_  = ~A167 & A169;
  assign \new_[52427]_  = ~A170 & \new_[52426]_ ;
  assign \new_[52431]_  = A200 & A199;
  assign \new_[52432]_  = ~A166 & \new_[52431]_ ;
  assign \new_[52433]_  = \new_[52432]_  & \new_[52427]_ ;
  assign \new_[52437]_  = ~A266 & ~A233;
  assign \new_[52438]_  = ~A232 & \new_[52437]_ ;
  assign \new_[52441]_  = ~A269 & ~A268;
  assign \new_[52444]_  = A299 & A298;
  assign \new_[52445]_  = \new_[52444]_  & \new_[52441]_ ;
  assign \new_[52446]_  = \new_[52445]_  & \new_[52438]_ ;
  assign \new_[52450]_  = ~A167 & A169;
  assign \new_[52451]_  = ~A170 & \new_[52450]_ ;
  assign \new_[52455]_  = A200 & A199;
  assign \new_[52456]_  = ~A166 & \new_[52455]_ ;
  assign \new_[52457]_  = \new_[52456]_  & \new_[52451]_ ;
  assign \new_[52461]_  = ~A266 & ~A233;
  assign \new_[52462]_  = ~A232 & \new_[52461]_ ;
  assign \new_[52465]_  = ~A269 & ~A268;
  assign \new_[52468]_  = ~A299 & ~A298;
  assign \new_[52469]_  = \new_[52468]_  & \new_[52465]_ ;
  assign \new_[52470]_  = \new_[52469]_  & \new_[52462]_ ;
  assign \new_[52474]_  = ~A167 & A169;
  assign \new_[52475]_  = ~A170 & \new_[52474]_ ;
  assign \new_[52479]_  = A200 & A199;
  assign \new_[52480]_  = ~A166 & \new_[52479]_ ;
  assign \new_[52481]_  = \new_[52480]_  & \new_[52475]_ ;
  assign \new_[52485]_  = ~A266 & ~A233;
  assign \new_[52486]_  = ~A232 & \new_[52485]_ ;
  assign \new_[52489]_  = A298 & ~A267;
  assign \new_[52492]_  = ~A302 & ~A301;
  assign \new_[52493]_  = \new_[52492]_  & \new_[52489]_ ;
  assign \new_[52494]_  = \new_[52493]_  & \new_[52486]_ ;
  assign \new_[52498]_  = ~A167 & A169;
  assign \new_[52499]_  = ~A170 & \new_[52498]_ ;
  assign \new_[52503]_  = A200 & A199;
  assign \new_[52504]_  = ~A166 & \new_[52503]_ ;
  assign \new_[52505]_  = \new_[52504]_  & \new_[52499]_ ;
  assign \new_[52509]_  = ~A265 & ~A233;
  assign \new_[52510]_  = ~A232 & \new_[52509]_ ;
  assign \new_[52513]_  = A298 & ~A266;
  assign \new_[52516]_  = ~A302 & ~A301;
  assign \new_[52517]_  = \new_[52516]_  & \new_[52513]_ ;
  assign \new_[52518]_  = \new_[52517]_  & \new_[52510]_ ;
  assign \new_[52522]_  = ~A167 & A169;
  assign \new_[52523]_  = ~A170 & \new_[52522]_ ;
  assign \new_[52527]_  = ~A202 & ~A200;
  assign \new_[52528]_  = ~A166 & \new_[52527]_ ;
  assign \new_[52529]_  = \new_[52528]_  & \new_[52523]_ ;
  assign \new_[52533]_  = A233 & A232;
  assign \new_[52534]_  = ~A203 & \new_[52533]_ ;
  assign \new_[52537]_  = ~A267 & A265;
  assign \new_[52540]_  = ~A300 & ~A299;
  assign \new_[52541]_  = \new_[52540]_  & \new_[52537]_ ;
  assign \new_[52542]_  = \new_[52541]_  & \new_[52534]_ ;
  assign \new_[52546]_  = ~A167 & A169;
  assign \new_[52547]_  = ~A170 & \new_[52546]_ ;
  assign \new_[52551]_  = ~A202 & ~A200;
  assign \new_[52552]_  = ~A166 & \new_[52551]_ ;
  assign \new_[52553]_  = \new_[52552]_  & \new_[52547]_ ;
  assign \new_[52557]_  = A233 & A232;
  assign \new_[52558]_  = ~A203 & \new_[52557]_ ;
  assign \new_[52561]_  = ~A267 & A265;
  assign \new_[52564]_  = A299 & A298;
  assign \new_[52565]_  = \new_[52564]_  & \new_[52561]_ ;
  assign \new_[52566]_  = \new_[52565]_  & \new_[52558]_ ;
  assign \new_[52570]_  = ~A167 & A169;
  assign \new_[52571]_  = ~A170 & \new_[52570]_ ;
  assign \new_[52575]_  = ~A202 & ~A200;
  assign \new_[52576]_  = ~A166 & \new_[52575]_ ;
  assign \new_[52577]_  = \new_[52576]_  & \new_[52571]_ ;
  assign \new_[52581]_  = A233 & A232;
  assign \new_[52582]_  = ~A203 & \new_[52581]_ ;
  assign \new_[52585]_  = ~A267 & A265;
  assign \new_[52588]_  = ~A299 & ~A298;
  assign \new_[52589]_  = \new_[52588]_  & \new_[52585]_ ;
  assign \new_[52590]_  = \new_[52589]_  & \new_[52582]_ ;
  assign \new_[52594]_  = ~A167 & A169;
  assign \new_[52595]_  = ~A170 & \new_[52594]_ ;
  assign \new_[52599]_  = ~A202 & ~A200;
  assign \new_[52600]_  = ~A166 & \new_[52599]_ ;
  assign \new_[52601]_  = \new_[52600]_  & \new_[52595]_ ;
  assign \new_[52605]_  = A233 & A232;
  assign \new_[52606]_  = ~A203 & \new_[52605]_ ;
  assign \new_[52609]_  = A266 & A265;
  assign \new_[52612]_  = ~A300 & ~A299;
  assign \new_[52613]_  = \new_[52612]_  & \new_[52609]_ ;
  assign \new_[52614]_  = \new_[52613]_  & \new_[52606]_ ;
  assign \new_[52618]_  = ~A167 & A169;
  assign \new_[52619]_  = ~A170 & \new_[52618]_ ;
  assign \new_[52623]_  = ~A202 & ~A200;
  assign \new_[52624]_  = ~A166 & \new_[52623]_ ;
  assign \new_[52625]_  = \new_[52624]_  & \new_[52619]_ ;
  assign \new_[52629]_  = A233 & A232;
  assign \new_[52630]_  = ~A203 & \new_[52629]_ ;
  assign \new_[52633]_  = A266 & A265;
  assign \new_[52636]_  = A299 & A298;
  assign \new_[52637]_  = \new_[52636]_  & \new_[52633]_ ;
  assign \new_[52638]_  = \new_[52637]_  & \new_[52630]_ ;
  assign \new_[52642]_  = ~A167 & A169;
  assign \new_[52643]_  = ~A170 & \new_[52642]_ ;
  assign \new_[52647]_  = ~A202 & ~A200;
  assign \new_[52648]_  = ~A166 & \new_[52647]_ ;
  assign \new_[52649]_  = \new_[52648]_  & \new_[52643]_ ;
  assign \new_[52653]_  = A233 & A232;
  assign \new_[52654]_  = ~A203 & \new_[52653]_ ;
  assign \new_[52657]_  = A266 & A265;
  assign \new_[52660]_  = ~A299 & ~A298;
  assign \new_[52661]_  = \new_[52660]_  & \new_[52657]_ ;
  assign \new_[52662]_  = \new_[52661]_  & \new_[52654]_ ;
  assign \new_[52666]_  = ~A167 & A169;
  assign \new_[52667]_  = ~A170 & \new_[52666]_ ;
  assign \new_[52671]_  = ~A202 & ~A200;
  assign \new_[52672]_  = ~A166 & \new_[52671]_ ;
  assign \new_[52673]_  = \new_[52672]_  & \new_[52667]_ ;
  assign \new_[52677]_  = A233 & A232;
  assign \new_[52678]_  = ~A203 & \new_[52677]_ ;
  assign \new_[52681]_  = ~A266 & ~A265;
  assign \new_[52684]_  = ~A300 & ~A299;
  assign \new_[52685]_  = \new_[52684]_  & \new_[52681]_ ;
  assign \new_[52686]_  = \new_[52685]_  & \new_[52678]_ ;
  assign \new_[52690]_  = ~A167 & A169;
  assign \new_[52691]_  = ~A170 & \new_[52690]_ ;
  assign \new_[52695]_  = ~A202 & ~A200;
  assign \new_[52696]_  = ~A166 & \new_[52695]_ ;
  assign \new_[52697]_  = \new_[52696]_  & \new_[52691]_ ;
  assign \new_[52701]_  = A233 & A232;
  assign \new_[52702]_  = ~A203 & \new_[52701]_ ;
  assign \new_[52705]_  = ~A266 & ~A265;
  assign \new_[52708]_  = A299 & A298;
  assign \new_[52709]_  = \new_[52708]_  & \new_[52705]_ ;
  assign \new_[52710]_  = \new_[52709]_  & \new_[52702]_ ;
  assign \new_[52714]_  = ~A167 & A169;
  assign \new_[52715]_  = ~A170 & \new_[52714]_ ;
  assign \new_[52719]_  = ~A202 & ~A200;
  assign \new_[52720]_  = ~A166 & \new_[52719]_ ;
  assign \new_[52721]_  = \new_[52720]_  & \new_[52715]_ ;
  assign \new_[52725]_  = A233 & A232;
  assign \new_[52726]_  = ~A203 & \new_[52725]_ ;
  assign \new_[52729]_  = ~A266 & ~A265;
  assign \new_[52732]_  = ~A299 & ~A298;
  assign \new_[52733]_  = \new_[52732]_  & \new_[52729]_ ;
  assign \new_[52734]_  = \new_[52733]_  & \new_[52726]_ ;
  assign \new_[52738]_  = ~A167 & A169;
  assign \new_[52739]_  = ~A170 & \new_[52738]_ ;
  assign \new_[52743]_  = ~A202 & ~A200;
  assign \new_[52744]_  = ~A166 & \new_[52743]_ ;
  assign \new_[52745]_  = \new_[52744]_  & \new_[52739]_ ;
  assign \new_[52749]_  = A233 & ~A232;
  assign \new_[52750]_  = ~A203 & \new_[52749]_ ;
  assign \new_[52753]_  = ~A299 & A298;
  assign \new_[52756]_  = A301 & A300;
  assign \new_[52757]_  = \new_[52756]_  & \new_[52753]_ ;
  assign \new_[52758]_  = \new_[52757]_  & \new_[52750]_ ;
  assign \new_[52762]_  = ~A167 & A169;
  assign \new_[52763]_  = ~A170 & \new_[52762]_ ;
  assign \new_[52767]_  = ~A202 & ~A200;
  assign \new_[52768]_  = ~A166 & \new_[52767]_ ;
  assign \new_[52769]_  = \new_[52768]_  & \new_[52763]_ ;
  assign \new_[52773]_  = A233 & ~A232;
  assign \new_[52774]_  = ~A203 & \new_[52773]_ ;
  assign \new_[52777]_  = ~A299 & A298;
  assign \new_[52780]_  = A302 & A300;
  assign \new_[52781]_  = \new_[52780]_  & \new_[52777]_ ;
  assign \new_[52782]_  = \new_[52781]_  & \new_[52774]_ ;
  assign \new_[52786]_  = ~A167 & A169;
  assign \new_[52787]_  = ~A170 & \new_[52786]_ ;
  assign \new_[52791]_  = ~A202 & ~A200;
  assign \new_[52792]_  = ~A166 & \new_[52791]_ ;
  assign \new_[52793]_  = \new_[52792]_  & \new_[52787]_ ;
  assign \new_[52797]_  = A233 & ~A232;
  assign \new_[52798]_  = ~A203 & \new_[52797]_ ;
  assign \new_[52801]_  = ~A266 & A265;
  assign \new_[52804]_  = A268 & A267;
  assign \new_[52805]_  = \new_[52804]_  & \new_[52801]_ ;
  assign \new_[52806]_  = \new_[52805]_  & \new_[52798]_ ;
  assign \new_[52810]_  = ~A167 & A169;
  assign \new_[52811]_  = ~A170 & \new_[52810]_ ;
  assign \new_[52815]_  = ~A202 & ~A200;
  assign \new_[52816]_  = ~A166 & \new_[52815]_ ;
  assign \new_[52817]_  = \new_[52816]_  & \new_[52811]_ ;
  assign \new_[52821]_  = A233 & ~A232;
  assign \new_[52822]_  = ~A203 & \new_[52821]_ ;
  assign \new_[52825]_  = ~A266 & A265;
  assign \new_[52828]_  = A269 & A267;
  assign \new_[52829]_  = \new_[52828]_  & \new_[52825]_ ;
  assign \new_[52830]_  = \new_[52829]_  & \new_[52822]_ ;
  assign \new_[52834]_  = ~A167 & A169;
  assign \new_[52835]_  = ~A170 & \new_[52834]_ ;
  assign \new_[52839]_  = ~A202 & ~A200;
  assign \new_[52840]_  = ~A166 & \new_[52839]_ ;
  assign \new_[52841]_  = \new_[52840]_  & \new_[52835]_ ;
  assign \new_[52845]_  = ~A234 & ~A233;
  assign \new_[52846]_  = ~A203 & \new_[52845]_ ;
  assign \new_[52849]_  = A266 & A265;
  assign \new_[52852]_  = ~A300 & A298;
  assign \new_[52853]_  = \new_[52852]_  & \new_[52849]_ ;
  assign \new_[52854]_  = \new_[52853]_  & \new_[52846]_ ;
  assign \new_[52858]_  = ~A167 & A169;
  assign \new_[52859]_  = ~A170 & \new_[52858]_ ;
  assign \new_[52863]_  = ~A202 & ~A200;
  assign \new_[52864]_  = ~A166 & \new_[52863]_ ;
  assign \new_[52865]_  = \new_[52864]_  & \new_[52859]_ ;
  assign \new_[52869]_  = ~A234 & ~A233;
  assign \new_[52870]_  = ~A203 & \new_[52869]_ ;
  assign \new_[52873]_  = A266 & A265;
  assign \new_[52876]_  = A299 & A298;
  assign \new_[52877]_  = \new_[52876]_  & \new_[52873]_ ;
  assign \new_[52878]_  = \new_[52877]_  & \new_[52870]_ ;
  assign \new_[52882]_  = ~A167 & A169;
  assign \new_[52883]_  = ~A170 & \new_[52882]_ ;
  assign \new_[52887]_  = ~A202 & ~A200;
  assign \new_[52888]_  = ~A166 & \new_[52887]_ ;
  assign \new_[52889]_  = \new_[52888]_  & \new_[52883]_ ;
  assign \new_[52893]_  = ~A234 & ~A233;
  assign \new_[52894]_  = ~A203 & \new_[52893]_ ;
  assign \new_[52897]_  = A266 & A265;
  assign \new_[52900]_  = ~A299 & ~A298;
  assign \new_[52901]_  = \new_[52900]_  & \new_[52897]_ ;
  assign \new_[52902]_  = \new_[52901]_  & \new_[52894]_ ;
  assign \new_[52906]_  = ~A167 & A169;
  assign \new_[52907]_  = ~A170 & \new_[52906]_ ;
  assign \new_[52911]_  = ~A202 & ~A200;
  assign \new_[52912]_  = ~A166 & \new_[52911]_ ;
  assign \new_[52913]_  = \new_[52912]_  & \new_[52907]_ ;
  assign \new_[52917]_  = ~A234 & ~A233;
  assign \new_[52918]_  = ~A203 & \new_[52917]_ ;
  assign \new_[52921]_  = ~A267 & ~A266;
  assign \new_[52924]_  = ~A300 & A298;
  assign \new_[52925]_  = \new_[52924]_  & \new_[52921]_ ;
  assign \new_[52926]_  = \new_[52925]_  & \new_[52918]_ ;
  assign \new_[52930]_  = ~A167 & A169;
  assign \new_[52931]_  = ~A170 & \new_[52930]_ ;
  assign \new_[52935]_  = ~A202 & ~A200;
  assign \new_[52936]_  = ~A166 & \new_[52935]_ ;
  assign \new_[52937]_  = \new_[52936]_  & \new_[52931]_ ;
  assign \new_[52941]_  = ~A234 & ~A233;
  assign \new_[52942]_  = ~A203 & \new_[52941]_ ;
  assign \new_[52945]_  = ~A267 & ~A266;
  assign \new_[52948]_  = A299 & A298;
  assign \new_[52949]_  = \new_[52948]_  & \new_[52945]_ ;
  assign \new_[52950]_  = \new_[52949]_  & \new_[52942]_ ;
  assign \new_[52954]_  = ~A167 & A169;
  assign \new_[52955]_  = ~A170 & \new_[52954]_ ;
  assign \new_[52959]_  = ~A202 & ~A200;
  assign \new_[52960]_  = ~A166 & \new_[52959]_ ;
  assign \new_[52961]_  = \new_[52960]_  & \new_[52955]_ ;
  assign \new_[52965]_  = ~A234 & ~A233;
  assign \new_[52966]_  = ~A203 & \new_[52965]_ ;
  assign \new_[52969]_  = ~A267 & ~A266;
  assign \new_[52972]_  = ~A299 & ~A298;
  assign \new_[52973]_  = \new_[52972]_  & \new_[52969]_ ;
  assign \new_[52974]_  = \new_[52973]_  & \new_[52966]_ ;
  assign \new_[52978]_  = ~A167 & A169;
  assign \new_[52979]_  = ~A170 & \new_[52978]_ ;
  assign \new_[52983]_  = ~A202 & ~A200;
  assign \new_[52984]_  = ~A166 & \new_[52983]_ ;
  assign \new_[52985]_  = \new_[52984]_  & \new_[52979]_ ;
  assign \new_[52989]_  = ~A234 & ~A233;
  assign \new_[52990]_  = ~A203 & \new_[52989]_ ;
  assign \new_[52993]_  = ~A266 & ~A265;
  assign \new_[52996]_  = ~A300 & A298;
  assign \new_[52997]_  = \new_[52996]_  & \new_[52993]_ ;
  assign \new_[52998]_  = \new_[52997]_  & \new_[52990]_ ;
  assign \new_[53002]_  = ~A167 & A169;
  assign \new_[53003]_  = ~A170 & \new_[53002]_ ;
  assign \new_[53007]_  = ~A202 & ~A200;
  assign \new_[53008]_  = ~A166 & \new_[53007]_ ;
  assign \new_[53009]_  = \new_[53008]_  & \new_[53003]_ ;
  assign \new_[53013]_  = ~A234 & ~A233;
  assign \new_[53014]_  = ~A203 & \new_[53013]_ ;
  assign \new_[53017]_  = ~A266 & ~A265;
  assign \new_[53020]_  = A299 & A298;
  assign \new_[53021]_  = \new_[53020]_  & \new_[53017]_ ;
  assign \new_[53022]_  = \new_[53021]_  & \new_[53014]_ ;
  assign \new_[53026]_  = ~A167 & A169;
  assign \new_[53027]_  = ~A170 & \new_[53026]_ ;
  assign \new_[53031]_  = ~A202 & ~A200;
  assign \new_[53032]_  = ~A166 & \new_[53031]_ ;
  assign \new_[53033]_  = \new_[53032]_  & \new_[53027]_ ;
  assign \new_[53037]_  = ~A234 & ~A233;
  assign \new_[53038]_  = ~A203 & \new_[53037]_ ;
  assign \new_[53041]_  = ~A266 & ~A265;
  assign \new_[53044]_  = ~A299 & ~A298;
  assign \new_[53045]_  = \new_[53044]_  & \new_[53041]_ ;
  assign \new_[53046]_  = \new_[53045]_  & \new_[53038]_ ;
  assign \new_[53050]_  = ~A167 & A169;
  assign \new_[53051]_  = ~A170 & \new_[53050]_ ;
  assign \new_[53055]_  = ~A202 & ~A200;
  assign \new_[53056]_  = ~A166 & \new_[53055]_ ;
  assign \new_[53057]_  = \new_[53056]_  & \new_[53051]_ ;
  assign \new_[53061]_  = ~A233 & A232;
  assign \new_[53062]_  = ~A203 & \new_[53061]_ ;
  assign \new_[53065]_  = A235 & A234;
  assign \new_[53068]_  = A299 & ~A298;
  assign \new_[53069]_  = \new_[53068]_  & \new_[53065]_ ;
  assign \new_[53070]_  = \new_[53069]_  & \new_[53062]_ ;
  assign \new_[53074]_  = ~A167 & A169;
  assign \new_[53075]_  = ~A170 & \new_[53074]_ ;
  assign \new_[53079]_  = ~A202 & ~A200;
  assign \new_[53080]_  = ~A166 & \new_[53079]_ ;
  assign \new_[53081]_  = \new_[53080]_  & \new_[53075]_ ;
  assign \new_[53085]_  = ~A233 & A232;
  assign \new_[53086]_  = ~A203 & \new_[53085]_ ;
  assign \new_[53089]_  = A235 & A234;
  assign \new_[53092]_  = A266 & ~A265;
  assign \new_[53093]_  = \new_[53092]_  & \new_[53089]_ ;
  assign \new_[53094]_  = \new_[53093]_  & \new_[53086]_ ;
  assign \new_[53098]_  = ~A167 & A169;
  assign \new_[53099]_  = ~A170 & \new_[53098]_ ;
  assign \new_[53103]_  = ~A202 & ~A200;
  assign \new_[53104]_  = ~A166 & \new_[53103]_ ;
  assign \new_[53105]_  = \new_[53104]_  & \new_[53099]_ ;
  assign \new_[53109]_  = ~A233 & A232;
  assign \new_[53110]_  = ~A203 & \new_[53109]_ ;
  assign \new_[53113]_  = A236 & A234;
  assign \new_[53116]_  = A299 & ~A298;
  assign \new_[53117]_  = \new_[53116]_  & \new_[53113]_ ;
  assign \new_[53118]_  = \new_[53117]_  & \new_[53110]_ ;
  assign \new_[53122]_  = ~A167 & A169;
  assign \new_[53123]_  = ~A170 & \new_[53122]_ ;
  assign \new_[53127]_  = ~A202 & ~A200;
  assign \new_[53128]_  = ~A166 & \new_[53127]_ ;
  assign \new_[53129]_  = \new_[53128]_  & \new_[53123]_ ;
  assign \new_[53133]_  = ~A233 & A232;
  assign \new_[53134]_  = ~A203 & \new_[53133]_ ;
  assign \new_[53137]_  = A236 & A234;
  assign \new_[53140]_  = A266 & ~A265;
  assign \new_[53141]_  = \new_[53140]_  & \new_[53137]_ ;
  assign \new_[53142]_  = \new_[53141]_  & \new_[53134]_ ;
  assign \new_[53146]_  = ~A167 & A169;
  assign \new_[53147]_  = ~A170 & \new_[53146]_ ;
  assign \new_[53151]_  = ~A202 & ~A200;
  assign \new_[53152]_  = ~A166 & \new_[53151]_ ;
  assign \new_[53153]_  = \new_[53152]_  & \new_[53147]_ ;
  assign \new_[53157]_  = ~A233 & ~A232;
  assign \new_[53158]_  = ~A203 & \new_[53157]_ ;
  assign \new_[53161]_  = A266 & A265;
  assign \new_[53164]_  = ~A300 & A298;
  assign \new_[53165]_  = \new_[53164]_  & \new_[53161]_ ;
  assign \new_[53166]_  = \new_[53165]_  & \new_[53158]_ ;
  assign \new_[53170]_  = ~A167 & A169;
  assign \new_[53171]_  = ~A170 & \new_[53170]_ ;
  assign \new_[53175]_  = ~A202 & ~A200;
  assign \new_[53176]_  = ~A166 & \new_[53175]_ ;
  assign \new_[53177]_  = \new_[53176]_  & \new_[53171]_ ;
  assign \new_[53181]_  = ~A233 & ~A232;
  assign \new_[53182]_  = ~A203 & \new_[53181]_ ;
  assign \new_[53185]_  = A266 & A265;
  assign \new_[53188]_  = A299 & A298;
  assign \new_[53189]_  = \new_[53188]_  & \new_[53185]_ ;
  assign \new_[53190]_  = \new_[53189]_  & \new_[53182]_ ;
  assign \new_[53194]_  = ~A167 & A169;
  assign \new_[53195]_  = ~A170 & \new_[53194]_ ;
  assign \new_[53199]_  = ~A202 & ~A200;
  assign \new_[53200]_  = ~A166 & \new_[53199]_ ;
  assign \new_[53201]_  = \new_[53200]_  & \new_[53195]_ ;
  assign \new_[53205]_  = ~A233 & ~A232;
  assign \new_[53206]_  = ~A203 & \new_[53205]_ ;
  assign \new_[53209]_  = A266 & A265;
  assign \new_[53212]_  = ~A299 & ~A298;
  assign \new_[53213]_  = \new_[53212]_  & \new_[53209]_ ;
  assign \new_[53214]_  = \new_[53213]_  & \new_[53206]_ ;
  assign \new_[53218]_  = ~A167 & A169;
  assign \new_[53219]_  = ~A170 & \new_[53218]_ ;
  assign \new_[53223]_  = ~A202 & ~A200;
  assign \new_[53224]_  = ~A166 & \new_[53223]_ ;
  assign \new_[53225]_  = \new_[53224]_  & \new_[53219]_ ;
  assign \new_[53229]_  = ~A233 & ~A232;
  assign \new_[53230]_  = ~A203 & \new_[53229]_ ;
  assign \new_[53233]_  = ~A267 & ~A266;
  assign \new_[53236]_  = ~A300 & A298;
  assign \new_[53237]_  = \new_[53236]_  & \new_[53233]_ ;
  assign \new_[53238]_  = \new_[53237]_  & \new_[53230]_ ;
  assign \new_[53242]_  = ~A167 & A169;
  assign \new_[53243]_  = ~A170 & \new_[53242]_ ;
  assign \new_[53247]_  = ~A202 & ~A200;
  assign \new_[53248]_  = ~A166 & \new_[53247]_ ;
  assign \new_[53249]_  = \new_[53248]_  & \new_[53243]_ ;
  assign \new_[53253]_  = ~A233 & ~A232;
  assign \new_[53254]_  = ~A203 & \new_[53253]_ ;
  assign \new_[53257]_  = ~A267 & ~A266;
  assign \new_[53260]_  = A299 & A298;
  assign \new_[53261]_  = \new_[53260]_  & \new_[53257]_ ;
  assign \new_[53262]_  = \new_[53261]_  & \new_[53254]_ ;
  assign \new_[53266]_  = ~A167 & A169;
  assign \new_[53267]_  = ~A170 & \new_[53266]_ ;
  assign \new_[53271]_  = ~A202 & ~A200;
  assign \new_[53272]_  = ~A166 & \new_[53271]_ ;
  assign \new_[53273]_  = \new_[53272]_  & \new_[53267]_ ;
  assign \new_[53277]_  = ~A233 & ~A232;
  assign \new_[53278]_  = ~A203 & \new_[53277]_ ;
  assign \new_[53281]_  = ~A267 & ~A266;
  assign \new_[53284]_  = ~A299 & ~A298;
  assign \new_[53285]_  = \new_[53284]_  & \new_[53281]_ ;
  assign \new_[53286]_  = \new_[53285]_  & \new_[53278]_ ;
  assign \new_[53290]_  = ~A167 & A169;
  assign \new_[53291]_  = ~A170 & \new_[53290]_ ;
  assign \new_[53295]_  = ~A202 & ~A200;
  assign \new_[53296]_  = ~A166 & \new_[53295]_ ;
  assign \new_[53297]_  = \new_[53296]_  & \new_[53291]_ ;
  assign \new_[53301]_  = ~A233 & ~A232;
  assign \new_[53302]_  = ~A203 & \new_[53301]_ ;
  assign \new_[53305]_  = ~A266 & ~A265;
  assign \new_[53308]_  = ~A300 & A298;
  assign \new_[53309]_  = \new_[53308]_  & \new_[53305]_ ;
  assign \new_[53310]_  = \new_[53309]_  & \new_[53302]_ ;
  assign \new_[53314]_  = ~A167 & A169;
  assign \new_[53315]_  = ~A170 & \new_[53314]_ ;
  assign \new_[53319]_  = ~A202 & ~A200;
  assign \new_[53320]_  = ~A166 & \new_[53319]_ ;
  assign \new_[53321]_  = \new_[53320]_  & \new_[53315]_ ;
  assign \new_[53325]_  = ~A233 & ~A232;
  assign \new_[53326]_  = ~A203 & \new_[53325]_ ;
  assign \new_[53329]_  = ~A266 & ~A265;
  assign \new_[53332]_  = A299 & A298;
  assign \new_[53333]_  = \new_[53332]_  & \new_[53329]_ ;
  assign \new_[53334]_  = \new_[53333]_  & \new_[53326]_ ;
  assign \new_[53338]_  = ~A167 & A169;
  assign \new_[53339]_  = ~A170 & \new_[53338]_ ;
  assign \new_[53343]_  = ~A202 & ~A200;
  assign \new_[53344]_  = ~A166 & \new_[53343]_ ;
  assign \new_[53345]_  = \new_[53344]_  & \new_[53339]_ ;
  assign \new_[53349]_  = ~A233 & ~A232;
  assign \new_[53350]_  = ~A203 & \new_[53349]_ ;
  assign \new_[53353]_  = ~A266 & ~A265;
  assign \new_[53356]_  = ~A299 & ~A298;
  assign \new_[53357]_  = \new_[53356]_  & \new_[53353]_ ;
  assign \new_[53358]_  = \new_[53357]_  & \new_[53350]_ ;
  assign \new_[53362]_  = ~A167 & A169;
  assign \new_[53363]_  = ~A170 & \new_[53362]_ ;
  assign \new_[53367]_  = ~A201 & ~A200;
  assign \new_[53368]_  = ~A166 & \new_[53367]_ ;
  assign \new_[53369]_  = \new_[53368]_  & \new_[53363]_ ;
  assign \new_[53373]_  = A265 & A233;
  assign \new_[53374]_  = A232 & \new_[53373]_ ;
  assign \new_[53377]_  = ~A269 & ~A268;
  assign \new_[53380]_  = ~A300 & ~A299;
  assign \new_[53381]_  = \new_[53380]_  & \new_[53377]_ ;
  assign \new_[53382]_  = \new_[53381]_  & \new_[53374]_ ;
  assign \new_[53386]_  = ~A167 & A169;
  assign \new_[53387]_  = ~A170 & \new_[53386]_ ;
  assign \new_[53391]_  = ~A201 & ~A200;
  assign \new_[53392]_  = ~A166 & \new_[53391]_ ;
  assign \new_[53393]_  = \new_[53392]_  & \new_[53387]_ ;
  assign \new_[53397]_  = A265 & A233;
  assign \new_[53398]_  = A232 & \new_[53397]_ ;
  assign \new_[53401]_  = ~A269 & ~A268;
  assign \new_[53404]_  = A299 & A298;
  assign \new_[53405]_  = \new_[53404]_  & \new_[53401]_ ;
  assign \new_[53406]_  = \new_[53405]_  & \new_[53398]_ ;
  assign \new_[53410]_  = ~A167 & A169;
  assign \new_[53411]_  = ~A170 & \new_[53410]_ ;
  assign \new_[53415]_  = ~A201 & ~A200;
  assign \new_[53416]_  = ~A166 & \new_[53415]_ ;
  assign \new_[53417]_  = \new_[53416]_  & \new_[53411]_ ;
  assign \new_[53421]_  = A265 & A233;
  assign \new_[53422]_  = A232 & \new_[53421]_ ;
  assign \new_[53425]_  = ~A269 & ~A268;
  assign \new_[53428]_  = ~A299 & ~A298;
  assign \new_[53429]_  = \new_[53428]_  & \new_[53425]_ ;
  assign \new_[53430]_  = \new_[53429]_  & \new_[53422]_ ;
  assign \new_[53434]_  = ~A167 & A169;
  assign \new_[53435]_  = ~A170 & \new_[53434]_ ;
  assign \new_[53439]_  = ~A201 & ~A200;
  assign \new_[53440]_  = ~A166 & \new_[53439]_ ;
  assign \new_[53441]_  = \new_[53440]_  & \new_[53435]_ ;
  assign \new_[53445]_  = A265 & A233;
  assign \new_[53446]_  = A232 & \new_[53445]_ ;
  assign \new_[53449]_  = ~A299 & ~A267;
  assign \new_[53452]_  = ~A302 & ~A301;
  assign \new_[53453]_  = \new_[53452]_  & \new_[53449]_ ;
  assign \new_[53454]_  = \new_[53453]_  & \new_[53446]_ ;
  assign \new_[53458]_  = ~A167 & A169;
  assign \new_[53459]_  = ~A170 & \new_[53458]_ ;
  assign \new_[53463]_  = ~A201 & ~A200;
  assign \new_[53464]_  = ~A166 & \new_[53463]_ ;
  assign \new_[53465]_  = \new_[53464]_  & \new_[53459]_ ;
  assign \new_[53469]_  = A265 & A233;
  assign \new_[53470]_  = A232 & \new_[53469]_ ;
  assign \new_[53473]_  = ~A299 & A266;
  assign \new_[53476]_  = ~A302 & ~A301;
  assign \new_[53477]_  = \new_[53476]_  & \new_[53473]_ ;
  assign \new_[53478]_  = \new_[53477]_  & \new_[53470]_ ;
  assign \new_[53482]_  = ~A167 & A169;
  assign \new_[53483]_  = ~A170 & \new_[53482]_ ;
  assign \new_[53487]_  = ~A201 & ~A200;
  assign \new_[53488]_  = ~A166 & \new_[53487]_ ;
  assign \new_[53489]_  = \new_[53488]_  & \new_[53483]_ ;
  assign \new_[53493]_  = ~A265 & A233;
  assign \new_[53494]_  = A232 & \new_[53493]_ ;
  assign \new_[53497]_  = ~A299 & ~A266;
  assign \new_[53500]_  = ~A302 & ~A301;
  assign \new_[53501]_  = \new_[53500]_  & \new_[53497]_ ;
  assign \new_[53502]_  = \new_[53501]_  & \new_[53494]_ ;
  assign \new_[53506]_  = ~A167 & A169;
  assign \new_[53507]_  = ~A170 & \new_[53506]_ ;
  assign \new_[53511]_  = ~A201 & ~A200;
  assign \new_[53512]_  = ~A166 & \new_[53511]_ ;
  assign \new_[53513]_  = \new_[53512]_  & \new_[53507]_ ;
  assign \new_[53517]_  = ~A236 & ~A235;
  assign \new_[53518]_  = ~A233 & \new_[53517]_ ;
  assign \new_[53521]_  = A266 & A265;
  assign \new_[53524]_  = ~A300 & A298;
  assign \new_[53525]_  = \new_[53524]_  & \new_[53521]_ ;
  assign \new_[53526]_  = \new_[53525]_  & \new_[53518]_ ;
  assign \new_[53530]_  = ~A167 & A169;
  assign \new_[53531]_  = ~A170 & \new_[53530]_ ;
  assign \new_[53535]_  = ~A201 & ~A200;
  assign \new_[53536]_  = ~A166 & \new_[53535]_ ;
  assign \new_[53537]_  = \new_[53536]_  & \new_[53531]_ ;
  assign \new_[53541]_  = ~A236 & ~A235;
  assign \new_[53542]_  = ~A233 & \new_[53541]_ ;
  assign \new_[53545]_  = A266 & A265;
  assign \new_[53548]_  = A299 & A298;
  assign \new_[53549]_  = \new_[53548]_  & \new_[53545]_ ;
  assign \new_[53550]_  = \new_[53549]_  & \new_[53542]_ ;
  assign \new_[53554]_  = ~A167 & A169;
  assign \new_[53555]_  = ~A170 & \new_[53554]_ ;
  assign \new_[53559]_  = ~A201 & ~A200;
  assign \new_[53560]_  = ~A166 & \new_[53559]_ ;
  assign \new_[53561]_  = \new_[53560]_  & \new_[53555]_ ;
  assign \new_[53565]_  = ~A236 & ~A235;
  assign \new_[53566]_  = ~A233 & \new_[53565]_ ;
  assign \new_[53569]_  = A266 & A265;
  assign \new_[53572]_  = ~A299 & ~A298;
  assign \new_[53573]_  = \new_[53572]_  & \new_[53569]_ ;
  assign \new_[53574]_  = \new_[53573]_  & \new_[53566]_ ;
  assign \new_[53578]_  = ~A167 & A169;
  assign \new_[53579]_  = ~A170 & \new_[53578]_ ;
  assign \new_[53583]_  = ~A201 & ~A200;
  assign \new_[53584]_  = ~A166 & \new_[53583]_ ;
  assign \new_[53585]_  = \new_[53584]_  & \new_[53579]_ ;
  assign \new_[53589]_  = ~A236 & ~A235;
  assign \new_[53590]_  = ~A233 & \new_[53589]_ ;
  assign \new_[53593]_  = ~A267 & ~A266;
  assign \new_[53596]_  = ~A300 & A298;
  assign \new_[53597]_  = \new_[53596]_  & \new_[53593]_ ;
  assign \new_[53598]_  = \new_[53597]_  & \new_[53590]_ ;
  assign \new_[53602]_  = ~A167 & A169;
  assign \new_[53603]_  = ~A170 & \new_[53602]_ ;
  assign \new_[53607]_  = ~A201 & ~A200;
  assign \new_[53608]_  = ~A166 & \new_[53607]_ ;
  assign \new_[53609]_  = \new_[53608]_  & \new_[53603]_ ;
  assign \new_[53613]_  = ~A236 & ~A235;
  assign \new_[53614]_  = ~A233 & \new_[53613]_ ;
  assign \new_[53617]_  = ~A267 & ~A266;
  assign \new_[53620]_  = A299 & A298;
  assign \new_[53621]_  = \new_[53620]_  & \new_[53617]_ ;
  assign \new_[53622]_  = \new_[53621]_  & \new_[53614]_ ;
  assign \new_[53626]_  = ~A167 & A169;
  assign \new_[53627]_  = ~A170 & \new_[53626]_ ;
  assign \new_[53631]_  = ~A201 & ~A200;
  assign \new_[53632]_  = ~A166 & \new_[53631]_ ;
  assign \new_[53633]_  = \new_[53632]_  & \new_[53627]_ ;
  assign \new_[53637]_  = ~A236 & ~A235;
  assign \new_[53638]_  = ~A233 & \new_[53637]_ ;
  assign \new_[53641]_  = ~A267 & ~A266;
  assign \new_[53644]_  = ~A299 & ~A298;
  assign \new_[53645]_  = \new_[53644]_  & \new_[53641]_ ;
  assign \new_[53646]_  = \new_[53645]_  & \new_[53638]_ ;
  assign \new_[53650]_  = ~A167 & A169;
  assign \new_[53651]_  = ~A170 & \new_[53650]_ ;
  assign \new_[53655]_  = ~A201 & ~A200;
  assign \new_[53656]_  = ~A166 & \new_[53655]_ ;
  assign \new_[53657]_  = \new_[53656]_  & \new_[53651]_ ;
  assign \new_[53661]_  = ~A236 & ~A235;
  assign \new_[53662]_  = ~A233 & \new_[53661]_ ;
  assign \new_[53665]_  = ~A266 & ~A265;
  assign \new_[53668]_  = ~A300 & A298;
  assign \new_[53669]_  = \new_[53668]_  & \new_[53665]_ ;
  assign \new_[53670]_  = \new_[53669]_  & \new_[53662]_ ;
  assign \new_[53674]_  = ~A167 & A169;
  assign \new_[53675]_  = ~A170 & \new_[53674]_ ;
  assign \new_[53679]_  = ~A201 & ~A200;
  assign \new_[53680]_  = ~A166 & \new_[53679]_ ;
  assign \new_[53681]_  = \new_[53680]_  & \new_[53675]_ ;
  assign \new_[53685]_  = ~A236 & ~A235;
  assign \new_[53686]_  = ~A233 & \new_[53685]_ ;
  assign \new_[53689]_  = ~A266 & ~A265;
  assign \new_[53692]_  = A299 & A298;
  assign \new_[53693]_  = \new_[53692]_  & \new_[53689]_ ;
  assign \new_[53694]_  = \new_[53693]_  & \new_[53686]_ ;
  assign \new_[53698]_  = ~A167 & A169;
  assign \new_[53699]_  = ~A170 & \new_[53698]_ ;
  assign \new_[53703]_  = ~A201 & ~A200;
  assign \new_[53704]_  = ~A166 & \new_[53703]_ ;
  assign \new_[53705]_  = \new_[53704]_  & \new_[53699]_ ;
  assign \new_[53709]_  = ~A236 & ~A235;
  assign \new_[53710]_  = ~A233 & \new_[53709]_ ;
  assign \new_[53713]_  = ~A266 & ~A265;
  assign \new_[53716]_  = ~A299 & ~A298;
  assign \new_[53717]_  = \new_[53716]_  & \new_[53713]_ ;
  assign \new_[53718]_  = \new_[53717]_  & \new_[53710]_ ;
  assign \new_[53722]_  = ~A167 & A169;
  assign \new_[53723]_  = ~A170 & \new_[53722]_ ;
  assign \new_[53727]_  = ~A201 & ~A200;
  assign \new_[53728]_  = ~A166 & \new_[53727]_ ;
  assign \new_[53729]_  = \new_[53728]_  & \new_[53723]_ ;
  assign \new_[53733]_  = A265 & ~A234;
  assign \new_[53734]_  = ~A233 & \new_[53733]_ ;
  assign \new_[53737]_  = A298 & A266;
  assign \new_[53740]_  = ~A302 & ~A301;
  assign \new_[53741]_  = \new_[53740]_  & \new_[53737]_ ;
  assign \new_[53742]_  = \new_[53741]_  & \new_[53734]_ ;
  assign \new_[53746]_  = ~A167 & A169;
  assign \new_[53747]_  = ~A170 & \new_[53746]_ ;
  assign \new_[53751]_  = ~A201 & ~A200;
  assign \new_[53752]_  = ~A166 & \new_[53751]_ ;
  assign \new_[53753]_  = \new_[53752]_  & \new_[53747]_ ;
  assign \new_[53757]_  = ~A266 & ~A234;
  assign \new_[53758]_  = ~A233 & \new_[53757]_ ;
  assign \new_[53761]_  = ~A269 & ~A268;
  assign \new_[53764]_  = ~A300 & A298;
  assign \new_[53765]_  = \new_[53764]_  & \new_[53761]_ ;
  assign \new_[53766]_  = \new_[53765]_  & \new_[53758]_ ;
  assign \new_[53770]_  = ~A167 & A169;
  assign \new_[53771]_  = ~A170 & \new_[53770]_ ;
  assign \new_[53775]_  = ~A201 & ~A200;
  assign \new_[53776]_  = ~A166 & \new_[53775]_ ;
  assign \new_[53777]_  = \new_[53776]_  & \new_[53771]_ ;
  assign \new_[53781]_  = ~A266 & ~A234;
  assign \new_[53782]_  = ~A233 & \new_[53781]_ ;
  assign \new_[53785]_  = ~A269 & ~A268;
  assign \new_[53788]_  = A299 & A298;
  assign \new_[53789]_  = \new_[53788]_  & \new_[53785]_ ;
  assign \new_[53790]_  = \new_[53789]_  & \new_[53782]_ ;
  assign \new_[53794]_  = ~A167 & A169;
  assign \new_[53795]_  = ~A170 & \new_[53794]_ ;
  assign \new_[53799]_  = ~A201 & ~A200;
  assign \new_[53800]_  = ~A166 & \new_[53799]_ ;
  assign \new_[53801]_  = \new_[53800]_  & \new_[53795]_ ;
  assign \new_[53805]_  = ~A266 & ~A234;
  assign \new_[53806]_  = ~A233 & \new_[53805]_ ;
  assign \new_[53809]_  = ~A269 & ~A268;
  assign \new_[53812]_  = ~A299 & ~A298;
  assign \new_[53813]_  = \new_[53812]_  & \new_[53809]_ ;
  assign \new_[53814]_  = \new_[53813]_  & \new_[53806]_ ;
  assign \new_[53818]_  = ~A167 & A169;
  assign \new_[53819]_  = ~A170 & \new_[53818]_ ;
  assign \new_[53823]_  = ~A201 & ~A200;
  assign \new_[53824]_  = ~A166 & \new_[53823]_ ;
  assign \new_[53825]_  = \new_[53824]_  & \new_[53819]_ ;
  assign \new_[53829]_  = ~A266 & ~A234;
  assign \new_[53830]_  = ~A233 & \new_[53829]_ ;
  assign \new_[53833]_  = A298 & ~A267;
  assign \new_[53836]_  = ~A302 & ~A301;
  assign \new_[53837]_  = \new_[53836]_  & \new_[53833]_ ;
  assign \new_[53838]_  = \new_[53837]_  & \new_[53830]_ ;
  assign \new_[53842]_  = ~A167 & A169;
  assign \new_[53843]_  = ~A170 & \new_[53842]_ ;
  assign \new_[53847]_  = ~A201 & ~A200;
  assign \new_[53848]_  = ~A166 & \new_[53847]_ ;
  assign \new_[53849]_  = \new_[53848]_  & \new_[53843]_ ;
  assign \new_[53853]_  = ~A265 & ~A234;
  assign \new_[53854]_  = ~A233 & \new_[53853]_ ;
  assign \new_[53857]_  = A298 & ~A266;
  assign \new_[53860]_  = ~A302 & ~A301;
  assign \new_[53861]_  = \new_[53860]_  & \new_[53857]_ ;
  assign \new_[53862]_  = \new_[53861]_  & \new_[53854]_ ;
  assign \new_[53866]_  = ~A167 & A169;
  assign \new_[53867]_  = ~A170 & \new_[53866]_ ;
  assign \new_[53871]_  = ~A201 & ~A200;
  assign \new_[53872]_  = ~A166 & \new_[53871]_ ;
  assign \new_[53873]_  = \new_[53872]_  & \new_[53867]_ ;
  assign \new_[53877]_  = A265 & ~A233;
  assign \new_[53878]_  = ~A232 & \new_[53877]_ ;
  assign \new_[53881]_  = A298 & A266;
  assign \new_[53884]_  = ~A302 & ~A301;
  assign \new_[53885]_  = \new_[53884]_  & \new_[53881]_ ;
  assign \new_[53886]_  = \new_[53885]_  & \new_[53878]_ ;
  assign \new_[53890]_  = ~A167 & A169;
  assign \new_[53891]_  = ~A170 & \new_[53890]_ ;
  assign \new_[53895]_  = ~A201 & ~A200;
  assign \new_[53896]_  = ~A166 & \new_[53895]_ ;
  assign \new_[53897]_  = \new_[53896]_  & \new_[53891]_ ;
  assign \new_[53901]_  = ~A266 & ~A233;
  assign \new_[53902]_  = ~A232 & \new_[53901]_ ;
  assign \new_[53905]_  = ~A269 & ~A268;
  assign \new_[53908]_  = ~A300 & A298;
  assign \new_[53909]_  = \new_[53908]_  & \new_[53905]_ ;
  assign \new_[53910]_  = \new_[53909]_  & \new_[53902]_ ;
  assign \new_[53914]_  = ~A167 & A169;
  assign \new_[53915]_  = ~A170 & \new_[53914]_ ;
  assign \new_[53919]_  = ~A201 & ~A200;
  assign \new_[53920]_  = ~A166 & \new_[53919]_ ;
  assign \new_[53921]_  = \new_[53920]_  & \new_[53915]_ ;
  assign \new_[53925]_  = ~A266 & ~A233;
  assign \new_[53926]_  = ~A232 & \new_[53925]_ ;
  assign \new_[53929]_  = ~A269 & ~A268;
  assign \new_[53932]_  = A299 & A298;
  assign \new_[53933]_  = \new_[53932]_  & \new_[53929]_ ;
  assign \new_[53934]_  = \new_[53933]_  & \new_[53926]_ ;
  assign \new_[53938]_  = ~A167 & A169;
  assign \new_[53939]_  = ~A170 & \new_[53938]_ ;
  assign \new_[53943]_  = ~A201 & ~A200;
  assign \new_[53944]_  = ~A166 & \new_[53943]_ ;
  assign \new_[53945]_  = \new_[53944]_  & \new_[53939]_ ;
  assign \new_[53949]_  = ~A266 & ~A233;
  assign \new_[53950]_  = ~A232 & \new_[53949]_ ;
  assign \new_[53953]_  = ~A269 & ~A268;
  assign \new_[53956]_  = ~A299 & ~A298;
  assign \new_[53957]_  = \new_[53956]_  & \new_[53953]_ ;
  assign \new_[53958]_  = \new_[53957]_  & \new_[53950]_ ;
  assign \new_[53962]_  = ~A167 & A169;
  assign \new_[53963]_  = ~A170 & \new_[53962]_ ;
  assign \new_[53967]_  = ~A201 & ~A200;
  assign \new_[53968]_  = ~A166 & \new_[53967]_ ;
  assign \new_[53969]_  = \new_[53968]_  & \new_[53963]_ ;
  assign \new_[53973]_  = ~A266 & ~A233;
  assign \new_[53974]_  = ~A232 & \new_[53973]_ ;
  assign \new_[53977]_  = A298 & ~A267;
  assign \new_[53980]_  = ~A302 & ~A301;
  assign \new_[53981]_  = \new_[53980]_  & \new_[53977]_ ;
  assign \new_[53982]_  = \new_[53981]_  & \new_[53974]_ ;
  assign \new_[53986]_  = ~A167 & A169;
  assign \new_[53987]_  = ~A170 & \new_[53986]_ ;
  assign \new_[53991]_  = ~A201 & ~A200;
  assign \new_[53992]_  = ~A166 & \new_[53991]_ ;
  assign \new_[53993]_  = \new_[53992]_  & \new_[53987]_ ;
  assign \new_[53997]_  = ~A265 & ~A233;
  assign \new_[53998]_  = ~A232 & \new_[53997]_ ;
  assign \new_[54001]_  = A298 & ~A266;
  assign \new_[54004]_  = ~A302 & ~A301;
  assign \new_[54005]_  = \new_[54004]_  & \new_[54001]_ ;
  assign \new_[54006]_  = \new_[54005]_  & \new_[53998]_ ;
  assign \new_[54010]_  = ~A167 & A169;
  assign \new_[54011]_  = ~A170 & \new_[54010]_ ;
  assign \new_[54015]_  = ~A200 & ~A199;
  assign \new_[54016]_  = ~A166 & \new_[54015]_ ;
  assign \new_[54017]_  = \new_[54016]_  & \new_[54011]_ ;
  assign \new_[54021]_  = A265 & A233;
  assign \new_[54022]_  = A232 & \new_[54021]_ ;
  assign \new_[54025]_  = ~A269 & ~A268;
  assign \new_[54028]_  = ~A300 & ~A299;
  assign \new_[54029]_  = \new_[54028]_  & \new_[54025]_ ;
  assign \new_[54030]_  = \new_[54029]_  & \new_[54022]_ ;
  assign \new_[54034]_  = ~A167 & A169;
  assign \new_[54035]_  = ~A170 & \new_[54034]_ ;
  assign \new_[54039]_  = ~A200 & ~A199;
  assign \new_[54040]_  = ~A166 & \new_[54039]_ ;
  assign \new_[54041]_  = \new_[54040]_  & \new_[54035]_ ;
  assign \new_[54045]_  = A265 & A233;
  assign \new_[54046]_  = A232 & \new_[54045]_ ;
  assign \new_[54049]_  = ~A269 & ~A268;
  assign \new_[54052]_  = A299 & A298;
  assign \new_[54053]_  = \new_[54052]_  & \new_[54049]_ ;
  assign \new_[54054]_  = \new_[54053]_  & \new_[54046]_ ;
  assign \new_[54058]_  = ~A167 & A169;
  assign \new_[54059]_  = ~A170 & \new_[54058]_ ;
  assign \new_[54063]_  = ~A200 & ~A199;
  assign \new_[54064]_  = ~A166 & \new_[54063]_ ;
  assign \new_[54065]_  = \new_[54064]_  & \new_[54059]_ ;
  assign \new_[54069]_  = A265 & A233;
  assign \new_[54070]_  = A232 & \new_[54069]_ ;
  assign \new_[54073]_  = ~A269 & ~A268;
  assign \new_[54076]_  = ~A299 & ~A298;
  assign \new_[54077]_  = \new_[54076]_  & \new_[54073]_ ;
  assign \new_[54078]_  = \new_[54077]_  & \new_[54070]_ ;
  assign \new_[54082]_  = ~A167 & A169;
  assign \new_[54083]_  = ~A170 & \new_[54082]_ ;
  assign \new_[54087]_  = ~A200 & ~A199;
  assign \new_[54088]_  = ~A166 & \new_[54087]_ ;
  assign \new_[54089]_  = \new_[54088]_  & \new_[54083]_ ;
  assign \new_[54093]_  = A265 & A233;
  assign \new_[54094]_  = A232 & \new_[54093]_ ;
  assign \new_[54097]_  = ~A299 & ~A267;
  assign \new_[54100]_  = ~A302 & ~A301;
  assign \new_[54101]_  = \new_[54100]_  & \new_[54097]_ ;
  assign \new_[54102]_  = \new_[54101]_  & \new_[54094]_ ;
  assign \new_[54106]_  = ~A167 & A169;
  assign \new_[54107]_  = ~A170 & \new_[54106]_ ;
  assign \new_[54111]_  = ~A200 & ~A199;
  assign \new_[54112]_  = ~A166 & \new_[54111]_ ;
  assign \new_[54113]_  = \new_[54112]_  & \new_[54107]_ ;
  assign \new_[54117]_  = A265 & A233;
  assign \new_[54118]_  = A232 & \new_[54117]_ ;
  assign \new_[54121]_  = ~A299 & A266;
  assign \new_[54124]_  = ~A302 & ~A301;
  assign \new_[54125]_  = \new_[54124]_  & \new_[54121]_ ;
  assign \new_[54126]_  = \new_[54125]_  & \new_[54118]_ ;
  assign \new_[54130]_  = ~A167 & A169;
  assign \new_[54131]_  = ~A170 & \new_[54130]_ ;
  assign \new_[54135]_  = ~A200 & ~A199;
  assign \new_[54136]_  = ~A166 & \new_[54135]_ ;
  assign \new_[54137]_  = \new_[54136]_  & \new_[54131]_ ;
  assign \new_[54141]_  = ~A265 & A233;
  assign \new_[54142]_  = A232 & \new_[54141]_ ;
  assign \new_[54145]_  = ~A299 & ~A266;
  assign \new_[54148]_  = ~A302 & ~A301;
  assign \new_[54149]_  = \new_[54148]_  & \new_[54145]_ ;
  assign \new_[54150]_  = \new_[54149]_  & \new_[54142]_ ;
  assign \new_[54154]_  = ~A167 & A169;
  assign \new_[54155]_  = ~A170 & \new_[54154]_ ;
  assign \new_[54159]_  = ~A200 & ~A199;
  assign \new_[54160]_  = ~A166 & \new_[54159]_ ;
  assign \new_[54161]_  = \new_[54160]_  & \new_[54155]_ ;
  assign \new_[54165]_  = ~A236 & ~A235;
  assign \new_[54166]_  = ~A233 & \new_[54165]_ ;
  assign \new_[54169]_  = A266 & A265;
  assign \new_[54172]_  = ~A300 & A298;
  assign \new_[54173]_  = \new_[54172]_  & \new_[54169]_ ;
  assign \new_[54174]_  = \new_[54173]_  & \new_[54166]_ ;
  assign \new_[54178]_  = ~A167 & A169;
  assign \new_[54179]_  = ~A170 & \new_[54178]_ ;
  assign \new_[54183]_  = ~A200 & ~A199;
  assign \new_[54184]_  = ~A166 & \new_[54183]_ ;
  assign \new_[54185]_  = \new_[54184]_  & \new_[54179]_ ;
  assign \new_[54189]_  = ~A236 & ~A235;
  assign \new_[54190]_  = ~A233 & \new_[54189]_ ;
  assign \new_[54193]_  = A266 & A265;
  assign \new_[54196]_  = A299 & A298;
  assign \new_[54197]_  = \new_[54196]_  & \new_[54193]_ ;
  assign \new_[54198]_  = \new_[54197]_  & \new_[54190]_ ;
  assign \new_[54202]_  = ~A167 & A169;
  assign \new_[54203]_  = ~A170 & \new_[54202]_ ;
  assign \new_[54207]_  = ~A200 & ~A199;
  assign \new_[54208]_  = ~A166 & \new_[54207]_ ;
  assign \new_[54209]_  = \new_[54208]_  & \new_[54203]_ ;
  assign \new_[54213]_  = ~A236 & ~A235;
  assign \new_[54214]_  = ~A233 & \new_[54213]_ ;
  assign \new_[54217]_  = A266 & A265;
  assign \new_[54220]_  = ~A299 & ~A298;
  assign \new_[54221]_  = \new_[54220]_  & \new_[54217]_ ;
  assign \new_[54222]_  = \new_[54221]_  & \new_[54214]_ ;
  assign \new_[54226]_  = ~A167 & A169;
  assign \new_[54227]_  = ~A170 & \new_[54226]_ ;
  assign \new_[54231]_  = ~A200 & ~A199;
  assign \new_[54232]_  = ~A166 & \new_[54231]_ ;
  assign \new_[54233]_  = \new_[54232]_  & \new_[54227]_ ;
  assign \new_[54237]_  = ~A236 & ~A235;
  assign \new_[54238]_  = ~A233 & \new_[54237]_ ;
  assign \new_[54241]_  = ~A267 & ~A266;
  assign \new_[54244]_  = ~A300 & A298;
  assign \new_[54245]_  = \new_[54244]_  & \new_[54241]_ ;
  assign \new_[54246]_  = \new_[54245]_  & \new_[54238]_ ;
  assign \new_[54250]_  = ~A167 & A169;
  assign \new_[54251]_  = ~A170 & \new_[54250]_ ;
  assign \new_[54255]_  = ~A200 & ~A199;
  assign \new_[54256]_  = ~A166 & \new_[54255]_ ;
  assign \new_[54257]_  = \new_[54256]_  & \new_[54251]_ ;
  assign \new_[54261]_  = ~A236 & ~A235;
  assign \new_[54262]_  = ~A233 & \new_[54261]_ ;
  assign \new_[54265]_  = ~A267 & ~A266;
  assign \new_[54268]_  = A299 & A298;
  assign \new_[54269]_  = \new_[54268]_  & \new_[54265]_ ;
  assign \new_[54270]_  = \new_[54269]_  & \new_[54262]_ ;
  assign \new_[54274]_  = ~A167 & A169;
  assign \new_[54275]_  = ~A170 & \new_[54274]_ ;
  assign \new_[54279]_  = ~A200 & ~A199;
  assign \new_[54280]_  = ~A166 & \new_[54279]_ ;
  assign \new_[54281]_  = \new_[54280]_  & \new_[54275]_ ;
  assign \new_[54285]_  = ~A236 & ~A235;
  assign \new_[54286]_  = ~A233 & \new_[54285]_ ;
  assign \new_[54289]_  = ~A267 & ~A266;
  assign \new_[54292]_  = ~A299 & ~A298;
  assign \new_[54293]_  = \new_[54292]_  & \new_[54289]_ ;
  assign \new_[54294]_  = \new_[54293]_  & \new_[54286]_ ;
  assign \new_[54298]_  = ~A167 & A169;
  assign \new_[54299]_  = ~A170 & \new_[54298]_ ;
  assign \new_[54303]_  = ~A200 & ~A199;
  assign \new_[54304]_  = ~A166 & \new_[54303]_ ;
  assign \new_[54305]_  = \new_[54304]_  & \new_[54299]_ ;
  assign \new_[54309]_  = ~A236 & ~A235;
  assign \new_[54310]_  = ~A233 & \new_[54309]_ ;
  assign \new_[54313]_  = ~A266 & ~A265;
  assign \new_[54316]_  = ~A300 & A298;
  assign \new_[54317]_  = \new_[54316]_  & \new_[54313]_ ;
  assign \new_[54318]_  = \new_[54317]_  & \new_[54310]_ ;
  assign \new_[54322]_  = ~A167 & A169;
  assign \new_[54323]_  = ~A170 & \new_[54322]_ ;
  assign \new_[54327]_  = ~A200 & ~A199;
  assign \new_[54328]_  = ~A166 & \new_[54327]_ ;
  assign \new_[54329]_  = \new_[54328]_  & \new_[54323]_ ;
  assign \new_[54333]_  = ~A236 & ~A235;
  assign \new_[54334]_  = ~A233 & \new_[54333]_ ;
  assign \new_[54337]_  = ~A266 & ~A265;
  assign \new_[54340]_  = A299 & A298;
  assign \new_[54341]_  = \new_[54340]_  & \new_[54337]_ ;
  assign \new_[54342]_  = \new_[54341]_  & \new_[54334]_ ;
  assign \new_[54346]_  = ~A167 & A169;
  assign \new_[54347]_  = ~A170 & \new_[54346]_ ;
  assign \new_[54351]_  = ~A200 & ~A199;
  assign \new_[54352]_  = ~A166 & \new_[54351]_ ;
  assign \new_[54353]_  = \new_[54352]_  & \new_[54347]_ ;
  assign \new_[54357]_  = ~A236 & ~A235;
  assign \new_[54358]_  = ~A233 & \new_[54357]_ ;
  assign \new_[54361]_  = ~A266 & ~A265;
  assign \new_[54364]_  = ~A299 & ~A298;
  assign \new_[54365]_  = \new_[54364]_  & \new_[54361]_ ;
  assign \new_[54366]_  = \new_[54365]_  & \new_[54358]_ ;
  assign \new_[54370]_  = ~A167 & A169;
  assign \new_[54371]_  = ~A170 & \new_[54370]_ ;
  assign \new_[54375]_  = ~A200 & ~A199;
  assign \new_[54376]_  = ~A166 & \new_[54375]_ ;
  assign \new_[54377]_  = \new_[54376]_  & \new_[54371]_ ;
  assign \new_[54381]_  = A265 & ~A234;
  assign \new_[54382]_  = ~A233 & \new_[54381]_ ;
  assign \new_[54385]_  = A298 & A266;
  assign \new_[54388]_  = ~A302 & ~A301;
  assign \new_[54389]_  = \new_[54388]_  & \new_[54385]_ ;
  assign \new_[54390]_  = \new_[54389]_  & \new_[54382]_ ;
  assign \new_[54394]_  = ~A167 & A169;
  assign \new_[54395]_  = ~A170 & \new_[54394]_ ;
  assign \new_[54399]_  = ~A200 & ~A199;
  assign \new_[54400]_  = ~A166 & \new_[54399]_ ;
  assign \new_[54401]_  = \new_[54400]_  & \new_[54395]_ ;
  assign \new_[54405]_  = ~A266 & ~A234;
  assign \new_[54406]_  = ~A233 & \new_[54405]_ ;
  assign \new_[54409]_  = ~A269 & ~A268;
  assign \new_[54412]_  = ~A300 & A298;
  assign \new_[54413]_  = \new_[54412]_  & \new_[54409]_ ;
  assign \new_[54414]_  = \new_[54413]_  & \new_[54406]_ ;
  assign \new_[54418]_  = ~A167 & A169;
  assign \new_[54419]_  = ~A170 & \new_[54418]_ ;
  assign \new_[54423]_  = ~A200 & ~A199;
  assign \new_[54424]_  = ~A166 & \new_[54423]_ ;
  assign \new_[54425]_  = \new_[54424]_  & \new_[54419]_ ;
  assign \new_[54429]_  = ~A266 & ~A234;
  assign \new_[54430]_  = ~A233 & \new_[54429]_ ;
  assign \new_[54433]_  = ~A269 & ~A268;
  assign \new_[54436]_  = A299 & A298;
  assign \new_[54437]_  = \new_[54436]_  & \new_[54433]_ ;
  assign \new_[54438]_  = \new_[54437]_  & \new_[54430]_ ;
  assign \new_[54442]_  = ~A167 & A169;
  assign \new_[54443]_  = ~A170 & \new_[54442]_ ;
  assign \new_[54447]_  = ~A200 & ~A199;
  assign \new_[54448]_  = ~A166 & \new_[54447]_ ;
  assign \new_[54449]_  = \new_[54448]_  & \new_[54443]_ ;
  assign \new_[54453]_  = ~A266 & ~A234;
  assign \new_[54454]_  = ~A233 & \new_[54453]_ ;
  assign \new_[54457]_  = ~A269 & ~A268;
  assign \new_[54460]_  = ~A299 & ~A298;
  assign \new_[54461]_  = \new_[54460]_  & \new_[54457]_ ;
  assign \new_[54462]_  = \new_[54461]_  & \new_[54454]_ ;
  assign \new_[54466]_  = ~A167 & A169;
  assign \new_[54467]_  = ~A170 & \new_[54466]_ ;
  assign \new_[54471]_  = ~A200 & ~A199;
  assign \new_[54472]_  = ~A166 & \new_[54471]_ ;
  assign \new_[54473]_  = \new_[54472]_  & \new_[54467]_ ;
  assign \new_[54477]_  = ~A266 & ~A234;
  assign \new_[54478]_  = ~A233 & \new_[54477]_ ;
  assign \new_[54481]_  = A298 & ~A267;
  assign \new_[54484]_  = ~A302 & ~A301;
  assign \new_[54485]_  = \new_[54484]_  & \new_[54481]_ ;
  assign \new_[54486]_  = \new_[54485]_  & \new_[54478]_ ;
  assign \new_[54490]_  = ~A167 & A169;
  assign \new_[54491]_  = ~A170 & \new_[54490]_ ;
  assign \new_[54495]_  = ~A200 & ~A199;
  assign \new_[54496]_  = ~A166 & \new_[54495]_ ;
  assign \new_[54497]_  = \new_[54496]_  & \new_[54491]_ ;
  assign \new_[54501]_  = ~A265 & ~A234;
  assign \new_[54502]_  = ~A233 & \new_[54501]_ ;
  assign \new_[54505]_  = A298 & ~A266;
  assign \new_[54508]_  = ~A302 & ~A301;
  assign \new_[54509]_  = \new_[54508]_  & \new_[54505]_ ;
  assign \new_[54510]_  = \new_[54509]_  & \new_[54502]_ ;
  assign \new_[54514]_  = ~A167 & A169;
  assign \new_[54515]_  = ~A170 & \new_[54514]_ ;
  assign \new_[54519]_  = ~A200 & ~A199;
  assign \new_[54520]_  = ~A166 & \new_[54519]_ ;
  assign \new_[54521]_  = \new_[54520]_  & \new_[54515]_ ;
  assign \new_[54525]_  = A265 & ~A233;
  assign \new_[54526]_  = ~A232 & \new_[54525]_ ;
  assign \new_[54529]_  = A298 & A266;
  assign \new_[54532]_  = ~A302 & ~A301;
  assign \new_[54533]_  = \new_[54532]_  & \new_[54529]_ ;
  assign \new_[54534]_  = \new_[54533]_  & \new_[54526]_ ;
  assign \new_[54538]_  = ~A167 & A169;
  assign \new_[54539]_  = ~A170 & \new_[54538]_ ;
  assign \new_[54543]_  = ~A200 & ~A199;
  assign \new_[54544]_  = ~A166 & \new_[54543]_ ;
  assign \new_[54545]_  = \new_[54544]_  & \new_[54539]_ ;
  assign \new_[54549]_  = ~A266 & ~A233;
  assign \new_[54550]_  = ~A232 & \new_[54549]_ ;
  assign \new_[54553]_  = ~A269 & ~A268;
  assign \new_[54556]_  = ~A300 & A298;
  assign \new_[54557]_  = \new_[54556]_  & \new_[54553]_ ;
  assign \new_[54558]_  = \new_[54557]_  & \new_[54550]_ ;
  assign \new_[54562]_  = ~A167 & A169;
  assign \new_[54563]_  = ~A170 & \new_[54562]_ ;
  assign \new_[54567]_  = ~A200 & ~A199;
  assign \new_[54568]_  = ~A166 & \new_[54567]_ ;
  assign \new_[54569]_  = \new_[54568]_  & \new_[54563]_ ;
  assign \new_[54573]_  = ~A266 & ~A233;
  assign \new_[54574]_  = ~A232 & \new_[54573]_ ;
  assign \new_[54577]_  = ~A269 & ~A268;
  assign \new_[54580]_  = A299 & A298;
  assign \new_[54581]_  = \new_[54580]_  & \new_[54577]_ ;
  assign \new_[54582]_  = \new_[54581]_  & \new_[54574]_ ;
  assign \new_[54586]_  = ~A167 & A169;
  assign \new_[54587]_  = ~A170 & \new_[54586]_ ;
  assign \new_[54591]_  = ~A200 & ~A199;
  assign \new_[54592]_  = ~A166 & \new_[54591]_ ;
  assign \new_[54593]_  = \new_[54592]_  & \new_[54587]_ ;
  assign \new_[54597]_  = ~A266 & ~A233;
  assign \new_[54598]_  = ~A232 & \new_[54597]_ ;
  assign \new_[54601]_  = ~A269 & ~A268;
  assign \new_[54604]_  = ~A299 & ~A298;
  assign \new_[54605]_  = \new_[54604]_  & \new_[54601]_ ;
  assign \new_[54606]_  = \new_[54605]_  & \new_[54598]_ ;
  assign \new_[54610]_  = ~A167 & A169;
  assign \new_[54611]_  = ~A170 & \new_[54610]_ ;
  assign \new_[54615]_  = ~A200 & ~A199;
  assign \new_[54616]_  = ~A166 & \new_[54615]_ ;
  assign \new_[54617]_  = \new_[54616]_  & \new_[54611]_ ;
  assign \new_[54621]_  = ~A266 & ~A233;
  assign \new_[54622]_  = ~A232 & \new_[54621]_ ;
  assign \new_[54625]_  = A298 & ~A267;
  assign \new_[54628]_  = ~A302 & ~A301;
  assign \new_[54629]_  = \new_[54628]_  & \new_[54625]_ ;
  assign \new_[54630]_  = \new_[54629]_  & \new_[54622]_ ;
  assign \new_[54634]_  = ~A167 & A169;
  assign \new_[54635]_  = ~A170 & \new_[54634]_ ;
  assign \new_[54639]_  = ~A200 & ~A199;
  assign \new_[54640]_  = ~A166 & \new_[54639]_ ;
  assign \new_[54641]_  = \new_[54640]_  & \new_[54635]_ ;
  assign \new_[54645]_  = ~A265 & ~A233;
  assign \new_[54646]_  = ~A232 & \new_[54645]_ ;
  assign \new_[54649]_  = A298 & ~A266;
  assign \new_[54652]_  = ~A302 & ~A301;
  assign \new_[54653]_  = \new_[54652]_  & \new_[54649]_ ;
  assign \new_[54654]_  = \new_[54653]_  & \new_[54646]_ ;
  assign \new_[54658]_  = ~A166 & ~A167;
  assign \new_[54659]_  = ~A169 & \new_[54658]_ ;
  assign \new_[54663]_  = A232 & A200;
  assign \new_[54664]_  = ~A199 & \new_[54663]_ ;
  assign \new_[54665]_  = \new_[54664]_  & \new_[54659]_ ;
  assign \new_[54669]_  = ~A268 & A265;
  assign \new_[54670]_  = A233 & \new_[54669]_ ;
  assign \new_[54673]_  = ~A299 & ~A269;
  assign \new_[54676]_  = ~A302 & ~A301;
  assign \new_[54677]_  = \new_[54676]_  & \new_[54673]_ ;
  assign \new_[54678]_  = \new_[54677]_  & \new_[54670]_ ;
  assign \new_[54682]_  = ~A166 & ~A167;
  assign \new_[54683]_  = ~A169 & \new_[54682]_ ;
  assign \new_[54687]_  = ~A233 & A200;
  assign \new_[54688]_  = ~A199 & \new_[54687]_ ;
  assign \new_[54689]_  = \new_[54688]_  & \new_[54683]_ ;
  assign \new_[54693]_  = A265 & ~A236;
  assign \new_[54694]_  = ~A235 & \new_[54693]_ ;
  assign \new_[54697]_  = A298 & A266;
  assign \new_[54700]_  = ~A302 & ~A301;
  assign \new_[54701]_  = \new_[54700]_  & \new_[54697]_ ;
  assign \new_[54702]_  = \new_[54701]_  & \new_[54694]_ ;
  assign \new_[54706]_  = ~A166 & ~A167;
  assign \new_[54707]_  = ~A169 & \new_[54706]_ ;
  assign \new_[54711]_  = ~A233 & A200;
  assign \new_[54712]_  = ~A199 & \new_[54711]_ ;
  assign \new_[54713]_  = \new_[54712]_  & \new_[54707]_ ;
  assign \new_[54717]_  = ~A266 & ~A236;
  assign \new_[54718]_  = ~A235 & \new_[54717]_ ;
  assign \new_[54721]_  = ~A269 & ~A268;
  assign \new_[54724]_  = ~A300 & A298;
  assign \new_[54725]_  = \new_[54724]_  & \new_[54721]_ ;
  assign \new_[54726]_  = \new_[54725]_  & \new_[54718]_ ;
  assign \new_[54730]_  = ~A166 & ~A167;
  assign \new_[54731]_  = ~A169 & \new_[54730]_ ;
  assign \new_[54735]_  = ~A233 & A200;
  assign \new_[54736]_  = ~A199 & \new_[54735]_ ;
  assign \new_[54737]_  = \new_[54736]_  & \new_[54731]_ ;
  assign \new_[54741]_  = ~A266 & ~A236;
  assign \new_[54742]_  = ~A235 & \new_[54741]_ ;
  assign \new_[54745]_  = ~A269 & ~A268;
  assign \new_[54748]_  = A299 & A298;
  assign \new_[54749]_  = \new_[54748]_  & \new_[54745]_ ;
  assign \new_[54750]_  = \new_[54749]_  & \new_[54742]_ ;
  assign \new_[54754]_  = ~A166 & ~A167;
  assign \new_[54755]_  = ~A169 & \new_[54754]_ ;
  assign \new_[54759]_  = ~A233 & A200;
  assign \new_[54760]_  = ~A199 & \new_[54759]_ ;
  assign \new_[54761]_  = \new_[54760]_  & \new_[54755]_ ;
  assign \new_[54765]_  = ~A266 & ~A236;
  assign \new_[54766]_  = ~A235 & \new_[54765]_ ;
  assign \new_[54769]_  = ~A269 & ~A268;
  assign \new_[54772]_  = ~A299 & ~A298;
  assign \new_[54773]_  = \new_[54772]_  & \new_[54769]_ ;
  assign \new_[54774]_  = \new_[54773]_  & \new_[54766]_ ;
  assign \new_[54778]_  = ~A166 & ~A167;
  assign \new_[54779]_  = ~A169 & \new_[54778]_ ;
  assign \new_[54783]_  = ~A233 & A200;
  assign \new_[54784]_  = ~A199 & \new_[54783]_ ;
  assign \new_[54785]_  = \new_[54784]_  & \new_[54779]_ ;
  assign \new_[54789]_  = ~A266 & ~A236;
  assign \new_[54790]_  = ~A235 & \new_[54789]_ ;
  assign \new_[54793]_  = A298 & ~A267;
  assign \new_[54796]_  = ~A302 & ~A301;
  assign \new_[54797]_  = \new_[54796]_  & \new_[54793]_ ;
  assign \new_[54798]_  = \new_[54797]_  & \new_[54790]_ ;
  assign \new_[54802]_  = ~A166 & ~A167;
  assign \new_[54803]_  = ~A169 & \new_[54802]_ ;
  assign \new_[54807]_  = ~A233 & A200;
  assign \new_[54808]_  = ~A199 & \new_[54807]_ ;
  assign \new_[54809]_  = \new_[54808]_  & \new_[54803]_ ;
  assign \new_[54813]_  = ~A265 & ~A236;
  assign \new_[54814]_  = ~A235 & \new_[54813]_ ;
  assign \new_[54817]_  = A298 & ~A266;
  assign \new_[54820]_  = ~A302 & ~A301;
  assign \new_[54821]_  = \new_[54820]_  & \new_[54817]_ ;
  assign \new_[54822]_  = \new_[54821]_  & \new_[54814]_ ;
  assign \new_[54826]_  = ~A166 & ~A167;
  assign \new_[54827]_  = ~A169 & \new_[54826]_ ;
  assign \new_[54831]_  = ~A233 & A200;
  assign \new_[54832]_  = ~A199 & \new_[54831]_ ;
  assign \new_[54833]_  = \new_[54832]_  & \new_[54827]_ ;
  assign \new_[54837]_  = ~A268 & ~A266;
  assign \new_[54838]_  = ~A234 & \new_[54837]_ ;
  assign \new_[54841]_  = A298 & ~A269;
  assign \new_[54844]_  = ~A302 & ~A301;
  assign \new_[54845]_  = \new_[54844]_  & \new_[54841]_ ;
  assign \new_[54846]_  = \new_[54845]_  & \new_[54838]_ ;
  assign \new_[54850]_  = ~A166 & ~A167;
  assign \new_[54851]_  = ~A169 & \new_[54850]_ ;
  assign \new_[54855]_  = A232 & A200;
  assign \new_[54856]_  = ~A199 & \new_[54855]_ ;
  assign \new_[54857]_  = \new_[54856]_  & \new_[54851]_ ;
  assign \new_[54861]_  = A235 & A234;
  assign \new_[54862]_  = ~A233 & \new_[54861]_ ;
  assign \new_[54865]_  = ~A299 & A298;
  assign \new_[54868]_  = A301 & A300;
  assign \new_[54869]_  = \new_[54868]_  & \new_[54865]_ ;
  assign \new_[54870]_  = \new_[54869]_  & \new_[54862]_ ;
  assign \new_[54874]_  = ~A166 & ~A167;
  assign \new_[54875]_  = ~A169 & \new_[54874]_ ;
  assign \new_[54879]_  = A232 & A200;
  assign \new_[54880]_  = ~A199 & \new_[54879]_ ;
  assign \new_[54881]_  = \new_[54880]_  & \new_[54875]_ ;
  assign \new_[54885]_  = A235 & A234;
  assign \new_[54886]_  = ~A233 & \new_[54885]_ ;
  assign \new_[54889]_  = ~A299 & A298;
  assign \new_[54892]_  = A302 & A300;
  assign \new_[54893]_  = \new_[54892]_  & \new_[54889]_ ;
  assign \new_[54894]_  = \new_[54893]_  & \new_[54886]_ ;
  assign \new_[54898]_  = ~A166 & ~A167;
  assign \new_[54899]_  = ~A169 & \new_[54898]_ ;
  assign \new_[54903]_  = A232 & A200;
  assign \new_[54904]_  = ~A199 & \new_[54903]_ ;
  assign \new_[54905]_  = \new_[54904]_  & \new_[54899]_ ;
  assign \new_[54909]_  = A235 & A234;
  assign \new_[54910]_  = ~A233 & \new_[54909]_ ;
  assign \new_[54913]_  = ~A266 & A265;
  assign \new_[54916]_  = A268 & A267;
  assign \new_[54917]_  = \new_[54916]_  & \new_[54913]_ ;
  assign \new_[54918]_  = \new_[54917]_  & \new_[54910]_ ;
  assign \new_[54922]_  = ~A166 & ~A167;
  assign \new_[54923]_  = ~A169 & \new_[54922]_ ;
  assign \new_[54927]_  = A232 & A200;
  assign \new_[54928]_  = ~A199 & \new_[54927]_ ;
  assign \new_[54929]_  = \new_[54928]_  & \new_[54923]_ ;
  assign \new_[54933]_  = A235 & A234;
  assign \new_[54934]_  = ~A233 & \new_[54933]_ ;
  assign \new_[54937]_  = ~A266 & A265;
  assign \new_[54940]_  = A269 & A267;
  assign \new_[54941]_  = \new_[54940]_  & \new_[54937]_ ;
  assign \new_[54942]_  = \new_[54941]_  & \new_[54934]_ ;
  assign \new_[54946]_  = ~A166 & ~A167;
  assign \new_[54947]_  = ~A169 & \new_[54946]_ ;
  assign \new_[54951]_  = A232 & A200;
  assign \new_[54952]_  = ~A199 & \new_[54951]_ ;
  assign \new_[54953]_  = \new_[54952]_  & \new_[54947]_ ;
  assign \new_[54957]_  = A236 & A234;
  assign \new_[54958]_  = ~A233 & \new_[54957]_ ;
  assign \new_[54961]_  = ~A299 & A298;
  assign \new_[54964]_  = A301 & A300;
  assign \new_[54965]_  = \new_[54964]_  & \new_[54961]_ ;
  assign \new_[54966]_  = \new_[54965]_  & \new_[54958]_ ;
  assign \new_[54970]_  = ~A166 & ~A167;
  assign \new_[54971]_  = ~A169 & \new_[54970]_ ;
  assign \new_[54975]_  = A232 & A200;
  assign \new_[54976]_  = ~A199 & \new_[54975]_ ;
  assign \new_[54977]_  = \new_[54976]_  & \new_[54971]_ ;
  assign \new_[54981]_  = A236 & A234;
  assign \new_[54982]_  = ~A233 & \new_[54981]_ ;
  assign \new_[54985]_  = ~A299 & A298;
  assign \new_[54988]_  = A302 & A300;
  assign \new_[54989]_  = \new_[54988]_  & \new_[54985]_ ;
  assign \new_[54990]_  = \new_[54989]_  & \new_[54982]_ ;
  assign \new_[54994]_  = ~A166 & ~A167;
  assign \new_[54995]_  = ~A169 & \new_[54994]_ ;
  assign \new_[54999]_  = A232 & A200;
  assign \new_[55000]_  = ~A199 & \new_[54999]_ ;
  assign \new_[55001]_  = \new_[55000]_  & \new_[54995]_ ;
  assign \new_[55005]_  = A236 & A234;
  assign \new_[55006]_  = ~A233 & \new_[55005]_ ;
  assign \new_[55009]_  = ~A266 & A265;
  assign \new_[55012]_  = A268 & A267;
  assign \new_[55013]_  = \new_[55012]_  & \new_[55009]_ ;
  assign \new_[55014]_  = \new_[55013]_  & \new_[55006]_ ;
  assign \new_[55018]_  = ~A166 & ~A167;
  assign \new_[55019]_  = ~A169 & \new_[55018]_ ;
  assign \new_[55023]_  = A232 & A200;
  assign \new_[55024]_  = ~A199 & \new_[55023]_ ;
  assign \new_[55025]_  = \new_[55024]_  & \new_[55019]_ ;
  assign \new_[55029]_  = A236 & A234;
  assign \new_[55030]_  = ~A233 & \new_[55029]_ ;
  assign \new_[55033]_  = ~A266 & A265;
  assign \new_[55036]_  = A269 & A267;
  assign \new_[55037]_  = \new_[55036]_  & \new_[55033]_ ;
  assign \new_[55038]_  = \new_[55037]_  & \new_[55030]_ ;
  assign \new_[55042]_  = ~A166 & ~A167;
  assign \new_[55043]_  = ~A169 & \new_[55042]_ ;
  assign \new_[55047]_  = ~A232 & A200;
  assign \new_[55048]_  = ~A199 & \new_[55047]_ ;
  assign \new_[55049]_  = \new_[55048]_  & \new_[55043]_ ;
  assign \new_[55053]_  = ~A268 & ~A266;
  assign \new_[55054]_  = ~A233 & \new_[55053]_ ;
  assign \new_[55057]_  = A298 & ~A269;
  assign \new_[55060]_  = ~A302 & ~A301;
  assign \new_[55061]_  = \new_[55060]_  & \new_[55057]_ ;
  assign \new_[55062]_  = \new_[55061]_  & \new_[55054]_ ;
  assign \new_[55066]_  = ~A166 & ~A167;
  assign \new_[55067]_  = ~A169 & \new_[55066]_ ;
  assign \new_[55071]_  = A201 & ~A200;
  assign \new_[55072]_  = A199 & \new_[55071]_ ;
  assign \new_[55073]_  = \new_[55072]_  & \new_[55067]_ ;
  assign \new_[55077]_  = A233 & A232;
  assign \new_[55078]_  = A202 & \new_[55077]_ ;
  assign \new_[55081]_  = ~A267 & A265;
  assign \new_[55084]_  = ~A300 & ~A299;
  assign \new_[55085]_  = \new_[55084]_  & \new_[55081]_ ;
  assign \new_[55086]_  = \new_[55085]_  & \new_[55078]_ ;
  assign \new_[55090]_  = ~A166 & ~A167;
  assign \new_[55091]_  = ~A169 & \new_[55090]_ ;
  assign \new_[55095]_  = A201 & ~A200;
  assign \new_[55096]_  = A199 & \new_[55095]_ ;
  assign \new_[55097]_  = \new_[55096]_  & \new_[55091]_ ;
  assign \new_[55101]_  = A233 & A232;
  assign \new_[55102]_  = A202 & \new_[55101]_ ;
  assign \new_[55105]_  = ~A267 & A265;
  assign \new_[55108]_  = A299 & A298;
  assign \new_[55109]_  = \new_[55108]_  & \new_[55105]_ ;
  assign \new_[55110]_  = \new_[55109]_  & \new_[55102]_ ;
  assign \new_[55114]_  = ~A166 & ~A167;
  assign \new_[55115]_  = ~A169 & \new_[55114]_ ;
  assign \new_[55119]_  = A201 & ~A200;
  assign \new_[55120]_  = A199 & \new_[55119]_ ;
  assign \new_[55121]_  = \new_[55120]_  & \new_[55115]_ ;
  assign \new_[55125]_  = A233 & A232;
  assign \new_[55126]_  = A202 & \new_[55125]_ ;
  assign \new_[55129]_  = ~A267 & A265;
  assign \new_[55132]_  = ~A299 & ~A298;
  assign \new_[55133]_  = \new_[55132]_  & \new_[55129]_ ;
  assign \new_[55134]_  = \new_[55133]_  & \new_[55126]_ ;
  assign \new_[55138]_  = ~A166 & ~A167;
  assign \new_[55139]_  = ~A169 & \new_[55138]_ ;
  assign \new_[55143]_  = A201 & ~A200;
  assign \new_[55144]_  = A199 & \new_[55143]_ ;
  assign \new_[55145]_  = \new_[55144]_  & \new_[55139]_ ;
  assign \new_[55149]_  = A233 & A232;
  assign \new_[55150]_  = A202 & \new_[55149]_ ;
  assign \new_[55153]_  = A266 & A265;
  assign \new_[55156]_  = ~A300 & ~A299;
  assign \new_[55157]_  = \new_[55156]_  & \new_[55153]_ ;
  assign \new_[55158]_  = \new_[55157]_  & \new_[55150]_ ;
  assign \new_[55162]_  = ~A166 & ~A167;
  assign \new_[55163]_  = ~A169 & \new_[55162]_ ;
  assign \new_[55167]_  = A201 & ~A200;
  assign \new_[55168]_  = A199 & \new_[55167]_ ;
  assign \new_[55169]_  = \new_[55168]_  & \new_[55163]_ ;
  assign \new_[55173]_  = A233 & A232;
  assign \new_[55174]_  = A202 & \new_[55173]_ ;
  assign \new_[55177]_  = A266 & A265;
  assign \new_[55180]_  = A299 & A298;
  assign \new_[55181]_  = \new_[55180]_  & \new_[55177]_ ;
  assign \new_[55182]_  = \new_[55181]_  & \new_[55174]_ ;
  assign \new_[55186]_  = ~A166 & ~A167;
  assign \new_[55187]_  = ~A169 & \new_[55186]_ ;
  assign \new_[55191]_  = A201 & ~A200;
  assign \new_[55192]_  = A199 & \new_[55191]_ ;
  assign \new_[55193]_  = \new_[55192]_  & \new_[55187]_ ;
  assign \new_[55197]_  = A233 & A232;
  assign \new_[55198]_  = A202 & \new_[55197]_ ;
  assign \new_[55201]_  = A266 & A265;
  assign \new_[55204]_  = ~A299 & ~A298;
  assign \new_[55205]_  = \new_[55204]_  & \new_[55201]_ ;
  assign \new_[55206]_  = \new_[55205]_  & \new_[55198]_ ;
  assign \new_[55210]_  = ~A166 & ~A167;
  assign \new_[55211]_  = ~A169 & \new_[55210]_ ;
  assign \new_[55215]_  = A201 & ~A200;
  assign \new_[55216]_  = A199 & \new_[55215]_ ;
  assign \new_[55217]_  = \new_[55216]_  & \new_[55211]_ ;
  assign \new_[55221]_  = A233 & A232;
  assign \new_[55222]_  = A202 & \new_[55221]_ ;
  assign \new_[55225]_  = ~A266 & ~A265;
  assign \new_[55228]_  = ~A300 & ~A299;
  assign \new_[55229]_  = \new_[55228]_  & \new_[55225]_ ;
  assign \new_[55230]_  = \new_[55229]_  & \new_[55222]_ ;
  assign \new_[55234]_  = ~A166 & ~A167;
  assign \new_[55235]_  = ~A169 & \new_[55234]_ ;
  assign \new_[55239]_  = A201 & ~A200;
  assign \new_[55240]_  = A199 & \new_[55239]_ ;
  assign \new_[55241]_  = \new_[55240]_  & \new_[55235]_ ;
  assign \new_[55245]_  = A233 & A232;
  assign \new_[55246]_  = A202 & \new_[55245]_ ;
  assign \new_[55249]_  = ~A266 & ~A265;
  assign \new_[55252]_  = A299 & A298;
  assign \new_[55253]_  = \new_[55252]_  & \new_[55249]_ ;
  assign \new_[55254]_  = \new_[55253]_  & \new_[55246]_ ;
  assign \new_[55258]_  = ~A166 & ~A167;
  assign \new_[55259]_  = ~A169 & \new_[55258]_ ;
  assign \new_[55263]_  = A201 & ~A200;
  assign \new_[55264]_  = A199 & \new_[55263]_ ;
  assign \new_[55265]_  = \new_[55264]_  & \new_[55259]_ ;
  assign \new_[55269]_  = A233 & A232;
  assign \new_[55270]_  = A202 & \new_[55269]_ ;
  assign \new_[55273]_  = ~A266 & ~A265;
  assign \new_[55276]_  = ~A299 & ~A298;
  assign \new_[55277]_  = \new_[55276]_  & \new_[55273]_ ;
  assign \new_[55278]_  = \new_[55277]_  & \new_[55270]_ ;
  assign \new_[55282]_  = ~A166 & ~A167;
  assign \new_[55283]_  = ~A169 & \new_[55282]_ ;
  assign \new_[55287]_  = A201 & ~A200;
  assign \new_[55288]_  = A199 & \new_[55287]_ ;
  assign \new_[55289]_  = \new_[55288]_  & \new_[55283]_ ;
  assign \new_[55293]_  = A233 & ~A232;
  assign \new_[55294]_  = A202 & \new_[55293]_ ;
  assign \new_[55297]_  = ~A299 & A298;
  assign \new_[55300]_  = A301 & A300;
  assign \new_[55301]_  = \new_[55300]_  & \new_[55297]_ ;
  assign \new_[55302]_  = \new_[55301]_  & \new_[55294]_ ;
  assign \new_[55306]_  = ~A166 & ~A167;
  assign \new_[55307]_  = ~A169 & \new_[55306]_ ;
  assign \new_[55311]_  = A201 & ~A200;
  assign \new_[55312]_  = A199 & \new_[55311]_ ;
  assign \new_[55313]_  = \new_[55312]_  & \new_[55307]_ ;
  assign \new_[55317]_  = A233 & ~A232;
  assign \new_[55318]_  = A202 & \new_[55317]_ ;
  assign \new_[55321]_  = ~A299 & A298;
  assign \new_[55324]_  = A302 & A300;
  assign \new_[55325]_  = \new_[55324]_  & \new_[55321]_ ;
  assign \new_[55326]_  = \new_[55325]_  & \new_[55318]_ ;
  assign \new_[55330]_  = ~A166 & ~A167;
  assign \new_[55331]_  = ~A169 & \new_[55330]_ ;
  assign \new_[55335]_  = A201 & ~A200;
  assign \new_[55336]_  = A199 & \new_[55335]_ ;
  assign \new_[55337]_  = \new_[55336]_  & \new_[55331]_ ;
  assign \new_[55341]_  = A233 & ~A232;
  assign \new_[55342]_  = A202 & \new_[55341]_ ;
  assign \new_[55345]_  = ~A266 & A265;
  assign \new_[55348]_  = A268 & A267;
  assign \new_[55349]_  = \new_[55348]_  & \new_[55345]_ ;
  assign \new_[55350]_  = \new_[55349]_  & \new_[55342]_ ;
  assign \new_[55354]_  = ~A166 & ~A167;
  assign \new_[55355]_  = ~A169 & \new_[55354]_ ;
  assign \new_[55359]_  = A201 & ~A200;
  assign \new_[55360]_  = A199 & \new_[55359]_ ;
  assign \new_[55361]_  = \new_[55360]_  & \new_[55355]_ ;
  assign \new_[55365]_  = A233 & ~A232;
  assign \new_[55366]_  = A202 & \new_[55365]_ ;
  assign \new_[55369]_  = ~A266 & A265;
  assign \new_[55372]_  = A269 & A267;
  assign \new_[55373]_  = \new_[55372]_  & \new_[55369]_ ;
  assign \new_[55374]_  = \new_[55373]_  & \new_[55366]_ ;
  assign \new_[55378]_  = ~A166 & ~A167;
  assign \new_[55379]_  = ~A169 & \new_[55378]_ ;
  assign \new_[55383]_  = A201 & ~A200;
  assign \new_[55384]_  = A199 & \new_[55383]_ ;
  assign \new_[55385]_  = \new_[55384]_  & \new_[55379]_ ;
  assign \new_[55389]_  = ~A234 & ~A233;
  assign \new_[55390]_  = A202 & \new_[55389]_ ;
  assign \new_[55393]_  = A266 & A265;
  assign \new_[55396]_  = ~A300 & A298;
  assign \new_[55397]_  = \new_[55396]_  & \new_[55393]_ ;
  assign \new_[55398]_  = \new_[55397]_  & \new_[55390]_ ;
  assign \new_[55402]_  = ~A166 & ~A167;
  assign \new_[55403]_  = ~A169 & \new_[55402]_ ;
  assign \new_[55407]_  = A201 & ~A200;
  assign \new_[55408]_  = A199 & \new_[55407]_ ;
  assign \new_[55409]_  = \new_[55408]_  & \new_[55403]_ ;
  assign \new_[55413]_  = ~A234 & ~A233;
  assign \new_[55414]_  = A202 & \new_[55413]_ ;
  assign \new_[55417]_  = A266 & A265;
  assign \new_[55420]_  = A299 & A298;
  assign \new_[55421]_  = \new_[55420]_  & \new_[55417]_ ;
  assign \new_[55422]_  = \new_[55421]_  & \new_[55414]_ ;
  assign \new_[55426]_  = ~A166 & ~A167;
  assign \new_[55427]_  = ~A169 & \new_[55426]_ ;
  assign \new_[55431]_  = A201 & ~A200;
  assign \new_[55432]_  = A199 & \new_[55431]_ ;
  assign \new_[55433]_  = \new_[55432]_  & \new_[55427]_ ;
  assign \new_[55437]_  = ~A234 & ~A233;
  assign \new_[55438]_  = A202 & \new_[55437]_ ;
  assign \new_[55441]_  = A266 & A265;
  assign \new_[55444]_  = ~A299 & ~A298;
  assign \new_[55445]_  = \new_[55444]_  & \new_[55441]_ ;
  assign \new_[55446]_  = \new_[55445]_  & \new_[55438]_ ;
  assign \new_[55450]_  = ~A166 & ~A167;
  assign \new_[55451]_  = ~A169 & \new_[55450]_ ;
  assign \new_[55455]_  = A201 & ~A200;
  assign \new_[55456]_  = A199 & \new_[55455]_ ;
  assign \new_[55457]_  = \new_[55456]_  & \new_[55451]_ ;
  assign \new_[55461]_  = ~A234 & ~A233;
  assign \new_[55462]_  = A202 & \new_[55461]_ ;
  assign \new_[55465]_  = ~A267 & ~A266;
  assign \new_[55468]_  = ~A300 & A298;
  assign \new_[55469]_  = \new_[55468]_  & \new_[55465]_ ;
  assign \new_[55470]_  = \new_[55469]_  & \new_[55462]_ ;
  assign \new_[55474]_  = ~A166 & ~A167;
  assign \new_[55475]_  = ~A169 & \new_[55474]_ ;
  assign \new_[55479]_  = A201 & ~A200;
  assign \new_[55480]_  = A199 & \new_[55479]_ ;
  assign \new_[55481]_  = \new_[55480]_  & \new_[55475]_ ;
  assign \new_[55485]_  = ~A234 & ~A233;
  assign \new_[55486]_  = A202 & \new_[55485]_ ;
  assign \new_[55489]_  = ~A267 & ~A266;
  assign \new_[55492]_  = A299 & A298;
  assign \new_[55493]_  = \new_[55492]_  & \new_[55489]_ ;
  assign \new_[55494]_  = \new_[55493]_  & \new_[55486]_ ;
  assign \new_[55498]_  = ~A166 & ~A167;
  assign \new_[55499]_  = ~A169 & \new_[55498]_ ;
  assign \new_[55503]_  = A201 & ~A200;
  assign \new_[55504]_  = A199 & \new_[55503]_ ;
  assign \new_[55505]_  = \new_[55504]_  & \new_[55499]_ ;
  assign \new_[55509]_  = ~A234 & ~A233;
  assign \new_[55510]_  = A202 & \new_[55509]_ ;
  assign \new_[55513]_  = ~A267 & ~A266;
  assign \new_[55516]_  = ~A299 & ~A298;
  assign \new_[55517]_  = \new_[55516]_  & \new_[55513]_ ;
  assign \new_[55518]_  = \new_[55517]_  & \new_[55510]_ ;
  assign \new_[55522]_  = ~A166 & ~A167;
  assign \new_[55523]_  = ~A169 & \new_[55522]_ ;
  assign \new_[55527]_  = A201 & ~A200;
  assign \new_[55528]_  = A199 & \new_[55527]_ ;
  assign \new_[55529]_  = \new_[55528]_  & \new_[55523]_ ;
  assign \new_[55533]_  = ~A234 & ~A233;
  assign \new_[55534]_  = A202 & \new_[55533]_ ;
  assign \new_[55537]_  = ~A266 & ~A265;
  assign \new_[55540]_  = ~A300 & A298;
  assign \new_[55541]_  = \new_[55540]_  & \new_[55537]_ ;
  assign \new_[55542]_  = \new_[55541]_  & \new_[55534]_ ;
  assign \new_[55546]_  = ~A166 & ~A167;
  assign \new_[55547]_  = ~A169 & \new_[55546]_ ;
  assign \new_[55551]_  = A201 & ~A200;
  assign \new_[55552]_  = A199 & \new_[55551]_ ;
  assign \new_[55553]_  = \new_[55552]_  & \new_[55547]_ ;
  assign \new_[55557]_  = ~A234 & ~A233;
  assign \new_[55558]_  = A202 & \new_[55557]_ ;
  assign \new_[55561]_  = ~A266 & ~A265;
  assign \new_[55564]_  = A299 & A298;
  assign \new_[55565]_  = \new_[55564]_  & \new_[55561]_ ;
  assign \new_[55566]_  = \new_[55565]_  & \new_[55558]_ ;
  assign \new_[55570]_  = ~A166 & ~A167;
  assign \new_[55571]_  = ~A169 & \new_[55570]_ ;
  assign \new_[55575]_  = A201 & ~A200;
  assign \new_[55576]_  = A199 & \new_[55575]_ ;
  assign \new_[55577]_  = \new_[55576]_  & \new_[55571]_ ;
  assign \new_[55581]_  = ~A234 & ~A233;
  assign \new_[55582]_  = A202 & \new_[55581]_ ;
  assign \new_[55585]_  = ~A266 & ~A265;
  assign \new_[55588]_  = ~A299 & ~A298;
  assign \new_[55589]_  = \new_[55588]_  & \new_[55585]_ ;
  assign \new_[55590]_  = \new_[55589]_  & \new_[55582]_ ;
  assign \new_[55594]_  = ~A166 & ~A167;
  assign \new_[55595]_  = ~A169 & \new_[55594]_ ;
  assign \new_[55599]_  = A201 & ~A200;
  assign \new_[55600]_  = A199 & \new_[55599]_ ;
  assign \new_[55601]_  = \new_[55600]_  & \new_[55595]_ ;
  assign \new_[55605]_  = ~A233 & A232;
  assign \new_[55606]_  = A202 & \new_[55605]_ ;
  assign \new_[55609]_  = A235 & A234;
  assign \new_[55612]_  = A299 & ~A298;
  assign \new_[55613]_  = \new_[55612]_  & \new_[55609]_ ;
  assign \new_[55614]_  = \new_[55613]_  & \new_[55606]_ ;
  assign \new_[55618]_  = ~A166 & ~A167;
  assign \new_[55619]_  = ~A169 & \new_[55618]_ ;
  assign \new_[55623]_  = A201 & ~A200;
  assign \new_[55624]_  = A199 & \new_[55623]_ ;
  assign \new_[55625]_  = \new_[55624]_  & \new_[55619]_ ;
  assign \new_[55629]_  = ~A233 & A232;
  assign \new_[55630]_  = A202 & \new_[55629]_ ;
  assign \new_[55633]_  = A235 & A234;
  assign \new_[55636]_  = A266 & ~A265;
  assign \new_[55637]_  = \new_[55636]_  & \new_[55633]_ ;
  assign \new_[55638]_  = \new_[55637]_  & \new_[55630]_ ;
  assign \new_[55642]_  = ~A166 & ~A167;
  assign \new_[55643]_  = ~A169 & \new_[55642]_ ;
  assign \new_[55647]_  = A201 & ~A200;
  assign \new_[55648]_  = A199 & \new_[55647]_ ;
  assign \new_[55649]_  = \new_[55648]_  & \new_[55643]_ ;
  assign \new_[55653]_  = ~A233 & A232;
  assign \new_[55654]_  = A202 & \new_[55653]_ ;
  assign \new_[55657]_  = A236 & A234;
  assign \new_[55660]_  = A299 & ~A298;
  assign \new_[55661]_  = \new_[55660]_  & \new_[55657]_ ;
  assign \new_[55662]_  = \new_[55661]_  & \new_[55654]_ ;
  assign \new_[55666]_  = ~A166 & ~A167;
  assign \new_[55667]_  = ~A169 & \new_[55666]_ ;
  assign \new_[55671]_  = A201 & ~A200;
  assign \new_[55672]_  = A199 & \new_[55671]_ ;
  assign \new_[55673]_  = \new_[55672]_  & \new_[55667]_ ;
  assign \new_[55677]_  = ~A233 & A232;
  assign \new_[55678]_  = A202 & \new_[55677]_ ;
  assign \new_[55681]_  = A236 & A234;
  assign \new_[55684]_  = A266 & ~A265;
  assign \new_[55685]_  = \new_[55684]_  & \new_[55681]_ ;
  assign \new_[55686]_  = \new_[55685]_  & \new_[55678]_ ;
  assign \new_[55690]_  = ~A166 & ~A167;
  assign \new_[55691]_  = ~A169 & \new_[55690]_ ;
  assign \new_[55695]_  = A201 & ~A200;
  assign \new_[55696]_  = A199 & \new_[55695]_ ;
  assign \new_[55697]_  = \new_[55696]_  & \new_[55691]_ ;
  assign \new_[55701]_  = ~A233 & ~A232;
  assign \new_[55702]_  = A202 & \new_[55701]_ ;
  assign \new_[55705]_  = A266 & A265;
  assign \new_[55708]_  = ~A300 & A298;
  assign \new_[55709]_  = \new_[55708]_  & \new_[55705]_ ;
  assign \new_[55710]_  = \new_[55709]_  & \new_[55702]_ ;
  assign \new_[55714]_  = ~A166 & ~A167;
  assign \new_[55715]_  = ~A169 & \new_[55714]_ ;
  assign \new_[55719]_  = A201 & ~A200;
  assign \new_[55720]_  = A199 & \new_[55719]_ ;
  assign \new_[55721]_  = \new_[55720]_  & \new_[55715]_ ;
  assign \new_[55725]_  = ~A233 & ~A232;
  assign \new_[55726]_  = A202 & \new_[55725]_ ;
  assign \new_[55729]_  = A266 & A265;
  assign \new_[55732]_  = A299 & A298;
  assign \new_[55733]_  = \new_[55732]_  & \new_[55729]_ ;
  assign \new_[55734]_  = \new_[55733]_  & \new_[55726]_ ;
  assign \new_[55738]_  = ~A166 & ~A167;
  assign \new_[55739]_  = ~A169 & \new_[55738]_ ;
  assign \new_[55743]_  = A201 & ~A200;
  assign \new_[55744]_  = A199 & \new_[55743]_ ;
  assign \new_[55745]_  = \new_[55744]_  & \new_[55739]_ ;
  assign \new_[55749]_  = ~A233 & ~A232;
  assign \new_[55750]_  = A202 & \new_[55749]_ ;
  assign \new_[55753]_  = A266 & A265;
  assign \new_[55756]_  = ~A299 & ~A298;
  assign \new_[55757]_  = \new_[55756]_  & \new_[55753]_ ;
  assign \new_[55758]_  = \new_[55757]_  & \new_[55750]_ ;
  assign \new_[55762]_  = ~A166 & ~A167;
  assign \new_[55763]_  = ~A169 & \new_[55762]_ ;
  assign \new_[55767]_  = A201 & ~A200;
  assign \new_[55768]_  = A199 & \new_[55767]_ ;
  assign \new_[55769]_  = \new_[55768]_  & \new_[55763]_ ;
  assign \new_[55773]_  = ~A233 & ~A232;
  assign \new_[55774]_  = A202 & \new_[55773]_ ;
  assign \new_[55777]_  = ~A267 & ~A266;
  assign \new_[55780]_  = ~A300 & A298;
  assign \new_[55781]_  = \new_[55780]_  & \new_[55777]_ ;
  assign \new_[55782]_  = \new_[55781]_  & \new_[55774]_ ;
  assign \new_[55786]_  = ~A166 & ~A167;
  assign \new_[55787]_  = ~A169 & \new_[55786]_ ;
  assign \new_[55791]_  = A201 & ~A200;
  assign \new_[55792]_  = A199 & \new_[55791]_ ;
  assign \new_[55793]_  = \new_[55792]_  & \new_[55787]_ ;
  assign \new_[55797]_  = ~A233 & ~A232;
  assign \new_[55798]_  = A202 & \new_[55797]_ ;
  assign \new_[55801]_  = ~A267 & ~A266;
  assign \new_[55804]_  = A299 & A298;
  assign \new_[55805]_  = \new_[55804]_  & \new_[55801]_ ;
  assign \new_[55806]_  = \new_[55805]_  & \new_[55798]_ ;
  assign \new_[55810]_  = ~A166 & ~A167;
  assign \new_[55811]_  = ~A169 & \new_[55810]_ ;
  assign \new_[55815]_  = A201 & ~A200;
  assign \new_[55816]_  = A199 & \new_[55815]_ ;
  assign \new_[55817]_  = \new_[55816]_  & \new_[55811]_ ;
  assign \new_[55821]_  = ~A233 & ~A232;
  assign \new_[55822]_  = A202 & \new_[55821]_ ;
  assign \new_[55825]_  = ~A267 & ~A266;
  assign \new_[55828]_  = ~A299 & ~A298;
  assign \new_[55829]_  = \new_[55828]_  & \new_[55825]_ ;
  assign \new_[55830]_  = \new_[55829]_  & \new_[55822]_ ;
  assign \new_[55834]_  = ~A166 & ~A167;
  assign \new_[55835]_  = ~A169 & \new_[55834]_ ;
  assign \new_[55839]_  = A201 & ~A200;
  assign \new_[55840]_  = A199 & \new_[55839]_ ;
  assign \new_[55841]_  = \new_[55840]_  & \new_[55835]_ ;
  assign \new_[55845]_  = ~A233 & ~A232;
  assign \new_[55846]_  = A202 & \new_[55845]_ ;
  assign \new_[55849]_  = ~A266 & ~A265;
  assign \new_[55852]_  = ~A300 & A298;
  assign \new_[55853]_  = \new_[55852]_  & \new_[55849]_ ;
  assign \new_[55854]_  = \new_[55853]_  & \new_[55846]_ ;
  assign \new_[55858]_  = ~A166 & ~A167;
  assign \new_[55859]_  = ~A169 & \new_[55858]_ ;
  assign \new_[55863]_  = A201 & ~A200;
  assign \new_[55864]_  = A199 & \new_[55863]_ ;
  assign \new_[55865]_  = \new_[55864]_  & \new_[55859]_ ;
  assign \new_[55869]_  = ~A233 & ~A232;
  assign \new_[55870]_  = A202 & \new_[55869]_ ;
  assign \new_[55873]_  = ~A266 & ~A265;
  assign \new_[55876]_  = A299 & A298;
  assign \new_[55877]_  = \new_[55876]_  & \new_[55873]_ ;
  assign \new_[55878]_  = \new_[55877]_  & \new_[55870]_ ;
  assign \new_[55882]_  = ~A166 & ~A167;
  assign \new_[55883]_  = ~A169 & \new_[55882]_ ;
  assign \new_[55887]_  = A201 & ~A200;
  assign \new_[55888]_  = A199 & \new_[55887]_ ;
  assign \new_[55889]_  = \new_[55888]_  & \new_[55883]_ ;
  assign \new_[55893]_  = ~A233 & ~A232;
  assign \new_[55894]_  = A202 & \new_[55893]_ ;
  assign \new_[55897]_  = ~A266 & ~A265;
  assign \new_[55900]_  = ~A299 & ~A298;
  assign \new_[55901]_  = \new_[55900]_  & \new_[55897]_ ;
  assign \new_[55902]_  = \new_[55901]_  & \new_[55894]_ ;
  assign \new_[55906]_  = ~A166 & ~A167;
  assign \new_[55907]_  = ~A169 & \new_[55906]_ ;
  assign \new_[55911]_  = A201 & ~A200;
  assign \new_[55912]_  = A199 & \new_[55911]_ ;
  assign \new_[55913]_  = \new_[55912]_  & \new_[55907]_ ;
  assign \new_[55917]_  = A233 & A232;
  assign \new_[55918]_  = A203 & \new_[55917]_ ;
  assign \new_[55921]_  = ~A267 & A265;
  assign \new_[55924]_  = ~A300 & ~A299;
  assign \new_[55925]_  = \new_[55924]_  & \new_[55921]_ ;
  assign \new_[55926]_  = \new_[55925]_  & \new_[55918]_ ;
  assign \new_[55930]_  = ~A166 & ~A167;
  assign \new_[55931]_  = ~A169 & \new_[55930]_ ;
  assign \new_[55935]_  = A201 & ~A200;
  assign \new_[55936]_  = A199 & \new_[55935]_ ;
  assign \new_[55937]_  = \new_[55936]_  & \new_[55931]_ ;
  assign \new_[55941]_  = A233 & A232;
  assign \new_[55942]_  = A203 & \new_[55941]_ ;
  assign \new_[55945]_  = ~A267 & A265;
  assign \new_[55948]_  = A299 & A298;
  assign \new_[55949]_  = \new_[55948]_  & \new_[55945]_ ;
  assign \new_[55950]_  = \new_[55949]_  & \new_[55942]_ ;
  assign \new_[55954]_  = ~A166 & ~A167;
  assign \new_[55955]_  = ~A169 & \new_[55954]_ ;
  assign \new_[55959]_  = A201 & ~A200;
  assign \new_[55960]_  = A199 & \new_[55959]_ ;
  assign \new_[55961]_  = \new_[55960]_  & \new_[55955]_ ;
  assign \new_[55965]_  = A233 & A232;
  assign \new_[55966]_  = A203 & \new_[55965]_ ;
  assign \new_[55969]_  = ~A267 & A265;
  assign \new_[55972]_  = ~A299 & ~A298;
  assign \new_[55973]_  = \new_[55972]_  & \new_[55969]_ ;
  assign \new_[55974]_  = \new_[55973]_  & \new_[55966]_ ;
  assign \new_[55978]_  = ~A166 & ~A167;
  assign \new_[55979]_  = ~A169 & \new_[55978]_ ;
  assign \new_[55983]_  = A201 & ~A200;
  assign \new_[55984]_  = A199 & \new_[55983]_ ;
  assign \new_[55985]_  = \new_[55984]_  & \new_[55979]_ ;
  assign \new_[55989]_  = A233 & A232;
  assign \new_[55990]_  = A203 & \new_[55989]_ ;
  assign \new_[55993]_  = A266 & A265;
  assign \new_[55996]_  = ~A300 & ~A299;
  assign \new_[55997]_  = \new_[55996]_  & \new_[55993]_ ;
  assign \new_[55998]_  = \new_[55997]_  & \new_[55990]_ ;
  assign \new_[56002]_  = ~A166 & ~A167;
  assign \new_[56003]_  = ~A169 & \new_[56002]_ ;
  assign \new_[56007]_  = A201 & ~A200;
  assign \new_[56008]_  = A199 & \new_[56007]_ ;
  assign \new_[56009]_  = \new_[56008]_  & \new_[56003]_ ;
  assign \new_[56013]_  = A233 & A232;
  assign \new_[56014]_  = A203 & \new_[56013]_ ;
  assign \new_[56017]_  = A266 & A265;
  assign \new_[56020]_  = A299 & A298;
  assign \new_[56021]_  = \new_[56020]_  & \new_[56017]_ ;
  assign \new_[56022]_  = \new_[56021]_  & \new_[56014]_ ;
  assign \new_[56026]_  = ~A166 & ~A167;
  assign \new_[56027]_  = ~A169 & \new_[56026]_ ;
  assign \new_[56031]_  = A201 & ~A200;
  assign \new_[56032]_  = A199 & \new_[56031]_ ;
  assign \new_[56033]_  = \new_[56032]_  & \new_[56027]_ ;
  assign \new_[56037]_  = A233 & A232;
  assign \new_[56038]_  = A203 & \new_[56037]_ ;
  assign \new_[56041]_  = A266 & A265;
  assign \new_[56044]_  = ~A299 & ~A298;
  assign \new_[56045]_  = \new_[56044]_  & \new_[56041]_ ;
  assign \new_[56046]_  = \new_[56045]_  & \new_[56038]_ ;
  assign \new_[56050]_  = ~A166 & ~A167;
  assign \new_[56051]_  = ~A169 & \new_[56050]_ ;
  assign \new_[56055]_  = A201 & ~A200;
  assign \new_[56056]_  = A199 & \new_[56055]_ ;
  assign \new_[56057]_  = \new_[56056]_  & \new_[56051]_ ;
  assign \new_[56061]_  = A233 & A232;
  assign \new_[56062]_  = A203 & \new_[56061]_ ;
  assign \new_[56065]_  = ~A266 & ~A265;
  assign \new_[56068]_  = ~A300 & ~A299;
  assign \new_[56069]_  = \new_[56068]_  & \new_[56065]_ ;
  assign \new_[56070]_  = \new_[56069]_  & \new_[56062]_ ;
  assign \new_[56074]_  = ~A166 & ~A167;
  assign \new_[56075]_  = ~A169 & \new_[56074]_ ;
  assign \new_[56079]_  = A201 & ~A200;
  assign \new_[56080]_  = A199 & \new_[56079]_ ;
  assign \new_[56081]_  = \new_[56080]_  & \new_[56075]_ ;
  assign \new_[56085]_  = A233 & A232;
  assign \new_[56086]_  = A203 & \new_[56085]_ ;
  assign \new_[56089]_  = ~A266 & ~A265;
  assign \new_[56092]_  = A299 & A298;
  assign \new_[56093]_  = \new_[56092]_  & \new_[56089]_ ;
  assign \new_[56094]_  = \new_[56093]_  & \new_[56086]_ ;
  assign \new_[56098]_  = ~A166 & ~A167;
  assign \new_[56099]_  = ~A169 & \new_[56098]_ ;
  assign \new_[56103]_  = A201 & ~A200;
  assign \new_[56104]_  = A199 & \new_[56103]_ ;
  assign \new_[56105]_  = \new_[56104]_  & \new_[56099]_ ;
  assign \new_[56109]_  = A233 & A232;
  assign \new_[56110]_  = A203 & \new_[56109]_ ;
  assign \new_[56113]_  = ~A266 & ~A265;
  assign \new_[56116]_  = ~A299 & ~A298;
  assign \new_[56117]_  = \new_[56116]_  & \new_[56113]_ ;
  assign \new_[56118]_  = \new_[56117]_  & \new_[56110]_ ;
  assign \new_[56122]_  = ~A166 & ~A167;
  assign \new_[56123]_  = ~A169 & \new_[56122]_ ;
  assign \new_[56127]_  = A201 & ~A200;
  assign \new_[56128]_  = A199 & \new_[56127]_ ;
  assign \new_[56129]_  = \new_[56128]_  & \new_[56123]_ ;
  assign \new_[56133]_  = A233 & ~A232;
  assign \new_[56134]_  = A203 & \new_[56133]_ ;
  assign \new_[56137]_  = ~A299 & A298;
  assign \new_[56140]_  = A301 & A300;
  assign \new_[56141]_  = \new_[56140]_  & \new_[56137]_ ;
  assign \new_[56142]_  = \new_[56141]_  & \new_[56134]_ ;
  assign \new_[56146]_  = ~A166 & ~A167;
  assign \new_[56147]_  = ~A169 & \new_[56146]_ ;
  assign \new_[56151]_  = A201 & ~A200;
  assign \new_[56152]_  = A199 & \new_[56151]_ ;
  assign \new_[56153]_  = \new_[56152]_  & \new_[56147]_ ;
  assign \new_[56157]_  = A233 & ~A232;
  assign \new_[56158]_  = A203 & \new_[56157]_ ;
  assign \new_[56161]_  = ~A299 & A298;
  assign \new_[56164]_  = A302 & A300;
  assign \new_[56165]_  = \new_[56164]_  & \new_[56161]_ ;
  assign \new_[56166]_  = \new_[56165]_  & \new_[56158]_ ;
  assign \new_[56170]_  = ~A166 & ~A167;
  assign \new_[56171]_  = ~A169 & \new_[56170]_ ;
  assign \new_[56175]_  = A201 & ~A200;
  assign \new_[56176]_  = A199 & \new_[56175]_ ;
  assign \new_[56177]_  = \new_[56176]_  & \new_[56171]_ ;
  assign \new_[56181]_  = A233 & ~A232;
  assign \new_[56182]_  = A203 & \new_[56181]_ ;
  assign \new_[56185]_  = ~A266 & A265;
  assign \new_[56188]_  = A268 & A267;
  assign \new_[56189]_  = \new_[56188]_  & \new_[56185]_ ;
  assign \new_[56190]_  = \new_[56189]_  & \new_[56182]_ ;
  assign \new_[56194]_  = ~A166 & ~A167;
  assign \new_[56195]_  = ~A169 & \new_[56194]_ ;
  assign \new_[56199]_  = A201 & ~A200;
  assign \new_[56200]_  = A199 & \new_[56199]_ ;
  assign \new_[56201]_  = \new_[56200]_  & \new_[56195]_ ;
  assign \new_[56205]_  = A233 & ~A232;
  assign \new_[56206]_  = A203 & \new_[56205]_ ;
  assign \new_[56209]_  = ~A266 & A265;
  assign \new_[56212]_  = A269 & A267;
  assign \new_[56213]_  = \new_[56212]_  & \new_[56209]_ ;
  assign \new_[56214]_  = \new_[56213]_  & \new_[56206]_ ;
  assign \new_[56218]_  = ~A166 & ~A167;
  assign \new_[56219]_  = ~A169 & \new_[56218]_ ;
  assign \new_[56223]_  = A201 & ~A200;
  assign \new_[56224]_  = A199 & \new_[56223]_ ;
  assign \new_[56225]_  = \new_[56224]_  & \new_[56219]_ ;
  assign \new_[56229]_  = ~A234 & ~A233;
  assign \new_[56230]_  = A203 & \new_[56229]_ ;
  assign \new_[56233]_  = A266 & A265;
  assign \new_[56236]_  = ~A300 & A298;
  assign \new_[56237]_  = \new_[56236]_  & \new_[56233]_ ;
  assign \new_[56238]_  = \new_[56237]_  & \new_[56230]_ ;
  assign \new_[56242]_  = ~A166 & ~A167;
  assign \new_[56243]_  = ~A169 & \new_[56242]_ ;
  assign \new_[56247]_  = A201 & ~A200;
  assign \new_[56248]_  = A199 & \new_[56247]_ ;
  assign \new_[56249]_  = \new_[56248]_  & \new_[56243]_ ;
  assign \new_[56253]_  = ~A234 & ~A233;
  assign \new_[56254]_  = A203 & \new_[56253]_ ;
  assign \new_[56257]_  = A266 & A265;
  assign \new_[56260]_  = A299 & A298;
  assign \new_[56261]_  = \new_[56260]_  & \new_[56257]_ ;
  assign \new_[56262]_  = \new_[56261]_  & \new_[56254]_ ;
  assign \new_[56266]_  = ~A166 & ~A167;
  assign \new_[56267]_  = ~A169 & \new_[56266]_ ;
  assign \new_[56271]_  = A201 & ~A200;
  assign \new_[56272]_  = A199 & \new_[56271]_ ;
  assign \new_[56273]_  = \new_[56272]_  & \new_[56267]_ ;
  assign \new_[56277]_  = ~A234 & ~A233;
  assign \new_[56278]_  = A203 & \new_[56277]_ ;
  assign \new_[56281]_  = A266 & A265;
  assign \new_[56284]_  = ~A299 & ~A298;
  assign \new_[56285]_  = \new_[56284]_  & \new_[56281]_ ;
  assign \new_[56286]_  = \new_[56285]_  & \new_[56278]_ ;
  assign \new_[56290]_  = ~A166 & ~A167;
  assign \new_[56291]_  = ~A169 & \new_[56290]_ ;
  assign \new_[56295]_  = A201 & ~A200;
  assign \new_[56296]_  = A199 & \new_[56295]_ ;
  assign \new_[56297]_  = \new_[56296]_  & \new_[56291]_ ;
  assign \new_[56301]_  = ~A234 & ~A233;
  assign \new_[56302]_  = A203 & \new_[56301]_ ;
  assign \new_[56305]_  = ~A267 & ~A266;
  assign \new_[56308]_  = ~A300 & A298;
  assign \new_[56309]_  = \new_[56308]_  & \new_[56305]_ ;
  assign \new_[56310]_  = \new_[56309]_  & \new_[56302]_ ;
  assign \new_[56314]_  = ~A166 & ~A167;
  assign \new_[56315]_  = ~A169 & \new_[56314]_ ;
  assign \new_[56319]_  = A201 & ~A200;
  assign \new_[56320]_  = A199 & \new_[56319]_ ;
  assign \new_[56321]_  = \new_[56320]_  & \new_[56315]_ ;
  assign \new_[56325]_  = ~A234 & ~A233;
  assign \new_[56326]_  = A203 & \new_[56325]_ ;
  assign \new_[56329]_  = ~A267 & ~A266;
  assign \new_[56332]_  = A299 & A298;
  assign \new_[56333]_  = \new_[56332]_  & \new_[56329]_ ;
  assign \new_[56334]_  = \new_[56333]_  & \new_[56326]_ ;
  assign \new_[56338]_  = ~A166 & ~A167;
  assign \new_[56339]_  = ~A169 & \new_[56338]_ ;
  assign \new_[56343]_  = A201 & ~A200;
  assign \new_[56344]_  = A199 & \new_[56343]_ ;
  assign \new_[56345]_  = \new_[56344]_  & \new_[56339]_ ;
  assign \new_[56349]_  = ~A234 & ~A233;
  assign \new_[56350]_  = A203 & \new_[56349]_ ;
  assign \new_[56353]_  = ~A267 & ~A266;
  assign \new_[56356]_  = ~A299 & ~A298;
  assign \new_[56357]_  = \new_[56356]_  & \new_[56353]_ ;
  assign \new_[56358]_  = \new_[56357]_  & \new_[56350]_ ;
  assign \new_[56362]_  = ~A166 & ~A167;
  assign \new_[56363]_  = ~A169 & \new_[56362]_ ;
  assign \new_[56367]_  = A201 & ~A200;
  assign \new_[56368]_  = A199 & \new_[56367]_ ;
  assign \new_[56369]_  = \new_[56368]_  & \new_[56363]_ ;
  assign \new_[56373]_  = ~A234 & ~A233;
  assign \new_[56374]_  = A203 & \new_[56373]_ ;
  assign \new_[56377]_  = ~A266 & ~A265;
  assign \new_[56380]_  = ~A300 & A298;
  assign \new_[56381]_  = \new_[56380]_  & \new_[56377]_ ;
  assign \new_[56382]_  = \new_[56381]_  & \new_[56374]_ ;
  assign \new_[56386]_  = ~A166 & ~A167;
  assign \new_[56387]_  = ~A169 & \new_[56386]_ ;
  assign \new_[56391]_  = A201 & ~A200;
  assign \new_[56392]_  = A199 & \new_[56391]_ ;
  assign \new_[56393]_  = \new_[56392]_  & \new_[56387]_ ;
  assign \new_[56397]_  = ~A234 & ~A233;
  assign \new_[56398]_  = A203 & \new_[56397]_ ;
  assign \new_[56401]_  = ~A266 & ~A265;
  assign \new_[56404]_  = A299 & A298;
  assign \new_[56405]_  = \new_[56404]_  & \new_[56401]_ ;
  assign \new_[56406]_  = \new_[56405]_  & \new_[56398]_ ;
  assign \new_[56410]_  = ~A166 & ~A167;
  assign \new_[56411]_  = ~A169 & \new_[56410]_ ;
  assign \new_[56415]_  = A201 & ~A200;
  assign \new_[56416]_  = A199 & \new_[56415]_ ;
  assign \new_[56417]_  = \new_[56416]_  & \new_[56411]_ ;
  assign \new_[56421]_  = ~A234 & ~A233;
  assign \new_[56422]_  = A203 & \new_[56421]_ ;
  assign \new_[56425]_  = ~A266 & ~A265;
  assign \new_[56428]_  = ~A299 & ~A298;
  assign \new_[56429]_  = \new_[56428]_  & \new_[56425]_ ;
  assign \new_[56430]_  = \new_[56429]_  & \new_[56422]_ ;
  assign \new_[56434]_  = ~A166 & ~A167;
  assign \new_[56435]_  = ~A169 & \new_[56434]_ ;
  assign \new_[56439]_  = A201 & ~A200;
  assign \new_[56440]_  = A199 & \new_[56439]_ ;
  assign \new_[56441]_  = \new_[56440]_  & \new_[56435]_ ;
  assign \new_[56445]_  = ~A233 & A232;
  assign \new_[56446]_  = A203 & \new_[56445]_ ;
  assign \new_[56449]_  = A235 & A234;
  assign \new_[56452]_  = A299 & ~A298;
  assign \new_[56453]_  = \new_[56452]_  & \new_[56449]_ ;
  assign \new_[56454]_  = \new_[56453]_  & \new_[56446]_ ;
  assign \new_[56458]_  = ~A166 & ~A167;
  assign \new_[56459]_  = ~A169 & \new_[56458]_ ;
  assign \new_[56463]_  = A201 & ~A200;
  assign \new_[56464]_  = A199 & \new_[56463]_ ;
  assign \new_[56465]_  = \new_[56464]_  & \new_[56459]_ ;
  assign \new_[56469]_  = ~A233 & A232;
  assign \new_[56470]_  = A203 & \new_[56469]_ ;
  assign \new_[56473]_  = A235 & A234;
  assign \new_[56476]_  = A266 & ~A265;
  assign \new_[56477]_  = \new_[56476]_  & \new_[56473]_ ;
  assign \new_[56478]_  = \new_[56477]_  & \new_[56470]_ ;
  assign \new_[56482]_  = ~A166 & ~A167;
  assign \new_[56483]_  = ~A169 & \new_[56482]_ ;
  assign \new_[56487]_  = A201 & ~A200;
  assign \new_[56488]_  = A199 & \new_[56487]_ ;
  assign \new_[56489]_  = \new_[56488]_  & \new_[56483]_ ;
  assign \new_[56493]_  = ~A233 & A232;
  assign \new_[56494]_  = A203 & \new_[56493]_ ;
  assign \new_[56497]_  = A236 & A234;
  assign \new_[56500]_  = A299 & ~A298;
  assign \new_[56501]_  = \new_[56500]_  & \new_[56497]_ ;
  assign \new_[56502]_  = \new_[56501]_  & \new_[56494]_ ;
  assign \new_[56506]_  = ~A166 & ~A167;
  assign \new_[56507]_  = ~A169 & \new_[56506]_ ;
  assign \new_[56511]_  = A201 & ~A200;
  assign \new_[56512]_  = A199 & \new_[56511]_ ;
  assign \new_[56513]_  = \new_[56512]_  & \new_[56507]_ ;
  assign \new_[56517]_  = ~A233 & A232;
  assign \new_[56518]_  = A203 & \new_[56517]_ ;
  assign \new_[56521]_  = A236 & A234;
  assign \new_[56524]_  = A266 & ~A265;
  assign \new_[56525]_  = \new_[56524]_  & \new_[56521]_ ;
  assign \new_[56526]_  = \new_[56525]_  & \new_[56518]_ ;
  assign \new_[56530]_  = ~A166 & ~A167;
  assign \new_[56531]_  = ~A169 & \new_[56530]_ ;
  assign \new_[56535]_  = A201 & ~A200;
  assign \new_[56536]_  = A199 & \new_[56535]_ ;
  assign \new_[56537]_  = \new_[56536]_  & \new_[56531]_ ;
  assign \new_[56541]_  = ~A233 & ~A232;
  assign \new_[56542]_  = A203 & \new_[56541]_ ;
  assign \new_[56545]_  = A266 & A265;
  assign \new_[56548]_  = ~A300 & A298;
  assign \new_[56549]_  = \new_[56548]_  & \new_[56545]_ ;
  assign \new_[56550]_  = \new_[56549]_  & \new_[56542]_ ;
  assign \new_[56554]_  = ~A166 & ~A167;
  assign \new_[56555]_  = ~A169 & \new_[56554]_ ;
  assign \new_[56559]_  = A201 & ~A200;
  assign \new_[56560]_  = A199 & \new_[56559]_ ;
  assign \new_[56561]_  = \new_[56560]_  & \new_[56555]_ ;
  assign \new_[56565]_  = ~A233 & ~A232;
  assign \new_[56566]_  = A203 & \new_[56565]_ ;
  assign \new_[56569]_  = A266 & A265;
  assign \new_[56572]_  = A299 & A298;
  assign \new_[56573]_  = \new_[56572]_  & \new_[56569]_ ;
  assign \new_[56574]_  = \new_[56573]_  & \new_[56566]_ ;
  assign \new_[56578]_  = ~A166 & ~A167;
  assign \new_[56579]_  = ~A169 & \new_[56578]_ ;
  assign \new_[56583]_  = A201 & ~A200;
  assign \new_[56584]_  = A199 & \new_[56583]_ ;
  assign \new_[56585]_  = \new_[56584]_  & \new_[56579]_ ;
  assign \new_[56589]_  = ~A233 & ~A232;
  assign \new_[56590]_  = A203 & \new_[56589]_ ;
  assign \new_[56593]_  = A266 & A265;
  assign \new_[56596]_  = ~A299 & ~A298;
  assign \new_[56597]_  = \new_[56596]_  & \new_[56593]_ ;
  assign \new_[56598]_  = \new_[56597]_  & \new_[56590]_ ;
  assign \new_[56602]_  = ~A166 & ~A167;
  assign \new_[56603]_  = ~A169 & \new_[56602]_ ;
  assign \new_[56607]_  = A201 & ~A200;
  assign \new_[56608]_  = A199 & \new_[56607]_ ;
  assign \new_[56609]_  = \new_[56608]_  & \new_[56603]_ ;
  assign \new_[56613]_  = ~A233 & ~A232;
  assign \new_[56614]_  = A203 & \new_[56613]_ ;
  assign \new_[56617]_  = ~A267 & ~A266;
  assign \new_[56620]_  = ~A300 & A298;
  assign \new_[56621]_  = \new_[56620]_  & \new_[56617]_ ;
  assign \new_[56622]_  = \new_[56621]_  & \new_[56614]_ ;
  assign \new_[56626]_  = ~A166 & ~A167;
  assign \new_[56627]_  = ~A169 & \new_[56626]_ ;
  assign \new_[56631]_  = A201 & ~A200;
  assign \new_[56632]_  = A199 & \new_[56631]_ ;
  assign \new_[56633]_  = \new_[56632]_  & \new_[56627]_ ;
  assign \new_[56637]_  = ~A233 & ~A232;
  assign \new_[56638]_  = A203 & \new_[56637]_ ;
  assign \new_[56641]_  = ~A267 & ~A266;
  assign \new_[56644]_  = A299 & A298;
  assign \new_[56645]_  = \new_[56644]_  & \new_[56641]_ ;
  assign \new_[56646]_  = \new_[56645]_  & \new_[56638]_ ;
  assign \new_[56650]_  = ~A166 & ~A167;
  assign \new_[56651]_  = ~A169 & \new_[56650]_ ;
  assign \new_[56655]_  = A201 & ~A200;
  assign \new_[56656]_  = A199 & \new_[56655]_ ;
  assign \new_[56657]_  = \new_[56656]_  & \new_[56651]_ ;
  assign \new_[56661]_  = ~A233 & ~A232;
  assign \new_[56662]_  = A203 & \new_[56661]_ ;
  assign \new_[56665]_  = ~A267 & ~A266;
  assign \new_[56668]_  = ~A299 & ~A298;
  assign \new_[56669]_  = \new_[56668]_  & \new_[56665]_ ;
  assign \new_[56670]_  = \new_[56669]_  & \new_[56662]_ ;
  assign \new_[56674]_  = ~A166 & ~A167;
  assign \new_[56675]_  = ~A169 & \new_[56674]_ ;
  assign \new_[56679]_  = A201 & ~A200;
  assign \new_[56680]_  = A199 & \new_[56679]_ ;
  assign \new_[56681]_  = \new_[56680]_  & \new_[56675]_ ;
  assign \new_[56685]_  = ~A233 & ~A232;
  assign \new_[56686]_  = A203 & \new_[56685]_ ;
  assign \new_[56689]_  = ~A266 & ~A265;
  assign \new_[56692]_  = ~A300 & A298;
  assign \new_[56693]_  = \new_[56692]_  & \new_[56689]_ ;
  assign \new_[56694]_  = \new_[56693]_  & \new_[56686]_ ;
  assign \new_[56698]_  = ~A166 & ~A167;
  assign \new_[56699]_  = ~A169 & \new_[56698]_ ;
  assign \new_[56703]_  = A201 & ~A200;
  assign \new_[56704]_  = A199 & \new_[56703]_ ;
  assign \new_[56705]_  = \new_[56704]_  & \new_[56699]_ ;
  assign \new_[56709]_  = ~A233 & ~A232;
  assign \new_[56710]_  = A203 & \new_[56709]_ ;
  assign \new_[56713]_  = ~A266 & ~A265;
  assign \new_[56716]_  = A299 & A298;
  assign \new_[56717]_  = \new_[56716]_  & \new_[56713]_ ;
  assign \new_[56718]_  = \new_[56717]_  & \new_[56710]_ ;
  assign \new_[56722]_  = ~A166 & ~A167;
  assign \new_[56723]_  = ~A169 & \new_[56722]_ ;
  assign \new_[56727]_  = A201 & ~A200;
  assign \new_[56728]_  = A199 & \new_[56727]_ ;
  assign \new_[56729]_  = \new_[56728]_  & \new_[56723]_ ;
  assign \new_[56733]_  = ~A233 & ~A232;
  assign \new_[56734]_  = A203 & \new_[56733]_ ;
  assign \new_[56737]_  = ~A266 & ~A265;
  assign \new_[56740]_  = ~A299 & ~A298;
  assign \new_[56741]_  = \new_[56740]_  & \new_[56737]_ ;
  assign \new_[56742]_  = \new_[56741]_  & \new_[56734]_ ;
  assign \new_[56746]_  = A167 & ~A168;
  assign \new_[56747]_  = ~A169 & \new_[56746]_ ;
  assign \new_[56751]_  = A200 & ~A199;
  assign \new_[56752]_  = A166 & \new_[56751]_ ;
  assign \new_[56753]_  = \new_[56752]_  & \new_[56747]_ ;
  assign \new_[56757]_  = A265 & A233;
  assign \new_[56758]_  = A232 & \new_[56757]_ ;
  assign \new_[56761]_  = ~A269 & ~A268;
  assign \new_[56764]_  = ~A300 & ~A299;
  assign \new_[56765]_  = \new_[56764]_  & \new_[56761]_ ;
  assign \new_[56766]_  = \new_[56765]_  & \new_[56758]_ ;
  assign \new_[56770]_  = A167 & ~A168;
  assign \new_[56771]_  = ~A169 & \new_[56770]_ ;
  assign \new_[56775]_  = A200 & ~A199;
  assign \new_[56776]_  = A166 & \new_[56775]_ ;
  assign \new_[56777]_  = \new_[56776]_  & \new_[56771]_ ;
  assign \new_[56781]_  = A265 & A233;
  assign \new_[56782]_  = A232 & \new_[56781]_ ;
  assign \new_[56785]_  = ~A269 & ~A268;
  assign \new_[56788]_  = A299 & A298;
  assign \new_[56789]_  = \new_[56788]_  & \new_[56785]_ ;
  assign \new_[56790]_  = \new_[56789]_  & \new_[56782]_ ;
  assign \new_[56794]_  = A167 & ~A168;
  assign \new_[56795]_  = ~A169 & \new_[56794]_ ;
  assign \new_[56799]_  = A200 & ~A199;
  assign \new_[56800]_  = A166 & \new_[56799]_ ;
  assign \new_[56801]_  = \new_[56800]_  & \new_[56795]_ ;
  assign \new_[56805]_  = A265 & A233;
  assign \new_[56806]_  = A232 & \new_[56805]_ ;
  assign \new_[56809]_  = ~A269 & ~A268;
  assign \new_[56812]_  = ~A299 & ~A298;
  assign \new_[56813]_  = \new_[56812]_  & \new_[56809]_ ;
  assign \new_[56814]_  = \new_[56813]_  & \new_[56806]_ ;
  assign \new_[56818]_  = A167 & ~A168;
  assign \new_[56819]_  = ~A169 & \new_[56818]_ ;
  assign \new_[56823]_  = A200 & ~A199;
  assign \new_[56824]_  = A166 & \new_[56823]_ ;
  assign \new_[56825]_  = \new_[56824]_  & \new_[56819]_ ;
  assign \new_[56829]_  = A265 & A233;
  assign \new_[56830]_  = A232 & \new_[56829]_ ;
  assign \new_[56833]_  = ~A299 & ~A267;
  assign \new_[56836]_  = ~A302 & ~A301;
  assign \new_[56837]_  = \new_[56836]_  & \new_[56833]_ ;
  assign \new_[56838]_  = \new_[56837]_  & \new_[56830]_ ;
  assign \new_[56842]_  = A167 & ~A168;
  assign \new_[56843]_  = ~A169 & \new_[56842]_ ;
  assign \new_[56847]_  = A200 & ~A199;
  assign \new_[56848]_  = A166 & \new_[56847]_ ;
  assign \new_[56849]_  = \new_[56848]_  & \new_[56843]_ ;
  assign \new_[56853]_  = A265 & A233;
  assign \new_[56854]_  = A232 & \new_[56853]_ ;
  assign \new_[56857]_  = ~A299 & A266;
  assign \new_[56860]_  = ~A302 & ~A301;
  assign \new_[56861]_  = \new_[56860]_  & \new_[56857]_ ;
  assign \new_[56862]_  = \new_[56861]_  & \new_[56854]_ ;
  assign \new_[56866]_  = A167 & ~A168;
  assign \new_[56867]_  = ~A169 & \new_[56866]_ ;
  assign \new_[56871]_  = A200 & ~A199;
  assign \new_[56872]_  = A166 & \new_[56871]_ ;
  assign \new_[56873]_  = \new_[56872]_  & \new_[56867]_ ;
  assign \new_[56877]_  = ~A265 & A233;
  assign \new_[56878]_  = A232 & \new_[56877]_ ;
  assign \new_[56881]_  = ~A299 & ~A266;
  assign \new_[56884]_  = ~A302 & ~A301;
  assign \new_[56885]_  = \new_[56884]_  & \new_[56881]_ ;
  assign \new_[56886]_  = \new_[56885]_  & \new_[56878]_ ;
  assign \new_[56890]_  = A167 & ~A168;
  assign \new_[56891]_  = ~A169 & \new_[56890]_ ;
  assign \new_[56895]_  = A200 & ~A199;
  assign \new_[56896]_  = A166 & \new_[56895]_ ;
  assign \new_[56897]_  = \new_[56896]_  & \new_[56891]_ ;
  assign \new_[56901]_  = ~A236 & ~A235;
  assign \new_[56902]_  = ~A233 & \new_[56901]_ ;
  assign \new_[56905]_  = A266 & A265;
  assign \new_[56908]_  = ~A300 & A298;
  assign \new_[56909]_  = \new_[56908]_  & \new_[56905]_ ;
  assign \new_[56910]_  = \new_[56909]_  & \new_[56902]_ ;
  assign \new_[56914]_  = A167 & ~A168;
  assign \new_[56915]_  = ~A169 & \new_[56914]_ ;
  assign \new_[56919]_  = A200 & ~A199;
  assign \new_[56920]_  = A166 & \new_[56919]_ ;
  assign \new_[56921]_  = \new_[56920]_  & \new_[56915]_ ;
  assign \new_[56925]_  = ~A236 & ~A235;
  assign \new_[56926]_  = ~A233 & \new_[56925]_ ;
  assign \new_[56929]_  = A266 & A265;
  assign \new_[56932]_  = A299 & A298;
  assign \new_[56933]_  = \new_[56932]_  & \new_[56929]_ ;
  assign \new_[56934]_  = \new_[56933]_  & \new_[56926]_ ;
  assign \new_[56938]_  = A167 & ~A168;
  assign \new_[56939]_  = ~A169 & \new_[56938]_ ;
  assign \new_[56943]_  = A200 & ~A199;
  assign \new_[56944]_  = A166 & \new_[56943]_ ;
  assign \new_[56945]_  = \new_[56944]_  & \new_[56939]_ ;
  assign \new_[56949]_  = ~A236 & ~A235;
  assign \new_[56950]_  = ~A233 & \new_[56949]_ ;
  assign \new_[56953]_  = A266 & A265;
  assign \new_[56956]_  = ~A299 & ~A298;
  assign \new_[56957]_  = \new_[56956]_  & \new_[56953]_ ;
  assign \new_[56958]_  = \new_[56957]_  & \new_[56950]_ ;
  assign \new_[56962]_  = A167 & ~A168;
  assign \new_[56963]_  = ~A169 & \new_[56962]_ ;
  assign \new_[56967]_  = A200 & ~A199;
  assign \new_[56968]_  = A166 & \new_[56967]_ ;
  assign \new_[56969]_  = \new_[56968]_  & \new_[56963]_ ;
  assign \new_[56973]_  = ~A236 & ~A235;
  assign \new_[56974]_  = ~A233 & \new_[56973]_ ;
  assign \new_[56977]_  = ~A267 & ~A266;
  assign \new_[56980]_  = ~A300 & A298;
  assign \new_[56981]_  = \new_[56980]_  & \new_[56977]_ ;
  assign \new_[56982]_  = \new_[56981]_  & \new_[56974]_ ;
  assign \new_[56986]_  = A167 & ~A168;
  assign \new_[56987]_  = ~A169 & \new_[56986]_ ;
  assign \new_[56991]_  = A200 & ~A199;
  assign \new_[56992]_  = A166 & \new_[56991]_ ;
  assign \new_[56993]_  = \new_[56992]_  & \new_[56987]_ ;
  assign \new_[56997]_  = ~A236 & ~A235;
  assign \new_[56998]_  = ~A233 & \new_[56997]_ ;
  assign \new_[57001]_  = ~A267 & ~A266;
  assign \new_[57004]_  = A299 & A298;
  assign \new_[57005]_  = \new_[57004]_  & \new_[57001]_ ;
  assign \new_[57006]_  = \new_[57005]_  & \new_[56998]_ ;
  assign \new_[57010]_  = A167 & ~A168;
  assign \new_[57011]_  = ~A169 & \new_[57010]_ ;
  assign \new_[57015]_  = A200 & ~A199;
  assign \new_[57016]_  = A166 & \new_[57015]_ ;
  assign \new_[57017]_  = \new_[57016]_  & \new_[57011]_ ;
  assign \new_[57021]_  = ~A236 & ~A235;
  assign \new_[57022]_  = ~A233 & \new_[57021]_ ;
  assign \new_[57025]_  = ~A267 & ~A266;
  assign \new_[57028]_  = ~A299 & ~A298;
  assign \new_[57029]_  = \new_[57028]_  & \new_[57025]_ ;
  assign \new_[57030]_  = \new_[57029]_  & \new_[57022]_ ;
  assign \new_[57034]_  = A167 & ~A168;
  assign \new_[57035]_  = ~A169 & \new_[57034]_ ;
  assign \new_[57039]_  = A200 & ~A199;
  assign \new_[57040]_  = A166 & \new_[57039]_ ;
  assign \new_[57041]_  = \new_[57040]_  & \new_[57035]_ ;
  assign \new_[57045]_  = ~A236 & ~A235;
  assign \new_[57046]_  = ~A233 & \new_[57045]_ ;
  assign \new_[57049]_  = ~A266 & ~A265;
  assign \new_[57052]_  = ~A300 & A298;
  assign \new_[57053]_  = \new_[57052]_  & \new_[57049]_ ;
  assign \new_[57054]_  = \new_[57053]_  & \new_[57046]_ ;
  assign \new_[57058]_  = A167 & ~A168;
  assign \new_[57059]_  = ~A169 & \new_[57058]_ ;
  assign \new_[57063]_  = A200 & ~A199;
  assign \new_[57064]_  = A166 & \new_[57063]_ ;
  assign \new_[57065]_  = \new_[57064]_  & \new_[57059]_ ;
  assign \new_[57069]_  = ~A236 & ~A235;
  assign \new_[57070]_  = ~A233 & \new_[57069]_ ;
  assign \new_[57073]_  = ~A266 & ~A265;
  assign \new_[57076]_  = A299 & A298;
  assign \new_[57077]_  = \new_[57076]_  & \new_[57073]_ ;
  assign \new_[57078]_  = \new_[57077]_  & \new_[57070]_ ;
  assign \new_[57082]_  = A167 & ~A168;
  assign \new_[57083]_  = ~A169 & \new_[57082]_ ;
  assign \new_[57087]_  = A200 & ~A199;
  assign \new_[57088]_  = A166 & \new_[57087]_ ;
  assign \new_[57089]_  = \new_[57088]_  & \new_[57083]_ ;
  assign \new_[57093]_  = ~A236 & ~A235;
  assign \new_[57094]_  = ~A233 & \new_[57093]_ ;
  assign \new_[57097]_  = ~A266 & ~A265;
  assign \new_[57100]_  = ~A299 & ~A298;
  assign \new_[57101]_  = \new_[57100]_  & \new_[57097]_ ;
  assign \new_[57102]_  = \new_[57101]_  & \new_[57094]_ ;
  assign \new_[57106]_  = A167 & ~A168;
  assign \new_[57107]_  = ~A169 & \new_[57106]_ ;
  assign \new_[57111]_  = A200 & ~A199;
  assign \new_[57112]_  = A166 & \new_[57111]_ ;
  assign \new_[57113]_  = \new_[57112]_  & \new_[57107]_ ;
  assign \new_[57117]_  = A265 & ~A234;
  assign \new_[57118]_  = ~A233 & \new_[57117]_ ;
  assign \new_[57121]_  = A298 & A266;
  assign \new_[57124]_  = ~A302 & ~A301;
  assign \new_[57125]_  = \new_[57124]_  & \new_[57121]_ ;
  assign \new_[57126]_  = \new_[57125]_  & \new_[57118]_ ;
  assign \new_[57130]_  = A167 & ~A168;
  assign \new_[57131]_  = ~A169 & \new_[57130]_ ;
  assign \new_[57135]_  = A200 & ~A199;
  assign \new_[57136]_  = A166 & \new_[57135]_ ;
  assign \new_[57137]_  = \new_[57136]_  & \new_[57131]_ ;
  assign \new_[57141]_  = ~A266 & ~A234;
  assign \new_[57142]_  = ~A233 & \new_[57141]_ ;
  assign \new_[57145]_  = ~A269 & ~A268;
  assign \new_[57148]_  = ~A300 & A298;
  assign \new_[57149]_  = \new_[57148]_  & \new_[57145]_ ;
  assign \new_[57150]_  = \new_[57149]_  & \new_[57142]_ ;
  assign \new_[57154]_  = A167 & ~A168;
  assign \new_[57155]_  = ~A169 & \new_[57154]_ ;
  assign \new_[57159]_  = A200 & ~A199;
  assign \new_[57160]_  = A166 & \new_[57159]_ ;
  assign \new_[57161]_  = \new_[57160]_  & \new_[57155]_ ;
  assign \new_[57165]_  = ~A266 & ~A234;
  assign \new_[57166]_  = ~A233 & \new_[57165]_ ;
  assign \new_[57169]_  = ~A269 & ~A268;
  assign \new_[57172]_  = A299 & A298;
  assign \new_[57173]_  = \new_[57172]_  & \new_[57169]_ ;
  assign \new_[57174]_  = \new_[57173]_  & \new_[57166]_ ;
  assign \new_[57178]_  = A167 & ~A168;
  assign \new_[57179]_  = ~A169 & \new_[57178]_ ;
  assign \new_[57183]_  = A200 & ~A199;
  assign \new_[57184]_  = A166 & \new_[57183]_ ;
  assign \new_[57185]_  = \new_[57184]_  & \new_[57179]_ ;
  assign \new_[57189]_  = ~A266 & ~A234;
  assign \new_[57190]_  = ~A233 & \new_[57189]_ ;
  assign \new_[57193]_  = ~A269 & ~A268;
  assign \new_[57196]_  = ~A299 & ~A298;
  assign \new_[57197]_  = \new_[57196]_  & \new_[57193]_ ;
  assign \new_[57198]_  = \new_[57197]_  & \new_[57190]_ ;
  assign \new_[57202]_  = A167 & ~A168;
  assign \new_[57203]_  = ~A169 & \new_[57202]_ ;
  assign \new_[57207]_  = A200 & ~A199;
  assign \new_[57208]_  = A166 & \new_[57207]_ ;
  assign \new_[57209]_  = \new_[57208]_  & \new_[57203]_ ;
  assign \new_[57213]_  = ~A266 & ~A234;
  assign \new_[57214]_  = ~A233 & \new_[57213]_ ;
  assign \new_[57217]_  = A298 & ~A267;
  assign \new_[57220]_  = ~A302 & ~A301;
  assign \new_[57221]_  = \new_[57220]_  & \new_[57217]_ ;
  assign \new_[57222]_  = \new_[57221]_  & \new_[57214]_ ;
  assign \new_[57226]_  = A167 & ~A168;
  assign \new_[57227]_  = ~A169 & \new_[57226]_ ;
  assign \new_[57231]_  = A200 & ~A199;
  assign \new_[57232]_  = A166 & \new_[57231]_ ;
  assign \new_[57233]_  = \new_[57232]_  & \new_[57227]_ ;
  assign \new_[57237]_  = ~A265 & ~A234;
  assign \new_[57238]_  = ~A233 & \new_[57237]_ ;
  assign \new_[57241]_  = A298 & ~A266;
  assign \new_[57244]_  = ~A302 & ~A301;
  assign \new_[57245]_  = \new_[57244]_  & \new_[57241]_ ;
  assign \new_[57246]_  = \new_[57245]_  & \new_[57238]_ ;
  assign \new_[57250]_  = A167 & ~A168;
  assign \new_[57251]_  = ~A169 & \new_[57250]_ ;
  assign \new_[57255]_  = A200 & ~A199;
  assign \new_[57256]_  = A166 & \new_[57255]_ ;
  assign \new_[57257]_  = \new_[57256]_  & \new_[57251]_ ;
  assign \new_[57261]_  = A265 & ~A233;
  assign \new_[57262]_  = ~A232 & \new_[57261]_ ;
  assign \new_[57265]_  = A298 & A266;
  assign \new_[57268]_  = ~A302 & ~A301;
  assign \new_[57269]_  = \new_[57268]_  & \new_[57265]_ ;
  assign \new_[57270]_  = \new_[57269]_  & \new_[57262]_ ;
  assign \new_[57274]_  = A167 & ~A168;
  assign \new_[57275]_  = ~A169 & \new_[57274]_ ;
  assign \new_[57279]_  = A200 & ~A199;
  assign \new_[57280]_  = A166 & \new_[57279]_ ;
  assign \new_[57281]_  = \new_[57280]_  & \new_[57275]_ ;
  assign \new_[57285]_  = ~A266 & ~A233;
  assign \new_[57286]_  = ~A232 & \new_[57285]_ ;
  assign \new_[57289]_  = ~A269 & ~A268;
  assign \new_[57292]_  = ~A300 & A298;
  assign \new_[57293]_  = \new_[57292]_  & \new_[57289]_ ;
  assign \new_[57294]_  = \new_[57293]_  & \new_[57286]_ ;
  assign \new_[57298]_  = A167 & ~A168;
  assign \new_[57299]_  = ~A169 & \new_[57298]_ ;
  assign \new_[57303]_  = A200 & ~A199;
  assign \new_[57304]_  = A166 & \new_[57303]_ ;
  assign \new_[57305]_  = \new_[57304]_  & \new_[57299]_ ;
  assign \new_[57309]_  = ~A266 & ~A233;
  assign \new_[57310]_  = ~A232 & \new_[57309]_ ;
  assign \new_[57313]_  = ~A269 & ~A268;
  assign \new_[57316]_  = A299 & A298;
  assign \new_[57317]_  = \new_[57316]_  & \new_[57313]_ ;
  assign \new_[57318]_  = \new_[57317]_  & \new_[57310]_ ;
  assign \new_[57322]_  = A167 & ~A168;
  assign \new_[57323]_  = ~A169 & \new_[57322]_ ;
  assign \new_[57327]_  = A200 & ~A199;
  assign \new_[57328]_  = A166 & \new_[57327]_ ;
  assign \new_[57329]_  = \new_[57328]_  & \new_[57323]_ ;
  assign \new_[57333]_  = ~A266 & ~A233;
  assign \new_[57334]_  = ~A232 & \new_[57333]_ ;
  assign \new_[57337]_  = ~A269 & ~A268;
  assign \new_[57340]_  = ~A299 & ~A298;
  assign \new_[57341]_  = \new_[57340]_  & \new_[57337]_ ;
  assign \new_[57342]_  = \new_[57341]_  & \new_[57334]_ ;
  assign \new_[57346]_  = A167 & ~A168;
  assign \new_[57347]_  = ~A169 & \new_[57346]_ ;
  assign \new_[57351]_  = A200 & ~A199;
  assign \new_[57352]_  = A166 & \new_[57351]_ ;
  assign \new_[57353]_  = \new_[57352]_  & \new_[57347]_ ;
  assign \new_[57357]_  = ~A266 & ~A233;
  assign \new_[57358]_  = ~A232 & \new_[57357]_ ;
  assign \new_[57361]_  = A298 & ~A267;
  assign \new_[57364]_  = ~A302 & ~A301;
  assign \new_[57365]_  = \new_[57364]_  & \new_[57361]_ ;
  assign \new_[57366]_  = \new_[57365]_  & \new_[57358]_ ;
  assign \new_[57370]_  = A167 & ~A168;
  assign \new_[57371]_  = ~A169 & \new_[57370]_ ;
  assign \new_[57375]_  = A200 & ~A199;
  assign \new_[57376]_  = A166 & \new_[57375]_ ;
  assign \new_[57377]_  = \new_[57376]_  & \new_[57371]_ ;
  assign \new_[57381]_  = ~A265 & ~A233;
  assign \new_[57382]_  = ~A232 & \new_[57381]_ ;
  assign \new_[57385]_  = A298 & ~A266;
  assign \new_[57388]_  = ~A302 & ~A301;
  assign \new_[57389]_  = \new_[57388]_  & \new_[57385]_ ;
  assign \new_[57390]_  = \new_[57389]_  & \new_[57382]_ ;
  assign \new_[57394]_  = A167 & ~A169;
  assign \new_[57395]_  = A170 & \new_[57394]_ ;
  assign \new_[57399]_  = A200 & A199;
  assign \new_[57400]_  = ~A166 & \new_[57399]_ ;
  assign \new_[57401]_  = \new_[57400]_  & \new_[57395]_ ;
  assign \new_[57405]_  = A265 & A233;
  assign \new_[57406]_  = A232 & \new_[57405]_ ;
  assign \new_[57409]_  = ~A269 & ~A268;
  assign \new_[57412]_  = ~A300 & ~A299;
  assign \new_[57413]_  = \new_[57412]_  & \new_[57409]_ ;
  assign \new_[57414]_  = \new_[57413]_  & \new_[57406]_ ;
  assign \new_[57418]_  = A167 & ~A169;
  assign \new_[57419]_  = A170 & \new_[57418]_ ;
  assign \new_[57423]_  = A200 & A199;
  assign \new_[57424]_  = ~A166 & \new_[57423]_ ;
  assign \new_[57425]_  = \new_[57424]_  & \new_[57419]_ ;
  assign \new_[57429]_  = A265 & A233;
  assign \new_[57430]_  = A232 & \new_[57429]_ ;
  assign \new_[57433]_  = ~A269 & ~A268;
  assign \new_[57436]_  = A299 & A298;
  assign \new_[57437]_  = \new_[57436]_  & \new_[57433]_ ;
  assign \new_[57438]_  = \new_[57437]_  & \new_[57430]_ ;
  assign \new_[57442]_  = A167 & ~A169;
  assign \new_[57443]_  = A170 & \new_[57442]_ ;
  assign \new_[57447]_  = A200 & A199;
  assign \new_[57448]_  = ~A166 & \new_[57447]_ ;
  assign \new_[57449]_  = \new_[57448]_  & \new_[57443]_ ;
  assign \new_[57453]_  = A265 & A233;
  assign \new_[57454]_  = A232 & \new_[57453]_ ;
  assign \new_[57457]_  = ~A269 & ~A268;
  assign \new_[57460]_  = ~A299 & ~A298;
  assign \new_[57461]_  = \new_[57460]_  & \new_[57457]_ ;
  assign \new_[57462]_  = \new_[57461]_  & \new_[57454]_ ;
  assign \new_[57466]_  = A167 & ~A169;
  assign \new_[57467]_  = A170 & \new_[57466]_ ;
  assign \new_[57471]_  = A200 & A199;
  assign \new_[57472]_  = ~A166 & \new_[57471]_ ;
  assign \new_[57473]_  = \new_[57472]_  & \new_[57467]_ ;
  assign \new_[57477]_  = A265 & A233;
  assign \new_[57478]_  = A232 & \new_[57477]_ ;
  assign \new_[57481]_  = ~A299 & ~A267;
  assign \new_[57484]_  = ~A302 & ~A301;
  assign \new_[57485]_  = \new_[57484]_  & \new_[57481]_ ;
  assign \new_[57486]_  = \new_[57485]_  & \new_[57478]_ ;
  assign \new_[57490]_  = A167 & ~A169;
  assign \new_[57491]_  = A170 & \new_[57490]_ ;
  assign \new_[57495]_  = A200 & A199;
  assign \new_[57496]_  = ~A166 & \new_[57495]_ ;
  assign \new_[57497]_  = \new_[57496]_  & \new_[57491]_ ;
  assign \new_[57501]_  = A265 & A233;
  assign \new_[57502]_  = A232 & \new_[57501]_ ;
  assign \new_[57505]_  = ~A299 & A266;
  assign \new_[57508]_  = ~A302 & ~A301;
  assign \new_[57509]_  = \new_[57508]_  & \new_[57505]_ ;
  assign \new_[57510]_  = \new_[57509]_  & \new_[57502]_ ;
  assign \new_[57514]_  = A167 & ~A169;
  assign \new_[57515]_  = A170 & \new_[57514]_ ;
  assign \new_[57519]_  = A200 & A199;
  assign \new_[57520]_  = ~A166 & \new_[57519]_ ;
  assign \new_[57521]_  = \new_[57520]_  & \new_[57515]_ ;
  assign \new_[57525]_  = ~A265 & A233;
  assign \new_[57526]_  = A232 & \new_[57525]_ ;
  assign \new_[57529]_  = ~A299 & ~A266;
  assign \new_[57532]_  = ~A302 & ~A301;
  assign \new_[57533]_  = \new_[57532]_  & \new_[57529]_ ;
  assign \new_[57534]_  = \new_[57533]_  & \new_[57526]_ ;
  assign \new_[57538]_  = A167 & ~A169;
  assign \new_[57539]_  = A170 & \new_[57538]_ ;
  assign \new_[57543]_  = A200 & A199;
  assign \new_[57544]_  = ~A166 & \new_[57543]_ ;
  assign \new_[57545]_  = \new_[57544]_  & \new_[57539]_ ;
  assign \new_[57549]_  = ~A236 & ~A235;
  assign \new_[57550]_  = ~A233 & \new_[57549]_ ;
  assign \new_[57553]_  = A266 & A265;
  assign \new_[57556]_  = ~A300 & A298;
  assign \new_[57557]_  = \new_[57556]_  & \new_[57553]_ ;
  assign \new_[57558]_  = \new_[57557]_  & \new_[57550]_ ;
  assign \new_[57562]_  = A167 & ~A169;
  assign \new_[57563]_  = A170 & \new_[57562]_ ;
  assign \new_[57567]_  = A200 & A199;
  assign \new_[57568]_  = ~A166 & \new_[57567]_ ;
  assign \new_[57569]_  = \new_[57568]_  & \new_[57563]_ ;
  assign \new_[57573]_  = ~A236 & ~A235;
  assign \new_[57574]_  = ~A233 & \new_[57573]_ ;
  assign \new_[57577]_  = A266 & A265;
  assign \new_[57580]_  = A299 & A298;
  assign \new_[57581]_  = \new_[57580]_  & \new_[57577]_ ;
  assign \new_[57582]_  = \new_[57581]_  & \new_[57574]_ ;
  assign \new_[57586]_  = A167 & ~A169;
  assign \new_[57587]_  = A170 & \new_[57586]_ ;
  assign \new_[57591]_  = A200 & A199;
  assign \new_[57592]_  = ~A166 & \new_[57591]_ ;
  assign \new_[57593]_  = \new_[57592]_  & \new_[57587]_ ;
  assign \new_[57597]_  = ~A236 & ~A235;
  assign \new_[57598]_  = ~A233 & \new_[57597]_ ;
  assign \new_[57601]_  = A266 & A265;
  assign \new_[57604]_  = ~A299 & ~A298;
  assign \new_[57605]_  = \new_[57604]_  & \new_[57601]_ ;
  assign \new_[57606]_  = \new_[57605]_  & \new_[57598]_ ;
  assign \new_[57610]_  = A167 & ~A169;
  assign \new_[57611]_  = A170 & \new_[57610]_ ;
  assign \new_[57615]_  = A200 & A199;
  assign \new_[57616]_  = ~A166 & \new_[57615]_ ;
  assign \new_[57617]_  = \new_[57616]_  & \new_[57611]_ ;
  assign \new_[57621]_  = ~A236 & ~A235;
  assign \new_[57622]_  = ~A233 & \new_[57621]_ ;
  assign \new_[57625]_  = ~A267 & ~A266;
  assign \new_[57628]_  = ~A300 & A298;
  assign \new_[57629]_  = \new_[57628]_  & \new_[57625]_ ;
  assign \new_[57630]_  = \new_[57629]_  & \new_[57622]_ ;
  assign \new_[57634]_  = A167 & ~A169;
  assign \new_[57635]_  = A170 & \new_[57634]_ ;
  assign \new_[57639]_  = A200 & A199;
  assign \new_[57640]_  = ~A166 & \new_[57639]_ ;
  assign \new_[57641]_  = \new_[57640]_  & \new_[57635]_ ;
  assign \new_[57645]_  = ~A236 & ~A235;
  assign \new_[57646]_  = ~A233 & \new_[57645]_ ;
  assign \new_[57649]_  = ~A267 & ~A266;
  assign \new_[57652]_  = A299 & A298;
  assign \new_[57653]_  = \new_[57652]_  & \new_[57649]_ ;
  assign \new_[57654]_  = \new_[57653]_  & \new_[57646]_ ;
  assign \new_[57658]_  = A167 & ~A169;
  assign \new_[57659]_  = A170 & \new_[57658]_ ;
  assign \new_[57663]_  = A200 & A199;
  assign \new_[57664]_  = ~A166 & \new_[57663]_ ;
  assign \new_[57665]_  = \new_[57664]_  & \new_[57659]_ ;
  assign \new_[57669]_  = ~A236 & ~A235;
  assign \new_[57670]_  = ~A233 & \new_[57669]_ ;
  assign \new_[57673]_  = ~A267 & ~A266;
  assign \new_[57676]_  = ~A299 & ~A298;
  assign \new_[57677]_  = \new_[57676]_  & \new_[57673]_ ;
  assign \new_[57678]_  = \new_[57677]_  & \new_[57670]_ ;
  assign \new_[57682]_  = A167 & ~A169;
  assign \new_[57683]_  = A170 & \new_[57682]_ ;
  assign \new_[57687]_  = A200 & A199;
  assign \new_[57688]_  = ~A166 & \new_[57687]_ ;
  assign \new_[57689]_  = \new_[57688]_  & \new_[57683]_ ;
  assign \new_[57693]_  = ~A236 & ~A235;
  assign \new_[57694]_  = ~A233 & \new_[57693]_ ;
  assign \new_[57697]_  = ~A266 & ~A265;
  assign \new_[57700]_  = ~A300 & A298;
  assign \new_[57701]_  = \new_[57700]_  & \new_[57697]_ ;
  assign \new_[57702]_  = \new_[57701]_  & \new_[57694]_ ;
  assign \new_[57706]_  = A167 & ~A169;
  assign \new_[57707]_  = A170 & \new_[57706]_ ;
  assign \new_[57711]_  = A200 & A199;
  assign \new_[57712]_  = ~A166 & \new_[57711]_ ;
  assign \new_[57713]_  = \new_[57712]_  & \new_[57707]_ ;
  assign \new_[57717]_  = ~A236 & ~A235;
  assign \new_[57718]_  = ~A233 & \new_[57717]_ ;
  assign \new_[57721]_  = ~A266 & ~A265;
  assign \new_[57724]_  = A299 & A298;
  assign \new_[57725]_  = \new_[57724]_  & \new_[57721]_ ;
  assign \new_[57726]_  = \new_[57725]_  & \new_[57718]_ ;
  assign \new_[57730]_  = A167 & ~A169;
  assign \new_[57731]_  = A170 & \new_[57730]_ ;
  assign \new_[57735]_  = A200 & A199;
  assign \new_[57736]_  = ~A166 & \new_[57735]_ ;
  assign \new_[57737]_  = \new_[57736]_  & \new_[57731]_ ;
  assign \new_[57741]_  = ~A236 & ~A235;
  assign \new_[57742]_  = ~A233 & \new_[57741]_ ;
  assign \new_[57745]_  = ~A266 & ~A265;
  assign \new_[57748]_  = ~A299 & ~A298;
  assign \new_[57749]_  = \new_[57748]_  & \new_[57745]_ ;
  assign \new_[57750]_  = \new_[57749]_  & \new_[57742]_ ;
  assign \new_[57754]_  = A167 & ~A169;
  assign \new_[57755]_  = A170 & \new_[57754]_ ;
  assign \new_[57759]_  = A200 & A199;
  assign \new_[57760]_  = ~A166 & \new_[57759]_ ;
  assign \new_[57761]_  = \new_[57760]_  & \new_[57755]_ ;
  assign \new_[57765]_  = A265 & ~A234;
  assign \new_[57766]_  = ~A233 & \new_[57765]_ ;
  assign \new_[57769]_  = A298 & A266;
  assign \new_[57772]_  = ~A302 & ~A301;
  assign \new_[57773]_  = \new_[57772]_  & \new_[57769]_ ;
  assign \new_[57774]_  = \new_[57773]_  & \new_[57766]_ ;
  assign \new_[57778]_  = A167 & ~A169;
  assign \new_[57779]_  = A170 & \new_[57778]_ ;
  assign \new_[57783]_  = A200 & A199;
  assign \new_[57784]_  = ~A166 & \new_[57783]_ ;
  assign \new_[57785]_  = \new_[57784]_  & \new_[57779]_ ;
  assign \new_[57789]_  = ~A266 & ~A234;
  assign \new_[57790]_  = ~A233 & \new_[57789]_ ;
  assign \new_[57793]_  = ~A269 & ~A268;
  assign \new_[57796]_  = ~A300 & A298;
  assign \new_[57797]_  = \new_[57796]_  & \new_[57793]_ ;
  assign \new_[57798]_  = \new_[57797]_  & \new_[57790]_ ;
  assign \new_[57802]_  = A167 & ~A169;
  assign \new_[57803]_  = A170 & \new_[57802]_ ;
  assign \new_[57807]_  = A200 & A199;
  assign \new_[57808]_  = ~A166 & \new_[57807]_ ;
  assign \new_[57809]_  = \new_[57808]_  & \new_[57803]_ ;
  assign \new_[57813]_  = ~A266 & ~A234;
  assign \new_[57814]_  = ~A233 & \new_[57813]_ ;
  assign \new_[57817]_  = ~A269 & ~A268;
  assign \new_[57820]_  = A299 & A298;
  assign \new_[57821]_  = \new_[57820]_  & \new_[57817]_ ;
  assign \new_[57822]_  = \new_[57821]_  & \new_[57814]_ ;
  assign \new_[57826]_  = A167 & ~A169;
  assign \new_[57827]_  = A170 & \new_[57826]_ ;
  assign \new_[57831]_  = A200 & A199;
  assign \new_[57832]_  = ~A166 & \new_[57831]_ ;
  assign \new_[57833]_  = \new_[57832]_  & \new_[57827]_ ;
  assign \new_[57837]_  = ~A266 & ~A234;
  assign \new_[57838]_  = ~A233 & \new_[57837]_ ;
  assign \new_[57841]_  = ~A269 & ~A268;
  assign \new_[57844]_  = ~A299 & ~A298;
  assign \new_[57845]_  = \new_[57844]_  & \new_[57841]_ ;
  assign \new_[57846]_  = \new_[57845]_  & \new_[57838]_ ;
  assign \new_[57850]_  = A167 & ~A169;
  assign \new_[57851]_  = A170 & \new_[57850]_ ;
  assign \new_[57855]_  = A200 & A199;
  assign \new_[57856]_  = ~A166 & \new_[57855]_ ;
  assign \new_[57857]_  = \new_[57856]_  & \new_[57851]_ ;
  assign \new_[57861]_  = ~A266 & ~A234;
  assign \new_[57862]_  = ~A233 & \new_[57861]_ ;
  assign \new_[57865]_  = A298 & ~A267;
  assign \new_[57868]_  = ~A302 & ~A301;
  assign \new_[57869]_  = \new_[57868]_  & \new_[57865]_ ;
  assign \new_[57870]_  = \new_[57869]_  & \new_[57862]_ ;
  assign \new_[57874]_  = A167 & ~A169;
  assign \new_[57875]_  = A170 & \new_[57874]_ ;
  assign \new_[57879]_  = A200 & A199;
  assign \new_[57880]_  = ~A166 & \new_[57879]_ ;
  assign \new_[57881]_  = \new_[57880]_  & \new_[57875]_ ;
  assign \new_[57885]_  = ~A265 & ~A234;
  assign \new_[57886]_  = ~A233 & \new_[57885]_ ;
  assign \new_[57889]_  = A298 & ~A266;
  assign \new_[57892]_  = ~A302 & ~A301;
  assign \new_[57893]_  = \new_[57892]_  & \new_[57889]_ ;
  assign \new_[57894]_  = \new_[57893]_  & \new_[57886]_ ;
  assign \new_[57898]_  = A167 & ~A169;
  assign \new_[57899]_  = A170 & \new_[57898]_ ;
  assign \new_[57903]_  = A200 & A199;
  assign \new_[57904]_  = ~A166 & \new_[57903]_ ;
  assign \new_[57905]_  = \new_[57904]_  & \new_[57899]_ ;
  assign \new_[57909]_  = A265 & ~A233;
  assign \new_[57910]_  = ~A232 & \new_[57909]_ ;
  assign \new_[57913]_  = A298 & A266;
  assign \new_[57916]_  = ~A302 & ~A301;
  assign \new_[57917]_  = \new_[57916]_  & \new_[57913]_ ;
  assign \new_[57918]_  = \new_[57917]_  & \new_[57910]_ ;
  assign \new_[57922]_  = A167 & ~A169;
  assign \new_[57923]_  = A170 & \new_[57922]_ ;
  assign \new_[57927]_  = A200 & A199;
  assign \new_[57928]_  = ~A166 & \new_[57927]_ ;
  assign \new_[57929]_  = \new_[57928]_  & \new_[57923]_ ;
  assign \new_[57933]_  = ~A266 & ~A233;
  assign \new_[57934]_  = ~A232 & \new_[57933]_ ;
  assign \new_[57937]_  = ~A269 & ~A268;
  assign \new_[57940]_  = ~A300 & A298;
  assign \new_[57941]_  = \new_[57940]_  & \new_[57937]_ ;
  assign \new_[57942]_  = \new_[57941]_  & \new_[57934]_ ;
  assign \new_[57946]_  = A167 & ~A169;
  assign \new_[57947]_  = A170 & \new_[57946]_ ;
  assign \new_[57951]_  = A200 & A199;
  assign \new_[57952]_  = ~A166 & \new_[57951]_ ;
  assign \new_[57953]_  = \new_[57952]_  & \new_[57947]_ ;
  assign \new_[57957]_  = ~A266 & ~A233;
  assign \new_[57958]_  = ~A232 & \new_[57957]_ ;
  assign \new_[57961]_  = ~A269 & ~A268;
  assign \new_[57964]_  = A299 & A298;
  assign \new_[57965]_  = \new_[57964]_  & \new_[57961]_ ;
  assign \new_[57966]_  = \new_[57965]_  & \new_[57958]_ ;
  assign \new_[57970]_  = A167 & ~A169;
  assign \new_[57971]_  = A170 & \new_[57970]_ ;
  assign \new_[57975]_  = A200 & A199;
  assign \new_[57976]_  = ~A166 & \new_[57975]_ ;
  assign \new_[57977]_  = \new_[57976]_  & \new_[57971]_ ;
  assign \new_[57981]_  = ~A266 & ~A233;
  assign \new_[57982]_  = ~A232 & \new_[57981]_ ;
  assign \new_[57985]_  = ~A269 & ~A268;
  assign \new_[57988]_  = ~A299 & ~A298;
  assign \new_[57989]_  = \new_[57988]_  & \new_[57985]_ ;
  assign \new_[57990]_  = \new_[57989]_  & \new_[57982]_ ;
  assign \new_[57994]_  = A167 & ~A169;
  assign \new_[57995]_  = A170 & \new_[57994]_ ;
  assign \new_[57999]_  = A200 & A199;
  assign \new_[58000]_  = ~A166 & \new_[57999]_ ;
  assign \new_[58001]_  = \new_[58000]_  & \new_[57995]_ ;
  assign \new_[58005]_  = ~A266 & ~A233;
  assign \new_[58006]_  = ~A232 & \new_[58005]_ ;
  assign \new_[58009]_  = A298 & ~A267;
  assign \new_[58012]_  = ~A302 & ~A301;
  assign \new_[58013]_  = \new_[58012]_  & \new_[58009]_ ;
  assign \new_[58014]_  = \new_[58013]_  & \new_[58006]_ ;
  assign \new_[58018]_  = A167 & ~A169;
  assign \new_[58019]_  = A170 & \new_[58018]_ ;
  assign \new_[58023]_  = A200 & A199;
  assign \new_[58024]_  = ~A166 & \new_[58023]_ ;
  assign \new_[58025]_  = \new_[58024]_  & \new_[58019]_ ;
  assign \new_[58029]_  = ~A265 & ~A233;
  assign \new_[58030]_  = ~A232 & \new_[58029]_ ;
  assign \new_[58033]_  = A298 & ~A266;
  assign \new_[58036]_  = ~A302 & ~A301;
  assign \new_[58037]_  = \new_[58036]_  & \new_[58033]_ ;
  assign \new_[58038]_  = \new_[58037]_  & \new_[58030]_ ;
  assign \new_[58042]_  = A167 & ~A169;
  assign \new_[58043]_  = A170 & \new_[58042]_ ;
  assign \new_[58047]_  = ~A202 & ~A200;
  assign \new_[58048]_  = ~A166 & \new_[58047]_ ;
  assign \new_[58049]_  = \new_[58048]_  & \new_[58043]_ ;
  assign \new_[58053]_  = A233 & A232;
  assign \new_[58054]_  = ~A203 & \new_[58053]_ ;
  assign \new_[58057]_  = ~A267 & A265;
  assign \new_[58060]_  = ~A300 & ~A299;
  assign \new_[58061]_  = \new_[58060]_  & \new_[58057]_ ;
  assign \new_[58062]_  = \new_[58061]_  & \new_[58054]_ ;
  assign \new_[58066]_  = A167 & ~A169;
  assign \new_[58067]_  = A170 & \new_[58066]_ ;
  assign \new_[58071]_  = ~A202 & ~A200;
  assign \new_[58072]_  = ~A166 & \new_[58071]_ ;
  assign \new_[58073]_  = \new_[58072]_  & \new_[58067]_ ;
  assign \new_[58077]_  = A233 & A232;
  assign \new_[58078]_  = ~A203 & \new_[58077]_ ;
  assign \new_[58081]_  = ~A267 & A265;
  assign \new_[58084]_  = A299 & A298;
  assign \new_[58085]_  = \new_[58084]_  & \new_[58081]_ ;
  assign \new_[58086]_  = \new_[58085]_  & \new_[58078]_ ;
  assign \new_[58090]_  = A167 & ~A169;
  assign \new_[58091]_  = A170 & \new_[58090]_ ;
  assign \new_[58095]_  = ~A202 & ~A200;
  assign \new_[58096]_  = ~A166 & \new_[58095]_ ;
  assign \new_[58097]_  = \new_[58096]_  & \new_[58091]_ ;
  assign \new_[58101]_  = A233 & A232;
  assign \new_[58102]_  = ~A203 & \new_[58101]_ ;
  assign \new_[58105]_  = ~A267 & A265;
  assign \new_[58108]_  = ~A299 & ~A298;
  assign \new_[58109]_  = \new_[58108]_  & \new_[58105]_ ;
  assign \new_[58110]_  = \new_[58109]_  & \new_[58102]_ ;
  assign \new_[58114]_  = A167 & ~A169;
  assign \new_[58115]_  = A170 & \new_[58114]_ ;
  assign \new_[58119]_  = ~A202 & ~A200;
  assign \new_[58120]_  = ~A166 & \new_[58119]_ ;
  assign \new_[58121]_  = \new_[58120]_  & \new_[58115]_ ;
  assign \new_[58125]_  = A233 & A232;
  assign \new_[58126]_  = ~A203 & \new_[58125]_ ;
  assign \new_[58129]_  = A266 & A265;
  assign \new_[58132]_  = ~A300 & ~A299;
  assign \new_[58133]_  = \new_[58132]_  & \new_[58129]_ ;
  assign \new_[58134]_  = \new_[58133]_  & \new_[58126]_ ;
  assign \new_[58138]_  = A167 & ~A169;
  assign \new_[58139]_  = A170 & \new_[58138]_ ;
  assign \new_[58143]_  = ~A202 & ~A200;
  assign \new_[58144]_  = ~A166 & \new_[58143]_ ;
  assign \new_[58145]_  = \new_[58144]_  & \new_[58139]_ ;
  assign \new_[58149]_  = A233 & A232;
  assign \new_[58150]_  = ~A203 & \new_[58149]_ ;
  assign \new_[58153]_  = A266 & A265;
  assign \new_[58156]_  = A299 & A298;
  assign \new_[58157]_  = \new_[58156]_  & \new_[58153]_ ;
  assign \new_[58158]_  = \new_[58157]_  & \new_[58150]_ ;
  assign \new_[58162]_  = A167 & ~A169;
  assign \new_[58163]_  = A170 & \new_[58162]_ ;
  assign \new_[58167]_  = ~A202 & ~A200;
  assign \new_[58168]_  = ~A166 & \new_[58167]_ ;
  assign \new_[58169]_  = \new_[58168]_  & \new_[58163]_ ;
  assign \new_[58173]_  = A233 & A232;
  assign \new_[58174]_  = ~A203 & \new_[58173]_ ;
  assign \new_[58177]_  = A266 & A265;
  assign \new_[58180]_  = ~A299 & ~A298;
  assign \new_[58181]_  = \new_[58180]_  & \new_[58177]_ ;
  assign \new_[58182]_  = \new_[58181]_  & \new_[58174]_ ;
  assign \new_[58186]_  = A167 & ~A169;
  assign \new_[58187]_  = A170 & \new_[58186]_ ;
  assign \new_[58191]_  = ~A202 & ~A200;
  assign \new_[58192]_  = ~A166 & \new_[58191]_ ;
  assign \new_[58193]_  = \new_[58192]_  & \new_[58187]_ ;
  assign \new_[58197]_  = A233 & A232;
  assign \new_[58198]_  = ~A203 & \new_[58197]_ ;
  assign \new_[58201]_  = ~A266 & ~A265;
  assign \new_[58204]_  = ~A300 & ~A299;
  assign \new_[58205]_  = \new_[58204]_  & \new_[58201]_ ;
  assign \new_[58206]_  = \new_[58205]_  & \new_[58198]_ ;
  assign \new_[58210]_  = A167 & ~A169;
  assign \new_[58211]_  = A170 & \new_[58210]_ ;
  assign \new_[58215]_  = ~A202 & ~A200;
  assign \new_[58216]_  = ~A166 & \new_[58215]_ ;
  assign \new_[58217]_  = \new_[58216]_  & \new_[58211]_ ;
  assign \new_[58221]_  = A233 & A232;
  assign \new_[58222]_  = ~A203 & \new_[58221]_ ;
  assign \new_[58225]_  = ~A266 & ~A265;
  assign \new_[58228]_  = A299 & A298;
  assign \new_[58229]_  = \new_[58228]_  & \new_[58225]_ ;
  assign \new_[58230]_  = \new_[58229]_  & \new_[58222]_ ;
  assign \new_[58234]_  = A167 & ~A169;
  assign \new_[58235]_  = A170 & \new_[58234]_ ;
  assign \new_[58239]_  = ~A202 & ~A200;
  assign \new_[58240]_  = ~A166 & \new_[58239]_ ;
  assign \new_[58241]_  = \new_[58240]_  & \new_[58235]_ ;
  assign \new_[58245]_  = A233 & A232;
  assign \new_[58246]_  = ~A203 & \new_[58245]_ ;
  assign \new_[58249]_  = ~A266 & ~A265;
  assign \new_[58252]_  = ~A299 & ~A298;
  assign \new_[58253]_  = \new_[58252]_  & \new_[58249]_ ;
  assign \new_[58254]_  = \new_[58253]_  & \new_[58246]_ ;
  assign \new_[58258]_  = A167 & ~A169;
  assign \new_[58259]_  = A170 & \new_[58258]_ ;
  assign \new_[58263]_  = ~A202 & ~A200;
  assign \new_[58264]_  = ~A166 & \new_[58263]_ ;
  assign \new_[58265]_  = \new_[58264]_  & \new_[58259]_ ;
  assign \new_[58269]_  = A233 & ~A232;
  assign \new_[58270]_  = ~A203 & \new_[58269]_ ;
  assign \new_[58273]_  = ~A299 & A298;
  assign \new_[58276]_  = A301 & A300;
  assign \new_[58277]_  = \new_[58276]_  & \new_[58273]_ ;
  assign \new_[58278]_  = \new_[58277]_  & \new_[58270]_ ;
  assign \new_[58282]_  = A167 & ~A169;
  assign \new_[58283]_  = A170 & \new_[58282]_ ;
  assign \new_[58287]_  = ~A202 & ~A200;
  assign \new_[58288]_  = ~A166 & \new_[58287]_ ;
  assign \new_[58289]_  = \new_[58288]_  & \new_[58283]_ ;
  assign \new_[58293]_  = A233 & ~A232;
  assign \new_[58294]_  = ~A203 & \new_[58293]_ ;
  assign \new_[58297]_  = ~A299 & A298;
  assign \new_[58300]_  = A302 & A300;
  assign \new_[58301]_  = \new_[58300]_  & \new_[58297]_ ;
  assign \new_[58302]_  = \new_[58301]_  & \new_[58294]_ ;
  assign \new_[58306]_  = A167 & ~A169;
  assign \new_[58307]_  = A170 & \new_[58306]_ ;
  assign \new_[58311]_  = ~A202 & ~A200;
  assign \new_[58312]_  = ~A166 & \new_[58311]_ ;
  assign \new_[58313]_  = \new_[58312]_  & \new_[58307]_ ;
  assign \new_[58317]_  = A233 & ~A232;
  assign \new_[58318]_  = ~A203 & \new_[58317]_ ;
  assign \new_[58321]_  = ~A266 & A265;
  assign \new_[58324]_  = A268 & A267;
  assign \new_[58325]_  = \new_[58324]_  & \new_[58321]_ ;
  assign \new_[58326]_  = \new_[58325]_  & \new_[58318]_ ;
  assign \new_[58330]_  = A167 & ~A169;
  assign \new_[58331]_  = A170 & \new_[58330]_ ;
  assign \new_[58335]_  = ~A202 & ~A200;
  assign \new_[58336]_  = ~A166 & \new_[58335]_ ;
  assign \new_[58337]_  = \new_[58336]_  & \new_[58331]_ ;
  assign \new_[58341]_  = A233 & ~A232;
  assign \new_[58342]_  = ~A203 & \new_[58341]_ ;
  assign \new_[58345]_  = ~A266 & A265;
  assign \new_[58348]_  = A269 & A267;
  assign \new_[58349]_  = \new_[58348]_  & \new_[58345]_ ;
  assign \new_[58350]_  = \new_[58349]_  & \new_[58342]_ ;
  assign \new_[58354]_  = A167 & ~A169;
  assign \new_[58355]_  = A170 & \new_[58354]_ ;
  assign \new_[58359]_  = ~A202 & ~A200;
  assign \new_[58360]_  = ~A166 & \new_[58359]_ ;
  assign \new_[58361]_  = \new_[58360]_  & \new_[58355]_ ;
  assign \new_[58365]_  = ~A234 & ~A233;
  assign \new_[58366]_  = ~A203 & \new_[58365]_ ;
  assign \new_[58369]_  = A266 & A265;
  assign \new_[58372]_  = ~A300 & A298;
  assign \new_[58373]_  = \new_[58372]_  & \new_[58369]_ ;
  assign \new_[58374]_  = \new_[58373]_  & \new_[58366]_ ;
  assign \new_[58378]_  = A167 & ~A169;
  assign \new_[58379]_  = A170 & \new_[58378]_ ;
  assign \new_[58383]_  = ~A202 & ~A200;
  assign \new_[58384]_  = ~A166 & \new_[58383]_ ;
  assign \new_[58385]_  = \new_[58384]_  & \new_[58379]_ ;
  assign \new_[58389]_  = ~A234 & ~A233;
  assign \new_[58390]_  = ~A203 & \new_[58389]_ ;
  assign \new_[58393]_  = A266 & A265;
  assign \new_[58396]_  = A299 & A298;
  assign \new_[58397]_  = \new_[58396]_  & \new_[58393]_ ;
  assign \new_[58398]_  = \new_[58397]_  & \new_[58390]_ ;
  assign \new_[58402]_  = A167 & ~A169;
  assign \new_[58403]_  = A170 & \new_[58402]_ ;
  assign \new_[58407]_  = ~A202 & ~A200;
  assign \new_[58408]_  = ~A166 & \new_[58407]_ ;
  assign \new_[58409]_  = \new_[58408]_  & \new_[58403]_ ;
  assign \new_[58413]_  = ~A234 & ~A233;
  assign \new_[58414]_  = ~A203 & \new_[58413]_ ;
  assign \new_[58417]_  = A266 & A265;
  assign \new_[58420]_  = ~A299 & ~A298;
  assign \new_[58421]_  = \new_[58420]_  & \new_[58417]_ ;
  assign \new_[58422]_  = \new_[58421]_  & \new_[58414]_ ;
  assign \new_[58426]_  = A167 & ~A169;
  assign \new_[58427]_  = A170 & \new_[58426]_ ;
  assign \new_[58431]_  = ~A202 & ~A200;
  assign \new_[58432]_  = ~A166 & \new_[58431]_ ;
  assign \new_[58433]_  = \new_[58432]_  & \new_[58427]_ ;
  assign \new_[58437]_  = ~A234 & ~A233;
  assign \new_[58438]_  = ~A203 & \new_[58437]_ ;
  assign \new_[58441]_  = ~A267 & ~A266;
  assign \new_[58444]_  = ~A300 & A298;
  assign \new_[58445]_  = \new_[58444]_  & \new_[58441]_ ;
  assign \new_[58446]_  = \new_[58445]_  & \new_[58438]_ ;
  assign \new_[58450]_  = A167 & ~A169;
  assign \new_[58451]_  = A170 & \new_[58450]_ ;
  assign \new_[58455]_  = ~A202 & ~A200;
  assign \new_[58456]_  = ~A166 & \new_[58455]_ ;
  assign \new_[58457]_  = \new_[58456]_  & \new_[58451]_ ;
  assign \new_[58461]_  = ~A234 & ~A233;
  assign \new_[58462]_  = ~A203 & \new_[58461]_ ;
  assign \new_[58465]_  = ~A267 & ~A266;
  assign \new_[58468]_  = A299 & A298;
  assign \new_[58469]_  = \new_[58468]_  & \new_[58465]_ ;
  assign \new_[58470]_  = \new_[58469]_  & \new_[58462]_ ;
  assign \new_[58474]_  = A167 & ~A169;
  assign \new_[58475]_  = A170 & \new_[58474]_ ;
  assign \new_[58479]_  = ~A202 & ~A200;
  assign \new_[58480]_  = ~A166 & \new_[58479]_ ;
  assign \new_[58481]_  = \new_[58480]_  & \new_[58475]_ ;
  assign \new_[58485]_  = ~A234 & ~A233;
  assign \new_[58486]_  = ~A203 & \new_[58485]_ ;
  assign \new_[58489]_  = ~A267 & ~A266;
  assign \new_[58492]_  = ~A299 & ~A298;
  assign \new_[58493]_  = \new_[58492]_  & \new_[58489]_ ;
  assign \new_[58494]_  = \new_[58493]_  & \new_[58486]_ ;
  assign \new_[58498]_  = A167 & ~A169;
  assign \new_[58499]_  = A170 & \new_[58498]_ ;
  assign \new_[58503]_  = ~A202 & ~A200;
  assign \new_[58504]_  = ~A166 & \new_[58503]_ ;
  assign \new_[58505]_  = \new_[58504]_  & \new_[58499]_ ;
  assign \new_[58509]_  = ~A234 & ~A233;
  assign \new_[58510]_  = ~A203 & \new_[58509]_ ;
  assign \new_[58513]_  = ~A266 & ~A265;
  assign \new_[58516]_  = ~A300 & A298;
  assign \new_[58517]_  = \new_[58516]_  & \new_[58513]_ ;
  assign \new_[58518]_  = \new_[58517]_  & \new_[58510]_ ;
  assign \new_[58522]_  = A167 & ~A169;
  assign \new_[58523]_  = A170 & \new_[58522]_ ;
  assign \new_[58527]_  = ~A202 & ~A200;
  assign \new_[58528]_  = ~A166 & \new_[58527]_ ;
  assign \new_[58529]_  = \new_[58528]_  & \new_[58523]_ ;
  assign \new_[58533]_  = ~A234 & ~A233;
  assign \new_[58534]_  = ~A203 & \new_[58533]_ ;
  assign \new_[58537]_  = ~A266 & ~A265;
  assign \new_[58540]_  = A299 & A298;
  assign \new_[58541]_  = \new_[58540]_  & \new_[58537]_ ;
  assign \new_[58542]_  = \new_[58541]_  & \new_[58534]_ ;
  assign \new_[58546]_  = A167 & ~A169;
  assign \new_[58547]_  = A170 & \new_[58546]_ ;
  assign \new_[58551]_  = ~A202 & ~A200;
  assign \new_[58552]_  = ~A166 & \new_[58551]_ ;
  assign \new_[58553]_  = \new_[58552]_  & \new_[58547]_ ;
  assign \new_[58557]_  = ~A234 & ~A233;
  assign \new_[58558]_  = ~A203 & \new_[58557]_ ;
  assign \new_[58561]_  = ~A266 & ~A265;
  assign \new_[58564]_  = ~A299 & ~A298;
  assign \new_[58565]_  = \new_[58564]_  & \new_[58561]_ ;
  assign \new_[58566]_  = \new_[58565]_  & \new_[58558]_ ;
  assign \new_[58570]_  = A167 & ~A169;
  assign \new_[58571]_  = A170 & \new_[58570]_ ;
  assign \new_[58575]_  = ~A202 & ~A200;
  assign \new_[58576]_  = ~A166 & \new_[58575]_ ;
  assign \new_[58577]_  = \new_[58576]_  & \new_[58571]_ ;
  assign \new_[58581]_  = ~A233 & A232;
  assign \new_[58582]_  = ~A203 & \new_[58581]_ ;
  assign \new_[58585]_  = A235 & A234;
  assign \new_[58588]_  = A299 & ~A298;
  assign \new_[58589]_  = \new_[58588]_  & \new_[58585]_ ;
  assign \new_[58590]_  = \new_[58589]_  & \new_[58582]_ ;
  assign \new_[58594]_  = A167 & ~A169;
  assign \new_[58595]_  = A170 & \new_[58594]_ ;
  assign \new_[58599]_  = ~A202 & ~A200;
  assign \new_[58600]_  = ~A166 & \new_[58599]_ ;
  assign \new_[58601]_  = \new_[58600]_  & \new_[58595]_ ;
  assign \new_[58605]_  = ~A233 & A232;
  assign \new_[58606]_  = ~A203 & \new_[58605]_ ;
  assign \new_[58609]_  = A235 & A234;
  assign \new_[58612]_  = A266 & ~A265;
  assign \new_[58613]_  = \new_[58612]_  & \new_[58609]_ ;
  assign \new_[58614]_  = \new_[58613]_  & \new_[58606]_ ;
  assign \new_[58618]_  = A167 & ~A169;
  assign \new_[58619]_  = A170 & \new_[58618]_ ;
  assign \new_[58623]_  = ~A202 & ~A200;
  assign \new_[58624]_  = ~A166 & \new_[58623]_ ;
  assign \new_[58625]_  = \new_[58624]_  & \new_[58619]_ ;
  assign \new_[58629]_  = ~A233 & A232;
  assign \new_[58630]_  = ~A203 & \new_[58629]_ ;
  assign \new_[58633]_  = A236 & A234;
  assign \new_[58636]_  = A299 & ~A298;
  assign \new_[58637]_  = \new_[58636]_  & \new_[58633]_ ;
  assign \new_[58638]_  = \new_[58637]_  & \new_[58630]_ ;
  assign \new_[58642]_  = A167 & ~A169;
  assign \new_[58643]_  = A170 & \new_[58642]_ ;
  assign \new_[58647]_  = ~A202 & ~A200;
  assign \new_[58648]_  = ~A166 & \new_[58647]_ ;
  assign \new_[58649]_  = \new_[58648]_  & \new_[58643]_ ;
  assign \new_[58653]_  = ~A233 & A232;
  assign \new_[58654]_  = ~A203 & \new_[58653]_ ;
  assign \new_[58657]_  = A236 & A234;
  assign \new_[58660]_  = A266 & ~A265;
  assign \new_[58661]_  = \new_[58660]_  & \new_[58657]_ ;
  assign \new_[58662]_  = \new_[58661]_  & \new_[58654]_ ;
  assign \new_[58666]_  = A167 & ~A169;
  assign \new_[58667]_  = A170 & \new_[58666]_ ;
  assign \new_[58671]_  = ~A202 & ~A200;
  assign \new_[58672]_  = ~A166 & \new_[58671]_ ;
  assign \new_[58673]_  = \new_[58672]_  & \new_[58667]_ ;
  assign \new_[58677]_  = ~A233 & ~A232;
  assign \new_[58678]_  = ~A203 & \new_[58677]_ ;
  assign \new_[58681]_  = A266 & A265;
  assign \new_[58684]_  = ~A300 & A298;
  assign \new_[58685]_  = \new_[58684]_  & \new_[58681]_ ;
  assign \new_[58686]_  = \new_[58685]_  & \new_[58678]_ ;
  assign \new_[58690]_  = A167 & ~A169;
  assign \new_[58691]_  = A170 & \new_[58690]_ ;
  assign \new_[58695]_  = ~A202 & ~A200;
  assign \new_[58696]_  = ~A166 & \new_[58695]_ ;
  assign \new_[58697]_  = \new_[58696]_  & \new_[58691]_ ;
  assign \new_[58701]_  = ~A233 & ~A232;
  assign \new_[58702]_  = ~A203 & \new_[58701]_ ;
  assign \new_[58705]_  = A266 & A265;
  assign \new_[58708]_  = A299 & A298;
  assign \new_[58709]_  = \new_[58708]_  & \new_[58705]_ ;
  assign \new_[58710]_  = \new_[58709]_  & \new_[58702]_ ;
  assign \new_[58714]_  = A167 & ~A169;
  assign \new_[58715]_  = A170 & \new_[58714]_ ;
  assign \new_[58719]_  = ~A202 & ~A200;
  assign \new_[58720]_  = ~A166 & \new_[58719]_ ;
  assign \new_[58721]_  = \new_[58720]_  & \new_[58715]_ ;
  assign \new_[58725]_  = ~A233 & ~A232;
  assign \new_[58726]_  = ~A203 & \new_[58725]_ ;
  assign \new_[58729]_  = A266 & A265;
  assign \new_[58732]_  = ~A299 & ~A298;
  assign \new_[58733]_  = \new_[58732]_  & \new_[58729]_ ;
  assign \new_[58734]_  = \new_[58733]_  & \new_[58726]_ ;
  assign \new_[58738]_  = A167 & ~A169;
  assign \new_[58739]_  = A170 & \new_[58738]_ ;
  assign \new_[58743]_  = ~A202 & ~A200;
  assign \new_[58744]_  = ~A166 & \new_[58743]_ ;
  assign \new_[58745]_  = \new_[58744]_  & \new_[58739]_ ;
  assign \new_[58749]_  = ~A233 & ~A232;
  assign \new_[58750]_  = ~A203 & \new_[58749]_ ;
  assign \new_[58753]_  = ~A267 & ~A266;
  assign \new_[58756]_  = ~A300 & A298;
  assign \new_[58757]_  = \new_[58756]_  & \new_[58753]_ ;
  assign \new_[58758]_  = \new_[58757]_  & \new_[58750]_ ;
  assign \new_[58762]_  = A167 & ~A169;
  assign \new_[58763]_  = A170 & \new_[58762]_ ;
  assign \new_[58767]_  = ~A202 & ~A200;
  assign \new_[58768]_  = ~A166 & \new_[58767]_ ;
  assign \new_[58769]_  = \new_[58768]_  & \new_[58763]_ ;
  assign \new_[58773]_  = ~A233 & ~A232;
  assign \new_[58774]_  = ~A203 & \new_[58773]_ ;
  assign \new_[58777]_  = ~A267 & ~A266;
  assign \new_[58780]_  = A299 & A298;
  assign \new_[58781]_  = \new_[58780]_  & \new_[58777]_ ;
  assign \new_[58782]_  = \new_[58781]_  & \new_[58774]_ ;
  assign \new_[58786]_  = A167 & ~A169;
  assign \new_[58787]_  = A170 & \new_[58786]_ ;
  assign \new_[58791]_  = ~A202 & ~A200;
  assign \new_[58792]_  = ~A166 & \new_[58791]_ ;
  assign \new_[58793]_  = \new_[58792]_  & \new_[58787]_ ;
  assign \new_[58797]_  = ~A233 & ~A232;
  assign \new_[58798]_  = ~A203 & \new_[58797]_ ;
  assign \new_[58801]_  = ~A267 & ~A266;
  assign \new_[58804]_  = ~A299 & ~A298;
  assign \new_[58805]_  = \new_[58804]_  & \new_[58801]_ ;
  assign \new_[58806]_  = \new_[58805]_  & \new_[58798]_ ;
  assign \new_[58810]_  = A167 & ~A169;
  assign \new_[58811]_  = A170 & \new_[58810]_ ;
  assign \new_[58815]_  = ~A202 & ~A200;
  assign \new_[58816]_  = ~A166 & \new_[58815]_ ;
  assign \new_[58817]_  = \new_[58816]_  & \new_[58811]_ ;
  assign \new_[58821]_  = ~A233 & ~A232;
  assign \new_[58822]_  = ~A203 & \new_[58821]_ ;
  assign \new_[58825]_  = ~A266 & ~A265;
  assign \new_[58828]_  = ~A300 & A298;
  assign \new_[58829]_  = \new_[58828]_  & \new_[58825]_ ;
  assign \new_[58830]_  = \new_[58829]_  & \new_[58822]_ ;
  assign \new_[58834]_  = A167 & ~A169;
  assign \new_[58835]_  = A170 & \new_[58834]_ ;
  assign \new_[58839]_  = ~A202 & ~A200;
  assign \new_[58840]_  = ~A166 & \new_[58839]_ ;
  assign \new_[58841]_  = \new_[58840]_  & \new_[58835]_ ;
  assign \new_[58845]_  = ~A233 & ~A232;
  assign \new_[58846]_  = ~A203 & \new_[58845]_ ;
  assign \new_[58849]_  = ~A266 & ~A265;
  assign \new_[58852]_  = A299 & A298;
  assign \new_[58853]_  = \new_[58852]_  & \new_[58849]_ ;
  assign \new_[58854]_  = \new_[58853]_  & \new_[58846]_ ;
  assign \new_[58858]_  = A167 & ~A169;
  assign \new_[58859]_  = A170 & \new_[58858]_ ;
  assign \new_[58863]_  = ~A202 & ~A200;
  assign \new_[58864]_  = ~A166 & \new_[58863]_ ;
  assign \new_[58865]_  = \new_[58864]_  & \new_[58859]_ ;
  assign \new_[58869]_  = ~A233 & ~A232;
  assign \new_[58870]_  = ~A203 & \new_[58869]_ ;
  assign \new_[58873]_  = ~A266 & ~A265;
  assign \new_[58876]_  = ~A299 & ~A298;
  assign \new_[58877]_  = \new_[58876]_  & \new_[58873]_ ;
  assign \new_[58878]_  = \new_[58877]_  & \new_[58870]_ ;
  assign \new_[58882]_  = A167 & ~A169;
  assign \new_[58883]_  = A170 & \new_[58882]_ ;
  assign \new_[58887]_  = ~A201 & ~A200;
  assign \new_[58888]_  = ~A166 & \new_[58887]_ ;
  assign \new_[58889]_  = \new_[58888]_  & \new_[58883]_ ;
  assign \new_[58893]_  = A265 & A233;
  assign \new_[58894]_  = A232 & \new_[58893]_ ;
  assign \new_[58897]_  = ~A269 & ~A268;
  assign \new_[58900]_  = ~A300 & ~A299;
  assign \new_[58901]_  = \new_[58900]_  & \new_[58897]_ ;
  assign \new_[58902]_  = \new_[58901]_  & \new_[58894]_ ;
  assign \new_[58906]_  = A167 & ~A169;
  assign \new_[58907]_  = A170 & \new_[58906]_ ;
  assign \new_[58911]_  = ~A201 & ~A200;
  assign \new_[58912]_  = ~A166 & \new_[58911]_ ;
  assign \new_[58913]_  = \new_[58912]_  & \new_[58907]_ ;
  assign \new_[58917]_  = A265 & A233;
  assign \new_[58918]_  = A232 & \new_[58917]_ ;
  assign \new_[58921]_  = ~A269 & ~A268;
  assign \new_[58924]_  = A299 & A298;
  assign \new_[58925]_  = \new_[58924]_  & \new_[58921]_ ;
  assign \new_[58926]_  = \new_[58925]_  & \new_[58918]_ ;
  assign \new_[58930]_  = A167 & ~A169;
  assign \new_[58931]_  = A170 & \new_[58930]_ ;
  assign \new_[58935]_  = ~A201 & ~A200;
  assign \new_[58936]_  = ~A166 & \new_[58935]_ ;
  assign \new_[58937]_  = \new_[58936]_  & \new_[58931]_ ;
  assign \new_[58941]_  = A265 & A233;
  assign \new_[58942]_  = A232 & \new_[58941]_ ;
  assign \new_[58945]_  = ~A269 & ~A268;
  assign \new_[58948]_  = ~A299 & ~A298;
  assign \new_[58949]_  = \new_[58948]_  & \new_[58945]_ ;
  assign \new_[58950]_  = \new_[58949]_  & \new_[58942]_ ;
  assign \new_[58954]_  = A167 & ~A169;
  assign \new_[58955]_  = A170 & \new_[58954]_ ;
  assign \new_[58959]_  = ~A201 & ~A200;
  assign \new_[58960]_  = ~A166 & \new_[58959]_ ;
  assign \new_[58961]_  = \new_[58960]_  & \new_[58955]_ ;
  assign \new_[58965]_  = A265 & A233;
  assign \new_[58966]_  = A232 & \new_[58965]_ ;
  assign \new_[58969]_  = ~A299 & ~A267;
  assign \new_[58972]_  = ~A302 & ~A301;
  assign \new_[58973]_  = \new_[58972]_  & \new_[58969]_ ;
  assign \new_[58974]_  = \new_[58973]_  & \new_[58966]_ ;
  assign \new_[58978]_  = A167 & ~A169;
  assign \new_[58979]_  = A170 & \new_[58978]_ ;
  assign \new_[58983]_  = ~A201 & ~A200;
  assign \new_[58984]_  = ~A166 & \new_[58983]_ ;
  assign \new_[58985]_  = \new_[58984]_  & \new_[58979]_ ;
  assign \new_[58989]_  = A265 & A233;
  assign \new_[58990]_  = A232 & \new_[58989]_ ;
  assign \new_[58993]_  = ~A299 & A266;
  assign \new_[58996]_  = ~A302 & ~A301;
  assign \new_[58997]_  = \new_[58996]_  & \new_[58993]_ ;
  assign \new_[58998]_  = \new_[58997]_  & \new_[58990]_ ;
  assign \new_[59002]_  = A167 & ~A169;
  assign \new_[59003]_  = A170 & \new_[59002]_ ;
  assign \new_[59007]_  = ~A201 & ~A200;
  assign \new_[59008]_  = ~A166 & \new_[59007]_ ;
  assign \new_[59009]_  = \new_[59008]_  & \new_[59003]_ ;
  assign \new_[59013]_  = ~A265 & A233;
  assign \new_[59014]_  = A232 & \new_[59013]_ ;
  assign \new_[59017]_  = ~A299 & ~A266;
  assign \new_[59020]_  = ~A302 & ~A301;
  assign \new_[59021]_  = \new_[59020]_  & \new_[59017]_ ;
  assign \new_[59022]_  = \new_[59021]_  & \new_[59014]_ ;
  assign \new_[59026]_  = A167 & ~A169;
  assign \new_[59027]_  = A170 & \new_[59026]_ ;
  assign \new_[59031]_  = ~A201 & ~A200;
  assign \new_[59032]_  = ~A166 & \new_[59031]_ ;
  assign \new_[59033]_  = \new_[59032]_  & \new_[59027]_ ;
  assign \new_[59037]_  = ~A236 & ~A235;
  assign \new_[59038]_  = ~A233 & \new_[59037]_ ;
  assign \new_[59041]_  = A266 & A265;
  assign \new_[59044]_  = ~A300 & A298;
  assign \new_[59045]_  = \new_[59044]_  & \new_[59041]_ ;
  assign \new_[59046]_  = \new_[59045]_  & \new_[59038]_ ;
  assign \new_[59050]_  = A167 & ~A169;
  assign \new_[59051]_  = A170 & \new_[59050]_ ;
  assign \new_[59055]_  = ~A201 & ~A200;
  assign \new_[59056]_  = ~A166 & \new_[59055]_ ;
  assign \new_[59057]_  = \new_[59056]_  & \new_[59051]_ ;
  assign \new_[59061]_  = ~A236 & ~A235;
  assign \new_[59062]_  = ~A233 & \new_[59061]_ ;
  assign \new_[59065]_  = A266 & A265;
  assign \new_[59068]_  = A299 & A298;
  assign \new_[59069]_  = \new_[59068]_  & \new_[59065]_ ;
  assign \new_[59070]_  = \new_[59069]_  & \new_[59062]_ ;
  assign \new_[59074]_  = A167 & ~A169;
  assign \new_[59075]_  = A170 & \new_[59074]_ ;
  assign \new_[59079]_  = ~A201 & ~A200;
  assign \new_[59080]_  = ~A166 & \new_[59079]_ ;
  assign \new_[59081]_  = \new_[59080]_  & \new_[59075]_ ;
  assign \new_[59085]_  = ~A236 & ~A235;
  assign \new_[59086]_  = ~A233 & \new_[59085]_ ;
  assign \new_[59089]_  = A266 & A265;
  assign \new_[59092]_  = ~A299 & ~A298;
  assign \new_[59093]_  = \new_[59092]_  & \new_[59089]_ ;
  assign \new_[59094]_  = \new_[59093]_  & \new_[59086]_ ;
  assign \new_[59098]_  = A167 & ~A169;
  assign \new_[59099]_  = A170 & \new_[59098]_ ;
  assign \new_[59103]_  = ~A201 & ~A200;
  assign \new_[59104]_  = ~A166 & \new_[59103]_ ;
  assign \new_[59105]_  = \new_[59104]_  & \new_[59099]_ ;
  assign \new_[59109]_  = ~A236 & ~A235;
  assign \new_[59110]_  = ~A233 & \new_[59109]_ ;
  assign \new_[59113]_  = ~A267 & ~A266;
  assign \new_[59116]_  = ~A300 & A298;
  assign \new_[59117]_  = \new_[59116]_  & \new_[59113]_ ;
  assign \new_[59118]_  = \new_[59117]_  & \new_[59110]_ ;
  assign \new_[59122]_  = A167 & ~A169;
  assign \new_[59123]_  = A170 & \new_[59122]_ ;
  assign \new_[59127]_  = ~A201 & ~A200;
  assign \new_[59128]_  = ~A166 & \new_[59127]_ ;
  assign \new_[59129]_  = \new_[59128]_  & \new_[59123]_ ;
  assign \new_[59133]_  = ~A236 & ~A235;
  assign \new_[59134]_  = ~A233 & \new_[59133]_ ;
  assign \new_[59137]_  = ~A267 & ~A266;
  assign \new_[59140]_  = A299 & A298;
  assign \new_[59141]_  = \new_[59140]_  & \new_[59137]_ ;
  assign \new_[59142]_  = \new_[59141]_  & \new_[59134]_ ;
  assign \new_[59146]_  = A167 & ~A169;
  assign \new_[59147]_  = A170 & \new_[59146]_ ;
  assign \new_[59151]_  = ~A201 & ~A200;
  assign \new_[59152]_  = ~A166 & \new_[59151]_ ;
  assign \new_[59153]_  = \new_[59152]_  & \new_[59147]_ ;
  assign \new_[59157]_  = ~A236 & ~A235;
  assign \new_[59158]_  = ~A233 & \new_[59157]_ ;
  assign \new_[59161]_  = ~A267 & ~A266;
  assign \new_[59164]_  = ~A299 & ~A298;
  assign \new_[59165]_  = \new_[59164]_  & \new_[59161]_ ;
  assign \new_[59166]_  = \new_[59165]_  & \new_[59158]_ ;
  assign \new_[59170]_  = A167 & ~A169;
  assign \new_[59171]_  = A170 & \new_[59170]_ ;
  assign \new_[59175]_  = ~A201 & ~A200;
  assign \new_[59176]_  = ~A166 & \new_[59175]_ ;
  assign \new_[59177]_  = \new_[59176]_  & \new_[59171]_ ;
  assign \new_[59181]_  = ~A236 & ~A235;
  assign \new_[59182]_  = ~A233 & \new_[59181]_ ;
  assign \new_[59185]_  = ~A266 & ~A265;
  assign \new_[59188]_  = ~A300 & A298;
  assign \new_[59189]_  = \new_[59188]_  & \new_[59185]_ ;
  assign \new_[59190]_  = \new_[59189]_  & \new_[59182]_ ;
  assign \new_[59194]_  = A167 & ~A169;
  assign \new_[59195]_  = A170 & \new_[59194]_ ;
  assign \new_[59199]_  = ~A201 & ~A200;
  assign \new_[59200]_  = ~A166 & \new_[59199]_ ;
  assign \new_[59201]_  = \new_[59200]_  & \new_[59195]_ ;
  assign \new_[59205]_  = ~A236 & ~A235;
  assign \new_[59206]_  = ~A233 & \new_[59205]_ ;
  assign \new_[59209]_  = ~A266 & ~A265;
  assign \new_[59212]_  = A299 & A298;
  assign \new_[59213]_  = \new_[59212]_  & \new_[59209]_ ;
  assign \new_[59214]_  = \new_[59213]_  & \new_[59206]_ ;
  assign \new_[59218]_  = A167 & ~A169;
  assign \new_[59219]_  = A170 & \new_[59218]_ ;
  assign \new_[59223]_  = ~A201 & ~A200;
  assign \new_[59224]_  = ~A166 & \new_[59223]_ ;
  assign \new_[59225]_  = \new_[59224]_  & \new_[59219]_ ;
  assign \new_[59229]_  = ~A236 & ~A235;
  assign \new_[59230]_  = ~A233 & \new_[59229]_ ;
  assign \new_[59233]_  = ~A266 & ~A265;
  assign \new_[59236]_  = ~A299 & ~A298;
  assign \new_[59237]_  = \new_[59236]_  & \new_[59233]_ ;
  assign \new_[59238]_  = \new_[59237]_  & \new_[59230]_ ;
  assign \new_[59242]_  = A167 & ~A169;
  assign \new_[59243]_  = A170 & \new_[59242]_ ;
  assign \new_[59247]_  = ~A201 & ~A200;
  assign \new_[59248]_  = ~A166 & \new_[59247]_ ;
  assign \new_[59249]_  = \new_[59248]_  & \new_[59243]_ ;
  assign \new_[59253]_  = A265 & ~A234;
  assign \new_[59254]_  = ~A233 & \new_[59253]_ ;
  assign \new_[59257]_  = A298 & A266;
  assign \new_[59260]_  = ~A302 & ~A301;
  assign \new_[59261]_  = \new_[59260]_  & \new_[59257]_ ;
  assign \new_[59262]_  = \new_[59261]_  & \new_[59254]_ ;
  assign \new_[59266]_  = A167 & ~A169;
  assign \new_[59267]_  = A170 & \new_[59266]_ ;
  assign \new_[59271]_  = ~A201 & ~A200;
  assign \new_[59272]_  = ~A166 & \new_[59271]_ ;
  assign \new_[59273]_  = \new_[59272]_  & \new_[59267]_ ;
  assign \new_[59277]_  = ~A266 & ~A234;
  assign \new_[59278]_  = ~A233 & \new_[59277]_ ;
  assign \new_[59281]_  = ~A269 & ~A268;
  assign \new_[59284]_  = ~A300 & A298;
  assign \new_[59285]_  = \new_[59284]_  & \new_[59281]_ ;
  assign \new_[59286]_  = \new_[59285]_  & \new_[59278]_ ;
  assign \new_[59290]_  = A167 & ~A169;
  assign \new_[59291]_  = A170 & \new_[59290]_ ;
  assign \new_[59295]_  = ~A201 & ~A200;
  assign \new_[59296]_  = ~A166 & \new_[59295]_ ;
  assign \new_[59297]_  = \new_[59296]_  & \new_[59291]_ ;
  assign \new_[59301]_  = ~A266 & ~A234;
  assign \new_[59302]_  = ~A233 & \new_[59301]_ ;
  assign \new_[59305]_  = ~A269 & ~A268;
  assign \new_[59308]_  = A299 & A298;
  assign \new_[59309]_  = \new_[59308]_  & \new_[59305]_ ;
  assign \new_[59310]_  = \new_[59309]_  & \new_[59302]_ ;
  assign \new_[59314]_  = A167 & ~A169;
  assign \new_[59315]_  = A170 & \new_[59314]_ ;
  assign \new_[59319]_  = ~A201 & ~A200;
  assign \new_[59320]_  = ~A166 & \new_[59319]_ ;
  assign \new_[59321]_  = \new_[59320]_  & \new_[59315]_ ;
  assign \new_[59325]_  = ~A266 & ~A234;
  assign \new_[59326]_  = ~A233 & \new_[59325]_ ;
  assign \new_[59329]_  = ~A269 & ~A268;
  assign \new_[59332]_  = ~A299 & ~A298;
  assign \new_[59333]_  = \new_[59332]_  & \new_[59329]_ ;
  assign \new_[59334]_  = \new_[59333]_  & \new_[59326]_ ;
  assign \new_[59338]_  = A167 & ~A169;
  assign \new_[59339]_  = A170 & \new_[59338]_ ;
  assign \new_[59343]_  = ~A201 & ~A200;
  assign \new_[59344]_  = ~A166 & \new_[59343]_ ;
  assign \new_[59345]_  = \new_[59344]_  & \new_[59339]_ ;
  assign \new_[59349]_  = ~A266 & ~A234;
  assign \new_[59350]_  = ~A233 & \new_[59349]_ ;
  assign \new_[59353]_  = A298 & ~A267;
  assign \new_[59356]_  = ~A302 & ~A301;
  assign \new_[59357]_  = \new_[59356]_  & \new_[59353]_ ;
  assign \new_[59358]_  = \new_[59357]_  & \new_[59350]_ ;
  assign \new_[59362]_  = A167 & ~A169;
  assign \new_[59363]_  = A170 & \new_[59362]_ ;
  assign \new_[59367]_  = ~A201 & ~A200;
  assign \new_[59368]_  = ~A166 & \new_[59367]_ ;
  assign \new_[59369]_  = \new_[59368]_  & \new_[59363]_ ;
  assign \new_[59373]_  = ~A265 & ~A234;
  assign \new_[59374]_  = ~A233 & \new_[59373]_ ;
  assign \new_[59377]_  = A298 & ~A266;
  assign \new_[59380]_  = ~A302 & ~A301;
  assign \new_[59381]_  = \new_[59380]_  & \new_[59377]_ ;
  assign \new_[59382]_  = \new_[59381]_  & \new_[59374]_ ;
  assign \new_[59386]_  = A167 & ~A169;
  assign \new_[59387]_  = A170 & \new_[59386]_ ;
  assign \new_[59391]_  = ~A201 & ~A200;
  assign \new_[59392]_  = ~A166 & \new_[59391]_ ;
  assign \new_[59393]_  = \new_[59392]_  & \new_[59387]_ ;
  assign \new_[59397]_  = A265 & ~A233;
  assign \new_[59398]_  = ~A232 & \new_[59397]_ ;
  assign \new_[59401]_  = A298 & A266;
  assign \new_[59404]_  = ~A302 & ~A301;
  assign \new_[59405]_  = \new_[59404]_  & \new_[59401]_ ;
  assign \new_[59406]_  = \new_[59405]_  & \new_[59398]_ ;
  assign \new_[59410]_  = A167 & ~A169;
  assign \new_[59411]_  = A170 & \new_[59410]_ ;
  assign \new_[59415]_  = ~A201 & ~A200;
  assign \new_[59416]_  = ~A166 & \new_[59415]_ ;
  assign \new_[59417]_  = \new_[59416]_  & \new_[59411]_ ;
  assign \new_[59421]_  = ~A266 & ~A233;
  assign \new_[59422]_  = ~A232 & \new_[59421]_ ;
  assign \new_[59425]_  = ~A269 & ~A268;
  assign \new_[59428]_  = ~A300 & A298;
  assign \new_[59429]_  = \new_[59428]_  & \new_[59425]_ ;
  assign \new_[59430]_  = \new_[59429]_  & \new_[59422]_ ;
  assign \new_[59434]_  = A167 & ~A169;
  assign \new_[59435]_  = A170 & \new_[59434]_ ;
  assign \new_[59439]_  = ~A201 & ~A200;
  assign \new_[59440]_  = ~A166 & \new_[59439]_ ;
  assign \new_[59441]_  = \new_[59440]_  & \new_[59435]_ ;
  assign \new_[59445]_  = ~A266 & ~A233;
  assign \new_[59446]_  = ~A232 & \new_[59445]_ ;
  assign \new_[59449]_  = ~A269 & ~A268;
  assign \new_[59452]_  = A299 & A298;
  assign \new_[59453]_  = \new_[59452]_  & \new_[59449]_ ;
  assign \new_[59454]_  = \new_[59453]_  & \new_[59446]_ ;
  assign \new_[59458]_  = A167 & ~A169;
  assign \new_[59459]_  = A170 & \new_[59458]_ ;
  assign \new_[59463]_  = ~A201 & ~A200;
  assign \new_[59464]_  = ~A166 & \new_[59463]_ ;
  assign \new_[59465]_  = \new_[59464]_  & \new_[59459]_ ;
  assign \new_[59469]_  = ~A266 & ~A233;
  assign \new_[59470]_  = ~A232 & \new_[59469]_ ;
  assign \new_[59473]_  = ~A269 & ~A268;
  assign \new_[59476]_  = ~A299 & ~A298;
  assign \new_[59477]_  = \new_[59476]_  & \new_[59473]_ ;
  assign \new_[59478]_  = \new_[59477]_  & \new_[59470]_ ;
  assign \new_[59482]_  = A167 & ~A169;
  assign \new_[59483]_  = A170 & \new_[59482]_ ;
  assign \new_[59487]_  = ~A201 & ~A200;
  assign \new_[59488]_  = ~A166 & \new_[59487]_ ;
  assign \new_[59489]_  = \new_[59488]_  & \new_[59483]_ ;
  assign \new_[59493]_  = ~A266 & ~A233;
  assign \new_[59494]_  = ~A232 & \new_[59493]_ ;
  assign \new_[59497]_  = A298 & ~A267;
  assign \new_[59500]_  = ~A302 & ~A301;
  assign \new_[59501]_  = \new_[59500]_  & \new_[59497]_ ;
  assign \new_[59502]_  = \new_[59501]_  & \new_[59494]_ ;
  assign \new_[59506]_  = A167 & ~A169;
  assign \new_[59507]_  = A170 & \new_[59506]_ ;
  assign \new_[59511]_  = ~A201 & ~A200;
  assign \new_[59512]_  = ~A166 & \new_[59511]_ ;
  assign \new_[59513]_  = \new_[59512]_  & \new_[59507]_ ;
  assign \new_[59517]_  = ~A265 & ~A233;
  assign \new_[59518]_  = ~A232 & \new_[59517]_ ;
  assign \new_[59521]_  = A298 & ~A266;
  assign \new_[59524]_  = ~A302 & ~A301;
  assign \new_[59525]_  = \new_[59524]_  & \new_[59521]_ ;
  assign \new_[59526]_  = \new_[59525]_  & \new_[59518]_ ;
  assign \new_[59530]_  = A167 & ~A169;
  assign \new_[59531]_  = A170 & \new_[59530]_ ;
  assign \new_[59535]_  = ~A200 & ~A199;
  assign \new_[59536]_  = ~A166 & \new_[59535]_ ;
  assign \new_[59537]_  = \new_[59536]_  & \new_[59531]_ ;
  assign \new_[59541]_  = A265 & A233;
  assign \new_[59542]_  = A232 & \new_[59541]_ ;
  assign \new_[59545]_  = ~A269 & ~A268;
  assign \new_[59548]_  = ~A300 & ~A299;
  assign \new_[59549]_  = \new_[59548]_  & \new_[59545]_ ;
  assign \new_[59550]_  = \new_[59549]_  & \new_[59542]_ ;
  assign \new_[59554]_  = A167 & ~A169;
  assign \new_[59555]_  = A170 & \new_[59554]_ ;
  assign \new_[59559]_  = ~A200 & ~A199;
  assign \new_[59560]_  = ~A166 & \new_[59559]_ ;
  assign \new_[59561]_  = \new_[59560]_  & \new_[59555]_ ;
  assign \new_[59565]_  = A265 & A233;
  assign \new_[59566]_  = A232 & \new_[59565]_ ;
  assign \new_[59569]_  = ~A269 & ~A268;
  assign \new_[59572]_  = A299 & A298;
  assign \new_[59573]_  = \new_[59572]_  & \new_[59569]_ ;
  assign \new_[59574]_  = \new_[59573]_  & \new_[59566]_ ;
  assign \new_[59578]_  = A167 & ~A169;
  assign \new_[59579]_  = A170 & \new_[59578]_ ;
  assign \new_[59583]_  = ~A200 & ~A199;
  assign \new_[59584]_  = ~A166 & \new_[59583]_ ;
  assign \new_[59585]_  = \new_[59584]_  & \new_[59579]_ ;
  assign \new_[59589]_  = A265 & A233;
  assign \new_[59590]_  = A232 & \new_[59589]_ ;
  assign \new_[59593]_  = ~A269 & ~A268;
  assign \new_[59596]_  = ~A299 & ~A298;
  assign \new_[59597]_  = \new_[59596]_  & \new_[59593]_ ;
  assign \new_[59598]_  = \new_[59597]_  & \new_[59590]_ ;
  assign \new_[59602]_  = A167 & ~A169;
  assign \new_[59603]_  = A170 & \new_[59602]_ ;
  assign \new_[59607]_  = ~A200 & ~A199;
  assign \new_[59608]_  = ~A166 & \new_[59607]_ ;
  assign \new_[59609]_  = \new_[59608]_  & \new_[59603]_ ;
  assign \new_[59613]_  = A265 & A233;
  assign \new_[59614]_  = A232 & \new_[59613]_ ;
  assign \new_[59617]_  = ~A299 & ~A267;
  assign \new_[59620]_  = ~A302 & ~A301;
  assign \new_[59621]_  = \new_[59620]_  & \new_[59617]_ ;
  assign \new_[59622]_  = \new_[59621]_  & \new_[59614]_ ;
  assign \new_[59626]_  = A167 & ~A169;
  assign \new_[59627]_  = A170 & \new_[59626]_ ;
  assign \new_[59631]_  = ~A200 & ~A199;
  assign \new_[59632]_  = ~A166 & \new_[59631]_ ;
  assign \new_[59633]_  = \new_[59632]_  & \new_[59627]_ ;
  assign \new_[59637]_  = A265 & A233;
  assign \new_[59638]_  = A232 & \new_[59637]_ ;
  assign \new_[59641]_  = ~A299 & A266;
  assign \new_[59644]_  = ~A302 & ~A301;
  assign \new_[59645]_  = \new_[59644]_  & \new_[59641]_ ;
  assign \new_[59646]_  = \new_[59645]_  & \new_[59638]_ ;
  assign \new_[59650]_  = A167 & ~A169;
  assign \new_[59651]_  = A170 & \new_[59650]_ ;
  assign \new_[59655]_  = ~A200 & ~A199;
  assign \new_[59656]_  = ~A166 & \new_[59655]_ ;
  assign \new_[59657]_  = \new_[59656]_  & \new_[59651]_ ;
  assign \new_[59661]_  = ~A265 & A233;
  assign \new_[59662]_  = A232 & \new_[59661]_ ;
  assign \new_[59665]_  = ~A299 & ~A266;
  assign \new_[59668]_  = ~A302 & ~A301;
  assign \new_[59669]_  = \new_[59668]_  & \new_[59665]_ ;
  assign \new_[59670]_  = \new_[59669]_  & \new_[59662]_ ;
  assign \new_[59674]_  = A167 & ~A169;
  assign \new_[59675]_  = A170 & \new_[59674]_ ;
  assign \new_[59679]_  = ~A200 & ~A199;
  assign \new_[59680]_  = ~A166 & \new_[59679]_ ;
  assign \new_[59681]_  = \new_[59680]_  & \new_[59675]_ ;
  assign \new_[59685]_  = ~A236 & ~A235;
  assign \new_[59686]_  = ~A233 & \new_[59685]_ ;
  assign \new_[59689]_  = A266 & A265;
  assign \new_[59692]_  = ~A300 & A298;
  assign \new_[59693]_  = \new_[59692]_  & \new_[59689]_ ;
  assign \new_[59694]_  = \new_[59693]_  & \new_[59686]_ ;
  assign \new_[59698]_  = A167 & ~A169;
  assign \new_[59699]_  = A170 & \new_[59698]_ ;
  assign \new_[59703]_  = ~A200 & ~A199;
  assign \new_[59704]_  = ~A166 & \new_[59703]_ ;
  assign \new_[59705]_  = \new_[59704]_  & \new_[59699]_ ;
  assign \new_[59709]_  = ~A236 & ~A235;
  assign \new_[59710]_  = ~A233 & \new_[59709]_ ;
  assign \new_[59713]_  = A266 & A265;
  assign \new_[59716]_  = A299 & A298;
  assign \new_[59717]_  = \new_[59716]_  & \new_[59713]_ ;
  assign \new_[59718]_  = \new_[59717]_  & \new_[59710]_ ;
  assign \new_[59722]_  = A167 & ~A169;
  assign \new_[59723]_  = A170 & \new_[59722]_ ;
  assign \new_[59727]_  = ~A200 & ~A199;
  assign \new_[59728]_  = ~A166 & \new_[59727]_ ;
  assign \new_[59729]_  = \new_[59728]_  & \new_[59723]_ ;
  assign \new_[59733]_  = ~A236 & ~A235;
  assign \new_[59734]_  = ~A233 & \new_[59733]_ ;
  assign \new_[59737]_  = A266 & A265;
  assign \new_[59740]_  = ~A299 & ~A298;
  assign \new_[59741]_  = \new_[59740]_  & \new_[59737]_ ;
  assign \new_[59742]_  = \new_[59741]_  & \new_[59734]_ ;
  assign \new_[59746]_  = A167 & ~A169;
  assign \new_[59747]_  = A170 & \new_[59746]_ ;
  assign \new_[59751]_  = ~A200 & ~A199;
  assign \new_[59752]_  = ~A166 & \new_[59751]_ ;
  assign \new_[59753]_  = \new_[59752]_  & \new_[59747]_ ;
  assign \new_[59757]_  = ~A236 & ~A235;
  assign \new_[59758]_  = ~A233 & \new_[59757]_ ;
  assign \new_[59761]_  = ~A267 & ~A266;
  assign \new_[59764]_  = ~A300 & A298;
  assign \new_[59765]_  = \new_[59764]_  & \new_[59761]_ ;
  assign \new_[59766]_  = \new_[59765]_  & \new_[59758]_ ;
  assign \new_[59770]_  = A167 & ~A169;
  assign \new_[59771]_  = A170 & \new_[59770]_ ;
  assign \new_[59775]_  = ~A200 & ~A199;
  assign \new_[59776]_  = ~A166 & \new_[59775]_ ;
  assign \new_[59777]_  = \new_[59776]_  & \new_[59771]_ ;
  assign \new_[59781]_  = ~A236 & ~A235;
  assign \new_[59782]_  = ~A233 & \new_[59781]_ ;
  assign \new_[59785]_  = ~A267 & ~A266;
  assign \new_[59788]_  = A299 & A298;
  assign \new_[59789]_  = \new_[59788]_  & \new_[59785]_ ;
  assign \new_[59790]_  = \new_[59789]_  & \new_[59782]_ ;
  assign \new_[59794]_  = A167 & ~A169;
  assign \new_[59795]_  = A170 & \new_[59794]_ ;
  assign \new_[59799]_  = ~A200 & ~A199;
  assign \new_[59800]_  = ~A166 & \new_[59799]_ ;
  assign \new_[59801]_  = \new_[59800]_  & \new_[59795]_ ;
  assign \new_[59805]_  = ~A236 & ~A235;
  assign \new_[59806]_  = ~A233 & \new_[59805]_ ;
  assign \new_[59809]_  = ~A267 & ~A266;
  assign \new_[59812]_  = ~A299 & ~A298;
  assign \new_[59813]_  = \new_[59812]_  & \new_[59809]_ ;
  assign \new_[59814]_  = \new_[59813]_  & \new_[59806]_ ;
  assign \new_[59818]_  = A167 & ~A169;
  assign \new_[59819]_  = A170 & \new_[59818]_ ;
  assign \new_[59823]_  = ~A200 & ~A199;
  assign \new_[59824]_  = ~A166 & \new_[59823]_ ;
  assign \new_[59825]_  = \new_[59824]_  & \new_[59819]_ ;
  assign \new_[59829]_  = ~A236 & ~A235;
  assign \new_[59830]_  = ~A233 & \new_[59829]_ ;
  assign \new_[59833]_  = ~A266 & ~A265;
  assign \new_[59836]_  = ~A300 & A298;
  assign \new_[59837]_  = \new_[59836]_  & \new_[59833]_ ;
  assign \new_[59838]_  = \new_[59837]_  & \new_[59830]_ ;
  assign \new_[59842]_  = A167 & ~A169;
  assign \new_[59843]_  = A170 & \new_[59842]_ ;
  assign \new_[59847]_  = ~A200 & ~A199;
  assign \new_[59848]_  = ~A166 & \new_[59847]_ ;
  assign \new_[59849]_  = \new_[59848]_  & \new_[59843]_ ;
  assign \new_[59853]_  = ~A236 & ~A235;
  assign \new_[59854]_  = ~A233 & \new_[59853]_ ;
  assign \new_[59857]_  = ~A266 & ~A265;
  assign \new_[59860]_  = A299 & A298;
  assign \new_[59861]_  = \new_[59860]_  & \new_[59857]_ ;
  assign \new_[59862]_  = \new_[59861]_  & \new_[59854]_ ;
  assign \new_[59866]_  = A167 & ~A169;
  assign \new_[59867]_  = A170 & \new_[59866]_ ;
  assign \new_[59871]_  = ~A200 & ~A199;
  assign \new_[59872]_  = ~A166 & \new_[59871]_ ;
  assign \new_[59873]_  = \new_[59872]_  & \new_[59867]_ ;
  assign \new_[59877]_  = ~A236 & ~A235;
  assign \new_[59878]_  = ~A233 & \new_[59877]_ ;
  assign \new_[59881]_  = ~A266 & ~A265;
  assign \new_[59884]_  = ~A299 & ~A298;
  assign \new_[59885]_  = \new_[59884]_  & \new_[59881]_ ;
  assign \new_[59886]_  = \new_[59885]_  & \new_[59878]_ ;
  assign \new_[59890]_  = A167 & ~A169;
  assign \new_[59891]_  = A170 & \new_[59890]_ ;
  assign \new_[59895]_  = ~A200 & ~A199;
  assign \new_[59896]_  = ~A166 & \new_[59895]_ ;
  assign \new_[59897]_  = \new_[59896]_  & \new_[59891]_ ;
  assign \new_[59901]_  = A265 & ~A234;
  assign \new_[59902]_  = ~A233 & \new_[59901]_ ;
  assign \new_[59905]_  = A298 & A266;
  assign \new_[59908]_  = ~A302 & ~A301;
  assign \new_[59909]_  = \new_[59908]_  & \new_[59905]_ ;
  assign \new_[59910]_  = \new_[59909]_  & \new_[59902]_ ;
  assign \new_[59914]_  = A167 & ~A169;
  assign \new_[59915]_  = A170 & \new_[59914]_ ;
  assign \new_[59919]_  = ~A200 & ~A199;
  assign \new_[59920]_  = ~A166 & \new_[59919]_ ;
  assign \new_[59921]_  = \new_[59920]_  & \new_[59915]_ ;
  assign \new_[59925]_  = ~A266 & ~A234;
  assign \new_[59926]_  = ~A233 & \new_[59925]_ ;
  assign \new_[59929]_  = ~A269 & ~A268;
  assign \new_[59932]_  = ~A300 & A298;
  assign \new_[59933]_  = \new_[59932]_  & \new_[59929]_ ;
  assign \new_[59934]_  = \new_[59933]_  & \new_[59926]_ ;
  assign \new_[59938]_  = A167 & ~A169;
  assign \new_[59939]_  = A170 & \new_[59938]_ ;
  assign \new_[59943]_  = ~A200 & ~A199;
  assign \new_[59944]_  = ~A166 & \new_[59943]_ ;
  assign \new_[59945]_  = \new_[59944]_  & \new_[59939]_ ;
  assign \new_[59949]_  = ~A266 & ~A234;
  assign \new_[59950]_  = ~A233 & \new_[59949]_ ;
  assign \new_[59953]_  = ~A269 & ~A268;
  assign \new_[59956]_  = A299 & A298;
  assign \new_[59957]_  = \new_[59956]_  & \new_[59953]_ ;
  assign \new_[59958]_  = \new_[59957]_  & \new_[59950]_ ;
  assign \new_[59962]_  = A167 & ~A169;
  assign \new_[59963]_  = A170 & \new_[59962]_ ;
  assign \new_[59967]_  = ~A200 & ~A199;
  assign \new_[59968]_  = ~A166 & \new_[59967]_ ;
  assign \new_[59969]_  = \new_[59968]_  & \new_[59963]_ ;
  assign \new_[59973]_  = ~A266 & ~A234;
  assign \new_[59974]_  = ~A233 & \new_[59973]_ ;
  assign \new_[59977]_  = ~A269 & ~A268;
  assign \new_[59980]_  = ~A299 & ~A298;
  assign \new_[59981]_  = \new_[59980]_  & \new_[59977]_ ;
  assign \new_[59982]_  = \new_[59981]_  & \new_[59974]_ ;
  assign \new_[59986]_  = A167 & ~A169;
  assign \new_[59987]_  = A170 & \new_[59986]_ ;
  assign \new_[59991]_  = ~A200 & ~A199;
  assign \new_[59992]_  = ~A166 & \new_[59991]_ ;
  assign \new_[59993]_  = \new_[59992]_  & \new_[59987]_ ;
  assign \new_[59997]_  = ~A266 & ~A234;
  assign \new_[59998]_  = ~A233 & \new_[59997]_ ;
  assign \new_[60001]_  = A298 & ~A267;
  assign \new_[60004]_  = ~A302 & ~A301;
  assign \new_[60005]_  = \new_[60004]_  & \new_[60001]_ ;
  assign \new_[60006]_  = \new_[60005]_  & \new_[59998]_ ;
  assign \new_[60010]_  = A167 & ~A169;
  assign \new_[60011]_  = A170 & \new_[60010]_ ;
  assign \new_[60015]_  = ~A200 & ~A199;
  assign \new_[60016]_  = ~A166 & \new_[60015]_ ;
  assign \new_[60017]_  = \new_[60016]_  & \new_[60011]_ ;
  assign \new_[60021]_  = ~A265 & ~A234;
  assign \new_[60022]_  = ~A233 & \new_[60021]_ ;
  assign \new_[60025]_  = A298 & ~A266;
  assign \new_[60028]_  = ~A302 & ~A301;
  assign \new_[60029]_  = \new_[60028]_  & \new_[60025]_ ;
  assign \new_[60030]_  = \new_[60029]_  & \new_[60022]_ ;
  assign \new_[60034]_  = A167 & ~A169;
  assign \new_[60035]_  = A170 & \new_[60034]_ ;
  assign \new_[60039]_  = ~A200 & ~A199;
  assign \new_[60040]_  = ~A166 & \new_[60039]_ ;
  assign \new_[60041]_  = \new_[60040]_  & \new_[60035]_ ;
  assign \new_[60045]_  = A265 & ~A233;
  assign \new_[60046]_  = ~A232 & \new_[60045]_ ;
  assign \new_[60049]_  = A298 & A266;
  assign \new_[60052]_  = ~A302 & ~A301;
  assign \new_[60053]_  = \new_[60052]_  & \new_[60049]_ ;
  assign \new_[60054]_  = \new_[60053]_  & \new_[60046]_ ;
  assign \new_[60058]_  = A167 & ~A169;
  assign \new_[60059]_  = A170 & \new_[60058]_ ;
  assign \new_[60063]_  = ~A200 & ~A199;
  assign \new_[60064]_  = ~A166 & \new_[60063]_ ;
  assign \new_[60065]_  = \new_[60064]_  & \new_[60059]_ ;
  assign \new_[60069]_  = ~A266 & ~A233;
  assign \new_[60070]_  = ~A232 & \new_[60069]_ ;
  assign \new_[60073]_  = ~A269 & ~A268;
  assign \new_[60076]_  = ~A300 & A298;
  assign \new_[60077]_  = \new_[60076]_  & \new_[60073]_ ;
  assign \new_[60078]_  = \new_[60077]_  & \new_[60070]_ ;
  assign \new_[60082]_  = A167 & ~A169;
  assign \new_[60083]_  = A170 & \new_[60082]_ ;
  assign \new_[60087]_  = ~A200 & ~A199;
  assign \new_[60088]_  = ~A166 & \new_[60087]_ ;
  assign \new_[60089]_  = \new_[60088]_  & \new_[60083]_ ;
  assign \new_[60093]_  = ~A266 & ~A233;
  assign \new_[60094]_  = ~A232 & \new_[60093]_ ;
  assign \new_[60097]_  = ~A269 & ~A268;
  assign \new_[60100]_  = A299 & A298;
  assign \new_[60101]_  = \new_[60100]_  & \new_[60097]_ ;
  assign \new_[60102]_  = \new_[60101]_  & \new_[60094]_ ;
  assign \new_[60106]_  = A167 & ~A169;
  assign \new_[60107]_  = A170 & \new_[60106]_ ;
  assign \new_[60111]_  = ~A200 & ~A199;
  assign \new_[60112]_  = ~A166 & \new_[60111]_ ;
  assign \new_[60113]_  = \new_[60112]_  & \new_[60107]_ ;
  assign \new_[60117]_  = ~A266 & ~A233;
  assign \new_[60118]_  = ~A232 & \new_[60117]_ ;
  assign \new_[60121]_  = ~A269 & ~A268;
  assign \new_[60124]_  = ~A299 & ~A298;
  assign \new_[60125]_  = \new_[60124]_  & \new_[60121]_ ;
  assign \new_[60126]_  = \new_[60125]_  & \new_[60118]_ ;
  assign \new_[60130]_  = A167 & ~A169;
  assign \new_[60131]_  = A170 & \new_[60130]_ ;
  assign \new_[60135]_  = ~A200 & ~A199;
  assign \new_[60136]_  = ~A166 & \new_[60135]_ ;
  assign \new_[60137]_  = \new_[60136]_  & \new_[60131]_ ;
  assign \new_[60141]_  = ~A266 & ~A233;
  assign \new_[60142]_  = ~A232 & \new_[60141]_ ;
  assign \new_[60145]_  = A298 & ~A267;
  assign \new_[60148]_  = ~A302 & ~A301;
  assign \new_[60149]_  = \new_[60148]_  & \new_[60145]_ ;
  assign \new_[60150]_  = \new_[60149]_  & \new_[60142]_ ;
  assign \new_[60154]_  = A167 & ~A169;
  assign \new_[60155]_  = A170 & \new_[60154]_ ;
  assign \new_[60159]_  = ~A200 & ~A199;
  assign \new_[60160]_  = ~A166 & \new_[60159]_ ;
  assign \new_[60161]_  = \new_[60160]_  & \new_[60155]_ ;
  assign \new_[60165]_  = ~A265 & ~A233;
  assign \new_[60166]_  = ~A232 & \new_[60165]_ ;
  assign \new_[60169]_  = A298 & ~A266;
  assign \new_[60172]_  = ~A302 & ~A301;
  assign \new_[60173]_  = \new_[60172]_  & \new_[60169]_ ;
  assign \new_[60174]_  = \new_[60173]_  & \new_[60166]_ ;
  assign \new_[60178]_  = ~A167 & ~A169;
  assign \new_[60179]_  = A170 & \new_[60178]_ ;
  assign \new_[60183]_  = A200 & A199;
  assign \new_[60184]_  = A166 & \new_[60183]_ ;
  assign \new_[60185]_  = \new_[60184]_  & \new_[60179]_ ;
  assign \new_[60189]_  = A265 & A233;
  assign \new_[60190]_  = A232 & \new_[60189]_ ;
  assign \new_[60193]_  = ~A269 & ~A268;
  assign \new_[60196]_  = ~A300 & ~A299;
  assign \new_[60197]_  = \new_[60196]_  & \new_[60193]_ ;
  assign \new_[60198]_  = \new_[60197]_  & \new_[60190]_ ;
  assign \new_[60202]_  = ~A167 & ~A169;
  assign \new_[60203]_  = A170 & \new_[60202]_ ;
  assign \new_[60207]_  = A200 & A199;
  assign \new_[60208]_  = A166 & \new_[60207]_ ;
  assign \new_[60209]_  = \new_[60208]_  & \new_[60203]_ ;
  assign \new_[60213]_  = A265 & A233;
  assign \new_[60214]_  = A232 & \new_[60213]_ ;
  assign \new_[60217]_  = ~A269 & ~A268;
  assign \new_[60220]_  = A299 & A298;
  assign \new_[60221]_  = \new_[60220]_  & \new_[60217]_ ;
  assign \new_[60222]_  = \new_[60221]_  & \new_[60214]_ ;
  assign \new_[60226]_  = ~A167 & ~A169;
  assign \new_[60227]_  = A170 & \new_[60226]_ ;
  assign \new_[60231]_  = A200 & A199;
  assign \new_[60232]_  = A166 & \new_[60231]_ ;
  assign \new_[60233]_  = \new_[60232]_  & \new_[60227]_ ;
  assign \new_[60237]_  = A265 & A233;
  assign \new_[60238]_  = A232 & \new_[60237]_ ;
  assign \new_[60241]_  = ~A269 & ~A268;
  assign \new_[60244]_  = ~A299 & ~A298;
  assign \new_[60245]_  = \new_[60244]_  & \new_[60241]_ ;
  assign \new_[60246]_  = \new_[60245]_  & \new_[60238]_ ;
  assign \new_[60250]_  = ~A167 & ~A169;
  assign \new_[60251]_  = A170 & \new_[60250]_ ;
  assign \new_[60255]_  = A200 & A199;
  assign \new_[60256]_  = A166 & \new_[60255]_ ;
  assign \new_[60257]_  = \new_[60256]_  & \new_[60251]_ ;
  assign \new_[60261]_  = A265 & A233;
  assign \new_[60262]_  = A232 & \new_[60261]_ ;
  assign \new_[60265]_  = ~A299 & ~A267;
  assign \new_[60268]_  = ~A302 & ~A301;
  assign \new_[60269]_  = \new_[60268]_  & \new_[60265]_ ;
  assign \new_[60270]_  = \new_[60269]_  & \new_[60262]_ ;
  assign \new_[60274]_  = ~A167 & ~A169;
  assign \new_[60275]_  = A170 & \new_[60274]_ ;
  assign \new_[60279]_  = A200 & A199;
  assign \new_[60280]_  = A166 & \new_[60279]_ ;
  assign \new_[60281]_  = \new_[60280]_  & \new_[60275]_ ;
  assign \new_[60285]_  = A265 & A233;
  assign \new_[60286]_  = A232 & \new_[60285]_ ;
  assign \new_[60289]_  = ~A299 & A266;
  assign \new_[60292]_  = ~A302 & ~A301;
  assign \new_[60293]_  = \new_[60292]_  & \new_[60289]_ ;
  assign \new_[60294]_  = \new_[60293]_  & \new_[60286]_ ;
  assign \new_[60298]_  = ~A167 & ~A169;
  assign \new_[60299]_  = A170 & \new_[60298]_ ;
  assign \new_[60303]_  = A200 & A199;
  assign \new_[60304]_  = A166 & \new_[60303]_ ;
  assign \new_[60305]_  = \new_[60304]_  & \new_[60299]_ ;
  assign \new_[60309]_  = ~A265 & A233;
  assign \new_[60310]_  = A232 & \new_[60309]_ ;
  assign \new_[60313]_  = ~A299 & ~A266;
  assign \new_[60316]_  = ~A302 & ~A301;
  assign \new_[60317]_  = \new_[60316]_  & \new_[60313]_ ;
  assign \new_[60318]_  = \new_[60317]_  & \new_[60310]_ ;
  assign \new_[60322]_  = ~A167 & ~A169;
  assign \new_[60323]_  = A170 & \new_[60322]_ ;
  assign \new_[60327]_  = A200 & A199;
  assign \new_[60328]_  = A166 & \new_[60327]_ ;
  assign \new_[60329]_  = \new_[60328]_  & \new_[60323]_ ;
  assign \new_[60333]_  = ~A236 & ~A235;
  assign \new_[60334]_  = ~A233 & \new_[60333]_ ;
  assign \new_[60337]_  = A266 & A265;
  assign \new_[60340]_  = ~A300 & A298;
  assign \new_[60341]_  = \new_[60340]_  & \new_[60337]_ ;
  assign \new_[60342]_  = \new_[60341]_  & \new_[60334]_ ;
  assign \new_[60346]_  = ~A167 & ~A169;
  assign \new_[60347]_  = A170 & \new_[60346]_ ;
  assign \new_[60351]_  = A200 & A199;
  assign \new_[60352]_  = A166 & \new_[60351]_ ;
  assign \new_[60353]_  = \new_[60352]_  & \new_[60347]_ ;
  assign \new_[60357]_  = ~A236 & ~A235;
  assign \new_[60358]_  = ~A233 & \new_[60357]_ ;
  assign \new_[60361]_  = A266 & A265;
  assign \new_[60364]_  = A299 & A298;
  assign \new_[60365]_  = \new_[60364]_  & \new_[60361]_ ;
  assign \new_[60366]_  = \new_[60365]_  & \new_[60358]_ ;
  assign \new_[60370]_  = ~A167 & ~A169;
  assign \new_[60371]_  = A170 & \new_[60370]_ ;
  assign \new_[60375]_  = A200 & A199;
  assign \new_[60376]_  = A166 & \new_[60375]_ ;
  assign \new_[60377]_  = \new_[60376]_  & \new_[60371]_ ;
  assign \new_[60381]_  = ~A236 & ~A235;
  assign \new_[60382]_  = ~A233 & \new_[60381]_ ;
  assign \new_[60385]_  = A266 & A265;
  assign \new_[60388]_  = ~A299 & ~A298;
  assign \new_[60389]_  = \new_[60388]_  & \new_[60385]_ ;
  assign \new_[60390]_  = \new_[60389]_  & \new_[60382]_ ;
  assign \new_[60394]_  = ~A167 & ~A169;
  assign \new_[60395]_  = A170 & \new_[60394]_ ;
  assign \new_[60399]_  = A200 & A199;
  assign \new_[60400]_  = A166 & \new_[60399]_ ;
  assign \new_[60401]_  = \new_[60400]_  & \new_[60395]_ ;
  assign \new_[60405]_  = ~A236 & ~A235;
  assign \new_[60406]_  = ~A233 & \new_[60405]_ ;
  assign \new_[60409]_  = ~A267 & ~A266;
  assign \new_[60412]_  = ~A300 & A298;
  assign \new_[60413]_  = \new_[60412]_  & \new_[60409]_ ;
  assign \new_[60414]_  = \new_[60413]_  & \new_[60406]_ ;
  assign \new_[60418]_  = ~A167 & ~A169;
  assign \new_[60419]_  = A170 & \new_[60418]_ ;
  assign \new_[60423]_  = A200 & A199;
  assign \new_[60424]_  = A166 & \new_[60423]_ ;
  assign \new_[60425]_  = \new_[60424]_  & \new_[60419]_ ;
  assign \new_[60429]_  = ~A236 & ~A235;
  assign \new_[60430]_  = ~A233 & \new_[60429]_ ;
  assign \new_[60433]_  = ~A267 & ~A266;
  assign \new_[60436]_  = A299 & A298;
  assign \new_[60437]_  = \new_[60436]_  & \new_[60433]_ ;
  assign \new_[60438]_  = \new_[60437]_  & \new_[60430]_ ;
  assign \new_[60442]_  = ~A167 & ~A169;
  assign \new_[60443]_  = A170 & \new_[60442]_ ;
  assign \new_[60447]_  = A200 & A199;
  assign \new_[60448]_  = A166 & \new_[60447]_ ;
  assign \new_[60449]_  = \new_[60448]_  & \new_[60443]_ ;
  assign \new_[60453]_  = ~A236 & ~A235;
  assign \new_[60454]_  = ~A233 & \new_[60453]_ ;
  assign \new_[60457]_  = ~A267 & ~A266;
  assign \new_[60460]_  = ~A299 & ~A298;
  assign \new_[60461]_  = \new_[60460]_  & \new_[60457]_ ;
  assign \new_[60462]_  = \new_[60461]_  & \new_[60454]_ ;
  assign \new_[60466]_  = ~A167 & ~A169;
  assign \new_[60467]_  = A170 & \new_[60466]_ ;
  assign \new_[60471]_  = A200 & A199;
  assign \new_[60472]_  = A166 & \new_[60471]_ ;
  assign \new_[60473]_  = \new_[60472]_  & \new_[60467]_ ;
  assign \new_[60477]_  = ~A236 & ~A235;
  assign \new_[60478]_  = ~A233 & \new_[60477]_ ;
  assign \new_[60481]_  = ~A266 & ~A265;
  assign \new_[60484]_  = ~A300 & A298;
  assign \new_[60485]_  = \new_[60484]_  & \new_[60481]_ ;
  assign \new_[60486]_  = \new_[60485]_  & \new_[60478]_ ;
  assign \new_[60490]_  = ~A167 & ~A169;
  assign \new_[60491]_  = A170 & \new_[60490]_ ;
  assign \new_[60495]_  = A200 & A199;
  assign \new_[60496]_  = A166 & \new_[60495]_ ;
  assign \new_[60497]_  = \new_[60496]_  & \new_[60491]_ ;
  assign \new_[60501]_  = ~A236 & ~A235;
  assign \new_[60502]_  = ~A233 & \new_[60501]_ ;
  assign \new_[60505]_  = ~A266 & ~A265;
  assign \new_[60508]_  = A299 & A298;
  assign \new_[60509]_  = \new_[60508]_  & \new_[60505]_ ;
  assign \new_[60510]_  = \new_[60509]_  & \new_[60502]_ ;
  assign \new_[60514]_  = ~A167 & ~A169;
  assign \new_[60515]_  = A170 & \new_[60514]_ ;
  assign \new_[60519]_  = A200 & A199;
  assign \new_[60520]_  = A166 & \new_[60519]_ ;
  assign \new_[60521]_  = \new_[60520]_  & \new_[60515]_ ;
  assign \new_[60525]_  = ~A236 & ~A235;
  assign \new_[60526]_  = ~A233 & \new_[60525]_ ;
  assign \new_[60529]_  = ~A266 & ~A265;
  assign \new_[60532]_  = ~A299 & ~A298;
  assign \new_[60533]_  = \new_[60532]_  & \new_[60529]_ ;
  assign \new_[60534]_  = \new_[60533]_  & \new_[60526]_ ;
  assign \new_[60538]_  = ~A167 & ~A169;
  assign \new_[60539]_  = A170 & \new_[60538]_ ;
  assign \new_[60543]_  = A200 & A199;
  assign \new_[60544]_  = A166 & \new_[60543]_ ;
  assign \new_[60545]_  = \new_[60544]_  & \new_[60539]_ ;
  assign \new_[60549]_  = A265 & ~A234;
  assign \new_[60550]_  = ~A233 & \new_[60549]_ ;
  assign \new_[60553]_  = A298 & A266;
  assign \new_[60556]_  = ~A302 & ~A301;
  assign \new_[60557]_  = \new_[60556]_  & \new_[60553]_ ;
  assign \new_[60558]_  = \new_[60557]_  & \new_[60550]_ ;
  assign \new_[60562]_  = ~A167 & ~A169;
  assign \new_[60563]_  = A170 & \new_[60562]_ ;
  assign \new_[60567]_  = A200 & A199;
  assign \new_[60568]_  = A166 & \new_[60567]_ ;
  assign \new_[60569]_  = \new_[60568]_  & \new_[60563]_ ;
  assign \new_[60573]_  = ~A266 & ~A234;
  assign \new_[60574]_  = ~A233 & \new_[60573]_ ;
  assign \new_[60577]_  = ~A269 & ~A268;
  assign \new_[60580]_  = ~A300 & A298;
  assign \new_[60581]_  = \new_[60580]_  & \new_[60577]_ ;
  assign \new_[60582]_  = \new_[60581]_  & \new_[60574]_ ;
  assign \new_[60586]_  = ~A167 & ~A169;
  assign \new_[60587]_  = A170 & \new_[60586]_ ;
  assign \new_[60591]_  = A200 & A199;
  assign \new_[60592]_  = A166 & \new_[60591]_ ;
  assign \new_[60593]_  = \new_[60592]_  & \new_[60587]_ ;
  assign \new_[60597]_  = ~A266 & ~A234;
  assign \new_[60598]_  = ~A233 & \new_[60597]_ ;
  assign \new_[60601]_  = ~A269 & ~A268;
  assign \new_[60604]_  = A299 & A298;
  assign \new_[60605]_  = \new_[60604]_  & \new_[60601]_ ;
  assign \new_[60606]_  = \new_[60605]_  & \new_[60598]_ ;
  assign \new_[60610]_  = ~A167 & ~A169;
  assign \new_[60611]_  = A170 & \new_[60610]_ ;
  assign \new_[60615]_  = A200 & A199;
  assign \new_[60616]_  = A166 & \new_[60615]_ ;
  assign \new_[60617]_  = \new_[60616]_  & \new_[60611]_ ;
  assign \new_[60621]_  = ~A266 & ~A234;
  assign \new_[60622]_  = ~A233 & \new_[60621]_ ;
  assign \new_[60625]_  = ~A269 & ~A268;
  assign \new_[60628]_  = ~A299 & ~A298;
  assign \new_[60629]_  = \new_[60628]_  & \new_[60625]_ ;
  assign \new_[60630]_  = \new_[60629]_  & \new_[60622]_ ;
  assign \new_[60634]_  = ~A167 & ~A169;
  assign \new_[60635]_  = A170 & \new_[60634]_ ;
  assign \new_[60639]_  = A200 & A199;
  assign \new_[60640]_  = A166 & \new_[60639]_ ;
  assign \new_[60641]_  = \new_[60640]_  & \new_[60635]_ ;
  assign \new_[60645]_  = ~A266 & ~A234;
  assign \new_[60646]_  = ~A233 & \new_[60645]_ ;
  assign \new_[60649]_  = A298 & ~A267;
  assign \new_[60652]_  = ~A302 & ~A301;
  assign \new_[60653]_  = \new_[60652]_  & \new_[60649]_ ;
  assign \new_[60654]_  = \new_[60653]_  & \new_[60646]_ ;
  assign \new_[60658]_  = ~A167 & ~A169;
  assign \new_[60659]_  = A170 & \new_[60658]_ ;
  assign \new_[60663]_  = A200 & A199;
  assign \new_[60664]_  = A166 & \new_[60663]_ ;
  assign \new_[60665]_  = \new_[60664]_  & \new_[60659]_ ;
  assign \new_[60669]_  = ~A265 & ~A234;
  assign \new_[60670]_  = ~A233 & \new_[60669]_ ;
  assign \new_[60673]_  = A298 & ~A266;
  assign \new_[60676]_  = ~A302 & ~A301;
  assign \new_[60677]_  = \new_[60676]_  & \new_[60673]_ ;
  assign \new_[60678]_  = \new_[60677]_  & \new_[60670]_ ;
  assign \new_[60682]_  = ~A167 & ~A169;
  assign \new_[60683]_  = A170 & \new_[60682]_ ;
  assign \new_[60687]_  = A200 & A199;
  assign \new_[60688]_  = A166 & \new_[60687]_ ;
  assign \new_[60689]_  = \new_[60688]_  & \new_[60683]_ ;
  assign \new_[60693]_  = A265 & ~A233;
  assign \new_[60694]_  = ~A232 & \new_[60693]_ ;
  assign \new_[60697]_  = A298 & A266;
  assign \new_[60700]_  = ~A302 & ~A301;
  assign \new_[60701]_  = \new_[60700]_  & \new_[60697]_ ;
  assign \new_[60702]_  = \new_[60701]_  & \new_[60694]_ ;
  assign \new_[60706]_  = ~A167 & ~A169;
  assign \new_[60707]_  = A170 & \new_[60706]_ ;
  assign \new_[60711]_  = A200 & A199;
  assign \new_[60712]_  = A166 & \new_[60711]_ ;
  assign \new_[60713]_  = \new_[60712]_  & \new_[60707]_ ;
  assign \new_[60717]_  = ~A266 & ~A233;
  assign \new_[60718]_  = ~A232 & \new_[60717]_ ;
  assign \new_[60721]_  = ~A269 & ~A268;
  assign \new_[60724]_  = ~A300 & A298;
  assign \new_[60725]_  = \new_[60724]_  & \new_[60721]_ ;
  assign \new_[60726]_  = \new_[60725]_  & \new_[60718]_ ;
  assign \new_[60730]_  = ~A167 & ~A169;
  assign \new_[60731]_  = A170 & \new_[60730]_ ;
  assign \new_[60735]_  = A200 & A199;
  assign \new_[60736]_  = A166 & \new_[60735]_ ;
  assign \new_[60737]_  = \new_[60736]_  & \new_[60731]_ ;
  assign \new_[60741]_  = ~A266 & ~A233;
  assign \new_[60742]_  = ~A232 & \new_[60741]_ ;
  assign \new_[60745]_  = ~A269 & ~A268;
  assign \new_[60748]_  = A299 & A298;
  assign \new_[60749]_  = \new_[60748]_  & \new_[60745]_ ;
  assign \new_[60750]_  = \new_[60749]_  & \new_[60742]_ ;
  assign \new_[60754]_  = ~A167 & ~A169;
  assign \new_[60755]_  = A170 & \new_[60754]_ ;
  assign \new_[60759]_  = A200 & A199;
  assign \new_[60760]_  = A166 & \new_[60759]_ ;
  assign \new_[60761]_  = \new_[60760]_  & \new_[60755]_ ;
  assign \new_[60765]_  = ~A266 & ~A233;
  assign \new_[60766]_  = ~A232 & \new_[60765]_ ;
  assign \new_[60769]_  = ~A269 & ~A268;
  assign \new_[60772]_  = ~A299 & ~A298;
  assign \new_[60773]_  = \new_[60772]_  & \new_[60769]_ ;
  assign \new_[60774]_  = \new_[60773]_  & \new_[60766]_ ;
  assign \new_[60778]_  = ~A167 & ~A169;
  assign \new_[60779]_  = A170 & \new_[60778]_ ;
  assign \new_[60783]_  = A200 & A199;
  assign \new_[60784]_  = A166 & \new_[60783]_ ;
  assign \new_[60785]_  = \new_[60784]_  & \new_[60779]_ ;
  assign \new_[60789]_  = ~A266 & ~A233;
  assign \new_[60790]_  = ~A232 & \new_[60789]_ ;
  assign \new_[60793]_  = A298 & ~A267;
  assign \new_[60796]_  = ~A302 & ~A301;
  assign \new_[60797]_  = \new_[60796]_  & \new_[60793]_ ;
  assign \new_[60798]_  = \new_[60797]_  & \new_[60790]_ ;
  assign \new_[60802]_  = ~A167 & ~A169;
  assign \new_[60803]_  = A170 & \new_[60802]_ ;
  assign \new_[60807]_  = A200 & A199;
  assign \new_[60808]_  = A166 & \new_[60807]_ ;
  assign \new_[60809]_  = \new_[60808]_  & \new_[60803]_ ;
  assign \new_[60813]_  = ~A265 & ~A233;
  assign \new_[60814]_  = ~A232 & \new_[60813]_ ;
  assign \new_[60817]_  = A298 & ~A266;
  assign \new_[60820]_  = ~A302 & ~A301;
  assign \new_[60821]_  = \new_[60820]_  & \new_[60817]_ ;
  assign \new_[60822]_  = \new_[60821]_  & \new_[60814]_ ;
  assign \new_[60826]_  = ~A167 & ~A169;
  assign \new_[60827]_  = A170 & \new_[60826]_ ;
  assign \new_[60831]_  = ~A202 & ~A200;
  assign \new_[60832]_  = A166 & \new_[60831]_ ;
  assign \new_[60833]_  = \new_[60832]_  & \new_[60827]_ ;
  assign \new_[60837]_  = A233 & A232;
  assign \new_[60838]_  = ~A203 & \new_[60837]_ ;
  assign \new_[60841]_  = ~A267 & A265;
  assign \new_[60844]_  = ~A300 & ~A299;
  assign \new_[60845]_  = \new_[60844]_  & \new_[60841]_ ;
  assign \new_[60846]_  = \new_[60845]_  & \new_[60838]_ ;
  assign \new_[60850]_  = ~A167 & ~A169;
  assign \new_[60851]_  = A170 & \new_[60850]_ ;
  assign \new_[60855]_  = ~A202 & ~A200;
  assign \new_[60856]_  = A166 & \new_[60855]_ ;
  assign \new_[60857]_  = \new_[60856]_  & \new_[60851]_ ;
  assign \new_[60861]_  = A233 & A232;
  assign \new_[60862]_  = ~A203 & \new_[60861]_ ;
  assign \new_[60865]_  = ~A267 & A265;
  assign \new_[60868]_  = A299 & A298;
  assign \new_[60869]_  = \new_[60868]_  & \new_[60865]_ ;
  assign \new_[60870]_  = \new_[60869]_  & \new_[60862]_ ;
  assign \new_[60874]_  = ~A167 & ~A169;
  assign \new_[60875]_  = A170 & \new_[60874]_ ;
  assign \new_[60879]_  = ~A202 & ~A200;
  assign \new_[60880]_  = A166 & \new_[60879]_ ;
  assign \new_[60881]_  = \new_[60880]_  & \new_[60875]_ ;
  assign \new_[60885]_  = A233 & A232;
  assign \new_[60886]_  = ~A203 & \new_[60885]_ ;
  assign \new_[60889]_  = ~A267 & A265;
  assign \new_[60892]_  = ~A299 & ~A298;
  assign \new_[60893]_  = \new_[60892]_  & \new_[60889]_ ;
  assign \new_[60894]_  = \new_[60893]_  & \new_[60886]_ ;
  assign \new_[60898]_  = ~A167 & ~A169;
  assign \new_[60899]_  = A170 & \new_[60898]_ ;
  assign \new_[60903]_  = ~A202 & ~A200;
  assign \new_[60904]_  = A166 & \new_[60903]_ ;
  assign \new_[60905]_  = \new_[60904]_  & \new_[60899]_ ;
  assign \new_[60909]_  = A233 & A232;
  assign \new_[60910]_  = ~A203 & \new_[60909]_ ;
  assign \new_[60913]_  = A266 & A265;
  assign \new_[60916]_  = ~A300 & ~A299;
  assign \new_[60917]_  = \new_[60916]_  & \new_[60913]_ ;
  assign \new_[60918]_  = \new_[60917]_  & \new_[60910]_ ;
  assign \new_[60922]_  = ~A167 & ~A169;
  assign \new_[60923]_  = A170 & \new_[60922]_ ;
  assign \new_[60927]_  = ~A202 & ~A200;
  assign \new_[60928]_  = A166 & \new_[60927]_ ;
  assign \new_[60929]_  = \new_[60928]_  & \new_[60923]_ ;
  assign \new_[60933]_  = A233 & A232;
  assign \new_[60934]_  = ~A203 & \new_[60933]_ ;
  assign \new_[60937]_  = A266 & A265;
  assign \new_[60940]_  = A299 & A298;
  assign \new_[60941]_  = \new_[60940]_  & \new_[60937]_ ;
  assign \new_[60942]_  = \new_[60941]_  & \new_[60934]_ ;
  assign \new_[60946]_  = ~A167 & ~A169;
  assign \new_[60947]_  = A170 & \new_[60946]_ ;
  assign \new_[60951]_  = ~A202 & ~A200;
  assign \new_[60952]_  = A166 & \new_[60951]_ ;
  assign \new_[60953]_  = \new_[60952]_  & \new_[60947]_ ;
  assign \new_[60957]_  = A233 & A232;
  assign \new_[60958]_  = ~A203 & \new_[60957]_ ;
  assign \new_[60961]_  = A266 & A265;
  assign \new_[60964]_  = ~A299 & ~A298;
  assign \new_[60965]_  = \new_[60964]_  & \new_[60961]_ ;
  assign \new_[60966]_  = \new_[60965]_  & \new_[60958]_ ;
  assign \new_[60970]_  = ~A167 & ~A169;
  assign \new_[60971]_  = A170 & \new_[60970]_ ;
  assign \new_[60975]_  = ~A202 & ~A200;
  assign \new_[60976]_  = A166 & \new_[60975]_ ;
  assign \new_[60977]_  = \new_[60976]_  & \new_[60971]_ ;
  assign \new_[60981]_  = A233 & A232;
  assign \new_[60982]_  = ~A203 & \new_[60981]_ ;
  assign \new_[60985]_  = ~A266 & ~A265;
  assign \new_[60988]_  = ~A300 & ~A299;
  assign \new_[60989]_  = \new_[60988]_  & \new_[60985]_ ;
  assign \new_[60990]_  = \new_[60989]_  & \new_[60982]_ ;
  assign \new_[60994]_  = ~A167 & ~A169;
  assign \new_[60995]_  = A170 & \new_[60994]_ ;
  assign \new_[60999]_  = ~A202 & ~A200;
  assign \new_[61000]_  = A166 & \new_[60999]_ ;
  assign \new_[61001]_  = \new_[61000]_  & \new_[60995]_ ;
  assign \new_[61005]_  = A233 & A232;
  assign \new_[61006]_  = ~A203 & \new_[61005]_ ;
  assign \new_[61009]_  = ~A266 & ~A265;
  assign \new_[61012]_  = A299 & A298;
  assign \new_[61013]_  = \new_[61012]_  & \new_[61009]_ ;
  assign \new_[61014]_  = \new_[61013]_  & \new_[61006]_ ;
  assign \new_[61018]_  = ~A167 & ~A169;
  assign \new_[61019]_  = A170 & \new_[61018]_ ;
  assign \new_[61023]_  = ~A202 & ~A200;
  assign \new_[61024]_  = A166 & \new_[61023]_ ;
  assign \new_[61025]_  = \new_[61024]_  & \new_[61019]_ ;
  assign \new_[61029]_  = A233 & A232;
  assign \new_[61030]_  = ~A203 & \new_[61029]_ ;
  assign \new_[61033]_  = ~A266 & ~A265;
  assign \new_[61036]_  = ~A299 & ~A298;
  assign \new_[61037]_  = \new_[61036]_  & \new_[61033]_ ;
  assign \new_[61038]_  = \new_[61037]_  & \new_[61030]_ ;
  assign \new_[61042]_  = ~A167 & ~A169;
  assign \new_[61043]_  = A170 & \new_[61042]_ ;
  assign \new_[61047]_  = ~A202 & ~A200;
  assign \new_[61048]_  = A166 & \new_[61047]_ ;
  assign \new_[61049]_  = \new_[61048]_  & \new_[61043]_ ;
  assign \new_[61053]_  = A233 & ~A232;
  assign \new_[61054]_  = ~A203 & \new_[61053]_ ;
  assign \new_[61057]_  = ~A299 & A298;
  assign \new_[61060]_  = A301 & A300;
  assign \new_[61061]_  = \new_[61060]_  & \new_[61057]_ ;
  assign \new_[61062]_  = \new_[61061]_  & \new_[61054]_ ;
  assign \new_[61066]_  = ~A167 & ~A169;
  assign \new_[61067]_  = A170 & \new_[61066]_ ;
  assign \new_[61071]_  = ~A202 & ~A200;
  assign \new_[61072]_  = A166 & \new_[61071]_ ;
  assign \new_[61073]_  = \new_[61072]_  & \new_[61067]_ ;
  assign \new_[61077]_  = A233 & ~A232;
  assign \new_[61078]_  = ~A203 & \new_[61077]_ ;
  assign \new_[61081]_  = ~A299 & A298;
  assign \new_[61084]_  = A302 & A300;
  assign \new_[61085]_  = \new_[61084]_  & \new_[61081]_ ;
  assign \new_[61086]_  = \new_[61085]_  & \new_[61078]_ ;
  assign \new_[61090]_  = ~A167 & ~A169;
  assign \new_[61091]_  = A170 & \new_[61090]_ ;
  assign \new_[61095]_  = ~A202 & ~A200;
  assign \new_[61096]_  = A166 & \new_[61095]_ ;
  assign \new_[61097]_  = \new_[61096]_  & \new_[61091]_ ;
  assign \new_[61101]_  = A233 & ~A232;
  assign \new_[61102]_  = ~A203 & \new_[61101]_ ;
  assign \new_[61105]_  = ~A266 & A265;
  assign \new_[61108]_  = A268 & A267;
  assign \new_[61109]_  = \new_[61108]_  & \new_[61105]_ ;
  assign \new_[61110]_  = \new_[61109]_  & \new_[61102]_ ;
  assign \new_[61114]_  = ~A167 & ~A169;
  assign \new_[61115]_  = A170 & \new_[61114]_ ;
  assign \new_[61119]_  = ~A202 & ~A200;
  assign \new_[61120]_  = A166 & \new_[61119]_ ;
  assign \new_[61121]_  = \new_[61120]_  & \new_[61115]_ ;
  assign \new_[61125]_  = A233 & ~A232;
  assign \new_[61126]_  = ~A203 & \new_[61125]_ ;
  assign \new_[61129]_  = ~A266 & A265;
  assign \new_[61132]_  = A269 & A267;
  assign \new_[61133]_  = \new_[61132]_  & \new_[61129]_ ;
  assign \new_[61134]_  = \new_[61133]_  & \new_[61126]_ ;
  assign \new_[61138]_  = ~A167 & ~A169;
  assign \new_[61139]_  = A170 & \new_[61138]_ ;
  assign \new_[61143]_  = ~A202 & ~A200;
  assign \new_[61144]_  = A166 & \new_[61143]_ ;
  assign \new_[61145]_  = \new_[61144]_  & \new_[61139]_ ;
  assign \new_[61149]_  = ~A234 & ~A233;
  assign \new_[61150]_  = ~A203 & \new_[61149]_ ;
  assign \new_[61153]_  = A266 & A265;
  assign \new_[61156]_  = ~A300 & A298;
  assign \new_[61157]_  = \new_[61156]_  & \new_[61153]_ ;
  assign \new_[61158]_  = \new_[61157]_  & \new_[61150]_ ;
  assign \new_[61162]_  = ~A167 & ~A169;
  assign \new_[61163]_  = A170 & \new_[61162]_ ;
  assign \new_[61167]_  = ~A202 & ~A200;
  assign \new_[61168]_  = A166 & \new_[61167]_ ;
  assign \new_[61169]_  = \new_[61168]_  & \new_[61163]_ ;
  assign \new_[61173]_  = ~A234 & ~A233;
  assign \new_[61174]_  = ~A203 & \new_[61173]_ ;
  assign \new_[61177]_  = A266 & A265;
  assign \new_[61180]_  = A299 & A298;
  assign \new_[61181]_  = \new_[61180]_  & \new_[61177]_ ;
  assign \new_[61182]_  = \new_[61181]_  & \new_[61174]_ ;
  assign \new_[61186]_  = ~A167 & ~A169;
  assign \new_[61187]_  = A170 & \new_[61186]_ ;
  assign \new_[61191]_  = ~A202 & ~A200;
  assign \new_[61192]_  = A166 & \new_[61191]_ ;
  assign \new_[61193]_  = \new_[61192]_  & \new_[61187]_ ;
  assign \new_[61197]_  = ~A234 & ~A233;
  assign \new_[61198]_  = ~A203 & \new_[61197]_ ;
  assign \new_[61201]_  = A266 & A265;
  assign \new_[61204]_  = ~A299 & ~A298;
  assign \new_[61205]_  = \new_[61204]_  & \new_[61201]_ ;
  assign \new_[61206]_  = \new_[61205]_  & \new_[61198]_ ;
  assign \new_[61210]_  = ~A167 & ~A169;
  assign \new_[61211]_  = A170 & \new_[61210]_ ;
  assign \new_[61215]_  = ~A202 & ~A200;
  assign \new_[61216]_  = A166 & \new_[61215]_ ;
  assign \new_[61217]_  = \new_[61216]_  & \new_[61211]_ ;
  assign \new_[61221]_  = ~A234 & ~A233;
  assign \new_[61222]_  = ~A203 & \new_[61221]_ ;
  assign \new_[61225]_  = ~A267 & ~A266;
  assign \new_[61228]_  = ~A300 & A298;
  assign \new_[61229]_  = \new_[61228]_  & \new_[61225]_ ;
  assign \new_[61230]_  = \new_[61229]_  & \new_[61222]_ ;
  assign \new_[61234]_  = ~A167 & ~A169;
  assign \new_[61235]_  = A170 & \new_[61234]_ ;
  assign \new_[61239]_  = ~A202 & ~A200;
  assign \new_[61240]_  = A166 & \new_[61239]_ ;
  assign \new_[61241]_  = \new_[61240]_  & \new_[61235]_ ;
  assign \new_[61245]_  = ~A234 & ~A233;
  assign \new_[61246]_  = ~A203 & \new_[61245]_ ;
  assign \new_[61249]_  = ~A267 & ~A266;
  assign \new_[61252]_  = A299 & A298;
  assign \new_[61253]_  = \new_[61252]_  & \new_[61249]_ ;
  assign \new_[61254]_  = \new_[61253]_  & \new_[61246]_ ;
  assign \new_[61258]_  = ~A167 & ~A169;
  assign \new_[61259]_  = A170 & \new_[61258]_ ;
  assign \new_[61263]_  = ~A202 & ~A200;
  assign \new_[61264]_  = A166 & \new_[61263]_ ;
  assign \new_[61265]_  = \new_[61264]_  & \new_[61259]_ ;
  assign \new_[61269]_  = ~A234 & ~A233;
  assign \new_[61270]_  = ~A203 & \new_[61269]_ ;
  assign \new_[61273]_  = ~A267 & ~A266;
  assign \new_[61276]_  = ~A299 & ~A298;
  assign \new_[61277]_  = \new_[61276]_  & \new_[61273]_ ;
  assign \new_[61278]_  = \new_[61277]_  & \new_[61270]_ ;
  assign \new_[61282]_  = ~A167 & ~A169;
  assign \new_[61283]_  = A170 & \new_[61282]_ ;
  assign \new_[61287]_  = ~A202 & ~A200;
  assign \new_[61288]_  = A166 & \new_[61287]_ ;
  assign \new_[61289]_  = \new_[61288]_  & \new_[61283]_ ;
  assign \new_[61293]_  = ~A234 & ~A233;
  assign \new_[61294]_  = ~A203 & \new_[61293]_ ;
  assign \new_[61297]_  = ~A266 & ~A265;
  assign \new_[61300]_  = ~A300 & A298;
  assign \new_[61301]_  = \new_[61300]_  & \new_[61297]_ ;
  assign \new_[61302]_  = \new_[61301]_  & \new_[61294]_ ;
  assign \new_[61306]_  = ~A167 & ~A169;
  assign \new_[61307]_  = A170 & \new_[61306]_ ;
  assign \new_[61311]_  = ~A202 & ~A200;
  assign \new_[61312]_  = A166 & \new_[61311]_ ;
  assign \new_[61313]_  = \new_[61312]_  & \new_[61307]_ ;
  assign \new_[61317]_  = ~A234 & ~A233;
  assign \new_[61318]_  = ~A203 & \new_[61317]_ ;
  assign \new_[61321]_  = ~A266 & ~A265;
  assign \new_[61324]_  = A299 & A298;
  assign \new_[61325]_  = \new_[61324]_  & \new_[61321]_ ;
  assign \new_[61326]_  = \new_[61325]_  & \new_[61318]_ ;
  assign \new_[61330]_  = ~A167 & ~A169;
  assign \new_[61331]_  = A170 & \new_[61330]_ ;
  assign \new_[61335]_  = ~A202 & ~A200;
  assign \new_[61336]_  = A166 & \new_[61335]_ ;
  assign \new_[61337]_  = \new_[61336]_  & \new_[61331]_ ;
  assign \new_[61341]_  = ~A234 & ~A233;
  assign \new_[61342]_  = ~A203 & \new_[61341]_ ;
  assign \new_[61345]_  = ~A266 & ~A265;
  assign \new_[61348]_  = ~A299 & ~A298;
  assign \new_[61349]_  = \new_[61348]_  & \new_[61345]_ ;
  assign \new_[61350]_  = \new_[61349]_  & \new_[61342]_ ;
  assign \new_[61354]_  = ~A167 & ~A169;
  assign \new_[61355]_  = A170 & \new_[61354]_ ;
  assign \new_[61359]_  = ~A202 & ~A200;
  assign \new_[61360]_  = A166 & \new_[61359]_ ;
  assign \new_[61361]_  = \new_[61360]_  & \new_[61355]_ ;
  assign \new_[61365]_  = ~A233 & A232;
  assign \new_[61366]_  = ~A203 & \new_[61365]_ ;
  assign \new_[61369]_  = A235 & A234;
  assign \new_[61372]_  = A299 & ~A298;
  assign \new_[61373]_  = \new_[61372]_  & \new_[61369]_ ;
  assign \new_[61374]_  = \new_[61373]_  & \new_[61366]_ ;
  assign \new_[61378]_  = ~A167 & ~A169;
  assign \new_[61379]_  = A170 & \new_[61378]_ ;
  assign \new_[61383]_  = ~A202 & ~A200;
  assign \new_[61384]_  = A166 & \new_[61383]_ ;
  assign \new_[61385]_  = \new_[61384]_  & \new_[61379]_ ;
  assign \new_[61389]_  = ~A233 & A232;
  assign \new_[61390]_  = ~A203 & \new_[61389]_ ;
  assign \new_[61393]_  = A235 & A234;
  assign \new_[61396]_  = A266 & ~A265;
  assign \new_[61397]_  = \new_[61396]_  & \new_[61393]_ ;
  assign \new_[61398]_  = \new_[61397]_  & \new_[61390]_ ;
  assign \new_[61402]_  = ~A167 & ~A169;
  assign \new_[61403]_  = A170 & \new_[61402]_ ;
  assign \new_[61407]_  = ~A202 & ~A200;
  assign \new_[61408]_  = A166 & \new_[61407]_ ;
  assign \new_[61409]_  = \new_[61408]_  & \new_[61403]_ ;
  assign \new_[61413]_  = ~A233 & A232;
  assign \new_[61414]_  = ~A203 & \new_[61413]_ ;
  assign \new_[61417]_  = A236 & A234;
  assign \new_[61420]_  = A299 & ~A298;
  assign \new_[61421]_  = \new_[61420]_  & \new_[61417]_ ;
  assign \new_[61422]_  = \new_[61421]_  & \new_[61414]_ ;
  assign \new_[61426]_  = ~A167 & ~A169;
  assign \new_[61427]_  = A170 & \new_[61426]_ ;
  assign \new_[61431]_  = ~A202 & ~A200;
  assign \new_[61432]_  = A166 & \new_[61431]_ ;
  assign \new_[61433]_  = \new_[61432]_  & \new_[61427]_ ;
  assign \new_[61437]_  = ~A233 & A232;
  assign \new_[61438]_  = ~A203 & \new_[61437]_ ;
  assign \new_[61441]_  = A236 & A234;
  assign \new_[61444]_  = A266 & ~A265;
  assign \new_[61445]_  = \new_[61444]_  & \new_[61441]_ ;
  assign \new_[61446]_  = \new_[61445]_  & \new_[61438]_ ;
  assign \new_[61450]_  = ~A167 & ~A169;
  assign \new_[61451]_  = A170 & \new_[61450]_ ;
  assign \new_[61455]_  = ~A202 & ~A200;
  assign \new_[61456]_  = A166 & \new_[61455]_ ;
  assign \new_[61457]_  = \new_[61456]_  & \new_[61451]_ ;
  assign \new_[61461]_  = ~A233 & ~A232;
  assign \new_[61462]_  = ~A203 & \new_[61461]_ ;
  assign \new_[61465]_  = A266 & A265;
  assign \new_[61468]_  = ~A300 & A298;
  assign \new_[61469]_  = \new_[61468]_  & \new_[61465]_ ;
  assign \new_[61470]_  = \new_[61469]_  & \new_[61462]_ ;
  assign \new_[61474]_  = ~A167 & ~A169;
  assign \new_[61475]_  = A170 & \new_[61474]_ ;
  assign \new_[61479]_  = ~A202 & ~A200;
  assign \new_[61480]_  = A166 & \new_[61479]_ ;
  assign \new_[61481]_  = \new_[61480]_  & \new_[61475]_ ;
  assign \new_[61485]_  = ~A233 & ~A232;
  assign \new_[61486]_  = ~A203 & \new_[61485]_ ;
  assign \new_[61489]_  = A266 & A265;
  assign \new_[61492]_  = A299 & A298;
  assign \new_[61493]_  = \new_[61492]_  & \new_[61489]_ ;
  assign \new_[61494]_  = \new_[61493]_  & \new_[61486]_ ;
  assign \new_[61498]_  = ~A167 & ~A169;
  assign \new_[61499]_  = A170 & \new_[61498]_ ;
  assign \new_[61503]_  = ~A202 & ~A200;
  assign \new_[61504]_  = A166 & \new_[61503]_ ;
  assign \new_[61505]_  = \new_[61504]_  & \new_[61499]_ ;
  assign \new_[61509]_  = ~A233 & ~A232;
  assign \new_[61510]_  = ~A203 & \new_[61509]_ ;
  assign \new_[61513]_  = A266 & A265;
  assign \new_[61516]_  = ~A299 & ~A298;
  assign \new_[61517]_  = \new_[61516]_  & \new_[61513]_ ;
  assign \new_[61518]_  = \new_[61517]_  & \new_[61510]_ ;
  assign \new_[61522]_  = ~A167 & ~A169;
  assign \new_[61523]_  = A170 & \new_[61522]_ ;
  assign \new_[61527]_  = ~A202 & ~A200;
  assign \new_[61528]_  = A166 & \new_[61527]_ ;
  assign \new_[61529]_  = \new_[61528]_  & \new_[61523]_ ;
  assign \new_[61533]_  = ~A233 & ~A232;
  assign \new_[61534]_  = ~A203 & \new_[61533]_ ;
  assign \new_[61537]_  = ~A267 & ~A266;
  assign \new_[61540]_  = ~A300 & A298;
  assign \new_[61541]_  = \new_[61540]_  & \new_[61537]_ ;
  assign \new_[61542]_  = \new_[61541]_  & \new_[61534]_ ;
  assign \new_[61546]_  = ~A167 & ~A169;
  assign \new_[61547]_  = A170 & \new_[61546]_ ;
  assign \new_[61551]_  = ~A202 & ~A200;
  assign \new_[61552]_  = A166 & \new_[61551]_ ;
  assign \new_[61553]_  = \new_[61552]_  & \new_[61547]_ ;
  assign \new_[61557]_  = ~A233 & ~A232;
  assign \new_[61558]_  = ~A203 & \new_[61557]_ ;
  assign \new_[61561]_  = ~A267 & ~A266;
  assign \new_[61564]_  = A299 & A298;
  assign \new_[61565]_  = \new_[61564]_  & \new_[61561]_ ;
  assign \new_[61566]_  = \new_[61565]_  & \new_[61558]_ ;
  assign \new_[61570]_  = ~A167 & ~A169;
  assign \new_[61571]_  = A170 & \new_[61570]_ ;
  assign \new_[61575]_  = ~A202 & ~A200;
  assign \new_[61576]_  = A166 & \new_[61575]_ ;
  assign \new_[61577]_  = \new_[61576]_  & \new_[61571]_ ;
  assign \new_[61581]_  = ~A233 & ~A232;
  assign \new_[61582]_  = ~A203 & \new_[61581]_ ;
  assign \new_[61585]_  = ~A267 & ~A266;
  assign \new_[61588]_  = ~A299 & ~A298;
  assign \new_[61589]_  = \new_[61588]_  & \new_[61585]_ ;
  assign \new_[61590]_  = \new_[61589]_  & \new_[61582]_ ;
  assign \new_[61594]_  = ~A167 & ~A169;
  assign \new_[61595]_  = A170 & \new_[61594]_ ;
  assign \new_[61599]_  = ~A202 & ~A200;
  assign \new_[61600]_  = A166 & \new_[61599]_ ;
  assign \new_[61601]_  = \new_[61600]_  & \new_[61595]_ ;
  assign \new_[61605]_  = ~A233 & ~A232;
  assign \new_[61606]_  = ~A203 & \new_[61605]_ ;
  assign \new_[61609]_  = ~A266 & ~A265;
  assign \new_[61612]_  = ~A300 & A298;
  assign \new_[61613]_  = \new_[61612]_  & \new_[61609]_ ;
  assign \new_[61614]_  = \new_[61613]_  & \new_[61606]_ ;
  assign \new_[61618]_  = ~A167 & ~A169;
  assign \new_[61619]_  = A170 & \new_[61618]_ ;
  assign \new_[61623]_  = ~A202 & ~A200;
  assign \new_[61624]_  = A166 & \new_[61623]_ ;
  assign \new_[61625]_  = \new_[61624]_  & \new_[61619]_ ;
  assign \new_[61629]_  = ~A233 & ~A232;
  assign \new_[61630]_  = ~A203 & \new_[61629]_ ;
  assign \new_[61633]_  = ~A266 & ~A265;
  assign \new_[61636]_  = A299 & A298;
  assign \new_[61637]_  = \new_[61636]_  & \new_[61633]_ ;
  assign \new_[61638]_  = \new_[61637]_  & \new_[61630]_ ;
  assign \new_[61642]_  = ~A167 & ~A169;
  assign \new_[61643]_  = A170 & \new_[61642]_ ;
  assign \new_[61647]_  = ~A202 & ~A200;
  assign \new_[61648]_  = A166 & \new_[61647]_ ;
  assign \new_[61649]_  = \new_[61648]_  & \new_[61643]_ ;
  assign \new_[61653]_  = ~A233 & ~A232;
  assign \new_[61654]_  = ~A203 & \new_[61653]_ ;
  assign \new_[61657]_  = ~A266 & ~A265;
  assign \new_[61660]_  = ~A299 & ~A298;
  assign \new_[61661]_  = \new_[61660]_  & \new_[61657]_ ;
  assign \new_[61662]_  = \new_[61661]_  & \new_[61654]_ ;
  assign \new_[61666]_  = ~A167 & ~A169;
  assign \new_[61667]_  = A170 & \new_[61666]_ ;
  assign \new_[61671]_  = ~A201 & ~A200;
  assign \new_[61672]_  = A166 & \new_[61671]_ ;
  assign \new_[61673]_  = \new_[61672]_  & \new_[61667]_ ;
  assign \new_[61677]_  = A265 & A233;
  assign \new_[61678]_  = A232 & \new_[61677]_ ;
  assign \new_[61681]_  = ~A269 & ~A268;
  assign \new_[61684]_  = ~A300 & ~A299;
  assign \new_[61685]_  = \new_[61684]_  & \new_[61681]_ ;
  assign \new_[61686]_  = \new_[61685]_  & \new_[61678]_ ;
  assign \new_[61690]_  = ~A167 & ~A169;
  assign \new_[61691]_  = A170 & \new_[61690]_ ;
  assign \new_[61695]_  = ~A201 & ~A200;
  assign \new_[61696]_  = A166 & \new_[61695]_ ;
  assign \new_[61697]_  = \new_[61696]_  & \new_[61691]_ ;
  assign \new_[61701]_  = A265 & A233;
  assign \new_[61702]_  = A232 & \new_[61701]_ ;
  assign \new_[61705]_  = ~A269 & ~A268;
  assign \new_[61708]_  = A299 & A298;
  assign \new_[61709]_  = \new_[61708]_  & \new_[61705]_ ;
  assign \new_[61710]_  = \new_[61709]_  & \new_[61702]_ ;
  assign \new_[61714]_  = ~A167 & ~A169;
  assign \new_[61715]_  = A170 & \new_[61714]_ ;
  assign \new_[61719]_  = ~A201 & ~A200;
  assign \new_[61720]_  = A166 & \new_[61719]_ ;
  assign \new_[61721]_  = \new_[61720]_  & \new_[61715]_ ;
  assign \new_[61725]_  = A265 & A233;
  assign \new_[61726]_  = A232 & \new_[61725]_ ;
  assign \new_[61729]_  = ~A269 & ~A268;
  assign \new_[61732]_  = ~A299 & ~A298;
  assign \new_[61733]_  = \new_[61732]_  & \new_[61729]_ ;
  assign \new_[61734]_  = \new_[61733]_  & \new_[61726]_ ;
  assign \new_[61738]_  = ~A167 & ~A169;
  assign \new_[61739]_  = A170 & \new_[61738]_ ;
  assign \new_[61743]_  = ~A201 & ~A200;
  assign \new_[61744]_  = A166 & \new_[61743]_ ;
  assign \new_[61745]_  = \new_[61744]_  & \new_[61739]_ ;
  assign \new_[61749]_  = A265 & A233;
  assign \new_[61750]_  = A232 & \new_[61749]_ ;
  assign \new_[61753]_  = ~A299 & ~A267;
  assign \new_[61756]_  = ~A302 & ~A301;
  assign \new_[61757]_  = \new_[61756]_  & \new_[61753]_ ;
  assign \new_[61758]_  = \new_[61757]_  & \new_[61750]_ ;
  assign \new_[61762]_  = ~A167 & ~A169;
  assign \new_[61763]_  = A170 & \new_[61762]_ ;
  assign \new_[61767]_  = ~A201 & ~A200;
  assign \new_[61768]_  = A166 & \new_[61767]_ ;
  assign \new_[61769]_  = \new_[61768]_  & \new_[61763]_ ;
  assign \new_[61773]_  = A265 & A233;
  assign \new_[61774]_  = A232 & \new_[61773]_ ;
  assign \new_[61777]_  = ~A299 & A266;
  assign \new_[61780]_  = ~A302 & ~A301;
  assign \new_[61781]_  = \new_[61780]_  & \new_[61777]_ ;
  assign \new_[61782]_  = \new_[61781]_  & \new_[61774]_ ;
  assign \new_[61786]_  = ~A167 & ~A169;
  assign \new_[61787]_  = A170 & \new_[61786]_ ;
  assign \new_[61791]_  = ~A201 & ~A200;
  assign \new_[61792]_  = A166 & \new_[61791]_ ;
  assign \new_[61793]_  = \new_[61792]_  & \new_[61787]_ ;
  assign \new_[61797]_  = ~A265 & A233;
  assign \new_[61798]_  = A232 & \new_[61797]_ ;
  assign \new_[61801]_  = ~A299 & ~A266;
  assign \new_[61804]_  = ~A302 & ~A301;
  assign \new_[61805]_  = \new_[61804]_  & \new_[61801]_ ;
  assign \new_[61806]_  = \new_[61805]_  & \new_[61798]_ ;
  assign \new_[61810]_  = ~A167 & ~A169;
  assign \new_[61811]_  = A170 & \new_[61810]_ ;
  assign \new_[61815]_  = ~A201 & ~A200;
  assign \new_[61816]_  = A166 & \new_[61815]_ ;
  assign \new_[61817]_  = \new_[61816]_  & \new_[61811]_ ;
  assign \new_[61821]_  = ~A236 & ~A235;
  assign \new_[61822]_  = ~A233 & \new_[61821]_ ;
  assign \new_[61825]_  = A266 & A265;
  assign \new_[61828]_  = ~A300 & A298;
  assign \new_[61829]_  = \new_[61828]_  & \new_[61825]_ ;
  assign \new_[61830]_  = \new_[61829]_  & \new_[61822]_ ;
  assign \new_[61834]_  = ~A167 & ~A169;
  assign \new_[61835]_  = A170 & \new_[61834]_ ;
  assign \new_[61839]_  = ~A201 & ~A200;
  assign \new_[61840]_  = A166 & \new_[61839]_ ;
  assign \new_[61841]_  = \new_[61840]_  & \new_[61835]_ ;
  assign \new_[61845]_  = ~A236 & ~A235;
  assign \new_[61846]_  = ~A233 & \new_[61845]_ ;
  assign \new_[61849]_  = A266 & A265;
  assign \new_[61852]_  = A299 & A298;
  assign \new_[61853]_  = \new_[61852]_  & \new_[61849]_ ;
  assign \new_[61854]_  = \new_[61853]_  & \new_[61846]_ ;
  assign \new_[61858]_  = ~A167 & ~A169;
  assign \new_[61859]_  = A170 & \new_[61858]_ ;
  assign \new_[61863]_  = ~A201 & ~A200;
  assign \new_[61864]_  = A166 & \new_[61863]_ ;
  assign \new_[61865]_  = \new_[61864]_  & \new_[61859]_ ;
  assign \new_[61869]_  = ~A236 & ~A235;
  assign \new_[61870]_  = ~A233 & \new_[61869]_ ;
  assign \new_[61873]_  = A266 & A265;
  assign \new_[61876]_  = ~A299 & ~A298;
  assign \new_[61877]_  = \new_[61876]_  & \new_[61873]_ ;
  assign \new_[61878]_  = \new_[61877]_  & \new_[61870]_ ;
  assign \new_[61882]_  = ~A167 & ~A169;
  assign \new_[61883]_  = A170 & \new_[61882]_ ;
  assign \new_[61887]_  = ~A201 & ~A200;
  assign \new_[61888]_  = A166 & \new_[61887]_ ;
  assign \new_[61889]_  = \new_[61888]_  & \new_[61883]_ ;
  assign \new_[61893]_  = ~A236 & ~A235;
  assign \new_[61894]_  = ~A233 & \new_[61893]_ ;
  assign \new_[61897]_  = ~A267 & ~A266;
  assign \new_[61900]_  = ~A300 & A298;
  assign \new_[61901]_  = \new_[61900]_  & \new_[61897]_ ;
  assign \new_[61902]_  = \new_[61901]_  & \new_[61894]_ ;
  assign \new_[61906]_  = ~A167 & ~A169;
  assign \new_[61907]_  = A170 & \new_[61906]_ ;
  assign \new_[61911]_  = ~A201 & ~A200;
  assign \new_[61912]_  = A166 & \new_[61911]_ ;
  assign \new_[61913]_  = \new_[61912]_  & \new_[61907]_ ;
  assign \new_[61917]_  = ~A236 & ~A235;
  assign \new_[61918]_  = ~A233 & \new_[61917]_ ;
  assign \new_[61921]_  = ~A267 & ~A266;
  assign \new_[61924]_  = A299 & A298;
  assign \new_[61925]_  = \new_[61924]_  & \new_[61921]_ ;
  assign \new_[61926]_  = \new_[61925]_  & \new_[61918]_ ;
  assign \new_[61930]_  = ~A167 & ~A169;
  assign \new_[61931]_  = A170 & \new_[61930]_ ;
  assign \new_[61935]_  = ~A201 & ~A200;
  assign \new_[61936]_  = A166 & \new_[61935]_ ;
  assign \new_[61937]_  = \new_[61936]_  & \new_[61931]_ ;
  assign \new_[61941]_  = ~A236 & ~A235;
  assign \new_[61942]_  = ~A233 & \new_[61941]_ ;
  assign \new_[61945]_  = ~A267 & ~A266;
  assign \new_[61948]_  = ~A299 & ~A298;
  assign \new_[61949]_  = \new_[61948]_  & \new_[61945]_ ;
  assign \new_[61950]_  = \new_[61949]_  & \new_[61942]_ ;
  assign \new_[61954]_  = ~A167 & ~A169;
  assign \new_[61955]_  = A170 & \new_[61954]_ ;
  assign \new_[61959]_  = ~A201 & ~A200;
  assign \new_[61960]_  = A166 & \new_[61959]_ ;
  assign \new_[61961]_  = \new_[61960]_  & \new_[61955]_ ;
  assign \new_[61965]_  = ~A236 & ~A235;
  assign \new_[61966]_  = ~A233 & \new_[61965]_ ;
  assign \new_[61969]_  = ~A266 & ~A265;
  assign \new_[61972]_  = ~A300 & A298;
  assign \new_[61973]_  = \new_[61972]_  & \new_[61969]_ ;
  assign \new_[61974]_  = \new_[61973]_  & \new_[61966]_ ;
  assign \new_[61978]_  = ~A167 & ~A169;
  assign \new_[61979]_  = A170 & \new_[61978]_ ;
  assign \new_[61983]_  = ~A201 & ~A200;
  assign \new_[61984]_  = A166 & \new_[61983]_ ;
  assign \new_[61985]_  = \new_[61984]_  & \new_[61979]_ ;
  assign \new_[61989]_  = ~A236 & ~A235;
  assign \new_[61990]_  = ~A233 & \new_[61989]_ ;
  assign \new_[61993]_  = ~A266 & ~A265;
  assign \new_[61996]_  = A299 & A298;
  assign \new_[61997]_  = \new_[61996]_  & \new_[61993]_ ;
  assign \new_[61998]_  = \new_[61997]_  & \new_[61990]_ ;
  assign \new_[62002]_  = ~A167 & ~A169;
  assign \new_[62003]_  = A170 & \new_[62002]_ ;
  assign \new_[62007]_  = ~A201 & ~A200;
  assign \new_[62008]_  = A166 & \new_[62007]_ ;
  assign \new_[62009]_  = \new_[62008]_  & \new_[62003]_ ;
  assign \new_[62013]_  = ~A236 & ~A235;
  assign \new_[62014]_  = ~A233 & \new_[62013]_ ;
  assign \new_[62017]_  = ~A266 & ~A265;
  assign \new_[62020]_  = ~A299 & ~A298;
  assign \new_[62021]_  = \new_[62020]_  & \new_[62017]_ ;
  assign \new_[62022]_  = \new_[62021]_  & \new_[62014]_ ;
  assign \new_[62026]_  = ~A167 & ~A169;
  assign \new_[62027]_  = A170 & \new_[62026]_ ;
  assign \new_[62031]_  = ~A201 & ~A200;
  assign \new_[62032]_  = A166 & \new_[62031]_ ;
  assign \new_[62033]_  = \new_[62032]_  & \new_[62027]_ ;
  assign \new_[62037]_  = A265 & ~A234;
  assign \new_[62038]_  = ~A233 & \new_[62037]_ ;
  assign \new_[62041]_  = A298 & A266;
  assign \new_[62044]_  = ~A302 & ~A301;
  assign \new_[62045]_  = \new_[62044]_  & \new_[62041]_ ;
  assign \new_[62046]_  = \new_[62045]_  & \new_[62038]_ ;
  assign \new_[62050]_  = ~A167 & ~A169;
  assign \new_[62051]_  = A170 & \new_[62050]_ ;
  assign \new_[62055]_  = ~A201 & ~A200;
  assign \new_[62056]_  = A166 & \new_[62055]_ ;
  assign \new_[62057]_  = \new_[62056]_  & \new_[62051]_ ;
  assign \new_[62061]_  = ~A266 & ~A234;
  assign \new_[62062]_  = ~A233 & \new_[62061]_ ;
  assign \new_[62065]_  = ~A269 & ~A268;
  assign \new_[62068]_  = ~A300 & A298;
  assign \new_[62069]_  = \new_[62068]_  & \new_[62065]_ ;
  assign \new_[62070]_  = \new_[62069]_  & \new_[62062]_ ;
  assign \new_[62074]_  = ~A167 & ~A169;
  assign \new_[62075]_  = A170 & \new_[62074]_ ;
  assign \new_[62079]_  = ~A201 & ~A200;
  assign \new_[62080]_  = A166 & \new_[62079]_ ;
  assign \new_[62081]_  = \new_[62080]_  & \new_[62075]_ ;
  assign \new_[62085]_  = ~A266 & ~A234;
  assign \new_[62086]_  = ~A233 & \new_[62085]_ ;
  assign \new_[62089]_  = ~A269 & ~A268;
  assign \new_[62092]_  = A299 & A298;
  assign \new_[62093]_  = \new_[62092]_  & \new_[62089]_ ;
  assign \new_[62094]_  = \new_[62093]_  & \new_[62086]_ ;
  assign \new_[62098]_  = ~A167 & ~A169;
  assign \new_[62099]_  = A170 & \new_[62098]_ ;
  assign \new_[62103]_  = ~A201 & ~A200;
  assign \new_[62104]_  = A166 & \new_[62103]_ ;
  assign \new_[62105]_  = \new_[62104]_  & \new_[62099]_ ;
  assign \new_[62109]_  = ~A266 & ~A234;
  assign \new_[62110]_  = ~A233 & \new_[62109]_ ;
  assign \new_[62113]_  = ~A269 & ~A268;
  assign \new_[62116]_  = ~A299 & ~A298;
  assign \new_[62117]_  = \new_[62116]_  & \new_[62113]_ ;
  assign \new_[62118]_  = \new_[62117]_  & \new_[62110]_ ;
  assign \new_[62122]_  = ~A167 & ~A169;
  assign \new_[62123]_  = A170 & \new_[62122]_ ;
  assign \new_[62127]_  = ~A201 & ~A200;
  assign \new_[62128]_  = A166 & \new_[62127]_ ;
  assign \new_[62129]_  = \new_[62128]_  & \new_[62123]_ ;
  assign \new_[62133]_  = ~A266 & ~A234;
  assign \new_[62134]_  = ~A233 & \new_[62133]_ ;
  assign \new_[62137]_  = A298 & ~A267;
  assign \new_[62140]_  = ~A302 & ~A301;
  assign \new_[62141]_  = \new_[62140]_  & \new_[62137]_ ;
  assign \new_[62142]_  = \new_[62141]_  & \new_[62134]_ ;
  assign \new_[62146]_  = ~A167 & ~A169;
  assign \new_[62147]_  = A170 & \new_[62146]_ ;
  assign \new_[62151]_  = ~A201 & ~A200;
  assign \new_[62152]_  = A166 & \new_[62151]_ ;
  assign \new_[62153]_  = \new_[62152]_  & \new_[62147]_ ;
  assign \new_[62157]_  = ~A265 & ~A234;
  assign \new_[62158]_  = ~A233 & \new_[62157]_ ;
  assign \new_[62161]_  = A298 & ~A266;
  assign \new_[62164]_  = ~A302 & ~A301;
  assign \new_[62165]_  = \new_[62164]_  & \new_[62161]_ ;
  assign \new_[62166]_  = \new_[62165]_  & \new_[62158]_ ;
  assign \new_[62170]_  = ~A167 & ~A169;
  assign \new_[62171]_  = A170 & \new_[62170]_ ;
  assign \new_[62175]_  = ~A201 & ~A200;
  assign \new_[62176]_  = A166 & \new_[62175]_ ;
  assign \new_[62177]_  = \new_[62176]_  & \new_[62171]_ ;
  assign \new_[62181]_  = A265 & ~A233;
  assign \new_[62182]_  = ~A232 & \new_[62181]_ ;
  assign \new_[62185]_  = A298 & A266;
  assign \new_[62188]_  = ~A302 & ~A301;
  assign \new_[62189]_  = \new_[62188]_  & \new_[62185]_ ;
  assign \new_[62190]_  = \new_[62189]_  & \new_[62182]_ ;
  assign \new_[62194]_  = ~A167 & ~A169;
  assign \new_[62195]_  = A170 & \new_[62194]_ ;
  assign \new_[62199]_  = ~A201 & ~A200;
  assign \new_[62200]_  = A166 & \new_[62199]_ ;
  assign \new_[62201]_  = \new_[62200]_  & \new_[62195]_ ;
  assign \new_[62205]_  = ~A266 & ~A233;
  assign \new_[62206]_  = ~A232 & \new_[62205]_ ;
  assign \new_[62209]_  = ~A269 & ~A268;
  assign \new_[62212]_  = ~A300 & A298;
  assign \new_[62213]_  = \new_[62212]_  & \new_[62209]_ ;
  assign \new_[62214]_  = \new_[62213]_  & \new_[62206]_ ;
  assign \new_[62218]_  = ~A167 & ~A169;
  assign \new_[62219]_  = A170 & \new_[62218]_ ;
  assign \new_[62223]_  = ~A201 & ~A200;
  assign \new_[62224]_  = A166 & \new_[62223]_ ;
  assign \new_[62225]_  = \new_[62224]_  & \new_[62219]_ ;
  assign \new_[62229]_  = ~A266 & ~A233;
  assign \new_[62230]_  = ~A232 & \new_[62229]_ ;
  assign \new_[62233]_  = ~A269 & ~A268;
  assign \new_[62236]_  = A299 & A298;
  assign \new_[62237]_  = \new_[62236]_  & \new_[62233]_ ;
  assign \new_[62238]_  = \new_[62237]_  & \new_[62230]_ ;
  assign \new_[62242]_  = ~A167 & ~A169;
  assign \new_[62243]_  = A170 & \new_[62242]_ ;
  assign \new_[62247]_  = ~A201 & ~A200;
  assign \new_[62248]_  = A166 & \new_[62247]_ ;
  assign \new_[62249]_  = \new_[62248]_  & \new_[62243]_ ;
  assign \new_[62253]_  = ~A266 & ~A233;
  assign \new_[62254]_  = ~A232 & \new_[62253]_ ;
  assign \new_[62257]_  = ~A269 & ~A268;
  assign \new_[62260]_  = ~A299 & ~A298;
  assign \new_[62261]_  = \new_[62260]_  & \new_[62257]_ ;
  assign \new_[62262]_  = \new_[62261]_  & \new_[62254]_ ;
  assign \new_[62266]_  = ~A167 & ~A169;
  assign \new_[62267]_  = A170 & \new_[62266]_ ;
  assign \new_[62271]_  = ~A201 & ~A200;
  assign \new_[62272]_  = A166 & \new_[62271]_ ;
  assign \new_[62273]_  = \new_[62272]_  & \new_[62267]_ ;
  assign \new_[62277]_  = ~A266 & ~A233;
  assign \new_[62278]_  = ~A232 & \new_[62277]_ ;
  assign \new_[62281]_  = A298 & ~A267;
  assign \new_[62284]_  = ~A302 & ~A301;
  assign \new_[62285]_  = \new_[62284]_  & \new_[62281]_ ;
  assign \new_[62286]_  = \new_[62285]_  & \new_[62278]_ ;
  assign \new_[62290]_  = ~A167 & ~A169;
  assign \new_[62291]_  = A170 & \new_[62290]_ ;
  assign \new_[62295]_  = ~A201 & ~A200;
  assign \new_[62296]_  = A166 & \new_[62295]_ ;
  assign \new_[62297]_  = \new_[62296]_  & \new_[62291]_ ;
  assign \new_[62301]_  = ~A265 & ~A233;
  assign \new_[62302]_  = ~A232 & \new_[62301]_ ;
  assign \new_[62305]_  = A298 & ~A266;
  assign \new_[62308]_  = ~A302 & ~A301;
  assign \new_[62309]_  = \new_[62308]_  & \new_[62305]_ ;
  assign \new_[62310]_  = \new_[62309]_  & \new_[62302]_ ;
  assign \new_[62314]_  = ~A167 & ~A169;
  assign \new_[62315]_  = A170 & \new_[62314]_ ;
  assign \new_[62319]_  = ~A200 & ~A199;
  assign \new_[62320]_  = A166 & \new_[62319]_ ;
  assign \new_[62321]_  = \new_[62320]_  & \new_[62315]_ ;
  assign \new_[62325]_  = A265 & A233;
  assign \new_[62326]_  = A232 & \new_[62325]_ ;
  assign \new_[62329]_  = ~A269 & ~A268;
  assign \new_[62332]_  = ~A300 & ~A299;
  assign \new_[62333]_  = \new_[62332]_  & \new_[62329]_ ;
  assign \new_[62334]_  = \new_[62333]_  & \new_[62326]_ ;
  assign \new_[62338]_  = ~A167 & ~A169;
  assign \new_[62339]_  = A170 & \new_[62338]_ ;
  assign \new_[62343]_  = ~A200 & ~A199;
  assign \new_[62344]_  = A166 & \new_[62343]_ ;
  assign \new_[62345]_  = \new_[62344]_  & \new_[62339]_ ;
  assign \new_[62349]_  = A265 & A233;
  assign \new_[62350]_  = A232 & \new_[62349]_ ;
  assign \new_[62353]_  = ~A269 & ~A268;
  assign \new_[62356]_  = A299 & A298;
  assign \new_[62357]_  = \new_[62356]_  & \new_[62353]_ ;
  assign \new_[62358]_  = \new_[62357]_  & \new_[62350]_ ;
  assign \new_[62362]_  = ~A167 & ~A169;
  assign \new_[62363]_  = A170 & \new_[62362]_ ;
  assign \new_[62367]_  = ~A200 & ~A199;
  assign \new_[62368]_  = A166 & \new_[62367]_ ;
  assign \new_[62369]_  = \new_[62368]_  & \new_[62363]_ ;
  assign \new_[62373]_  = A265 & A233;
  assign \new_[62374]_  = A232 & \new_[62373]_ ;
  assign \new_[62377]_  = ~A269 & ~A268;
  assign \new_[62380]_  = ~A299 & ~A298;
  assign \new_[62381]_  = \new_[62380]_  & \new_[62377]_ ;
  assign \new_[62382]_  = \new_[62381]_  & \new_[62374]_ ;
  assign \new_[62386]_  = ~A167 & ~A169;
  assign \new_[62387]_  = A170 & \new_[62386]_ ;
  assign \new_[62391]_  = ~A200 & ~A199;
  assign \new_[62392]_  = A166 & \new_[62391]_ ;
  assign \new_[62393]_  = \new_[62392]_  & \new_[62387]_ ;
  assign \new_[62397]_  = A265 & A233;
  assign \new_[62398]_  = A232 & \new_[62397]_ ;
  assign \new_[62401]_  = ~A299 & ~A267;
  assign \new_[62404]_  = ~A302 & ~A301;
  assign \new_[62405]_  = \new_[62404]_  & \new_[62401]_ ;
  assign \new_[62406]_  = \new_[62405]_  & \new_[62398]_ ;
  assign \new_[62410]_  = ~A167 & ~A169;
  assign \new_[62411]_  = A170 & \new_[62410]_ ;
  assign \new_[62415]_  = ~A200 & ~A199;
  assign \new_[62416]_  = A166 & \new_[62415]_ ;
  assign \new_[62417]_  = \new_[62416]_  & \new_[62411]_ ;
  assign \new_[62421]_  = A265 & A233;
  assign \new_[62422]_  = A232 & \new_[62421]_ ;
  assign \new_[62425]_  = ~A299 & A266;
  assign \new_[62428]_  = ~A302 & ~A301;
  assign \new_[62429]_  = \new_[62428]_  & \new_[62425]_ ;
  assign \new_[62430]_  = \new_[62429]_  & \new_[62422]_ ;
  assign \new_[62434]_  = ~A167 & ~A169;
  assign \new_[62435]_  = A170 & \new_[62434]_ ;
  assign \new_[62439]_  = ~A200 & ~A199;
  assign \new_[62440]_  = A166 & \new_[62439]_ ;
  assign \new_[62441]_  = \new_[62440]_  & \new_[62435]_ ;
  assign \new_[62445]_  = ~A265 & A233;
  assign \new_[62446]_  = A232 & \new_[62445]_ ;
  assign \new_[62449]_  = ~A299 & ~A266;
  assign \new_[62452]_  = ~A302 & ~A301;
  assign \new_[62453]_  = \new_[62452]_  & \new_[62449]_ ;
  assign \new_[62454]_  = \new_[62453]_  & \new_[62446]_ ;
  assign \new_[62458]_  = ~A167 & ~A169;
  assign \new_[62459]_  = A170 & \new_[62458]_ ;
  assign \new_[62463]_  = ~A200 & ~A199;
  assign \new_[62464]_  = A166 & \new_[62463]_ ;
  assign \new_[62465]_  = \new_[62464]_  & \new_[62459]_ ;
  assign \new_[62469]_  = ~A236 & ~A235;
  assign \new_[62470]_  = ~A233 & \new_[62469]_ ;
  assign \new_[62473]_  = A266 & A265;
  assign \new_[62476]_  = ~A300 & A298;
  assign \new_[62477]_  = \new_[62476]_  & \new_[62473]_ ;
  assign \new_[62478]_  = \new_[62477]_  & \new_[62470]_ ;
  assign \new_[62482]_  = ~A167 & ~A169;
  assign \new_[62483]_  = A170 & \new_[62482]_ ;
  assign \new_[62487]_  = ~A200 & ~A199;
  assign \new_[62488]_  = A166 & \new_[62487]_ ;
  assign \new_[62489]_  = \new_[62488]_  & \new_[62483]_ ;
  assign \new_[62493]_  = ~A236 & ~A235;
  assign \new_[62494]_  = ~A233 & \new_[62493]_ ;
  assign \new_[62497]_  = A266 & A265;
  assign \new_[62500]_  = A299 & A298;
  assign \new_[62501]_  = \new_[62500]_  & \new_[62497]_ ;
  assign \new_[62502]_  = \new_[62501]_  & \new_[62494]_ ;
  assign \new_[62506]_  = ~A167 & ~A169;
  assign \new_[62507]_  = A170 & \new_[62506]_ ;
  assign \new_[62511]_  = ~A200 & ~A199;
  assign \new_[62512]_  = A166 & \new_[62511]_ ;
  assign \new_[62513]_  = \new_[62512]_  & \new_[62507]_ ;
  assign \new_[62517]_  = ~A236 & ~A235;
  assign \new_[62518]_  = ~A233 & \new_[62517]_ ;
  assign \new_[62521]_  = A266 & A265;
  assign \new_[62524]_  = ~A299 & ~A298;
  assign \new_[62525]_  = \new_[62524]_  & \new_[62521]_ ;
  assign \new_[62526]_  = \new_[62525]_  & \new_[62518]_ ;
  assign \new_[62530]_  = ~A167 & ~A169;
  assign \new_[62531]_  = A170 & \new_[62530]_ ;
  assign \new_[62535]_  = ~A200 & ~A199;
  assign \new_[62536]_  = A166 & \new_[62535]_ ;
  assign \new_[62537]_  = \new_[62536]_  & \new_[62531]_ ;
  assign \new_[62541]_  = ~A236 & ~A235;
  assign \new_[62542]_  = ~A233 & \new_[62541]_ ;
  assign \new_[62545]_  = ~A267 & ~A266;
  assign \new_[62548]_  = ~A300 & A298;
  assign \new_[62549]_  = \new_[62548]_  & \new_[62545]_ ;
  assign \new_[62550]_  = \new_[62549]_  & \new_[62542]_ ;
  assign \new_[62554]_  = ~A167 & ~A169;
  assign \new_[62555]_  = A170 & \new_[62554]_ ;
  assign \new_[62559]_  = ~A200 & ~A199;
  assign \new_[62560]_  = A166 & \new_[62559]_ ;
  assign \new_[62561]_  = \new_[62560]_  & \new_[62555]_ ;
  assign \new_[62565]_  = ~A236 & ~A235;
  assign \new_[62566]_  = ~A233 & \new_[62565]_ ;
  assign \new_[62569]_  = ~A267 & ~A266;
  assign \new_[62572]_  = A299 & A298;
  assign \new_[62573]_  = \new_[62572]_  & \new_[62569]_ ;
  assign \new_[62574]_  = \new_[62573]_  & \new_[62566]_ ;
  assign \new_[62578]_  = ~A167 & ~A169;
  assign \new_[62579]_  = A170 & \new_[62578]_ ;
  assign \new_[62583]_  = ~A200 & ~A199;
  assign \new_[62584]_  = A166 & \new_[62583]_ ;
  assign \new_[62585]_  = \new_[62584]_  & \new_[62579]_ ;
  assign \new_[62589]_  = ~A236 & ~A235;
  assign \new_[62590]_  = ~A233 & \new_[62589]_ ;
  assign \new_[62593]_  = ~A267 & ~A266;
  assign \new_[62596]_  = ~A299 & ~A298;
  assign \new_[62597]_  = \new_[62596]_  & \new_[62593]_ ;
  assign \new_[62598]_  = \new_[62597]_  & \new_[62590]_ ;
  assign \new_[62602]_  = ~A167 & ~A169;
  assign \new_[62603]_  = A170 & \new_[62602]_ ;
  assign \new_[62607]_  = ~A200 & ~A199;
  assign \new_[62608]_  = A166 & \new_[62607]_ ;
  assign \new_[62609]_  = \new_[62608]_  & \new_[62603]_ ;
  assign \new_[62613]_  = ~A236 & ~A235;
  assign \new_[62614]_  = ~A233 & \new_[62613]_ ;
  assign \new_[62617]_  = ~A266 & ~A265;
  assign \new_[62620]_  = ~A300 & A298;
  assign \new_[62621]_  = \new_[62620]_  & \new_[62617]_ ;
  assign \new_[62622]_  = \new_[62621]_  & \new_[62614]_ ;
  assign \new_[62626]_  = ~A167 & ~A169;
  assign \new_[62627]_  = A170 & \new_[62626]_ ;
  assign \new_[62631]_  = ~A200 & ~A199;
  assign \new_[62632]_  = A166 & \new_[62631]_ ;
  assign \new_[62633]_  = \new_[62632]_  & \new_[62627]_ ;
  assign \new_[62637]_  = ~A236 & ~A235;
  assign \new_[62638]_  = ~A233 & \new_[62637]_ ;
  assign \new_[62641]_  = ~A266 & ~A265;
  assign \new_[62644]_  = A299 & A298;
  assign \new_[62645]_  = \new_[62644]_  & \new_[62641]_ ;
  assign \new_[62646]_  = \new_[62645]_  & \new_[62638]_ ;
  assign \new_[62650]_  = ~A167 & ~A169;
  assign \new_[62651]_  = A170 & \new_[62650]_ ;
  assign \new_[62655]_  = ~A200 & ~A199;
  assign \new_[62656]_  = A166 & \new_[62655]_ ;
  assign \new_[62657]_  = \new_[62656]_  & \new_[62651]_ ;
  assign \new_[62661]_  = ~A236 & ~A235;
  assign \new_[62662]_  = ~A233 & \new_[62661]_ ;
  assign \new_[62665]_  = ~A266 & ~A265;
  assign \new_[62668]_  = ~A299 & ~A298;
  assign \new_[62669]_  = \new_[62668]_  & \new_[62665]_ ;
  assign \new_[62670]_  = \new_[62669]_  & \new_[62662]_ ;
  assign \new_[62674]_  = ~A167 & ~A169;
  assign \new_[62675]_  = A170 & \new_[62674]_ ;
  assign \new_[62679]_  = ~A200 & ~A199;
  assign \new_[62680]_  = A166 & \new_[62679]_ ;
  assign \new_[62681]_  = \new_[62680]_  & \new_[62675]_ ;
  assign \new_[62685]_  = A265 & ~A234;
  assign \new_[62686]_  = ~A233 & \new_[62685]_ ;
  assign \new_[62689]_  = A298 & A266;
  assign \new_[62692]_  = ~A302 & ~A301;
  assign \new_[62693]_  = \new_[62692]_  & \new_[62689]_ ;
  assign \new_[62694]_  = \new_[62693]_  & \new_[62686]_ ;
  assign \new_[62698]_  = ~A167 & ~A169;
  assign \new_[62699]_  = A170 & \new_[62698]_ ;
  assign \new_[62703]_  = ~A200 & ~A199;
  assign \new_[62704]_  = A166 & \new_[62703]_ ;
  assign \new_[62705]_  = \new_[62704]_  & \new_[62699]_ ;
  assign \new_[62709]_  = ~A266 & ~A234;
  assign \new_[62710]_  = ~A233 & \new_[62709]_ ;
  assign \new_[62713]_  = ~A269 & ~A268;
  assign \new_[62716]_  = ~A300 & A298;
  assign \new_[62717]_  = \new_[62716]_  & \new_[62713]_ ;
  assign \new_[62718]_  = \new_[62717]_  & \new_[62710]_ ;
  assign \new_[62722]_  = ~A167 & ~A169;
  assign \new_[62723]_  = A170 & \new_[62722]_ ;
  assign \new_[62727]_  = ~A200 & ~A199;
  assign \new_[62728]_  = A166 & \new_[62727]_ ;
  assign \new_[62729]_  = \new_[62728]_  & \new_[62723]_ ;
  assign \new_[62733]_  = ~A266 & ~A234;
  assign \new_[62734]_  = ~A233 & \new_[62733]_ ;
  assign \new_[62737]_  = ~A269 & ~A268;
  assign \new_[62740]_  = A299 & A298;
  assign \new_[62741]_  = \new_[62740]_  & \new_[62737]_ ;
  assign \new_[62742]_  = \new_[62741]_  & \new_[62734]_ ;
  assign \new_[62746]_  = ~A167 & ~A169;
  assign \new_[62747]_  = A170 & \new_[62746]_ ;
  assign \new_[62751]_  = ~A200 & ~A199;
  assign \new_[62752]_  = A166 & \new_[62751]_ ;
  assign \new_[62753]_  = \new_[62752]_  & \new_[62747]_ ;
  assign \new_[62757]_  = ~A266 & ~A234;
  assign \new_[62758]_  = ~A233 & \new_[62757]_ ;
  assign \new_[62761]_  = ~A269 & ~A268;
  assign \new_[62764]_  = ~A299 & ~A298;
  assign \new_[62765]_  = \new_[62764]_  & \new_[62761]_ ;
  assign \new_[62766]_  = \new_[62765]_  & \new_[62758]_ ;
  assign \new_[62770]_  = ~A167 & ~A169;
  assign \new_[62771]_  = A170 & \new_[62770]_ ;
  assign \new_[62775]_  = ~A200 & ~A199;
  assign \new_[62776]_  = A166 & \new_[62775]_ ;
  assign \new_[62777]_  = \new_[62776]_  & \new_[62771]_ ;
  assign \new_[62781]_  = ~A266 & ~A234;
  assign \new_[62782]_  = ~A233 & \new_[62781]_ ;
  assign \new_[62785]_  = A298 & ~A267;
  assign \new_[62788]_  = ~A302 & ~A301;
  assign \new_[62789]_  = \new_[62788]_  & \new_[62785]_ ;
  assign \new_[62790]_  = \new_[62789]_  & \new_[62782]_ ;
  assign \new_[62794]_  = ~A167 & ~A169;
  assign \new_[62795]_  = A170 & \new_[62794]_ ;
  assign \new_[62799]_  = ~A200 & ~A199;
  assign \new_[62800]_  = A166 & \new_[62799]_ ;
  assign \new_[62801]_  = \new_[62800]_  & \new_[62795]_ ;
  assign \new_[62805]_  = ~A265 & ~A234;
  assign \new_[62806]_  = ~A233 & \new_[62805]_ ;
  assign \new_[62809]_  = A298 & ~A266;
  assign \new_[62812]_  = ~A302 & ~A301;
  assign \new_[62813]_  = \new_[62812]_  & \new_[62809]_ ;
  assign \new_[62814]_  = \new_[62813]_  & \new_[62806]_ ;
  assign \new_[62818]_  = ~A167 & ~A169;
  assign \new_[62819]_  = A170 & \new_[62818]_ ;
  assign \new_[62823]_  = ~A200 & ~A199;
  assign \new_[62824]_  = A166 & \new_[62823]_ ;
  assign \new_[62825]_  = \new_[62824]_  & \new_[62819]_ ;
  assign \new_[62829]_  = A265 & ~A233;
  assign \new_[62830]_  = ~A232 & \new_[62829]_ ;
  assign \new_[62833]_  = A298 & A266;
  assign \new_[62836]_  = ~A302 & ~A301;
  assign \new_[62837]_  = \new_[62836]_  & \new_[62833]_ ;
  assign \new_[62838]_  = \new_[62837]_  & \new_[62830]_ ;
  assign \new_[62842]_  = ~A167 & ~A169;
  assign \new_[62843]_  = A170 & \new_[62842]_ ;
  assign \new_[62847]_  = ~A200 & ~A199;
  assign \new_[62848]_  = A166 & \new_[62847]_ ;
  assign \new_[62849]_  = \new_[62848]_  & \new_[62843]_ ;
  assign \new_[62853]_  = ~A266 & ~A233;
  assign \new_[62854]_  = ~A232 & \new_[62853]_ ;
  assign \new_[62857]_  = ~A269 & ~A268;
  assign \new_[62860]_  = ~A300 & A298;
  assign \new_[62861]_  = \new_[62860]_  & \new_[62857]_ ;
  assign \new_[62862]_  = \new_[62861]_  & \new_[62854]_ ;
  assign \new_[62866]_  = ~A167 & ~A169;
  assign \new_[62867]_  = A170 & \new_[62866]_ ;
  assign \new_[62871]_  = ~A200 & ~A199;
  assign \new_[62872]_  = A166 & \new_[62871]_ ;
  assign \new_[62873]_  = \new_[62872]_  & \new_[62867]_ ;
  assign \new_[62877]_  = ~A266 & ~A233;
  assign \new_[62878]_  = ~A232 & \new_[62877]_ ;
  assign \new_[62881]_  = ~A269 & ~A268;
  assign \new_[62884]_  = A299 & A298;
  assign \new_[62885]_  = \new_[62884]_  & \new_[62881]_ ;
  assign \new_[62886]_  = \new_[62885]_  & \new_[62878]_ ;
  assign \new_[62890]_  = ~A167 & ~A169;
  assign \new_[62891]_  = A170 & \new_[62890]_ ;
  assign \new_[62895]_  = ~A200 & ~A199;
  assign \new_[62896]_  = A166 & \new_[62895]_ ;
  assign \new_[62897]_  = \new_[62896]_  & \new_[62891]_ ;
  assign \new_[62901]_  = ~A266 & ~A233;
  assign \new_[62902]_  = ~A232 & \new_[62901]_ ;
  assign \new_[62905]_  = ~A269 & ~A268;
  assign \new_[62908]_  = ~A299 & ~A298;
  assign \new_[62909]_  = \new_[62908]_  & \new_[62905]_ ;
  assign \new_[62910]_  = \new_[62909]_  & \new_[62902]_ ;
  assign \new_[62914]_  = ~A167 & ~A169;
  assign \new_[62915]_  = A170 & \new_[62914]_ ;
  assign \new_[62919]_  = ~A200 & ~A199;
  assign \new_[62920]_  = A166 & \new_[62919]_ ;
  assign \new_[62921]_  = \new_[62920]_  & \new_[62915]_ ;
  assign \new_[62925]_  = ~A266 & ~A233;
  assign \new_[62926]_  = ~A232 & \new_[62925]_ ;
  assign \new_[62929]_  = A298 & ~A267;
  assign \new_[62932]_  = ~A302 & ~A301;
  assign \new_[62933]_  = \new_[62932]_  & \new_[62929]_ ;
  assign \new_[62934]_  = \new_[62933]_  & \new_[62926]_ ;
  assign \new_[62938]_  = ~A167 & ~A169;
  assign \new_[62939]_  = A170 & \new_[62938]_ ;
  assign \new_[62943]_  = ~A200 & ~A199;
  assign \new_[62944]_  = A166 & \new_[62943]_ ;
  assign \new_[62945]_  = \new_[62944]_  & \new_[62939]_ ;
  assign \new_[62949]_  = ~A265 & ~A233;
  assign \new_[62950]_  = ~A232 & \new_[62949]_ ;
  assign \new_[62953]_  = A298 & ~A266;
  assign \new_[62956]_  = ~A302 & ~A301;
  assign \new_[62957]_  = \new_[62956]_  & \new_[62953]_ ;
  assign \new_[62958]_  = \new_[62957]_  & \new_[62950]_ ;
  assign \new_[62962]_  = ~A168 & ~A169;
  assign \new_[62963]_  = ~A170 & \new_[62962]_ ;
  assign \new_[62967]_  = A201 & ~A200;
  assign \new_[62968]_  = A199 & \new_[62967]_ ;
  assign \new_[62969]_  = \new_[62968]_  & \new_[62963]_ ;
  assign \new_[62973]_  = A233 & A232;
  assign \new_[62974]_  = A202 & \new_[62973]_ ;
  assign \new_[62977]_  = ~A267 & A265;
  assign \new_[62980]_  = ~A300 & ~A299;
  assign \new_[62981]_  = \new_[62980]_  & \new_[62977]_ ;
  assign \new_[62982]_  = \new_[62981]_  & \new_[62974]_ ;
  assign \new_[62986]_  = ~A168 & ~A169;
  assign \new_[62987]_  = ~A170 & \new_[62986]_ ;
  assign \new_[62991]_  = A201 & ~A200;
  assign \new_[62992]_  = A199 & \new_[62991]_ ;
  assign \new_[62993]_  = \new_[62992]_  & \new_[62987]_ ;
  assign \new_[62997]_  = A233 & A232;
  assign \new_[62998]_  = A202 & \new_[62997]_ ;
  assign \new_[63001]_  = ~A267 & A265;
  assign \new_[63004]_  = A299 & A298;
  assign \new_[63005]_  = \new_[63004]_  & \new_[63001]_ ;
  assign \new_[63006]_  = \new_[63005]_  & \new_[62998]_ ;
  assign \new_[63010]_  = ~A168 & ~A169;
  assign \new_[63011]_  = ~A170 & \new_[63010]_ ;
  assign \new_[63015]_  = A201 & ~A200;
  assign \new_[63016]_  = A199 & \new_[63015]_ ;
  assign \new_[63017]_  = \new_[63016]_  & \new_[63011]_ ;
  assign \new_[63021]_  = A233 & A232;
  assign \new_[63022]_  = A202 & \new_[63021]_ ;
  assign \new_[63025]_  = ~A267 & A265;
  assign \new_[63028]_  = ~A299 & ~A298;
  assign \new_[63029]_  = \new_[63028]_  & \new_[63025]_ ;
  assign \new_[63030]_  = \new_[63029]_  & \new_[63022]_ ;
  assign \new_[63034]_  = ~A168 & ~A169;
  assign \new_[63035]_  = ~A170 & \new_[63034]_ ;
  assign \new_[63039]_  = A201 & ~A200;
  assign \new_[63040]_  = A199 & \new_[63039]_ ;
  assign \new_[63041]_  = \new_[63040]_  & \new_[63035]_ ;
  assign \new_[63045]_  = A233 & A232;
  assign \new_[63046]_  = A202 & \new_[63045]_ ;
  assign \new_[63049]_  = A266 & A265;
  assign \new_[63052]_  = ~A300 & ~A299;
  assign \new_[63053]_  = \new_[63052]_  & \new_[63049]_ ;
  assign \new_[63054]_  = \new_[63053]_  & \new_[63046]_ ;
  assign \new_[63058]_  = ~A168 & ~A169;
  assign \new_[63059]_  = ~A170 & \new_[63058]_ ;
  assign \new_[63063]_  = A201 & ~A200;
  assign \new_[63064]_  = A199 & \new_[63063]_ ;
  assign \new_[63065]_  = \new_[63064]_  & \new_[63059]_ ;
  assign \new_[63069]_  = A233 & A232;
  assign \new_[63070]_  = A202 & \new_[63069]_ ;
  assign \new_[63073]_  = A266 & A265;
  assign \new_[63076]_  = A299 & A298;
  assign \new_[63077]_  = \new_[63076]_  & \new_[63073]_ ;
  assign \new_[63078]_  = \new_[63077]_  & \new_[63070]_ ;
  assign \new_[63082]_  = ~A168 & ~A169;
  assign \new_[63083]_  = ~A170 & \new_[63082]_ ;
  assign \new_[63087]_  = A201 & ~A200;
  assign \new_[63088]_  = A199 & \new_[63087]_ ;
  assign \new_[63089]_  = \new_[63088]_  & \new_[63083]_ ;
  assign \new_[63093]_  = A233 & A232;
  assign \new_[63094]_  = A202 & \new_[63093]_ ;
  assign \new_[63097]_  = A266 & A265;
  assign \new_[63100]_  = ~A299 & ~A298;
  assign \new_[63101]_  = \new_[63100]_  & \new_[63097]_ ;
  assign \new_[63102]_  = \new_[63101]_  & \new_[63094]_ ;
  assign \new_[63106]_  = ~A168 & ~A169;
  assign \new_[63107]_  = ~A170 & \new_[63106]_ ;
  assign \new_[63111]_  = A201 & ~A200;
  assign \new_[63112]_  = A199 & \new_[63111]_ ;
  assign \new_[63113]_  = \new_[63112]_  & \new_[63107]_ ;
  assign \new_[63117]_  = A233 & A232;
  assign \new_[63118]_  = A202 & \new_[63117]_ ;
  assign \new_[63121]_  = ~A266 & ~A265;
  assign \new_[63124]_  = ~A300 & ~A299;
  assign \new_[63125]_  = \new_[63124]_  & \new_[63121]_ ;
  assign \new_[63126]_  = \new_[63125]_  & \new_[63118]_ ;
  assign \new_[63130]_  = ~A168 & ~A169;
  assign \new_[63131]_  = ~A170 & \new_[63130]_ ;
  assign \new_[63135]_  = A201 & ~A200;
  assign \new_[63136]_  = A199 & \new_[63135]_ ;
  assign \new_[63137]_  = \new_[63136]_  & \new_[63131]_ ;
  assign \new_[63141]_  = A233 & A232;
  assign \new_[63142]_  = A202 & \new_[63141]_ ;
  assign \new_[63145]_  = ~A266 & ~A265;
  assign \new_[63148]_  = A299 & A298;
  assign \new_[63149]_  = \new_[63148]_  & \new_[63145]_ ;
  assign \new_[63150]_  = \new_[63149]_  & \new_[63142]_ ;
  assign \new_[63154]_  = ~A168 & ~A169;
  assign \new_[63155]_  = ~A170 & \new_[63154]_ ;
  assign \new_[63159]_  = A201 & ~A200;
  assign \new_[63160]_  = A199 & \new_[63159]_ ;
  assign \new_[63161]_  = \new_[63160]_  & \new_[63155]_ ;
  assign \new_[63165]_  = A233 & A232;
  assign \new_[63166]_  = A202 & \new_[63165]_ ;
  assign \new_[63169]_  = ~A266 & ~A265;
  assign \new_[63172]_  = ~A299 & ~A298;
  assign \new_[63173]_  = \new_[63172]_  & \new_[63169]_ ;
  assign \new_[63174]_  = \new_[63173]_  & \new_[63166]_ ;
  assign \new_[63178]_  = ~A168 & ~A169;
  assign \new_[63179]_  = ~A170 & \new_[63178]_ ;
  assign \new_[63183]_  = A201 & ~A200;
  assign \new_[63184]_  = A199 & \new_[63183]_ ;
  assign \new_[63185]_  = \new_[63184]_  & \new_[63179]_ ;
  assign \new_[63189]_  = A233 & ~A232;
  assign \new_[63190]_  = A202 & \new_[63189]_ ;
  assign \new_[63193]_  = ~A299 & A298;
  assign \new_[63196]_  = A301 & A300;
  assign \new_[63197]_  = \new_[63196]_  & \new_[63193]_ ;
  assign \new_[63198]_  = \new_[63197]_  & \new_[63190]_ ;
  assign \new_[63202]_  = ~A168 & ~A169;
  assign \new_[63203]_  = ~A170 & \new_[63202]_ ;
  assign \new_[63207]_  = A201 & ~A200;
  assign \new_[63208]_  = A199 & \new_[63207]_ ;
  assign \new_[63209]_  = \new_[63208]_  & \new_[63203]_ ;
  assign \new_[63213]_  = A233 & ~A232;
  assign \new_[63214]_  = A202 & \new_[63213]_ ;
  assign \new_[63217]_  = ~A299 & A298;
  assign \new_[63220]_  = A302 & A300;
  assign \new_[63221]_  = \new_[63220]_  & \new_[63217]_ ;
  assign \new_[63222]_  = \new_[63221]_  & \new_[63214]_ ;
  assign \new_[63226]_  = ~A168 & ~A169;
  assign \new_[63227]_  = ~A170 & \new_[63226]_ ;
  assign \new_[63231]_  = A201 & ~A200;
  assign \new_[63232]_  = A199 & \new_[63231]_ ;
  assign \new_[63233]_  = \new_[63232]_  & \new_[63227]_ ;
  assign \new_[63237]_  = A233 & ~A232;
  assign \new_[63238]_  = A202 & \new_[63237]_ ;
  assign \new_[63241]_  = ~A266 & A265;
  assign \new_[63244]_  = A268 & A267;
  assign \new_[63245]_  = \new_[63244]_  & \new_[63241]_ ;
  assign \new_[63246]_  = \new_[63245]_  & \new_[63238]_ ;
  assign \new_[63250]_  = ~A168 & ~A169;
  assign \new_[63251]_  = ~A170 & \new_[63250]_ ;
  assign \new_[63255]_  = A201 & ~A200;
  assign \new_[63256]_  = A199 & \new_[63255]_ ;
  assign \new_[63257]_  = \new_[63256]_  & \new_[63251]_ ;
  assign \new_[63261]_  = A233 & ~A232;
  assign \new_[63262]_  = A202 & \new_[63261]_ ;
  assign \new_[63265]_  = ~A266 & A265;
  assign \new_[63268]_  = A269 & A267;
  assign \new_[63269]_  = \new_[63268]_  & \new_[63265]_ ;
  assign \new_[63270]_  = \new_[63269]_  & \new_[63262]_ ;
  assign \new_[63274]_  = ~A168 & ~A169;
  assign \new_[63275]_  = ~A170 & \new_[63274]_ ;
  assign \new_[63279]_  = A201 & ~A200;
  assign \new_[63280]_  = A199 & \new_[63279]_ ;
  assign \new_[63281]_  = \new_[63280]_  & \new_[63275]_ ;
  assign \new_[63285]_  = ~A234 & ~A233;
  assign \new_[63286]_  = A202 & \new_[63285]_ ;
  assign \new_[63289]_  = A266 & A265;
  assign \new_[63292]_  = ~A300 & A298;
  assign \new_[63293]_  = \new_[63292]_  & \new_[63289]_ ;
  assign \new_[63294]_  = \new_[63293]_  & \new_[63286]_ ;
  assign \new_[63298]_  = ~A168 & ~A169;
  assign \new_[63299]_  = ~A170 & \new_[63298]_ ;
  assign \new_[63303]_  = A201 & ~A200;
  assign \new_[63304]_  = A199 & \new_[63303]_ ;
  assign \new_[63305]_  = \new_[63304]_  & \new_[63299]_ ;
  assign \new_[63309]_  = ~A234 & ~A233;
  assign \new_[63310]_  = A202 & \new_[63309]_ ;
  assign \new_[63313]_  = A266 & A265;
  assign \new_[63316]_  = A299 & A298;
  assign \new_[63317]_  = \new_[63316]_  & \new_[63313]_ ;
  assign \new_[63318]_  = \new_[63317]_  & \new_[63310]_ ;
  assign \new_[63322]_  = ~A168 & ~A169;
  assign \new_[63323]_  = ~A170 & \new_[63322]_ ;
  assign \new_[63327]_  = A201 & ~A200;
  assign \new_[63328]_  = A199 & \new_[63327]_ ;
  assign \new_[63329]_  = \new_[63328]_  & \new_[63323]_ ;
  assign \new_[63333]_  = ~A234 & ~A233;
  assign \new_[63334]_  = A202 & \new_[63333]_ ;
  assign \new_[63337]_  = A266 & A265;
  assign \new_[63340]_  = ~A299 & ~A298;
  assign \new_[63341]_  = \new_[63340]_  & \new_[63337]_ ;
  assign \new_[63342]_  = \new_[63341]_  & \new_[63334]_ ;
  assign \new_[63346]_  = ~A168 & ~A169;
  assign \new_[63347]_  = ~A170 & \new_[63346]_ ;
  assign \new_[63351]_  = A201 & ~A200;
  assign \new_[63352]_  = A199 & \new_[63351]_ ;
  assign \new_[63353]_  = \new_[63352]_  & \new_[63347]_ ;
  assign \new_[63357]_  = ~A234 & ~A233;
  assign \new_[63358]_  = A202 & \new_[63357]_ ;
  assign \new_[63361]_  = ~A267 & ~A266;
  assign \new_[63364]_  = ~A300 & A298;
  assign \new_[63365]_  = \new_[63364]_  & \new_[63361]_ ;
  assign \new_[63366]_  = \new_[63365]_  & \new_[63358]_ ;
  assign \new_[63370]_  = ~A168 & ~A169;
  assign \new_[63371]_  = ~A170 & \new_[63370]_ ;
  assign \new_[63375]_  = A201 & ~A200;
  assign \new_[63376]_  = A199 & \new_[63375]_ ;
  assign \new_[63377]_  = \new_[63376]_  & \new_[63371]_ ;
  assign \new_[63381]_  = ~A234 & ~A233;
  assign \new_[63382]_  = A202 & \new_[63381]_ ;
  assign \new_[63385]_  = ~A267 & ~A266;
  assign \new_[63388]_  = A299 & A298;
  assign \new_[63389]_  = \new_[63388]_  & \new_[63385]_ ;
  assign \new_[63390]_  = \new_[63389]_  & \new_[63382]_ ;
  assign \new_[63394]_  = ~A168 & ~A169;
  assign \new_[63395]_  = ~A170 & \new_[63394]_ ;
  assign \new_[63399]_  = A201 & ~A200;
  assign \new_[63400]_  = A199 & \new_[63399]_ ;
  assign \new_[63401]_  = \new_[63400]_  & \new_[63395]_ ;
  assign \new_[63405]_  = ~A234 & ~A233;
  assign \new_[63406]_  = A202 & \new_[63405]_ ;
  assign \new_[63409]_  = ~A267 & ~A266;
  assign \new_[63412]_  = ~A299 & ~A298;
  assign \new_[63413]_  = \new_[63412]_  & \new_[63409]_ ;
  assign \new_[63414]_  = \new_[63413]_  & \new_[63406]_ ;
  assign \new_[63418]_  = ~A168 & ~A169;
  assign \new_[63419]_  = ~A170 & \new_[63418]_ ;
  assign \new_[63423]_  = A201 & ~A200;
  assign \new_[63424]_  = A199 & \new_[63423]_ ;
  assign \new_[63425]_  = \new_[63424]_  & \new_[63419]_ ;
  assign \new_[63429]_  = ~A234 & ~A233;
  assign \new_[63430]_  = A202 & \new_[63429]_ ;
  assign \new_[63433]_  = ~A266 & ~A265;
  assign \new_[63436]_  = ~A300 & A298;
  assign \new_[63437]_  = \new_[63436]_  & \new_[63433]_ ;
  assign \new_[63438]_  = \new_[63437]_  & \new_[63430]_ ;
  assign \new_[63442]_  = ~A168 & ~A169;
  assign \new_[63443]_  = ~A170 & \new_[63442]_ ;
  assign \new_[63447]_  = A201 & ~A200;
  assign \new_[63448]_  = A199 & \new_[63447]_ ;
  assign \new_[63449]_  = \new_[63448]_  & \new_[63443]_ ;
  assign \new_[63453]_  = ~A234 & ~A233;
  assign \new_[63454]_  = A202 & \new_[63453]_ ;
  assign \new_[63457]_  = ~A266 & ~A265;
  assign \new_[63460]_  = A299 & A298;
  assign \new_[63461]_  = \new_[63460]_  & \new_[63457]_ ;
  assign \new_[63462]_  = \new_[63461]_  & \new_[63454]_ ;
  assign \new_[63466]_  = ~A168 & ~A169;
  assign \new_[63467]_  = ~A170 & \new_[63466]_ ;
  assign \new_[63471]_  = A201 & ~A200;
  assign \new_[63472]_  = A199 & \new_[63471]_ ;
  assign \new_[63473]_  = \new_[63472]_  & \new_[63467]_ ;
  assign \new_[63477]_  = ~A234 & ~A233;
  assign \new_[63478]_  = A202 & \new_[63477]_ ;
  assign \new_[63481]_  = ~A266 & ~A265;
  assign \new_[63484]_  = ~A299 & ~A298;
  assign \new_[63485]_  = \new_[63484]_  & \new_[63481]_ ;
  assign \new_[63486]_  = \new_[63485]_  & \new_[63478]_ ;
  assign \new_[63490]_  = ~A168 & ~A169;
  assign \new_[63491]_  = ~A170 & \new_[63490]_ ;
  assign \new_[63495]_  = A201 & ~A200;
  assign \new_[63496]_  = A199 & \new_[63495]_ ;
  assign \new_[63497]_  = \new_[63496]_  & \new_[63491]_ ;
  assign \new_[63501]_  = ~A233 & A232;
  assign \new_[63502]_  = A202 & \new_[63501]_ ;
  assign \new_[63505]_  = A235 & A234;
  assign \new_[63508]_  = A299 & ~A298;
  assign \new_[63509]_  = \new_[63508]_  & \new_[63505]_ ;
  assign \new_[63510]_  = \new_[63509]_  & \new_[63502]_ ;
  assign \new_[63514]_  = ~A168 & ~A169;
  assign \new_[63515]_  = ~A170 & \new_[63514]_ ;
  assign \new_[63519]_  = A201 & ~A200;
  assign \new_[63520]_  = A199 & \new_[63519]_ ;
  assign \new_[63521]_  = \new_[63520]_  & \new_[63515]_ ;
  assign \new_[63525]_  = ~A233 & A232;
  assign \new_[63526]_  = A202 & \new_[63525]_ ;
  assign \new_[63529]_  = A235 & A234;
  assign \new_[63532]_  = A266 & ~A265;
  assign \new_[63533]_  = \new_[63532]_  & \new_[63529]_ ;
  assign \new_[63534]_  = \new_[63533]_  & \new_[63526]_ ;
  assign \new_[63538]_  = ~A168 & ~A169;
  assign \new_[63539]_  = ~A170 & \new_[63538]_ ;
  assign \new_[63543]_  = A201 & ~A200;
  assign \new_[63544]_  = A199 & \new_[63543]_ ;
  assign \new_[63545]_  = \new_[63544]_  & \new_[63539]_ ;
  assign \new_[63549]_  = ~A233 & A232;
  assign \new_[63550]_  = A202 & \new_[63549]_ ;
  assign \new_[63553]_  = A236 & A234;
  assign \new_[63556]_  = A299 & ~A298;
  assign \new_[63557]_  = \new_[63556]_  & \new_[63553]_ ;
  assign \new_[63558]_  = \new_[63557]_  & \new_[63550]_ ;
  assign \new_[63562]_  = ~A168 & ~A169;
  assign \new_[63563]_  = ~A170 & \new_[63562]_ ;
  assign \new_[63567]_  = A201 & ~A200;
  assign \new_[63568]_  = A199 & \new_[63567]_ ;
  assign \new_[63569]_  = \new_[63568]_  & \new_[63563]_ ;
  assign \new_[63573]_  = ~A233 & A232;
  assign \new_[63574]_  = A202 & \new_[63573]_ ;
  assign \new_[63577]_  = A236 & A234;
  assign \new_[63580]_  = A266 & ~A265;
  assign \new_[63581]_  = \new_[63580]_  & \new_[63577]_ ;
  assign \new_[63582]_  = \new_[63581]_  & \new_[63574]_ ;
  assign \new_[63586]_  = ~A168 & ~A169;
  assign \new_[63587]_  = ~A170 & \new_[63586]_ ;
  assign \new_[63591]_  = A201 & ~A200;
  assign \new_[63592]_  = A199 & \new_[63591]_ ;
  assign \new_[63593]_  = \new_[63592]_  & \new_[63587]_ ;
  assign \new_[63597]_  = ~A233 & ~A232;
  assign \new_[63598]_  = A202 & \new_[63597]_ ;
  assign \new_[63601]_  = A266 & A265;
  assign \new_[63604]_  = ~A300 & A298;
  assign \new_[63605]_  = \new_[63604]_  & \new_[63601]_ ;
  assign \new_[63606]_  = \new_[63605]_  & \new_[63598]_ ;
  assign \new_[63610]_  = ~A168 & ~A169;
  assign \new_[63611]_  = ~A170 & \new_[63610]_ ;
  assign \new_[63615]_  = A201 & ~A200;
  assign \new_[63616]_  = A199 & \new_[63615]_ ;
  assign \new_[63617]_  = \new_[63616]_  & \new_[63611]_ ;
  assign \new_[63621]_  = ~A233 & ~A232;
  assign \new_[63622]_  = A202 & \new_[63621]_ ;
  assign \new_[63625]_  = A266 & A265;
  assign \new_[63628]_  = A299 & A298;
  assign \new_[63629]_  = \new_[63628]_  & \new_[63625]_ ;
  assign \new_[63630]_  = \new_[63629]_  & \new_[63622]_ ;
  assign \new_[63634]_  = ~A168 & ~A169;
  assign \new_[63635]_  = ~A170 & \new_[63634]_ ;
  assign \new_[63639]_  = A201 & ~A200;
  assign \new_[63640]_  = A199 & \new_[63639]_ ;
  assign \new_[63641]_  = \new_[63640]_  & \new_[63635]_ ;
  assign \new_[63645]_  = ~A233 & ~A232;
  assign \new_[63646]_  = A202 & \new_[63645]_ ;
  assign \new_[63649]_  = A266 & A265;
  assign \new_[63652]_  = ~A299 & ~A298;
  assign \new_[63653]_  = \new_[63652]_  & \new_[63649]_ ;
  assign \new_[63654]_  = \new_[63653]_  & \new_[63646]_ ;
  assign \new_[63658]_  = ~A168 & ~A169;
  assign \new_[63659]_  = ~A170 & \new_[63658]_ ;
  assign \new_[63663]_  = A201 & ~A200;
  assign \new_[63664]_  = A199 & \new_[63663]_ ;
  assign \new_[63665]_  = \new_[63664]_  & \new_[63659]_ ;
  assign \new_[63669]_  = ~A233 & ~A232;
  assign \new_[63670]_  = A202 & \new_[63669]_ ;
  assign \new_[63673]_  = ~A267 & ~A266;
  assign \new_[63676]_  = ~A300 & A298;
  assign \new_[63677]_  = \new_[63676]_  & \new_[63673]_ ;
  assign \new_[63678]_  = \new_[63677]_  & \new_[63670]_ ;
  assign \new_[63682]_  = ~A168 & ~A169;
  assign \new_[63683]_  = ~A170 & \new_[63682]_ ;
  assign \new_[63687]_  = A201 & ~A200;
  assign \new_[63688]_  = A199 & \new_[63687]_ ;
  assign \new_[63689]_  = \new_[63688]_  & \new_[63683]_ ;
  assign \new_[63693]_  = ~A233 & ~A232;
  assign \new_[63694]_  = A202 & \new_[63693]_ ;
  assign \new_[63697]_  = ~A267 & ~A266;
  assign \new_[63700]_  = A299 & A298;
  assign \new_[63701]_  = \new_[63700]_  & \new_[63697]_ ;
  assign \new_[63702]_  = \new_[63701]_  & \new_[63694]_ ;
  assign \new_[63706]_  = ~A168 & ~A169;
  assign \new_[63707]_  = ~A170 & \new_[63706]_ ;
  assign \new_[63711]_  = A201 & ~A200;
  assign \new_[63712]_  = A199 & \new_[63711]_ ;
  assign \new_[63713]_  = \new_[63712]_  & \new_[63707]_ ;
  assign \new_[63717]_  = ~A233 & ~A232;
  assign \new_[63718]_  = A202 & \new_[63717]_ ;
  assign \new_[63721]_  = ~A267 & ~A266;
  assign \new_[63724]_  = ~A299 & ~A298;
  assign \new_[63725]_  = \new_[63724]_  & \new_[63721]_ ;
  assign \new_[63726]_  = \new_[63725]_  & \new_[63718]_ ;
  assign \new_[63730]_  = ~A168 & ~A169;
  assign \new_[63731]_  = ~A170 & \new_[63730]_ ;
  assign \new_[63735]_  = A201 & ~A200;
  assign \new_[63736]_  = A199 & \new_[63735]_ ;
  assign \new_[63737]_  = \new_[63736]_  & \new_[63731]_ ;
  assign \new_[63741]_  = ~A233 & ~A232;
  assign \new_[63742]_  = A202 & \new_[63741]_ ;
  assign \new_[63745]_  = ~A266 & ~A265;
  assign \new_[63748]_  = ~A300 & A298;
  assign \new_[63749]_  = \new_[63748]_  & \new_[63745]_ ;
  assign \new_[63750]_  = \new_[63749]_  & \new_[63742]_ ;
  assign \new_[63754]_  = ~A168 & ~A169;
  assign \new_[63755]_  = ~A170 & \new_[63754]_ ;
  assign \new_[63759]_  = A201 & ~A200;
  assign \new_[63760]_  = A199 & \new_[63759]_ ;
  assign \new_[63761]_  = \new_[63760]_  & \new_[63755]_ ;
  assign \new_[63765]_  = ~A233 & ~A232;
  assign \new_[63766]_  = A202 & \new_[63765]_ ;
  assign \new_[63769]_  = ~A266 & ~A265;
  assign \new_[63772]_  = A299 & A298;
  assign \new_[63773]_  = \new_[63772]_  & \new_[63769]_ ;
  assign \new_[63774]_  = \new_[63773]_  & \new_[63766]_ ;
  assign \new_[63778]_  = ~A168 & ~A169;
  assign \new_[63779]_  = ~A170 & \new_[63778]_ ;
  assign \new_[63783]_  = A201 & ~A200;
  assign \new_[63784]_  = A199 & \new_[63783]_ ;
  assign \new_[63785]_  = \new_[63784]_  & \new_[63779]_ ;
  assign \new_[63789]_  = ~A233 & ~A232;
  assign \new_[63790]_  = A202 & \new_[63789]_ ;
  assign \new_[63793]_  = ~A266 & ~A265;
  assign \new_[63796]_  = ~A299 & ~A298;
  assign \new_[63797]_  = \new_[63796]_  & \new_[63793]_ ;
  assign \new_[63798]_  = \new_[63797]_  & \new_[63790]_ ;
  assign \new_[63802]_  = ~A168 & ~A169;
  assign \new_[63803]_  = ~A170 & \new_[63802]_ ;
  assign \new_[63807]_  = A201 & ~A200;
  assign \new_[63808]_  = A199 & \new_[63807]_ ;
  assign \new_[63809]_  = \new_[63808]_  & \new_[63803]_ ;
  assign \new_[63813]_  = A233 & A232;
  assign \new_[63814]_  = A203 & \new_[63813]_ ;
  assign \new_[63817]_  = ~A267 & A265;
  assign \new_[63820]_  = ~A300 & ~A299;
  assign \new_[63821]_  = \new_[63820]_  & \new_[63817]_ ;
  assign \new_[63822]_  = \new_[63821]_  & \new_[63814]_ ;
  assign \new_[63826]_  = ~A168 & ~A169;
  assign \new_[63827]_  = ~A170 & \new_[63826]_ ;
  assign \new_[63831]_  = A201 & ~A200;
  assign \new_[63832]_  = A199 & \new_[63831]_ ;
  assign \new_[63833]_  = \new_[63832]_  & \new_[63827]_ ;
  assign \new_[63837]_  = A233 & A232;
  assign \new_[63838]_  = A203 & \new_[63837]_ ;
  assign \new_[63841]_  = ~A267 & A265;
  assign \new_[63844]_  = A299 & A298;
  assign \new_[63845]_  = \new_[63844]_  & \new_[63841]_ ;
  assign \new_[63846]_  = \new_[63845]_  & \new_[63838]_ ;
  assign \new_[63850]_  = ~A168 & ~A169;
  assign \new_[63851]_  = ~A170 & \new_[63850]_ ;
  assign \new_[63855]_  = A201 & ~A200;
  assign \new_[63856]_  = A199 & \new_[63855]_ ;
  assign \new_[63857]_  = \new_[63856]_  & \new_[63851]_ ;
  assign \new_[63861]_  = A233 & A232;
  assign \new_[63862]_  = A203 & \new_[63861]_ ;
  assign \new_[63865]_  = ~A267 & A265;
  assign \new_[63868]_  = ~A299 & ~A298;
  assign \new_[63869]_  = \new_[63868]_  & \new_[63865]_ ;
  assign \new_[63870]_  = \new_[63869]_  & \new_[63862]_ ;
  assign \new_[63874]_  = ~A168 & ~A169;
  assign \new_[63875]_  = ~A170 & \new_[63874]_ ;
  assign \new_[63879]_  = A201 & ~A200;
  assign \new_[63880]_  = A199 & \new_[63879]_ ;
  assign \new_[63881]_  = \new_[63880]_  & \new_[63875]_ ;
  assign \new_[63885]_  = A233 & A232;
  assign \new_[63886]_  = A203 & \new_[63885]_ ;
  assign \new_[63889]_  = A266 & A265;
  assign \new_[63892]_  = ~A300 & ~A299;
  assign \new_[63893]_  = \new_[63892]_  & \new_[63889]_ ;
  assign \new_[63894]_  = \new_[63893]_  & \new_[63886]_ ;
  assign \new_[63898]_  = ~A168 & ~A169;
  assign \new_[63899]_  = ~A170 & \new_[63898]_ ;
  assign \new_[63903]_  = A201 & ~A200;
  assign \new_[63904]_  = A199 & \new_[63903]_ ;
  assign \new_[63905]_  = \new_[63904]_  & \new_[63899]_ ;
  assign \new_[63909]_  = A233 & A232;
  assign \new_[63910]_  = A203 & \new_[63909]_ ;
  assign \new_[63913]_  = A266 & A265;
  assign \new_[63916]_  = A299 & A298;
  assign \new_[63917]_  = \new_[63916]_  & \new_[63913]_ ;
  assign \new_[63918]_  = \new_[63917]_  & \new_[63910]_ ;
  assign \new_[63922]_  = ~A168 & ~A169;
  assign \new_[63923]_  = ~A170 & \new_[63922]_ ;
  assign \new_[63927]_  = A201 & ~A200;
  assign \new_[63928]_  = A199 & \new_[63927]_ ;
  assign \new_[63929]_  = \new_[63928]_  & \new_[63923]_ ;
  assign \new_[63933]_  = A233 & A232;
  assign \new_[63934]_  = A203 & \new_[63933]_ ;
  assign \new_[63937]_  = A266 & A265;
  assign \new_[63940]_  = ~A299 & ~A298;
  assign \new_[63941]_  = \new_[63940]_  & \new_[63937]_ ;
  assign \new_[63942]_  = \new_[63941]_  & \new_[63934]_ ;
  assign \new_[63946]_  = ~A168 & ~A169;
  assign \new_[63947]_  = ~A170 & \new_[63946]_ ;
  assign \new_[63951]_  = A201 & ~A200;
  assign \new_[63952]_  = A199 & \new_[63951]_ ;
  assign \new_[63953]_  = \new_[63952]_  & \new_[63947]_ ;
  assign \new_[63957]_  = A233 & A232;
  assign \new_[63958]_  = A203 & \new_[63957]_ ;
  assign \new_[63961]_  = ~A266 & ~A265;
  assign \new_[63964]_  = ~A300 & ~A299;
  assign \new_[63965]_  = \new_[63964]_  & \new_[63961]_ ;
  assign \new_[63966]_  = \new_[63965]_  & \new_[63958]_ ;
  assign \new_[63970]_  = ~A168 & ~A169;
  assign \new_[63971]_  = ~A170 & \new_[63970]_ ;
  assign \new_[63975]_  = A201 & ~A200;
  assign \new_[63976]_  = A199 & \new_[63975]_ ;
  assign \new_[63977]_  = \new_[63976]_  & \new_[63971]_ ;
  assign \new_[63981]_  = A233 & A232;
  assign \new_[63982]_  = A203 & \new_[63981]_ ;
  assign \new_[63985]_  = ~A266 & ~A265;
  assign \new_[63988]_  = A299 & A298;
  assign \new_[63989]_  = \new_[63988]_  & \new_[63985]_ ;
  assign \new_[63990]_  = \new_[63989]_  & \new_[63982]_ ;
  assign \new_[63994]_  = ~A168 & ~A169;
  assign \new_[63995]_  = ~A170 & \new_[63994]_ ;
  assign \new_[63999]_  = A201 & ~A200;
  assign \new_[64000]_  = A199 & \new_[63999]_ ;
  assign \new_[64001]_  = \new_[64000]_  & \new_[63995]_ ;
  assign \new_[64005]_  = A233 & A232;
  assign \new_[64006]_  = A203 & \new_[64005]_ ;
  assign \new_[64009]_  = ~A266 & ~A265;
  assign \new_[64012]_  = ~A299 & ~A298;
  assign \new_[64013]_  = \new_[64012]_  & \new_[64009]_ ;
  assign \new_[64014]_  = \new_[64013]_  & \new_[64006]_ ;
  assign \new_[64018]_  = ~A168 & ~A169;
  assign \new_[64019]_  = ~A170 & \new_[64018]_ ;
  assign \new_[64023]_  = A201 & ~A200;
  assign \new_[64024]_  = A199 & \new_[64023]_ ;
  assign \new_[64025]_  = \new_[64024]_  & \new_[64019]_ ;
  assign \new_[64029]_  = A233 & ~A232;
  assign \new_[64030]_  = A203 & \new_[64029]_ ;
  assign \new_[64033]_  = ~A299 & A298;
  assign \new_[64036]_  = A301 & A300;
  assign \new_[64037]_  = \new_[64036]_  & \new_[64033]_ ;
  assign \new_[64038]_  = \new_[64037]_  & \new_[64030]_ ;
  assign \new_[64042]_  = ~A168 & ~A169;
  assign \new_[64043]_  = ~A170 & \new_[64042]_ ;
  assign \new_[64047]_  = A201 & ~A200;
  assign \new_[64048]_  = A199 & \new_[64047]_ ;
  assign \new_[64049]_  = \new_[64048]_  & \new_[64043]_ ;
  assign \new_[64053]_  = A233 & ~A232;
  assign \new_[64054]_  = A203 & \new_[64053]_ ;
  assign \new_[64057]_  = ~A299 & A298;
  assign \new_[64060]_  = A302 & A300;
  assign \new_[64061]_  = \new_[64060]_  & \new_[64057]_ ;
  assign \new_[64062]_  = \new_[64061]_  & \new_[64054]_ ;
  assign \new_[64066]_  = ~A168 & ~A169;
  assign \new_[64067]_  = ~A170 & \new_[64066]_ ;
  assign \new_[64071]_  = A201 & ~A200;
  assign \new_[64072]_  = A199 & \new_[64071]_ ;
  assign \new_[64073]_  = \new_[64072]_  & \new_[64067]_ ;
  assign \new_[64077]_  = A233 & ~A232;
  assign \new_[64078]_  = A203 & \new_[64077]_ ;
  assign \new_[64081]_  = ~A266 & A265;
  assign \new_[64084]_  = A268 & A267;
  assign \new_[64085]_  = \new_[64084]_  & \new_[64081]_ ;
  assign \new_[64086]_  = \new_[64085]_  & \new_[64078]_ ;
  assign \new_[64090]_  = ~A168 & ~A169;
  assign \new_[64091]_  = ~A170 & \new_[64090]_ ;
  assign \new_[64095]_  = A201 & ~A200;
  assign \new_[64096]_  = A199 & \new_[64095]_ ;
  assign \new_[64097]_  = \new_[64096]_  & \new_[64091]_ ;
  assign \new_[64101]_  = A233 & ~A232;
  assign \new_[64102]_  = A203 & \new_[64101]_ ;
  assign \new_[64105]_  = ~A266 & A265;
  assign \new_[64108]_  = A269 & A267;
  assign \new_[64109]_  = \new_[64108]_  & \new_[64105]_ ;
  assign \new_[64110]_  = \new_[64109]_  & \new_[64102]_ ;
  assign \new_[64114]_  = ~A168 & ~A169;
  assign \new_[64115]_  = ~A170 & \new_[64114]_ ;
  assign \new_[64119]_  = A201 & ~A200;
  assign \new_[64120]_  = A199 & \new_[64119]_ ;
  assign \new_[64121]_  = \new_[64120]_  & \new_[64115]_ ;
  assign \new_[64125]_  = ~A234 & ~A233;
  assign \new_[64126]_  = A203 & \new_[64125]_ ;
  assign \new_[64129]_  = A266 & A265;
  assign \new_[64132]_  = ~A300 & A298;
  assign \new_[64133]_  = \new_[64132]_  & \new_[64129]_ ;
  assign \new_[64134]_  = \new_[64133]_  & \new_[64126]_ ;
  assign \new_[64138]_  = ~A168 & ~A169;
  assign \new_[64139]_  = ~A170 & \new_[64138]_ ;
  assign \new_[64143]_  = A201 & ~A200;
  assign \new_[64144]_  = A199 & \new_[64143]_ ;
  assign \new_[64145]_  = \new_[64144]_  & \new_[64139]_ ;
  assign \new_[64149]_  = ~A234 & ~A233;
  assign \new_[64150]_  = A203 & \new_[64149]_ ;
  assign \new_[64153]_  = A266 & A265;
  assign \new_[64156]_  = A299 & A298;
  assign \new_[64157]_  = \new_[64156]_  & \new_[64153]_ ;
  assign \new_[64158]_  = \new_[64157]_  & \new_[64150]_ ;
  assign \new_[64162]_  = ~A168 & ~A169;
  assign \new_[64163]_  = ~A170 & \new_[64162]_ ;
  assign \new_[64167]_  = A201 & ~A200;
  assign \new_[64168]_  = A199 & \new_[64167]_ ;
  assign \new_[64169]_  = \new_[64168]_  & \new_[64163]_ ;
  assign \new_[64173]_  = ~A234 & ~A233;
  assign \new_[64174]_  = A203 & \new_[64173]_ ;
  assign \new_[64177]_  = A266 & A265;
  assign \new_[64180]_  = ~A299 & ~A298;
  assign \new_[64181]_  = \new_[64180]_  & \new_[64177]_ ;
  assign \new_[64182]_  = \new_[64181]_  & \new_[64174]_ ;
  assign \new_[64186]_  = ~A168 & ~A169;
  assign \new_[64187]_  = ~A170 & \new_[64186]_ ;
  assign \new_[64191]_  = A201 & ~A200;
  assign \new_[64192]_  = A199 & \new_[64191]_ ;
  assign \new_[64193]_  = \new_[64192]_  & \new_[64187]_ ;
  assign \new_[64197]_  = ~A234 & ~A233;
  assign \new_[64198]_  = A203 & \new_[64197]_ ;
  assign \new_[64201]_  = ~A267 & ~A266;
  assign \new_[64204]_  = ~A300 & A298;
  assign \new_[64205]_  = \new_[64204]_  & \new_[64201]_ ;
  assign \new_[64206]_  = \new_[64205]_  & \new_[64198]_ ;
  assign \new_[64210]_  = ~A168 & ~A169;
  assign \new_[64211]_  = ~A170 & \new_[64210]_ ;
  assign \new_[64215]_  = A201 & ~A200;
  assign \new_[64216]_  = A199 & \new_[64215]_ ;
  assign \new_[64217]_  = \new_[64216]_  & \new_[64211]_ ;
  assign \new_[64221]_  = ~A234 & ~A233;
  assign \new_[64222]_  = A203 & \new_[64221]_ ;
  assign \new_[64225]_  = ~A267 & ~A266;
  assign \new_[64228]_  = A299 & A298;
  assign \new_[64229]_  = \new_[64228]_  & \new_[64225]_ ;
  assign \new_[64230]_  = \new_[64229]_  & \new_[64222]_ ;
  assign \new_[64234]_  = ~A168 & ~A169;
  assign \new_[64235]_  = ~A170 & \new_[64234]_ ;
  assign \new_[64239]_  = A201 & ~A200;
  assign \new_[64240]_  = A199 & \new_[64239]_ ;
  assign \new_[64241]_  = \new_[64240]_  & \new_[64235]_ ;
  assign \new_[64245]_  = ~A234 & ~A233;
  assign \new_[64246]_  = A203 & \new_[64245]_ ;
  assign \new_[64249]_  = ~A267 & ~A266;
  assign \new_[64252]_  = ~A299 & ~A298;
  assign \new_[64253]_  = \new_[64252]_  & \new_[64249]_ ;
  assign \new_[64254]_  = \new_[64253]_  & \new_[64246]_ ;
  assign \new_[64258]_  = ~A168 & ~A169;
  assign \new_[64259]_  = ~A170 & \new_[64258]_ ;
  assign \new_[64263]_  = A201 & ~A200;
  assign \new_[64264]_  = A199 & \new_[64263]_ ;
  assign \new_[64265]_  = \new_[64264]_  & \new_[64259]_ ;
  assign \new_[64269]_  = ~A234 & ~A233;
  assign \new_[64270]_  = A203 & \new_[64269]_ ;
  assign \new_[64273]_  = ~A266 & ~A265;
  assign \new_[64276]_  = ~A300 & A298;
  assign \new_[64277]_  = \new_[64276]_  & \new_[64273]_ ;
  assign \new_[64278]_  = \new_[64277]_  & \new_[64270]_ ;
  assign \new_[64282]_  = ~A168 & ~A169;
  assign \new_[64283]_  = ~A170 & \new_[64282]_ ;
  assign \new_[64287]_  = A201 & ~A200;
  assign \new_[64288]_  = A199 & \new_[64287]_ ;
  assign \new_[64289]_  = \new_[64288]_  & \new_[64283]_ ;
  assign \new_[64293]_  = ~A234 & ~A233;
  assign \new_[64294]_  = A203 & \new_[64293]_ ;
  assign \new_[64297]_  = ~A266 & ~A265;
  assign \new_[64300]_  = A299 & A298;
  assign \new_[64301]_  = \new_[64300]_  & \new_[64297]_ ;
  assign \new_[64302]_  = \new_[64301]_  & \new_[64294]_ ;
  assign \new_[64306]_  = ~A168 & ~A169;
  assign \new_[64307]_  = ~A170 & \new_[64306]_ ;
  assign \new_[64311]_  = A201 & ~A200;
  assign \new_[64312]_  = A199 & \new_[64311]_ ;
  assign \new_[64313]_  = \new_[64312]_  & \new_[64307]_ ;
  assign \new_[64317]_  = ~A234 & ~A233;
  assign \new_[64318]_  = A203 & \new_[64317]_ ;
  assign \new_[64321]_  = ~A266 & ~A265;
  assign \new_[64324]_  = ~A299 & ~A298;
  assign \new_[64325]_  = \new_[64324]_  & \new_[64321]_ ;
  assign \new_[64326]_  = \new_[64325]_  & \new_[64318]_ ;
  assign \new_[64330]_  = ~A168 & ~A169;
  assign \new_[64331]_  = ~A170 & \new_[64330]_ ;
  assign \new_[64335]_  = A201 & ~A200;
  assign \new_[64336]_  = A199 & \new_[64335]_ ;
  assign \new_[64337]_  = \new_[64336]_  & \new_[64331]_ ;
  assign \new_[64341]_  = ~A233 & A232;
  assign \new_[64342]_  = A203 & \new_[64341]_ ;
  assign \new_[64345]_  = A235 & A234;
  assign \new_[64348]_  = A299 & ~A298;
  assign \new_[64349]_  = \new_[64348]_  & \new_[64345]_ ;
  assign \new_[64350]_  = \new_[64349]_  & \new_[64342]_ ;
  assign \new_[64354]_  = ~A168 & ~A169;
  assign \new_[64355]_  = ~A170 & \new_[64354]_ ;
  assign \new_[64359]_  = A201 & ~A200;
  assign \new_[64360]_  = A199 & \new_[64359]_ ;
  assign \new_[64361]_  = \new_[64360]_  & \new_[64355]_ ;
  assign \new_[64365]_  = ~A233 & A232;
  assign \new_[64366]_  = A203 & \new_[64365]_ ;
  assign \new_[64369]_  = A235 & A234;
  assign \new_[64372]_  = A266 & ~A265;
  assign \new_[64373]_  = \new_[64372]_  & \new_[64369]_ ;
  assign \new_[64374]_  = \new_[64373]_  & \new_[64366]_ ;
  assign \new_[64378]_  = ~A168 & ~A169;
  assign \new_[64379]_  = ~A170 & \new_[64378]_ ;
  assign \new_[64383]_  = A201 & ~A200;
  assign \new_[64384]_  = A199 & \new_[64383]_ ;
  assign \new_[64385]_  = \new_[64384]_  & \new_[64379]_ ;
  assign \new_[64389]_  = ~A233 & A232;
  assign \new_[64390]_  = A203 & \new_[64389]_ ;
  assign \new_[64393]_  = A236 & A234;
  assign \new_[64396]_  = A299 & ~A298;
  assign \new_[64397]_  = \new_[64396]_  & \new_[64393]_ ;
  assign \new_[64398]_  = \new_[64397]_  & \new_[64390]_ ;
  assign \new_[64402]_  = ~A168 & ~A169;
  assign \new_[64403]_  = ~A170 & \new_[64402]_ ;
  assign \new_[64407]_  = A201 & ~A200;
  assign \new_[64408]_  = A199 & \new_[64407]_ ;
  assign \new_[64409]_  = \new_[64408]_  & \new_[64403]_ ;
  assign \new_[64413]_  = ~A233 & A232;
  assign \new_[64414]_  = A203 & \new_[64413]_ ;
  assign \new_[64417]_  = A236 & A234;
  assign \new_[64420]_  = A266 & ~A265;
  assign \new_[64421]_  = \new_[64420]_  & \new_[64417]_ ;
  assign \new_[64422]_  = \new_[64421]_  & \new_[64414]_ ;
  assign \new_[64426]_  = ~A168 & ~A169;
  assign \new_[64427]_  = ~A170 & \new_[64426]_ ;
  assign \new_[64431]_  = A201 & ~A200;
  assign \new_[64432]_  = A199 & \new_[64431]_ ;
  assign \new_[64433]_  = \new_[64432]_  & \new_[64427]_ ;
  assign \new_[64437]_  = ~A233 & ~A232;
  assign \new_[64438]_  = A203 & \new_[64437]_ ;
  assign \new_[64441]_  = A266 & A265;
  assign \new_[64444]_  = ~A300 & A298;
  assign \new_[64445]_  = \new_[64444]_  & \new_[64441]_ ;
  assign \new_[64446]_  = \new_[64445]_  & \new_[64438]_ ;
  assign \new_[64450]_  = ~A168 & ~A169;
  assign \new_[64451]_  = ~A170 & \new_[64450]_ ;
  assign \new_[64455]_  = A201 & ~A200;
  assign \new_[64456]_  = A199 & \new_[64455]_ ;
  assign \new_[64457]_  = \new_[64456]_  & \new_[64451]_ ;
  assign \new_[64461]_  = ~A233 & ~A232;
  assign \new_[64462]_  = A203 & \new_[64461]_ ;
  assign \new_[64465]_  = A266 & A265;
  assign \new_[64468]_  = A299 & A298;
  assign \new_[64469]_  = \new_[64468]_  & \new_[64465]_ ;
  assign \new_[64470]_  = \new_[64469]_  & \new_[64462]_ ;
  assign \new_[64474]_  = ~A168 & ~A169;
  assign \new_[64475]_  = ~A170 & \new_[64474]_ ;
  assign \new_[64479]_  = A201 & ~A200;
  assign \new_[64480]_  = A199 & \new_[64479]_ ;
  assign \new_[64481]_  = \new_[64480]_  & \new_[64475]_ ;
  assign \new_[64485]_  = ~A233 & ~A232;
  assign \new_[64486]_  = A203 & \new_[64485]_ ;
  assign \new_[64489]_  = A266 & A265;
  assign \new_[64492]_  = ~A299 & ~A298;
  assign \new_[64493]_  = \new_[64492]_  & \new_[64489]_ ;
  assign \new_[64494]_  = \new_[64493]_  & \new_[64486]_ ;
  assign \new_[64498]_  = ~A168 & ~A169;
  assign \new_[64499]_  = ~A170 & \new_[64498]_ ;
  assign \new_[64503]_  = A201 & ~A200;
  assign \new_[64504]_  = A199 & \new_[64503]_ ;
  assign \new_[64505]_  = \new_[64504]_  & \new_[64499]_ ;
  assign \new_[64509]_  = ~A233 & ~A232;
  assign \new_[64510]_  = A203 & \new_[64509]_ ;
  assign \new_[64513]_  = ~A267 & ~A266;
  assign \new_[64516]_  = ~A300 & A298;
  assign \new_[64517]_  = \new_[64516]_  & \new_[64513]_ ;
  assign \new_[64518]_  = \new_[64517]_  & \new_[64510]_ ;
  assign \new_[64522]_  = ~A168 & ~A169;
  assign \new_[64523]_  = ~A170 & \new_[64522]_ ;
  assign \new_[64527]_  = A201 & ~A200;
  assign \new_[64528]_  = A199 & \new_[64527]_ ;
  assign \new_[64529]_  = \new_[64528]_  & \new_[64523]_ ;
  assign \new_[64533]_  = ~A233 & ~A232;
  assign \new_[64534]_  = A203 & \new_[64533]_ ;
  assign \new_[64537]_  = ~A267 & ~A266;
  assign \new_[64540]_  = A299 & A298;
  assign \new_[64541]_  = \new_[64540]_  & \new_[64537]_ ;
  assign \new_[64542]_  = \new_[64541]_  & \new_[64534]_ ;
  assign \new_[64546]_  = ~A168 & ~A169;
  assign \new_[64547]_  = ~A170 & \new_[64546]_ ;
  assign \new_[64551]_  = A201 & ~A200;
  assign \new_[64552]_  = A199 & \new_[64551]_ ;
  assign \new_[64553]_  = \new_[64552]_  & \new_[64547]_ ;
  assign \new_[64557]_  = ~A233 & ~A232;
  assign \new_[64558]_  = A203 & \new_[64557]_ ;
  assign \new_[64561]_  = ~A267 & ~A266;
  assign \new_[64564]_  = ~A299 & ~A298;
  assign \new_[64565]_  = \new_[64564]_  & \new_[64561]_ ;
  assign \new_[64566]_  = \new_[64565]_  & \new_[64558]_ ;
  assign \new_[64570]_  = ~A168 & ~A169;
  assign \new_[64571]_  = ~A170 & \new_[64570]_ ;
  assign \new_[64575]_  = A201 & ~A200;
  assign \new_[64576]_  = A199 & \new_[64575]_ ;
  assign \new_[64577]_  = \new_[64576]_  & \new_[64571]_ ;
  assign \new_[64581]_  = ~A233 & ~A232;
  assign \new_[64582]_  = A203 & \new_[64581]_ ;
  assign \new_[64585]_  = ~A266 & ~A265;
  assign \new_[64588]_  = ~A300 & A298;
  assign \new_[64589]_  = \new_[64588]_  & \new_[64585]_ ;
  assign \new_[64590]_  = \new_[64589]_  & \new_[64582]_ ;
  assign \new_[64594]_  = ~A168 & ~A169;
  assign \new_[64595]_  = ~A170 & \new_[64594]_ ;
  assign \new_[64599]_  = A201 & ~A200;
  assign \new_[64600]_  = A199 & \new_[64599]_ ;
  assign \new_[64601]_  = \new_[64600]_  & \new_[64595]_ ;
  assign \new_[64605]_  = ~A233 & ~A232;
  assign \new_[64606]_  = A203 & \new_[64605]_ ;
  assign \new_[64609]_  = ~A266 & ~A265;
  assign \new_[64612]_  = A299 & A298;
  assign \new_[64613]_  = \new_[64612]_  & \new_[64609]_ ;
  assign \new_[64614]_  = \new_[64613]_  & \new_[64606]_ ;
  assign \new_[64618]_  = ~A168 & ~A169;
  assign \new_[64619]_  = ~A170 & \new_[64618]_ ;
  assign \new_[64623]_  = A201 & ~A200;
  assign \new_[64624]_  = A199 & \new_[64623]_ ;
  assign \new_[64625]_  = \new_[64624]_  & \new_[64619]_ ;
  assign \new_[64629]_  = ~A233 & ~A232;
  assign \new_[64630]_  = A203 & \new_[64629]_ ;
  assign \new_[64633]_  = ~A266 & ~A265;
  assign \new_[64636]_  = ~A299 & ~A298;
  assign \new_[64637]_  = \new_[64636]_  & \new_[64633]_ ;
  assign \new_[64638]_  = \new_[64637]_  & \new_[64630]_ ;
  assign \new_[64642]_  = ~A200 & A166;
  assign \new_[64643]_  = A168 & \new_[64642]_ ;
  assign \new_[64646]_  = ~A203 & ~A202;
  assign \new_[64649]_  = ~A235 & ~A233;
  assign \new_[64650]_  = \new_[64649]_  & \new_[64646]_ ;
  assign \new_[64651]_  = \new_[64650]_  & \new_[64643]_ ;
  assign \new_[64655]_  = ~A268 & ~A266;
  assign \new_[64656]_  = ~A236 & \new_[64655]_ ;
  assign \new_[64659]_  = A298 & ~A269;
  assign \new_[64662]_  = ~A302 & ~A301;
  assign \new_[64663]_  = \new_[64662]_  & \new_[64659]_ ;
  assign \new_[64664]_  = \new_[64663]_  & \new_[64656]_ ;
  assign \new_[64668]_  = ~A200 & A167;
  assign \new_[64669]_  = A168 & \new_[64668]_ ;
  assign \new_[64672]_  = ~A203 & ~A202;
  assign \new_[64675]_  = ~A235 & ~A233;
  assign \new_[64676]_  = \new_[64675]_  & \new_[64672]_ ;
  assign \new_[64677]_  = \new_[64676]_  & \new_[64669]_ ;
  assign \new_[64681]_  = ~A268 & ~A266;
  assign \new_[64682]_  = ~A236 & \new_[64681]_ ;
  assign \new_[64685]_  = A298 & ~A269;
  assign \new_[64688]_  = ~A302 & ~A301;
  assign \new_[64689]_  = \new_[64688]_  & \new_[64685]_ ;
  assign \new_[64690]_  = \new_[64689]_  & \new_[64682]_ ;
  assign \new_[64694]_  = ~A166 & ~A167;
  assign \new_[64695]_  = A170 & \new_[64694]_ ;
  assign \new_[64698]_  = A200 & ~A199;
  assign \new_[64701]_  = ~A235 & ~A233;
  assign \new_[64702]_  = \new_[64701]_  & \new_[64698]_ ;
  assign \new_[64703]_  = \new_[64702]_  & \new_[64695]_ ;
  assign \new_[64707]_  = ~A268 & ~A266;
  assign \new_[64708]_  = ~A236 & \new_[64707]_ ;
  assign \new_[64711]_  = A298 & ~A269;
  assign \new_[64714]_  = ~A302 & ~A301;
  assign \new_[64715]_  = \new_[64714]_  & \new_[64711]_ ;
  assign \new_[64716]_  = \new_[64715]_  & \new_[64708]_ ;
  assign \new_[64720]_  = ~A166 & ~A167;
  assign \new_[64721]_  = A170 & \new_[64720]_ ;
  assign \new_[64724]_  = ~A200 & A199;
  assign \new_[64727]_  = A202 & A201;
  assign \new_[64728]_  = \new_[64727]_  & \new_[64724]_ ;
  assign \new_[64729]_  = \new_[64728]_  & \new_[64721]_ ;
  assign \new_[64733]_  = A265 & A233;
  assign \new_[64734]_  = A232 & \new_[64733]_ ;
  assign \new_[64737]_  = ~A269 & ~A268;
  assign \new_[64740]_  = ~A300 & ~A299;
  assign \new_[64741]_  = \new_[64740]_  & \new_[64737]_ ;
  assign \new_[64742]_  = \new_[64741]_  & \new_[64734]_ ;
  assign \new_[64746]_  = ~A166 & ~A167;
  assign \new_[64747]_  = A170 & \new_[64746]_ ;
  assign \new_[64750]_  = ~A200 & A199;
  assign \new_[64753]_  = A202 & A201;
  assign \new_[64754]_  = \new_[64753]_  & \new_[64750]_ ;
  assign \new_[64755]_  = \new_[64754]_  & \new_[64747]_ ;
  assign \new_[64759]_  = A265 & A233;
  assign \new_[64760]_  = A232 & \new_[64759]_ ;
  assign \new_[64763]_  = ~A269 & ~A268;
  assign \new_[64766]_  = A299 & A298;
  assign \new_[64767]_  = \new_[64766]_  & \new_[64763]_ ;
  assign \new_[64768]_  = \new_[64767]_  & \new_[64760]_ ;
  assign \new_[64772]_  = ~A166 & ~A167;
  assign \new_[64773]_  = A170 & \new_[64772]_ ;
  assign \new_[64776]_  = ~A200 & A199;
  assign \new_[64779]_  = A202 & A201;
  assign \new_[64780]_  = \new_[64779]_  & \new_[64776]_ ;
  assign \new_[64781]_  = \new_[64780]_  & \new_[64773]_ ;
  assign \new_[64785]_  = A265 & A233;
  assign \new_[64786]_  = A232 & \new_[64785]_ ;
  assign \new_[64789]_  = ~A269 & ~A268;
  assign \new_[64792]_  = ~A299 & ~A298;
  assign \new_[64793]_  = \new_[64792]_  & \new_[64789]_ ;
  assign \new_[64794]_  = \new_[64793]_  & \new_[64786]_ ;
  assign \new_[64798]_  = ~A166 & ~A167;
  assign \new_[64799]_  = A170 & \new_[64798]_ ;
  assign \new_[64802]_  = ~A200 & A199;
  assign \new_[64805]_  = A202 & A201;
  assign \new_[64806]_  = \new_[64805]_  & \new_[64802]_ ;
  assign \new_[64807]_  = \new_[64806]_  & \new_[64799]_ ;
  assign \new_[64811]_  = A265 & A233;
  assign \new_[64812]_  = A232 & \new_[64811]_ ;
  assign \new_[64815]_  = ~A299 & ~A267;
  assign \new_[64818]_  = ~A302 & ~A301;
  assign \new_[64819]_  = \new_[64818]_  & \new_[64815]_ ;
  assign \new_[64820]_  = \new_[64819]_  & \new_[64812]_ ;
  assign \new_[64824]_  = ~A166 & ~A167;
  assign \new_[64825]_  = A170 & \new_[64824]_ ;
  assign \new_[64828]_  = ~A200 & A199;
  assign \new_[64831]_  = A202 & A201;
  assign \new_[64832]_  = \new_[64831]_  & \new_[64828]_ ;
  assign \new_[64833]_  = \new_[64832]_  & \new_[64825]_ ;
  assign \new_[64837]_  = A265 & A233;
  assign \new_[64838]_  = A232 & \new_[64837]_ ;
  assign \new_[64841]_  = ~A299 & A266;
  assign \new_[64844]_  = ~A302 & ~A301;
  assign \new_[64845]_  = \new_[64844]_  & \new_[64841]_ ;
  assign \new_[64846]_  = \new_[64845]_  & \new_[64838]_ ;
  assign \new_[64850]_  = ~A166 & ~A167;
  assign \new_[64851]_  = A170 & \new_[64850]_ ;
  assign \new_[64854]_  = ~A200 & A199;
  assign \new_[64857]_  = A202 & A201;
  assign \new_[64858]_  = \new_[64857]_  & \new_[64854]_ ;
  assign \new_[64859]_  = \new_[64858]_  & \new_[64851]_ ;
  assign \new_[64863]_  = ~A265 & A233;
  assign \new_[64864]_  = A232 & \new_[64863]_ ;
  assign \new_[64867]_  = ~A299 & ~A266;
  assign \new_[64870]_  = ~A302 & ~A301;
  assign \new_[64871]_  = \new_[64870]_  & \new_[64867]_ ;
  assign \new_[64872]_  = \new_[64871]_  & \new_[64864]_ ;
  assign \new_[64876]_  = ~A166 & ~A167;
  assign \new_[64877]_  = A170 & \new_[64876]_ ;
  assign \new_[64880]_  = ~A200 & A199;
  assign \new_[64883]_  = A202 & A201;
  assign \new_[64884]_  = \new_[64883]_  & \new_[64880]_ ;
  assign \new_[64885]_  = \new_[64884]_  & \new_[64877]_ ;
  assign \new_[64889]_  = ~A236 & ~A235;
  assign \new_[64890]_  = ~A233 & \new_[64889]_ ;
  assign \new_[64893]_  = A266 & A265;
  assign \new_[64896]_  = ~A300 & A298;
  assign \new_[64897]_  = \new_[64896]_  & \new_[64893]_ ;
  assign \new_[64898]_  = \new_[64897]_  & \new_[64890]_ ;
  assign \new_[64902]_  = ~A166 & ~A167;
  assign \new_[64903]_  = A170 & \new_[64902]_ ;
  assign \new_[64906]_  = ~A200 & A199;
  assign \new_[64909]_  = A202 & A201;
  assign \new_[64910]_  = \new_[64909]_  & \new_[64906]_ ;
  assign \new_[64911]_  = \new_[64910]_  & \new_[64903]_ ;
  assign \new_[64915]_  = ~A236 & ~A235;
  assign \new_[64916]_  = ~A233 & \new_[64915]_ ;
  assign \new_[64919]_  = A266 & A265;
  assign \new_[64922]_  = A299 & A298;
  assign \new_[64923]_  = \new_[64922]_  & \new_[64919]_ ;
  assign \new_[64924]_  = \new_[64923]_  & \new_[64916]_ ;
  assign \new_[64928]_  = ~A166 & ~A167;
  assign \new_[64929]_  = A170 & \new_[64928]_ ;
  assign \new_[64932]_  = ~A200 & A199;
  assign \new_[64935]_  = A202 & A201;
  assign \new_[64936]_  = \new_[64935]_  & \new_[64932]_ ;
  assign \new_[64937]_  = \new_[64936]_  & \new_[64929]_ ;
  assign \new_[64941]_  = ~A236 & ~A235;
  assign \new_[64942]_  = ~A233 & \new_[64941]_ ;
  assign \new_[64945]_  = A266 & A265;
  assign \new_[64948]_  = ~A299 & ~A298;
  assign \new_[64949]_  = \new_[64948]_  & \new_[64945]_ ;
  assign \new_[64950]_  = \new_[64949]_  & \new_[64942]_ ;
  assign \new_[64954]_  = ~A166 & ~A167;
  assign \new_[64955]_  = A170 & \new_[64954]_ ;
  assign \new_[64958]_  = ~A200 & A199;
  assign \new_[64961]_  = A202 & A201;
  assign \new_[64962]_  = \new_[64961]_  & \new_[64958]_ ;
  assign \new_[64963]_  = \new_[64962]_  & \new_[64955]_ ;
  assign \new_[64967]_  = ~A236 & ~A235;
  assign \new_[64968]_  = ~A233 & \new_[64967]_ ;
  assign \new_[64971]_  = ~A267 & ~A266;
  assign \new_[64974]_  = ~A300 & A298;
  assign \new_[64975]_  = \new_[64974]_  & \new_[64971]_ ;
  assign \new_[64976]_  = \new_[64975]_  & \new_[64968]_ ;
  assign \new_[64980]_  = ~A166 & ~A167;
  assign \new_[64981]_  = A170 & \new_[64980]_ ;
  assign \new_[64984]_  = ~A200 & A199;
  assign \new_[64987]_  = A202 & A201;
  assign \new_[64988]_  = \new_[64987]_  & \new_[64984]_ ;
  assign \new_[64989]_  = \new_[64988]_  & \new_[64981]_ ;
  assign \new_[64993]_  = ~A236 & ~A235;
  assign \new_[64994]_  = ~A233 & \new_[64993]_ ;
  assign \new_[64997]_  = ~A267 & ~A266;
  assign \new_[65000]_  = A299 & A298;
  assign \new_[65001]_  = \new_[65000]_  & \new_[64997]_ ;
  assign \new_[65002]_  = \new_[65001]_  & \new_[64994]_ ;
  assign \new_[65006]_  = ~A166 & ~A167;
  assign \new_[65007]_  = A170 & \new_[65006]_ ;
  assign \new_[65010]_  = ~A200 & A199;
  assign \new_[65013]_  = A202 & A201;
  assign \new_[65014]_  = \new_[65013]_  & \new_[65010]_ ;
  assign \new_[65015]_  = \new_[65014]_  & \new_[65007]_ ;
  assign \new_[65019]_  = ~A236 & ~A235;
  assign \new_[65020]_  = ~A233 & \new_[65019]_ ;
  assign \new_[65023]_  = ~A267 & ~A266;
  assign \new_[65026]_  = ~A299 & ~A298;
  assign \new_[65027]_  = \new_[65026]_  & \new_[65023]_ ;
  assign \new_[65028]_  = \new_[65027]_  & \new_[65020]_ ;
  assign \new_[65032]_  = ~A166 & ~A167;
  assign \new_[65033]_  = A170 & \new_[65032]_ ;
  assign \new_[65036]_  = ~A200 & A199;
  assign \new_[65039]_  = A202 & A201;
  assign \new_[65040]_  = \new_[65039]_  & \new_[65036]_ ;
  assign \new_[65041]_  = \new_[65040]_  & \new_[65033]_ ;
  assign \new_[65045]_  = ~A236 & ~A235;
  assign \new_[65046]_  = ~A233 & \new_[65045]_ ;
  assign \new_[65049]_  = ~A266 & ~A265;
  assign \new_[65052]_  = ~A300 & A298;
  assign \new_[65053]_  = \new_[65052]_  & \new_[65049]_ ;
  assign \new_[65054]_  = \new_[65053]_  & \new_[65046]_ ;
  assign \new_[65058]_  = ~A166 & ~A167;
  assign \new_[65059]_  = A170 & \new_[65058]_ ;
  assign \new_[65062]_  = ~A200 & A199;
  assign \new_[65065]_  = A202 & A201;
  assign \new_[65066]_  = \new_[65065]_  & \new_[65062]_ ;
  assign \new_[65067]_  = \new_[65066]_  & \new_[65059]_ ;
  assign \new_[65071]_  = ~A236 & ~A235;
  assign \new_[65072]_  = ~A233 & \new_[65071]_ ;
  assign \new_[65075]_  = ~A266 & ~A265;
  assign \new_[65078]_  = A299 & A298;
  assign \new_[65079]_  = \new_[65078]_  & \new_[65075]_ ;
  assign \new_[65080]_  = \new_[65079]_  & \new_[65072]_ ;
  assign \new_[65084]_  = ~A166 & ~A167;
  assign \new_[65085]_  = A170 & \new_[65084]_ ;
  assign \new_[65088]_  = ~A200 & A199;
  assign \new_[65091]_  = A202 & A201;
  assign \new_[65092]_  = \new_[65091]_  & \new_[65088]_ ;
  assign \new_[65093]_  = \new_[65092]_  & \new_[65085]_ ;
  assign \new_[65097]_  = ~A236 & ~A235;
  assign \new_[65098]_  = ~A233 & \new_[65097]_ ;
  assign \new_[65101]_  = ~A266 & ~A265;
  assign \new_[65104]_  = ~A299 & ~A298;
  assign \new_[65105]_  = \new_[65104]_  & \new_[65101]_ ;
  assign \new_[65106]_  = \new_[65105]_  & \new_[65098]_ ;
  assign \new_[65110]_  = ~A166 & ~A167;
  assign \new_[65111]_  = A170 & \new_[65110]_ ;
  assign \new_[65114]_  = ~A200 & A199;
  assign \new_[65117]_  = A202 & A201;
  assign \new_[65118]_  = \new_[65117]_  & \new_[65114]_ ;
  assign \new_[65119]_  = \new_[65118]_  & \new_[65111]_ ;
  assign \new_[65123]_  = A265 & ~A234;
  assign \new_[65124]_  = ~A233 & \new_[65123]_ ;
  assign \new_[65127]_  = A298 & A266;
  assign \new_[65130]_  = ~A302 & ~A301;
  assign \new_[65131]_  = \new_[65130]_  & \new_[65127]_ ;
  assign \new_[65132]_  = \new_[65131]_  & \new_[65124]_ ;
  assign \new_[65136]_  = ~A166 & ~A167;
  assign \new_[65137]_  = A170 & \new_[65136]_ ;
  assign \new_[65140]_  = ~A200 & A199;
  assign \new_[65143]_  = A202 & A201;
  assign \new_[65144]_  = \new_[65143]_  & \new_[65140]_ ;
  assign \new_[65145]_  = \new_[65144]_  & \new_[65137]_ ;
  assign \new_[65149]_  = ~A266 & ~A234;
  assign \new_[65150]_  = ~A233 & \new_[65149]_ ;
  assign \new_[65153]_  = ~A269 & ~A268;
  assign \new_[65156]_  = ~A300 & A298;
  assign \new_[65157]_  = \new_[65156]_  & \new_[65153]_ ;
  assign \new_[65158]_  = \new_[65157]_  & \new_[65150]_ ;
  assign \new_[65162]_  = ~A166 & ~A167;
  assign \new_[65163]_  = A170 & \new_[65162]_ ;
  assign \new_[65166]_  = ~A200 & A199;
  assign \new_[65169]_  = A202 & A201;
  assign \new_[65170]_  = \new_[65169]_  & \new_[65166]_ ;
  assign \new_[65171]_  = \new_[65170]_  & \new_[65163]_ ;
  assign \new_[65175]_  = ~A266 & ~A234;
  assign \new_[65176]_  = ~A233 & \new_[65175]_ ;
  assign \new_[65179]_  = ~A269 & ~A268;
  assign \new_[65182]_  = A299 & A298;
  assign \new_[65183]_  = \new_[65182]_  & \new_[65179]_ ;
  assign \new_[65184]_  = \new_[65183]_  & \new_[65176]_ ;
  assign \new_[65188]_  = ~A166 & ~A167;
  assign \new_[65189]_  = A170 & \new_[65188]_ ;
  assign \new_[65192]_  = ~A200 & A199;
  assign \new_[65195]_  = A202 & A201;
  assign \new_[65196]_  = \new_[65195]_  & \new_[65192]_ ;
  assign \new_[65197]_  = \new_[65196]_  & \new_[65189]_ ;
  assign \new_[65201]_  = ~A266 & ~A234;
  assign \new_[65202]_  = ~A233 & \new_[65201]_ ;
  assign \new_[65205]_  = ~A269 & ~A268;
  assign \new_[65208]_  = ~A299 & ~A298;
  assign \new_[65209]_  = \new_[65208]_  & \new_[65205]_ ;
  assign \new_[65210]_  = \new_[65209]_  & \new_[65202]_ ;
  assign \new_[65214]_  = ~A166 & ~A167;
  assign \new_[65215]_  = A170 & \new_[65214]_ ;
  assign \new_[65218]_  = ~A200 & A199;
  assign \new_[65221]_  = A202 & A201;
  assign \new_[65222]_  = \new_[65221]_  & \new_[65218]_ ;
  assign \new_[65223]_  = \new_[65222]_  & \new_[65215]_ ;
  assign \new_[65227]_  = ~A266 & ~A234;
  assign \new_[65228]_  = ~A233 & \new_[65227]_ ;
  assign \new_[65231]_  = A298 & ~A267;
  assign \new_[65234]_  = ~A302 & ~A301;
  assign \new_[65235]_  = \new_[65234]_  & \new_[65231]_ ;
  assign \new_[65236]_  = \new_[65235]_  & \new_[65228]_ ;
  assign \new_[65240]_  = ~A166 & ~A167;
  assign \new_[65241]_  = A170 & \new_[65240]_ ;
  assign \new_[65244]_  = ~A200 & A199;
  assign \new_[65247]_  = A202 & A201;
  assign \new_[65248]_  = \new_[65247]_  & \new_[65244]_ ;
  assign \new_[65249]_  = \new_[65248]_  & \new_[65241]_ ;
  assign \new_[65253]_  = ~A265 & ~A234;
  assign \new_[65254]_  = ~A233 & \new_[65253]_ ;
  assign \new_[65257]_  = A298 & ~A266;
  assign \new_[65260]_  = ~A302 & ~A301;
  assign \new_[65261]_  = \new_[65260]_  & \new_[65257]_ ;
  assign \new_[65262]_  = \new_[65261]_  & \new_[65254]_ ;
  assign \new_[65266]_  = ~A166 & ~A167;
  assign \new_[65267]_  = A170 & \new_[65266]_ ;
  assign \new_[65270]_  = ~A200 & A199;
  assign \new_[65273]_  = A202 & A201;
  assign \new_[65274]_  = \new_[65273]_  & \new_[65270]_ ;
  assign \new_[65275]_  = \new_[65274]_  & \new_[65267]_ ;
  assign \new_[65279]_  = A265 & ~A233;
  assign \new_[65280]_  = ~A232 & \new_[65279]_ ;
  assign \new_[65283]_  = A298 & A266;
  assign \new_[65286]_  = ~A302 & ~A301;
  assign \new_[65287]_  = \new_[65286]_  & \new_[65283]_ ;
  assign \new_[65288]_  = \new_[65287]_  & \new_[65280]_ ;
  assign \new_[65292]_  = ~A166 & ~A167;
  assign \new_[65293]_  = A170 & \new_[65292]_ ;
  assign \new_[65296]_  = ~A200 & A199;
  assign \new_[65299]_  = A202 & A201;
  assign \new_[65300]_  = \new_[65299]_  & \new_[65296]_ ;
  assign \new_[65301]_  = \new_[65300]_  & \new_[65293]_ ;
  assign \new_[65305]_  = ~A266 & ~A233;
  assign \new_[65306]_  = ~A232 & \new_[65305]_ ;
  assign \new_[65309]_  = ~A269 & ~A268;
  assign \new_[65312]_  = ~A300 & A298;
  assign \new_[65313]_  = \new_[65312]_  & \new_[65309]_ ;
  assign \new_[65314]_  = \new_[65313]_  & \new_[65306]_ ;
  assign \new_[65318]_  = ~A166 & ~A167;
  assign \new_[65319]_  = A170 & \new_[65318]_ ;
  assign \new_[65322]_  = ~A200 & A199;
  assign \new_[65325]_  = A202 & A201;
  assign \new_[65326]_  = \new_[65325]_  & \new_[65322]_ ;
  assign \new_[65327]_  = \new_[65326]_  & \new_[65319]_ ;
  assign \new_[65331]_  = ~A266 & ~A233;
  assign \new_[65332]_  = ~A232 & \new_[65331]_ ;
  assign \new_[65335]_  = ~A269 & ~A268;
  assign \new_[65338]_  = A299 & A298;
  assign \new_[65339]_  = \new_[65338]_  & \new_[65335]_ ;
  assign \new_[65340]_  = \new_[65339]_  & \new_[65332]_ ;
  assign \new_[65344]_  = ~A166 & ~A167;
  assign \new_[65345]_  = A170 & \new_[65344]_ ;
  assign \new_[65348]_  = ~A200 & A199;
  assign \new_[65351]_  = A202 & A201;
  assign \new_[65352]_  = \new_[65351]_  & \new_[65348]_ ;
  assign \new_[65353]_  = \new_[65352]_  & \new_[65345]_ ;
  assign \new_[65357]_  = ~A266 & ~A233;
  assign \new_[65358]_  = ~A232 & \new_[65357]_ ;
  assign \new_[65361]_  = ~A269 & ~A268;
  assign \new_[65364]_  = ~A299 & ~A298;
  assign \new_[65365]_  = \new_[65364]_  & \new_[65361]_ ;
  assign \new_[65366]_  = \new_[65365]_  & \new_[65358]_ ;
  assign \new_[65370]_  = ~A166 & ~A167;
  assign \new_[65371]_  = A170 & \new_[65370]_ ;
  assign \new_[65374]_  = ~A200 & A199;
  assign \new_[65377]_  = A202 & A201;
  assign \new_[65378]_  = \new_[65377]_  & \new_[65374]_ ;
  assign \new_[65379]_  = \new_[65378]_  & \new_[65371]_ ;
  assign \new_[65383]_  = ~A266 & ~A233;
  assign \new_[65384]_  = ~A232 & \new_[65383]_ ;
  assign \new_[65387]_  = A298 & ~A267;
  assign \new_[65390]_  = ~A302 & ~A301;
  assign \new_[65391]_  = \new_[65390]_  & \new_[65387]_ ;
  assign \new_[65392]_  = \new_[65391]_  & \new_[65384]_ ;
  assign \new_[65396]_  = ~A166 & ~A167;
  assign \new_[65397]_  = A170 & \new_[65396]_ ;
  assign \new_[65400]_  = ~A200 & A199;
  assign \new_[65403]_  = A202 & A201;
  assign \new_[65404]_  = \new_[65403]_  & \new_[65400]_ ;
  assign \new_[65405]_  = \new_[65404]_  & \new_[65397]_ ;
  assign \new_[65409]_  = ~A265 & ~A233;
  assign \new_[65410]_  = ~A232 & \new_[65409]_ ;
  assign \new_[65413]_  = A298 & ~A266;
  assign \new_[65416]_  = ~A302 & ~A301;
  assign \new_[65417]_  = \new_[65416]_  & \new_[65413]_ ;
  assign \new_[65418]_  = \new_[65417]_  & \new_[65410]_ ;
  assign \new_[65422]_  = ~A166 & ~A167;
  assign \new_[65423]_  = A170 & \new_[65422]_ ;
  assign \new_[65426]_  = ~A200 & A199;
  assign \new_[65429]_  = A203 & A201;
  assign \new_[65430]_  = \new_[65429]_  & \new_[65426]_ ;
  assign \new_[65431]_  = \new_[65430]_  & \new_[65423]_ ;
  assign \new_[65435]_  = A265 & A233;
  assign \new_[65436]_  = A232 & \new_[65435]_ ;
  assign \new_[65439]_  = ~A269 & ~A268;
  assign \new_[65442]_  = ~A300 & ~A299;
  assign \new_[65443]_  = \new_[65442]_  & \new_[65439]_ ;
  assign \new_[65444]_  = \new_[65443]_  & \new_[65436]_ ;
  assign \new_[65448]_  = ~A166 & ~A167;
  assign \new_[65449]_  = A170 & \new_[65448]_ ;
  assign \new_[65452]_  = ~A200 & A199;
  assign \new_[65455]_  = A203 & A201;
  assign \new_[65456]_  = \new_[65455]_  & \new_[65452]_ ;
  assign \new_[65457]_  = \new_[65456]_  & \new_[65449]_ ;
  assign \new_[65461]_  = A265 & A233;
  assign \new_[65462]_  = A232 & \new_[65461]_ ;
  assign \new_[65465]_  = ~A269 & ~A268;
  assign \new_[65468]_  = A299 & A298;
  assign \new_[65469]_  = \new_[65468]_  & \new_[65465]_ ;
  assign \new_[65470]_  = \new_[65469]_  & \new_[65462]_ ;
  assign \new_[65474]_  = ~A166 & ~A167;
  assign \new_[65475]_  = A170 & \new_[65474]_ ;
  assign \new_[65478]_  = ~A200 & A199;
  assign \new_[65481]_  = A203 & A201;
  assign \new_[65482]_  = \new_[65481]_  & \new_[65478]_ ;
  assign \new_[65483]_  = \new_[65482]_  & \new_[65475]_ ;
  assign \new_[65487]_  = A265 & A233;
  assign \new_[65488]_  = A232 & \new_[65487]_ ;
  assign \new_[65491]_  = ~A269 & ~A268;
  assign \new_[65494]_  = ~A299 & ~A298;
  assign \new_[65495]_  = \new_[65494]_  & \new_[65491]_ ;
  assign \new_[65496]_  = \new_[65495]_  & \new_[65488]_ ;
  assign \new_[65500]_  = ~A166 & ~A167;
  assign \new_[65501]_  = A170 & \new_[65500]_ ;
  assign \new_[65504]_  = ~A200 & A199;
  assign \new_[65507]_  = A203 & A201;
  assign \new_[65508]_  = \new_[65507]_  & \new_[65504]_ ;
  assign \new_[65509]_  = \new_[65508]_  & \new_[65501]_ ;
  assign \new_[65513]_  = A265 & A233;
  assign \new_[65514]_  = A232 & \new_[65513]_ ;
  assign \new_[65517]_  = ~A299 & ~A267;
  assign \new_[65520]_  = ~A302 & ~A301;
  assign \new_[65521]_  = \new_[65520]_  & \new_[65517]_ ;
  assign \new_[65522]_  = \new_[65521]_  & \new_[65514]_ ;
  assign \new_[65526]_  = ~A166 & ~A167;
  assign \new_[65527]_  = A170 & \new_[65526]_ ;
  assign \new_[65530]_  = ~A200 & A199;
  assign \new_[65533]_  = A203 & A201;
  assign \new_[65534]_  = \new_[65533]_  & \new_[65530]_ ;
  assign \new_[65535]_  = \new_[65534]_  & \new_[65527]_ ;
  assign \new_[65539]_  = A265 & A233;
  assign \new_[65540]_  = A232 & \new_[65539]_ ;
  assign \new_[65543]_  = ~A299 & A266;
  assign \new_[65546]_  = ~A302 & ~A301;
  assign \new_[65547]_  = \new_[65546]_  & \new_[65543]_ ;
  assign \new_[65548]_  = \new_[65547]_  & \new_[65540]_ ;
  assign \new_[65552]_  = ~A166 & ~A167;
  assign \new_[65553]_  = A170 & \new_[65552]_ ;
  assign \new_[65556]_  = ~A200 & A199;
  assign \new_[65559]_  = A203 & A201;
  assign \new_[65560]_  = \new_[65559]_  & \new_[65556]_ ;
  assign \new_[65561]_  = \new_[65560]_  & \new_[65553]_ ;
  assign \new_[65565]_  = ~A265 & A233;
  assign \new_[65566]_  = A232 & \new_[65565]_ ;
  assign \new_[65569]_  = ~A299 & ~A266;
  assign \new_[65572]_  = ~A302 & ~A301;
  assign \new_[65573]_  = \new_[65572]_  & \new_[65569]_ ;
  assign \new_[65574]_  = \new_[65573]_  & \new_[65566]_ ;
  assign \new_[65578]_  = ~A166 & ~A167;
  assign \new_[65579]_  = A170 & \new_[65578]_ ;
  assign \new_[65582]_  = ~A200 & A199;
  assign \new_[65585]_  = A203 & A201;
  assign \new_[65586]_  = \new_[65585]_  & \new_[65582]_ ;
  assign \new_[65587]_  = \new_[65586]_  & \new_[65579]_ ;
  assign \new_[65591]_  = ~A236 & ~A235;
  assign \new_[65592]_  = ~A233 & \new_[65591]_ ;
  assign \new_[65595]_  = A266 & A265;
  assign \new_[65598]_  = ~A300 & A298;
  assign \new_[65599]_  = \new_[65598]_  & \new_[65595]_ ;
  assign \new_[65600]_  = \new_[65599]_  & \new_[65592]_ ;
  assign \new_[65604]_  = ~A166 & ~A167;
  assign \new_[65605]_  = A170 & \new_[65604]_ ;
  assign \new_[65608]_  = ~A200 & A199;
  assign \new_[65611]_  = A203 & A201;
  assign \new_[65612]_  = \new_[65611]_  & \new_[65608]_ ;
  assign \new_[65613]_  = \new_[65612]_  & \new_[65605]_ ;
  assign \new_[65617]_  = ~A236 & ~A235;
  assign \new_[65618]_  = ~A233 & \new_[65617]_ ;
  assign \new_[65621]_  = A266 & A265;
  assign \new_[65624]_  = A299 & A298;
  assign \new_[65625]_  = \new_[65624]_  & \new_[65621]_ ;
  assign \new_[65626]_  = \new_[65625]_  & \new_[65618]_ ;
  assign \new_[65630]_  = ~A166 & ~A167;
  assign \new_[65631]_  = A170 & \new_[65630]_ ;
  assign \new_[65634]_  = ~A200 & A199;
  assign \new_[65637]_  = A203 & A201;
  assign \new_[65638]_  = \new_[65637]_  & \new_[65634]_ ;
  assign \new_[65639]_  = \new_[65638]_  & \new_[65631]_ ;
  assign \new_[65643]_  = ~A236 & ~A235;
  assign \new_[65644]_  = ~A233 & \new_[65643]_ ;
  assign \new_[65647]_  = A266 & A265;
  assign \new_[65650]_  = ~A299 & ~A298;
  assign \new_[65651]_  = \new_[65650]_  & \new_[65647]_ ;
  assign \new_[65652]_  = \new_[65651]_  & \new_[65644]_ ;
  assign \new_[65656]_  = ~A166 & ~A167;
  assign \new_[65657]_  = A170 & \new_[65656]_ ;
  assign \new_[65660]_  = ~A200 & A199;
  assign \new_[65663]_  = A203 & A201;
  assign \new_[65664]_  = \new_[65663]_  & \new_[65660]_ ;
  assign \new_[65665]_  = \new_[65664]_  & \new_[65657]_ ;
  assign \new_[65669]_  = ~A236 & ~A235;
  assign \new_[65670]_  = ~A233 & \new_[65669]_ ;
  assign \new_[65673]_  = ~A267 & ~A266;
  assign \new_[65676]_  = ~A300 & A298;
  assign \new_[65677]_  = \new_[65676]_  & \new_[65673]_ ;
  assign \new_[65678]_  = \new_[65677]_  & \new_[65670]_ ;
  assign \new_[65682]_  = ~A166 & ~A167;
  assign \new_[65683]_  = A170 & \new_[65682]_ ;
  assign \new_[65686]_  = ~A200 & A199;
  assign \new_[65689]_  = A203 & A201;
  assign \new_[65690]_  = \new_[65689]_  & \new_[65686]_ ;
  assign \new_[65691]_  = \new_[65690]_  & \new_[65683]_ ;
  assign \new_[65695]_  = ~A236 & ~A235;
  assign \new_[65696]_  = ~A233 & \new_[65695]_ ;
  assign \new_[65699]_  = ~A267 & ~A266;
  assign \new_[65702]_  = A299 & A298;
  assign \new_[65703]_  = \new_[65702]_  & \new_[65699]_ ;
  assign \new_[65704]_  = \new_[65703]_  & \new_[65696]_ ;
  assign \new_[65708]_  = ~A166 & ~A167;
  assign \new_[65709]_  = A170 & \new_[65708]_ ;
  assign \new_[65712]_  = ~A200 & A199;
  assign \new_[65715]_  = A203 & A201;
  assign \new_[65716]_  = \new_[65715]_  & \new_[65712]_ ;
  assign \new_[65717]_  = \new_[65716]_  & \new_[65709]_ ;
  assign \new_[65721]_  = ~A236 & ~A235;
  assign \new_[65722]_  = ~A233 & \new_[65721]_ ;
  assign \new_[65725]_  = ~A267 & ~A266;
  assign \new_[65728]_  = ~A299 & ~A298;
  assign \new_[65729]_  = \new_[65728]_  & \new_[65725]_ ;
  assign \new_[65730]_  = \new_[65729]_  & \new_[65722]_ ;
  assign \new_[65734]_  = ~A166 & ~A167;
  assign \new_[65735]_  = A170 & \new_[65734]_ ;
  assign \new_[65738]_  = ~A200 & A199;
  assign \new_[65741]_  = A203 & A201;
  assign \new_[65742]_  = \new_[65741]_  & \new_[65738]_ ;
  assign \new_[65743]_  = \new_[65742]_  & \new_[65735]_ ;
  assign \new_[65747]_  = ~A236 & ~A235;
  assign \new_[65748]_  = ~A233 & \new_[65747]_ ;
  assign \new_[65751]_  = ~A266 & ~A265;
  assign \new_[65754]_  = ~A300 & A298;
  assign \new_[65755]_  = \new_[65754]_  & \new_[65751]_ ;
  assign \new_[65756]_  = \new_[65755]_  & \new_[65748]_ ;
  assign \new_[65760]_  = ~A166 & ~A167;
  assign \new_[65761]_  = A170 & \new_[65760]_ ;
  assign \new_[65764]_  = ~A200 & A199;
  assign \new_[65767]_  = A203 & A201;
  assign \new_[65768]_  = \new_[65767]_  & \new_[65764]_ ;
  assign \new_[65769]_  = \new_[65768]_  & \new_[65761]_ ;
  assign \new_[65773]_  = ~A236 & ~A235;
  assign \new_[65774]_  = ~A233 & \new_[65773]_ ;
  assign \new_[65777]_  = ~A266 & ~A265;
  assign \new_[65780]_  = A299 & A298;
  assign \new_[65781]_  = \new_[65780]_  & \new_[65777]_ ;
  assign \new_[65782]_  = \new_[65781]_  & \new_[65774]_ ;
  assign \new_[65786]_  = ~A166 & ~A167;
  assign \new_[65787]_  = A170 & \new_[65786]_ ;
  assign \new_[65790]_  = ~A200 & A199;
  assign \new_[65793]_  = A203 & A201;
  assign \new_[65794]_  = \new_[65793]_  & \new_[65790]_ ;
  assign \new_[65795]_  = \new_[65794]_  & \new_[65787]_ ;
  assign \new_[65799]_  = ~A236 & ~A235;
  assign \new_[65800]_  = ~A233 & \new_[65799]_ ;
  assign \new_[65803]_  = ~A266 & ~A265;
  assign \new_[65806]_  = ~A299 & ~A298;
  assign \new_[65807]_  = \new_[65806]_  & \new_[65803]_ ;
  assign \new_[65808]_  = \new_[65807]_  & \new_[65800]_ ;
  assign \new_[65812]_  = ~A166 & ~A167;
  assign \new_[65813]_  = A170 & \new_[65812]_ ;
  assign \new_[65816]_  = ~A200 & A199;
  assign \new_[65819]_  = A203 & A201;
  assign \new_[65820]_  = \new_[65819]_  & \new_[65816]_ ;
  assign \new_[65821]_  = \new_[65820]_  & \new_[65813]_ ;
  assign \new_[65825]_  = A265 & ~A234;
  assign \new_[65826]_  = ~A233 & \new_[65825]_ ;
  assign \new_[65829]_  = A298 & A266;
  assign \new_[65832]_  = ~A302 & ~A301;
  assign \new_[65833]_  = \new_[65832]_  & \new_[65829]_ ;
  assign \new_[65834]_  = \new_[65833]_  & \new_[65826]_ ;
  assign \new_[65838]_  = ~A166 & ~A167;
  assign \new_[65839]_  = A170 & \new_[65838]_ ;
  assign \new_[65842]_  = ~A200 & A199;
  assign \new_[65845]_  = A203 & A201;
  assign \new_[65846]_  = \new_[65845]_  & \new_[65842]_ ;
  assign \new_[65847]_  = \new_[65846]_  & \new_[65839]_ ;
  assign \new_[65851]_  = ~A266 & ~A234;
  assign \new_[65852]_  = ~A233 & \new_[65851]_ ;
  assign \new_[65855]_  = ~A269 & ~A268;
  assign \new_[65858]_  = ~A300 & A298;
  assign \new_[65859]_  = \new_[65858]_  & \new_[65855]_ ;
  assign \new_[65860]_  = \new_[65859]_  & \new_[65852]_ ;
  assign \new_[65864]_  = ~A166 & ~A167;
  assign \new_[65865]_  = A170 & \new_[65864]_ ;
  assign \new_[65868]_  = ~A200 & A199;
  assign \new_[65871]_  = A203 & A201;
  assign \new_[65872]_  = \new_[65871]_  & \new_[65868]_ ;
  assign \new_[65873]_  = \new_[65872]_  & \new_[65865]_ ;
  assign \new_[65877]_  = ~A266 & ~A234;
  assign \new_[65878]_  = ~A233 & \new_[65877]_ ;
  assign \new_[65881]_  = ~A269 & ~A268;
  assign \new_[65884]_  = A299 & A298;
  assign \new_[65885]_  = \new_[65884]_  & \new_[65881]_ ;
  assign \new_[65886]_  = \new_[65885]_  & \new_[65878]_ ;
  assign \new_[65890]_  = ~A166 & ~A167;
  assign \new_[65891]_  = A170 & \new_[65890]_ ;
  assign \new_[65894]_  = ~A200 & A199;
  assign \new_[65897]_  = A203 & A201;
  assign \new_[65898]_  = \new_[65897]_  & \new_[65894]_ ;
  assign \new_[65899]_  = \new_[65898]_  & \new_[65891]_ ;
  assign \new_[65903]_  = ~A266 & ~A234;
  assign \new_[65904]_  = ~A233 & \new_[65903]_ ;
  assign \new_[65907]_  = ~A269 & ~A268;
  assign \new_[65910]_  = ~A299 & ~A298;
  assign \new_[65911]_  = \new_[65910]_  & \new_[65907]_ ;
  assign \new_[65912]_  = \new_[65911]_  & \new_[65904]_ ;
  assign \new_[65916]_  = ~A166 & ~A167;
  assign \new_[65917]_  = A170 & \new_[65916]_ ;
  assign \new_[65920]_  = ~A200 & A199;
  assign \new_[65923]_  = A203 & A201;
  assign \new_[65924]_  = \new_[65923]_  & \new_[65920]_ ;
  assign \new_[65925]_  = \new_[65924]_  & \new_[65917]_ ;
  assign \new_[65929]_  = ~A266 & ~A234;
  assign \new_[65930]_  = ~A233 & \new_[65929]_ ;
  assign \new_[65933]_  = A298 & ~A267;
  assign \new_[65936]_  = ~A302 & ~A301;
  assign \new_[65937]_  = \new_[65936]_  & \new_[65933]_ ;
  assign \new_[65938]_  = \new_[65937]_  & \new_[65930]_ ;
  assign \new_[65942]_  = ~A166 & ~A167;
  assign \new_[65943]_  = A170 & \new_[65942]_ ;
  assign \new_[65946]_  = ~A200 & A199;
  assign \new_[65949]_  = A203 & A201;
  assign \new_[65950]_  = \new_[65949]_  & \new_[65946]_ ;
  assign \new_[65951]_  = \new_[65950]_  & \new_[65943]_ ;
  assign \new_[65955]_  = ~A265 & ~A234;
  assign \new_[65956]_  = ~A233 & \new_[65955]_ ;
  assign \new_[65959]_  = A298 & ~A266;
  assign \new_[65962]_  = ~A302 & ~A301;
  assign \new_[65963]_  = \new_[65962]_  & \new_[65959]_ ;
  assign \new_[65964]_  = \new_[65963]_  & \new_[65956]_ ;
  assign \new_[65968]_  = ~A166 & ~A167;
  assign \new_[65969]_  = A170 & \new_[65968]_ ;
  assign \new_[65972]_  = ~A200 & A199;
  assign \new_[65975]_  = A203 & A201;
  assign \new_[65976]_  = \new_[65975]_  & \new_[65972]_ ;
  assign \new_[65977]_  = \new_[65976]_  & \new_[65969]_ ;
  assign \new_[65981]_  = A265 & ~A233;
  assign \new_[65982]_  = ~A232 & \new_[65981]_ ;
  assign \new_[65985]_  = A298 & A266;
  assign \new_[65988]_  = ~A302 & ~A301;
  assign \new_[65989]_  = \new_[65988]_  & \new_[65985]_ ;
  assign \new_[65990]_  = \new_[65989]_  & \new_[65982]_ ;
  assign \new_[65994]_  = ~A166 & ~A167;
  assign \new_[65995]_  = A170 & \new_[65994]_ ;
  assign \new_[65998]_  = ~A200 & A199;
  assign \new_[66001]_  = A203 & A201;
  assign \new_[66002]_  = \new_[66001]_  & \new_[65998]_ ;
  assign \new_[66003]_  = \new_[66002]_  & \new_[65995]_ ;
  assign \new_[66007]_  = ~A266 & ~A233;
  assign \new_[66008]_  = ~A232 & \new_[66007]_ ;
  assign \new_[66011]_  = ~A269 & ~A268;
  assign \new_[66014]_  = ~A300 & A298;
  assign \new_[66015]_  = \new_[66014]_  & \new_[66011]_ ;
  assign \new_[66016]_  = \new_[66015]_  & \new_[66008]_ ;
  assign \new_[66020]_  = ~A166 & ~A167;
  assign \new_[66021]_  = A170 & \new_[66020]_ ;
  assign \new_[66024]_  = ~A200 & A199;
  assign \new_[66027]_  = A203 & A201;
  assign \new_[66028]_  = \new_[66027]_  & \new_[66024]_ ;
  assign \new_[66029]_  = \new_[66028]_  & \new_[66021]_ ;
  assign \new_[66033]_  = ~A266 & ~A233;
  assign \new_[66034]_  = ~A232 & \new_[66033]_ ;
  assign \new_[66037]_  = ~A269 & ~A268;
  assign \new_[66040]_  = A299 & A298;
  assign \new_[66041]_  = \new_[66040]_  & \new_[66037]_ ;
  assign \new_[66042]_  = \new_[66041]_  & \new_[66034]_ ;
  assign \new_[66046]_  = ~A166 & ~A167;
  assign \new_[66047]_  = A170 & \new_[66046]_ ;
  assign \new_[66050]_  = ~A200 & A199;
  assign \new_[66053]_  = A203 & A201;
  assign \new_[66054]_  = \new_[66053]_  & \new_[66050]_ ;
  assign \new_[66055]_  = \new_[66054]_  & \new_[66047]_ ;
  assign \new_[66059]_  = ~A266 & ~A233;
  assign \new_[66060]_  = ~A232 & \new_[66059]_ ;
  assign \new_[66063]_  = ~A269 & ~A268;
  assign \new_[66066]_  = ~A299 & ~A298;
  assign \new_[66067]_  = \new_[66066]_  & \new_[66063]_ ;
  assign \new_[66068]_  = \new_[66067]_  & \new_[66060]_ ;
  assign \new_[66072]_  = ~A166 & ~A167;
  assign \new_[66073]_  = A170 & \new_[66072]_ ;
  assign \new_[66076]_  = ~A200 & A199;
  assign \new_[66079]_  = A203 & A201;
  assign \new_[66080]_  = \new_[66079]_  & \new_[66076]_ ;
  assign \new_[66081]_  = \new_[66080]_  & \new_[66073]_ ;
  assign \new_[66085]_  = ~A266 & ~A233;
  assign \new_[66086]_  = ~A232 & \new_[66085]_ ;
  assign \new_[66089]_  = A298 & ~A267;
  assign \new_[66092]_  = ~A302 & ~A301;
  assign \new_[66093]_  = \new_[66092]_  & \new_[66089]_ ;
  assign \new_[66094]_  = \new_[66093]_  & \new_[66086]_ ;
  assign \new_[66098]_  = ~A166 & ~A167;
  assign \new_[66099]_  = A170 & \new_[66098]_ ;
  assign \new_[66102]_  = ~A200 & A199;
  assign \new_[66105]_  = A203 & A201;
  assign \new_[66106]_  = \new_[66105]_  & \new_[66102]_ ;
  assign \new_[66107]_  = \new_[66106]_  & \new_[66099]_ ;
  assign \new_[66111]_  = ~A265 & ~A233;
  assign \new_[66112]_  = ~A232 & \new_[66111]_ ;
  assign \new_[66115]_  = A298 & ~A266;
  assign \new_[66118]_  = ~A302 & ~A301;
  assign \new_[66119]_  = \new_[66118]_  & \new_[66115]_ ;
  assign \new_[66120]_  = \new_[66119]_  & \new_[66112]_ ;
  assign \new_[66124]_  = A167 & ~A168;
  assign \new_[66125]_  = A170 & \new_[66124]_ ;
  assign \new_[66128]_  = ~A199 & A166;
  assign \new_[66131]_  = A232 & A200;
  assign \new_[66132]_  = \new_[66131]_  & \new_[66128]_ ;
  assign \new_[66133]_  = \new_[66132]_  & \new_[66125]_ ;
  assign \new_[66137]_  = ~A268 & A265;
  assign \new_[66138]_  = A233 & \new_[66137]_ ;
  assign \new_[66141]_  = ~A299 & ~A269;
  assign \new_[66144]_  = ~A302 & ~A301;
  assign \new_[66145]_  = \new_[66144]_  & \new_[66141]_ ;
  assign \new_[66146]_  = \new_[66145]_  & \new_[66138]_ ;
  assign \new_[66150]_  = A167 & ~A168;
  assign \new_[66151]_  = A170 & \new_[66150]_ ;
  assign \new_[66154]_  = ~A199 & A166;
  assign \new_[66157]_  = ~A233 & A200;
  assign \new_[66158]_  = \new_[66157]_  & \new_[66154]_ ;
  assign \new_[66159]_  = \new_[66158]_  & \new_[66151]_ ;
  assign \new_[66163]_  = A265 & ~A236;
  assign \new_[66164]_  = ~A235 & \new_[66163]_ ;
  assign \new_[66167]_  = A298 & A266;
  assign \new_[66170]_  = ~A302 & ~A301;
  assign \new_[66171]_  = \new_[66170]_  & \new_[66167]_ ;
  assign \new_[66172]_  = \new_[66171]_  & \new_[66164]_ ;
  assign \new_[66176]_  = A167 & ~A168;
  assign \new_[66177]_  = A170 & \new_[66176]_ ;
  assign \new_[66180]_  = ~A199 & A166;
  assign \new_[66183]_  = ~A233 & A200;
  assign \new_[66184]_  = \new_[66183]_  & \new_[66180]_ ;
  assign \new_[66185]_  = \new_[66184]_  & \new_[66177]_ ;
  assign \new_[66189]_  = ~A266 & ~A236;
  assign \new_[66190]_  = ~A235 & \new_[66189]_ ;
  assign \new_[66193]_  = ~A269 & ~A268;
  assign \new_[66196]_  = ~A300 & A298;
  assign \new_[66197]_  = \new_[66196]_  & \new_[66193]_ ;
  assign \new_[66198]_  = \new_[66197]_  & \new_[66190]_ ;
  assign \new_[66202]_  = A167 & ~A168;
  assign \new_[66203]_  = A170 & \new_[66202]_ ;
  assign \new_[66206]_  = ~A199 & A166;
  assign \new_[66209]_  = ~A233 & A200;
  assign \new_[66210]_  = \new_[66209]_  & \new_[66206]_ ;
  assign \new_[66211]_  = \new_[66210]_  & \new_[66203]_ ;
  assign \new_[66215]_  = ~A266 & ~A236;
  assign \new_[66216]_  = ~A235 & \new_[66215]_ ;
  assign \new_[66219]_  = ~A269 & ~A268;
  assign \new_[66222]_  = A299 & A298;
  assign \new_[66223]_  = \new_[66222]_  & \new_[66219]_ ;
  assign \new_[66224]_  = \new_[66223]_  & \new_[66216]_ ;
  assign \new_[66228]_  = A167 & ~A168;
  assign \new_[66229]_  = A170 & \new_[66228]_ ;
  assign \new_[66232]_  = ~A199 & A166;
  assign \new_[66235]_  = ~A233 & A200;
  assign \new_[66236]_  = \new_[66235]_  & \new_[66232]_ ;
  assign \new_[66237]_  = \new_[66236]_  & \new_[66229]_ ;
  assign \new_[66241]_  = ~A266 & ~A236;
  assign \new_[66242]_  = ~A235 & \new_[66241]_ ;
  assign \new_[66245]_  = ~A269 & ~A268;
  assign \new_[66248]_  = ~A299 & ~A298;
  assign \new_[66249]_  = \new_[66248]_  & \new_[66245]_ ;
  assign \new_[66250]_  = \new_[66249]_  & \new_[66242]_ ;
  assign \new_[66254]_  = A167 & ~A168;
  assign \new_[66255]_  = A170 & \new_[66254]_ ;
  assign \new_[66258]_  = ~A199 & A166;
  assign \new_[66261]_  = ~A233 & A200;
  assign \new_[66262]_  = \new_[66261]_  & \new_[66258]_ ;
  assign \new_[66263]_  = \new_[66262]_  & \new_[66255]_ ;
  assign \new_[66267]_  = ~A266 & ~A236;
  assign \new_[66268]_  = ~A235 & \new_[66267]_ ;
  assign \new_[66271]_  = A298 & ~A267;
  assign \new_[66274]_  = ~A302 & ~A301;
  assign \new_[66275]_  = \new_[66274]_  & \new_[66271]_ ;
  assign \new_[66276]_  = \new_[66275]_  & \new_[66268]_ ;
  assign \new_[66280]_  = A167 & ~A168;
  assign \new_[66281]_  = A170 & \new_[66280]_ ;
  assign \new_[66284]_  = ~A199 & A166;
  assign \new_[66287]_  = ~A233 & A200;
  assign \new_[66288]_  = \new_[66287]_  & \new_[66284]_ ;
  assign \new_[66289]_  = \new_[66288]_  & \new_[66281]_ ;
  assign \new_[66293]_  = ~A265 & ~A236;
  assign \new_[66294]_  = ~A235 & \new_[66293]_ ;
  assign \new_[66297]_  = A298 & ~A266;
  assign \new_[66300]_  = ~A302 & ~A301;
  assign \new_[66301]_  = \new_[66300]_  & \new_[66297]_ ;
  assign \new_[66302]_  = \new_[66301]_  & \new_[66294]_ ;
  assign \new_[66306]_  = A167 & ~A168;
  assign \new_[66307]_  = A170 & \new_[66306]_ ;
  assign \new_[66310]_  = ~A199 & A166;
  assign \new_[66313]_  = ~A233 & A200;
  assign \new_[66314]_  = \new_[66313]_  & \new_[66310]_ ;
  assign \new_[66315]_  = \new_[66314]_  & \new_[66307]_ ;
  assign \new_[66319]_  = ~A268 & ~A266;
  assign \new_[66320]_  = ~A234 & \new_[66319]_ ;
  assign \new_[66323]_  = A298 & ~A269;
  assign \new_[66326]_  = ~A302 & ~A301;
  assign \new_[66327]_  = \new_[66326]_  & \new_[66323]_ ;
  assign \new_[66328]_  = \new_[66327]_  & \new_[66320]_ ;
  assign \new_[66332]_  = A167 & ~A168;
  assign \new_[66333]_  = A170 & \new_[66332]_ ;
  assign \new_[66336]_  = ~A199 & A166;
  assign \new_[66339]_  = A232 & A200;
  assign \new_[66340]_  = \new_[66339]_  & \new_[66336]_ ;
  assign \new_[66341]_  = \new_[66340]_  & \new_[66333]_ ;
  assign \new_[66345]_  = A235 & A234;
  assign \new_[66346]_  = ~A233 & \new_[66345]_ ;
  assign \new_[66349]_  = ~A299 & A298;
  assign \new_[66352]_  = A301 & A300;
  assign \new_[66353]_  = \new_[66352]_  & \new_[66349]_ ;
  assign \new_[66354]_  = \new_[66353]_  & \new_[66346]_ ;
  assign \new_[66358]_  = A167 & ~A168;
  assign \new_[66359]_  = A170 & \new_[66358]_ ;
  assign \new_[66362]_  = ~A199 & A166;
  assign \new_[66365]_  = A232 & A200;
  assign \new_[66366]_  = \new_[66365]_  & \new_[66362]_ ;
  assign \new_[66367]_  = \new_[66366]_  & \new_[66359]_ ;
  assign \new_[66371]_  = A235 & A234;
  assign \new_[66372]_  = ~A233 & \new_[66371]_ ;
  assign \new_[66375]_  = ~A299 & A298;
  assign \new_[66378]_  = A302 & A300;
  assign \new_[66379]_  = \new_[66378]_  & \new_[66375]_ ;
  assign \new_[66380]_  = \new_[66379]_  & \new_[66372]_ ;
  assign \new_[66384]_  = A167 & ~A168;
  assign \new_[66385]_  = A170 & \new_[66384]_ ;
  assign \new_[66388]_  = ~A199 & A166;
  assign \new_[66391]_  = A232 & A200;
  assign \new_[66392]_  = \new_[66391]_  & \new_[66388]_ ;
  assign \new_[66393]_  = \new_[66392]_  & \new_[66385]_ ;
  assign \new_[66397]_  = A235 & A234;
  assign \new_[66398]_  = ~A233 & \new_[66397]_ ;
  assign \new_[66401]_  = ~A266 & A265;
  assign \new_[66404]_  = A268 & A267;
  assign \new_[66405]_  = \new_[66404]_  & \new_[66401]_ ;
  assign \new_[66406]_  = \new_[66405]_  & \new_[66398]_ ;
  assign \new_[66410]_  = A167 & ~A168;
  assign \new_[66411]_  = A170 & \new_[66410]_ ;
  assign \new_[66414]_  = ~A199 & A166;
  assign \new_[66417]_  = A232 & A200;
  assign \new_[66418]_  = \new_[66417]_  & \new_[66414]_ ;
  assign \new_[66419]_  = \new_[66418]_  & \new_[66411]_ ;
  assign \new_[66423]_  = A235 & A234;
  assign \new_[66424]_  = ~A233 & \new_[66423]_ ;
  assign \new_[66427]_  = ~A266 & A265;
  assign \new_[66430]_  = A269 & A267;
  assign \new_[66431]_  = \new_[66430]_  & \new_[66427]_ ;
  assign \new_[66432]_  = \new_[66431]_  & \new_[66424]_ ;
  assign \new_[66436]_  = A167 & ~A168;
  assign \new_[66437]_  = A170 & \new_[66436]_ ;
  assign \new_[66440]_  = ~A199 & A166;
  assign \new_[66443]_  = A232 & A200;
  assign \new_[66444]_  = \new_[66443]_  & \new_[66440]_ ;
  assign \new_[66445]_  = \new_[66444]_  & \new_[66437]_ ;
  assign \new_[66449]_  = A236 & A234;
  assign \new_[66450]_  = ~A233 & \new_[66449]_ ;
  assign \new_[66453]_  = ~A299 & A298;
  assign \new_[66456]_  = A301 & A300;
  assign \new_[66457]_  = \new_[66456]_  & \new_[66453]_ ;
  assign \new_[66458]_  = \new_[66457]_  & \new_[66450]_ ;
  assign \new_[66462]_  = A167 & ~A168;
  assign \new_[66463]_  = A170 & \new_[66462]_ ;
  assign \new_[66466]_  = ~A199 & A166;
  assign \new_[66469]_  = A232 & A200;
  assign \new_[66470]_  = \new_[66469]_  & \new_[66466]_ ;
  assign \new_[66471]_  = \new_[66470]_  & \new_[66463]_ ;
  assign \new_[66475]_  = A236 & A234;
  assign \new_[66476]_  = ~A233 & \new_[66475]_ ;
  assign \new_[66479]_  = ~A299 & A298;
  assign \new_[66482]_  = A302 & A300;
  assign \new_[66483]_  = \new_[66482]_  & \new_[66479]_ ;
  assign \new_[66484]_  = \new_[66483]_  & \new_[66476]_ ;
  assign \new_[66488]_  = A167 & ~A168;
  assign \new_[66489]_  = A170 & \new_[66488]_ ;
  assign \new_[66492]_  = ~A199 & A166;
  assign \new_[66495]_  = A232 & A200;
  assign \new_[66496]_  = \new_[66495]_  & \new_[66492]_ ;
  assign \new_[66497]_  = \new_[66496]_  & \new_[66489]_ ;
  assign \new_[66501]_  = A236 & A234;
  assign \new_[66502]_  = ~A233 & \new_[66501]_ ;
  assign \new_[66505]_  = ~A266 & A265;
  assign \new_[66508]_  = A268 & A267;
  assign \new_[66509]_  = \new_[66508]_  & \new_[66505]_ ;
  assign \new_[66510]_  = \new_[66509]_  & \new_[66502]_ ;
  assign \new_[66514]_  = A167 & ~A168;
  assign \new_[66515]_  = A170 & \new_[66514]_ ;
  assign \new_[66518]_  = ~A199 & A166;
  assign \new_[66521]_  = A232 & A200;
  assign \new_[66522]_  = \new_[66521]_  & \new_[66518]_ ;
  assign \new_[66523]_  = \new_[66522]_  & \new_[66515]_ ;
  assign \new_[66527]_  = A236 & A234;
  assign \new_[66528]_  = ~A233 & \new_[66527]_ ;
  assign \new_[66531]_  = ~A266 & A265;
  assign \new_[66534]_  = A269 & A267;
  assign \new_[66535]_  = \new_[66534]_  & \new_[66531]_ ;
  assign \new_[66536]_  = \new_[66535]_  & \new_[66528]_ ;
  assign \new_[66540]_  = A167 & ~A168;
  assign \new_[66541]_  = A170 & \new_[66540]_ ;
  assign \new_[66544]_  = ~A199 & A166;
  assign \new_[66547]_  = ~A232 & A200;
  assign \new_[66548]_  = \new_[66547]_  & \new_[66544]_ ;
  assign \new_[66549]_  = \new_[66548]_  & \new_[66541]_ ;
  assign \new_[66553]_  = ~A268 & ~A266;
  assign \new_[66554]_  = ~A233 & \new_[66553]_ ;
  assign \new_[66557]_  = A298 & ~A269;
  assign \new_[66560]_  = ~A302 & ~A301;
  assign \new_[66561]_  = \new_[66560]_  & \new_[66557]_ ;
  assign \new_[66562]_  = \new_[66561]_  & \new_[66554]_ ;
  assign \new_[66566]_  = A167 & ~A168;
  assign \new_[66567]_  = ~A170 & \new_[66566]_ ;
  assign \new_[66570]_  = ~A199 & ~A166;
  assign \new_[66573]_  = A232 & A200;
  assign \new_[66574]_  = \new_[66573]_  & \new_[66570]_ ;
  assign \new_[66575]_  = \new_[66574]_  & \new_[66567]_ ;
  assign \new_[66579]_  = ~A268 & A265;
  assign \new_[66580]_  = A233 & \new_[66579]_ ;
  assign \new_[66583]_  = ~A299 & ~A269;
  assign \new_[66586]_  = ~A302 & ~A301;
  assign \new_[66587]_  = \new_[66586]_  & \new_[66583]_ ;
  assign \new_[66588]_  = \new_[66587]_  & \new_[66580]_ ;
  assign \new_[66592]_  = A167 & ~A168;
  assign \new_[66593]_  = ~A170 & \new_[66592]_ ;
  assign \new_[66596]_  = ~A199 & ~A166;
  assign \new_[66599]_  = ~A233 & A200;
  assign \new_[66600]_  = \new_[66599]_  & \new_[66596]_ ;
  assign \new_[66601]_  = \new_[66600]_  & \new_[66593]_ ;
  assign \new_[66605]_  = A265 & ~A236;
  assign \new_[66606]_  = ~A235 & \new_[66605]_ ;
  assign \new_[66609]_  = A298 & A266;
  assign \new_[66612]_  = ~A302 & ~A301;
  assign \new_[66613]_  = \new_[66612]_  & \new_[66609]_ ;
  assign \new_[66614]_  = \new_[66613]_  & \new_[66606]_ ;
  assign \new_[66618]_  = A167 & ~A168;
  assign \new_[66619]_  = ~A170 & \new_[66618]_ ;
  assign \new_[66622]_  = ~A199 & ~A166;
  assign \new_[66625]_  = ~A233 & A200;
  assign \new_[66626]_  = \new_[66625]_  & \new_[66622]_ ;
  assign \new_[66627]_  = \new_[66626]_  & \new_[66619]_ ;
  assign \new_[66631]_  = ~A266 & ~A236;
  assign \new_[66632]_  = ~A235 & \new_[66631]_ ;
  assign \new_[66635]_  = ~A269 & ~A268;
  assign \new_[66638]_  = ~A300 & A298;
  assign \new_[66639]_  = \new_[66638]_  & \new_[66635]_ ;
  assign \new_[66640]_  = \new_[66639]_  & \new_[66632]_ ;
  assign \new_[66644]_  = A167 & ~A168;
  assign \new_[66645]_  = ~A170 & \new_[66644]_ ;
  assign \new_[66648]_  = ~A199 & ~A166;
  assign \new_[66651]_  = ~A233 & A200;
  assign \new_[66652]_  = \new_[66651]_  & \new_[66648]_ ;
  assign \new_[66653]_  = \new_[66652]_  & \new_[66645]_ ;
  assign \new_[66657]_  = ~A266 & ~A236;
  assign \new_[66658]_  = ~A235 & \new_[66657]_ ;
  assign \new_[66661]_  = ~A269 & ~A268;
  assign \new_[66664]_  = A299 & A298;
  assign \new_[66665]_  = \new_[66664]_  & \new_[66661]_ ;
  assign \new_[66666]_  = \new_[66665]_  & \new_[66658]_ ;
  assign \new_[66670]_  = A167 & ~A168;
  assign \new_[66671]_  = ~A170 & \new_[66670]_ ;
  assign \new_[66674]_  = ~A199 & ~A166;
  assign \new_[66677]_  = ~A233 & A200;
  assign \new_[66678]_  = \new_[66677]_  & \new_[66674]_ ;
  assign \new_[66679]_  = \new_[66678]_  & \new_[66671]_ ;
  assign \new_[66683]_  = ~A266 & ~A236;
  assign \new_[66684]_  = ~A235 & \new_[66683]_ ;
  assign \new_[66687]_  = ~A269 & ~A268;
  assign \new_[66690]_  = ~A299 & ~A298;
  assign \new_[66691]_  = \new_[66690]_  & \new_[66687]_ ;
  assign \new_[66692]_  = \new_[66691]_  & \new_[66684]_ ;
  assign \new_[66696]_  = A167 & ~A168;
  assign \new_[66697]_  = ~A170 & \new_[66696]_ ;
  assign \new_[66700]_  = ~A199 & ~A166;
  assign \new_[66703]_  = ~A233 & A200;
  assign \new_[66704]_  = \new_[66703]_  & \new_[66700]_ ;
  assign \new_[66705]_  = \new_[66704]_  & \new_[66697]_ ;
  assign \new_[66709]_  = ~A266 & ~A236;
  assign \new_[66710]_  = ~A235 & \new_[66709]_ ;
  assign \new_[66713]_  = A298 & ~A267;
  assign \new_[66716]_  = ~A302 & ~A301;
  assign \new_[66717]_  = \new_[66716]_  & \new_[66713]_ ;
  assign \new_[66718]_  = \new_[66717]_  & \new_[66710]_ ;
  assign \new_[66722]_  = A167 & ~A168;
  assign \new_[66723]_  = ~A170 & \new_[66722]_ ;
  assign \new_[66726]_  = ~A199 & ~A166;
  assign \new_[66729]_  = ~A233 & A200;
  assign \new_[66730]_  = \new_[66729]_  & \new_[66726]_ ;
  assign \new_[66731]_  = \new_[66730]_  & \new_[66723]_ ;
  assign \new_[66735]_  = ~A265 & ~A236;
  assign \new_[66736]_  = ~A235 & \new_[66735]_ ;
  assign \new_[66739]_  = A298 & ~A266;
  assign \new_[66742]_  = ~A302 & ~A301;
  assign \new_[66743]_  = \new_[66742]_  & \new_[66739]_ ;
  assign \new_[66744]_  = \new_[66743]_  & \new_[66736]_ ;
  assign \new_[66748]_  = A167 & ~A168;
  assign \new_[66749]_  = ~A170 & \new_[66748]_ ;
  assign \new_[66752]_  = ~A199 & ~A166;
  assign \new_[66755]_  = ~A233 & A200;
  assign \new_[66756]_  = \new_[66755]_  & \new_[66752]_ ;
  assign \new_[66757]_  = \new_[66756]_  & \new_[66749]_ ;
  assign \new_[66761]_  = ~A268 & ~A266;
  assign \new_[66762]_  = ~A234 & \new_[66761]_ ;
  assign \new_[66765]_  = A298 & ~A269;
  assign \new_[66768]_  = ~A302 & ~A301;
  assign \new_[66769]_  = \new_[66768]_  & \new_[66765]_ ;
  assign \new_[66770]_  = \new_[66769]_  & \new_[66762]_ ;
  assign \new_[66774]_  = A167 & ~A168;
  assign \new_[66775]_  = ~A170 & \new_[66774]_ ;
  assign \new_[66778]_  = ~A199 & ~A166;
  assign \new_[66781]_  = A232 & A200;
  assign \new_[66782]_  = \new_[66781]_  & \new_[66778]_ ;
  assign \new_[66783]_  = \new_[66782]_  & \new_[66775]_ ;
  assign \new_[66787]_  = A235 & A234;
  assign \new_[66788]_  = ~A233 & \new_[66787]_ ;
  assign \new_[66791]_  = ~A299 & A298;
  assign \new_[66794]_  = A301 & A300;
  assign \new_[66795]_  = \new_[66794]_  & \new_[66791]_ ;
  assign \new_[66796]_  = \new_[66795]_  & \new_[66788]_ ;
  assign \new_[66800]_  = A167 & ~A168;
  assign \new_[66801]_  = ~A170 & \new_[66800]_ ;
  assign \new_[66804]_  = ~A199 & ~A166;
  assign \new_[66807]_  = A232 & A200;
  assign \new_[66808]_  = \new_[66807]_  & \new_[66804]_ ;
  assign \new_[66809]_  = \new_[66808]_  & \new_[66801]_ ;
  assign \new_[66813]_  = A235 & A234;
  assign \new_[66814]_  = ~A233 & \new_[66813]_ ;
  assign \new_[66817]_  = ~A299 & A298;
  assign \new_[66820]_  = A302 & A300;
  assign \new_[66821]_  = \new_[66820]_  & \new_[66817]_ ;
  assign \new_[66822]_  = \new_[66821]_  & \new_[66814]_ ;
  assign \new_[66826]_  = A167 & ~A168;
  assign \new_[66827]_  = ~A170 & \new_[66826]_ ;
  assign \new_[66830]_  = ~A199 & ~A166;
  assign \new_[66833]_  = A232 & A200;
  assign \new_[66834]_  = \new_[66833]_  & \new_[66830]_ ;
  assign \new_[66835]_  = \new_[66834]_  & \new_[66827]_ ;
  assign \new_[66839]_  = A235 & A234;
  assign \new_[66840]_  = ~A233 & \new_[66839]_ ;
  assign \new_[66843]_  = ~A266 & A265;
  assign \new_[66846]_  = A268 & A267;
  assign \new_[66847]_  = \new_[66846]_  & \new_[66843]_ ;
  assign \new_[66848]_  = \new_[66847]_  & \new_[66840]_ ;
  assign \new_[66852]_  = A167 & ~A168;
  assign \new_[66853]_  = ~A170 & \new_[66852]_ ;
  assign \new_[66856]_  = ~A199 & ~A166;
  assign \new_[66859]_  = A232 & A200;
  assign \new_[66860]_  = \new_[66859]_  & \new_[66856]_ ;
  assign \new_[66861]_  = \new_[66860]_  & \new_[66853]_ ;
  assign \new_[66865]_  = A235 & A234;
  assign \new_[66866]_  = ~A233 & \new_[66865]_ ;
  assign \new_[66869]_  = ~A266 & A265;
  assign \new_[66872]_  = A269 & A267;
  assign \new_[66873]_  = \new_[66872]_  & \new_[66869]_ ;
  assign \new_[66874]_  = \new_[66873]_  & \new_[66866]_ ;
  assign \new_[66878]_  = A167 & ~A168;
  assign \new_[66879]_  = ~A170 & \new_[66878]_ ;
  assign \new_[66882]_  = ~A199 & ~A166;
  assign \new_[66885]_  = A232 & A200;
  assign \new_[66886]_  = \new_[66885]_  & \new_[66882]_ ;
  assign \new_[66887]_  = \new_[66886]_  & \new_[66879]_ ;
  assign \new_[66891]_  = A236 & A234;
  assign \new_[66892]_  = ~A233 & \new_[66891]_ ;
  assign \new_[66895]_  = ~A299 & A298;
  assign \new_[66898]_  = A301 & A300;
  assign \new_[66899]_  = \new_[66898]_  & \new_[66895]_ ;
  assign \new_[66900]_  = \new_[66899]_  & \new_[66892]_ ;
  assign \new_[66904]_  = A167 & ~A168;
  assign \new_[66905]_  = ~A170 & \new_[66904]_ ;
  assign \new_[66908]_  = ~A199 & ~A166;
  assign \new_[66911]_  = A232 & A200;
  assign \new_[66912]_  = \new_[66911]_  & \new_[66908]_ ;
  assign \new_[66913]_  = \new_[66912]_  & \new_[66905]_ ;
  assign \new_[66917]_  = A236 & A234;
  assign \new_[66918]_  = ~A233 & \new_[66917]_ ;
  assign \new_[66921]_  = ~A299 & A298;
  assign \new_[66924]_  = A302 & A300;
  assign \new_[66925]_  = \new_[66924]_  & \new_[66921]_ ;
  assign \new_[66926]_  = \new_[66925]_  & \new_[66918]_ ;
  assign \new_[66930]_  = A167 & ~A168;
  assign \new_[66931]_  = ~A170 & \new_[66930]_ ;
  assign \new_[66934]_  = ~A199 & ~A166;
  assign \new_[66937]_  = A232 & A200;
  assign \new_[66938]_  = \new_[66937]_  & \new_[66934]_ ;
  assign \new_[66939]_  = \new_[66938]_  & \new_[66931]_ ;
  assign \new_[66943]_  = A236 & A234;
  assign \new_[66944]_  = ~A233 & \new_[66943]_ ;
  assign \new_[66947]_  = ~A266 & A265;
  assign \new_[66950]_  = A268 & A267;
  assign \new_[66951]_  = \new_[66950]_  & \new_[66947]_ ;
  assign \new_[66952]_  = \new_[66951]_  & \new_[66944]_ ;
  assign \new_[66956]_  = A167 & ~A168;
  assign \new_[66957]_  = ~A170 & \new_[66956]_ ;
  assign \new_[66960]_  = ~A199 & ~A166;
  assign \new_[66963]_  = A232 & A200;
  assign \new_[66964]_  = \new_[66963]_  & \new_[66960]_ ;
  assign \new_[66965]_  = \new_[66964]_  & \new_[66957]_ ;
  assign \new_[66969]_  = A236 & A234;
  assign \new_[66970]_  = ~A233 & \new_[66969]_ ;
  assign \new_[66973]_  = ~A266 & A265;
  assign \new_[66976]_  = A269 & A267;
  assign \new_[66977]_  = \new_[66976]_  & \new_[66973]_ ;
  assign \new_[66978]_  = \new_[66977]_  & \new_[66970]_ ;
  assign \new_[66982]_  = A167 & ~A168;
  assign \new_[66983]_  = ~A170 & \new_[66982]_ ;
  assign \new_[66986]_  = ~A199 & ~A166;
  assign \new_[66989]_  = ~A232 & A200;
  assign \new_[66990]_  = \new_[66989]_  & \new_[66986]_ ;
  assign \new_[66991]_  = \new_[66990]_  & \new_[66983]_ ;
  assign \new_[66995]_  = ~A268 & ~A266;
  assign \new_[66996]_  = ~A233 & \new_[66995]_ ;
  assign \new_[66999]_  = A298 & ~A269;
  assign \new_[67002]_  = ~A302 & ~A301;
  assign \new_[67003]_  = \new_[67002]_  & \new_[66999]_ ;
  assign \new_[67004]_  = \new_[67003]_  & \new_[66996]_ ;
  assign \new_[67008]_  = ~A167 & ~A168;
  assign \new_[67009]_  = ~A170 & \new_[67008]_ ;
  assign \new_[67012]_  = ~A199 & A166;
  assign \new_[67015]_  = A232 & A200;
  assign \new_[67016]_  = \new_[67015]_  & \new_[67012]_ ;
  assign \new_[67017]_  = \new_[67016]_  & \new_[67009]_ ;
  assign \new_[67021]_  = ~A268 & A265;
  assign \new_[67022]_  = A233 & \new_[67021]_ ;
  assign \new_[67025]_  = ~A299 & ~A269;
  assign \new_[67028]_  = ~A302 & ~A301;
  assign \new_[67029]_  = \new_[67028]_  & \new_[67025]_ ;
  assign \new_[67030]_  = \new_[67029]_  & \new_[67022]_ ;
  assign \new_[67034]_  = ~A167 & ~A168;
  assign \new_[67035]_  = ~A170 & \new_[67034]_ ;
  assign \new_[67038]_  = ~A199 & A166;
  assign \new_[67041]_  = ~A233 & A200;
  assign \new_[67042]_  = \new_[67041]_  & \new_[67038]_ ;
  assign \new_[67043]_  = \new_[67042]_  & \new_[67035]_ ;
  assign \new_[67047]_  = A265 & ~A236;
  assign \new_[67048]_  = ~A235 & \new_[67047]_ ;
  assign \new_[67051]_  = A298 & A266;
  assign \new_[67054]_  = ~A302 & ~A301;
  assign \new_[67055]_  = \new_[67054]_  & \new_[67051]_ ;
  assign \new_[67056]_  = \new_[67055]_  & \new_[67048]_ ;
  assign \new_[67060]_  = ~A167 & ~A168;
  assign \new_[67061]_  = ~A170 & \new_[67060]_ ;
  assign \new_[67064]_  = ~A199 & A166;
  assign \new_[67067]_  = ~A233 & A200;
  assign \new_[67068]_  = \new_[67067]_  & \new_[67064]_ ;
  assign \new_[67069]_  = \new_[67068]_  & \new_[67061]_ ;
  assign \new_[67073]_  = ~A266 & ~A236;
  assign \new_[67074]_  = ~A235 & \new_[67073]_ ;
  assign \new_[67077]_  = ~A269 & ~A268;
  assign \new_[67080]_  = ~A300 & A298;
  assign \new_[67081]_  = \new_[67080]_  & \new_[67077]_ ;
  assign \new_[67082]_  = \new_[67081]_  & \new_[67074]_ ;
  assign \new_[67086]_  = ~A167 & ~A168;
  assign \new_[67087]_  = ~A170 & \new_[67086]_ ;
  assign \new_[67090]_  = ~A199 & A166;
  assign \new_[67093]_  = ~A233 & A200;
  assign \new_[67094]_  = \new_[67093]_  & \new_[67090]_ ;
  assign \new_[67095]_  = \new_[67094]_  & \new_[67087]_ ;
  assign \new_[67099]_  = ~A266 & ~A236;
  assign \new_[67100]_  = ~A235 & \new_[67099]_ ;
  assign \new_[67103]_  = ~A269 & ~A268;
  assign \new_[67106]_  = A299 & A298;
  assign \new_[67107]_  = \new_[67106]_  & \new_[67103]_ ;
  assign \new_[67108]_  = \new_[67107]_  & \new_[67100]_ ;
  assign \new_[67112]_  = ~A167 & ~A168;
  assign \new_[67113]_  = ~A170 & \new_[67112]_ ;
  assign \new_[67116]_  = ~A199 & A166;
  assign \new_[67119]_  = ~A233 & A200;
  assign \new_[67120]_  = \new_[67119]_  & \new_[67116]_ ;
  assign \new_[67121]_  = \new_[67120]_  & \new_[67113]_ ;
  assign \new_[67125]_  = ~A266 & ~A236;
  assign \new_[67126]_  = ~A235 & \new_[67125]_ ;
  assign \new_[67129]_  = ~A269 & ~A268;
  assign \new_[67132]_  = ~A299 & ~A298;
  assign \new_[67133]_  = \new_[67132]_  & \new_[67129]_ ;
  assign \new_[67134]_  = \new_[67133]_  & \new_[67126]_ ;
  assign \new_[67138]_  = ~A167 & ~A168;
  assign \new_[67139]_  = ~A170 & \new_[67138]_ ;
  assign \new_[67142]_  = ~A199 & A166;
  assign \new_[67145]_  = ~A233 & A200;
  assign \new_[67146]_  = \new_[67145]_  & \new_[67142]_ ;
  assign \new_[67147]_  = \new_[67146]_  & \new_[67139]_ ;
  assign \new_[67151]_  = ~A266 & ~A236;
  assign \new_[67152]_  = ~A235 & \new_[67151]_ ;
  assign \new_[67155]_  = A298 & ~A267;
  assign \new_[67158]_  = ~A302 & ~A301;
  assign \new_[67159]_  = \new_[67158]_  & \new_[67155]_ ;
  assign \new_[67160]_  = \new_[67159]_  & \new_[67152]_ ;
  assign \new_[67164]_  = ~A167 & ~A168;
  assign \new_[67165]_  = ~A170 & \new_[67164]_ ;
  assign \new_[67168]_  = ~A199 & A166;
  assign \new_[67171]_  = ~A233 & A200;
  assign \new_[67172]_  = \new_[67171]_  & \new_[67168]_ ;
  assign \new_[67173]_  = \new_[67172]_  & \new_[67165]_ ;
  assign \new_[67177]_  = ~A265 & ~A236;
  assign \new_[67178]_  = ~A235 & \new_[67177]_ ;
  assign \new_[67181]_  = A298 & ~A266;
  assign \new_[67184]_  = ~A302 & ~A301;
  assign \new_[67185]_  = \new_[67184]_  & \new_[67181]_ ;
  assign \new_[67186]_  = \new_[67185]_  & \new_[67178]_ ;
  assign \new_[67190]_  = ~A167 & ~A168;
  assign \new_[67191]_  = ~A170 & \new_[67190]_ ;
  assign \new_[67194]_  = ~A199 & A166;
  assign \new_[67197]_  = ~A233 & A200;
  assign \new_[67198]_  = \new_[67197]_  & \new_[67194]_ ;
  assign \new_[67199]_  = \new_[67198]_  & \new_[67191]_ ;
  assign \new_[67203]_  = ~A268 & ~A266;
  assign \new_[67204]_  = ~A234 & \new_[67203]_ ;
  assign \new_[67207]_  = A298 & ~A269;
  assign \new_[67210]_  = ~A302 & ~A301;
  assign \new_[67211]_  = \new_[67210]_  & \new_[67207]_ ;
  assign \new_[67212]_  = \new_[67211]_  & \new_[67204]_ ;
  assign \new_[67216]_  = ~A167 & ~A168;
  assign \new_[67217]_  = ~A170 & \new_[67216]_ ;
  assign \new_[67220]_  = ~A199 & A166;
  assign \new_[67223]_  = A232 & A200;
  assign \new_[67224]_  = \new_[67223]_  & \new_[67220]_ ;
  assign \new_[67225]_  = \new_[67224]_  & \new_[67217]_ ;
  assign \new_[67229]_  = A235 & A234;
  assign \new_[67230]_  = ~A233 & \new_[67229]_ ;
  assign \new_[67233]_  = ~A299 & A298;
  assign \new_[67236]_  = A301 & A300;
  assign \new_[67237]_  = \new_[67236]_  & \new_[67233]_ ;
  assign \new_[67238]_  = \new_[67237]_  & \new_[67230]_ ;
  assign \new_[67242]_  = ~A167 & ~A168;
  assign \new_[67243]_  = ~A170 & \new_[67242]_ ;
  assign \new_[67246]_  = ~A199 & A166;
  assign \new_[67249]_  = A232 & A200;
  assign \new_[67250]_  = \new_[67249]_  & \new_[67246]_ ;
  assign \new_[67251]_  = \new_[67250]_  & \new_[67243]_ ;
  assign \new_[67255]_  = A235 & A234;
  assign \new_[67256]_  = ~A233 & \new_[67255]_ ;
  assign \new_[67259]_  = ~A299 & A298;
  assign \new_[67262]_  = A302 & A300;
  assign \new_[67263]_  = \new_[67262]_  & \new_[67259]_ ;
  assign \new_[67264]_  = \new_[67263]_  & \new_[67256]_ ;
  assign \new_[67268]_  = ~A167 & ~A168;
  assign \new_[67269]_  = ~A170 & \new_[67268]_ ;
  assign \new_[67272]_  = ~A199 & A166;
  assign \new_[67275]_  = A232 & A200;
  assign \new_[67276]_  = \new_[67275]_  & \new_[67272]_ ;
  assign \new_[67277]_  = \new_[67276]_  & \new_[67269]_ ;
  assign \new_[67281]_  = A235 & A234;
  assign \new_[67282]_  = ~A233 & \new_[67281]_ ;
  assign \new_[67285]_  = ~A266 & A265;
  assign \new_[67288]_  = A268 & A267;
  assign \new_[67289]_  = \new_[67288]_  & \new_[67285]_ ;
  assign \new_[67290]_  = \new_[67289]_  & \new_[67282]_ ;
  assign \new_[67294]_  = ~A167 & ~A168;
  assign \new_[67295]_  = ~A170 & \new_[67294]_ ;
  assign \new_[67298]_  = ~A199 & A166;
  assign \new_[67301]_  = A232 & A200;
  assign \new_[67302]_  = \new_[67301]_  & \new_[67298]_ ;
  assign \new_[67303]_  = \new_[67302]_  & \new_[67295]_ ;
  assign \new_[67307]_  = A235 & A234;
  assign \new_[67308]_  = ~A233 & \new_[67307]_ ;
  assign \new_[67311]_  = ~A266 & A265;
  assign \new_[67314]_  = A269 & A267;
  assign \new_[67315]_  = \new_[67314]_  & \new_[67311]_ ;
  assign \new_[67316]_  = \new_[67315]_  & \new_[67308]_ ;
  assign \new_[67320]_  = ~A167 & ~A168;
  assign \new_[67321]_  = ~A170 & \new_[67320]_ ;
  assign \new_[67324]_  = ~A199 & A166;
  assign \new_[67327]_  = A232 & A200;
  assign \new_[67328]_  = \new_[67327]_  & \new_[67324]_ ;
  assign \new_[67329]_  = \new_[67328]_  & \new_[67321]_ ;
  assign \new_[67333]_  = A236 & A234;
  assign \new_[67334]_  = ~A233 & \new_[67333]_ ;
  assign \new_[67337]_  = ~A299 & A298;
  assign \new_[67340]_  = A301 & A300;
  assign \new_[67341]_  = \new_[67340]_  & \new_[67337]_ ;
  assign \new_[67342]_  = \new_[67341]_  & \new_[67334]_ ;
  assign \new_[67346]_  = ~A167 & ~A168;
  assign \new_[67347]_  = ~A170 & \new_[67346]_ ;
  assign \new_[67350]_  = ~A199 & A166;
  assign \new_[67353]_  = A232 & A200;
  assign \new_[67354]_  = \new_[67353]_  & \new_[67350]_ ;
  assign \new_[67355]_  = \new_[67354]_  & \new_[67347]_ ;
  assign \new_[67359]_  = A236 & A234;
  assign \new_[67360]_  = ~A233 & \new_[67359]_ ;
  assign \new_[67363]_  = ~A299 & A298;
  assign \new_[67366]_  = A302 & A300;
  assign \new_[67367]_  = \new_[67366]_  & \new_[67363]_ ;
  assign \new_[67368]_  = \new_[67367]_  & \new_[67360]_ ;
  assign \new_[67372]_  = ~A167 & ~A168;
  assign \new_[67373]_  = ~A170 & \new_[67372]_ ;
  assign \new_[67376]_  = ~A199 & A166;
  assign \new_[67379]_  = A232 & A200;
  assign \new_[67380]_  = \new_[67379]_  & \new_[67376]_ ;
  assign \new_[67381]_  = \new_[67380]_  & \new_[67373]_ ;
  assign \new_[67385]_  = A236 & A234;
  assign \new_[67386]_  = ~A233 & \new_[67385]_ ;
  assign \new_[67389]_  = ~A266 & A265;
  assign \new_[67392]_  = A268 & A267;
  assign \new_[67393]_  = \new_[67392]_  & \new_[67389]_ ;
  assign \new_[67394]_  = \new_[67393]_  & \new_[67386]_ ;
  assign \new_[67398]_  = ~A167 & ~A168;
  assign \new_[67399]_  = ~A170 & \new_[67398]_ ;
  assign \new_[67402]_  = ~A199 & A166;
  assign \new_[67405]_  = A232 & A200;
  assign \new_[67406]_  = \new_[67405]_  & \new_[67402]_ ;
  assign \new_[67407]_  = \new_[67406]_  & \new_[67399]_ ;
  assign \new_[67411]_  = A236 & A234;
  assign \new_[67412]_  = ~A233 & \new_[67411]_ ;
  assign \new_[67415]_  = ~A266 & A265;
  assign \new_[67418]_  = A269 & A267;
  assign \new_[67419]_  = \new_[67418]_  & \new_[67415]_ ;
  assign \new_[67420]_  = \new_[67419]_  & \new_[67412]_ ;
  assign \new_[67424]_  = ~A167 & ~A168;
  assign \new_[67425]_  = ~A170 & \new_[67424]_ ;
  assign \new_[67428]_  = ~A199 & A166;
  assign \new_[67431]_  = ~A232 & A200;
  assign \new_[67432]_  = \new_[67431]_  & \new_[67428]_ ;
  assign \new_[67433]_  = \new_[67432]_  & \new_[67425]_ ;
  assign \new_[67437]_  = ~A268 & ~A266;
  assign \new_[67438]_  = ~A233 & \new_[67437]_ ;
  assign \new_[67441]_  = A298 & ~A269;
  assign \new_[67444]_  = ~A302 & ~A301;
  assign \new_[67445]_  = \new_[67444]_  & \new_[67441]_ ;
  assign \new_[67446]_  = \new_[67445]_  & \new_[67438]_ ;
  assign \new_[67450]_  = A167 & ~A168;
  assign \new_[67451]_  = A169 & \new_[67450]_ ;
  assign \new_[67454]_  = ~A199 & ~A166;
  assign \new_[67457]_  = A232 & A200;
  assign \new_[67458]_  = \new_[67457]_  & \new_[67454]_ ;
  assign \new_[67459]_  = \new_[67458]_  & \new_[67451]_ ;
  assign \new_[67463]_  = ~A268 & A265;
  assign \new_[67464]_  = A233 & \new_[67463]_ ;
  assign \new_[67467]_  = ~A299 & ~A269;
  assign \new_[67470]_  = ~A302 & ~A301;
  assign \new_[67471]_  = \new_[67470]_  & \new_[67467]_ ;
  assign \new_[67472]_  = \new_[67471]_  & \new_[67464]_ ;
  assign \new_[67476]_  = A167 & ~A168;
  assign \new_[67477]_  = A169 & \new_[67476]_ ;
  assign \new_[67480]_  = ~A199 & ~A166;
  assign \new_[67483]_  = ~A233 & A200;
  assign \new_[67484]_  = \new_[67483]_  & \new_[67480]_ ;
  assign \new_[67485]_  = \new_[67484]_  & \new_[67477]_ ;
  assign \new_[67489]_  = A265 & ~A236;
  assign \new_[67490]_  = ~A235 & \new_[67489]_ ;
  assign \new_[67493]_  = A298 & A266;
  assign \new_[67496]_  = ~A302 & ~A301;
  assign \new_[67497]_  = \new_[67496]_  & \new_[67493]_ ;
  assign \new_[67498]_  = \new_[67497]_  & \new_[67490]_ ;
  assign \new_[67502]_  = A167 & ~A168;
  assign \new_[67503]_  = A169 & \new_[67502]_ ;
  assign \new_[67506]_  = ~A199 & ~A166;
  assign \new_[67509]_  = ~A233 & A200;
  assign \new_[67510]_  = \new_[67509]_  & \new_[67506]_ ;
  assign \new_[67511]_  = \new_[67510]_  & \new_[67503]_ ;
  assign \new_[67515]_  = ~A266 & ~A236;
  assign \new_[67516]_  = ~A235 & \new_[67515]_ ;
  assign \new_[67519]_  = ~A269 & ~A268;
  assign \new_[67522]_  = ~A300 & A298;
  assign \new_[67523]_  = \new_[67522]_  & \new_[67519]_ ;
  assign \new_[67524]_  = \new_[67523]_  & \new_[67516]_ ;
  assign \new_[67528]_  = A167 & ~A168;
  assign \new_[67529]_  = A169 & \new_[67528]_ ;
  assign \new_[67532]_  = ~A199 & ~A166;
  assign \new_[67535]_  = ~A233 & A200;
  assign \new_[67536]_  = \new_[67535]_  & \new_[67532]_ ;
  assign \new_[67537]_  = \new_[67536]_  & \new_[67529]_ ;
  assign \new_[67541]_  = ~A266 & ~A236;
  assign \new_[67542]_  = ~A235 & \new_[67541]_ ;
  assign \new_[67545]_  = ~A269 & ~A268;
  assign \new_[67548]_  = A299 & A298;
  assign \new_[67549]_  = \new_[67548]_  & \new_[67545]_ ;
  assign \new_[67550]_  = \new_[67549]_  & \new_[67542]_ ;
  assign \new_[67554]_  = A167 & ~A168;
  assign \new_[67555]_  = A169 & \new_[67554]_ ;
  assign \new_[67558]_  = ~A199 & ~A166;
  assign \new_[67561]_  = ~A233 & A200;
  assign \new_[67562]_  = \new_[67561]_  & \new_[67558]_ ;
  assign \new_[67563]_  = \new_[67562]_  & \new_[67555]_ ;
  assign \new_[67567]_  = ~A266 & ~A236;
  assign \new_[67568]_  = ~A235 & \new_[67567]_ ;
  assign \new_[67571]_  = ~A269 & ~A268;
  assign \new_[67574]_  = ~A299 & ~A298;
  assign \new_[67575]_  = \new_[67574]_  & \new_[67571]_ ;
  assign \new_[67576]_  = \new_[67575]_  & \new_[67568]_ ;
  assign \new_[67580]_  = A167 & ~A168;
  assign \new_[67581]_  = A169 & \new_[67580]_ ;
  assign \new_[67584]_  = ~A199 & ~A166;
  assign \new_[67587]_  = ~A233 & A200;
  assign \new_[67588]_  = \new_[67587]_  & \new_[67584]_ ;
  assign \new_[67589]_  = \new_[67588]_  & \new_[67581]_ ;
  assign \new_[67593]_  = ~A266 & ~A236;
  assign \new_[67594]_  = ~A235 & \new_[67593]_ ;
  assign \new_[67597]_  = A298 & ~A267;
  assign \new_[67600]_  = ~A302 & ~A301;
  assign \new_[67601]_  = \new_[67600]_  & \new_[67597]_ ;
  assign \new_[67602]_  = \new_[67601]_  & \new_[67594]_ ;
  assign \new_[67606]_  = A167 & ~A168;
  assign \new_[67607]_  = A169 & \new_[67606]_ ;
  assign \new_[67610]_  = ~A199 & ~A166;
  assign \new_[67613]_  = ~A233 & A200;
  assign \new_[67614]_  = \new_[67613]_  & \new_[67610]_ ;
  assign \new_[67615]_  = \new_[67614]_  & \new_[67607]_ ;
  assign \new_[67619]_  = ~A265 & ~A236;
  assign \new_[67620]_  = ~A235 & \new_[67619]_ ;
  assign \new_[67623]_  = A298 & ~A266;
  assign \new_[67626]_  = ~A302 & ~A301;
  assign \new_[67627]_  = \new_[67626]_  & \new_[67623]_ ;
  assign \new_[67628]_  = \new_[67627]_  & \new_[67620]_ ;
  assign \new_[67632]_  = A167 & ~A168;
  assign \new_[67633]_  = A169 & \new_[67632]_ ;
  assign \new_[67636]_  = ~A199 & ~A166;
  assign \new_[67639]_  = ~A233 & A200;
  assign \new_[67640]_  = \new_[67639]_  & \new_[67636]_ ;
  assign \new_[67641]_  = \new_[67640]_  & \new_[67633]_ ;
  assign \new_[67645]_  = ~A268 & ~A266;
  assign \new_[67646]_  = ~A234 & \new_[67645]_ ;
  assign \new_[67649]_  = A298 & ~A269;
  assign \new_[67652]_  = ~A302 & ~A301;
  assign \new_[67653]_  = \new_[67652]_  & \new_[67649]_ ;
  assign \new_[67654]_  = \new_[67653]_  & \new_[67646]_ ;
  assign \new_[67658]_  = A167 & ~A168;
  assign \new_[67659]_  = A169 & \new_[67658]_ ;
  assign \new_[67662]_  = ~A199 & ~A166;
  assign \new_[67665]_  = A232 & A200;
  assign \new_[67666]_  = \new_[67665]_  & \new_[67662]_ ;
  assign \new_[67667]_  = \new_[67666]_  & \new_[67659]_ ;
  assign \new_[67671]_  = A235 & A234;
  assign \new_[67672]_  = ~A233 & \new_[67671]_ ;
  assign \new_[67675]_  = ~A299 & A298;
  assign \new_[67678]_  = A301 & A300;
  assign \new_[67679]_  = \new_[67678]_  & \new_[67675]_ ;
  assign \new_[67680]_  = \new_[67679]_  & \new_[67672]_ ;
  assign \new_[67684]_  = A167 & ~A168;
  assign \new_[67685]_  = A169 & \new_[67684]_ ;
  assign \new_[67688]_  = ~A199 & ~A166;
  assign \new_[67691]_  = A232 & A200;
  assign \new_[67692]_  = \new_[67691]_  & \new_[67688]_ ;
  assign \new_[67693]_  = \new_[67692]_  & \new_[67685]_ ;
  assign \new_[67697]_  = A235 & A234;
  assign \new_[67698]_  = ~A233 & \new_[67697]_ ;
  assign \new_[67701]_  = ~A299 & A298;
  assign \new_[67704]_  = A302 & A300;
  assign \new_[67705]_  = \new_[67704]_  & \new_[67701]_ ;
  assign \new_[67706]_  = \new_[67705]_  & \new_[67698]_ ;
  assign \new_[67710]_  = A167 & ~A168;
  assign \new_[67711]_  = A169 & \new_[67710]_ ;
  assign \new_[67714]_  = ~A199 & ~A166;
  assign \new_[67717]_  = A232 & A200;
  assign \new_[67718]_  = \new_[67717]_  & \new_[67714]_ ;
  assign \new_[67719]_  = \new_[67718]_  & \new_[67711]_ ;
  assign \new_[67723]_  = A235 & A234;
  assign \new_[67724]_  = ~A233 & \new_[67723]_ ;
  assign \new_[67727]_  = ~A266 & A265;
  assign \new_[67730]_  = A268 & A267;
  assign \new_[67731]_  = \new_[67730]_  & \new_[67727]_ ;
  assign \new_[67732]_  = \new_[67731]_  & \new_[67724]_ ;
  assign \new_[67736]_  = A167 & ~A168;
  assign \new_[67737]_  = A169 & \new_[67736]_ ;
  assign \new_[67740]_  = ~A199 & ~A166;
  assign \new_[67743]_  = A232 & A200;
  assign \new_[67744]_  = \new_[67743]_  & \new_[67740]_ ;
  assign \new_[67745]_  = \new_[67744]_  & \new_[67737]_ ;
  assign \new_[67749]_  = A235 & A234;
  assign \new_[67750]_  = ~A233 & \new_[67749]_ ;
  assign \new_[67753]_  = ~A266 & A265;
  assign \new_[67756]_  = A269 & A267;
  assign \new_[67757]_  = \new_[67756]_  & \new_[67753]_ ;
  assign \new_[67758]_  = \new_[67757]_  & \new_[67750]_ ;
  assign \new_[67762]_  = A167 & ~A168;
  assign \new_[67763]_  = A169 & \new_[67762]_ ;
  assign \new_[67766]_  = ~A199 & ~A166;
  assign \new_[67769]_  = A232 & A200;
  assign \new_[67770]_  = \new_[67769]_  & \new_[67766]_ ;
  assign \new_[67771]_  = \new_[67770]_  & \new_[67763]_ ;
  assign \new_[67775]_  = A236 & A234;
  assign \new_[67776]_  = ~A233 & \new_[67775]_ ;
  assign \new_[67779]_  = ~A299 & A298;
  assign \new_[67782]_  = A301 & A300;
  assign \new_[67783]_  = \new_[67782]_  & \new_[67779]_ ;
  assign \new_[67784]_  = \new_[67783]_  & \new_[67776]_ ;
  assign \new_[67788]_  = A167 & ~A168;
  assign \new_[67789]_  = A169 & \new_[67788]_ ;
  assign \new_[67792]_  = ~A199 & ~A166;
  assign \new_[67795]_  = A232 & A200;
  assign \new_[67796]_  = \new_[67795]_  & \new_[67792]_ ;
  assign \new_[67797]_  = \new_[67796]_  & \new_[67789]_ ;
  assign \new_[67801]_  = A236 & A234;
  assign \new_[67802]_  = ~A233 & \new_[67801]_ ;
  assign \new_[67805]_  = ~A299 & A298;
  assign \new_[67808]_  = A302 & A300;
  assign \new_[67809]_  = \new_[67808]_  & \new_[67805]_ ;
  assign \new_[67810]_  = \new_[67809]_  & \new_[67802]_ ;
  assign \new_[67814]_  = A167 & ~A168;
  assign \new_[67815]_  = A169 & \new_[67814]_ ;
  assign \new_[67818]_  = ~A199 & ~A166;
  assign \new_[67821]_  = A232 & A200;
  assign \new_[67822]_  = \new_[67821]_  & \new_[67818]_ ;
  assign \new_[67823]_  = \new_[67822]_  & \new_[67815]_ ;
  assign \new_[67827]_  = A236 & A234;
  assign \new_[67828]_  = ~A233 & \new_[67827]_ ;
  assign \new_[67831]_  = ~A266 & A265;
  assign \new_[67834]_  = A268 & A267;
  assign \new_[67835]_  = \new_[67834]_  & \new_[67831]_ ;
  assign \new_[67836]_  = \new_[67835]_  & \new_[67828]_ ;
  assign \new_[67840]_  = A167 & ~A168;
  assign \new_[67841]_  = A169 & \new_[67840]_ ;
  assign \new_[67844]_  = ~A199 & ~A166;
  assign \new_[67847]_  = A232 & A200;
  assign \new_[67848]_  = \new_[67847]_  & \new_[67844]_ ;
  assign \new_[67849]_  = \new_[67848]_  & \new_[67841]_ ;
  assign \new_[67853]_  = A236 & A234;
  assign \new_[67854]_  = ~A233 & \new_[67853]_ ;
  assign \new_[67857]_  = ~A266 & A265;
  assign \new_[67860]_  = A269 & A267;
  assign \new_[67861]_  = \new_[67860]_  & \new_[67857]_ ;
  assign \new_[67862]_  = \new_[67861]_  & \new_[67854]_ ;
  assign \new_[67866]_  = A167 & ~A168;
  assign \new_[67867]_  = A169 & \new_[67866]_ ;
  assign \new_[67870]_  = ~A199 & ~A166;
  assign \new_[67873]_  = ~A232 & A200;
  assign \new_[67874]_  = \new_[67873]_  & \new_[67870]_ ;
  assign \new_[67875]_  = \new_[67874]_  & \new_[67867]_ ;
  assign \new_[67879]_  = ~A268 & ~A266;
  assign \new_[67880]_  = ~A233 & \new_[67879]_ ;
  assign \new_[67883]_  = A298 & ~A269;
  assign \new_[67886]_  = ~A302 & ~A301;
  assign \new_[67887]_  = \new_[67886]_  & \new_[67883]_ ;
  assign \new_[67888]_  = \new_[67887]_  & \new_[67880]_ ;
  assign \new_[67892]_  = A167 & ~A168;
  assign \new_[67893]_  = A169 & \new_[67892]_ ;
  assign \new_[67896]_  = A199 & ~A166;
  assign \new_[67899]_  = A201 & ~A200;
  assign \new_[67900]_  = \new_[67899]_  & \new_[67896]_ ;
  assign \new_[67901]_  = \new_[67900]_  & \new_[67893]_ ;
  assign \new_[67905]_  = A233 & A232;
  assign \new_[67906]_  = A202 & \new_[67905]_ ;
  assign \new_[67909]_  = ~A267 & A265;
  assign \new_[67912]_  = ~A300 & ~A299;
  assign \new_[67913]_  = \new_[67912]_  & \new_[67909]_ ;
  assign \new_[67914]_  = \new_[67913]_  & \new_[67906]_ ;
  assign \new_[67918]_  = A167 & ~A168;
  assign \new_[67919]_  = A169 & \new_[67918]_ ;
  assign \new_[67922]_  = A199 & ~A166;
  assign \new_[67925]_  = A201 & ~A200;
  assign \new_[67926]_  = \new_[67925]_  & \new_[67922]_ ;
  assign \new_[67927]_  = \new_[67926]_  & \new_[67919]_ ;
  assign \new_[67931]_  = A233 & A232;
  assign \new_[67932]_  = A202 & \new_[67931]_ ;
  assign \new_[67935]_  = ~A267 & A265;
  assign \new_[67938]_  = A299 & A298;
  assign \new_[67939]_  = \new_[67938]_  & \new_[67935]_ ;
  assign \new_[67940]_  = \new_[67939]_  & \new_[67932]_ ;
  assign \new_[67944]_  = A167 & ~A168;
  assign \new_[67945]_  = A169 & \new_[67944]_ ;
  assign \new_[67948]_  = A199 & ~A166;
  assign \new_[67951]_  = A201 & ~A200;
  assign \new_[67952]_  = \new_[67951]_  & \new_[67948]_ ;
  assign \new_[67953]_  = \new_[67952]_  & \new_[67945]_ ;
  assign \new_[67957]_  = A233 & A232;
  assign \new_[67958]_  = A202 & \new_[67957]_ ;
  assign \new_[67961]_  = ~A267 & A265;
  assign \new_[67964]_  = ~A299 & ~A298;
  assign \new_[67965]_  = \new_[67964]_  & \new_[67961]_ ;
  assign \new_[67966]_  = \new_[67965]_  & \new_[67958]_ ;
  assign \new_[67970]_  = A167 & ~A168;
  assign \new_[67971]_  = A169 & \new_[67970]_ ;
  assign \new_[67974]_  = A199 & ~A166;
  assign \new_[67977]_  = A201 & ~A200;
  assign \new_[67978]_  = \new_[67977]_  & \new_[67974]_ ;
  assign \new_[67979]_  = \new_[67978]_  & \new_[67971]_ ;
  assign \new_[67983]_  = A233 & A232;
  assign \new_[67984]_  = A202 & \new_[67983]_ ;
  assign \new_[67987]_  = A266 & A265;
  assign \new_[67990]_  = ~A300 & ~A299;
  assign \new_[67991]_  = \new_[67990]_  & \new_[67987]_ ;
  assign \new_[67992]_  = \new_[67991]_  & \new_[67984]_ ;
  assign \new_[67996]_  = A167 & ~A168;
  assign \new_[67997]_  = A169 & \new_[67996]_ ;
  assign \new_[68000]_  = A199 & ~A166;
  assign \new_[68003]_  = A201 & ~A200;
  assign \new_[68004]_  = \new_[68003]_  & \new_[68000]_ ;
  assign \new_[68005]_  = \new_[68004]_  & \new_[67997]_ ;
  assign \new_[68009]_  = A233 & A232;
  assign \new_[68010]_  = A202 & \new_[68009]_ ;
  assign \new_[68013]_  = A266 & A265;
  assign \new_[68016]_  = A299 & A298;
  assign \new_[68017]_  = \new_[68016]_  & \new_[68013]_ ;
  assign \new_[68018]_  = \new_[68017]_  & \new_[68010]_ ;
  assign \new_[68022]_  = A167 & ~A168;
  assign \new_[68023]_  = A169 & \new_[68022]_ ;
  assign \new_[68026]_  = A199 & ~A166;
  assign \new_[68029]_  = A201 & ~A200;
  assign \new_[68030]_  = \new_[68029]_  & \new_[68026]_ ;
  assign \new_[68031]_  = \new_[68030]_  & \new_[68023]_ ;
  assign \new_[68035]_  = A233 & A232;
  assign \new_[68036]_  = A202 & \new_[68035]_ ;
  assign \new_[68039]_  = A266 & A265;
  assign \new_[68042]_  = ~A299 & ~A298;
  assign \new_[68043]_  = \new_[68042]_  & \new_[68039]_ ;
  assign \new_[68044]_  = \new_[68043]_  & \new_[68036]_ ;
  assign \new_[68048]_  = A167 & ~A168;
  assign \new_[68049]_  = A169 & \new_[68048]_ ;
  assign \new_[68052]_  = A199 & ~A166;
  assign \new_[68055]_  = A201 & ~A200;
  assign \new_[68056]_  = \new_[68055]_  & \new_[68052]_ ;
  assign \new_[68057]_  = \new_[68056]_  & \new_[68049]_ ;
  assign \new_[68061]_  = A233 & A232;
  assign \new_[68062]_  = A202 & \new_[68061]_ ;
  assign \new_[68065]_  = ~A266 & ~A265;
  assign \new_[68068]_  = ~A300 & ~A299;
  assign \new_[68069]_  = \new_[68068]_  & \new_[68065]_ ;
  assign \new_[68070]_  = \new_[68069]_  & \new_[68062]_ ;
  assign \new_[68074]_  = A167 & ~A168;
  assign \new_[68075]_  = A169 & \new_[68074]_ ;
  assign \new_[68078]_  = A199 & ~A166;
  assign \new_[68081]_  = A201 & ~A200;
  assign \new_[68082]_  = \new_[68081]_  & \new_[68078]_ ;
  assign \new_[68083]_  = \new_[68082]_  & \new_[68075]_ ;
  assign \new_[68087]_  = A233 & A232;
  assign \new_[68088]_  = A202 & \new_[68087]_ ;
  assign \new_[68091]_  = ~A266 & ~A265;
  assign \new_[68094]_  = A299 & A298;
  assign \new_[68095]_  = \new_[68094]_  & \new_[68091]_ ;
  assign \new_[68096]_  = \new_[68095]_  & \new_[68088]_ ;
  assign \new_[68100]_  = A167 & ~A168;
  assign \new_[68101]_  = A169 & \new_[68100]_ ;
  assign \new_[68104]_  = A199 & ~A166;
  assign \new_[68107]_  = A201 & ~A200;
  assign \new_[68108]_  = \new_[68107]_  & \new_[68104]_ ;
  assign \new_[68109]_  = \new_[68108]_  & \new_[68101]_ ;
  assign \new_[68113]_  = A233 & A232;
  assign \new_[68114]_  = A202 & \new_[68113]_ ;
  assign \new_[68117]_  = ~A266 & ~A265;
  assign \new_[68120]_  = ~A299 & ~A298;
  assign \new_[68121]_  = \new_[68120]_  & \new_[68117]_ ;
  assign \new_[68122]_  = \new_[68121]_  & \new_[68114]_ ;
  assign \new_[68126]_  = A167 & ~A168;
  assign \new_[68127]_  = A169 & \new_[68126]_ ;
  assign \new_[68130]_  = A199 & ~A166;
  assign \new_[68133]_  = A201 & ~A200;
  assign \new_[68134]_  = \new_[68133]_  & \new_[68130]_ ;
  assign \new_[68135]_  = \new_[68134]_  & \new_[68127]_ ;
  assign \new_[68139]_  = A233 & ~A232;
  assign \new_[68140]_  = A202 & \new_[68139]_ ;
  assign \new_[68143]_  = ~A299 & A298;
  assign \new_[68146]_  = A301 & A300;
  assign \new_[68147]_  = \new_[68146]_  & \new_[68143]_ ;
  assign \new_[68148]_  = \new_[68147]_  & \new_[68140]_ ;
  assign \new_[68152]_  = A167 & ~A168;
  assign \new_[68153]_  = A169 & \new_[68152]_ ;
  assign \new_[68156]_  = A199 & ~A166;
  assign \new_[68159]_  = A201 & ~A200;
  assign \new_[68160]_  = \new_[68159]_  & \new_[68156]_ ;
  assign \new_[68161]_  = \new_[68160]_  & \new_[68153]_ ;
  assign \new_[68165]_  = A233 & ~A232;
  assign \new_[68166]_  = A202 & \new_[68165]_ ;
  assign \new_[68169]_  = ~A299 & A298;
  assign \new_[68172]_  = A302 & A300;
  assign \new_[68173]_  = \new_[68172]_  & \new_[68169]_ ;
  assign \new_[68174]_  = \new_[68173]_  & \new_[68166]_ ;
  assign \new_[68178]_  = A167 & ~A168;
  assign \new_[68179]_  = A169 & \new_[68178]_ ;
  assign \new_[68182]_  = A199 & ~A166;
  assign \new_[68185]_  = A201 & ~A200;
  assign \new_[68186]_  = \new_[68185]_  & \new_[68182]_ ;
  assign \new_[68187]_  = \new_[68186]_  & \new_[68179]_ ;
  assign \new_[68191]_  = A233 & ~A232;
  assign \new_[68192]_  = A202 & \new_[68191]_ ;
  assign \new_[68195]_  = ~A266 & A265;
  assign \new_[68198]_  = A268 & A267;
  assign \new_[68199]_  = \new_[68198]_  & \new_[68195]_ ;
  assign \new_[68200]_  = \new_[68199]_  & \new_[68192]_ ;
  assign \new_[68204]_  = A167 & ~A168;
  assign \new_[68205]_  = A169 & \new_[68204]_ ;
  assign \new_[68208]_  = A199 & ~A166;
  assign \new_[68211]_  = A201 & ~A200;
  assign \new_[68212]_  = \new_[68211]_  & \new_[68208]_ ;
  assign \new_[68213]_  = \new_[68212]_  & \new_[68205]_ ;
  assign \new_[68217]_  = A233 & ~A232;
  assign \new_[68218]_  = A202 & \new_[68217]_ ;
  assign \new_[68221]_  = ~A266 & A265;
  assign \new_[68224]_  = A269 & A267;
  assign \new_[68225]_  = \new_[68224]_  & \new_[68221]_ ;
  assign \new_[68226]_  = \new_[68225]_  & \new_[68218]_ ;
  assign \new_[68230]_  = A167 & ~A168;
  assign \new_[68231]_  = A169 & \new_[68230]_ ;
  assign \new_[68234]_  = A199 & ~A166;
  assign \new_[68237]_  = A201 & ~A200;
  assign \new_[68238]_  = \new_[68237]_  & \new_[68234]_ ;
  assign \new_[68239]_  = \new_[68238]_  & \new_[68231]_ ;
  assign \new_[68243]_  = ~A234 & ~A233;
  assign \new_[68244]_  = A202 & \new_[68243]_ ;
  assign \new_[68247]_  = A266 & A265;
  assign \new_[68250]_  = ~A300 & A298;
  assign \new_[68251]_  = \new_[68250]_  & \new_[68247]_ ;
  assign \new_[68252]_  = \new_[68251]_  & \new_[68244]_ ;
  assign \new_[68256]_  = A167 & ~A168;
  assign \new_[68257]_  = A169 & \new_[68256]_ ;
  assign \new_[68260]_  = A199 & ~A166;
  assign \new_[68263]_  = A201 & ~A200;
  assign \new_[68264]_  = \new_[68263]_  & \new_[68260]_ ;
  assign \new_[68265]_  = \new_[68264]_  & \new_[68257]_ ;
  assign \new_[68269]_  = ~A234 & ~A233;
  assign \new_[68270]_  = A202 & \new_[68269]_ ;
  assign \new_[68273]_  = A266 & A265;
  assign \new_[68276]_  = A299 & A298;
  assign \new_[68277]_  = \new_[68276]_  & \new_[68273]_ ;
  assign \new_[68278]_  = \new_[68277]_  & \new_[68270]_ ;
  assign \new_[68282]_  = A167 & ~A168;
  assign \new_[68283]_  = A169 & \new_[68282]_ ;
  assign \new_[68286]_  = A199 & ~A166;
  assign \new_[68289]_  = A201 & ~A200;
  assign \new_[68290]_  = \new_[68289]_  & \new_[68286]_ ;
  assign \new_[68291]_  = \new_[68290]_  & \new_[68283]_ ;
  assign \new_[68295]_  = ~A234 & ~A233;
  assign \new_[68296]_  = A202 & \new_[68295]_ ;
  assign \new_[68299]_  = A266 & A265;
  assign \new_[68302]_  = ~A299 & ~A298;
  assign \new_[68303]_  = \new_[68302]_  & \new_[68299]_ ;
  assign \new_[68304]_  = \new_[68303]_  & \new_[68296]_ ;
  assign \new_[68308]_  = A167 & ~A168;
  assign \new_[68309]_  = A169 & \new_[68308]_ ;
  assign \new_[68312]_  = A199 & ~A166;
  assign \new_[68315]_  = A201 & ~A200;
  assign \new_[68316]_  = \new_[68315]_  & \new_[68312]_ ;
  assign \new_[68317]_  = \new_[68316]_  & \new_[68309]_ ;
  assign \new_[68321]_  = ~A234 & ~A233;
  assign \new_[68322]_  = A202 & \new_[68321]_ ;
  assign \new_[68325]_  = ~A267 & ~A266;
  assign \new_[68328]_  = ~A300 & A298;
  assign \new_[68329]_  = \new_[68328]_  & \new_[68325]_ ;
  assign \new_[68330]_  = \new_[68329]_  & \new_[68322]_ ;
  assign \new_[68334]_  = A167 & ~A168;
  assign \new_[68335]_  = A169 & \new_[68334]_ ;
  assign \new_[68338]_  = A199 & ~A166;
  assign \new_[68341]_  = A201 & ~A200;
  assign \new_[68342]_  = \new_[68341]_  & \new_[68338]_ ;
  assign \new_[68343]_  = \new_[68342]_  & \new_[68335]_ ;
  assign \new_[68347]_  = ~A234 & ~A233;
  assign \new_[68348]_  = A202 & \new_[68347]_ ;
  assign \new_[68351]_  = ~A267 & ~A266;
  assign \new_[68354]_  = A299 & A298;
  assign \new_[68355]_  = \new_[68354]_  & \new_[68351]_ ;
  assign \new_[68356]_  = \new_[68355]_  & \new_[68348]_ ;
  assign \new_[68360]_  = A167 & ~A168;
  assign \new_[68361]_  = A169 & \new_[68360]_ ;
  assign \new_[68364]_  = A199 & ~A166;
  assign \new_[68367]_  = A201 & ~A200;
  assign \new_[68368]_  = \new_[68367]_  & \new_[68364]_ ;
  assign \new_[68369]_  = \new_[68368]_  & \new_[68361]_ ;
  assign \new_[68373]_  = ~A234 & ~A233;
  assign \new_[68374]_  = A202 & \new_[68373]_ ;
  assign \new_[68377]_  = ~A267 & ~A266;
  assign \new_[68380]_  = ~A299 & ~A298;
  assign \new_[68381]_  = \new_[68380]_  & \new_[68377]_ ;
  assign \new_[68382]_  = \new_[68381]_  & \new_[68374]_ ;
  assign \new_[68386]_  = A167 & ~A168;
  assign \new_[68387]_  = A169 & \new_[68386]_ ;
  assign \new_[68390]_  = A199 & ~A166;
  assign \new_[68393]_  = A201 & ~A200;
  assign \new_[68394]_  = \new_[68393]_  & \new_[68390]_ ;
  assign \new_[68395]_  = \new_[68394]_  & \new_[68387]_ ;
  assign \new_[68399]_  = ~A234 & ~A233;
  assign \new_[68400]_  = A202 & \new_[68399]_ ;
  assign \new_[68403]_  = ~A266 & ~A265;
  assign \new_[68406]_  = ~A300 & A298;
  assign \new_[68407]_  = \new_[68406]_  & \new_[68403]_ ;
  assign \new_[68408]_  = \new_[68407]_  & \new_[68400]_ ;
  assign \new_[68412]_  = A167 & ~A168;
  assign \new_[68413]_  = A169 & \new_[68412]_ ;
  assign \new_[68416]_  = A199 & ~A166;
  assign \new_[68419]_  = A201 & ~A200;
  assign \new_[68420]_  = \new_[68419]_  & \new_[68416]_ ;
  assign \new_[68421]_  = \new_[68420]_  & \new_[68413]_ ;
  assign \new_[68425]_  = ~A234 & ~A233;
  assign \new_[68426]_  = A202 & \new_[68425]_ ;
  assign \new_[68429]_  = ~A266 & ~A265;
  assign \new_[68432]_  = A299 & A298;
  assign \new_[68433]_  = \new_[68432]_  & \new_[68429]_ ;
  assign \new_[68434]_  = \new_[68433]_  & \new_[68426]_ ;
  assign \new_[68438]_  = A167 & ~A168;
  assign \new_[68439]_  = A169 & \new_[68438]_ ;
  assign \new_[68442]_  = A199 & ~A166;
  assign \new_[68445]_  = A201 & ~A200;
  assign \new_[68446]_  = \new_[68445]_  & \new_[68442]_ ;
  assign \new_[68447]_  = \new_[68446]_  & \new_[68439]_ ;
  assign \new_[68451]_  = ~A234 & ~A233;
  assign \new_[68452]_  = A202 & \new_[68451]_ ;
  assign \new_[68455]_  = ~A266 & ~A265;
  assign \new_[68458]_  = ~A299 & ~A298;
  assign \new_[68459]_  = \new_[68458]_  & \new_[68455]_ ;
  assign \new_[68460]_  = \new_[68459]_  & \new_[68452]_ ;
  assign \new_[68464]_  = A167 & ~A168;
  assign \new_[68465]_  = A169 & \new_[68464]_ ;
  assign \new_[68468]_  = A199 & ~A166;
  assign \new_[68471]_  = A201 & ~A200;
  assign \new_[68472]_  = \new_[68471]_  & \new_[68468]_ ;
  assign \new_[68473]_  = \new_[68472]_  & \new_[68465]_ ;
  assign \new_[68477]_  = ~A233 & A232;
  assign \new_[68478]_  = A202 & \new_[68477]_ ;
  assign \new_[68481]_  = A235 & A234;
  assign \new_[68484]_  = A299 & ~A298;
  assign \new_[68485]_  = \new_[68484]_  & \new_[68481]_ ;
  assign \new_[68486]_  = \new_[68485]_  & \new_[68478]_ ;
  assign \new_[68490]_  = A167 & ~A168;
  assign \new_[68491]_  = A169 & \new_[68490]_ ;
  assign \new_[68494]_  = A199 & ~A166;
  assign \new_[68497]_  = A201 & ~A200;
  assign \new_[68498]_  = \new_[68497]_  & \new_[68494]_ ;
  assign \new_[68499]_  = \new_[68498]_  & \new_[68491]_ ;
  assign \new_[68503]_  = ~A233 & A232;
  assign \new_[68504]_  = A202 & \new_[68503]_ ;
  assign \new_[68507]_  = A235 & A234;
  assign \new_[68510]_  = A266 & ~A265;
  assign \new_[68511]_  = \new_[68510]_  & \new_[68507]_ ;
  assign \new_[68512]_  = \new_[68511]_  & \new_[68504]_ ;
  assign \new_[68516]_  = A167 & ~A168;
  assign \new_[68517]_  = A169 & \new_[68516]_ ;
  assign \new_[68520]_  = A199 & ~A166;
  assign \new_[68523]_  = A201 & ~A200;
  assign \new_[68524]_  = \new_[68523]_  & \new_[68520]_ ;
  assign \new_[68525]_  = \new_[68524]_  & \new_[68517]_ ;
  assign \new_[68529]_  = ~A233 & A232;
  assign \new_[68530]_  = A202 & \new_[68529]_ ;
  assign \new_[68533]_  = A236 & A234;
  assign \new_[68536]_  = A299 & ~A298;
  assign \new_[68537]_  = \new_[68536]_  & \new_[68533]_ ;
  assign \new_[68538]_  = \new_[68537]_  & \new_[68530]_ ;
  assign \new_[68542]_  = A167 & ~A168;
  assign \new_[68543]_  = A169 & \new_[68542]_ ;
  assign \new_[68546]_  = A199 & ~A166;
  assign \new_[68549]_  = A201 & ~A200;
  assign \new_[68550]_  = \new_[68549]_  & \new_[68546]_ ;
  assign \new_[68551]_  = \new_[68550]_  & \new_[68543]_ ;
  assign \new_[68555]_  = ~A233 & A232;
  assign \new_[68556]_  = A202 & \new_[68555]_ ;
  assign \new_[68559]_  = A236 & A234;
  assign \new_[68562]_  = A266 & ~A265;
  assign \new_[68563]_  = \new_[68562]_  & \new_[68559]_ ;
  assign \new_[68564]_  = \new_[68563]_  & \new_[68556]_ ;
  assign \new_[68568]_  = A167 & ~A168;
  assign \new_[68569]_  = A169 & \new_[68568]_ ;
  assign \new_[68572]_  = A199 & ~A166;
  assign \new_[68575]_  = A201 & ~A200;
  assign \new_[68576]_  = \new_[68575]_  & \new_[68572]_ ;
  assign \new_[68577]_  = \new_[68576]_  & \new_[68569]_ ;
  assign \new_[68581]_  = ~A233 & ~A232;
  assign \new_[68582]_  = A202 & \new_[68581]_ ;
  assign \new_[68585]_  = A266 & A265;
  assign \new_[68588]_  = ~A300 & A298;
  assign \new_[68589]_  = \new_[68588]_  & \new_[68585]_ ;
  assign \new_[68590]_  = \new_[68589]_  & \new_[68582]_ ;
  assign \new_[68594]_  = A167 & ~A168;
  assign \new_[68595]_  = A169 & \new_[68594]_ ;
  assign \new_[68598]_  = A199 & ~A166;
  assign \new_[68601]_  = A201 & ~A200;
  assign \new_[68602]_  = \new_[68601]_  & \new_[68598]_ ;
  assign \new_[68603]_  = \new_[68602]_  & \new_[68595]_ ;
  assign \new_[68607]_  = ~A233 & ~A232;
  assign \new_[68608]_  = A202 & \new_[68607]_ ;
  assign \new_[68611]_  = A266 & A265;
  assign \new_[68614]_  = A299 & A298;
  assign \new_[68615]_  = \new_[68614]_  & \new_[68611]_ ;
  assign \new_[68616]_  = \new_[68615]_  & \new_[68608]_ ;
  assign \new_[68620]_  = A167 & ~A168;
  assign \new_[68621]_  = A169 & \new_[68620]_ ;
  assign \new_[68624]_  = A199 & ~A166;
  assign \new_[68627]_  = A201 & ~A200;
  assign \new_[68628]_  = \new_[68627]_  & \new_[68624]_ ;
  assign \new_[68629]_  = \new_[68628]_  & \new_[68621]_ ;
  assign \new_[68633]_  = ~A233 & ~A232;
  assign \new_[68634]_  = A202 & \new_[68633]_ ;
  assign \new_[68637]_  = A266 & A265;
  assign \new_[68640]_  = ~A299 & ~A298;
  assign \new_[68641]_  = \new_[68640]_  & \new_[68637]_ ;
  assign \new_[68642]_  = \new_[68641]_  & \new_[68634]_ ;
  assign \new_[68646]_  = A167 & ~A168;
  assign \new_[68647]_  = A169 & \new_[68646]_ ;
  assign \new_[68650]_  = A199 & ~A166;
  assign \new_[68653]_  = A201 & ~A200;
  assign \new_[68654]_  = \new_[68653]_  & \new_[68650]_ ;
  assign \new_[68655]_  = \new_[68654]_  & \new_[68647]_ ;
  assign \new_[68659]_  = ~A233 & ~A232;
  assign \new_[68660]_  = A202 & \new_[68659]_ ;
  assign \new_[68663]_  = ~A267 & ~A266;
  assign \new_[68666]_  = ~A300 & A298;
  assign \new_[68667]_  = \new_[68666]_  & \new_[68663]_ ;
  assign \new_[68668]_  = \new_[68667]_  & \new_[68660]_ ;
  assign \new_[68672]_  = A167 & ~A168;
  assign \new_[68673]_  = A169 & \new_[68672]_ ;
  assign \new_[68676]_  = A199 & ~A166;
  assign \new_[68679]_  = A201 & ~A200;
  assign \new_[68680]_  = \new_[68679]_  & \new_[68676]_ ;
  assign \new_[68681]_  = \new_[68680]_  & \new_[68673]_ ;
  assign \new_[68685]_  = ~A233 & ~A232;
  assign \new_[68686]_  = A202 & \new_[68685]_ ;
  assign \new_[68689]_  = ~A267 & ~A266;
  assign \new_[68692]_  = A299 & A298;
  assign \new_[68693]_  = \new_[68692]_  & \new_[68689]_ ;
  assign \new_[68694]_  = \new_[68693]_  & \new_[68686]_ ;
  assign \new_[68698]_  = A167 & ~A168;
  assign \new_[68699]_  = A169 & \new_[68698]_ ;
  assign \new_[68702]_  = A199 & ~A166;
  assign \new_[68705]_  = A201 & ~A200;
  assign \new_[68706]_  = \new_[68705]_  & \new_[68702]_ ;
  assign \new_[68707]_  = \new_[68706]_  & \new_[68699]_ ;
  assign \new_[68711]_  = ~A233 & ~A232;
  assign \new_[68712]_  = A202 & \new_[68711]_ ;
  assign \new_[68715]_  = ~A267 & ~A266;
  assign \new_[68718]_  = ~A299 & ~A298;
  assign \new_[68719]_  = \new_[68718]_  & \new_[68715]_ ;
  assign \new_[68720]_  = \new_[68719]_  & \new_[68712]_ ;
  assign \new_[68724]_  = A167 & ~A168;
  assign \new_[68725]_  = A169 & \new_[68724]_ ;
  assign \new_[68728]_  = A199 & ~A166;
  assign \new_[68731]_  = A201 & ~A200;
  assign \new_[68732]_  = \new_[68731]_  & \new_[68728]_ ;
  assign \new_[68733]_  = \new_[68732]_  & \new_[68725]_ ;
  assign \new_[68737]_  = ~A233 & ~A232;
  assign \new_[68738]_  = A202 & \new_[68737]_ ;
  assign \new_[68741]_  = ~A266 & ~A265;
  assign \new_[68744]_  = ~A300 & A298;
  assign \new_[68745]_  = \new_[68744]_  & \new_[68741]_ ;
  assign \new_[68746]_  = \new_[68745]_  & \new_[68738]_ ;
  assign \new_[68750]_  = A167 & ~A168;
  assign \new_[68751]_  = A169 & \new_[68750]_ ;
  assign \new_[68754]_  = A199 & ~A166;
  assign \new_[68757]_  = A201 & ~A200;
  assign \new_[68758]_  = \new_[68757]_  & \new_[68754]_ ;
  assign \new_[68759]_  = \new_[68758]_  & \new_[68751]_ ;
  assign \new_[68763]_  = ~A233 & ~A232;
  assign \new_[68764]_  = A202 & \new_[68763]_ ;
  assign \new_[68767]_  = ~A266 & ~A265;
  assign \new_[68770]_  = A299 & A298;
  assign \new_[68771]_  = \new_[68770]_  & \new_[68767]_ ;
  assign \new_[68772]_  = \new_[68771]_  & \new_[68764]_ ;
  assign \new_[68776]_  = A167 & ~A168;
  assign \new_[68777]_  = A169 & \new_[68776]_ ;
  assign \new_[68780]_  = A199 & ~A166;
  assign \new_[68783]_  = A201 & ~A200;
  assign \new_[68784]_  = \new_[68783]_  & \new_[68780]_ ;
  assign \new_[68785]_  = \new_[68784]_  & \new_[68777]_ ;
  assign \new_[68789]_  = ~A233 & ~A232;
  assign \new_[68790]_  = A202 & \new_[68789]_ ;
  assign \new_[68793]_  = ~A266 & ~A265;
  assign \new_[68796]_  = ~A299 & ~A298;
  assign \new_[68797]_  = \new_[68796]_  & \new_[68793]_ ;
  assign \new_[68798]_  = \new_[68797]_  & \new_[68790]_ ;
  assign \new_[68802]_  = A167 & ~A168;
  assign \new_[68803]_  = A169 & \new_[68802]_ ;
  assign \new_[68806]_  = A199 & ~A166;
  assign \new_[68809]_  = A201 & ~A200;
  assign \new_[68810]_  = \new_[68809]_  & \new_[68806]_ ;
  assign \new_[68811]_  = \new_[68810]_  & \new_[68803]_ ;
  assign \new_[68815]_  = A233 & A232;
  assign \new_[68816]_  = A203 & \new_[68815]_ ;
  assign \new_[68819]_  = ~A267 & A265;
  assign \new_[68822]_  = ~A300 & ~A299;
  assign \new_[68823]_  = \new_[68822]_  & \new_[68819]_ ;
  assign \new_[68824]_  = \new_[68823]_  & \new_[68816]_ ;
  assign \new_[68828]_  = A167 & ~A168;
  assign \new_[68829]_  = A169 & \new_[68828]_ ;
  assign \new_[68832]_  = A199 & ~A166;
  assign \new_[68835]_  = A201 & ~A200;
  assign \new_[68836]_  = \new_[68835]_  & \new_[68832]_ ;
  assign \new_[68837]_  = \new_[68836]_  & \new_[68829]_ ;
  assign \new_[68841]_  = A233 & A232;
  assign \new_[68842]_  = A203 & \new_[68841]_ ;
  assign \new_[68845]_  = ~A267 & A265;
  assign \new_[68848]_  = A299 & A298;
  assign \new_[68849]_  = \new_[68848]_  & \new_[68845]_ ;
  assign \new_[68850]_  = \new_[68849]_  & \new_[68842]_ ;
  assign \new_[68854]_  = A167 & ~A168;
  assign \new_[68855]_  = A169 & \new_[68854]_ ;
  assign \new_[68858]_  = A199 & ~A166;
  assign \new_[68861]_  = A201 & ~A200;
  assign \new_[68862]_  = \new_[68861]_  & \new_[68858]_ ;
  assign \new_[68863]_  = \new_[68862]_  & \new_[68855]_ ;
  assign \new_[68867]_  = A233 & A232;
  assign \new_[68868]_  = A203 & \new_[68867]_ ;
  assign \new_[68871]_  = ~A267 & A265;
  assign \new_[68874]_  = ~A299 & ~A298;
  assign \new_[68875]_  = \new_[68874]_  & \new_[68871]_ ;
  assign \new_[68876]_  = \new_[68875]_  & \new_[68868]_ ;
  assign \new_[68880]_  = A167 & ~A168;
  assign \new_[68881]_  = A169 & \new_[68880]_ ;
  assign \new_[68884]_  = A199 & ~A166;
  assign \new_[68887]_  = A201 & ~A200;
  assign \new_[68888]_  = \new_[68887]_  & \new_[68884]_ ;
  assign \new_[68889]_  = \new_[68888]_  & \new_[68881]_ ;
  assign \new_[68893]_  = A233 & A232;
  assign \new_[68894]_  = A203 & \new_[68893]_ ;
  assign \new_[68897]_  = A266 & A265;
  assign \new_[68900]_  = ~A300 & ~A299;
  assign \new_[68901]_  = \new_[68900]_  & \new_[68897]_ ;
  assign \new_[68902]_  = \new_[68901]_  & \new_[68894]_ ;
  assign \new_[68906]_  = A167 & ~A168;
  assign \new_[68907]_  = A169 & \new_[68906]_ ;
  assign \new_[68910]_  = A199 & ~A166;
  assign \new_[68913]_  = A201 & ~A200;
  assign \new_[68914]_  = \new_[68913]_  & \new_[68910]_ ;
  assign \new_[68915]_  = \new_[68914]_  & \new_[68907]_ ;
  assign \new_[68919]_  = A233 & A232;
  assign \new_[68920]_  = A203 & \new_[68919]_ ;
  assign \new_[68923]_  = A266 & A265;
  assign \new_[68926]_  = A299 & A298;
  assign \new_[68927]_  = \new_[68926]_  & \new_[68923]_ ;
  assign \new_[68928]_  = \new_[68927]_  & \new_[68920]_ ;
  assign \new_[68932]_  = A167 & ~A168;
  assign \new_[68933]_  = A169 & \new_[68932]_ ;
  assign \new_[68936]_  = A199 & ~A166;
  assign \new_[68939]_  = A201 & ~A200;
  assign \new_[68940]_  = \new_[68939]_  & \new_[68936]_ ;
  assign \new_[68941]_  = \new_[68940]_  & \new_[68933]_ ;
  assign \new_[68945]_  = A233 & A232;
  assign \new_[68946]_  = A203 & \new_[68945]_ ;
  assign \new_[68949]_  = A266 & A265;
  assign \new_[68952]_  = ~A299 & ~A298;
  assign \new_[68953]_  = \new_[68952]_  & \new_[68949]_ ;
  assign \new_[68954]_  = \new_[68953]_  & \new_[68946]_ ;
  assign \new_[68958]_  = A167 & ~A168;
  assign \new_[68959]_  = A169 & \new_[68958]_ ;
  assign \new_[68962]_  = A199 & ~A166;
  assign \new_[68965]_  = A201 & ~A200;
  assign \new_[68966]_  = \new_[68965]_  & \new_[68962]_ ;
  assign \new_[68967]_  = \new_[68966]_  & \new_[68959]_ ;
  assign \new_[68971]_  = A233 & A232;
  assign \new_[68972]_  = A203 & \new_[68971]_ ;
  assign \new_[68975]_  = ~A266 & ~A265;
  assign \new_[68978]_  = ~A300 & ~A299;
  assign \new_[68979]_  = \new_[68978]_  & \new_[68975]_ ;
  assign \new_[68980]_  = \new_[68979]_  & \new_[68972]_ ;
  assign \new_[68984]_  = A167 & ~A168;
  assign \new_[68985]_  = A169 & \new_[68984]_ ;
  assign \new_[68988]_  = A199 & ~A166;
  assign \new_[68991]_  = A201 & ~A200;
  assign \new_[68992]_  = \new_[68991]_  & \new_[68988]_ ;
  assign \new_[68993]_  = \new_[68992]_  & \new_[68985]_ ;
  assign \new_[68997]_  = A233 & A232;
  assign \new_[68998]_  = A203 & \new_[68997]_ ;
  assign \new_[69001]_  = ~A266 & ~A265;
  assign \new_[69004]_  = A299 & A298;
  assign \new_[69005]_  = \new_[69004]_  & \new_[69001]_ ;
  assign \new_[69006]_  = \new_[69005]_  & \new_[68998]_ ;
  assign \new_[69010]_  = A167 & ~A168;
  assign \new_[69011]_  = A169 & \new_[69010]_ ;
  assign \new_[69014]_  = A199 & ~A166;
  assign \new_[69017]_  = A201 & ~A200;
  assign \new_[69018]_  = \new_[69017]_  & \new_[69014]_ ;
  assign \new_[69019]_  = \new_[69018]_  & \new_[69011]_ ;
  assign \new_[69023]_  = A233 & A232;
  assign \new_[69024]_  = A203 & \new_[69023]_ ;
  assign \new_[69027]_  = ~A266 & ~A265;
  assign \new_[69030]_  = ~A299 & ~A298;
  assign \new_[69031]_  = \new_[69030]_  & \new_[69027]_ ;
  assign \new_[69032]_  = \new_[69031]_  & \new_[69024]_ ;
  assign \new_[69036]_  = A167 & ~A168;
  assign \new_[69037]_  = A169 & \new_[69036]_ ;
  assign \new_[69040]_  = A199 & ~A166;
  assign \new_[69043]_  = A201 & ~A200;
  assign \new_[69044]_  = \new_[69043]_  & \new_[69040]_ ;
  assign \new_[69045]_  = \new_[69044]_  & \new_[69037]_ ;
  assign \new_[69049]_  = A233 & ~A232;
  assign \new_[69050]_  = A203 & \new_[69049]_ ;
  assign \new_[69053]_  = ~A299 & A298;
  assign \new_[69056]_  = A301 & A300;
  assign \new_[69057]_  = \new_[69056]_  & \new_[69053]_ ;
  assign \new_[69058]_  = \new_[69057]_  & \new_[69050]_ ;
  assign \new_[69062]_  = A167 & ~A168;
  assign \new_[69063]_  = A169 & \new_[69062]_ ;
  assign \new_[69066]_  = A199 & ~A166;
  assign \new_[69069]_  = A201 & ~A200;
  assign \new_[69070]_  = \new_[69069]_  & \new_[69066]_ ;
  assign \new_[69071]_  = \new_[69070]_  & \new_[69063]_ ;
  assign \new_[69075]_  = A233 & ~A232;
  assign \new_[69076]_  = A203 & \new_[69075]_ ;
  assign \new_[69079]_  = ~A299 & A298;
  assign \new_[69082]_  = A302 & A300;
  assign \new_[69083]_  = \new_[69082]_  & \new_[69079]_ ;
  assign \new_[69084]_  = \new_[69083]_  & \new_[69076]_ ;
  assign \new_[69088]_  = A167 & ~A168;
  assign \new_[69089]_  = A169 & \new_[69088]_ ;
  assign \new_[69092]_  = A199 & ~A166;
  assign \new_[69095]_  = A201 & ~A200;
  assign \new_[69096]_  = \new_[69095]_  & \new_[69092]_ ;
  assign \new_[69097]_  = \new_[69096]_  & \new_[69089]_ ;
  assign \new_[69101]_  = A233 & ~A232;
  assign \new_[69102]_  = A203 & \new_[69101]_ ;
  assign \new_[69105]_  = ~A266 & A265;
  assign \new_[69108]_  = A268 & A267;
  assign \new_[69109]_  = \new_[69108]_  & \new_[69105]_ ;
  assign \new_[69110]_  = \new_[69109]_  & \new_[69102]_ ;
  assign \new_[69114]_  = A167 & ~A168;
  assign \new_[69115]_  = A169 & \new_[69114]_ ;
  assign \new_[69118]_  = A199 & ~A166;
  assign \new_[69121]_  = A201 & ~A200;
  assign \new_[69122]_  = \new_[69121]_  & \new_[69118]_ ;
  assign \new_[69123]_  = \new_[69122]_  & \new_[69115]_ ;
  assign \new_[69127]_  = A233 & ~A232;
  assign \new_[69128]_  = A203 & \new_[69127]_ ;
  assign \new_[69131]_  = ~A266 & A265;
  assign \new_[69134]_  = A269 & A267;
  assign \new_[69135]_  = \new_[69134]_  & \new_[69131]_ ;
  assign \new_[69136]_  = \new_[69135]_  & \new_[69128]_ ;
  assign \new_[69140]_  = A167 & ~A168;
  assign \new_[69141]_  = A169 & \new_[69140]_ ;
  assign \new_[69144]_  = A199 & ~A166;
  assign \new_[69147]_  = A201 & ~A200;
  assign \new_[69148]_  = \new_[69147]_  & \new_[69144]_ ;
  assign \new_[69149]_  = \new_[69148]_  & \new_[69141]_ ;
  assign \new_[69153]_  = ~A234 & ~A233;
  assign \new_[69154]_  = A203 & \new_[69153]_ ;
  assign \new_[69157]_  = A266 & A265;
  assign \new_[69160]_  = ~A300 & A298;
  assign \new_[69161]_  = \new_[69160]_  & \new_[69157]_ ;
  assign \new_[69162]_  = \new_[69161]_  & \new_[69154]_ ;
  assign \new_[69166]_  = A167 & ~A168;
  assign \new_[69167]_  = A169 & \new_[69166]_ ;
  assign \new_[69170]_  = A199 & ~A166;
  assign \new_[69173]_  = A201 & ~A200;
  assign \new_[69174]_  = \new_[69173]_  & \new_[69170]_ ;
  assign \new_[69175]_  = \new_[69174]_  & \new_[69167]_ ;
  assign \new_[69179]_  = ~A234 & ~A233;
  assign \new_[69180]_  = A203 & \new_[69179]_ ;
  assign \new_[69183]_  = A266 & A265;
  assign \new_[69186]_  = A299 & A298;
  assign \new_[69187]_  = \new_[69186]_  & \new_[69183]_ ;
  assign \new_[69188]_  = \new_[69187]_  & \new_[69180]_ ;
  assign \new_[69192]_  = A167 & ~A168;
  assign \new_[69193]_  = A169 & \new_[69192]_ ;
  assign \new_[69196]_  = A199 & ~A166;
  assign \new_[69199]_  = A201 & ~A200;
  assign \new_[69200]_  = \new_[69199]_  & \new_[69196]_ ;
  assign \new_[69201]_  = \new_[69200]_  & \new_[69193]_ ;
  assign \new_[69205]_  = ~A234 & ~A233;
  assign \new_[69206]_  = A203 & \new_[69205]_ ;
  assign \new_[69209]_  = A266 & A265;
  assign \new_[69212]_  = ~A299 & ~A298;
  assign \new_[69213]_  = \new_[69212]_  & \new_[69209]_ ;
  assign \new_[69214]_  = \new_[69213]_  & \new_[69206]_ ;
  assign \new_[69218]_  = A167 & ~A168;
  assign \new_[69219]_  = A169 & \new_[69218]_ ;
  assign \new_[69222]_  = A199 & ~A166;
  assign \new_[69225]_  = A201 & ~A200;
  assign \new_[69226]_  = \new_[69225]_  & \new_[69222]_ ;
  assign \new_[69227]_  = \new_[69226]_  & \new_[69219]_ ;
  assign \new_[69231]_  = ~A234 & ~A233;
  assign \new_[69232]_  = A203 & \new_[69231]_ ;
  assign \new_[69235]_  = ~A267 & ~A266;
  assign \new_[69238]_  = ~A300 & A298;
  assign \new_[69239]_  = \new_[69238]_  & \new_[69235]_ ;
  assign \new_[69240]_  = \new_[69239]_  & \new_[69232]_ ;
  assign \new_[69244]_  = A167 & ~A168;
  assign \new_[69245]_  = A169 & \new_[69244]_ ;
  assign \new_[69248]_  = A199 & ~A166;
  assign \new_[69251]_  = A201 & ~A200;
  assign \new_[69252]_  = \new_[69251]_  & \new_[69248]_ ;
  assign \new_[69253]_  = \new_[69252]_  & \new_[69245]_ ;
  assign \new_[69257]_  = ~A234 & ~A233;
  assign \new_[69258]_  = A203 & \new_[69257]_ ;
  assign \new_[69261]_  = ~A267 & ~A266;
  assign \new_[69264]_  = A299 & A298;
  assign \new_[69265]_  = \new_[69264]_  & \new_[69261]_ ;
  assign \new_[69266]_  = \new_[69265]_  & \new_[69258]_ ;
  assign \new_[69270]_  = A167 & ~A168;
  assign \new_[69271]_  = A169 & \new_[69270]_ ;
  assign \new_[69274]_  = A199 & ~A166;
  assign \new_[69277]_  = A201 & ~A200;
  assign \new_[69278]_  = \new_[69277]_  & \new_[69274]_ ;
  assign \new_[69279]_  = \new_[69278]_  & \new_[69271]_ ;
  assign \new_[69283]_  = ~A234 & ~A233;
  assign \new_[69284]_  = A203 & \new_[69283]_ ;
  assign \new_[69287]_  = ~A267 & ~A266;
  assign \new_[69290]_  = ~A299 & ~A298;
  assign \new_[69291]_  = \new_[69290]_  & \new_[69287]_ ;
  assign \new_[69292]_  = \new_[69291]_  & \new_[69284]_ ;
  assign \new_[69296]_  = A167 & ~A168;
  assign \new_[69297]_  = A169 & \new_[69296]_ ;
  assign \new_[69300]_  = A199 & ~A166;
  assign \new_[69303]_  = A201 & ~A200;
  assign \new_[69304]_  = \new_[69303]_  & \new_[69300]_ ;
  assign \new_[69305]_  = \new_[69304]_  & \new_[69297]_ ;
  assign \new_[69309]_  = ~A234 & ~A233;
  assign \new_[69310]_  = A203 & \new_[69309]_ ;
  assign \new_[69313]_  = ~A266 & ~A265;
  assign \new_[69316]_  = ~A300 & A298;
  assign \new_[69317]_  = \new_[69316]_  & \new_[69313]_ ;
  assign \new_[69318]_  = \new_[69317]_  & \new_[69310]_ ;
  assign \new_[69322]_  = A167 & ~A168;
  assign \new_[69323]_  = A169 & \new_[69322]_ ;
  assign \new_[69326]_  = A199 & ~A166;
  assign \new_[69329]_  = A201 & ~A200;
  assign \new_[69330]_  = \new_[69329]_  & \new_[69326]_ ;
  assign \new_[69331]_  = \new_[69330]_  & \new_[69323]_ ;
  assign \new_[69335]_  = ~A234 & ~A233;
  assign \new_[69336]_  = A203 & \new_[69335]_ ;
  assign \new_[69339]_  = ~A266 & ~A265;
  assign \new_[69342]_  = A299 & A298;
  assign \new_[69343]_  = \new_[69342]_  & \new_[69339]_ ;
  assign \new_[69344]_  = \new_[69343]_  & \new_[69336]_ ;
  assign \new_[69348]_  = A167 & ~A168;
  assign \new_[69349]_  = A169 & \new_[69348]_ ;
  assign \new_[69352]_  = A199 & ~A166;
  assign \new_[69355]_  = A201 & ~A200;
  assign \new_[69356]_  = \new_[69355]_  & \new_[69352]_ ;
  assign \new_[69357]_  = \new_[69356]_  & \new_[69349]_ ;
  assign \new_[69361]_  = ~A234 & ~A233;
  assign \new_[69362]_  = A203 & \new_[69361]_ ;
  assign \new_[69365]_  = ~A266 & ~A265;
  assign \new_[69368]_  = ~A299 & ~A298;
  assign \new_[69369]_  = \new_[69368]_  & \new_[69365]_ ;
  assign \new_[69370]_  = \new_[69369]_  & \new_[69362]_ ;
  assign \new_[69374]_  = A167 & ~A168;
  assign \new_[69375]_  = A169 & \new_[69374]_ ;
  assign \new_[69378]_  = A199 & ~A166;
  assign \new_[69381]_  = A201 & ~A200;
  assign \new_[69382]_  = \new_[69381]_  & \new_[69378]_ ;
  assign \new_[69383]_  = \new_[69382]_  & \new_[69375]_ ;
  assign \new_[69387]_  = ~A233 & A232;
  assign \new_[69388]_  = A203 & \new_[69387]_ ;
  assign \new_[69391]_  = A235 & A234;
  assign \new_[69394]_  = A299 & ~A298;
  assign \new_[69395]_  = \new_[69394]_  & \new_[69391]_ ;
  assign \new_[69396]_  = \new_[69395]_  & \new_[69388]_ ;
  assign \new_[69400]_  = A167 & ~A168;
  assign \new_[69401]_  = A169 & \new_[69400]_ ;
  assign \new_[69404]_  = A199 & ~A166;
  assign \new_[69407]_  = A201 & ~A200;
  assign \new_[69408]_  = \new_[69407]_  & \new_[69404]_ ;
  assign \new_[69409]_  = \new_[69408]_  & \new_[69401]_ ;
  assign \new_[69413]_  = ~A233 & A232;
  assign \new_[69414]_  = A203 & \new_[69413]_ ;
  assign \new_[69417]_  = A235 & A234;
  assign \new_[69420]_  = A266 & ~A265;
  assign \new_[69421]_  = \new_[69420]_  & \new_[69417]_ ;
  assign \new_[69422]_  = \new_[69421]_  & \new_[69414]_ ;
  assign \new_[69426]_  = A167 & ~A168;
  assign \new_[69427]_  = A169 & \new_[69426]_ ;
  assign \new_[69430]_  = A199 & ~A166;
  assign \new_[69433]_  = A201 & ~A200;
  assign \new_[69434]_  = \new_[69433]_  & \new_[69430]_ ;
  assign \new_[69435]_  = \new_[69434]_  & \new_[69427]_ ;
  assign \new_[69439]_  = ~A233 & A232;
  assign \new_[69440]_  = A203 & \new_[69439]_ ;
  assign \new_[69443]_  = A236 & A234;
  assign \new_[69446]_  = A299 & ~A298;
  assign \new_[69447]_  = \new_[69446]_  & \new_[69443]_ ;
  assign \new_[69448]_  = \new_[69447]_  & \new_[69440]_ ;
  assign \new_[69452]_  = A167 & ~A168;
  assign \new_[69453]_  = A169 & \new_[69452]_ ;
  assign \new_[69456]_  = A199 & ~A166;
  assign \new_[69459]_  = A201 & ~A200;
  assign \new_[69460]_  = \new_[69459]_  & \new_[69456]_ ;
  assign \new_[69461]_  = \new_[69460]_  & \new_[69453]_ ;
  assign \new_[69465]_  = ~A233 & A232;
  assign \new_[69466]_  = A203 & \new_[69465]_ ;
  assign \new_[69469]_  = A236 & A234;
  assign \new_[69472]_  = A266 & ~A265;
  assign \new_[69473]_  = \new_[69472]_  & \new_[69469]_ ;
  assign \new_[69474]_  = \new_[69473]_  & \new_[69466]_ ;
  assign \new_[69478]_  = A167 & ~A168;
  assign \new_[69479]_  = A169 & \new_[69478]_ ;
  assign \new_[69482]_  = A199 & ~A166;
  assign \new_[69485]_  = A201 & ~A200;
  assign \new_[69486]_  = \new_[69485]_  & \new_[69482]_ ;
  assign \new_[69487]_  = \new_[69486]_  & \new_[69479]_ ;
  assign \new_[69491]_  = ~A233 & ~A232;
  assign \new_[69492]_  = A203 & \new_[69491]_ ;
  assign \new_[69495]_  = A266 & A265;
  assign \new_[69498]_  = ~A300 & A298;
  assign \new_[69499]_  = \new_[69498]_  & \new_[69495]_ ;
  assign \new_[69500]_  = \new_[69499]_  & \new_[69492]_ ;
  assign \new_[69504]_  = A167 & ~A168;
  assign \new_[69505]_  = A169 & \new_[69504]_ ;
  assign \new_[69508]_  = A199 & ~A166;
  assign \new_[69511]_  = A201 & ~A200;
  assign \new_[69512]_  = \new_[69511]_  & \new_[69508]_ ;
  assign \new_[69513]_  = \new_[69512]_  & \new_[69505]_ ;
  assign \new_[69517]_  = ~A233 & ~A232;
  assign \new_[69518]_  = A203 & \new_[69517]_ ;
  assign \new_[69521]_  = A266 & A265;
  assign \new_[69524]_  = A299 & A298;
  assign \new_[69525]_  = \new_[69524]_  & \new_[69521]_ ;
  assign \new_[69526]_  = \new_[69525]_  & \new_[69518]_ ;
  assign \new_[69530]_  = A167 & ~A168;
  assign \new_[69531]_  = A169 & \new_[69530]_ ;
  assign \new_[69534]_  = A199 & ~A166;
  assign \new_[69537]_  = A201 & ~A200;
  assign \new_[69538]_  = \new_[69537]_  & \new_[69534]_ ;
  assign \new_[69539]_  = \new_[69538]_  & \new_[69531]_ ;
  assign \new_[69543]_  = ~A233 & ~A232;
  assign \new_[69544]_  = A203 & \new_[69543]_ ;
  assign \new_[69547]_  = A266 & A265;
  assign \new_[69550]_  = ~A299 & ~A298;
  assign \new_[69551]_  = \new_[69550]_  & \new_[69547]_ ;
  assign \new_[69552]_  = \new_[69551]_  & \new_[69544]_ ;
  assign \new_[69556]_  = A167 & ~A168;
  assign \new_[69557]_  = A169 & \new_[69556]_ ;
  assign \new_[69560]_  = A199 & ~A166;
  assign \new_[69563]_  = A201 & ~A200;
  assign \new_[69564]_  = \new_[69563]_  & \new_[69560]_ ;
  assign \new_[69565]_  = \new_[69564]_  & \new_[69557]_ ;
  assign \new_[69569]_  = ~A233 & ~A232;
  assign \new_[69570]_  = A203 & \new_[69569]_ ;
  assign \new_[69573]_  = ~A267 & ~A266;
  assign \new_[69576]_  = ~A300 & A298;
  assign \new_[69577]_  = \new_[69576]_  & \new_[69573]_ ;
  assign \new_[69578]_  = \new_[69577]_  & \new_[69570]_ ;
  assign \new_[69582]_  = A167 & ~A168;
  assign \new_[69583]_  = A169 & \new_[69582]_ ;
  assign \new_[69586]_  = A199 & ~A166;
  assign \new_[69589]_  = A201 & ~A200;
  assign \new_[69590]_  = \new_[69589]_  & \new_[69586]_ ;
  assign \new_[69591]_  = \new_[69590]_  & \new_[69583]_ ;
  assign \new_[69595]_  = ~A233 & ~A232;
  assign \new_[69596]_  = A203 & \new_[69595]_ ;
  assign \new_[69599]_  = ~A267 & ~A266;
  assign \new_[69602]_  = A299 & A298;
  assign \new_[69603]_  = \new_[69602]_  & \new_[69599]_ ;
  assign \new_[69604]_  = \new_[69603]_  & \new_[69596]_ ;
  assign \new_[69608]_  = A167 & ~A168;
  assign \new_[69609]_  = A169 & \new_[69608]_ ;
  assign \new_[69612]_  = A199 & ~A166;
  assign \new_[69615]_  = A201 & ~A200;
  assign \new_[69616]_  = \new_[69615]_  & \new_[69612]_ ;
  assign \new_[69617]_  = \new_[69616]_  & \new_[69609]_ ;
  assign \new_[69621]_  = ~A233 & ~A232;
  assign \new_[69622]_  = A203 & \new_[69621]_ ;
  assign \new_[69625]_  = ~A267 & ~A266;
  assign \new_[69628]_  = ~A299 & ~A298;
  assign \new_[69629]_  = \new_[69628]_  & \new_[69625]_ ;
  assign \new_[69630]_  = \new_[69629]_  & \new_[69622]_ ;
  assign \new_[69634]_  = A167 & ~A168;
  assign \new_[69635]_  = A169 & \new_[69634]_ ;
  assign \new_[69638]_  = A199 & ~A166;
  assign \new_[69641]_  = A201 & ~A200;
  assign \new_[69642]_  = \new_[69641]_  & \new_[69638]_ ;
  assign \new_[69643]_  = \new_[69642]_  & \new_[69635]_ ;
  assign \new_[69647]_  = ~A233 & ~A232;
  assign \new_[69648]_  = A203 & \new_[69647]_ ;
  assign \new_[69651]_  = ~A266 & ~A265;
  assign \new_[69654]_  = ~A300 & A298;
  assign \new_[69655]_  = \new_[69654]_  & \new_[69651]_ ;
  assign \new_[69656]_  = \new_[69655]_  & \new_[69648]_ ;
  assign \new_[69660]_  = A167 & ~A168;
  assign \new_[69661]_  = A169 & \new_[69660]_ ;
  assign \new_[69664]_  = A199 & ~A166;
  assign \new_[69667]_  = A201 & ~A200;
  assign \new_[69668]_  = \new_[69667]_  & \new_[69664]_ ;
  assign \new_[69669]_  = \new_[69668]_  & \new_[69661]_ ;
  assign \new_[69673]_  = ~A233 & ~A232;
  assign \new_[69674]_  = A203 & \new_[69673]_ ;
  assign \new_[69677]_  = ~A266 & ~A265;
  assign \new_[69680]_  = A299 & A298;
  assign \new_[69681]_  = \new_[69680]_  & \new_[69677]_ ;
  assign \new_[69682]_  = \new_[69681]_  & \new_[69674]_ ;
  assign \new_[69686]_  = A167 & ~A168;
  assign \new_[69687]_  = A169 & \new_[69686]_ ;
  assign \new_[69690]_  = A199 & ~A166;
  assign \new_[69693]_  = A201 & ~A200;
  assign \new_[69694]_  = \new_[69693]_  & \new_[69690]_ ;
  assign \new_[69695]_  = \new_[69694]_  & \new_[69687]_ ;
  assign \new_[69699]_  = ~A233 & ~A232;
  assign \new_[69700]_  = A203 & \new_[69699]_ ;
  assign \new_[69703]_  = ~A266 & ~A265;
  assign \new_[69706]_  = ~A299 & ~A298;
  assign \new_[69707]_  = \new_[69706]_  & \new_[69703]_ ;
  assign \new_[69708]_  = \new_[69707]_  & \new_[69700]_ ;
  assign \new_[69712]_  = ~A167 & ~A168;
  assign \new_[69713]_  = A169 & \new_[69712]_ ;
  assign \new_[69716]_  = ~A199 & A166;
  assign \new_[69719]_  = A232 & A200;
  assign \new_[69720]_  = \new_[69719]_  & \new_[69716]_ ;
  assign \new_[69721]_  = \new_[69720]_  & \new_[69713]_ ;
  assign \new_[69725]_  = ~A268 & A265;
  assign \new_[69726]_  = A233 & \new_[69725]_ ;
  assign \new_[69729]_  = ~A299 & ~A269;
  assign \new_[69732]_  = ~A302 & ~A301;
  assign \new_[69733]_  = \new_[69732]_  & \new_[69729]_ ;
  assign \new_[69734]_  = \new_[69733]_  & \new_[69726]_ ;
  assign \new_[69738]_  = ~A167 & ~A168;
  assign \new_[69739]_  = A169 & \new_[69738]_ ;
  assign \new_[69742]_  = ~A199 & A166;
  assign \new_[69745]_  = ~A233 & A200;
  assign \new_[69746]_  = \new_[69745]_  & \new_[69742]_ ;
  assign \new_[69747]_  = \new_[69746]_  & \new_[69739]_ ;
  assign \new_[69751]_  = A265 & ~A236;
  assign \new_[69752]_  = ~A235 & \new_[69751]_ ;
  assign \new_[69755]_  = A298 & A266;
  assign \new_[69758]_  = ~A302 & ~A301;
  assign \new_[69759]_  = \new_[69758]_  & \new_[69755]_ ;
  assign \new_[69760]_  = \new_[69759]_  & \new_[69752]_ ;
  assign \new_[69764]_  = ~A167 & ~A168;
  assign \new_[69765]_  = A169 & \new_[69764]_ ;
  assign \new_[69768]_  = ~A199 & A166;
  assign \new_[69771]_  = ~A233 & A200;
  assign \new_[69772]_  = \new_[69771]_  & \new_[69768]_ ;
  assign \new_[69773]_  = \new_[69772]_  & \new_[69765]_ ;
  assign \new_[69777]_  = ~A266 & ~A236;
  assign \new_[69778]_  = ~A235 & \new_[69777]_ ;
  assign \new_[69781]_  = ~A269 & ~A268;
  assign \new_[69784]_  = ~A300 & A298;
  assign \new_[69785]_  = \new_[69784]_  & \new_[69781]_ ;
  assign \new_[69786]_  = \new_[69785]_  & \new_[69778]_ ;
  assign \new_[69790]_  = ~A167 & ~A168;
  assign \new_[69791]_  = A169 & \new_[69790]_ ;
  assign \new_[69794]_  = ~A199 & A166;
  assign \new_[69797]_  = ~A233 & A200;
  assign \new_[69798]_  = \new_[69797]_  & \new_[69794]_ ;
  assign \new_[69799]_  = \new_[69798]_  & \new_[69791]_ ;
  assign \new_[69803]_  = ~A266 & ~A236;
  assign \new_[69804]_  = ~A235 & \new_[69803]_ ;
  assign \new_[69807]_  = ~A269 & ~A268;
  assign \new_[69810]_  = A299 & A298;
  assign \new_[69811]_  = \new_[69810]_  & \new_[69807]_ ;
  assign \new_[69812]_  = \new_[69811]_  & \new_[69804]_ ;
  assign \new_[69816]_  = ~A167 & ~A168;
  assign \new_[69817]_  = A169 & \new_[69816]_ ;
  assign \new_[69820]_  = ~A199 & A166;
  assign \new_[69823]_  = ~A233 & A200;
  assign \new_[69824]_  = \new_[69823]_  & \new_[69820]_ ;
  assign \new_[69825]_  = \new_[69824]_  & \new_[69817]_ ;
  assign \new_[69829]_  = ~A266 & ~A236;
  assign \new_[69830]_  = ~A235 & \new_[69829]_ ;
  assign \new_[69833]_  = ~A269 & ~A268;
  assign \new_[69836]_  = ~A299 & ~A298;
  assign \new_[69837]_  = \new_[69836]_  & \new_[69833]_ ;
  assign \new_[69838]_  = \new_[69837]_  & \new_[69830]_ ;
  assign \new_[69842]_  = ~A167 & ~A168;
  assign \new_[69843]_  = A169 & \new_[69842]_ ;
  assign \new_[69846]_  = ~A199 & A166;
  assign \new_[69849]_  = ~A233 & A200;
  assign \new_[69850]_  = \new_[69849]_  & \new_[69846]_ ;
  assign \new_[69851]_  = \new_[69850]_  & \new_[69843]_ ;
  assign \new_[69855]_  = ~A266 & ~A236;
  assign \new_[69856]_  = ~A235 & \new_[69855]_ ;
  assign \new_[69859]_  = A298 & ~A267;
  assign \new_[69862]_  = ~A302 & ~A301;
  assign \new_[69863]_  = \new_[69862]_  & \new_[69859]_ ;
  assign \new_[69864]_  = \new_[69863]_  & \new_[69856]_ ;
  assign \new_[69868]_  = ~A167 & ~A168;
  assign \new_[69869]_  = A169 & \new_[69868]_ ;
  assign \new_[69872]_  = ~A199 & A166;
  assign \new_[69875]_  = ~A233 & A200;
  assign \new_[69876]_  = \new_[69875]_  & \new_[69872]_ ;
  assign \new_[69877]_  = \new_[69876]_  & \new_[69869]_ ;
  assign \new_[69881]_  = ~A265 & ~A236;
  assign \new_[69882]_  = ~A235 & \new_[69881]_ ;
  assign \new_[69885]_  = A298 & ~A266;
  assign \new_[69888]_  = ~A302 & ~A301;
  assign \new_[69889]_  = \new_[69888]_  & \new_[69885]_ ;
  assign \new_[69890]_  = \new_[69889]_  & \new_[69882]_ ;
  assign \new_[69894]_  = ~A167 & ~A168;
  assign \new_[69895]_  = A169 & \new_[69894]_ ;
  assign \new_[69898]_  = ~A199 & A166;
  assign \new_[69901]_  = ~A233 & A200;
  assign \new_[69902]_  = \new_[69901]_  & \new_[69898]_ ;
  assign \new_[69903]_  = \new_[69902]_  & \new_[69895]_ ;
  assign \new_[69907]_  = ~A268 & ~A266;
  assign \new_[69908]_  = ~A234 & \new_[69907]_ ;
  assign \new_[69911]_  = A298 & ~A269;
  assign \new_[69914]_  = ~A302 & ~A301;
  assign \new_[69915]_  = \new_[69914]_  & \new_[69911]_ ;
  assign \new_[69916]_  = \new_[69915]_  & \new_[69908]_ ;
  assign \new_[69920]_  = ~A167 & ~A168;
  assign \new_[69921]_  = A169 & \new_[69920]_ ;
  assign \new_[69924]_  = ~A199 & A166;
  assign \new_[69927]_  = A232 & A200;
  assign \new_[69928]_  = \new_[69927]_  & \new_[69924]_ ;
  assign \new_[69929]_  = \new_[69928]_  & \new_[69921]_ ;
  assign \new_[69933]_  = A235 & A234;
  assign \new_[69934]_  = ~A233 & \new_[69933]_ ;
  assign \new_[69937]_  = ~A299 & A298;
  assign \new_[69940]_  = A301 & A300;
  assign \new_[69941]_  = \new_[69940]_  & \new_[69937]_ ;
  assign \new_[69942]_  = \new_[69941]_  & \new_[69934]_ ;
  assign \new_[69946]_  = ~A167 & ~A168;
  assign \new_[69947]_  = A169 & \new_[69946]_ ;
  assign \new_[69950]_  = ~A199 & A166;
  assign \new_[69953]_  = A232 & A200;
  assign \new_[69954]_  = \new_[69953]_  & \new_[69950]_ ;
  assign \new_[69955]_  = \new_[69954]_  & \new_[69947]_ ;
  assign \new_[69959]_  = A235 & A234;
  assign \new_[69960]_  = ~A233 & \new_[69959]_ ;
  assign \new_[69963]_  = ~A299 & A298;
  assign \new_[69966]_  = A302 & A300;
  assign \new_[69967]_  = \new_[69966]_  & \new_[69963]_ ;
  assign \new_[69968]_  = \new_[69967]_  & \new_[69960]_ ;
  assign \new_[69972]_  = ~A167 & ~A168;
  assign \new_[69973]_  = A169 & \new_[69972]_ ;
  assign \new_[69976]_  = ~A199 & A166;
  assign \new_[69979]_  = A232 & A200;
  assign \new_[69980]_  = \new_[69979]_  & \new_[69976]_ ;
  assign \new_[69981]_  = \new_[69980]_  & \new_[69973]_ ;
  assign \new_[69985]_  = A235 & A234;
  assign \new_[69986]_  = ~A233 & \new_[69985]_ ;
  assign \new_[69989]_  = ~A266 & A265;
  assign \new_[69992]_  = A268 & A267;
  assign \new_[69993]_  = \new_[69992]_  & \new_[69989]_ ;
  assign \new_[69994]_  = \new_[69993]_  & \new_[69986]_ ;
  assign \new_[69998]_  = ~A167 & ~A168;
  assign \new_[69999]_  = A169 & \new_[69998]_ ;
  assign \new_[70002]_  = ~A199 & A166;
  assign \new_[70005]_  = A232 & A200;
  assign \new_[70006]_  = \new_[70005]_  & \new_[70002]_ ;
  assign \new_[70007]_  = \new_[70006]_  & \new_[69999]_ ;
  assign \new_[70011]_  = A235 & A234;
  assign \new_[70012]_  = ~A233 & \new_[70011]_ ;
  assign \new_[70015]_  = ~A266 & A265;
  assign \new_[70018]_  = A269 & A267;
  assign \new_[70019]_  = \new_[70018]_  & \new_[70015]_ ;
  assign \new_[70020]_  = \new_[70019]_  & \new_[70012]_ ;
  assign \new_[70024]_  = ~A167 & ~A168;
  assign \new_[70025]_  = A169 & \new_[70024]_ ;
  assign \new_[70028]_  = ~A199 & A166;
  assign \new_[70031]_  = A232 & A200;
  assign \new_[70032]_  = \new_[70031]_  & \new_[70028]_ ;
  assign \new_[70033]_  = \new_[70032]_  & \new_[70025]_ ;
  assign \new_[70037]_  = A236 & A234;
  assign \new_[70038]_  = ~A233 & \new_[70037]_ ;
  assign \new_[70041]_  = ~A299 & A298;
  assign \new_[70044]_  = A301 & A300;
  assign \new_[70045]_  = \new_[70044]_  & \new_[70041]_ ;
  assign \new_[70046]_  = \new_[70045]_  & \new_[70038]_ ;
  assign \new_[70050]_  = ~A167 & ~A168;
  assign \new_[70051]_  = A169 & \new_[70050]_ ;
  assign \new_[70054]_  = ~A199 & A166;
  assign \new_[70057]_  = A232 & A200;
  assign \new_[70058]_  = \new_[70057]_  & \new_[70054]_ ;
  assign \new_[70059]_  = \new_[70058]_  & \new_[70051]_ ;
  assign \new_[70063]_  = A236 & A234;
  assign \new_[70064]_  = ~A233 & \new_[70063]_ ;
  assign \new_[70067]_  = ~A299 & A298;
  assign \new_[70070]_  = A302 & A300;
  assign \new_[70071]_  = \new_[70070]_  & \new_[70067]_ ;
  assign \new_[70072]_  = \new_[70071]_  & \new_[70064]_ ;
  assign \new_[70076]_  = ~A167 & ~A168;
  assign \new_[70077]_  = A169 & \new_[70076]_ ;
  assign \new_[70080]_  = ~A199 & A166;
  assign \new_[70083]_  = A232 & A200;
  assign \new_[70084]_  = \new_[70083]_  & \new_[70080]_ ;
  assign \new_[70085]_  = \new_[70084]_  & \new_[70077]_ ;
  assign \new_[70089]_  = A236 & A234;
  assign \new_[70090]_  = ~A233 & \new_[70089]_ ;
  assign \new_[70093]_  = ~A266 & A265;
  assign \new_[70096]_  = A268 & A267;
  assign \new_[70097]_  = \new_[70096]_  & \new_[70093]_ ;
  assign \new_[70098]_  = \new_[70097]_  & \new_[70090]_ ;
  assign \new_[70102]_  = ~A167 & ~A168;
  assign \new_[70103]_  = A169 & \new_[70102]_ ;
  assign \new_[70106]_  = ~A199 & A166;
  assign \new_[70109]_  = A232 & A200;
  assign \new_[70110]_  = \new_[70109]_  & \new_[70106]_ ;
  assign \new_[70111]_  = \new_[70110]_  & \new_[70103]_ ;
  assign \new_[70115]_  = A236 & A234;
  assign \new_[70116]_  = ~A233 & \new_[70115]_ ;
  assign \new_[70119]_  = ~A266 & A265;
  assign \new_[70122]_  = A269 & A267;
  assign \new_[70123]_  = \new_[70122]_  & \new_[70119]_ ;
  assign \new_[70124]_  = \new_[70123]_  & \new_[70116]_ ;
  assign \new_[70128]_  = ~A167 & ~A168;
  assign \new_[70129]_  = A169 & \new_[70128]_ ;
  assign \new_[70132]_  = ~A199 & A166;
  assign \new_[70135]_  = ~A232 & A200;
  assign \new_[70136]_  = \new_[70135]_  & \new_[70132]_ ;
  assign \new_[70137]_  = \new_[70136]_  & \new_[70129]_ ;
  assign \new_[70141]_  = ~A268 & ~A266;
  assign \new_[70142]_  = ~A233 & \new_[70141]_ ;
  assign \new_[70145]_  = A298 & ~A269;
  assign \new_[70148]_  = ~A302 & ~A301;
  assign \new_[70149]_  = \new_[70148]_  & \new_[70145]_ ;
  assign \new_[70150]_  = \new_[70149]_  & \new_[70142]_ ;
  assign \new_[70154]_  = ~A167 & ~A168;
  assign \new_[70155]_  = A169 & \new_[70154]_ ;
  assign \new_[70158]_  = A199 & A166;
  assign \new_[70161]_  = A201 & ~A200;
  assign \new_[70162]_  = \new_[70161]_  & \new_[70158]_ ;
  assign \new_[70163]_  = \new_[70162]_  & \new_[70155]_ ;
  assign \new_[70167]_  = A233 & A232;
  assign \new_[70168]_  = A202 & \new_[70167]_ ;
  assign \new_[70171]_  = ~A267 & A265;
  assign \new_[70174]_  = ~A300 & ~A299;
  assign \new_[70175]_  = \new_[70174]_  & \new_[70171]_ ;
  assign \new_[70176]_  = \new_[70175]_  & \new_[70168]_ ;
  assign \new_[70180]_  = ~A167 & ~A168;
  assign \new_[70181]_  = A169 & \new_[70180]_ ;
  assign \new_[70184]_  = A199 & A166;
  assign \new_[70187]_  = A201 & ~A200;
  assign \new_[70188]_  = \new_[70187]_  & \new_[70184]_ ;
  assign \new_[70189]_  = \new_[70188]_  & \new_[70181]_ ;
  assign \new_[70193]_  = A233 & A232;
  assign \new_[70194]_  = A202 & \new_[70193]_ ;
  assign \new_[70197]_  = ~A267 & A265;
  assign \new_[70200]_  = A299 & A298;
  assign \new_[70201]_  = \new_[70200]_  & \new_[70197]_ ;
  assign \new_[70202]_  = \new_[70201]_  & \new_[70194]_ ;
  assign \new_[70206]_  = ~A167 & ~A168;
  assign \new_[70207]_  = A169 & \new_[70206]_ ;
  assign \new_[70210]_  = A199 & A166;
  assign \new_[70213]_  = A201 & ~A200;
  assign \new_[70214]_  = \new_[70213]_  & \new_[70210]_ ;
  assign \new_[70215]_  = \new_[70214]_  & \new_[70207]_ ;
  assign \new_[70219]_  = A233 & A232;
  assign \new_[70220]_  = A202 & \new_[70219]_ ;
  assign \new_[70223]_  = ~A267 & A265;
  assign \new_[70226]_  = ~A299 & ~A298;
  assign \new_[70227]_  = \new_[70226]_  & \new_[70223]_ ;
  assign \new_[70228]_  = \new_[70227]_  & \new_[70220]_ ;
  assign \new_[70232]_  = ~A167 & ~A168;
  assign \new_[70233]_  = A169 & \new_[70232]_ ;
  assign \new_[70236]_  = A199 & A166;
  assign \new_[70239]_  = A201 & ~A200;
  assign \new_[70240]_  = \new_[70239]_  & \new_[70236]_ ;
  assign \new_[70241]_  = \new_[70240]_  & \new_[70233]_ ;
  assign \new_[70245]_  = A233 & A232;
  assign \new_[70246]_  = A202 & \new_[70245]_ ;
  assign \new_[70249]_  = A266 & A265;
  assign \new_[70252]_  = ~A300 & ~A299;
  assign \new_[70253]_  = \new_[70252]_  & \new_[70249]_ ;
  assign \new_[70254]_  = \new_[70253]_  & \new_[70246]_ ;
  assign \new_[70258]_  = ~A167 & ~A168;
  assign \new_[70259]_  = A169 & \new_[70258]_ ;
  assign \new_[70262]_  = A199 & A166;
  assign \new_[70265]_  = A201 & ~A200;
  assign \new_[70266]_  = \new_[70265]_  & \new_[70262]_ ;
  assign \new_[70267]_  = \new_[70266]_  & \new_[70259]_ ;
  assign \new_[70271]_  = A233 & A232;
  assign \new_[70272]_  = A202 & \new_[70271]_ ;
  assign \new_[70275]_  = A266 & A265;
  assign \new_[70278]_  = A299 & A298;
  assign \new_[70279]_  = \new_[70278]_  & \new_[70275]_ ;
  assign \new_[70280]_  = \new_[70279]_  & \new_[70272]_ ;
  assign \new_[70284]_  = ~A167 & ~A168;
  assign \new_[70285]_  = A169 & \new_[70284]_ ;
  assign \new_[70288]_  = A199 & A166;
  assign \new_[70291]_  = A201 & ~A200;
  assign \new_[70292]_  = \new_[70291]_  & \new_[70288]_ ;
  assign \new_[70293]_  = \new_[70292]_  & \new_[70285]_ ;
  assign \new_[70297]_  = A233 & A232;
  assign \new_[70298]_  = A202 & \new_[70297]_ ;
  assign \new_[70301]_  = A266 & A265;
  assign \new_[70304]_  = ~A299 & ~A298;
  assign \new_[70305]_  = \new_[70304]_  & \new_[70301]_ ;
  assign \new_[70306]_  = \new_[70305]_  & \new_[70298]_ ;
  assign \new_[70310]_  = ~A167 & ~A168;
  assign \new_[70311]_  = A169 & \new_[70310]_ ;
  assign \new_[70314]_  = A199 & A166;
  assign \new_[70317]_  = A201 & ~A200;
  assign \new_[70318]_  = \new_[70317]_  & \new_[70314]_ ;
  assign \new_[70319]_  = \new_[70318]_  & \new_[70311]_ ;
  assign \new_[70323]_  = A233 & A232;
  assign \new_[70324]_  = A202 & \new_[70323]_ ;
  assign \new_[70327]_  = ~A266 & ~A265;
  assign \new_[70330]_  = ~A300 & ~A299;
  assign \new_[70331]_  = \new_[70330]_  & \new_[70327]_ ;
  assign \new_[70332]_  = \new_[70331]_  & \new_[70324]_ ;
  assign \new_[70336]_  = ~A167 & ~A168;
  assign \new_[70337]_  = A169 & \new_[70336]_ ;
  assign \new_[70340]_  = A199 & A166;
  assign \new_[70343]_  = A201 & ~A200;
  assign \new_[70344]_  = \new_[70343]_  & \new_[70340]_ ;
  assign \new_[70345]_  = \new_[70344]_  & \new_[70337]_ ;
  assign \new_[70349]_  = A233 & A232;
  assign \new_[70350]_  = A202 & \new_[70349]_ ;
  assign \new_[70353]_  = ~A266 & ~A265;
  assign \new_[70356]_  = A299 & A298;
  assign \new_[70357]_  = \new_[70356]_  & \new_[70353]_ ;
  assign \new_[70358]_  = \new_[70357]_  & \new_[70350]_ ;
  assign \new_[70362]_  = ~A167 & ~A168;
  assign \new_[70363]_  = A169 & \new_[70362]_ ;
  assign \new_[70366]_  = A199 & A166;
  assign \new_[70369]_  = A201 & ~A200;
  assign \new_[70370]_  = \new_[70369]_  & \new_[70366]_ ;
  assign \new_[70371]_  = \new_[70370]_  & \new_[70363]_ ;
  assign \new_[70375]_  = A233 & A232;
  assign \new_[70376]_  = A202 & \new_[70375]_ ;
  assign \new_[70379]_  = ~A266 & ~A265;
  assign \new_[70382]_  = ~A299 & ~A298;
  assign \new_[70383]_  = \new_[70382]_  & \new_[70379]_ ;
  assign \new_[70384]_  = \new_[70383]_  & \new_[70376]_ ;
  assign \new_[70388]_  = ~A167 & ~A168;
  assign \new_[70389]_  = A169 & \new_[70388]_ ;
  assign \new_[70392]_  = A199 & A166;
  assign \new_[70395]_  = A201 & ~A200;
  assign \new_[70396]_  = \new_[70395]_  & \new_[70392]_ ;
  assign \new_[70397]_  = \new_[70396]_  & \new_[70389]_ ;
  assign \new_[70401]_  = A233 & ~A232;
  assign \new_[70402]_  = A202 & \new_[70401]_ ;
  assign \new_[70405]_  = ~A299 & A298;
  assign \new_[70408]_  = A301 & A300;
  assign \new_[70409]_  = \new_[70408]_  & \new_[70405]_ ;
  assign \new_[70410]_  = \new_[70409]_  & \new_[70402]_ ;
  assign \new_[70414]_  = ~A167 & ~A168;
  assign \new_[70415]_  = A169 & \new_[70414]_ ;
  assign \new_[70418]_  = A199 & A166;
  assign \new_[70421]_  = A201 & ~A200;
  assign \new_[70422]_  = \new_[70421]_  & \new_[70418]_ ;
  assign \new_[70423]_  = \new_[70422]_  & \new_[70415]_ ;
  assign \new_[70427]_  = A233 & ~A232;
  assign \new_[70428]_  = A202 & \new_[70427]_ ;
  assign \new_[70431]_  = ~A299 & A298;
  assign \new_[70434]_  = A302 & A300;
  assign \new_[70435]_  = \new_[70434]_  & \new_[70431]_ ;
  assign \new_[70436]_  = \new_[70435]_  & \new_[70428]_ ;
  assign \new_[70440]_  = ~A167 & ~A168;
  assign \new_[70441]_  = A169 & \new_[70440]_ ;
  assign \new_[70444]_  = A199 & A166;
  assign \new_[70447]_  = A201 & ~A200;
  assign \new_[70448]_  = \new_[70447]_  & \new_[70444]_ ;
  assign \new_[70449]_  = \new_[70448]_  & \new_[70441]_ ;
  assign \new_[70453]_  = A233 & ~A232;
  assign \new_[70454]_  = A202 & \new_[70453]_ ;
  assign \new_[70457]_  = ~A266 & A265;
  assign \new_[70460]_  = A268 & A267;
  assign \new_[70461]_  = \new_[70460]_  & \new_[70457]_ ;
  assign \new_[70462]_  = \new_[70461]_  & \new_[70454]_ ;
  assign \new_[70466]_  = ~A167 & ~A168;
  assign \new_[70467]_  = A169 & \new_[70466]_ ;
  assign \new_[70470]_  = A199 & A166;
  assign \new_[70473]_  = A201 & ~A200;
  assign \new_[70474]_  = \new_[70473]_  & \new_[70470]_ ;
  assign \new_[70475]_  = \new_[70474]_  & \new_[70467]_ ;
  assign \new_[70479]_  = A233 & ~A232;
  assign \new_[70480]_  = A202 & \new_[70479]_ ;
  assign \new_[70483]_  = ~A266 & A265;
  assign \new_[70486]_  = A269 & A267;
  assign \new_[70487]_  = \new_[70486]_  & \new_[70483]_ ;
  assign \new_[70488]_  = \new_[70487]_  & \new_[70480]_ ;
  assign \new_[70492]_  = ~A167 & ~A168;
  assign \new_[70493]_  = A169 & \new_[70492]_ ;
  assign \new_[70496]_  = A199 & A166;
  assign \new_[70499]_  = A201 & ~A200;
  assign \new_[70500]_  = \new_[70499]_  & \new_[70496]_ ;
  assign \new_[70501]_  = \new_[70500]_  & \new_[70493]_ ;
  assign \new_[70505]_  = ~A234 & ~A233;
  assign \new_[70506]_  = A202 & \new_[70505]_ ;
  assign \new_[70509]_  = A266 & A265;
  assign \new_[70512]_  = ~A300 & A298;
  assign \new_[70513]_  = \new_[70512]_  & \new_[70509]_ ;
  assign \new_[70514]_  = \new_[70513]_  & \new_[70506]_ ;
  assign \new_[70518]_  = ~A167 & ~A168;
  assign \new_[70519]_  = A169 & \new_[70518]_ ;
  assign \new_[70522]_  = A199 & A166;
  assign \new_[70525]_  = A201 & ~A200;
  assign \new_[70526]_  = \new_[70525]_  & \new_[70522]_ ;
  assign \new_[70527]_  = \new_[70526]_  & \new_[70519]_ ;
  assign \new_[70531]_  = ~A234 & ~A233;
  assign \new_[70532]_  = A202 & \new_[70531]_ ;
  assign \new_[70535]_  = A266 & A265;
  assign \new_[70538]_  = A299 & A298;
  assign \new_[70539]_  = \new_[70538]_  & \new_[70535]_ ;
  assign \new_[70540]_  = \new_[70539]_  & \new_[70532]_ ;
  assign \new_[70544]_  = ~A167 & ~A168;
  assign \new_[70545]_  = A169 & \new_[70544]_ ;
  assign \new_[70548]_  = A199 & A166;
  assign \new_[70551]_  = A201 & ~A200;
  assign \new_[70552]_  = \new_[70551]_  & \new_[70548]_ ;
  assign \new_[70553]_  = \new_[70552]_  & \new_[70545]_ ;
  assign \new_[70557]_  = ~A234 & ~A233;
  assign \new_[70558]_  = A202 & \new_[70557]_ ;
  assign \new_[70561]_  = A266 & A265;
  assign \new_[70564]_  = ~A299 & ~A298;
  assign \new_[70565]_  = \new_[70564]_  & \new_[70561]_ ;
  assign \new_[70566]_  = \new_[70565]_  & \new_[70558]_ ;
  assign \new_[70570]_  = ~A167 & ~A168;
  assign \new_[70571]_  = A169 & \new_[70570]_ ;
  assign \new_[70574]_  = A199 & A166;
  assign \new_[70577]_  = A201 & ~A200;
  assign \new_[70578]_  = \new_[70577]_  & \new_[70574]_ ;
  assign \new_[70579]_  = \new_[70578]_  & \new_[70571]_ ;
  assign \new_[70583]_  = ~A234 & ~A233;
  assign \new_[70584]_  = A202 & \new_[70583]_ ;
  assign \new_[70587]_  = ~A267 & ~A266;
  assign \new_[70590]_  = ~A300 & A298;
  assign \new_[70591]_  = \new_[70590]_  & \new_[70587]_ ;
  assign \new_[70592]_  = \new_[70591]_  & \new_[70584]_ ;
  assign \new_[70596]_  = ~A167 & ~A168;
  assign \new_[70597]_  = A169 & \new_[70596]_ ;
  assign \new_[70600]_  = A199 & A166;
  assign \new_[70603]_  = A201 & ~A200;
  assign \new_[70604]_  = \new_[70603]_  & \new_[70600]_ ;
  assign \new_[70605]_  = \new_[70604]_  & \new_[70597]_ ;
  assign \new_[70609]_  = ~A234 & ~A233;
  assign \new_[70610]_  = A202 & \new_[70609]_ ;
  assign \new_[70613]_  = ~A267 & ~A266;
  assign \new_[70616]_  = A299 & A298;
  assign \new_[70617]_  = \new_[70616]_  & \new_[70613]_ ;
  assign \new_[70618]_  = \new_[70617]_  & \new_[70610]_ ;
  assign \new_[70622]_  = ~A167 & ~A168;
  assign \new_[70623]_  = A169 & \new_[70622]_ ;
  assign \new_[70626]_  = A199 & A166;
  assign \new_[70629]_  = A201 & ~A200;
  assign \new_[70630]_  = \new_[70629]_  & \new_[70626]_ ;
  assign \new_[70631]_  = \new_[70630]_  & \new_[70623]_ ;
  assign \new_[70635]_  = ~A234 & ~A233;
  assign \new_[70636]_  = A202 & \new_[70635]_ ;
  assign \new_[70639]_  = ~A267 & ~A266;
  assign \new_[70642]_  = ~A299 & ~A298;
  assign \new_[70643]_  = \new_[70642]_  & \new_[70639]_ ;
  assign \new_[70644]_  = \new_[70643]_  & \new_[70636]_ ;
  assign \new_[70648]_  = ~A167 & ~A168;
  assign \new_[70649]_  = A169 & \new_[70648]_ ;
  assign \new_[70652]_  = A199 & A166;
  assign \new_[70655]_  = A201 & ~A200;
  assign \new_[70656]_  = \new_[70655]_  & \new_[70652]_ ;
  assign \new_[70657]_  = \new_[70656]_  & \new_[70649]_ ;
  assign \new_[70661]_  = ~A234 & ~A233;
  assign \new_[70662]_  = A202 & \new_[70661]_ ;
  assign \new_[70665]_  = ~A266 & ~A265;
  assign \new_[70668]_  = ~A300 & A298;
  assign \new_[70669]_  = \new_[70668]_  & \new_[70665]_ ;
  assign \new_[70670]_  = \new_[70669]_  & \new_[70662]_ ;
  assign \new_[70674]_  = ~A167 & ~A168;
  assign \new_[70675]_  = A169 & \new_[70674]_ ;
  assign \new_[70678]_  = A199 & A166;
  assign \new_[70681]_  = A201 & ~A200;
  assign \new_[70682]_  = \new_[70681]_  & \new_[70678]_ ;
  assign \new_[70683]_  = \new_[70682]_  & \new_[70675]_ ;
  assign \new_[70687]_  = ~A234 & ~A233;
  assign \new_[70688]_  = A202 & \new_[70687]_ ;
  assign \new_[70691]_  = ~A266 & ~A265;
  assign \new_[70694]_  = A299 & A298;
  assign \new_[70695]_  = \new_[70694]_  & \new_[70691]_ ;
  assign \new_[70696]_  = \new_[70695]_  & \new_[70688]_ ;
  assign \new_[70700]_  = ~A167 & ~A168;
  assign \new_[70701]_  = A169 & \new_[70700]_ ;
  assign \new_[70704]_  = A199 & A166;
  assign \new_[70707]_  = A201 & ~A200;
  assign \new_[70708]_  = \new_[70707]_  & \new_[70704]_ ;
  assign \new_[70709]_  = \new_[70708]_  & \new_[70701]_ ;
  assign \new_[70713]_  = ~A234 & ~A233;
  assign \new_[70714]_  = A202 & \new_[70713]_ ;
  assign \new_[70717]_  = ~A266 & ~A265;
  assign \new_[70720]_  = ~A299 & ~A298;
  assign \new_[70721]_  = \new_[70720]_  & \new_[70717]_ ;
  assign \new_[70722]_  = \new_[70721]_  & \new_[70714]_ ;
  assign \new_[70726]_  = ~A167 & ~A168;
  assign \new_[70727]_  = A169 & \new_[70726]_ ;
  assign \new_[70730]_  = A199 & A166;
  assign \new_[70733]_  = A201 & ~A200;
  assign \new_[70734]_  = \new_[70733]_  & \new_[70730]_ ;
  assign \new_[70735]_  = \new_[70734]_  & \new_[70727]_ ;
  assign \new_[70739]_  = ~A233 & A232;
  assign \new_[70740]_  = A202 & \new_[70739]_ ;
  assign \new_[70743]_  = A235 & A234;
  assign \new_[70746]_  = A299 & ~A298;
  assign \new_[70747]_  = \new_[70746]_  & \new_[70743]_ ;
  assign \new_[70748]_  = \new_[70747]_  & \new_[70740]_ ;
  assign \new_[70752]_  = ~A167 & ~A168;
  assign \new_[70753]_  = A169 & \new_[70752]_ ;
  assign \new_[70756]_  = A199 & A166;
  assign \new_[70759]_  = A201 & ~A200;
  assign \new_[70760]_  = \new_[70759]_  & \new_[70756]_ ;
  assign \new_[70761]_  = \new_[70760]_  & \new_[70753]_ ;
  assign \new_[70765]_  = ~A233 & A232;
  assign \new_[70766]_  = A202 & \new_[70765]_ ;
  assign \new_[70769]_  = A235 & A234;
  assign \new_[70772]_  = A266 & ~A265;
  assign \new_[70773]_  = \new_[70772]_  & \new_[70769]_ ;
  assign \new_[70774]_  = \new_[70773]_  & \new_[70766]_ ;
  assign \new_[70778]_  = ~A167 & ~A168;
  assign \new_[70779]_  = A169 & \new_[70778]_ ;
  assign \new_[70782]_  = A199 & A166;
  assign \new_[70785]_  = A201 & ~A200;
  assign \new_[70786]_  = \new_[70785]_  & \new_[70782]_ ;
  assign \new_[70787]_  = \new_[70786]_  & \new_[70779]_ ;
  assign \new_[70791]_  = ~A233 & A232;
  assign \new_[70792]_  = A202 & \new_[70791]_ ;
  assign \new_[70795]_  = A236 & A234;
  assign \new_[70798]_  = A299 & ~A298;
  assign \new_[70799]_  = \new_[70798]_  & \new_[70795]_ ;
  assign \new_[70800]_  = \new_[70799]_  & \new_[70792]_ ;
  assign \new_[70804]_  = ~A167 & ~A168;
  assign \new_[70805]_  = A169 & \new_[70804]_ ;
  assign \new_[70808]_  = A199 & A166;
  assign \new_[70811]_  = A201 & ~A200;
  assign \new_[70812]_  = \new_[70811]_  & \new_[70808]_ ;
  assign \new_[70813]_  = \new_[70812]_  & \new_[70805]_ ;
  assign \new_[70817]_  = ~A233 & A232;
  assign \new_[70818]_  = A202 & \new_[70817]_ ;
  assign \new_[70821]_  = A236 & A234;
  assign \new_[70824]_  = A266 & ~A265;
  assign \new_[70825]_  = \new_[70824]_  & \new_[70821]_ ;
  assign \new_[70826]_  = \new_[70825]_  & \new_[70818]_ ;
  assign \new_[70830]_  = ~A167 & ~A168;
  assign \new_[70831]_  = A169 & \new_[70830]_ ;
  assign \new_[70834]_  = A199 & A166;
  assign \new_[70837]_  = A201 & ~A200;
  assign \new_[70838]_  = \new_[70837]_  & \new_[70834]_ ;
  assign \new_[70839]_  = \new_[70838]_  & \new_[70831]_ ;
  assign \new_[70843]_  = ~A233 & ~A232;
  assign \new_[70844]_  = A202 & \new_[70843]_ ;
  assign \new_[70847]_  = A266 & A265;
  assign \new_[70850]_  = ~A300 & A298;
  assign \new_[70851]_  = \new_[70850]_  & \new_[70847]_ ;
  assign \new_[70852]_  = \new_[70851]_  & \new_[70844]_ ;
  assign \new_[70856]_  = ~A167 & ~A168;
  assign \new_[70857]_  = A169 & \new_[70856]_ ;
  assign \new_[70860]_  = A199 & A166;
  assign \new_[70863]_  = A201 & ~A200;
  assign \new_[70864]_  = \new_[70863]_  & \new_[70860]_ ;
  assign \new_[70865]_  = \new_[70864]_  & \new_[70857]_ ;
  assign \new_[70869]_  = ~A233 & ~A232;
  assign \new_[70870]_  = A202 & \new_[70869]_ ;
  assign \new_[70873]_  = A266 & A265;
  assign \new_[70876]_  = A299 & A298;
  assign \new_[70877]_  = \new_[70876]_  & \new_[70873]_ ;
  assign \new_[70878]_  = \new_[70877]_  & \new_[70870]_ ;
  assign \new_[70882]_  = ~A167 & ~A168;
  assign \new_[70883]_  = A169 & \new_[70882]_ ;
  assign \new_[70886]_  = A199 & A166;
  assign \new_[70889]_  = A201 & ~A200;
  assign \new_[70890]_  = \new_[70889]_  & \new_[70886]_ ;
  assign \new_[70891]_  = \new_[70890]_  & \new_[70883]_ ;
  assign \new_[70895]_  = ~A233 & ~A232;
  assign \new_[70896]_  = A202 & \new_[70895]_ ;
  assign \new_[70899]_  = A266 & A265;
  assign \new_[70902]_  = ~A299 & ~A298;
  assign \new_[70903]_  = \new_[70902]_  & \new_[70899]_ ;
  assign \new_[70904]_  = \new_[70903]_  & \new_[70896]_ ;
  assign \new_[70908]_  = ~A167 & ~A168;
  assign \new_[70909]_  = A169 & \new_[70908]_ ;
  assign \new_[70912]_  = A199 & A166;
  assign \new_[70915]_  = A201 & ~A200;
  assign \new_[70916]_  = \new_[70915]_  & \new_[70912]_ ;
  assign \new_[70917]_  = \new_[70916]_  & \new_[70909]_ ;
  assign \new_[70921]_  = ~A233 & ~A232;
  assign \new_[70922]_  = A202 & \new_[70921]_ ;
  assign \new_[70925]_  = ~A267 & ~A266;
  assign \new_[70928]_  = ~A300 & A298;
  assign \new_[70929]_  = \new_[70928]_  & \new_[70925]_ ;
  assign \new_[70930]_  = \new_[70929]_  & \new_[70922]_ ;
  assign \new_[70934]_  = ~A167 & ~A168;
  assign \new_[70935]_  = A169 & \new_[70934]_ ;
  assign \new_[70938]_  = A199 & A166;
  assign \new_[70941]_  = A201 & ~A200;
  assign \new_[70942]_  = \new_[70941]_  & \new_[70938]_ ;
  assign \new_[70943]_  = \new_[70942]_  & \new_[70935]_ ;
  assign \new_[70947]_  = ~A233 & ~A232;
  assign \new_[70948]_  = A202 & \new_[70947]_ ;
  assign \new_[70951]_  = ~A267 & ~A266;
  assign \new_[70954]_  = A299 & A298;
  assign \new_[70955]_  = \new_[70954]_  & \new_[70951]_ ;
  assign \new_[70956]_  = \new_[70955]_  & \new_[70948]_ ;
  assign \new_[70960]_  = ~A167 & ~A168;
  assign \new_[70961]_  = A169 & \new_[70960]_ ;
  assign \new_[70964]_  = A199 & A166;
  assign \new_[70967]_  = A201 & ~A200;
  assign \new_[70968]_  = \new_[70967]_  & \new_[70964]_ ;
  assign \new_[70969]_  = \new_[70968]_  & \new_[70961]_ ;
  assign \new_[70973]_  = ~A233 & ~A232;
  assign \new_[70974]_  = A202 & \new_[70973]_ ;
  assign \new_[70977]_  = ~A267 & ~A266;
  assign \new_[70980]_  = ~A299 & ~A298;
  assign \new_[70981]_  = \new_[70980]_  & \new_[70977]_ ;
  assign \new_[70982]_  = \new_[70981]_  & \new_[70974]_ ;
  assign \new_[70986]_  = ~A167 & ~A168;
  assign \new_[70987]_  = A169 & \new_[70986]_ ;
  assign \new_[70990]_  = A199 & A166;
  assign \new_[70993]_  = A201 & ~A200;
  assign \new_[70994]_  = \new_[70993]_  & \new_[70990]_ ;
  assign \new_[70995]_  = \new_[70994]_  & \new_[70987]_ ;
  assign \new_[70999]_  = ~A233 & ~A232;
  assign \new_[71000]_  = A202 & \new_[70999]_ ;
  assign \new_[71003]_  = ~A266 & ~A265;
  assign \new_[71006]_  = ~A300 & A298;
  assign \new_[71007]_  = \new_[71006]_  & \new_[71003]_ ;
  assign \new_[71008]_  = \new_[71007]_  & \new_[71000]_ ;
  assign \new_[71012]_  = ~A167 & ~A168;
  assign \new_[71013]_  = A169 & \new_[71012]_ ;
  assign \new_[71016]_  = A199 & A166;
  assign \new_[71019]_  = A201 & ~A200;
  assign \new_[71020]_  = \new_[71019]_  & \new_[71016]_ ;
  assign \new_[71021]_  = \new_[71020]_  & \new_[71013]_ ;
  assign \new_[71025]_  = ~A233 & ~A232;
  assign \new_[71026]_  = A202 & \new_[71025]_ ;
  assign \new_[71029]_  = ~A266 & ~A265;
  assign \new_[71032]_  = A299 & A298;
  assign \new_[71033]_  = \new_[71032]_  & \new_[71029]_ ;
  assign \new_[71034]_  = \new_[71033]_  & \new_[71026]_ ;
  assign \new_[71038]_  = ~A167 & ~A168;
  assign \new_[71039]_  = A169 & \new_[71038]_ ;
  assign \new_[71042]_  = A199 & A166;
  assign \new_[71045]_  = A201 & ~A200;
  assign \new_[71046]_  = \new_[71045]_  & \new_[71042]_ ;
  assign \new_[71047]_  = \new_[71046]_  & \new_[71039]_ ;
  assign \new_[71051]_  = ~A233 & ~A232;
  assign \new_[71052]_  = A202 & \new_[71051]_ ;
  assign \new_[71055]_  = ~A266 & ~A265;
  assign \new_[71058]_  = ~A299 & ~A298;
  assign \new_[71059]_  = \new_[71058]_  & \new_[71055]_ ;
  assign \new_[71060]_  = \new_[71059]_  & \new_[71052]_ ;
  assign \new_[71064]_  = ~A167 & ~A168;
  assign \new_[71065]_  = A169 & \new_[71064]_ ;
  assign \new_[71068]_  = A199 & A166;
  assign \new_[71071]_  = A201 & ~A200;
  assign \new_[71072]_  = \new_[71071]_  & \new_[71068]_ ;
  assign \new_[71073]_  = \new_[71072]_  & \new_[71065]_ ;
  assign \new_[71077]_  = A233 & A232;
  assign \new_[71078]_  = A203 & \new_[71077]_ ;
  assign \new_[71081]_  = ~A267 & A265;
  assign \new_[71084]_  = ~A300 & ~A299;
  assign \new_[71085]_  = \new_[71084]_  & \new_[71081]_ ;
  assign \new_[71086]_  = \new_[71085]_  & \new_[71078]_ ;
  assign \new_[71090]_  = ~A167 & ~A168;
  assign \new_[71091]_  = A169 & \new_[71090]_ ;
  assign \new_[71094]_  = A199 & A166;
  assign \new_[71097]_  = A201 & ~A200;
  assign \new_[71098]_  = \new_[71097]_  & \new_[71094]_ ;
  assign \new_[71099]_  = \new_[71098]_  & \new_[71091]_ ;
  assign \new_[71103]_  = A233 & A232;
  assign \new_[71104]_  = A203 & \new_[71103]_ ;
  assign \new_[71107]_  = ~A267 & A265;
  assign \new_[71110]_  = A299 & A298;
  assign \new_[71111]_  = \new_[71110]_  & \new_[71107]_ ;
  assign \new_[71112]_  = \new_[71111]_  & \new_[71104]_ ;
  assign \new_[71116]_  = ~A167 & ~A168;
  assign \new_[71117]_  = A169 & \new_[71116]_ ;
  assign \new_[71120]_  = A199 & A166;
  assign \new_[71123]_  = A201 & ~A200;
  assign \new_[71124]_  = \new_[71123]_  & \new_[71120]_ ;
  assign \new_[71125]_  = \new_[71124]_  & \new_[71117]_ ;
  assign \new_[71129]_  = A233 & A232;
  assign \new_[71130]_  = A203 & \new_[71129]_ ;
  assign \new_[71133]_  = ~A267 & A265;
  assign \new_[71136]_  = ~A299 & ~A298;
  assign \new_[71137]_  = \new_[71136]_  & \new_[71133]_ ;
  assign \new_[71138]_  = \new_[71137]_  & \new_[71130]_ ;
  assign \new_[71142]_  = ~A167 & ~A168;
  assign \new_[71143]_  = A169 & \new_[71142]_ ;
  assign \new_[71146]_  = A199 & A166;
  assign \new_[71149]_  = A201 & ~A200;
  assign \new_[71150]_  = \new_[71149]_  & \new_[71146]_ ;
  assign \new_[71151]_  = \new_[71150]_  & \new_[71143]_ ;
  assign \new_[71155]_  = A233 & A232;
  assign \new_[71156]_  = A203 & \new_[71155]_ ;
  assign \new_[71159]_  = A266 & A265;
  assign \new_[71162]_  = ~A300 & ~A299;
  assign \new_[71163]_  = \new_[71162]_  & \new_[71159]_ ;
  assign \new_[71164]_  = \new_[71163]_  & \new_[71156]_ ;
  assign \new_[71168]_  = ~A167 & ~A168;
  assign \new_[71169]_  = A169 & \new_[71168]_ ;
  assign \new_[71172]_  = A199 & A166;
  assign \new_[71175]_  = A201 & ~A200;
  assign \new_[71176]_  = \new_[71175]_  & \new_[71172]_ ;
  assign \new_[71177]_  = \new_[71176]_  & \new_[71169]_ ;
  assign \new_[71181]_  = A233 & A232;
  assign \new_[71182]_  = A203 & \new_[71181]_ ;
  assign \new_[71185]_  = A266 & A265;
  assign \new_[71188]_  = A299 & A298;
  assign \new_[71189]_  = \new_[71188]_  & \new_[71185]_ ;
  assign \new_[71190]_  = \new_[71189]_  & \new_[71182]_ ;
  assign \new_[71194]_  = ~A167 & ~A168;
  assign \new_[71195]_  = A169 & \new_[71194]_ ;
  assign \new_[71198]_  = A199 & A166;
  assign \new_[71201]_  = A201 & ~A200;
  assign \new_[71202]_  = \new_[71201]_  & \new_[71198]_ ;
  assign \new_[71203]_  = \new_[71202]_  & \new_[71195]_ ;
  assign \new_[71207]_  = A233 & A232;
  assign \new_[71208]_  = A203 & \new_[71207]_ ;
  assign \new_[71211]_  = A266 & A265;
  assign \new_[71214]_  = ~A299 & ~A298;
  assign \new_[71215]_  = \new_[71214]_  & \new_[71211]_ ;
  assign \new_[71216]_  = \new_[71215]_  & \new_[71208]_ ;
  assign \new_[71220]_  = ~A167 & ~A168;
  assign \new_[71221]_  = A169 & \new_[71220]_ ;
  assign \new_[71224]_  = A199 & A166;
  assign \new_[71227]_  = A201 & ~A200;
  assign \new_[71228]_  = \new_[71227]_  & \new_[71224]_ ;
  assign \new_[71229]_  = \new_[71228]_  & \new_[71221]_ ;
  assign \new_[71233]_  = A233 & A232;
  assign \new_[71234]_  = A203 & \new_[71233]_ ;
  assign \new_[71237]_  = ~A266 & ~A265;
  assign \new_[71240]_  = ~A300 & ~A299;
  assign \new_[71241]_  = \new_[71240]_  & \new_[71237]_ ;
  assign \new_[71242]_  = \new_[71241]_  & \new_[71234]_ ;
  assign \new_[71246]_  = ~A167 & ~A168;
  assign \new_[71247]_  = A169 & \new_[71246]_ ;
  assign \new_[71250]_  = A199 & A166;
  assign \new_[71253]_  = A201 & ~A200;
  assign \new_[71254]_  = \new_[71253]_  & \new_[71250]_ ;
  assign \new_[71255]_  = \new_[71254]_  & \new_[71247]_ ;
  assign \new_[71259]_  = A233 & A232;
  assign \new_[71260]_  = A203 & \new_[71259]_ ;
  assign \new_[71263]_  = ~A266 & ~A265;
  assign \new_[71266]_  = A299 & A298;
  assign \new_[71267]_  = \new_[71266]_  & \new_[71263]_ ;
  assign \new_[71268]_  = \new_[71267]_  & \new_[71260]_ ;
  assign \new_[71272]_  = ~A167 & ~A168;
  assign \new_[71273]_  = A169 & \new_[71272]_ ;
  assign \new_[71276]_  = A199 & A166;
  assign \new_[71279]_  = A201 & ~A200;
  assign \new_[71280]_  = \new_[71279]_  & \new_[71276]_ ;
  assign \new_[71281]_  = \new_[71280]_  & \new_[71273]_ ;
  assign \new_[71285]_  = A233 & A232;
  assign \new_[71286]_  = A203 & \new_[71285]_ ;
  assign \new_[71289]_  = ~A266 & ~A265;
  assign \new_[71292]_  = ~A299 & ~A298;
  assign \new_[71293]_  = \new_[71292]_  & \new_[71289]_ ;
  assign \new_[71294]_  = \new_[71293]_  & \new_[71286]_ ;
  assign \new_[71298]_  = ~A167 & ~A168;
  assign \new_[71299]_  = A169 & \new_[71298]_ ;
  assign \new_[71302]_  = A199 & A166;
  assign \new_[71305]_  = A201 & ~A200;
  assign \new_[71306]_  = \new_[71305]_  & \new_[71302]_ ;
  assign \new_[71307]_  = \new_[71306]_  & \new_[71299]_ ;
  assign \new_[71311]_  = A233 & ~A232;
  assign \new_[71312]_  = A203 & \new_[71311]_ ;
  assign \new_[71315]_  = ~A299 & A298;
  assign \new_[71318]_  = A301 & A300;
  assign \new_[71319]_  = \new_[71318]_  & \new_[71315]_ ;
  assign \new_[71320]_  = \new_[71319]_  & \new_[71312]_ ;
  assign \new_[71324]_  = ~A167 & ~A168;
  assign \new_[71325]_  = A169 & \new_[71324]_ ;
  assign \new_[71328]_  = A199 & A166;
  assign \new_[71331]_  = A201 & ~A200;
  assign \new_[71332]_  = \new_[71331]_  & \new_[71328]_ ;
  assign \new_[71333]_  = \new_[71332]_  & \new_[71325]_ ;
  assign \new_[71337]_  = A233 & ~A232;
  assign \new_[71338]_  = A203 & \new_[71337]_ ;
  assign \new_[71341]_  = ~A299 & A298;
  assign \new_[71344]_  = A302 & A300;
  assign \new_[71345]_  = \new_[71344]_  & \new_[71341]_ ;
  assign \new_[71346]_  = \new_[71345]_  & \new_[71338]_ ;
  assign \new_[71350]_  = ~A167 & ~A168;
  assign \new_[71351]_  = A169 & \new_[71350]_ ;
  assign \new_[71354]_  = A199 & A166;
  assign \new_[71357]_  = A201 & ~A200;
  assign \new_[71358]_  = \new_[71357]_  & \new_[71354]_ ;
  assign \new_[71359]_  = \new_[71358]_  & \new_[71351]_ ;
  assign \new_[71363]_  = A233 & ~A232;
  assign \new_[71364]_  = A203 & \new_[71363]_ ;
  assign \new_[71367]_  = ~A266 & A265;
  assign \new_[71370]_  = A268 & A267;
  assign \new_[71371]_  = \new_[71370]_  & \new_[71367]_ ;
  assign \new_[71372]_  = \new_[71371]_  & \new_[71364]_ ;
  assign \new_[71376]_  = ~A167 & ~A168;
  assign \new_[71377]_  = A169 & \new_[71376]_ ;
  assign \new_[71380]_  = A199 & A166;
  assign \new_[71383]_  = A201 & ~A200;
  assign \new_[71384]_  = \new_[71383]_  & \new_[71380]_ ;
  assign \new_[71385]_  = \new_[71384]_  & \new_[71377]_ ;
  assign \new_[71389]_  = A233 & ~A232;
  assign \new_[71390]_  = A203 & \new_[71389]_ ;
  assign \new_[71393]_  = ~A266 & A265;
  assign \new_[71396]_  = A269 & A267;
  assign \new_[71397]_  = \new_[71396]_  & \new_[71393]_ ;
  assign \new_[71398]_  = \new_[71397]_  & \new_[71390]_ ;
  assign \new_[71402]_  = ~A167 & ~A168;
  assign \new_[71403]_  = A169 & \new_[71402]_ ;
  assign \new_[71406]_  = A199 & A166;
  assign \new_[71409]_  = A201 & ~A200;
  assign \new_[71410]_  = \new_[71409]_  & \new_[71406]_ ;
  assign \new_[71411]_  = \new_[71410]_  & \new_[71403]_ ;
  assign \new_[71415]_  = ~A234 & ~A233;
  assign \new_[71416]_  = A203 & \new_[71415]_ ;
  assign \new_[71419]_  = A266 & A265;
  assign \new_[71422]_  = ~A300 & A298;
  assign \new_[71423]_  = \new_[71422]_  & \new_[71419]_ ;
  assign \new_[71424]_  = \new_[71423]_  & \new_[71416]_ ;
  assign \new_[71428]_  = ~A167 & ~A168;
  assign \new_[71429]_  = A169 & \new_[71428]_ ;
  assign \new_[71432]_  = A199 & A166;
  assign \new_[71435]_  = A201 & ~A200;
  assign \new_[71436]_  = \new_[71435]_  & \new_[71432]_ ;
  assign \new_[71437]_  = \new_[71436]_  & \new_[71429]_ ;
  assign \new_[71441]_  = ~A234 & ~A233;
  assign \new_[71442]_  = A203 & \new_[71441]_ ;
  assign \new_[71445]_  = A266 & A265;
  assign \new_[71448]_  = A299 & A298;
  assign \new_[71449]_  = \new_[71448]_  & \new_[71445]_ ;
  assign \new_[71450]_  = \new_[71449]_  & \new_[71442]_ ;
  assign \new_[71454]_  = ~A167 & ~A168;
  assign \new_[71455]_  = A169 & \new_[71454]_ ;
  assign \new_[71458]_  = A199 & A166;
  assign \new_[71461]_  = A201 & ~A200;
  assign \new_[71462]_  = \new_[71461]_  & \new_[71458]_ ;
  assign \new_[71463]_  = \new_[71462]_  & \new_[71455]_ ;
  assign \new_[71467]_  = ~A234 & ~A233;
  assign \new_[71468]_  = A203 & \new_[71467]_ ;
  assign \new_[71471]_  = A266 & A265;
  assign \new_[71474]_  = ~A299 & ~A298;
  assign \new_[71475]_  = \new_[71474]_  & \new_[71471]_ ;
  assign \new_[71476]_  = \new_[71475]_  & \new_[71468]_ ;
  assign \new_[71480]_  = ~A167 & ~A168;
  assign \new_[71481]_  = A169 & \new_[71480]_ ;
  assign \new_[71484]_  = A199 & A166;
  assign \new_[71487]_  = A201 & ~A200;
  assign \new_[71488]_  = \new_[71487]_  & \new_[71484]_ ;
  assign \new_[71489]_  = \new_[71488]_  & \new_[71481]_ ;
  assign \new_[71493]_  = ~A234 & ~A233;
  assign \new_[71494]_  = A203 & \new_[71493]_ ;
  assign \new_[71497]_  = ~A267 & ~A266;
  assign \new_[71500]_  = ~A300 & A298;
  assign \new_[71501]_  = \new_[71500]_  & \new_[71497]_ ;
  assign \new_[71502]_  = \new_[71501]_  & \new_[71494]_ ;
  assign \new_[71506]_  = ~A167 & ~A168;
  assign \new_[71507]_  = A169 & \new_[71506]_ ;
  assign \new_[71510]_  = A199 & A166;
  assign \new_[71513]_  = A201 & ~A200;
  assign \new_[71514]_  = \new_[71513]_  & \new_[71510]_ ;
  assign \new_[71515]_  = \new_[71514]_  & \new_[71507]_ ;
  assign \new_[71519]_  = ~A234 & ~A233;
  assign \new_[71520]_  = A203 & \new_[71519]_ ;
  assign \new_[71523]_  = ~A267 & ~A266;
  assign \new_[71526]_  = A299 & A298;
  assign \new_[71527]_  = \new_[71526]_  & \new_[71523]_ ;
  assign \new_[71528]_  = \new_[71527]_  & \new_[71520]_ ;
  assign \new_[71532]_  = ~A167 & ~A168;
  assign \new_[71533]_  = A169 & \new_[71532]_ ;
  assign \new_[71536]_  = A199 & A166;
  assign \new_[71539]_  = A201 & ~A200;
  assign \new_[71540]_  = \new_[71539]_  & \new_[71536]_ ;
  assign \new_[71541]_  = \new_[71540]_  & \new_[71533]_ ;
  assign \new_[71545]_  = ~A234 & ~A233;
  assign \new_[71546]_  = A203 & \new_[71545]_ ;
  assign \new_[71549]_  = ~A267 & ~A266;
  assign \new_[71552]_  = ~A299 & ~A298;
  assign \new_[71553]_  = \new_[71552]_  & \new_[71549]_ ;
  assign \new_[71554]_  = \new_[71553]_  & \new_[71546]_ ;
  assign \new_[71558]_  = ~A167 & ~A168;
  assign \new_[71559]_  = A169 & \new_[71558]_ ;
  assign \new_[71562]_  = A199 & A166;
  assign \new_[71565]_  = A201 & ~A200;
  assign \new_[71566]_  = \new_[71565]_  & \new_[71562]_ ;
  assign \new_[71567]_  = \new_[71566]_  & \new_[71559]_ ;
  assign \new_[71571]_  = ~A234 & ~A233;
  assign \new_[71572]_  = A203 & \new_[71571]_ ;
  assign \new_[71575]_  = ~A266 & ~A265;
  assign \new_[71578]_  = ~A300 & A298;
  assign \new_[71579]_  = \new_[71578]_  & \new_[71575]_ ;
  assign \new_[71580]_  = \new_[71579]_  & \new_[71572]_ ;
  assign \new_[71584]_  = ~A167 & ~A168;
  assign \new_[71585]_  = A169 & \new_[71584]_ ;
  assign \new_[71588]_  = A199 & A166;
  assign \new_[71591]_  = A201 & ~A200;
  assign \new_[71592]_  = \new_[71591]_  & \new_[71588]_ ;
  assign \new_[71593]_  = \new_[71592]_  & \new_[71585]_ ;
  assign \new_[71597]_  = ~A234 & ~A233;
  assign \new_[71598]_  = A203 & \new_[71597]_ ;
  assign \new_[71601]_  = ~A266 & ~A265;
  assign \new_[71604]_  = A299 & A298;
  assign \new_[71605]_  = \new_[71604]_  & \new_[71601]_ ;
  assign \new_[71606]_  = \new_[71605]_  & \new_[71598]_ ;
  assign \new_[71610]_  = ~A167 & ~A168;
  assign \new_[71611]_  = A169 & \new_[71610]_ ;
  assign \new_[71614]_  = A199 & A166;
  assign \new_[71617]_  = A201 & ~A200;
  assign \new_[71618]_  = \new_[71617]_  & \new_[71614]_ ;
  assign \new_[71619]_  = \new_[71618]_  & \new_[71611]_ ;
  assign \new_[71623]_  = ~A234 & ~A233;
  assign \new_[71624]_  = A203 & \new_[71623]_ ;
  assign \new_[71627]_  = ~A266 & ~A265;
  assign \new_[71630]_  = ~A299 & ~A298;
  assign \new_[71631]_  = \new_[71630]_  & \new_[71627]_ ;
  assign \new_[71632]_  = \new_[71631]_  & \new_[71624]_ ;
  assign \new_[71636]_  = ~A167 & ~A168;
  assign \new_[71637]_  = A169 & \new_[71636]_ ;
  assign \new_[71640]_  = A199 & A166;
  assign \new_[71643]_  = A201 & ~A200;
  assign \new_[71644]_  = \new_[71643]_  & \new_[71640]_ ;
  assign \new_[71645]_  = \new_[71644]_  & \new_[71637]_ ;
  assign \new_[71649]_  = ~A233 & A232;
  assign \new_[71650]_  = A203 & \new_[71649]_ ;
  assign \new_[71653]_  = A235 & A234;
  assign \new_[71656]_  = A299 & ~A298;
  assign \new_[71657]_  = \new_[71656]_  & \new_[71653]_ ;
  assign \new_[71658]_  = \new_[71657]_  & \new_[71650]_ ;
  assign \new_[71662]_  = ~A167 & ~A168;
  assign \new_[71663]_  = A169 & \new_[71662]_ ;
  assign \new_[71666]_  = A199 & A166;
  assign \new_[71669]_  = A201 & ~A200;
  assign \new_[71670]_  = \new_[71669]_  & \new_[71666]_ ;
  assign \new_[71671]_  = \new_[71670]_  & \new_[71663]_ ;
  assign \new_[71675]_  = ~A233 & A232;
  assign \new_[71676]_  = A203 & \new_[71675]_ ;
  assign \new_[71679]_  = A235 & A234;
  assign \new_[71682]_  = A266 & ~A265;
  assign \new_[71683]_  = \new_[71682]_  & \new_[71679]_ ;
  assign \new_[71684]_  = \new_[71683]_  & \new_[71676]_ ;
  assign \new_[71688]_  = ~A167 & ~A168;
  assign \new_[71689]_  = A169 & \new_[71688]_ ;
  assign \new_[71692]_  = A199 & A166;
  assign \new_[71695]_  = A201 & ~A200;
  assign \new_[71696]_  = \new_[71695]_  & \new_[71692]_ ;
  assign \new_[71697]_  = \new_[71696]_  & \new_[71689]_ ;
  assign \new_[71701]_  = ~A233 & A232;
  assign \new_[71702]_  = A203 & \new_[71701]_ ;
  assign \new_[71705]_  = A236 & A234;
  assign \new_[71708]_  = A299 & ~A298;
  assign \new_[71709]_  = \new_[71708]_  & \new_[71705]_ ;
  assign \new_[71710]_  = \new_[71709]_  & \new_[71702]_ ;
  assign \new_[71714]_  = ~A167 & ~A168;
  assign \new_[71715]_  = A169 & \new_[71714]_ ;
  assign \new_[71718]_  = A199 & A166;
  assign \new_[71721]_  = A201 & ~A200;
  assign \new_[71722]_  = \new_[71721]_  & \new_[71718]_ ;
  assign \new_[71723]_  = \new_[71722]_  & \new_[71715]_ ;
  assign \new_[71727]_  = ~A233 & A232;
  assign \new_[71728]_  = A203 & \new_[71727]_ ;
  assign \new_[71731]_  = A236 & A234;
  assign \new_[71734]_  = A266 & ~A265;
  assign \new_[71735]_  = \new_[71734]_  & \new_[71731]_ ;
  assign \new_[71736]_  = \new_[71735]_  & \new_[71728]_ ;
  assign \new_[71740]_  = ~A167 & ~A168;
  assign \new_[71741]_  = A169 & \new_[71740]_ ;
  assign \new_[71744]_  = A199 & A166;
  assign \new_[71747]_  = A201 & ~A200;
  assign \new_[71748]_  = \new_[71747]_  & \new_[71744]_ ;
  assign \new_[71749]_  = \new_[71748]_  & \new_[71741]_ ;
  assign \new_[71753]_  = ~A233 & ~A232;
  assign \new_[71754]_  = A203 & \new_[71753]_ ;
  assign \new_[71757]_  = A266 & A265;
  assign \new_[71760]_  = ~A300 & A298;
  assign \new_[71761]_  = \new_[71760]_  & \new_[71757]_ ;
  assign \new_[71762]_  = \new_[71761]_  & \new_[71754]_ ;
  assign \new_[71766]_  = ~A167 & ~A168;
  assign \new_[71767]_  = A169 & \new_[71766]_ ;
  assign \new_[71770]_  = A199 & A166;
  assign \new_[71773]_  = A201 & ~A200;
  assign \new_[71774]_  = \new_[71773]_  & \new_[71770]_ ;
  assign \new_[71775]_  = \new_[71774]_  & \new_[71767]_ ;
  assign \new_[71779]_  = ~A233 & ~A232;
  assign \new_[71780]_  = A203 & \new_[71779]_ ;
  assign \new_[71783]_  = A266 & A265;
  assign \new_[71786]_  = A299 & A298;
  assign \new_[71787]_  = \new_[71786]_  & \new_[71783]_ ;
  assign \new_[71788]_  = \new_[71787]_  & \new_[71780]_ ;
  assign \new_[71792]_  = ~A167 & ~A168;
  assign \new_[71793]_  = A169 & \new_[71792]_ ;
  assign \new_[71796]_  = A199 & A166;
  assign \new_[71799]_  = A201 & ~A200;
  assign \new_[71800]_  = \new_[71799]_  & \new_[71796]_ ;
  assign \new_[71801]_  = \new_[71800]_  & \new_[71793]_ ;
  assign \new_[71805]_  = ~A233 & ~A232;
  assign \new_[71806]_  = A203 & \new_[71805]_ ;
  assign \new_[71809]_  = A266 & A265;
  assign \new_[71812]_  = ~A299 & ~A298;
  assign \new_[71813]_  = \new_[71812]_  & \new_[71809]_ ;
  assign \new_[71814]_  = \new_[71813]_  & \new_[71806]_ ;
  assign \new_[71818]_  = ~A167 & ~A168;
  assign \new_[71819]_  = A169 & \new_[71818]_ ;
  assign \new_[71822]_  = A199 & A166;
  assign \new_[71825]_  = A201 & ~A200;
  assign \new_[71826]_  = \new_[71825]_  & \new_[71822]_ ;
  assign \new_[71827]_  = \new_[71826]_  & \new_[71819]_ ;
  assign \new_[71831]_  = ~A233 & ~A232;
  assign \new_[71832]_  = A203 & \new_[71831]_ ;
  assign \new_[71835]_  = ~A267 & ~A266;
  assign \new_[71838]_  = ~A300 & A298;
  assign \new_[71839]_  = \new_[71838]_  & \new_[71835]_ ;
  assign \new_[71840]_  = \new_[71839]_  & \new_[71832]_ ;
  assign \new_[71844]_  = ~A167 & ~A168;
  assign \new_[71845]_  = A169 & \new_[71844]_ ;
  assign \new_[71848]_  = A199 & A166;
  assign \new_[71851]_  = A201 & ~A200;
  assign \new_[71852]_  = \new_[71851]_  & \new_[71848]_ ;
  assign \new_[71853]_  = \new_[71852]_  & \new_[71845]_ ;
  assign \new_[71857]_  = ~A233 & ~A232;
  assign \new_[71858]_  = A203 & \new_[71857]_ ;
  assign \new_[71861]_  = ~A267 & ~A266;
  assign \new_[71864]_  = A299 & A298;
  assign \new_[71865]_  = \new_[71864]_  & \new_[71861]_ ;
  assign \new_[71866]_  = \new_[71865]_  & \new_[71858]_ ;
  assign \new_[71870]_  = ~A167 & ~A168;
  assign \new_[71871]_  = A169 & \new_[71870]_ ;
  assign \new_[71874]_  = A199 & A166;
  assign \new_[71877]_  = A201 & ~A200;
  assign \new_[71878]_  = \new_[71877]_  & \new_[71874]_ ;
  assign \new_[71879]_  = \new_[71878]_  & \new_[71871]_ ;
  assign \new_[71883]_  = ~A233 & ~A232;
  assign \new_[71884]_  = A203 & \new_[71883]_ ;
  assign \new_[71887]_  = ~A267 & ~A266;
  assign \new_[71890]_  = ~A299 & ~A298;
  assign \new_[71891]_  = \new_[71890]_  & \new_[71887]_ ;
  assign \new_[71892]_  = \new_[71891]_  & \new_[71884]_ ;
  assign \new_[71896]_  = ~A167 & ~A168;
  assign \new_[71897]_  = A169 & \new_[71896]_ ;
  assign \new_[71900]_  = A199 & A166;
  assign \new_[71903]_  = A201 & ~A200;
  assign \new_[71904]_  = \new_[71903]_  & \new_[71900]_ ;
  assign \new_[71905]_  = \new_[71904]_  & \new_[71897]_ ;
  assign \new_[71909]_  = ~A233 & ~A232;
  assign \new_[71910]_  = A203 & \new_[71909]_ ;
  assign \new_[71913]_  = ~A266 & ~A265;
  assign \new_[71916]_  = ~A300 & A298;
  assign \new_[71917]_  = \new_[71916]_  & \new_[71913]_ ;
  assign \new_[71918]_  = \new_[71917]_  & \new_[71910]_ ;
  assign \new_[71922]_  = ~A167 & ~A168;
  assign \new_[71923]_  = A169 & \new_[71922]_ ;
  assign \new_[71926]_  = A199 & A166;
  assign \new_[71929]_  = A201 & ~A200;
  assign \new_[71930]_  = \new_[71929]_  & \new_[71926]_ ;
  assign \new_[71931]_  = \new_[71930]_  & \new_[71923]_ ;
  assign \new_[71935]_  = ~A233 & ~A232;
  assign \new_[71936]_  = A203 & \new_[71935]_ ;
  assign \new_[71939]_  = ~A266 & ~A265;
  assign \new_[71942]_  = A299 & A298;
  assign \new_[71943]_  = \new_[71942]_  & \new_[71939]_ ;
  assign \new_[71944]_  = \new_[71943]_  & \new_[71936]_ ;
  assign \new_[71948]_  = ~A167 & ~A168;
  assign \new_[71949]_  = A169 & \new_[71948]_ ;
  assign \new_[71952]_  = A199 & A166;
  assign \new_[71955]_  = A201 & ~A200;
  assign \new_[71956]_  = \new_[71955]_  & \new_[71952]_ ;
  assign \new_[71957]_  = \new_[71956]_  & \new_[71949]_ ;
  assign \new_[71961]_  = ~A233 & ~A232;
  assign \new_[71962]_  = A203 & \new_[71961]_ ;
  assign \new_[71965]_  = ~A266 & ~A265;
  assign \new_[71968]_  = ~A299 & ~A298;
  assign \new_[71969]_  = \new_[71968]_  & \new_[71965]_ ;
  assign \new_[71970]_  = \new_[71969]_  & \new_[71962]_ ;
  assign \new_[71974]_  = ~A168 & A169;
  assign \new_[71975]_  = A170 & \new_[71974]_ ;
  assign \new_[71978]_  = ~A200 & A199;
  assign \new_[71981]_  = A202 & A201;
  assign \new_[71982]_  = \new_[71981]_  & \new_[71978]_ ;
  assign \new_[71983]_  = \new_[71982]_  & \new_[71975]_ ;
  assign \new_[71987]_  = A265 & A233;
  assign \new_[71988]_  = A232 & \new_[71987]_ ;
  assign \new_[71991]_  = ~A269 & ~A268;
  assign \new_[71994]_  = ~A300 & ~A299;
  assign \new_[71995]_  = \new_[71994]_  & \new_[71991]_ ;
  assign \new_[71996]_  = \new_[71995]_  & \new_[71988]_ ;
  assign \new_[72000]_  = ~A168 & A169;
  assign \new_[72001]_  = A170 & \new_[72000]_ ;
  assign \new_[72004]_  = ~A200 & A199;
  assign \new_[72007]_  = A202 & A201;
  assign \new_[72008]_  = \new_[72007]_  & \new_[72004]_ ;
  assign \new_[72009]_  = \new_[72008]_  & \new_[72001]_ ;
  assign \new_[72013]_  = A265 & A233;
  assign \new_[72014]_  = A232 & \new_[72013]_ ;
  assign \new_[72017]_  = ~A269 & ~A268;
  assign \new_[72020]_  = A299 & A298;
  assign \new_[72021]_  = \new_[72020]_  & \new_[72017]_ ;
  assign \new_[72022]_  = \new_[72021]_  & \new_[72014]_ ;
  assign \new_[72026]_  = ~A168 & A169;
  assign \new_[72027]_  = A170 & \new_[72026]_ ;
  assign \new_[72030]_  = ~A200 & A199;
  assign \new_[72033]_  = A202 & A201;
  assign \new_[72034]_  = \new_[72033]_  & \new_[72030]_ ;
  assign \new_[72035]_  = \new_[72034]_  & \new_[72027]_ ;
  assign \new_[72039]_  = A265 & A233;
  assign \new_[72040]_  = A232 & \new_[72039]_ ;
  assign \new_[72043]_  = ~A269 & ~A268;
  assign \new_[72046]_  = ~A299 & ~A298;
  assign \new_[72047]_  = \new_[72046]_  & \new_[72043]_ ;
  assign \new_[72048]_  = \new_[72047]_  & \new_[72040]_ ;
  assign \new_[72052]_  = ~A168 & A169;
  assign \new_[72053]_  = A170 & \new_[72052]_ ;
  assign \new_[72056]_  = ~A200 & A199;
  assign \new_[72059]_  = A202 & A201;
  assign \new_[72060]_  = \new_[72059]_  & \new_[72056]_ ;
  assign \new_[72061]_  = \new_[72060]_  & \new_[72053]_ ;
  assign \new_[72065]_  = A265 & A233;
  assign \new_[72066]_  = A232 & \new_[72065]_ ;
  assign \new_[72069]_  = ~A299 & ~A267;
  assign \new_[72072]_  = ~A302 & ~A301;
  assign \new_[72073]_  = \new_[72072]_  & \new_[72069]_ ;
  assign \new_[72074]_  = \new_[72073]_  & \new_[72066]_ ;
  assign \new_[72078]_  = ~A168 & A169;
  assign \new_[72079]_  = A170 & \new_[72078]_ ;
  assign \new_[72082]_  = ~A200 & A199;
  assign \new_[72085]_  = A202 & A201;
  assign \new_[72086]_  = \new_[72085]_  & \new_[72082]_ ;
  assign \new_[72087]_  = \new_[72086]_  & \new_[72079]_ ;
  assign \new_[72091]_  = A265 & A233;
  assign \new_[72092]_  = A232 & \new_[72091]_ ;
  assign \new_[72095]_  = ~A299 & A266;
  assign \new_[72098]_  = ~A302 & ~A301;
  assign \new_[72099]_  = \new_[72098]_  & \new_[72095]_ ;
  assign \new_[72100]_  = \new_[72099]_  & \new_[72092]_ ;
  assign \new_[72104]_  = ~A168 & A169;
  assign \new_[72105]_  = A170 & \new_[72104]_ ;
  assign \new_[72108]_  = ~A200 & A199;
  assign \new_[72111]_  = A202 & A201;
  assign \new_[72112]_  = \new_[72111]_  & \new_[72108]_ ;
  assign \new_[72113]_  = \new_[72112]_  & \new_[72105]_ ;
  assign \new_[72117]_  = ~A265 & A233;
  assign \new_[72118]_  = A232 & \new_[72117]_ ;
  assign \new_[72121]_  = ~A299 & ~A266;
  assign \new_[72124]_  = ~A302 & ~A301;
  assign \new_[72125]_  = \new_[72124]_  & \new_[72121]_ ;
  assign \new_[72126]_  = \new_[72125]_  & \new_[72118]_ ;
  assign \new_[72130]_  = ~A168 & A169;
  assign \new_[72131]_  = A170 & \new_[72130]_ ;
  assign \new_[72134]_  = ~A200 & A199;
  assign \new_[72137]_  = A202 & A201;
  assign \new_[72138]_  = \new_[72137]_  & \new_[72134]_ ;
  assign \new_[72139]_  = \new_[72138]_  & \new_[72131]_ ;
  assign \new_[72143]_  = ~A236 & ~A235;
  assign \new_[72144]_  = ~A233 & \new_[72143]_ ;
  assign \new_[72147]_  = A266 & A265;
  assign \new_[72150]_  = ~A300 & A298;
  assign \new_[72151]_  = \new_[72150]_  & \new_[72147]_ ;
  assign \new_[72152]_  = \new_[72151]_  & \new_[72144]_ ;
  assign \new_[72156]_  = ~A168 & A169;
  assign \new_[72157]_  = A170 & \new_[72156]_ ;
  assign \new_[72160]_  = ~A200 & A199;
  assign \new_[72163]_  = A202 & A201;
  assign \new_[72164]_  = \new_[72163]_  & \new_[72160]_ ;
  assign \new_[72165]_  = \new_[72164]_  & \new_[72157]_ ;
  assign \new_[72169]_  = ~A236 & ~A235;
  assign \new_[72170]_  = ~A233 & \new_[72169]_ ;
  assign \new_[72173]_  = A266 & A265;
  assign \new_[72176]_  = A299 & A298;
  assign \new_[72177]_  = \new_[72176]_  & \new_[72173]_ ;
  assign \new_[72178]_  = \new_[72177]_  & \new_[72170]_ ;
  assign \new_[72182]_  = ~A168 & A169;
  assign \new_[72183]_  = A170 & \new_[72182]_ ;
  assign \new_[72186]_  = ~A200 & A199;
  assign \new_[72189]_  = A202 & A201;
  assign \new_[72190]_  = \new_[72189]_  & \new_[72186]_ ;
  assign \new_[72191]_  = \new_[72190]_  & \new_[72183]_ ;
  assign \new_[72195]_  = ~A236 & ~A235;
  assign \new_[72196]_  = ~A233 & \new_[72195]_ ;
  assign \new_[72199]_  = A266 & A265;
  assign \new_[72202]_  = ~A299 & ~A298;
  assign \new_[72203]_  = \new_[72202]_  & \new_[72199]_ ;
  assign \new_[72204]_  = \new_[72203]_  & \new_[72196]_ ;
  assign \new_[72208]_  = ~A168 & A169;
  assign \new_[72209]_  = A170 & \new_[72208]_ ;
  assign \new_[72212]_  = ~A200 & A199;
  assign \new_[72215]_  = A202 & A201;
  assign \new_[72216]_  = \new_[72215]_  & \new_[72212]_ ;
  assign \new_[72217]_  = \new_[72216]_  & \new_[72209]_ ;
  assign \new_[72221]_  = ~A236 & ~A235;
  assign \new_[72222]_  = ~A233 & \new_[72221]_ ;
  assign \new_[72225]_  = ~A267 & ~A266;
  assign \new_[72228]_  = ~A300 & A298;
  assign \new_[72229]_  = \new_[72228]_  & \new_[72225]_ ;
  assign \new_[72230]_  = \new_[72229]_  & \new_[72222]_ ;
  assign \new_[72234]_  = ~A168 & A169;
  assign \new_[72235]_  = A170 & \new_[72234]_ ;
  assign \new_[72238]_  = ~A200 & A199;
  assign \new_[72241]_  = A202 & A201;
  assign \new_[72242]_  = \new_[72241]_  & \new_[72238]_ ;
  assign \new_[72243]_  = \new_[72242]_  & \new_[72235]_ ;
  assign \new_[72247]_  = ~A236 & ~A235;
  assign \new_[72248]_  = ~A233 & \new_[72247]_ ;
  assign \new_[72251]_  = ~A267 & ~A266;
  assign \new_[72254]_  = A299 & A298;
  assign \new_[72255]_  = \new_[72254]_  & \new_[72251]_ ;
  assign \new_[72256]_  = \new_[72255]_  & \new_[72248]_ ;
  assign \new_[72260]_  = ~A168 & A169;
  assign \new_[72261]_  = A170 & \new_[72260]_ ;
  assign \new_[72264]_  = ~A200 & A199;
  assign \new_[72267]_  = A202 & A201;
  assign \new_[72268]_  = \new_[72267]_  & \new_[72264]_ ;
  assign \new_[72269]_  = \new_[72268]_  & \new_[72261]_ ;
  assign \new_[72273]_  = ~A236 & ~A235;
  assign \new_[72274]_  = ~A233 & \new_[72273]_ ;
  assign \new_[72277]_  = ~A267 & ~A266;
  assign \new_[72280]_  = ~A299 & ~A298;
  assign \new_[72281]_  = \new_[72280]_  & \new_[72277]_ ;
  assign \new_[72282]_  = \new_[72281]_  & \new_[72274]_ ;
  assign \new_[72286]_  = ~A168 & A169;
  assign \new_[72287]_  = A170 & \new_[72286]_ ;
  assign \new_[72290]_  = ~A200 & A199;
  assign \new_[72293]_  = A202 & A201;
  assign \new_[72294]_  = \new_[72293]_  & \new_[72290]_ ;
  assign \new_[72295]_  = \new_[72294]_  & \new_[72287]_ ;
  assign \new_[72299]_  = ~A236 & ~A235;
  assign \new_[72300]_  = ~A233 & \new_[72299]_ ;
  assign \new_[72303]_  = ~A266 & ~A265;
  assign \new_[72306]_  = ~A300 & A298;
  assign \new_[72307]_  = \new_[72306]_  & \new_[72303]_ ;
  assign \new_[72308]_  = \new_[72307]_  & \new_[72300]_ ;
  assign \new_[72312]_  = ~A168 & A169;
  assign \new_[72313]_  = A170 & \new_[72312]_ ;
  assign \new_[72316]_  = ~A200 & A199;
  assign \new_[72319]_  = A202 & A201;
  assign \new_[72320]_  = \new_[72319]_  & \new_[72316]_ ;
  assign \new_[72321]_  = \new_[72320]_  & \new_[72313]_ ;
  assign \new_[72325]_  = ~A236 & ~A235;
  assign \new_[72326]_  = ~A233 & \new_[72325]_ ;
  assign \new_[72329]_  = ~A266 & ~A265;
  assign \new_[72332]_  = A299 & A298;
  assign \new_[72333]_  = \new_[72332]_  & \new_[72329]_ ;
  assign \new_[72334]_  = \new_[72333]_  & \new_[72326]_ ;
  assign \new_[72338]_  = ~A168 & A169;
  assign \new_[72339]_  = A170 & \new_[72338]_ ;
  assign \new_[72342]_  = ~A200 & A199;
  assign \new_[72345]_  = A202 & A201;
  assign \new_[72346]_  = \new_[72345]_  & \new_[72342]_ ;
  assign \new_[72347]_  = \new_[72346]_  & \new_[72339]_ ;
  assign \new_[72351]_  = ~A236 & ~A235;
  assign \new_[72352]_  = ~A233 & \new_[72351]_ ;
  assign \new_[72355]_  = ~A266 & ~A265;
  assign \new_[72358]_  = ~A299 & ~A298;
  assign \new_[72359]_  = \new_[72358]_  & \new_[72355]_ ;
  assign \new_[72360]_  = \new_[72359]_  & \new_[72352]_ ;
  assign \new_[72364]_  = ~A168 & A169;
  assign \new_[72365]_  = A170 & \new_[72364]_ ;
  assign \new_[72368]_  = ~A200 & A199;
  assign \new_[72371]_  = A202 & A201;
  assign \new_[72372]_  = \new_[72371]_  & \new_[72368]_ ;
  assign \new_[72373]_  = \new_[72372]_  & \new_[72365]_ ;
  assign \new_[72377]_  = A265 & ~A234;
  assign \new_[72378]_  = ~A233 & \new_[72377]_ ;
  assign \new_[72381]_  = A298 & A266;
  assign \new_[72384]_  = ~A302 & ~A301;
  assign \new_[72385]_  = \new_[72384]_  & \new_[72381]_ ;
  assign \new_[72386]_  = \new_[72385]_  & \new_[72378]_ ;
  assign \new_[72390]_  = ~A168 & A169;
  assign \new_[72391]_  = A170 & \new_[72390]_ ;
  assign \new_[72394]_  = ~A200 & A199;
  assign \new_[72397]_  = A202 & A201;
  assign \new_[72398]_  = \new_[72397]_  & \new_[72394]_ ;
  assign \new_[72399]_  = \new_[72398]_  & \new_[72391]_ ;
  assign \new_[72403]_  = ~A266 & ~A234;
  assign \new_[72404]_  = ~A233 & \new_[72403]_ ;
  assign \new_[72407]_  = ~A269 & ~A268;
  assign \new_[72410]_  = ~A300 & A298;
  assign \new_[72411]_  = \new_[72410]_  & \new_[72407]_ ;
  assign \new_[72412]_  = \new_[72411]_  & \new_[72404]_ ;
  assign \new_[72416]_  = ~A168 & A169;
  assign \new_[72417]_  = A170 & \new_[72416]_ ;
  assign \new_[72420]_  = ~A200 & A199;
  assign \new_[72423]_  = A202 & A201;
  assign \new_[72424]_  = \new_[72423]_  & \new_[72420]_ ;
  assign \new_[72425]_  = \new_[72424]_  & \new_[72417]_ ;
  assign \new_[72429]_  = ~A266 & ~A234;
  assign \new_[72430]_  = ~A233 & \new_[72429]_ ;
  assign \new_[72433]_  = ~A269 & ~A268;
  assign \new_[72436]_  = A299 & A298;
  assign \new_[72437]_  = \new_[72436]_  & \new_[72433]_ ;
  assign \new_[72438]_  = \new_[72437]_  & \new_[72430]_ ;
  assign \new_[72442]_  = ~A168 & A169;
  assign \new_[72443]_  = A170 & \new_[72442]_ ;
  assign \new_[72446]_  = ~A200 & A199;
  assign \new_[72449]_  = A202 & A201;
  assign \new_[72450]_  = \new_[72449]_  & \new_[72446]_ ;
  assign \new_[72451]_  = \new_[72450]_  & \new_[72443]_ ;
  assign \new_[72455]_  = ~A266 & ~A234;
  assign \new_[72456]_  = ~A233 & \new_[72455]_ ;
  assign \new_[72459]_  = ~A269 & ~A268;
  assign \new_[72462]_  = ~A299 & ~A298;
  assign \new_[72463]_  = \new_[72462]_  & \new_[72459]_ ;
  assign \new_[72464]_  = \new_[72463]_  & \new_[72456]_ ;
  assign \new_[72468]_  = ~A168 & A169;
  assign \new_[72469]_  = A170 & \new_[72468]_ ;
  assign \new_[72472]_  = ~A200 & A199;
  assign \new_[72475]_  = A202 & A201;
  assign \new_[72476]_  = \new_[72475]_  & \new_[72472]_ ;
  assign \new_[72477]_  = \new_[72476]_  & \new_[72469]_ ;
  assign \new_[72481]_  = ~A266 & ~A234;
  assign \new_[72482]_  = ~A233 & \new_[72481]_ ;
  assign \new_[72485]_  = A298 & ~A267;
  assign \new_[72488]_  = ~A302 & ~A301;
  assign \new_[72489]_  = \new_[72488]_  & \new_[72485]_ ;
  assign \new_[72490]_  = \new_[72489]_  & \new_[72482]_ ;
  assign \new_[72494]_  = ~A168 & A169;
  assign \new_[72495]_  = A170 & \new_[72494]_ ;
  assign \new_[72498]_  = ~A200 & A199;
  assign \new_[72501]_  = A202 & A201;
  assign \new_[72502]_  = \new_[72501]_  & \new_[72498]_ ;
  assign \new_[72503]_  = \new_[72502]_  & \new_[72495]_ ;
  assign \new_[72507]_  = ~A265 & ~A234;
  assign \new_[72508]_  = ~A233 & \new_[72507]_ ;
  assign \new_[72511]_  = A298 & ~A266;
  assign \new_[72514]_  = ~A302 & ~A301;
  assign \new_[72515]_  = \new_[72514]_  & \new_[72511]_ ;
  assign \new_[72516]_  = \new_[72515]_  & \new_[72508]_ ;
  assign \new_[72520]_  = ~A168 & A169;
  assign \new_[72521]_  = A170 & \new_[72520]_ ;
  assign \new_[72524]_  = ~A200 & A199;
  assign \new_[72527]_  = A202 & A201;
  assign \new_[72528]_  = \new_[72527]_  & \new_[72524]_ ;
  assign \new_[72529]_  = \new_[72528]_  & \new_[72521]_ ;
  assign \new_[72533]_  = A265 & ~A233;
  assign \new_[72534]_  = ~A232 & \new_[72533]_ ;
  assign \new_[72537]_  = A298 & A266;
  assign \new_[72540]_  = ~A302 & ~A301;
  assign \new_[72541]_  = \new_[72540]_  & \new_[72537]_ ;
  assign \new_[72542]_  = \new_[72541]_  & \new_[72534]_ ;
  assign \new_[72546]_  = ~A168 & A169;
  assign \new_[72547]_  = A170 & \new_[72546]_ ;
  assign \new_[72550]_  = ~A200 & A199;
  assign \new_[72553]_  = A202 & A201;
  assign \new_[72554]_  = \new_[72553]_  & \new_[72550]_ ;
  assign \new_[72555]_  = \new_[72554]_  & \new_[72547]_ ;
  assign \new_[72559]_  = ~A266 & ~A233;
  assign \new_[72560]_  = ~A232 & \new_[72559]_ ;
  assign \new_[72563]_  = ~A269 & ~A268;
  assign \new_[72566]_  = ~A300 & A298;
  assign \new_[72567]_  = \new_[72566]_  & \new_[72563]_ ;
  assign \new_[72568]_  = \new_[72567]_  & \new_[72560]_ ;
  assign \new_[72572]_  = ~A168 & A169;
  assign \new_[72573]_  = A170 & \new_[72572]_ ;
  assign \new_[72576]_  = ~A200 & A199;
  assign \new_[72579]_  = A202 & A201;
  assign \new_[72580]_  = \new_[72579]_  & \new_[72576]_ ;
  assign \new_[72581]_  = \new_[72580]_  & \new_[72573]_ ;
  assign \new_[72585]_  = ~A266 & ~A233;
  assign \new_[72586]_  = ~A232 & \new_[72585]_ ;
  assign \new_[72589]_  = ~A269 & ~A268;
  assign \new_[72592]_  = A299 & A298;
  assign \new_[72593]_  = \new_[72592]_  & \new_[72589]_ ;
  assign \new_[72594]_  = \new_[72593]_  & \new_[72586]_ ;
  assign \new_[72598]_  = ~A168 & A169;
  assign \new_[72599]_  = A170 & \new_[72598]_ ;
  assign \new_[72602]_  = ~A200 & A199;
  assign \new_[72605]_  = A202 & A201;
  assign \new_[72606]_  = \new_[72605]_  & \new_[72602]_ ;
  assign \new_[72607]_  = \new_[72606]_  & \new_[72599]_ ;
  assign \new_[72611]_  = ~A266 & ~A233;
  assign \new_[72612]_  = ~A232 & \new_[72611]_ ;
  assign \new_[72615]_  = ~A269 & ~A268;
  assign \new_[72618]_  = ~A299 & ~A298;
  assign \new_[72619]_  = \new_[72618]_  & \new_[72615]_ ;
  assign \new_[72620]_  = \new_[72619]_  & \new_[72612]_ ;
  assign \new_[72624]_  = ~A168 & A169;
  assign \new_[72625]_  = A170 & \new_[72624]_ ;
  assign \new_[72628]_  = ~A200 & A199;
  assign \new_[72631]_  = A202 & A201;
  assign \new_[72632]_  = \new_[72631]_  & \new_[72628]_ ;
  assign \new_[72633]_  = \new_[72632]_  & \new_[72625]_ ;
  assign \new_[72637]_  = ~A266 & ~A233;
  assign \new_[72638]_  = ~A232 & \new_[72637]_ ;
  assign \new_[72641]_  = A298 & ~A267;
  assign \new_[72644]_  = ~A302 & ~A301;
  assign \new_[72645]_  = \new_[72644]_  & \new_[72641]_ ;
  assign \new_[72646]_  = \new_[72645]_  & \new_[72638]_ ;
  assign \new_[72650]_  = ~A168 & A169;
  assign \new_[72651]_  = A170 & \new_[72650]_ ;
  assign \new_[72654]_  = ~A200 & A199;
  assign \new_[72657]_  = A202 & A201;
  assign \new_[72658]_  = \new_[72657]_  & \new_[72654]_ ;
  assign \new_[72659]_  = \new_[72658]_  & \new_[72651]_ ;
  assign \new_[72663]_  = ~A265 & ~A233;
  assign \new_[72664]_  = ~A232 & \new_[72663]_ ;
  assign \new_[72667]_  = A298 & ~A266;
  assign \new_[72670]_  = ~A302 & ~A301;
  assign \new_[72671]_  = \new_[72670]_  & \new_[72667]_ ;
  assign \new_[72672]_  = \new_[72671]_  & \new_[72664]_ ;
  assign \new_[72676]_  = ~A168 & A169;
  assign \new_[72677]_  = A170 & \new_[72676]_ ;
  assign \new_[72680]_  = ~A200 & A199;
  assign \new_[72683]_  = A203 & A201;
  assign \new_[72684]_  = \new_[72683]_  & \new_[72680]_ ;
  assign \new_[72685]_  = \new_[72684]_  & \new_[72677]_ ;
  assign \new_[72689]_  = A265 & A233;
  assign \new_[72690]_  = A232 & \new_[72689]_ ;
  assign \new_[72693]_  = ~A269 & ~A268;
  assign \new_[72696]_  = ~A300 & ~A299;
  assign \new_[72697]_  = \new_[72696]_  & \new_[72693]_ ;
  assign \new_[72698]_  = \new_[72697]_  & \new_[72690]_ ;
  assign \new_[72702]_  = ~A168 & A169;
  assign \new_[72703]_  = A170 & \new_[72702]_ ;
  assign \new_[72706]_  = ~A200 & A199;
  assign \new_[72709]_  = A203 & A201;
  assign \new_[72710]_  = \new_[72709]_  & \new_[72706]_ ;
  assign \new_[72711]_  = \new_[72710]_  & \new_[72703]_ ;
  assign \new_[72715]_  = A265 & A233;
  assign \new_[72716]_  = A232 & \new_[72715]_ ;
  assign \new_[72719]_  = ~A269 & ~A268;
  assign \new_[72722]_  = A299 & A298;
  assign \new_[72723]_  = \new_[72722]_  & \new_[72719]_ ;
  assign \new_[72724]_  = \new_[72723]_  & \new_[72716]_ ;
  assign \new_[72728]_  = ~A168 & A169;
  assign \new_[72729]_  = A170 & \new_[72728]_ ;
  assign \new_[72732]_  = ~A200 & A199;
  assign \new_[72735]_  = A203 & A201;
  assign \new_[72736]_  = \new_[72735]_  & \new_[72732]_ ;
  assign \new_[72737]_  = \new_[72736]_  & \new_[72729]_ ;
  assign \new_[72741]_  = A265 & A233;
  assign \new_[72742]_  = A232 & \new_[72741]_ ;
  assign \new_[72745]_  = ~A269 & ~A268;
  assign \new_[72748]_  = ~A299 & ~A298;
  assign \new_[72749]_  = \new_[72748]_  & \new_[72745]_ ;
  assign \new_[72750]_  = \new_[72749]_  & \new_[72742]_ ;
  assign \new_[72754]_  = ~A168 & A169;
  assign \new_[72755]_  = A170 & \new_[72754]_ ;
  assign \new_[72758]_  = ~A200 & A199;
  assign \new_[72761]_  = A203 & A201;
  assign \new_[72762]_  = \new_[72761]_  & \new_[72758]_ ;
  assign \new_[72763]_  = \new_[72762]_  & \new_[72755]_ ;
  assign \new_[72767]_  = A265 & A233;
  assign \new_[72768]_  = A232 & \new_[72767]_ ;
  assign \new_[72771]_  = ~A299 & ~A267;
  assign \new_[72774]_  = ~A302 & ~A301;
  assign \new_[72775]_  = \new_[72774]_  & \new_[72771]_ ;
  assign \new_[72776]_  = \new_[72775]_  & \new_[72768]_ ;
  assign \new_[72780]_  = ~A168 & A169;
  assign \new_[72781]_  = A170 & \new_[72780]_ ;
  assign \new_[72784]_  = ~A200 & A199;
  assign \new_[72787]_  = A203 & A201;
  assign \new_[72788]_  = \new_[72787]_  & \new_[72784]_ ;
  assign \new_[72789]_  = \new_[72788]_  & \new_[72781]_ ;
  assign \new_[72793]_  = A265 & A233;
  assign \new_[72794]_  = A232 & \new_[72793]_ ;
  assign \new_[72797]_  = ~A299 & A266;
  assign \new_[72800]_  = ~A302 & ~A301;
  assign \new_[72801]_  = \new_[72800]_  & \new_[72797]_ ;
  assign \new_[72802]_  = \new_[72801]_  & \new_[72794]_ ;
  assign \new_[72806]_  = ~A168 & A169;
  assign \new_[72807]_  = A170 & \new_[72806]_ ;
  assign \new_[72810]_  = ~A200 & A199;
  assign \new_[72813]_  = A203 & A201;
  assign \new_[72814]_  = \new_[72813]_  & \new_[72810]_ ;
  assign \new_[72815]_  = \new_[72814]_  & \new_[72807]_ ;
  assign \new_[72819]_  = ~A265 & A233;
  assign \new_[72820]_  = A232 & \new_[72819]_ ;
  assign \new_[72823]_  = ~A299 & ~A266;
  assign \new_[72826]_  = ~A302 & ~A301;
  assign \new_[72827]_  = \new_[72826]_  & \new_[72823]_ ;
  assign \new_[72828]_  = \new_[72827]_  & \new_[72820]_ ;
  assign \new_[72832]_  = ~A168 & A169;
  assign \new_[72833]_  = A170 & \new_[72832]_ ;
  assign \new_[72836]_  = ~A200 & A199;
  assign \new_[72839]_  = A203 & A201;
  assign \new_[72840]_  = \new_[72839]_  & \new_[72836]_ ;
  assign \new_[72841]_  = \new_[72840]_  & \new_[72833]_ ;
  assign \new_[72845]_  = ~A236 & ~A235;
  assign \new_[72846]_  = ~A233 & \new_[72845]_ ;
  assign \new_[72849]_  = A266 & A265;
  assign \new_[72852]_  = ~A300 & A298;
  assign \new_[72853]_  = \new_[72852]_  & \new_[72849]_ ;
  assign \new_[72854]_  = \new_[72853]_  & \new_[72846]_ ;
  assign \new_[72858]_  = ~A168 & A169;
  assign \new_[72859]_  = A170 & \new_[72858]_ ;
  assign \new_[72862]_  = ~A200 & A199;
  assign \new_[72865]_  = A203 & A201;
  assign \new_[72866]_  = \new_[72865]_  & \new_[72862]_ ;
  assign \new_[72867]_  = \new_[72866]_  & \new_[72859]_ ;
  assign \new_[72871]_  = ~A236 & ~A235;
  assign \new_[72872]_  = ~A233 & \new_[72871]_ ;
  assign \new_[72875]_  = A266 & A265;
  assign \new_[72878]_  = A299 & A298;
  assign \new_[72879]_  = \new_[72878]_  & \new_[72875]_ ;
  assign \new_[72880]_  = \new_[72879]_  & \new_[72872]_ ;
  assign \new_[72884]_  = ~A168 & A169;
  assign \new_[72885]_  = A170 & \new_[72884]_ ;
  assign \new_[72888]_  = ~A200 & A199;
  assign \new_[72891]_  = A203 & A201;
  assign \new_[72892]_  = \new_[72891]_  & \new_[72888]_ ;
  assign \new_[72893]_  = \new_[72892]_  & \new_[72885]_ ;
  assign \new_[72897]_  = ~A236 & ~A235;
  assign \new_[72898]_  = ~A233 & \new_[72897]_ ;
  assign \new_[72901]_  = A266 & A265;
  assign \new_[72904]_  = ~A299 & ~A298;
  assign \new_[72905]_  = \new_[72904]_  & \new_[72901]_ ;
  assign \new_[72906]_  = \new_[72905]_  & \new_[72898]_ ;
  assign \new_[72910]_  = ~A168 & A169;
  assign \new_[72911]_  = A170 & \new_[72910]_ ;
  assign \new_[72914]_  = ~A200 & A199;
  assign \new_[72917]_  = A203 & A201;
  assign \new_[72918]_  = \new_[72917]_  & \new_[72914]_ ;
  assign \new_[72919]_  = \new_[72918]_  & \new_[72911]_ ;
  assign \new_[72923]_  = ~A236 & ~A235;
  assign \new_[72924]_  = ~A233 & \new_[72923]_ ;
  assign \new_[72927]_  = ~A267 & ~A266;
  assign \new_[72930]_  = ~A300 & A298;
  assign \new_[72931]_  = \new_[72930]_  & \new_[72927]_ ;
  assign \new_[72932]_  = \new_[72931]_  & \new_[72924]_ ;
  assign \new_[72936]_  = ~A168 & A169;
  assign \new_[72937]_  = A170 & \new_[72936]_ ;
  assign \new_[72940]_  = ~A200 & A199;
  assign \new_[72943]_  = A203 & A201;
  assign \new_[72944]_  = \new_[72943]_  & \new_[72940]_ ;
  assign \new_[72945]_  = \new_[72944]_  & \new_[72937]_ ;
  assign \new_[72949]_  = ~A236 & ~A235;
  assign \new_[72950]_  = ~A233 & \new_[72949]_ ;
  assign \new_[72953]_  = ~A267 & ~A266;
  assign \new_[72956]_  = A299 & A298;
  assign \new_[72957]_  = \new_[72956]_  & \new_[72953]_ ;
  assign \new_[72958]_  = \new_[72957]_  & \new_[72950]_ ;
  assign \new_[72962]_  = ~A168 & A169;
  assign \new_[72963]_  = A170 & \new_[72962]_ ;
  assign \new_[72966]_  = ~A200 & A199;
  assign \new_[72969]_  = A203 & A201;
  assign \new_[72970]_  = \new_[72969]_  & \new_[72966]_ ;
  assign \new_[72971]_  = \new_[72970]_  & \new_[72963]_ ;
  assign \new_[72975]_  = ~A236 & ~A235;
  assign \new_[72976]_  = ~A233 & \new_[72975]_ ;
  assign \new_[72979]_  = ~A267 & ~A266;
  assign \new_[72982]_  = ~A299 & ~A298;
  assign \new_[72983]_  = \new_[72982]_  & \new_[72979]_ ;
  assign \new_[72984]_  = \new_[72983]_  & \new_[72976]_ ;
  assign \new_[72988]_  = ~A168 & A169;
  assign \new_[72989]_  = A170 & \new_[72988]_ ;
  assign \new_[72992]_  = ~A200 & A199;
  assign \new_[72995]_  = A203 & A201;
  assign \new_[72996]_  = \new_[72995]_  & \new_[72992]_ ;
  assign \new_[72997]_  = \new_[72996]_  & \new_[72989]_ ;
  assign \new_[73001]_  = ~A236 & ~A235;
  assign \new_[73002]_  = ~A233 & \new_[73001]_ ;
  assign \new_[73005]_  = ~A266 & ~A265;
  assign \new_[73008]_  = ~A300 & A298;
  assign \new_[73009]_  = \new_[73008]_  & \new_[73005]_ ;
  assign \new_[73010]_  = \new_[73009]_  & \new_[73002]_ ;
  assign \new_[73014]_  = ~A168 & A169;
  assign \new_[73015]_  = A170 & \new_[73014]_ ;
  assign \new_[73018]_  = ~A200 & A199;
  assign \new_[73021]_  = A203 & A201;
  assign \new_[73022]_  = \new_[73021]_  & \new_[73018]_ ;
  assign \new_[73023]_  = \new_[73022]_  & \new_[73015]_ ;
  assign \new_[73027]_  = ~A236 & ~A235;
  assign \new_[73028]_  = ~A233 & \new_[73027]_ ;
  assign \new_[73031]_  = ~A266 & ~A265;
  assign \new_[73034]_  = A299 & A298;
  assign \new_[73035]_  = \new_[73034]_  & \new_[73031]_ ;
  assign \new_[73036]_  = \new_[73035]_  & \new_[73028]_ ;
  assign \new_[73040]_  = ~A168 & A169;
  assign \new_[73041]_  = A170 & \new_[73040]_ ;
  assign \new_[73044]_  = ~A200 & A199;
  assign \new_[73047]_  = A203 & A201;
  assign \new_[73048]_  = \new_[73047]_  & \new_[73044]_ ;
  assign \new_[73049]_  = \new_[73048]_  & \new_[73041]_ ;
  assign \new_[73053]_  = ~A236 & ~A235;
  assign \new_[73054]_  = ~A233 & \new_[73053]_ ;
  assign \new_[73057]_  = ~A266 & ~A265;
  assign \new_[73060]_  = ~A299 & ~A298;
  assign \new_[73061]_  = \new_[73060]_  & \new_[73057]_ ;
  assign \new_[73062]_  = \new_[73061]_  & \new_[73054]_ ;
  assign \new_[73066]_  = ~A168 & A169;
  assign \new_[73067]_  = A170 & \new_[73066]_ ;
  assign \new_[73070]_  = ~A200 & A199;
  assign \new_[73073]_  = A203 & A201;
  assign \new_[73074]_  = \new_[73073]_  & \new_[73070]_ ;
  assign \new_[73075]_  = \new_[73074]_  & \new_[73067]_ ;
  assign \new_[73079]_  = A265 & ~A234;
  assign \new_[73080]_  = ~A233 & \new_[73079]_ ;
  assign \new_[73083]_  = A298 & A266;
  assign \new_[73086]_  = ~A302 & ~A301;
  assign \new_[73087]_  = \new_[73086]_  & \new_[73083]_ ;
  assign \new_[73088]_  = \new_[73087]_  & \new_[73080]_ ;
  assign \new_[73092]_  = ~A168 & A169;
  assign \new_[73093]_  = A170 & \new_[73092]_ ;
  assign \new_[73096]_  = ~A200 & A199;
  assign \new_[73099]_  = A203 & A201;
  assign \new_[73100]_  = \new_[73099]_  & \new_[73096]_ ;
  assign \new_[73101]_  = \new_[73100]_  & \new_[73093]_ ;
  assign \new_[73105]_  = ~A266 & ~A234;
  assign \new_[73106]_  = ~A233 & \new_[73105]_ ;
  assign \new_[73109]_  = ~A269 & ~A268;
  assign \new_[73112]_  = ~A300 & A298;
  assign \new_[73113]_  = \new_[73112]_  & \new_[73109]_ ;
  assign \new_[73114]_  = \new_[73113]_  & \new_[73106]_ ;
  assign \new_[73118]_  = ~A168 & A169;
  assign \new_[73119]_  = A170 & \new_[73118]_ ;
  assign \new_[73122]_  = ~A200 & A199;
  assign \new_[73125]_  = A203 & A201;
  assign \new_[73126]_  = \new_[73125]_  & \new_[73122]_ ;
  assign \new_[73127]_  = \new_[73126]_  & \new_[73119]_ ;
  assign \new_[73131]_  = ~A266 & ~A234;
  assign \new_[73132]_  = ~A233 & \new_[73131]_ ;
  assign \new_[73135]_  = ~A269 & ~A268;
  assign \new_[73138]_  = A299 & A298;
  assign \new_[73139]_  = \new_[73138]_  & \new_[73135]_ ;
  assign \new_[73140]_  = \new_[73139]_  & \new_[73132]_ ;
  assign \new_[73144]_  = ~A168 & A169;
  assign \new_[73145]_  = A170 & \new_[73144]_ ;
  assign \new_[73148]_  = ~A200 & A199;
  assign \new_[73151]_  = A203 & A201;
  assign \new_[73152]_  = \new_[73151]_  & \new_[73148]_ ;
  assign \new_[73153]_  = \new_[73152]_  & \new_[73145]_ ;
  assign \new_[73157]_  = ~A266 & ~A234;
  assign \new_[73158]_  = ~A233 & \new_[73157]_ ;
  assign \new_[73161]_  = ~A269 & ~A268;
  assign \new_[73164]_  = ~A299 & ~A298;
  assign \new_[73165]_  = \new_[73164]_  & \new_[73161]_ ;
  assign \new_[73166]_  = \new_[73165]_  & \new_[73158]_ ;
  assign \new_[73170]_  = ~A168 & A169;
  assign \new_[73171]_  = A170 & \new_[73170]_ ;
  assign \new_[73174]_  = ~A200 & A199;
  assign \new_[73177]_  = A203 & A201;
  assign \new_[73178]_  = \new_[73177]_  & \new_[73174]_ ;
  assign \new_[73179]_  = \new_[73178]_  & \new_[73171]_ ;
  assign \new_[73183]_  = ~A266 & ~A234;
  assign \new_[73184]_  = ~A233 & \new_[73183]_ ;
  assign \new_[73187]_  = A298 & ~A267;
  assign \new_[73190]_  = ~A302 & ~A301;
  assign \new_[73191]_  = \new_[73190]_  & \new_[73187]_ ;
  assign \new_[73192]_  = \new_[73191]_  & \new_[73184]_ ;
  assign \new_[73196]_  = ~A168 & A169;
  assign \new_[73197]_  = A170 & \new_[73196]_ ;
  assign \new_[73200]_  = ~A200 & A199;
  assign \new_[73203]_  = A203 & A201;
  assign \new_[73204]_  = \new_[73203]_  & \new_[73200]_ ;
  assign \new_[73205]_  = \new_[73204]_  & \new_[73197]_ ;
  assign \new_[73209]_  = ~A265 & ~A234;
  assign \new_[73210]_  = ~A233 & \new_[73209]_ ;
  assign \new_[73213]_  = A298 & ~A266;
  assign \new_[73216]_  = ~A302 & ~A301;
  assign \new_[73217]_  = \new_[73216]_  & \new_[73213]_ ;
  assign \new_[73218]_  = \new_[73217]_  & \new_[73210]_ ;
  assign \new_[73222]_  = ~A168 & A169;
  assign \new_[73223]_  = A170 & \new_[73222]_ ;
  assign \new_[73226]_  = ~A200 & A199;
  assign \new_[73229]_  = A203 & A201;
  assign \new_[73230]_  = \new_[73229]_  & \new_[73226]_ ;
  assign \new_[73231]_  = \new_[73230]_  & \new_[73223]_ ;
  assign \new_[73235]_  = A265 & ~A233;
  assign \new_[73236]_  = ~A232 & \new_[73235]_ ;
  assign \new_[73239]_  = A298 & A266;
  assign \new_[73242]_  = ~A302 & ~A301;
  assign \new_[73243]_  = \new_[73242]_  & \new_[73239]_ ;
  assign \new_[73244]_  = \new_[73243]_  & \new_[73236]_ ;
  assign \new_[73248]_  = ~A168 & A169;
  assign \new_[73249]_  = A170 & \new_[73248]_ ;
  assign \new_[73252]_  = ~A200 & A199;
  assign \new_[73255]_  = A203 & A201;
  assign \new_[73256]_  = \new_[73255]_  & \new_[73252]_ ;
  assign \new_[73257]_  = \new_[73256]_  & \new_[73249]_ ;
  assign \new_[73261]_  = ~A266 & ~A233;
  assign \new_[73262]_  = ~A232 & \new_[73261]_ ;
  assign \new_[73265]_  = ~A269 & ~A268;
  assign \new_[73268]_  = ~A300 & A298;
  assign \new_[73269]_  = \new_[73268]_  & \new_[73265]_ ;
  assign \new_[73270]_  = \new_[73269]_  & \new_[73262]_ ;
  assign \new_[73274]_  = ~A168 & A169;
  assign \new_[73275]_  = A170 & \new_[73274]_ ;
  assign \new_[73278]_  = ~A200 & A199;
  assign \new_[73281]_  = A203 & A201;
  assign \new_[73282]_  = \new_[73281]_  & \new_[73278]_ ;
  assign \new_[73283]_  = \new_[73282]_  & \new_[73275]_ ;
  assign \new_[73287]_  = ~A266 & ~A233;
  assign \new_[73288]_  = ~A232 & \new_[73287]_ ;
  assign \new_[73291]_  = ~A269 & ~A268;
  assign \new_[73294]_  = A299 & A298;
  assign \new_[73295]_  = \new_[73294]_  & \new_[73291]_ ;
  assign \new_[73296]_  = \new_[73295]_  & \new_[73288]_ ;
  assign \new_[73300]_  = ~A168 & A169;
  assign \new_[73301]_  = A170 & \new_[73300]_ ;
  assign \new_[73304]_  = ~A200 & A199;
  assign \new_[73307]_  = A203 & A201;
  assign \new_[73308]_  = \new_[73307]_  & \new_[73304]_ ;
  assign \new_[73309]_  = \new_[73308]_  & \new_[73301]_ ;
  assign \new_[73313]_  = ~A266 & ~A233;
  assign \new_[73314]_  = ~A232 & \new_[73313]_ ;
  assign \new_[73317]_  = ~A269 & ~A268;
  assign \new_[73320]_  = ~A299 & ~A298;
  assign \new_[73321]_  = \new_[73320]_  & \new_[73317]_ ;
  assign \new_[73322]_  = \new_[73321]_  & \new_[73314]_ ;
  assign \new_[73326]_  = ~A168 & A169;
  assign \new_[73327]_  = A170 & \new_[73326]_ ;
  assign \new_[73330]_  = ~A200 & A199;
  assign \new_[73333]_  = A203 & A201;
  assign \new_[73334]_  = \new_[73333]_  & \new_[73330]_ ;
  assign \new_[73335]_  = \new_[73334]_  & \new_[73327]_ ;
  assign \new_[73339]_  = ~A266 & ~A233;
  assign \new_[73340]_  = ~A232 & \new_[73339]_ ;
  assign \new_[73343]_  = A298 & ~A267;
  assign \new_[73346]_  = ~A302 & ~A301;
  assign \new_[73347]_  = \new_[73346]_  & \new_[73343]_ ;
  assign \new_[73348]_  = \new_[73347]_  & \new_[73340]_ ;
  assign \new_[73352]_  = ~A168 & A169;
  assign \new_[73353]_  = A170 & \new_[73352]_ ;
  assign \new_[73356]_  = ~A200 & A199;
  assign \new_[73359]_  = A203 & A201;
  assign \new_[73360]_  = \new_[73359]_  & \new_[73356]_ ;
  assign \new_[73361]_  = \new_[73360]_  & \new_[73353]_ ;
  assign \new_[73365]_  = ~A265 & ~A233;
  assign \new_[73366]_  = ~A232 & \new_[73365]_ ;
  assign \new_[73369]_  = A298 & ~A266;
  assign \new_[73372]_  = ~A302 & ~A301;
  assign \new_[73373]_  = \new_[73372]_  & \new_[73369]_ ;
  assign \new_[73374]_  = \new_[73373]_  & \new_[73366]_ ;
  assign \new_[73378]_  = ~A168 & A169;
  assign \new_[73379]_  = A170 & \new_[73378]_ ;
  assign \new_[73382]_  = A199 & A166;
  assign \new_[73385]_  = A201 & ~A200;
  assign \new_[73386]_  = \new_[73385]_  & \new_[73382]_ ;
  assign \new_[73387]_  = \new_[73386]_  & \new_[73379]_ ;
  assign \new_[73391]_  = A233 & ~A232;
  assign \new_[73392]_  = A202 & \new_[73391]_ ;
  assign \new_[73395]_  = ~A299 & A298;
  assign \new_[73398]_  = A301 & A300;
  assign \new_[73399]_  = \new_[73398]_  & \new_[73395]_ ;
  assign \new_[73400]_  = \new_[73399]_  & \new_[73392]_ ;
  assign \new_[73404]_  = ~A168 & A169;
  assign \new_[73405]_  = A170 & \new_[73404]_ ;
  assign \new_[73408]_  = A199 & A166;
  assign \new_[73411]_  = A201 & ~A200;
  assign \new_[73412]_  = \new_[73411]_  & \new_[73408]_ ;
  assign \new_[73413]_  = \new_[73412]_  & \new_[73405]_ ;
  assign \new_[73417]_  = A233 & ~A232;
  assign \new_[73418]_  = A202 & \new_[73417]_ ;
  assign \new_[73421]_  = ~A299 & A298;
  assign \new_[73424]_  = A302 & A300;
  assign \new_[73425]_  = \new_[73424]_  & \new_[73421]_ ;
  assign \new_[73426]_  = \new_[73425]_  & \new_[73418]_ ;
  assign \new_[73430]_  = ~A168 & A169;
  assign \new_[73431]_  = A170 & \new_[73430]_ ;
  assign \new_[73434]_  = A199 & A166;
  assign \new_[73437]_  = A201 & ~A200;
  assign \new_[73438]_  = \new_[73437]_  & \new_[73434]_ ;
  assign \new_[73439]_  = \new_[73438]_  & \new_[73431]_ ;
  assign \new_[73443]_  = A233 & ~A232;
  assign \new_[73444]_  = A202 & \new_[73443]_ ;
  assign \new_[73447]_  = ~A266 & A265;
  assign \new_[73450]_  = A268 & A267;
  assign \new_[73451]_  = \new_[73450]_  & \new_[73447]_ ;
  assign \new_[73452]_  = \new_[73451]_  & \new_[73444]_ ;
  assign \new_[73456]_  = ~A168 & A169;
  assign \new_[73457]_  = A170 & \new_[73456]_ ;
  assign \new_[73460]_  = A199 & A166;
  assign \new_[73463]_  = A201 & ~A200;
  assign \new_[73464]_  = \new_[73463]_  & \new_[73460]_ ;
  assign \new_[73465]_  = \new_[73464]_  & \new_[73457]_ ;
  assign \new_[73469]_  = A233 & ~A232;
  assign \new_[73470]_  = A202 & \new_[73469]_ ;
  assign \new_[73473]_  = ~A266 & A265;
  assign \new_[73476]_  = A269 & A267;
  assign \new_[73477]_  = \new_[73476]_  & \new_[73473]_ ;
  assign \new_[73478]_  = \new_[73477]_  & \new_[73470]_ ;
  assign \new_[73482]_  = ~A168 & A169;
  assign \new_[73483]_  = A170 & \new_[73482]_ ;
  assign \new_[73486]_  = A199 & A166;
  assign \new_[73489]_  = A201 & ~A200;
  assign \new_[73490]_  = \new_[73489]_  & \new_[73486]_ ;
  assign \new_[73491]_  = \new_[73490]_  & \new_[73483]_ ;
  assign \new_[73495]_  = A233 & ~A232;
  assign \new_[73496]_  = A203 & \new_[73495]_ ;
  assign \new_[73499]_  = ~A299 & A298;
  assign \new_[73502]_  = A301 & A300;
  assign \new_[73503]_  = \new_[73502]_  & \new_[73499]_ ;
  assign \new_[73504]_  = \new_[73503]_  & \new_[73496]_ ;
  assign \new_[73508]_  = ~A168 & A169;
  assign \new_[73509]_  = A170 & \new_[73508]_ ;
  assign \new_[73512]_  = A199 & A166;
  assign \new_[73515]_  = A201 & ~A200;
  assign \new_[73516]_  = \new_[73515]_  & \new_[73512]_ ;
  assign \new_[73517]_  = \new_[73516]_  & \new_[73509]_ ;
  assign \new_[73521]_  = A233 & ~A232;
  assign \new_[73522]_  = A203 & \new_[73521]_ ;
  assign \new_[73525]_  = ~A299 & A298;
  assign \new_[73528]_  = A302 & A300;
  assign \new_[73529]_  = \new_[73528]_  & \new_[73525]_ ;
  assign \new_[73530]_  = \new_[73529]_  & \new_[73522]_ ;
  assign \new_[73534]_  = ~A168 & A169;
  assign \new_[73535]_  = A170 & \new_[73534]_ ;
  assign \new_[73538]_  = A199 & A166;
  assign \new_[73541]_  = A201 & ~A200;
  assign \new_[73542]_  = \new_[73541]_  & \new_[73538]_ ;
  assign \new_[73543]_  = \new_[73542]_  & \new_[73535]_ ;
  assign \new_[73547]_  = A233 & ~A232;
  assign \new_[73548]_  = A203 & \new_[73547]_ ;
  assign \new_[73551]_  = ~A266 & A265;
  assign \new_[73554]_  = A268 & A267;
  assign \new_[73555]_  = \new_[73554]_  & \new_[73551]_ ;
  assign \new_[73556]_  = \new_[73555]_  & \new_[73548]_ ;
  assign \new_[73560]_  = ~A168 & A169;
  assign \new_[73561]_  = A170 & \new_[73560]_ ;
  assign \new_[73564]_  = A199 & A166;
  assign \new_[73567]_  = A201 & ~A200;
  assign \new_[73568]_  = \new_[73567]_  & \new_[73564]_ ;
  assign \new_[73569]_  = \new_[73568]_  & \new_[73561]_ ;
  assign \new_[73573]_  = A233 & ~A232;
  assign \new_[73574]_  = A203 & \new_[73573]_ ;
  assign \new_[73577]_  = ~A266 & A265;
  assign \new_[73580]_  = A269 & A267;
  assign \new_[73581]_  = \new_[73580]_  & \new_[73577]_ ;
  assign \new_[73582]_  = \new_[73581]_  & \new_[73574]_ ;
  assign \new_[73586]_  = A167 & A169;
  assign \new_[73587]_  = ~A170 & \new_[73586]_ ;
  assign \new_[73590]_  = A199 & A166;
  assign \new_[73593]_  = A232 & A200;
  assign \new_[73594]_  = \new_[73593]_  & \new_[73590]_ ;
  assign \new_[73595]_  = \new_[73594]_  & \new_[73587]_ ;
  assign \new_[73599]_  = ~A268 & A265;
  assign \new_[73600]_  = A233 & \new_[73599]_ ;
  assign \new_[73603]_  = ~A299 & ~A269;
  assign \new_[73606]_  = ~A302 & ~A301;
  assign \new_[73607]_  = \new_[73606]_  & \new_[73603]_ ;
  assign \new_[73608]_  = \new_[73607]_  & \new_[73600]_ ;
  assign \new_[73612]_  = A167 & A169;
  assign \new_[73613]_  = ~A170 & \new_[73612]_ ;
  assign \new_[73616]_  = A199 & A166;
  assign \new_[73619]_  = ~A233 & A200;
  assign \new_[73620]_  = \new_[73619]_  & \new_[73616]_ ;
  assign \new_[73621]_  = \new_[73620]_  & \new_[73613]_ ;
  assign \new_[73625]_  = A265 & ~A236;
  assign \new_[73626]_  = ~A235 & \new_[73625]_ ;
  assign \new_[73629]_  = A298 & A266;
  assign \new_[73632]_  = ~A302 & ~A301;
  assign \new_[73633]_  = \new_[73632]_  & \new_[73629]_ ;
  assign \new_[73634]_  = \new_[73633]_  & \new_[73626]_ ;
  assign \new_[73638]_  = A167 & A169;
  assign \new_[73639]_  = ~A170 & \new_[73638]_ ;
  assign \new_[73642]_  = A199 & A166;
  assign \new_[73645]_  = ~A233 & A200;
  assign \new_[73646]_  = \new_[73645]_  & \new_[73642]_ ;
  assign \new_[73647]_  = \new_[73646]_  & \new_[73639]_ ;
  assign \new_[73651]_  = ~A266 & ~A236;
  assign \new_[73652]_  = ~A235 & \new_[73651]_ ;
  assign \new_[73655]_  = ~A269 & ~A268;
  assign \new_[73658]_  = ~A300 & A298;
  assign \new_[73659]_  = \new_[73658]_  & \new_[73655]_ ;
  assign \new_[73660]_  = \new_[73659]_  & \new_[73652]_ ;
  assign \new_[73664]_  = A167 & A169;
  assign \new_[73665]_  = ~A170 & \new_[73664]_ ;
  assign \new_[73668]_  = A199 & A166;
  assign \new_[73671]_  = ~A233 & A200;
  assign \new_[73672]_  = \new_[73671]_  & \new_[73668]_ ;
  assign \new_[73673]_  = \new_[73672]_  & \new_[73665]_ ;
  assign \new_[73677]_  = ~A266 & ~A236;
  assign \new_[73678]_  = ~A235 & \new_[73677]_ ;
  assign \new_[73681]_  = ~A269 & ~A268;
  assign \new_[73684]_  = A299 & A298;
  assign \new_[73685]_  = \new_[73684]_  & \new_[73681]_ ;
  assign \new_[73686]_  = \new_[73685]_  & \new_[73678]_ ;
  assign \new_[73690]_  = A167 & A169;
  assign \new_[73691]_  = ~A170 & \new_[73690]_ ;
  assign \new_[73694]_  = A199 & A166;
  assign \new_[73697]_  = ~A233 & A200;
  assign \new_[73698]_  = \new_[73697]_  & \new_[73694]_ ;
  assign \new_[73699]_  = \new_[73698]_  & \new_[73691]_ ;
  assign \new_[73703]_  = ~A266 & ~A236;
  assign \new_[73704]_  = ~A235 & \new_[73703]_ ;
  assign \new_[73707]_  = ~A269 & ~A268;
  assign \new_[73710]_  = ~A299 & ~A298;
  assign \new_[73711]_  = \new_[73710]_  & \new_[73707]_ ;
  assign \new_[73712]_  = \new_[73711]_  & \new_[73704]_ ;
  assign \new_[73716]_  = A167 & A169;
  assign \new_[73717]_  = ~A170 & \new_[73716]_ ;
  assign \new_[73720]_  = A199 & A166;
  assign \new_[73723]_  = ~A233 & A200;
  assign \new_[73724]_  = \new_[73723]_  & \new_[73720]_ ;
  assign \new_[73725]_  = \new_[73724]_  & \new_[73717]_ ;
  assign \new_[73729]_  = ~A266 & ~A236;
  assign \new_[73730]_  = ~A235 & \new_[73729]_ ;
  assign \new_[73733]_  = A298 & ~A267;
  assign \new_[73736]_  = ~A302 & ~A301;
  assign \new_[73737]_  = \new_[73736]_  & \new_[73733]_ ;
  assign \new_[73738]_  = \new_[73737]_  & \new_[73730]_ ;
  assign \new_[73742]_  = A167 & A169;
  assign \new_[73743]_  = ~A170 & \new_[73742]_ ;
  assign \new_[73746]_  = A199 & A166;
  assign \new_[73749]_  = ~A233 & A200;
  assign \new_[73750]_  = \new_[73749]_  & \new_[73746]_ ;
  assign \new_[73751]_  = \new_[73750]_  & \new_[73743]_ ;
  assign \new_[73755]_  = ~A265 & ~A236;
  assign \new_[73756]_  = ~A235 & \new_[73755]_ ;
  assign \new_[73759]_  = A298 & ~A266;
  assign \new_[73762]_  = ~A302 & ~A301;
  assign \new_[73763]_  = \new_[73762]_  & \new_[73759]_ ;
  assign \new_[73764]_  = \new_[73763]_  & \new_[73756]_ ;
  assign \new_[73768]_  = A167 & A169;
  assign \new_[73769]_  = ~A170 & \new_[73768]_ ;
  assign \new_[73772]_  = A199 & A166;
  assign \new_[73775]_  = ~A233 & A200;
  assign \new_[73776]_  = \new_[73775]_  & \new_[73772]_ ;
  assign \new_[73777]_  = \new_[73776]_  & \new_[73769]_ ;
  assign \new_[73781]_  = ~A268 & ~A266;
  assign \new_[73782]_  = ~A234 & \new_[73781]_ ;
  assign \new_[73785]_  = A298 & ~A269;
  assign \new_[73788]_  = ~A302 & ~A301;
  assign \new_[73789]_  = \new_[73788]_  & \new_[73785]_ ;
  assign \new_[73790]_  = \new_[73789]_  & \new_[73782]_ ;
  assign \new_[73794]_  = A167 & A169;
  assign \new_[73795]_  = ~A170 & \new_[73794]_ ;
  assign \new_[73798]_  = A199 & A166;
  assign \new_[73801]_  = A232 & A200;
  assign \new_[73802]_  = \new_[73801]_  & \new_[73798]_ ;
  assign \new_[73803]_  = \new_[73802]_  & \new_[73795]_ ;
  assign \new_[73807]_  = A235 & A234;
  assign \new_[73808]_  = ~A233 & \new_[73807]_ ;
  assign \new_[73811]_  = ~A299 & A298;
  assign \new_[73814]_  = A301 & A300;
  assign \new_[73815]_  = \new_[73814]_  & \new_[73811]_ ;
  assign \new_[73816]_  = \new_[73815]_  & \new_[73808]_ ;
  assign \new_[73820]_  = A167 & A169;
  assign \new_[73821]_  = ~A170 & \new_[73820]_ ;
  assign \new_[73824]_  = A199 & A166;
  assign \new_[73827]_  = A232 & A200;
  assign \new_[73828]_  = \new_[73827]_  & \new_[73824]_ ;
  assign \new_[73829]_  = \new_[73828]_  & \new_[73821]_ ;
  assign \new_[73833]_  = A235 & A234;
  assign \new_[73834]_  = ~A233 & \new_[73833]_ ;
  assign \new_[73837]_  = ~A299 & A298;
  assign \new_[73840]_  = A302 & A300;
  assign \new_[73841]_  = \new_[73840]_  & \new_[73837]_ ;
  assign \new_[73842]_  = \new_[73841]_  & \new_[73834]_ ;
  assign \new_[73846]_  = A167 & A169;
  assign \new_[73847]_  = ~A170 & \new_[73846]_ ;
  assign \new_[73850]_  = A199 & A166;
  assign \new_[73853]_  = A232 & A200;
  assign \new_[73854]_  = \new_[73853]_  & \new_[73850]_ ;
  assign \new_[73855]_  = \new_[73854]_  & \new_[73847]_ ;
  assign \new_[73859]_  = A235 & A234;
  assign \new_[73860]_  = ~A233 & \new_[73859]_ ;
  assign \new_[73863]_  = ~A266 & A265;
  assign \new_[73866]_  = A268 & A267;
  assign \new_[73867]_  = \new_[73866]_  & \new_[73863]_ ;
  assign \new_[73868]_  = \new_[73867]_  & \new_[73860]_ ;
  assign \new_[73872]_  = A167 & A169;
  assign \new_[73873]_  = ~A170 & \new_[73872]_ ;
  assign \new_[73876]_  = A199 & A166;
  assign \new_[73879]_  = A232 & A200;
  assign \new_[73880]_  = \new_[73879]_  & \new_[73876]_ ;
  assign \new_[73881]_  = \new_[73880]_  & \new_[73873]_ ;
  assign \new_[73885]_  = A235 & A234;
  assign \new_[73886]_  = ~A233 & \new_[73885]_ ;
  assign \new_[73889]_  = ~A266 & A265;
  assign \new_[73892]_  = A269 & A267;
  assign \new_[73893]_  = \new_[73892]_  & \new_[73889]_ ;
  assign \new_[73894]_  = \new_[73893]_  & \new_[73886]_ ;
  assign \new_[73898]_  = A167 & A169;
  assign \new_[73899]_  = ~A170 & \new_[73898]_ ;
  assign \new_[73902]_  = A199 & A166;
  assign \new_[73905]_  = A232 & A200;
  assign \new_[73906]_  = \new_[73905]_  & \new_[73902]_ ;
  assign \new_[73907]_  = \new_[73906]_  & \new_[73899]_ ;
  assign \new_[73911]_  = A236 & A234;
  assign \new_[73912]_  = ~A233 & \new_[73911]_ ;
  assign \new_[73915]_  = ~A299 & A298;
  assign \new_[73918]_  = A301 & A300;
  assign \new_[73919]_  = \new_[73918]_  & \new_[73915]_ ;
  assign \new_[73920]_  = \new_[73919]_  & \new_[73912]_ ;
  assign \new_[73924]_  = A167 & A169;
  assign \new_[73925]_  = ~A170 & \new_[73924]_ ;
  assign \new_[73928]_  = A199 & A166;
  assign \new_[73931]_  = A232 & A200;
  assign \new_[73932]_  = \new_[73931]_  & \new_[73928]_ ;
  assign \new_[73933]_  = \new_[73932]_  & \new_[73925]_ ;
  assign \new_[73937]_  = A236 & A234;
  assign \new_[73938]_  = ~A233 & \new_[73937]_ ;
  assign \new_[73941]_  = ~A299 & A298;
  assign \new_[73944]_  = A302 & A300;
  assign \new_[73945]_  = \new_[73944]_  & \new_[73941]_ ;
  assign \new_[73946]_  = \new_[73945]_  & \new_[73938]_ ;
  assign \new_[73950]_  = A167 & A169;
  assign \new_[73951]_  = ~A170 & \new_[73950]_ ;
  assign \new_[73954]_  = A199 & A166;
  assign \new_[73957]_  = A232 & A200;
  assign \new_[73958]_  = \new_[73957]_  & \new_[73954]_ ;
  assign \new_[73959]_  = \new_[73958]_  & \new_[73951]_ ;
  assign \new_[73963]_  = A236 & A234;
  assign \new_[73964]_  = ~A233 & \new_[73963]_ ;
  assign \new_[73967]_  = ~A266 & A265;
  assign \new_[73970]_  = A268 & A267;
  assign \new_[73971]_  = \new_[73970]_  & \new_[73967]_ ;
  assign \new_[73972]_  = \new_[73971]_  & \new_[73964]_ ;
  assign \new_[73976]_  = A167 & A169;
  assign \new_[73977]_  = ~A170 & \new_[73976]_ ;
  assign \new_[73980]_  = A199 & A166;
  assign \new_[73983]_  = A232 & A200;
  assign \new_[73984]_  = \new_[73983]_  & \new_[73980]_ ;
  assign \new_[73985]_  = \new_[73984]_  & \new_[73977]_ ;
  assign \new_[73989]_  = A236 & A234;
  assign \new_[73990]_  = ~A233 & \new_[73989]_ ;
  assign \new_[73993]_  = ~A266 & A265;
  assign \new_[73996]_  = A269 & A267;
  assign \new_[73997]_  = \new_[73996]_  & \new_[73993]_ ;
  assign \new_[73998]_  = \new_[73997]_  & \new_[73990]_ ;
  assign \new_[74002]_  = A167 & A169;
  assign \new_[74003]_  = ~A170 & \new_[74002]_ ;
  assign \new_[74006]_  = A199 & A166;
  assign \new_[74009]_  = ~A232 & A200;
  assign \new_[74010]_  = \new_[74009]_  & \new_[74006]_ ;
  assign \new_[74011]_  = \new_[74010]_  & \new_[74003]_ ;
  assign \new_[74015]_  = ~A268 & ~A266;
  assign \new_[74016]_  = ~A233 & \new_[74015]_ ;
  assign \new_[74019]_  = A298 & ~A269;
  assign \new_[74022]_  = ~A302 & ~A301;
  assign \new_[74023]_  = \new_[74022]_  & \new_[74019]_ ;
  assign \new_[74024]_  = \new_[74023]_  & \new_[74016]_ ;
  assign \new_[74028]_  = A167 & A169;
  assign \new_[74029]_  = ~A170 & \new_[74028]_ ;
  assign \new_[74032]_  = ~A200 & A166;
  assign \new_[74035]_  = ~A203 & ~A202;
  assign \new_[74036]_  = \new_[74035]_  & \new_[74032]_ ;
  assign \new_[74037]_  = \new_[74036]_  & \new_[74029]_ ;
  assign \new_[74041]_  = A265 & A233;
  assign \new_[74042]_  = A232 & \new_[74041]_ ;
  assign \new_[74045]_  = ~A269 & ~A268;
  assign \new_[74048]_  = ~A300 & ~A299;
  assign \new_[74049]_  = \new_[74048]_  & \new_[74045]_ ;
  assign \new_[74050]_  = \new_[74049]_  & \new_[74042]_ ;
  assign \new_[74054]_  = A167 & A169;
  assign \new_[74055]_  = ~A170 & \new_[74054]_ ;
  assign \new_[74058]_  = ~A200 & A166;
  assign \new_[74061]_  = ~A203 & ~A202;
  assign \new_[74062]_  = \new_[74061]_  & \new_[74058]_ ;
  assign \new_[74063]_  = \new_[74062]_  & \new_[74055]_ ;
  assign \new_[74067]_  = A265 & A233;
  assign \new_[74068]_  = A232 & \new_[74067]_ ;
  assign \new_[74071]_  = ~A269 & ~A268;
  assign \new_[74074]_  = A299 & A298;
  assign \new_[74075]_  = \new_[74074]_  & \new_[74071]_ ;
  assign \new_[74076]_  = \new_[74075]_  & \new_[74068]_ ;
  assign \new_[74080]_  = A167 & A169;
  assign \new_[74081]_  = ~A170 & \new_[74080]_ ;
  assign \new_[74084]_  = ~A200 & A166;
  assign \new_[74087]_  = ~A203 & ~A202;
  assign \new_[74088]_  = \new_[74087]_  & \new_[74084]_ ;
  assign \new_[74089]_  = \new_[74088]_  & \new_[74081]_ ;
  assign \new_[74093]_  = A265 & A233;
  assign \new_[74094]_  = A232 & \new_[74093]_ ;
  assign \new_[74097]_  = ~A269 & ~A268;
  assign \new_[74100]_  = ~A299 & ~A298;
  assign \new_[74101]_  = \new_[74100]_  & \new_[74097]_ ;
  assign \new_[74102]_  = \new_[74101]_  & \new_[74094]_ ;
  assign \new_[74106]_  = A167 & A169;
  assign \new_[74107]_  = ~A170 & \new_[74106]_ ;
  assign \new_[74110]_  = ~A200 & A166;
  assign \new_[74113]_  = ~A203 & ~A202;
  assign \new_[74114]_  = \new_[74113]_  & \new_[74110]_ ;
  assign \new_[74115]_  = \new_[74114]_  & \new_[74107]_ ;
  assign \new_[74119]_  = A265 & A233;
  assign \new_[74120]_  = A232 & \new_[74119]_ ;
  assign \new_[74123]_  = ~A299 & ~A267;
  assign \new_[74126]_  = ~A302 & ~A301;
  assign \new_[74127]_  = \new_[74126]_  & \new_[74123]_ ;
  assign \new_[74128]_  = \new_[74127]_  & \new_[74120]_ ;
  assign \new_[74132]_  = A167 & A169;
  assign \new_[74133]_  = ~A170 & \new_[74132]_ ;
  assign \new_[74136]_  = ~A200 & A166;
  assign \new_[74139]_  = ~A203 & ~A202;
  assign \new_[74140]_  = \new_[74139]_  & \new_[74136]_ ;
  assign \new_[74141]_  = \new_[74140]_  & \new_[74133]_ ;
  assign \new_[74145]_  = A265 & A233;
  assign \new_[74146]_  = A232 & \new_[74145]_ ;
  assign \new_[74149]_  = ~A299 & A266;
  assign \new_[74152]_  = ~A302 & ~A301;
  assign \new_[74153]_  = \new_[74152]_  & \new_[74149]_ ;
  assign \new_[74154]_  = \new_[74153]_  & \new_[74146]_ ;
  assign \new_[74158]_  = A167 & A169;
  assign \new_[74159]_  = ~A170 & \new_[74158]_ ;
  assign \new_[74162]_  = ~A200 & A166;
  assign \new_[74165]_  = ~A203 & ~A202;
  assign \new_[74166]_  = \new_[74165]_  & \new_[74162]_ ;
  assign \new_[74167]_  = \new_[74166]_  & \new_[74159]_ ;
  assign \new_[74171]_  = ~A265 & A233;
  assign \new_[74172]_  = A232 & \new_[74171]_ ;
  assign \new_[74175]_  = ~A299 & ~A266;
  assign \new_[74178]_  = ~A302 & ~A301;
  assign \new_[74179]_  = \new_[74178]_  & \new_[74175]_ ;
  assign \new_[74180]_  = \new_[74179]_  & \new_[74172]_ ;
  assign \new_[74184]_  = A167 & A169;
  assign \new_[74185]_  = ~A170 & \new_[74184]_ ;
  assign \new_[74188]_  = ~A200 & A166;
  assign \new_[74191]_  = ~A203 & ~A202;
  assign \new_[74192]_  = \new_[74191]_  & \new_[74188]_ ;
  assign \new_[74193]_  = \new_[74192]_  & \new_[74185]_ ;
  assign \new_[74197]_  = ~A236 & ~A235;
  assign \new_[74198]_  = ~A233 & \new_[74197]_ ;
  assign \new_[74201]_  = A266 & A265;
  assign \new_[74204]_  = ~A300 & A298;
  assign \new_[74205]_  = \new_[74204]_  & \new_[74201]_ ;
  assign \new_[74206]_  = \new_[74205]_  & \new_[74198]_ ;
  assign \new_[74210]_  = A167 & A169;
  assign \new_[74211]_  = ~A170 & \new_[74210]_ ;
  assign \new_[74214]_  = ~A200 & A166;
  assign \new_[74217]_  = ~A203 & ~A202;
  assign \new_[74218]_  = \new_[74217]_  & \new_[74214]_ ;
  assign \new_[74219]_  = \new_[74218]_  & \new_[74211]_ ;
  assign \new_[74223]_  = ~A236 & ~A235;
  assign \new_[74224]_  = ~A233 & \new_[74223]_ ;
  assign \new_[74227]_  = A266 & A265;
  assign \new_[74230]_  = A299 & A298;
  assign \new_[74231]_  = \new_[74230]_  & \new_[74227]_ ;
  assign \new_[74232]_  = \new_[74231]_  & \new_[74224]_ ;
  assign \new_[74236]_  = A167 & A169;
  assign \new_[74237]_  = ~A170 & \new_[74236]_ ;
  assign \new_[74240]_  = ~A200 & A166;
  assign \new_[74243]_  = ~A203 & ~A202;
  assign \new_[74244]_  = \new_[74243]_  & \new_[74240]_ ;
  assign \new_[74245]_  = \new_[74244]_  & \new_[74237]_ ;
  assign \new_[74249]_  = ~A236 & ~A235;
  assign \new_[74250]_  = ~A233 & \new_[74249]_ ;
  assign \new_[74253]_  = A266 & A265;
  assign \new_[74256]_  = ~A299 & ~A298;
  assign \new_[74257]_  = \new_[74256]_  & \new_[74253]_ ;
  assign \new_[74258]_  = \new_[74257]_  & \new_[74250]_ ;
  assign \new_[74262]_  = A167 & A169;
  assign \new_[74263]_  = ~A170 & \new_[74262]_ ;
  assign \new_[74266]_  = ~A200 & A166;
  assign \new_[74269]_  = ~A203 & ~A202;
  assign \new_[74270]_  = \new_[74269]_  & \new_[74266]_ ;
  assign \new_[74271]_  = \new_[74270]_  & \new_[74263]_ ;
  assign \new_[74275]_  = ~A236 & ~A235;
  assign \new_[74276]_  = ~A233 & \new_[74275]_ ;
  assign \new_[74279]_  = ~A267 & ~A266;
  assign \new_[74282]_  = ~A300 & A298;
  assign \new_[74283]_  = \new_[74282]_  & \new_[74279]_ ;
  assign \new_[74284]_  = \new_[74283]_  & \new_[74276]_ ;
  assign \new_[74288]_  = A167 & A169;
  assign \new_[74289]_  = ~A170 & \new_[74288]_ ;
  assign \new_[74292]_  = ~A200 & A166;
  assign \new_[74295]_  = ~A203 & ~A202;
  assign \new_[74296]_  = \new_[74295]_  & \new_[74292]_ ;
  assign \new_[74297]_  = \new_[74296]_  & \new_[74289]_ ;
  assign \new_[74301]_  = ~A236 & ~A235;
  assign \new_[74302]_  = ~A233 & \new_[74301]_ ;
  assign \new_[74305]_  = ~A267 & ~A266;
  assign \new_[74308]_  = A299 & A298;
  assign \new_[74309]_  = \new_[74308]_  & \new_[74305]_ ;
  assign \new_[74310]_  = \new_[74309]_  & \new_[74302]_ ;
  assign \new_[74314]_  = A167 & A169;
  assign \new_[74315]_  = ~A170 & \new_[74314]_ ;
  assign \new_[74318]_  = ~A200 & A166;
  assign \new_[74321]_  = ~A203 & ~A202;
  assign \new_[74322]_  = \new_[74321]_  & \new_[74318]_ ;
  assign \new_[74323]_  = \new_[74322]_  & \new_[74315]_ ;
  assign \new_[74327]_  = ~A236 & ~A235;
  assign \new_[74328]_  = ~A233 & \new_[74327]_ ;
  assign \new_[74331]_  = ~A267 & ~A266;
  assign \new_[74334]_  = ~A299 & ~A298;
  assign \new_[74335]_  = \new_[74334]_  & \new_[74331]_ ;
  assign \new_[74336]_  = \new_[74335]_  & \new_[74328]_ ;
  assign \new_[74340]_  = A167 & A169;
  assign \new_[74341]_  = ~A170 & \new_[74340]_ ;
  assign \new_[74344]_  = ~A200 & A166;
  assign \new_[74347]_  = ~A203 & ~A202;
  assign \new_[74348]_  = \new_[74347]_  & \new_[74344]_ ;
  assign \new_[74349]_  = \new_[74348]_  & \new_[74341]_ ;
  assign \new_[74353]_  = ~A236 & ~A235;
  assign \new_[74354]_  = ~A233 & \new_[74353]_ ;
  assign \new_[74357]_  = ~A266 & ~A265;
  assign \new_[74360]_  = ~A300 & A298;
  assign \new_[74361]_  = \new_[74360]_  & \new_[74357]_ ;
  assign \new_[74362]_  = \new_[74361]_  & \new_[74354]_ ;
  assign \new_[74366]_  = A167 & A169;
  assign \new_[74367]_  = ~A170 & \new_[74366]_ ;
  assign \new_[74370]_  = ~A200 & A166;
  assign \new_[74373]_  = ~A203 & ~A202;
  assign \new_[74374]_  = \new_[74373]_  & \new_[74370]_ ;
  assign \new_[74375]_  = \new_[74374]_  & \new_[74367]_ ;
  assign \new_[74379]_  = ~A236 & ~A235;
  assign \new_[74380]_  = ~A233 & \new_[74379]_ ;
  assign \new_[74383]_  = ~A266 & ~A265;
  assign \new_[74386]_  = A299 & A298;
  assign \new_[74387]_  = \new_[74386]_  & \new_[74383]_ ;
  assign \new_[74388]_  = \new_[74387]_  & \new_[74380]_ ;
  assign \new_[74392]_  = A167 & A169;
  assign \new_[74393]_  = ~A170 & \new_[74392]_ ;
  assign \new_[74396]_  = ~A200 & A166;
  assign \new_[74399]_  = ~A203 & ~A202;
  assign \new_[74400]_  = \new_[74399]_  & \new_[74396]_ ;
  assign \new_[74401]_  = \new_[74400]_  & \new_[74393]_ ;
  assign \new_[74405]_  = ~A236 & ~A235;
  assign \new_[74406]_  = ~A233 & \new_[74405]_ ;
  assign \new_[74409]_  = ~A266 & ~A265;
  assign \new_[74412]_  = ~A299 & ~A298;
  assign \new_[74413]_  = \new_[74412]_  & \new_[74409]_ ;
  assign \new_[74414]_  = \new_[74413]_  & \new_[74406]_ ;
  assign \new_[74418]_  = A167 & A169;
  assign \new_[74419]_  = ~A170 & \new_[74418]_ ;
  assign \new_[74422]_  = ~A200 & A166;
  assign \new_[74425]_  = ~A203 & ~A202;
  assign \new_[74426]_  = \new_[74425]_  & \new_[74422]_ ;
  assign \new_[74427]_  = \new_[74426]_  & \new_[74419]_ ;
  assign \new_[74431]_  = A265 & ~A234;
  assign \new_[74432]_  = ~A233 & \new_[74431]_ ;
  assign \new_[74435]_  = A298 & A266;
  assign \new_[74438]_  = ~A302 & ~A301;
  assign \new_[74439]_  = \new_[74438]_  & \new_[74435]_ ;
  assign \new_[74440]_  = \new_[74439]_  & \new_[74432]_ ;
  assign \new_[74444]_  = A167 & A169;
  assign \new_[74445]_  = ~A170 & \new_[74444]_ ;
  assign \new_[74448]_  = ~A200 & A166;
  assign \new_[74451]_  = ~A203 & ~A202;
  assign \new_[74452]_  = \new_[74451]_  & \new_[74448]_ ;
  assign \new_[74453]_  = \new_[74452]_  & \new_[74445]_ ;
  assign \new_[74457]_  = ~A266 & ~A234;
  assign \new_[74458]_  = ~A233 & \new_[74457]_ ;
  assign \new_[74461]_  = ~A269 & ~A268;
  assign \new_[74464]_  = ~A300 & A298;
  assign \new_[74465]_  = \new_[74464]_  & \new_[74461]_ ;
  assign \new_[74466]_  = \new_[74465]_  & \new_[74458]_ ;
  assign \new_[74470]_  = A167 & A169;
  assign \new_[74471]_  = ~A170 & \new_[74470]_ ;
  assign \new_[74474]_  = ~A200 & A166;
  assign \new_[74477]_  = ~A203 & ~A202;
  assign \new_[74478]_  = \new_[74477]_  & \new_[74474]_ ;
  assign \new_[74479]_  = \new_[74478]_  & \new_[74471]_ ;
  assign \new_[74483]_  = ~A266 & ~A234;
  assign \new_[74484]_  = ~A233 & \new_[74483]_ ;
  assign \new_[74487]_  = ~A269 & ~A268;
  assign \new_[74490]_  = A299 & A298;
  assign \new_[74491]_  = \new_[74490]_  & \new_[74487]_ ;
  assign \new_[74492]_  = \new_[74491]_  & \new_[74484]_ ;
  assign \new_[74496]_  = A167 & A169;
  assign \new_[74497]_  = ~A170 & \new_[74496]_ ;
  assign \new_[74500]_  = ~A200 & A166;
  assign \new_[74503]_  = ~A203 & ~A202;
  assign \new_[74504]_  = \new_[74503]_  & \new_[74500]_ ;
  assign \new_[74505]_  = \new_[74504]_  & \new_[74497]_ ;
  assign \new_[74509]_  = ~A266 & ~A234;
  assign \new_[74510]_  = ~A233 & \new_[74509]_ ;
  assign \new_[74513]_  = ~A269 & ~A268;
  assign \new_[74516]_  = ~A299 & ~A298;
  assign \new_[74517]_  = \new_[74516]_  & \new_[74513]_ ;
  assign \new_[74518]_  = \new_[74517]_  & \new_[74510]_ ;
  assign \new_[74522]_  = A167 & A169;
  assign \new_[74523]_  = ~A170 & \new_[74522]_ ;
  assign \new_[74526]_  = ~A200 & A166;
  assign \new_[74529]_  = ~A203 & ~A202;
  assign \new_[74530]_  = \new_[74529]_  & \new_[74526]_ ;
  assign \new_[74531]_  = \new_[74530]_  & \new_[74523]_ ;
  assign \new_[74535]_  = ~A266 & ~A234;
  assign \new_[74536]_  = ~A233 & \new_[74535]_ ;
  assign \new_[74539]_  = A298 & ~A267;
  assign \new_[74542]_  = ~A302 & ~A301;
  assign \new_[74543]_  = \new_[74542]_  & \new_[74539]_ ;
  assign \new_[74544]_  = \new_[74543]_  & \new_[74536]_ ;
  assign \new_[74548]_  = A167 & A169;
  assign \new_[74549]_  = ~A170 & \new_[74548]_ ;
  assign \new_[74552]_  = ~A200 & A166;
  assign \new_[74555]_  = ~A203 & ~A202;
  assign \new_[74556]_  = \new_[74555]_  & \new_[74552]_ ;
  assign \new_[74557]_  = \new_[74556]_  & \new_[74549]_ ;
  assign \new_[74561]_  = ~A265 & ~A234;
  assign \new_[74562]_  = ~A233 & \new_[74561]_ ;
  assign \new_[74565]_  = A298 & ~A266;
  assign \new_[74568]_  = ~A302 & ~A301;
  assign \new_[74569]_  = \new_[74568]_  & \new_[74565]_ ;
  assign \new_[74570]_  = \new_[74569]_  & \new_[74562]_ ;
  assign \new_[74574]_  = A167 & A169;
  assign \new_[74575]_  = ~A170 & \new_[74574]_ ;
  assign \new_[74578]_  = ~A200 & A166;
  assign \new_[74581]_  = ~A203 & ~A202;
  assign \new_[74582]_  = \new_[74581]_  & \new_[74578]_ ;
  assign \new_[74583]_  = \new_[74582]_  & \new_[74575]_ ;
  assign \new_[74587]_  = A265 & ~A233;
  assign \new_[74588]_  = ~A232 & \new_[74587]_ ;
  assign \new_[74591]_  = A298 & A266;
  assign \new_[74594]_  = ~A302 & ~A301;
  assign \new_[74595]_  = \new_[74594]_  & \new_[74591]_ ;
  assign \new_[74596]_  = \new_[74595]_  & \new_[74588]_ ;
  assign \new_[74600]_  = A167 & A169;
  assign \new_[74601]_  = ~A170 & \new_[74600]_ ;
  assign \new_[74604]_  = ~A200 & A166;
  assign \new_[74607]_  = ~A203 & ~A202;
  assign \new_[74608]_  = \new_[74607]_  & \new_[74604]_ ;
  assign \new_[74609]_  = \new_[74608]_  & \new_[74601]_ ;
  assign \new_[74613]_  = ~A266 & ~A233;
  assign \new_[74614]_  = ~A232 & \new_[74613]_ ;
  assign \new_[74617]_  = ~A269 & ~A268;
  assign \new_[74620]_  = ~A300 & A298;
  assign \new_[74621]_  = \new_[74620]_  & \new_[74617]_ ;
  assign \new_[74622]_  = \new_[74621]_  & \new_[74614]_ ;
  assign \new_[74626]_  = A167 & A169;
  assign \new_[74627]_  = ~A170 & \new_[74626]_ ;
  assign \new_[74630]_  = ~A200 & A166;
  assign \new_[74633]_  = ~A203 & ~A202;
  assign \new_[74634]_  = \new_[74633]_  & \new_[74630]_ ;
  assign \new_[74635]_  = \new_[74634]_  & \new_[74627]_ ;
  assign \new_[74639]_  = ~A266 & ~A233;
  assign \new_[74640]_  = ~A232 & \new_[74639]_ ;
  assign \new_[74643]_  = ~A269 & ~A268;
  assign \new_[74646]_  = A299 & A298;
  assign \new_[74647]_  = \new_[74646]_  & \new_[74643]_ ;
  assign \new_[74648]_  = \new_[74647]_  & \new_[74640]_ ;
  assign \new_[74652]_  = A167 & A169;
  assign \new_[74653]_  = ~A170 & \new_[74652]_ ;
  assign \new_[74656]_  = ~A200 & A166;
  assign \new_[74659]_  = ~A203 & ~A202;
  assign \new_[74660]_  = \new_[74659]_  & \new_[74656]_ ;
  assign \new_[74661]_  = \new_[74660]_  & \new_[74653]_ ;
  assign \new_[74665]_  = ~A266 & ~A233;
  assign \new_[74666]_  = ~A232 & \new_[74665]_ ;
  assign \new_[74669]_  = ~A269 & ~A268;
  assign \new_[74672]_  = ~A299 & ~A298;
  assign \new_[74673]_  = \new_[74672]_  & \new_[74669]_ ;
  assign \new_[74674]_  = \new_[74673]_  & \new_[74666]_ ;
  assign \new_[74678]_  = A167 & A169;
  assign \new_[74679]_  = ~A170 & \new_[74678]_ ;
  assign \new_[74682]_  = ~A200 & A166;
  assign \new_[74685]_  = ~A203 & ~A202;
  assign \new_[74686]_  = \new_[74685]_  & \new_[74682]_ ;
  assign \new_[74687]_  = \new_[74686]_  & \new_[74679]_ ;
  assign \new_[74691]_  = ~A266 & ~A233;
  assign \new_[74692]_  = ~A232 & \new_[74691]_ ;
  assign \new_[74695]_  = A298 & ~A267;
  assign \new_[74698]_  = ~A302 & ~A301;
  assign \new_[74699]_  = \new_[74698]_  & \new_[74695]_ ;
  assign \new_[74700]_  = \new_[74699]_  & \new_[74692]_ ;
  assign \new_[74704]_  = A167 & A169;
  assign \new_[74705]_  = ~A170 & \new_[74704]_ ;
  assign \new_[74708]_  = ~A200 & A166;
  assign \new_[74711]_  = ~A203 & ~A202;
  assign \new_[74712]_  = \new_[74711]_  & \new_[74708]_ ;
  assign \new_[74713]_  = \new_[74712]_  & \new_[74705]_ ;
  assign \new_[74717]_  = ~A265 & ~A233;
  assign \new_[74718]_  = ~A232 & \new_[74717]_ ;
  assign \new_[74721]_  = A298 & ~A266;
  assign \new_[74724]_  = ~A302 & ~A301;
  assign \new_[74725]_  = \new_[74724]_  & \new_[74721]_ ;
  assign \new_[74726]_  = \new_[74725]_  & \new_[74718]_ ;
  assign \new_[74730]_  = A167 & A169;
  assign \new_[74731]_  = ~A170 & \new_[74730]_ ;
  assign \new_[74734]_  = ~A200 & A166;
  assign \new_[74737]_  = A232 & ~A201;
  assign \new_[74738]_  = \new_[74737]_  & \new_[74734]_ ;
  assign \new_[74739]_  = \new_[74738]_  & \new_[74731]_ ;
  assign \new_[74743]_  = ~A268 & A265;
  assign \new_[74744]_  = A233 & \new_[74743]_ ;
  assign \new_[74747]_  = ~A299 & ~A269;
  assign \new_[74750]_  = ~A302 & ~A301;
  assign \new_[74751]_  = \new_[74750]_  & \new_[74747]_ ;
  assign \new_[74752]_  = \new_[74751]_  & \new_[74744]_ ;
  assign \new_[74756]_  = A167 & A169;
  assign \new_[74757]_  = ~A170 & \new_[74756]_ ;
  assign \new_[74760]_  = ~A200 & A166;
  assign \new_[74763]_  = ~A233 & ~A201;
  assign \new_[74764]_  = \new_[74763]_  & \new_[74760]_ ;
  assign \new_[74765]_  = \new_[74764]_  & \new_[74757]_ ;
  assign \new_[74769]_  = A265 & ~A236;
  assign \new_[74770]_  = ~A235 & \new_[74769]_ ;
  assign \new_[74773]_  = A298 & A266;
  assign \new_[74776]_  = ~A302 & ~A301;
  assign \new_[74777]_  = \new_[74776]_  & \new_[74773]_ ;
  assign \new_[74778]_  = \new_[74777]_  & \new_[74770]_ ;
  assign \new_[74782]_  = A167 & A169;
  assign \new_[74783]_  = ~A170 & \new_[74782]_ ;
  assign \new_[74786]_  = ~A200 & A166;
  assign \new_[74789]_  = ~A233 & ~A201;
  assign \new_[74790]_  = \new_[74789]_  & \new_[74786]_ ;
  assign \new_[74791]_  = \new_[74790]_  & \new_[74783]_ ;
  assign \new_[74795]_  = ~A266 & ~A236;
  assign \new_[74796]_  = ~A235 & \new_[74795]_ ;
  assign \new_[74799]_  = ~A269 & ~A268;
  assign \new_[74802]_  = ~A300 & A298;
  assign \new_[74803]_  = \new_[74802]_  & \new_[74799]_ ;
  assign \new_[74804]_  = \new_[74803]_  & \new_[74796]_ ;
  assign \new_[74808]_  = A167 & A169;
  assign \new_[74809]_  = ~A170 & \new_[74808]_ ;
  assign \new_[74812]_  = ~A200 & A166;
  assign \new_[74815]_  = ~A233 & ~A201;
  assign \new_[74816]_  = \new_[74815]_  & \new_[74812]_ ;
  assign \new_[74817]_  = \new_[74816]_  & \new_[74809]_ ;
  assign \new_[74821]_  = ~A266 & ~A236;
  assign \new_[74822]_  = ~A235 & \new_[74821]_ ;
  assign \new_[74825]_  = ~A269 & ~A268;
  assign \new_[74828]_  = A299 & A298;
  assign \new_[74829]_  = \new_[74828]_  & \new_[74825]_ ;
  assign \new_[74830]_  = \new_[74829]_  & \new_[74822]_ ;
  assign \new_[74834]_  = A167 & A169;
  assign \new_[74835]_  = ~A170 & \new_[74834]_ ;
  assign \new_[74838]_  = ~A200 & A166;
  assign \new_[74841]_  = ~A233 & ~A201;
  assign \new_[74842]_  = \new_[74841]_  & \new_[74838]_ ;
  assign \new_[74843]_  = \new_[74842]_  & \new_[74835]_ ;
  assign \new_[74847]_  = ~A266 & ~A236;
  assign \new_[74848]_  = ~A235 & \new_[74847]_ ;
  assign \new_[74851]_  = ~A269 & ~A268;
  assign \new_[74854]_  = ~A299 & ~A298;
  assign \new_[74855]_  = \new_[74854]_  & \new_[74851]_ ;
  assign \new_[74856]_  = \new_[74855]_  & \new_[74848]_ ;
  assign \new_[74860]_  = A167 & A169;
  assign \new_[74861]_  = ~A170 & \new_[74860]_ ;
  assign \new_[74864]_  = ~A200 & A166;
  assign \new_[74867]_  = ~A233 & ~A201;
  assign \new_[74868]_  = \new_[74867]_  & \new_[74864]_ ;
  assign \new_[74869]_  = \new_[74868]_  & \new_[74861]_ ;
  assign \new_[74873]_  = ~A266 & ~A236;
  assign \new_[74874]_  = ~A235 & \new_[74873]_ ;
  assign \new_[74877]_  = A298 & ~A267;
  assign \new_[74880]_  = ~A302 & ~A301;
  assign \new_[74881]_  = \new_[74880]_  & \new_[74877]_ ;
  assign \new_[74882]_  = \new_[74881]_  & \new_[74874]_ ;
  assign \new_[74886]_  = A167 & A169;
  assign \new_[74887]_  = ~A170 & \new_[74886]_ ;
  assign \new_[74890]_  = ~A200 & A166;
  assign \new_[74893]_  = ~A233 & ~A201;
  assign \new_[74894]_  = \new_[74893]_  & \new_[74890]_ ;
  assign \new_[74895]_  = \new_[74894]_  & \new_[74887]_ ;
  assign \new_[74899]_  = ~A265 & ~A236;
  assign \new_[74900]_  = ~A235 & \new_[74899]_ ;
  assign \new_[74903]_  = A298 & ~A266;
  assign \new_[74906]_  = ~A302 & ~A301;
  assign \new_[74907]_  = \new_[74906]_  & \new_[74903]_ ;
  assign \new_[74908]_  = \new_[74907]_  & \new_[74900]_ ;
  assign \new_[74912]_  = A167 & A169;
  assign \new_[74913]_  = ~A170 & \new_[74912]_ ;
  assign \new_[74916]_  = ~A200 & A166;
  assign \new_[74919]_  = ~A233 & ~A201;
  assign \new_[74920]_  = \new_[74919]_  & \new_[74916]_ ;
  assign \new_[74921]_  = \new_[74920]_  & \new_[74913]_ ;
  assign \new_[74925]_  = ~A268 & ~A266;
  assign \new_[74926]_  = ~A234 & \new_[74925]_ ;
  assign \new_[74929]_  = A298 & ~A269;
  assign \new_[74932]_  = ~A302 & ~A301;
  assign \new_[74933]_  = \new_[74932]_  & \new_[74929]_ ;
  assign \new_[74934]_  = \new_[74933]_  & \new_[74926]_ ;
  assign \new_[74938]_  = A167 & A169;
  assign \new_[74939]_  = ~A170 & \new_[74938]_ ;
  assign \new_[74942]_  = ~A200 & A166;
  assign \new_[74945]_  = A232 & ~A201;
  assign \new_[74946]_  = \new_[74945]_  & \new_[74942]_ ;
  assign \new_[74947]_  = \new_[74946]_  & \new_[74939]_ ;
  assign \new_[74951]_  = A235 & A234;
  assign \new_[74952]_  = ~A233 & \new_[74951]_ ;
  assign \new_[74955]_  = ~A299 & A298;
  assign \new_[74958]_  = A301 & A300;
  assign \new_[74959]_  = \new_[74958]_  & \new_[74955]_ ;
  assign \new_[74960]_  = \new_[74959]_  & \new_[74952]_ ;
  assign \new_[74964]_  = A167 & A169;
  assign \new_[74965]_  = ~A170 & \new_[74964]_ ;
  assign \new_[74968]_  = ~A200 & A166;
  assign \new_[74971]_  = A232 & ~A201;
  assign \new_[74972]_  = \new_[74971]_  & \new_[74968]_ ;
  assign \new_[74973]_  = \new_[74972]_  & \new_[74965]_ ;
  assign \new_[74977]_  = A235 & A234;
  assign \new_[74978]_  = ~A233 & \new_[74977]_ ;
  assign \new_[74981]_  = ~A299 & A298;
  assign \new_[74984]_  = A302 & A300;
  assign \new_[74985]_  = \new_[74984]_  & \new_[74981]_ ;
  assign \new_[74986]_  = \new_[74985]_  & \new_[74978]_ ;
  assign \new_[74990]_  = A167 & A169;
  assign \new_[74991]_  = ~A170 & \new_[74990]_ ;
  assign \new_[74994]_  = ~A200 & A166;
  assign \new_[74997]_  = A232 & ~A201;
  assign \new_[74998]_  = \new_[74997]_  & \new_[74994]_ ;
  assign \new_[74999]_  = \new_[74998]_  & \new_[74991]_ ;
  assign \new_[75003]_  = A235 & A234;
  assign \new_[75004]_  = ~A233 & \new_[75003]_ ;
  assign \new_[75007]_  = ~A266 & A265;
  assign \new_[75010]_  = A268 & A267;
  assign \new_[75011]_  = \new_[75010]_  & \new_[75007]_ ;
  assign \new_[75012]_  = \new_[75011]_  & \new_[75004]_ ;
  assign \new_[75016]_  = A167 & A169;
  assign \new_[75017]_  = ~A170 & \new_[75016]_ ;
  assign \new_[75020]_  = ~A200 & A166;
  assign \new_[75023]_  = A232 & ~A201;
  assign \new_[75024]_  = \new_[75023]_  & \new_[75020]_ ;
  assign \new_[75025]_  = \new_[75024]_  & \new_[75017]_ ;
  assign \new_[75029]_  = A235 & A234;
  assign \new_[75030]_  = ~A233 & \new_[75029]_ ;
  assign \new_[75033]_  = ~A266 & A265;
  assign \new_[75036]_  = A269 & A267;
  assign \new_[75037]_  = \new_[75036]_  & \new_[75033]_ ;
  assign \new_[75038]_  = \new_[75037]_  & \new_[75030]_ ;
  assign \new_[75042]_  = A167 & A169;
  assign \new_[75043]_  = ~A170 & \new_[75042]_ ;
  assign \new_[75046]_  = ~A200 & A166;
  assign \new_[75049]_  = A232 & ~A201;
  assign \new_[75050]_  = \new_[75049]_  & \new_[75046]_ ;
  assign \new_[75051]_  = \new_[75050]_  & \new_[75043]_ ;
  assign \new_[75055]_  = A236 & A234;
  assign \new_[75056]_  = ~A233 & \new_[75055]_ ;
  assign \new_[75059]_  = ~A299 & A298;
  assign \new_[75062]_  = A301 & A300;
  assign \new_[75063]_  = \new_[75062]_  & \new_[75059]_ ;
  assign \new_[75064]_  = \new_[75063]_  & \new_[75056]_ ;
  assign \new_[75068]_  = A167 & A169;
  assign \new_[75069]_  = ~A170 & \new_[75068]_ ;
  assign \new_[75072]_  = ~A200 & A166;
  assign \new_[75075]_  = A232 & ~A201;
  assign \new_[75076]_  = \new_[75075]_  & \new_[75072]_ ;
  assign \new_[75077]_  = \new_[75076]_  & \new_[75069]_ ;
  assign \new_[75081]_  = A236 & A234;
  assign \new_[75082]_  = ~A233 & \new_[75081]_ ;
  assign \new_[75085]_  = ~A299 & A298;
  assign \new_[75088]_  = A302 & A300;
  assign \new_[75089]_  = \new_[75088]_  & \new_[75085]_ ;
  assign \new_[75090]_  = \new_[75089]_  & \new_[75082]_ ;
  assign \new_[75094]_  = A167 & A169;
  assign \new_[75095]_  = ~A170 & \new_[75094]_ ;
  assign \new_[75098]_  = ~A200 & A166;
  assign \new_[75101]_  = A232 & ~A201;
  assign \new_[75102]_  = \new_[75101]_  & \new_[75098]_ ;
  assign \new_[75103]_  = \new_[75102]_  & \new_[75095]_ ;
  assign \new_[75107]_  = A236 & A234;
  assign \new_[75108]_  = ~A233 & \new_[75107]_ ;
  assign \new_[75111]_  = ~A266 & A265;
  assign \new_[75114]_  = A268 & A267;
  assign \new_[75115]_  = \new_[75114]_  & \new_[75111]_ ;
  assign \new_[75116]_  = \new_[75115]_  & \new_[75108]_ ;
  assign \new_[75120]_  = A167 & A169;
  assign \new_[75121]_  = ~A170 & \new_[75120]_ ;
  assign \new_[75124]_  = ~A200 & A166;
  assign \new_[75127]_  = A232 & ~A201;
  assign \new_[75128]_  = \new_[75127]_  & \new_[75124]_ ;
  assign \new_[75129]_  = \new_[75128]_  & \new_[75121]_ ;
  assign \new_[75133]_  = A236 & A234;
  assign \new_[75134]_  = ~A233 & \new_[75133]_ ;
  assign \new_[75137]_  = ~A266 & A265;
  assign \new_[75140]_  = A269 & A267;
  assign \new_[75141]_  = \new_[75140]_  & \new_[75137]_ ;
  assign \new_[75142]_  = \new_[75141]_  & \new_[75134]_ ;
  assign \new_[75146]_  = A167 & A169;
  assign \new_[75147]_  = ~A170 & \new_[75146]_ ;
  assign \new_[75150]_  = ~A200 & A166;
  assign \new_[75153]_  = ~A232 & ~A201;
  assign \new_[75154]_  = \new_[75153]_  & \new_[75150]_ ;
  assign \new_[75155]_  = \new_[75154]_  & \new_[75147]_ ;
  assign \new_[75159]_  = ~A268 & ~A266;
  assign \new_[75160]_  = ~A233 & \new_[75159]_ ;
  assign \new_[75163]_  = A298 & ~A269;
  assign \new_[75166]_  = ~A302 & ~A301;
  assign \new_[75167]_  = \new_[75166]_  & \new_[75163]_ ;
  assign \new_[75168]_  = \new_[75167]_  & \new_[75160]_ ;
  assign \new_[75172]_  = A167 & A169;
  assign \new_[75173]_  = ~A170 & \new_[75172]_ ;
  assign \new_[75176]_  = ~A199 & A166;
  assign \new_[75179]_  = A232 & ~A200;
  assign \new_[75180]_  = \new_[75179]_  & \new_[75176]_ ;
  assign \new_[75181]_  = \new_[75180]_  & \new_[75173]_ ;
  assign \new_[75185]_  = ~A268 & A265;
  assign \new_[75186]_  = A233 & \new_[75185]_ ;
  assign \new_[75189]_  = ~A299 & ~A269;
  assign \new_[75192]_  = ~A302 & ~A301;
  assign \new_[75193]_  = \new_[75192]_  & \new_[75189]_ ;
  assign \new_[75194]_  = \new_[75193]_  & \new_[75186]_ ;
  assign \new_[75198]_  = A167 & A169;
  assign \new_[75199]_  = ~A170 & \new_[75198]_ ;
  assign \new_[75202]_  = ~A199 & A166;
  assign \new_[75205]_  = ~A233 & ~A200;
  assign \new_[75206]_  = \new_[75205]_  & \new_[75202]_ ;
  assign \new_[75207]_  = \new_[75206]_  & \new_[75199]_ ;
  assign \new_[75211]_  = A265 & ~A236;
  assign \new_[75212]_  = ~A235 & \new_[75211]_ ;
  assign \new_[75215]_  = A298 & A266;
  assign \new_[75218]_  = ~A302 & ~A301;
  assign \new_[75219]_  = \new_[75218]_  & \new_[75215]_ ;
  assign \new_[75220]_  = \new_[75219]_  & \new_[75212]_ ;
  assign \new_[75224]_  = A167 & A169;
  assign \new_[75225]_  = ~A170 & \new_[75224]_ ;
  assign \new_[75228]_  = ~A199 & A166;
  assign \new_[75231]_  = ~A233 & ~A200;
  assign \new_[75232]_  = \new_[75231]_  & \new_[75228]_ ;
  assign \new_[75233]_  = \new_[75232]_  & \new_[75225]_ ;
  assign \new_[75237]_  = ~A266 & ~A236;
  assign \new_[75238]_  = ~A235 & \new_[75237]_ ;
  assign \new_[75241]_  = ~A269 & ~A268;
  assign \new_[75244]_  = ~A300 & A298;
  assign \new_[75245]_  = \new_[75244]_  & \new_[75241]_ ;
  assign \new_[75246]_  = \new_[75245]_  & \new_[75238]_ ;
  assign \new_[75250]_  = A167 & A169;
  assign \new_[75251]_  = ~A170 & \new_[75250]_ ;
  assign \new_[75254]_  = ~A199 & A166;
  assign \new_[75257]_  = ~A233 & ~A200;
  assign \new_[75258]_  = \new_[75257]_  & \new_[75254]_ ;
  assign \new_[75259]_  = \new_[75258]_  & \new_[75251]_ ;
  assign \new_[75263]_  = ~A266 & ~A236;
  assign \new_[75264]_  = ~A235 & \new_[75263]_ ;
  assign \new_[75267]_  = ~A269 & ~A268;
  assign \new_[75270]_  = A299 & A298;
  assign \new_[75271]_  = \new_[75270]_  & \new_[75267]_ ;
  assign \new_[75272]_  = \new_[75271]_  & \new_[75264]_ ;
  assign \new_[75276]_  = A167 & A169;
  assign \new_[75277]_  = ~A170 & \new_[75276]_ ;
  assign \new_[75280]_  = ~A199 & A166;
  assign \new_[75283]_  = ~A233 & ~A200;
  assign \new_[75284]_  = \new_[75283]_  & \new_[75280]_ ;
  assign \new_[75285]_  = \new_[75284]_  & \new_[75277]_ ;
  assign \new_[75289]_  = ~A266 & ~A236;
  assign \new_[75290]_  = ~A235 & \new_[75289]_ ;
  assign \new_[75293]_  = ~A269 & ~A268;
  assign \new_[75296]_  = ~A299 & ~A298;
  assign \new_[75297]_  = \new_[75296]_  & \new_[75293]_ ;
  assign \new_[75298]_  = \new_[75297]_  & \new_[75290]_ ;
  assign \new_[75302]_  = A167 & A169;
  assign \new_[75303]_  = ~A170 & \new_[75302]_ ;
  assign \new_[75306]_  = ~A199 & A166;
  assign \new_[75309]_  = ~A233 & ~A200;
  assign \new_[75310]_  = \new_[75309]_  & \new_[75306]_ ;
  assign \new_[75311]_  = \new_[75310]_  & \new_[75303]_ ;
  assign \new_[75315]_  = ~A266 & ~A236;
  assign \new_[75316]_  = ~A235 & \new_[75315]_ ;
  assign \new_[75319]_  = A298 & ~A267;
  assign \new_[75322]_  = ~A302 & ~A301;
  assign \new_[75323]_  = \new_[75322]_  & \new_[75319]_ ;
  assign \new_[75324]_  = \new_[75323]_  & \new_[75316]_ ;
  assign \new_[75328]_  = A167 & A169;
  assign \new_[75329]_  = ~A170 & \new_[75328]_ ;
  assign \new_[75332]_  = ~A199 & A166;
  assign \new_[75335]_  = ~A233 & ~A200;
  assign \new_[75336]_  = \new_[75335]_  & \new_[75332]_ ;
  assign \new_[75337]_  = \new_[75336]_  & \new_[75329]_ ;
  assign \new_[75341]_  = ~A265 & ~A236;
  assign \new_[75342]_  = ~A235 & \new_[75341]_ ;
  assign \new_[75345]_  = A298 & ~A266;
  assign \new_[75348]_  = ~A302 & ~A301;
  assign \new_[75349]_  = \new_[75348]_  & \new_[75345]_ ;
  assign \new_[75350]_  = \new_[75349]_  & \new_[75342]_ ;
  assign \new_[75354]_  = A167 & A169;
  assign \new_[75355]_  = ~A170 & \new_[75354]_ ;
  assign \new_[75358]_  = ~A199 & A166;
  assign \new_[75361]_  = ~A233 & ~A200;
  assign \new_[75362]_  = \new_[75361]_  & \new_[75358]_ ;
  assign \new_[75363]_  = \new_[75362]_  & \new_[75355]_ ;
  assign \new_[75367]_  = ~A268 & ~A266;
  assign \new_[75368]_  = ~A234 & \new_[75367]_ ;
  assign \new_[75371]_  = A298 & ~A269;
  assign \new_[75374]_  = ~A302 & ~A301;
  assign \new_[75375]_  = \new_[75374]_  & \new_[75371]_ ;
  assign \new_[75376]_  = \new_[75375]_  & \new_[75368]_ ;
  assign \new_[75380]_  = A167 & A169;
  assign \new_[75381]_  = ~A170 & \new_[75380]_ ;
  assign \new_[75384]_  = ~A199 & A166;
  assign \new_[75387]_  = A232 & ~A200;
  assign \new_[75388]_  = \new_[75387]_  & \new_[75384]_ ;
  assign \new_[75389]_  = \new_[75388]_  & \new_[75381]_ ;
  assign \new_[75393]_  = A235 & A234;
  assign \new_[75394]_  = ~A233 & \new_[75393]_ ;
  assign \new_[75397]_  = ~A299 & A298;
  assign \new_[75400]_  = A301 & A300;
  assign \new_[75401]_  = \new_[75400]_  & \new_[75397]_ ;
  assign \new_[75402]_  = \new_[75401]_  & \new_[75394]_ ;
  assign \new_[75406]_  = A167 & A169;
  assign \new_[75407]_  = ~A170 & \new_[75406]_ ;
  assign \new_[75410]_  = ~A199 & A166;
  assign \new_[75413]_  = A232 & ~A200;
  assign \new_[75414]_  = \new_[75413]_  & \new_[75410]_ ;
  assign \new_[75415]_  = \new_[75414]_  & \new_[75407]_ ;
  assign \new_[75419]_  = A235 & A234;
  assign \new_[75420]_  = ~A233 & \new_[75419]_ ;
  assign \new_[75423]_  = ~A299 & A298;
  assign \new_[75426]_  = A302 & A300;
  assign \new_[75427]_  = \new_[75426]_  & \new_[75423]_ ;
  assign \new_[75428]_  = \new_[75427]_  & \new_[75420]_ ;
  assign \new_[75432]_  = A167 & A169;
  assign \new_[75433]_  = ~A170 & \new_[75432]_ ;
  assign \new_[75436]_  = ~A199 & A166;
  assign \new_[75439]_  = A232 & ~A200;
  assign \new_[75440]_  = \new_[75439]_  & \new_[75436]_ ;
  assign \new_[75441]_  = \new_[75440]_  & \new_[75433]_ ;
  assign \new_[75445]_  = A235 & A234;
  assign \new_[75446]_  = ~A233 & \new_[75445]_ ;
  assign \new_[75449]_  = ~A266 & A265;
  assign \new_[75452]_  = A268 & A267;
  assign \new_[75453]_  = \new_[75452]_  & \new_[75449]_ ;
  assign \new_[75454]_  = \new_[75453]_  & \new_[75446]_ ;
  assign \new_[75458]_  = A167 & A169;
  assign \new_[75459]_  = ~A170 & \new_[75458]_ ;
  assign \new_[75462]_  = ~A199 & A166;
  assign \new_[75465]_  = A232 & ~A200;
  assign \new_[75466]_  = \new_[75465]_  & \new_[75462]_ ;
  assign \new_[75467]_  = \new_[75466]_  & \new_[75459]_ ;
  assign \new_[75471]_  = A235 & A234;
  assign \new_[75472]_  = ~A233 & \new_[75471]_ ;
  assign \new_[75475]_  = ~A266 & A265;
  assign \new_[75478]_  = A269 & A267;
  assign \new_[75479]_  = \new_[75478]_  & \new_[75475]_ ;
  assign \new_[75480]_  = \new_[75479]_  & \new_[75472]_ ;
  assign \new_[75484]_  = A167 & A169;
  assign \new_[75485]_  = ~A170 & \new_[75484]_ ;
  assign \new_[75488]_  = ~A199 & A166;
  assign \new_[75491]_  = A232 & ~A200;
  assign \new_[75492]_  = \new_[75491]_  & \new_[75488]_ ;
  assign \new_[75493]_  = \new_[75492]_  & \new_[75485]_ ;
  assign \new_[75497]_  = A236 & A234;
  assign \new_[75498]_  = ~A233 & \new_[75497]_ ;
  assign \new_[75501]_  = ~A299 & A298;
  assign \new_[75504]_  = A301 & A300;
  assign \new_[75505]_  = \new_[75504]_  & \new_[75501]_ ;
  assign \new_[75506]_  = \new_[75505]_  & \new_[75498]_ ;
  assign \new_[75510]_  = A167 & A169;
  assign \new_[75511]_  = ~A170 & \new_[75510]_ ;
  assign \new_[75514]_  = ~A199 & A166;
  assign \new_[75517]_  = A232 & ~A200;
  assign \new_[75518]_  = \new_[75517]_  & \new_[75514]_ ;
  assign \new_[75519]_  = \new_[75518]_  & \new_[75511]_ ;
  assign \new_[75523]_  = A236 & A234;
  assign \new_[75524]_  = ~A233 & \new_[75523]_ ;
  assign \new_[75527]_  = ~A299 & A298;
  assign \new_[75530]_  = A302 & A300;
  assign \new_[75531]_  = \new_[75530]_  & \new_[75527]_ ;
  assign \new_[75532]_  = \new_[75531]_  & \new_[75524]_ ;
  assign \new_[75536]_  = A167 & A169;
  assign \new_[75537]_  = ~A170 & \new_[75536]_ ;
  assign \new_[75540]_  = ~A199 & A166;
  assign \new_[75543]_  = A232 & ~A200;
  assign \new_[75544]_  = \new_[75543]_  & \new_[75540]_ ;
  assign \new_[75545]_  = \new_[75544]_  & \new_[75537]_ ;
  assign \new_[75549]_  = A236 & A234;
  assign \new_[75550]_  = ~A233 & \new_[75549]_ ;
  assign \new_[75553]_  = ~A266 & A265;
  assign \new_[75556]_  = A268 & A267;
  assign \new_[75557]_  = \new_[75556]_  & \new_[75553]_ ;
  assign \new_[75558]_  = \new_[75557]_  & \new_[75550]_ ;
  assign \new_[75562]_  = A167 & A169;
  assign \new_[75563]_  = ~A170 & \new_[75562]_ ;
  assign \new_[75566]_  = ~A199 & A166;
  assign \new_[75569]_  = A232 & ~A200;
  assign \new_[75570]_  = \new_[75569]_  & \new_[75566]_ ;
  assign \new_[75571]_  = \new_[75570]_  & \new_[75563]_ ;
  assign \new_[75575]_  = A236 & A234;
  assign \new_[75576]_  = ~A233 & \new_[75575]_ ;
  assign \new_[75579]_  = ~A266 & A265;
  assign \new_[75582]_  = A269 & A267;
  assign \new_[75583]_  = \new_[75582]_  & \new_[75579]_ ;
  assign \new_[75584]_  = \new_[75583]_  & \new_[75576]_ ;
  assign \new_[75588]_  = A167 & A169;
  assign \new_[75589]_  = ~A170 & \new_[75588]_ ;
  assign \new_[75592]_  = ~A199 & A166;
  assign \new_[75595]_  = ~A232 & ~A200;
  assign \new_[75596]_  = \new_[75595]_  & \new_[75592]_ ;
  assign \new_[75597]_  = \new_[75596]_  & \new_[75589]_ ;
  assign \new_[75601]_  = ~A268 & ~A266;
  assign \new_[75602]_  = ~A233 & \new_[75601]_ ;
  assign \new_[75605]_  = A298 & ~A269;
  assign \new_[75608]_  = ~A302 & ~A301;
  assign \new_[75609]_  = \new_[75608]_  & \new_[75605]_ ;
  assign \new_[75610]_  = \new_[75609]_  & \new_[75602]_ ;
  assign \new_[75614]_  = ~A167 & A169;
  assign \new_[75615]_  = ~A170 & \new_[75614]_ ;
  assign \new_[75618]_  = A199 & ~A166;
  assign \new_[75621]_  = A232 & A200;
  assign \new_[75622]_  = \new_[75621]_  & \new_[75618]_ ;
  assign \new_[75623]_  = \new_[75622]_  & \new_[75615]_ ;
  assign \new_[75627]_  = ~A268 & A265;
  assign \new_[75628]_  = A233 & \new_[75627]_ ;
  assign \new_[75631]_  = ~A299 & ~A269;
  assign \new_[75634]_  = ~A302 & ~A301;
  assign \new_[75635]_  = \new_[75634]_  & \new_[75631]_ ;
  assign \new_[75636]_  = \new_[75635]_  & \new_[75628]_ ;
  assign \new_[75640]_  = ~A167 & A169;
  assign \new_[75641]_  = ~A170 & \new_[75640]_ ;
  assign \new_[75644]_  = A199 & ~A166;
  assign \new_[75647]_  = ~A233 & A200;
  assign \new_[75648]_  = \new_[75647]_  & \new_[75644]_ ;
  assign \new_[75649]_  = \new_[75648]_  & \new_[75641]_ ;
  assign \new_[75653]_  = A265 & ~A236;
  assign \new_[75654]_  = ~A235 & \new_[75653]_ ;
  assign \new_[75657]_  = A298 & A266;
  assign \new_[75660]_  = ~A302 & ~A301;
  assign \new_[75661]_  = \new_[75660]_  & \new_[75657]_ ;
  assign \new_[75662]_  = \new_[75661]_  & \new_[75654]_ ;
  assign \new_[75666]_  = ~A167 & A169;
  assign \new_[75667]_  = ~A170 & \new_[75666]_ ;
  assign \new_[75670]_  = A199 & ~A166;
  assign \new_[75673]_  = ~A233 & A200;
  assign \new_[75674]_  = \new_[75673]_  & \new_[75670]_ ;
  assign \new_[75675]_  = \new_[75674]_  & \new_[75667]_ ;
  assign \new_[75679]_  = ~A266 & ~A236;
  assign \new_[75680]_  = ~A235 & \new_[75679]_ ;
  assign \new_[75683]_  = ~A269 & ~A268;
  assign \new_[75686]_  = ~A300 & A298;
  assign \new_[75687]_  = \new_[75686]_  & \new_[75683]_ ;
  assign \new_[75688]_  = \new_[75687]_  & \new_[75680]_ ;
  assign \new_[75692]_  = ~A167 & A169;
  assign \new_[75693]_  = ~A170 & \new_[75692]_ ;
  assign \new_[75696]_  = A199 & ~A166;
  assign \new_[75699]_  = ~A233 & A200;
  assign \new_[75700]_  = \new_[75699]_  & \new_[75696]_ ;
  assign \new_[75701]_  = \new_[75700]_  & \new_[75693]_ ;
  assign \new_[75705]_  = ~A266 & ~A236;
  assign \new_[75706]_  = ~A235 & \new_[75705]_ ;
  assign \new_[75709]_  = ~A269 & ~A268;
  assign \new_[75712]_  = A299 & A298;
  assign \new_[75713]_  = \new_[75712]_  & \new_[75709]_ ;
  assign \new_[75714]_  = \new_[75713]_  & \new_[75706]_ ;
  assign \new_[75718]_  = ~A167 & A169;
  assign \new_[75719]_  = ~A170 & \new_[75718]_ ;
  assign \new_[75722]_  = A199 & ~A166;
  assign \new_[75725]_  = ~A233 & A200;
  assign \new_[75726]_  = \new_[75725]_  & \new_[75722]_ ;
  assign \new_[75727]_  = \new_[75726]_  & \new_[75719]_ ;
  assign \new_[75731]_  = ~A266 & ~A236;
  assign \new_[75732]_  = ~A235 & \new_[75731]_ ;
  assign \new_[75735]_  = ~A269 & ~A268;
  assign \new_[75738]_  = ~A299 & ~A298;
  assign \new_[75739]_  = \new_[75738]_  & \new_[75735]_ ;
  assign \new_[75740]_  = \new_[75739]_  & \new_[75732]_ ;
  assign \new_[75744]_  = ~A167 & A169;
  assign \new_[75745]_  = ~A170 & \new_[75744]_ ;
  assign \new_[75748]_  = A199 & ~A166;
  assign \new_[75751]_  = ~A233 & A200;
  assign \new_[75752]_  = \new_[75751]_  & \new_[75748]_ ;
  assign \new_[75753]_  = \new_[75752]_  & \new_[75745]_ ;
  assign \new_[75757]_  = ~A266 & ~A236;
  assign \new_[75758]_  = ~A235 & \new_[75757]_ ;
  assign \new_[75761]_  = A298 & ~A267;
  assign \new_[75764]_  = ~A302 & ~A301;
  assign \new_[75765]_  = \new_[75764]_  & \new_[75761]_ ;
  assign \new_[75766]_  = \new_[75765]_  & \new_[75758]_ ;
  assign \new_[75770]_  = ~A167 & A169;
  assign \new_[75771]_  = ~A170 & \new_[75770]_ ;
  assign \new_[75774]_  = A199 & ~A166;
  assign \new_[75777]_  = ~A233 & A200;
  assign \new_[75778]_  = \new_[75777]_  & \new_[75774]_ ;
  assign \new_[75779]_  = \new_[75778]_  & \new_[75771]_ ;
  assign \new_[75783]_  = ~A265 & ~A236;
  assign \new_[75784]_  = ~A235 & \new_[75783]_ ;
  assign \new_[75787]_  = A298 & ~A266;
  assign \new_[75790]_  = ~A302 & ~A301;
  assign \new_[75791]_  = \new_[75790]_  & \new_[75787]_ ;
  assign \new_[75792]_  = \new_[75791]_  & \new_[75784]_ ;
  assign \new_[75796]_  = ~A167 & A169;
  assign \new_[75797]_  = ~A170 & \new_[75796]_ ;
  assign \new_[75800]_  = A199 & ~A166;
  assign \new_[75803]_  = ~A233 & A200;
  assign \new_[75804]_  = \new_[75803]_  & \new_[75800]_ ;
  assign \new_[75805]_  = \new_[75804]_  & \new_[75797]_ ;
  assign \new_[75809]_  = ~A268 & ~A266;
  assign \new_[75810]_  = ~A234 & \new_[75809]_ ;
  assign \new_[75813]_  = A298 & ~A269;
  assign \new_[75816]_  = ~A302 & ~A301;
  assign \new_[75817]_  = \new_[75816]_  & \new_[75813]_ ;
  assign \new_[75818]_  = \new_[75817]_  & \new_[75810]_ ;
  assign \new_[75822]_  = ~A167 & A169;
  assign \new_[75823]_  = ~A170 & \new_[75822]_ ;
  assign \new_[75826]_  = A199 & ~A166;
  assign \new_[75829]_  = A232 & A200;
  assign \new_[75830]_  = \new_[75829]_  & \new_[75826]_ ;
  assign \new_[75831]_  = \new_[75830]_  & \new_[75823]_ ;
  assign \new_[75835]_  = A235 & A234;
  assign \new_[75836]_  = ~A233 & \new_[75835]_ ;
  assign \new_[75839]_  = ~A299 & A298;
  assign \new_[75842]_  = A301 & A300;
  assign \new_[75843]_  = \new_[75842]_  & \new_[75839]_ ;
  assign \new_[75844]_  = \new_[75843]_  & \new_[75836]_ ;
  assign \new_[75848]_  = ~A167 & A169;
  assign \new_[75849]_  = ~A170 & \new_[75848]_ ;
  assign \new_[75852]_  = A199 & ~A166;
  assign \new_[75855]_  = A232 & A200;
  assign \new_[75856]_  = \new_[75855]_  & \new_[75852]_ ;
  assign \new_[75857]_  = \new_[75856]_  & \new_[75849]_ ;
  assign \new_[75861]_  = A235 & A234;
  assign \new_[75862]_  = ~A233 & \new_[75861]_ ;
  assign \new_[75865]_  = ~A299 & A298;
  assign \new_[75868]_  = A302 & A300;
  assign \new_[75869]_  = \new_[75868]_  & \new_[75865]_ ;
  assign \new_[75870]_  = \new_[75869]_  & \new_[75862]_ ;
  assign \new_[75874]_  = ~A167 & A169;
  assign \new_[75875]_  = ~A170 & \new_[75874]_ ;
  assign \new_[75878]_  = A199 & ~A166;
  assign \new_[75881]_  = A232 & A200;
  assign \new_[75882]_  = \new_[75881]_  & \new_[75878]_ ;
  assign \new_[75883]_  = \new_[75882]_  & \new_[75875]_ ;
  assign \new_[75887]_  = A235 & A234;
  assign \new_[75888]_  = ~A233 & \new_[75887]_ ;
  assign \new_[75891]_  = ~A266 & A265;
  assign \new_[75894]_  = A268 & A267;
  assign \new_[75895]_  = \new_[75894]_  & \new_[75891]_ ;
  assign \new_[75896]_  = \new_[75895]_  & \new_[75888]_ ;
  assign \new_[75900]_  = ~A167 & A169;
  assign \new_[75901]_  = ~A170 & \new_[75900]_ ;
  assign \new_[75904]_  = A199 & ~A166;
  assign \new_[75907]_  = A232 & A200;
  assign \new_[75908]_  = \new_[75907]_  & \new_[75904]_ ;
  assign \new_[75909]_  = \new_[75908]_  & \new_[75901]_ ;
  assign \new_[75913]_  = A235 & A234;
  assign \new_[75914]_  = ~A233 & \new_[75913]_ ;
  assign \new_[75917]_  = ~A266 & A265;
  assign \new_[75920]_  = A269 & A267;
  assign \new_[75921]_  = \new_[75920]_  & \new_[75917]_ ;
  assign \new_[75922]_  = \new_[75921]_  & \new_[75914]_ ;
  assign \new_[75926]_  = ~A167 & A169;
  assign \new_[75927]_  = ~A170 & \new_[75926]_ ;
  assign \new_[75930]_  = A199 & ~A166;
  assign \new_[75933]_  = A232 & A200;
  assign \new_[75934]_  = \new_[75933]_  & \new_[75930]_ ;
  assign \new_[75935]_  = \new_[75934]_  & \new_[75927]_ ;
  assign \new_[75939]_  = A236 & A234;
  assign \new_[75940]_  = ~A233 & \new_[75939]_ ;
  assign \new_[75943]_  = ~A299 & A298;
  assign \new_[75946]_  = A301 & A300;
  assign \new_[75947]_  = \new_[75946]_  & \new_[75943]_ ;
  assign \new_[75948]_  = \new_[75947]_  & \new_[75940]_ ;
  assign \new_[75952]_  = ~A167 & A169;
  assign \new_[75953]_  = ~A170 & \new_[75952]_ ;
  assign \new_[75956]_  = A199 & ~A166;
  assign \new_[75959]_  = A232 & A200;
  assign \new_[75960]_  = \new_[75959]_  & \new_[75956]_ ;
  assign \new_[75961]_  = \new_[75960]_  & \new_[75953]_ ;
  assign \new_[75965]_  = A236 & A234;
  assign \new_[75966]_  = ~A233 & \new_[75965]_ ;
  assign \new_[75969]_  = ~A299 & A298;
  assign \new_[75972]_  = A302 & A300;
  assign \new_[75973]_  = \new_[75972]_  & \new_[75969]_ ;
  assign \new_[75974]_  = \new_[75973]_  & \new_[75966]_ ;
  assign \new_[75978]_  = ~A167 & A169;
  assign \new_[75979]_  = ~A170 & \new_[75978]_ ;
  assign \new_[75982]_  = A199 & ~A166;
  assign \new_[75985]_  = A232 & A200;
  assign \new_[75986]_  = \new_[75985]_  & \new_[75982]_ ;
  assign \new_[75987]_  = \new_[75986]_  & \new_[75979]_ ;
  assign \new_[75991]_  = A236 & A234;
  assign \new_[75992]_  = ~A233 & \new_[75991]_ ;
  assign \new_[75995]_  = ~A266 & A265;
  assign \new_[75998]_  = A268 & A267;
  assign \new_[75999]_  = \new_[75998]_  & \new_[75995]_ ;
  assign \new_[76000]_  = \new_[75999]_  & \new_[75992]_ ;
  assign \new_[76004]_  = ~A167 & A169;
  assign \new_[76005]_  = ~A170 & \new_[76004]_ ;
  assign \new_[76008]_  = A199 & ~A166;
  assign \new_[76011]_  = A232 & A200;
  assign \new_[76012]_  = \new_[76011]_  & \new_[76008]_ ;
  assign \new_[76013]_  = \new_[76012]_  & \new_[76005]_ ;
  assign \new_[76017]_  = A236 & A234;
  assign \new_[76018]_  = ~A233 & \new_[76017]_ ;
  assign \new_[76021]_  = ~A266 & A265;
  assign \new_[76024]_  = A269 & A267;
  assign \new_[76025]_  = \new_[76024]_  & \new_[76021]_ ;
  assign \new_[76026]_  = \new_[76025]_  & \new_[76018]_ ;
  assign \new_[76030]_  = ~A167 & A169;
  assign \new_[76031]_  = ~A170 & \new_[76030]_ ;
  assign \new_[76034]_  = A199 & ~A166;
  assign \new_[76037]_  = ~A232 & A200;
  assign \new_[76038]_  = \new_[76037]_  & \new_[76034]_ ;
  assign \new_[76039]_  = \new_[76038]_  & \new_[76031]_ ;
  assign \new_[76043]_  = ~A268 & ~A266;
  assign \new_[76044]_  = ~A233 & \new_[76043]_ ;
  assign \new_[76047]_  = A298 & ~A269;
  assign \new_[76050]_  = ~A302 & ~A301;
  assign \new_[76051]_  = \new_[76050]_  & \new_[76047]_ ;
  assign \new_[76052]_  = \new_[76051]_  & \new_[76044]_ ;
  assign \new_[76056]_  = ~A167 & A169;
  assign \new_[76057]_  = ~A170 & \new_[76056]_ ;
  assign \new_[76060]_  = ~A200 & ~A166;
  assign \new_[76063]_  = ~A203 & ~A202;
  assign \new_[76064]_  = \new_[76063]_  & \new_[76060]_ ;
  assign \new_[76065]_  = \new_[76064]_  & \new_[76057]_ ;
  assign \new_[76069]_  = A265 & A233;
  assign \new_[76070]_  = A232 & \new_[76069]_ ;
  assign \new_[76073]_  = ~A269 & ~A268;
  assign \new_[76076]_  = ~A300 & ~A299;
  assign \new_[76077]_  = \new_[76076]_  & \new_[76073]_ ;
  assign \new_[76078]_  = \new_[76077]_  & \new_[76070]_ ;
  assign \new_[76082]_  = ~A167 & A169;
  assign \new_[76083]_  = ~A170 & \new_[76082]_ ;
  assign \new_[76086]_  = ~A200 & ~A166;
  assign \new_[76089]_  = ~A203 & ~A202;
  assign \new_[76090]_  = \new_[76089]_  & \new_[76086]_ ;
  assign \new_[76091]_  = \new_[76090]_  & \new_[76083]_ ;
  assign \new_[76095]_  = A265 & A233;
  assign \new_[76096]_  = A232 & \new_[76095]_ ;
  assign \new_[76099]_  = ~A269 & ~A268;
  assign \new_[76102]_  = A299 & A298;
  assign \new_[76103]_  = \new_[76102]_  & \new_[76099]_ ;
  assign \new_[76104]_  = \new_[76103]_  & \new_[76096]_ ;
  assign \new_[76108]_  = ~A167 & A169;
  assign \new_[76109]_  = ~A170 & \new_[76108]_ ;
  assign \new_[76112]_  = ~A200 & ~A166;
  assign \new_[76115]_  = ~A203 & ~A202;
  assign \new_[76116]_  = \new_[76115]_  & \new_[76112]_ ;
  assign \new_[76117]_  = \new_[76116]_  & \new_[76109]_ ;
  assign \new_[76121]_  = A265 & A233;
  assign \new_[76122]_  = A232 & \new_[76121]_ ;
  assign \new_[76125]_  = ~A269 & ~A268;
  assign \new_[76128]_  = ~A299 & ~A298;
  assign \new_[76129]_  = \new_[76128]_  & \new_[76125]_ ;
  assign \new_[76130]_  = \new_[76129]_  & \new_[76122]_ ;
  assign \new_[76134]_  = ~A167 & A169;
  assign \new_[76135]_  = ~A170 & \new_[76134]_ ;
  assign \new_[76138]_  = ~A200 & ~A166;
  assign \new_[76141]_  = ~A203 & ~A202;
  assign \new_[76142]_  = \new_[76141]_  & \new_[76138]_ ;
  assign \new_[76143]_  = \new_[76142]_  & \new_[76135]_ ;
  assign \new_[76147]_  = A265 & A233;
  assign \new_[76148]_  = A232 & \new_[76147]_ ;
  assign \new_[76151]_  = ~A299 & ~A267;
  assign \new_[76154]_  = ~A302 & ~A301;
  assign \new_[76155]_  = \new_[76154]_  & \new_[76151]_ ;
  assign \new_[76156]_  = \new_[76155]_  & \new_[76148]_ ;
  assign \new_[76160]_  = ~A167 & A169;
  assign \new_[76161]_  = ~A170 & \new_[76160]_ ;
  assign \new_[76164]_  = ~A200 & ~A166;
  assign \new_[76167]_  = ~A203 & ~A202;
  assign \new_[76168]_  = \new_[76167]_  & \new_[76164]_ ;
  assign \new_[76169]_  = \new_[76168]_  & \new_[76161]_ ;
  assign \new_[76173]_  = A265 & A233;
  assign \new_[76174]_  = A232 & \new_[76173]_ ;
  assign \new_[76177]_  = ~A299 & A266;
  assign \new_[76180]_  = ~A302 & ~A301;
  assign \new_[76181]_  = \new_[76180]_  & \new_[76177]_ ;
  assign \new_[76182]_  = \new_[76181]_  & \new_[76174]_ ;
  assign \new_[76186]_  = ~A167 & A169;
  assign \new_[76187]_  = ~A170 & \new_[76186]_ ;
  assign \new_[76190]_  = ~A200 & ~A166;
  assign \new_[76193]_  = ~A203 & ~A202;
  assign \new_[76194]_  = \new_[76193]_  & \new_[76190]_ ;
  assign \new_[76195]_  = \new_[76194]_  & \new_[76187]_ ;
  assign \new_[76199]_  = ~A265 & A233;
  assign \new_[76200]_  = A232 & \new_[76199]_ ;
  assign \new_[76203]_  = ~A299 & ~A266;
  assign \new_[76206]_  = ~A302 & ~A301;
  assign \new_[76207]_  = \new_[76206]_  & \new_[76203]_ ;
  assign \new_[76208]_  = \new_[76207]_  & \new_[76200]_ ;
  assign \new_[76212]_  = ~A167 & A169;
  assign \new_[76213]_  = ~A170 & \new_[76212]_ ;
  assign \new_[76216]_  = ~A200 & ~A166;
  assign \new_[76219]_  = ~A203 & ~A202;
  assign \new_[76220]_  = \new_[76219]_  & \new_[76216]_ ;
  assign \new_[76221]_  = \new_[76220]_  & \new_[76213]_ ;
  assign \new_[76225]_  = ~A236 & ~A235;
  assign \new_[76226]_  = ~A233 & \new_[76225]_ ;
  assign \new_[76229]_  = A266 & A265;
  assign \new_[76232]_  = ~A300 & A298;
  assign \new_[76233]_  = \new_[76232]_  & \new_[76229]_ ;
  assign \new_[76234]_  = \new_[76233]_  & \new_[76226]_ ;
  assign \new_[76238]_  = ~A167 & A169;
  assign \new_[76239]_  = ~A170 & \new_[76238]_ ;
  assign \new_[76242]_  = ~A200 & ~A166;
  assign \new_[76245]_  = ~A203 & ~A202;
  assign \new_[76246]_  = \new_[76245]_  & \new_[76242]_ ;
  assign \new_[76247]_  = \new_[76246]_  & \new_[76239]_ ;
  assign \new_[76251]_  = ~A236 & ~A235;
  assign \new_[76252]_  = ~A233 & \new_[76251]_ ;
  assign \new_[76255]_  = A266 & A265;
  assign \new_[76258]_  = A299 & A298;
  assign \new_[76259]_  = \new_[76258]_  & \new_[76255]_ ;
  assign \new_[76260]_  = \new_[76259]_  & \new_[76252]_ ;
  assign \new_[76264]_  = ~A167 & A169;
  assign \new_[76265]_  = ~A170 & \new_[76264]_ ;
  assign \new_[76268]_  = ~A200 & ~A166;
  assign \new_[76271]_  = ~A203 & ~A202;
  assign \new_[76272]_  = \new_[76271]_  & \new_[76268]_ ;
  assign \new_[76273]_  = \new_[76272]_  & \new_[76265]_ ;
  assign \new_[76277]_  = ~A236 & ~A235;
  assign \new_[76278]_  = ~A233 & \new_[76277]_ ;
  assign \new_[76281]_  = A266 & A265;
  assign \new_[76284]_  = ~A299 & ~A298;
  assign \new_[76285]_  = \new_[76284]_  & \new_[76281]_ ;
  assign \new_[76286]_  = \new_[76285]_  & \new_[76278]_ ;
  assign \new_[76290]_  = ~A167 & A169;
  assign \new_[76291]_  = ~A170 & \new_[76290]_ ;
  assign \new_[76294]_  = ~A200 & ~A166;
  assign \new_[76297]_  = ~A203 & ~A202;
  assign \new_[76298]_  = \new_[76297]_  & \new_[76294]_ ;
  assign \new_[76299]_  = \new_[76298]_  & \new_[76291]_ ;
  assign \new_[76303]_  = ~A236 & ~A235;
  assign \new_[76304]_  = ~A233 & \new_[76303]_ ;
  assign \new_[76307]_  = ~A267 & ~A266;
  assign \new_[76310]_  = ~A300 & A298;
  assign \new_[76311]_  = \new_[76310]_  & \new_[76307]_ ;
  assign \new_[76312]_  = \new_[76311]_  & \new_[76304]_ ;
  assign \new_[76316]_  = ~A167 & A169;
  assign \new_[76317]_  = ~A170 & \new_[76316]_ ;
  assign \new_[76320]_  = ~A200 & ~A166;
  assign \new_[76323]_  = ~A203 & ~A202;
  assign \new_[76324]_  = \new_[76323]_  & \new_[76320]_ ;
  assign \new_[76325]_  = \new_[76324]_  & \new_[76317]_ ;
  assign \new_[76329]_  = ~A236 & ~A235;
  assign \new_[76330]_  = ~A233 & \new_[76329]_ ;
  assign \new_[76333]_  = ~A267 & ~A266;
  assign \new_[76336]_  = A299 & A298;
  assign \new_[76337]_  = \new_[76336]_  & \new_[76333]_ ;
  assign \new_[76338]_  = \new_[76337]_  & \new_[76330]_ ;
  assign \new_[76342]_  = ~A167 & A169;
  assign \new_[76343]_  = ~A170 & \new_[76342]_ ;
  assign \new_[76346]_  = ~A200 & ~A166;
  assign \new_[76349]_  = ~A203 & ~A202;
  assign \new_[76350]_  = \new_[76349]_  & \new_[76346]_ ;
  assign \new_[76351]_  = \new_[76350]_  & \new_[76343]_ ;
  assign \new_[76355]_  = ~A236 & ~A235;
  assign \new_[76356]_  = ~A233 & \new_[76355]_ ;
  assign \new_[76359]_  = ~A267 & ~A266;
  assign \new_[76362]_  = ~A299 & ~A298;
  assign \new_[76363]_  = \new_[76362]_  & \new_[76359]_ ;
  assign \new_[76364]_  = \new_[76363]_  & \new_[76356]_ ;
  assign \new_[76368]_  = ~A167 & A169;
  assign \new_[76369]_  = ~A170 & \new_[76368]_ ;
  assign \new_[76372]_  = ~A200 & ~A166;
  assign \new_[76375]_  = ~A203 & ~A202;
  assign \new_[76376]_  = \new_[76375]_  & \new_[76372]_ ;
  assign \new_[76377]_  = \new_[76376]_  & \new_[76369]_ ;
  assign \new_[76381]_  = ~A236 & ~A235;
  assign \new_[76382]_  = ~A233 & \new_[76381]_ ;
  assign \new_[76385]_  = ~A266 & ~A265;
  assign \new_[76388]_  = ~A300 & A298;
  assign \new_[76389]_  = \new_[76388]_  & \new_[76385]_ ;
  assign \new_[76390]_  = \new_[76389]_  & \new_[76382]_ ;
  assign \new_[76394]_  = ~A167 & A169;
  assign \new_[76395]_  = ~A170 & \new_[76394]_ ;
  assign \new_[76398]_  = ~A200 & ~A166;
  assign \new_[76401]_  = ~A203 & ~A202;
  assign \new_[76402]_  = \new_[76401]_  & \new_[76398]_ ;
  assign \new_[76403]_  = \new_[76402]_  & \new_[76395]_ ;
  assign \new_[76407]_  = ~A236 & ~A235;
  assign \new_[76408]_  = ~A233 & \new_[76407]_ ;
  assign \new_[76411]_  = ~A266 & ~A265;
  assign \new_[76414]_  = A299 & A298;
  assign \new_[76415]_  = \new_[76414]_  & \new_[76411]_ ;
  assign \new_[76416]_  = \new_[76415]_  & \new_[76408]_ ;
  assign \new_[76420]_  = ~A167 & A169;
  assign \new_[76421]_  = ~A170 & \new_[76420]_ ;
  assign \new_[76424]_  = ~A200 & ~A166;
  assign \new_[76427]_  = ~A203 & ~A202;
  assign \new_[76428]_  = \new_[76427]_  & \new_[76424]_ ;
  assign \new_[76429]_  = \new_[76428]_  & \new_[76421]_ ;
  assign \new_[76433]_  = ~A236 & ~A235;
  assign \new_[76434]_  = ~A233 & \new_[76433]_ ;
  assign \new_[76437]_  = ~A266 & ~A265;
  assign \new_[76440]_  = ~A299 & ~A298;
  assign \new_[76441]_  = \new_[76440]_  & \new_[76437]_ ;
  assign \new_[76442]_  = \new_[76441]_  & \new_[76434]_ ;
  assign \new_[76446]_  = ~A167 & A169;
  assign \new_[76447]_  = ~A170 & \new_[76446]_ ;
  assign \new_[76450]_  = ~A200 & ~A166;
  assign \new_[76453]_  = ~A203 & ~A202;
  assign \new_[76454]_  = \new_[76453]_  & \new_[76450]_ ;
  assign \new_[76455]_  = \new_[76454]_  & \new_[76447]_ ;
  assign \new_[76459]_  = A265 & ~A234;
  assign \new_[76460]_  = ~A233 & \new_[76459]_ ;
  assign \new_[76463]_  = A298 & A266;
  assign \new_[76466]_  = ~A302 & ~A301;
  assign \new_[76467]_  = \new_[76466]_  & \new_[76463]_ ;
  assign \new_[76468]_  = \new_[76467]_  & \new_[76460]_ ;
  assign \new_[76472]_  = ~A167 & A169;
  assign \new_[76473]_  = ~A170 & \new_[76472]_ ;
  assign \new_[76476]_  = ~A200 & ~A166;
  assign \new_[76479]_  = ~A203 & ~A202;
  assign \new_[76480]_  = \new_[76479]_  & \new_[76476]_ ;
  assign \new_[76481]_  = \new_[76480]_  & \new_[76473]_ ;
  assign \new_[76485]_  = ~A266 & ~A234;
  assign \new_[76486]_  = ~A233 & \new_[76485]_ ;
  assign \new_[76489]_  = ~A269 & ~A268;
  assign \new_[76492]_  = ~A300 & A298;
  assign \new_[76493]_  = \new_[76492]_  & \new_[76489]_ ;
  assign \new_[76494]_  = \new_[76493]_  & \new_[76486]_ ;
  assign \new_[76498]_  = ~A167 & A169;
  assign \new_[76499]_  = ~A170 & \new_[76498]_ ;
  assign \new_[76502]_  = ~A200 & ~A166;
  assign \new_[76505]_  = ~A203 & ~A202;
  assign \new_[76506]_  = \new_[76505]_  & \new_[76502]_ ;
  assign \new_[76507]_  = \new_[76506]_  & \new_[76499]_ ;
  assign \new_[76511]_  = ~A266 & ~A234;
  assign \new_[76512]_  = ~A233 & \new_[76511]_ ;
  assign \new_[76515]_  = ~A269 & ~A268;
  assign \new_[76518]_  = A299 & A298;
  assign \new_[76519]_  = \new_[76518]_  & \new_[76515]_ ;
  assign \new_[76520]_  = \new_[76519]_  & \new_[76512]_ ;
  assign \new_[76524]_  = ~A167 & A169;
  assign \new_[76525]_  = ~A170 & \new_[76524]_ ;
  assign \new_[76528]_  = ~A200 & ~A166;
  assign \new_[76531]_  = ~A203 & ~A202;
  assign \new_[76532]_  = \new_[76531]_  & \new_[76528]_ ;
  assign \new_[76533]_  = \new_[76532]_  & \new_[76525]_ ;
  assign \new_[76537]_  = ~A266 & ~A234;
  assign \new_[76538]_  = ~A233 & \new_[76537]_ ;
  assign \new_[76541]_  = ~A269 & ~A268;
  assign \new_[76544]_  = ~A299 & ~A298;
  assign \new_[76545]_  = \new_[76544]_  & \new_[76541]_ ;
  assign \new_[76546]_  = \new_[76545]_  & \new_[76538]_ ;
  assign \new_[76550]_  = ~A167 & A169;
  assign \new_[76551]_  = ~A170 & \new_[76550]_ ;
  assign \new_[76554]_  = ~A200 & ~A166;
  assign \new_[76557]_  = ~A203 & ~A202;
  assign \new_[76558]_  = \new_[76557]_  & \new_[76554]_ ;
  assign \new_[76559]_  = \new_[76558]_  & \new_[76551]_ ;
  assign \new_[76563]_  = ~A266 & ~A234;
  assign \new_[76564]_  = ~A233 & \new_[76563]_ ;
  assign \new_[76567]_  = A298 & ~A267;
  assign \new_[76570]_  = ~A302 & ~A301;
  assign \new_[76571]_  = \new_[76570]_  & \new_[76567]_ ;
  assign \new_[76572]_  = \new_[76571]_  & \new_[76564]_ ;
  assign \new_[76576]_  = ~A167 & A169;
  assign \new_[76577]_  = ~A170 & \new_[76576]_ ;
  assign \new_[76580]_  = ~A200 & ~A166;
  assign \new_[76583]_  = ~A203 & ~A202;
  assign \new_[76584]_  = \new_[76583]_  & \new_[76580]_ ;
  assign \new_[76585]_  = \new_[76584]_  & \new_[76577]_ ;
  assign \new_[76589]_  = ~A265 & ~A234;
  assign \new_[76590]_  = ~A233 & \new_[76589]_ ;
  assign \new_[76593]_  = A298 & ~A266;
  assign \new_[76596]_  = ~A302 & ~A301;
  assign \new_[76597]_  = \new_[76596]_  & \new_[76593]_ ;
  assign \new_[76598]_  = \new_[76597]_  & \new_[76590]_ ;
  assign \new_[76602]_  = ~A167 & A169;
  assign \new_[76603]_  = ~A170 & \new_[76602]_ ;
  assign \new_[76606]_  = ~A200 & ~A166;
  assign \new_[76609]_  = ~A203 & ~A202;
  assign \new_[76610]_  = \new_[76609]_  & \new_[76606]_ ;
  assign \new_[76611]_  = \new_[76610]_  & \new_[76603]_ ;
  assign \new_[76615]_  = A265 & ~A233;
  assign \new_[76616]_  = ~A232 & \new_[76615]_ ;
  assign \new_[76619]_  = A298 & A266;
  assign \new_[76622]_  = ~A302 & ~A301;
  assign \new_[76623]_  = \new_[76622]_  & \new_[76619]_ ;
  assign \new_[76624]_  = \new_[76623]_  & \new_[76616]_ ;
  assign \new_[76628]_  = ~A167 & A169;
  assign \new_[76629]_  = ~A170 & \new_[76628]_ ;
  assign \new_[76632]_  = ~A200 & ~A166;
  assign \new_[76635]_  = ~A203 & ~A202;
  assign \new_[76636]_  = \new_[76635]_  & \new_[76632]_ ;
  assign \new_[76637]_  = \new_[76636]_  & \new_[76629]_ ;
  assign \new_[76641]_  = ~A266 & ~A233;
  assign \new_[76642]_  = ~A232 & \new_[76641]_ ;
  assign \new_[76645]_  = ~A269 & ~A268;
  assign \new_[76648]_  = ~A300 & A298;
  assign \new_[76649]_  = \new_[76648]_  & \new_[76645]_ ;
  assign \new_[76650]_  = \new_[76649]_  & \new_[76642]_ ;
  assign \new_[76654]_  = ~A167 & A169;
  assign \new_[76655]_  = ~A170 & \new_[76654]_ ;
  assign \new_[76658]_  = ~A200 & ~A166;
  assign \new_[76661]_  = ~A203 & ~A202;
  assign \new_[76662]_  = \new_[76661]_  & \new_[76658]_ ;
  assign \new_[76663]_  = \new_[76662]_  & \new_[76655]_ ;
  assign \new_[76667]_  = ~A266 & ~A233;
  assign \new_[76668]_  = ~A232 & \new_[76667]_ ;
  assign \new_[76671]_  = ~A269 & ~A268;
  assign \new_[76674]_  = A299 & A298;
  assign \new_[76675]_  = \new_[76674]_  & \new_[76671]_ ;
  assign \new_[76676]_  = \new_[76675]_  & \new_[76668]_ ;
  assign \new_[76680]_  = ~A167 & A169;
  assign \new_[76681]_  = ~A170 & \new_[76680]_ ;
  assign \new_[76684]_  = ~A200 & ~A166;
  assign \new_[76687]_  = ~A203 & ~A202;
  assign \new_[76688]_  = \new_[76687]_  & \new_[76684]_ ;
  assign \new_[76689]_  = \new_[76688]_  & \new_[76681]_ ;
  assign \new_[76693]_  = ~A266 & ~A233;
  assign \new_[76694]_  = ~A232 & \new_[76693]_ ;
  assign \new_[76697]_  = ~A269 & ~A268;
  assign \new_[76700]_  = ~A299 & ~A298;
  assign \new_[76701]_  = \new_[76700]_  & \new_[76697]_ ;
  assign \new_[76702]_  = \new_[76701]_  & \new_[76694]_ ;
  assign \new_[76706]_  = ~A167 & A169;
  assign \new_[76707]_  = ~A170 & \new_[76706]_ ;
  assign \new_[76710]_  = ~A200 & ~A166;
  assign \new_[76713]_  = ~A203 & ~A202;
  assign \new_[76714]_  = \new_[76713]_  & \new_[76710]_ ;
  assign \new_[76715]_  = \new_[76714]_  & \new_[76707]_ ;
  assign \new_[76719]_  = ~A266 & ~A233;
  assign \new_[76720]_  = ~A232 & \new_[76719]_ ;
  assign \new_[76723]_  = A298 & ~A267;
  assign \new_[76726]_  = ~A302 & ~A301;
  assign \new_[76727]_  = \new_[76726]_  & \new_[76723]_ ;
  assign \new_[76728]_  = \new_[76727]_  & \new_[76720]_ ;
  assign \new_[76732]_  = ~A167 & A169;
  assign \new_[76733]_  = ~A170 & \new_[76732]_ ;
  assign \new_[76736]_  = ~A200 & ~A166;
  assign \new_[76739]_  = ~A203 & ~A202;
  assign \new_[76740]_  = \new_[76739]_  & \new_[76736]_ ;
  assign \new_[76741]_  = \new_[76740]_  & \new_[76733]_ ;
  assign \new_[76745]_  = ~A265 & ~A233;
  assign \new_[76746]_  = ~A232 & \new_[76745]_ ;
  assign \new_[76749]_  = A298 & ~A266;
  assign \new_[76752]_  = ~A302 & ~A301;
  assign \new_[76753]_  = \new_[76752]_  & \new_[76749]_ ;
  assign \new_[76754]_  = \new_[76753]_  & \new_[76746]_ ;
  assign \new_[76758]_  = ~A167 & A169;
  assign \new_[76759]_  = ~A170 & \new_[76758]_ ;
  assign \new_[76762]_  = ~A200 & ~A166;
  assign \new_[76765]_  = A232 & ~A201;
  assign \new_[76766]_  = \new_[76765]_  & \new_[76762]_ ;
  assign \new_[76767]_  = \new_[76766]_  & \new_[76759]_ ;
  assign \new_[76771]_  = ~A268 & A265;
  assign \new_[76772]_  = A233 & \new_[76771]_ ;
  assign \new_[76775]_  = ~A299 & ~A269;
  assign \new_[76778]_  = ~A302 & ~A301;
  assign \new_[76779]_  = \new_[76778]_  & \new_[76775]_ ;
  assign \new_[76780]_  = \new_[76779]_  & \new_[76772]_ ;
  assign \new_[76784]_  = ~A167 & A169;
  assign \new_[76785]_  = ~A170 & \new_[76784]_ ;
  assign \new_[76788]_  = ~A200 & ~A166;
  assign \new_[76791]_  = ~A233 & ~A201;
  assign \new_[76792]_  = \new_[76791]_  & \new_[76788]_ ;
  assign \new_[76793]_  = \new_[76792]_  & \new_[76785]_ ;
  assign \new_[76797]_  = A265 & ~A236;
  assign \new_[76798]_  = ~A235 & \new_[76797]_ ;
  assign \new_[76801]_  = A298 & A266;
  assign \new_[76804]_  = ~A302 & ~A301;
  assign \new_[76805]_  = \new_[76804]_  & \new_[76801]_ ;
  assign \new_[76806]_  = \new_[76805]_  & \new_[76798]_ ;
  assign \new_[76810]_  = ~A167 & A169;
  assign \new_[76811]_  = ~A170 & \new_[76810]_ ;
  assign \new_[76814]_  = ~A200 & ~A166;
  assign \new_[76817]_  = ~A233 & ~A201;
  assign \new_[76818]_  = \new_[76817]_  & \new_[76814]_ ;
  assign \new_[76819]_  = \new_[76818]_  & \new_[76811]_ ;
  assign \new_[76823]_  = ~A266 & ~A236;
  assign \new_[76824]_  = ~A235 & \new_[76823]_ ;
  assign \new_[76827]_  = ~A269 & ~A268;
  assign \new_[76830]_  = ~A300 & A298;
  assign \new_[76831]_  = \new_[76830]_  & \new_[76827]_ ;
  assign \new_[76832]_  = \new_[76831]_  & \new_[76824]_ ;
  assign \new_[76836]_  = ~A167 & A169;
  assign \new_[76837]_  = ~A170 & \new_[76836]_ ;
  assign \new_[76840]_  = ~A200 & ~A166;
  assign \new_[76843]_  = ~A233 & ~A201;
  assign \new_[76844]_  = \new_[76843]_  & \new_[76840]_ ;
  assign \new_[76845]_  = \new_[76844]_  & \new_[76837]_ ;
  assign \new_[76849]_  = ~A266 & ~A236;
  assign \new_[76850]_  = ~A235 & \new_[76849]_ ;
  assign \new_[76853]_  = ~A269 & ~A268;
  assign \new_[76856]_  = A299 & A298;
  assign \new_[76857]_  = \new_[76856]_  & \new_[76853]_ ;
  assign \new_[76858]_  = \new_[76857]_  & \new_[76850]_ ;
  assign \new_[76862]_  = ~A167 & A169;
  assign \new_[76863]_  = ~A170 & \new_[76862]_ ;
  assign \new_[76866]_  = ~A200 & ~A166;
  assign \new_[76869]_  = ~A233 & ~A201;
  assign \new_[76870]_  = \new_[76869]_  & \new_[76866]_ ;
  assign \new_[76871]_  = \new_[76870]_  & \new_[76863]_ ;
  assign \new_[76875]_  = ~A266 & ~A236;
  assign \new_[76876]_  = ~A235 & \new_[76875]_ ;
  assign \new_[76879]_  = ~A269 & ~A268;
  assign \new_[76882]_  = ~A299 & ~A298;
  assign \new_[76883]_  = \new_[76882]_  & \new_[76879]_ ;
  assign \new_[76884]_  = \new_[76883]_  & \new_[76876]_ ;
  assign \new_[76888]_  = ~A167 & A169;
  assign \new_[76889]_  = ~A170 & \new_[76888]_ ;
  assign \new_[76892]_  = ~A200 & ~A166;
  assign \new_[76895]_  = ~A233 & ~A201;
  assign \new_[76896]_  = \new_[76895]_  & \new_[76892]_ ;
  assign \new_[76897]_  = \new_[76896]_  & \new_[76889]_ ;
  assign \new_[76901]_  = ~A266 & ~A236;
  assign \new_[76902]_  = ~A235 & \new_[76901]_ ;
  assign \new_[76905]_  = A298 & ~A267;
  assign \new_[76908]_  = ~A302 & ~A301;
  assign \new_[76909]_  = \new_[76908]_  & \new_[76905]_ ;
  assign \new_[76910]_  = \new_[76909]_  & \new_[76902]_ ;
  assign \new_[76914]_  = ~A167 & A169;
  assign \new_[76915]_  = ~A170 & \new_[76914]_ ;
  assign \new_[76918]_  = ~A200 & ~A166;
  assign \new_[76921]_  = ~A233 & ~A201;
  assign \new_[76922]_  = \new_[76921]_  & \new_[76918]_ ;
  assign \new_[76923]_  = \new_[76922]_  & \new_[76915]_ ;
  assign \new_[76927]_  = ~A265 & ~A236;
  assign \new_[76928]_  = ~A235 & \new_[76927]_ ;
  assign \new_[76931]_  = A298 & ~A266;
  assign \new_[76934]_  = ~A302 & ~A301;
  assign \new_[76935]_  = \new_[76934]_  & \new_[76931]_ ;
  assign \new_[76936]_  = \new_[76935]_  & \new_[76928]_ ;
  assign \new_[76940]_  = ~A167 & A169;
  assign \new_[76941]_  = ~A170 & \new_[76940]_ ;
  assign \new_[76944]_  = ~A200 & ~A166;
  assign \new_[76947]_  = ~A233 & ~A201;
  assign \new_[76948]_  = \new_[76947]_  & \new_[76944]_ ;
  assign \new_[76949]_  = \new_[76948]_  & \new_[76941]_ ;
  assign \new_[76953]_  = ~A268 & ~A266;
  assign \new_[76954]_  = ~A234 & \new_[76953]_ ;
  assign \new_[76957]_  = A298 & ~A269;
  assign \new_[76960]_  = ~A302 & ~A301;
  assign \new_[76961]_  = \new_[76960]_  & \new_[76957]_ ;
  assign \new_[76962]_  = \new_[76961]_  & \new_[76954]_ ;
  assign \new_[76966]_  = ~A167 & A169;
  assign \new_[76967]_  = ~A170 & \new_[76966]_ ;
  assign \new_[76970]_  = ~A200 & ~A166;
  assign \new_[76973]_  = A232 & ~A201;
  assign \new_[76974]_  = \new_[76973]_  & \new_[76970]_ ;
  assign \new_[76975]_  = \new_[76974]_  & \new_[76967]_ ;
  assign \new_[76979]_  = A235 & A234;
  assign \new_[76980]_  = ~A233 & \new_[76979]_ ;
  assign \new_[76983]_  = ~A299 & A298;
  assign \new_[76986]_  = A301 & A300;
  assign \new_[76987]_  = \new_[76986]_  & \new_[76983]_ ;
  assign \new_[76988]_  = \new_[76987]_  & \new_[76980]_ ;
  assign \new_[76992]_  = ~A167 & A169;
  assign \new_[76993]_  = ~A170 & \new_[76992]_ ;
  assign \new_[76996]_  = ~A200 & ~A166;
  assign \new_[76999]_  = A232 & ~A201;
  assign \new_[77000]_  = \new_[76999]_  & \new_[76996]_ ;
  assign \new_[77001]_  = \new_[77000]_  & \new_[76993]_ ;
  assign \new_[77005]_  = A235 & A234;
  assign \new_[77006]_  = ~A233 & \new_[77005]_ ;
  assign \new_[77009]_  = ~A299 & A298;
  assign \new_[77012]_  = A302 & A300;
  assign \new_[77013]_  = \new_[77012]_  & \new_[77009]_ ;
  assign \new_[77014]_  = \new_[77013]_  & \new_[77006]_ ;
  assign \new_[77018]_  = ~A167 & A169;
  assign \new_[77019]_  = ~A170 & \new_[77018]_ ;
  assign \new_[77022]_  = ~A200 & ~A166;
  assign \new_[77025]_  = A232 & ~A201;
  assign \new_[77026]_  = \new_[77025]_  & \new_[77022]_ ;
  assign \new_[77027]_  = \new_[77026]_  & \new_[77019]_ ;
  assign \new_[77031]_  = A235 & A234;
  assign \new_[77032]_  = ~A233 & \new_[77031]_ ;
  assign \new_[77035]_  = ~A266 & A265;
  assign \new_[77038]_  = A268 & A267;
  assign \new_[77039]_  = \new_[77038]_  & \new_[77035]_ ;
  assign \new_[77040]_  = \new_[77039]_  & \new_[77032]_ ;
  assign \new_[77044]_  = ~A167 & A169;
  assign \new_[77045]_  = ~A170 & \new_[77044]_ ;
  assign \new_[77048]_  = ~A200 & ~A166;
  assign \new_[77051]_  = A232 & ~A201;
  assign \new_[77052]_  = \new_[77051]_  & \new_[77048]_ ;
  assign \new_[77053]_  = \new_[77052]_  & \new_[77045]_ ;
  assign \new_[77057]_  = A235 & A234;
  assign \new_[77058]_  = ~A233 & \new_[77057]_ ;
  assign \new_[77061]_  = ~A266 & A265;
  assign \new_[77064]_  = A269 & A267;
  assign \new_[77065]_  = \new_[77064]_  & \new_[77061]_ ;
  assign \new_[77066]_  = \new_[77065]_  & \new_[77058]_ ;
  assign \new_[77070]_  = ~A167 & A169;
  assign \new_[77071]_  = ~A170 & \new_[77070]_ ;
  assign \new_[77074]_  = ~A200 & ~A166;
  assign \new_[77077]_  = A232 & ~A201;
  assign \new_[77078]_  = \new_[77077]_  & \new_[77074]_ ;
  assign \new_[77079]_  = \new_[77078]_  & \new_[77071]_ ;
  assign \new_[77083]_  = A236 & A234;
  assign \new_[77084]_  = ~A233 & \new_[77083]_ ;
  assign \new_[77087]_  = ~A299 & A298;
  assign \new_[77090]_  = A301 & A300;
  assign \new_[77091]_  = \new_[77090]_  & \new_[77087]_ ;
  assign \new_[77092]_  = \new_[77091]_  & \new_[77084]_ ;
  assign \new_[77096]_  = ~A167 & A169;
  assign \new_[77097]_  = ~A170 & \new_[77096]_ ;
  assign \new_[77100]_  = ~A200 & ~A166;
  assign \new_[77103]_  = A232 & ~A201;
  assign \new_[77104]_  = \new_[77103]_  & \new_[77100]_ ;
  assign \new_[77105]_  = \new_[77104]_  & \new_[77097]_ ;
  assign \new_[77109]_  = A236 & A234;
  assign \new_[77110]_  = ~A233 & \new_[77109]_ ;
  assign \new_[77113]_  = ~A299 & A298;
  assign \new_[77116]_  = A302 & A300;
  assign \new_[77117]_  = \new_[77116]_  & \new_[77113]_ ;
  assign \new_[77118]_  = \new_[77117]_  & \new_[77110]_ ;
  assign \new_[77122]_  = ~A167 & A169;
  assign \new_[77123]_  = ~A170 & \new_[77122]_ ;
  assign \new_[77126]_  = ~A200 & ~A166;
  assign \new_[77129]_  = A232 & ~A201;
  assign \new_[77130]_  = \new_[77129]_  & \new_[77126]_ ;
  assign \new_[77131]_  = \new_[77130]_  & \new_[77123]_ ;
  assign \new_[77135]_  = A236 & A234;
  assign \new_[77136]_  = ~A233 & \new_[77135]_ ;
  assign \new_[77139]_  = ~A266 & A265;
  assign \new_[77142]_  = A268 & A267;
  assign \new_[77143]_  = \new_[77142]_  & \new_[77139]_ ;
  assign \new_[77144]_  = \new_[77143]_  & \new_[77136]_ ;
  assign \new_[77148]_  = ~A167 & A169;
  assign \new_[77149]_  = ~A170 & \new_[77148]_ ;
  assign \new_[77152]_  = ~A200 & ~A166;
  assign \new_[77155]_  = A232 & ~A201;
  assign \new_[77156]_  = \new_[77155]_  & \new_[77152]_ ;
  assign \new_[77157]_  = \new_[77156]_  & \new_[77149]_ ;
  assign \new_[77161]_  = A236 & A234;
  assign \new_[77162]_  = ~A233 & \new_[77161]_ ;
  assign \new_[77165]_  = ~A266 & A265;
  assign \new_[77168]_  = A269 & A267;
  assign \new_[77169]_  = \new_[77168]_  & \new_[77165]_ ;
  assign \new_[77170]_  = \new_[77169]_  & \new_[77162]_ ;
  assign \new_[77174]_  = ~A167 & A169;
  assign \new_[77175]_  = ~A170 & \new_[77174]_ ;
  assign \new_[77178]_  = ~A200 & ~A166;
  assign \new_[77181]_  = ~A232 & ~A201;
  assign \new_[77182]_  = \new_[77181]_  & \new_[77178]_ ;
  assign \new_[77183]_  = \new_[77182]_  & \new_[77175]_ ;
  assign \new_[77187]_  = ~A268 & ~A266;
  assign \new_[77188]_  = ~A233 & \new_[77187]_ ;
  assign \new_[77191]_  = A298 & ~A269;
  assign \new_[77194]_  = ~A302 & ~A301;
  assign \new_[77195]_  = \new_[77194]_  & \new_[77191]_ ;
  assign \new_[77196]_  = \new_[77195]_  & \new_[77188]_ ;
  assign \new_[77200]_  = ~A167 & A169;
  assign \new_[77201]_  = ~A170 & \new_[77200]_ ;
  assign \new_[77204]_  = ~A199 & ~A166;
  assign \new_[77207]_  = A232 & ~A200;
  assign \new_[77208]_  = \new_[77207]_  & \new_[77204]_ ;
  assign \new_[77209]_  = \new_[77208]_  & \new_[77201]_ ;
  assign \new_[77213]_  = ~A268 & A265;
  assign \new_[77214]_  = A233 & \new_[77213]_ ;
  assign \new_[77217]_  = ~A299 & ~A269;
  assign \new_[77220]_  = ~A302 & ~A301;
  assign \new_[77221]_  = \new_[77220]_  & \new_[77217]_ ;
  assign \new_[77222]_  = \new_[77221]_  & \new_[77214]_ ;
  assign \new_[77226]_  = ~A167 & A169;
  assign \new_[77227]_  = ~A170 & \new_[77226]_ ;
  assign \new_[77230]_  = ~A199 & ~A166;
  assign \new_[77233]_  = ~A233 & ~A200;
  assign \new_[77234]_  = \new_[77233]_  & \new_[77230]_ ;
  assign \new_[77235]_  = \new_[77234]_  & \new_[77227]_ ;
  assign \new_[77239]_  = A265 & ~A236;
  assign \new_[77240]_  = ~A235 & \new_[77239]_ ;
  assign \new_[77243]_  = A298 & A266;
  assign \new_[77246]_  = ~A302 & ~A301;
  assign \new_[77247]_  = \new_[77246]_  & \new_[77243]_ ;
  assign \new_[77248]_  = \new_[77247]_  & \new_[77240]_ ;
  assign \new_[77252]_  = ~A167 & A169;
  assign \new_[77253]_  = ~A170 & \new_[77252]_ ;
  assign \new_[77256]_  = ~A199 & ~A166;
  assign \new_[77259]_  = ~A233 & ~A200;
  assign \new_[77260]_  = \new_[77259]_  & \new_[77256]_ ;
  assign \new_[77261]_  = \new_[77260]_  & \new_[77253]_ ;
  assign \new_[77265]_  = ~A266 & ~A236;
  assign \new_[77266]_  = ~A235 & \new_[77265]_ ;
  assign \new_[77269]_  = ~A269 & ~A268;
  assign \new_[77272]_  = ~A300 & A298;
  assign \new_[77273]_  = \new_[77272]_  & \new_[77269]_ ;
  assign \new_[77274]_  = \new_[77273]_  & \new_[77266]_ ;
  assign \new_[77278]_  = ~A167 & A169;
  assign \new_[77279]_  = ~A170 & \new_[77278]_ ;
  assign \new_[77282]_  = ~A199 & ~A166;
  assign \new_[77285]_  = ~A233 & ~A200;
  assign \new_[77286]_  = \new_[77285]_  & \new_[77282]_ ;
  assign \new_[77287]_  = \new_[77286]_  & \new_[77279]_ ;
  assign \new_[77291]_  = ~A266 & ~A236;
  assign \new_[77292]_  = ~A235 & \new_[77291]_ ;
  assign \new_[77295]_  = ~A269 & ~A268;
  assign \new_[77298]_  = A299 & A298;
  assign \new_[77299]_  = \new_[77298]_  & \new_[77295]_ ;
  assign \new_[77300]_  = \new_[77299]_  & \new_[77292]_ ;
  assign \new_[77304]_  = ~A167 & A169;
  assign \new_[77305]_  = ~A170 & \new_[77304]_ ;
  assign \new_[77308]_  = ~A199 & ~A166;
  assign \new_[77311]_  = ~A233 & ~A200;
  assign \new_[77312]_  = \new_[77311]_  & \new_[77308]_ ;
  assign \new_[77313]_  = \new_[77312]_  & \new_[77305]_ ;
  assign \new_[77317]_  = ~A266 & ~A236;
  assign \new_[77318]_  = ~A235 & \new_[77317]_ ;
  assign \new_[77321]_  = ~A269 & ~A268;
  assign \new_[77324]_  = ~A299 & ~A298;
  assign \new_[77325]_  = \new_[77324]_  & \new_[77321]_ ;
  assign \new_[77326]_  = \new_[77325]_  & \new_[77318]_ ;
  assign \new_[77330]_  = ~A167 & A169;
  assign \new_[77331]_  = ~A170 & \new_[77330]_ ;
  assign \new_[77334]_  = ~A199 & ~A166;
  assign \new_[77337]_  = ~A233 & ~A200;
  assign \new_[77338]_  = \new_[77337]_  & \new_[77334]_ ;
  assign \new_[77339]_  = \new_[77338]_  & \new_[77331]_ ;
  assign \new_[77343]_  = ~A266 & ~A236;
  assign \new_[77344]_  = ~A235 & \new_[77343]_ ;
  assign \new_[77347]_  = A298 & ~A267;
  assign \new_[77350]_  = ~A302 & ~A301;
  assign \new_[77351]_  = \new_[77350]_  & \new_[77347]_ ;
  assign \new_[77352]_  = \new_[77351]_  & \new_[77344]_ ;
  assign \new_[77356]_  = ~A167 & A169;
  assign \new_[77357]_  = ~A170 & \new_[77356]_ ;
  assign \new_[77360]_  = ~A199 & ~A166;
  assign \new_[77363]_  = ~A233 & ~A200;
  assign \new_[77364]_  = \new_[77363]_  & \new_[77360]_ ;
  assign \new_[77365]_  = \new_[77364]_  & \new_[77357]_ ;
  assign \new_[77369]_  = ~A265 & ~A236;
  assign \new_[77370]_  = ~A235 & \new_[77369]_ ;
  assign \new_[77373]_  = A298 & ~A266;
  assign \new_[77376]_  = ~A302 & ~A301;
  assign \new_[77377]_  = \new_[77376]_  & \new_[77373]_ ;
  assign \new_[77378]_  = \new_[77377]_  & \new_[77370]_ ;
  assign \new_[77382]_  = ~A167 & A169;
  assign \new_[77383]_  = ~A170 & \new_[77382]_ ;
  assign \new_[77386]_  = ~A199 & ~A166;
  assign \new_[77389]_  = ~A233 & ~A200;
  assign \new_[77390]_  = \new_[77389]_  & \new_[77386]_ ;
  assign \new_[77391]_  = \new_[77390]_  & \new_[77383]_ ;
  assign \new_[77395]_  = ~A268 & ~A266;
  assign \new_[77396]_  = ~A234 & \new_[77395]_ ;
  assign \new_[77399]_  = A298 & ~A269;
  assign \new_[77402]_  = ~A302 & ~A301;
  assign \new_[77403]_  = \new_[77402]_  & \new_[77399]_ ;
  assign \new_[77404]_  = \new_[77403]_  & \new_[77396]_ ;
  assign \new_[77408]_  = ~A167 & A169;
  assign \new_[77409]_  = ~A170 & \new_[77408]_ ;
  assign \new_[77412]_  = ~A199 & ~A166;
  assign \new_[77415]_  = A232 & ~A200;
  assign \new_[77416]_  = \new_[77415]_  & \new_[77412]_ ;
  assign \new_[77417]_  = \new_[77416]_  & \new_[77409]_ ;
  assign \new_[77421]_  = A235 & A234;
  assign \new_[77422]_  = ~A233 & \new_[77421]_ ;
  assign \new_[77425]_  = ~A299 & A298;
  assign \new_[77428]_  = A301 & A300;
  assign \new_[77429]_  = \new_[77428]_  & \new_[77425]_ ;
  assign \new_[77430]_  = \new_[77429]_  & \new_[77422]_ ;
  assign \new_[77434]_  = ~A167 & A169;
  assign \new_[77435]_  = ~A170 & \new_[77434]_ ;
  assign \new_[77438]_  = ~A199 & ~A166;
  assign \new_[77441]_  = A232 & ~A200;
  assign \new_[77442]_  = \new_[77441]_  & \new_[77438]_ ;
  assign \new_[77443]_  = \new_[77442]_  & \new_[77435]_ ;
  assign \new_[77447]_  = A235 & A234;
  assign \new_[77448]_  = ~A233 & \new_[77447]_ ;
  assign \new_[77451]_  = ~A299 & A298;
  assign \new_[77454]_  = A302 & A300;
  assign \new_[77455]_  = \new_[77454]_  & \new_[77451]_ ;
  assign \new_[77456]_  = \new_[77455]_  & \new_[77448]_ ;
  assign \new_[77460]_  = ~A167 & A169;
  assign \new_[77461]_  = ~A170 & \new_[77460]_ ;
  assign \new_[77464]_  = ~A199 & ~A166;
  assign \new_[77467]_  = A232 & ~A200;
  assign \new_[77468]_  = \new_[77467]_  & \new_[77464]_ ;
  assign \new_[77469]_  = \new_[77468]_  & \new_[77461]_ ;
  assign \new_[77473]_  = A235 & A234;
  assign \new_[77474]_  = ~A233 & \new_[77473]_ ;
  assign \new_[77477]_  = ~A266 & A265;
  assign \new_[77480]_  = A268 & A267;
  assign \new_[77481]_  = \new_[77480]_  & \new_[77477]_ ;
  assign \new_[77482]_  = \new_[77481]_  & \new_[77474]_ ;
  assign \new_[77486]_  = ~A167 & A169;
  assign \new_[77487]_  = ~A170 & \new_[77486]_ ;
  assign \new_[77490]_  = ~A199 & ~A166;
  assign \new_[77493]_  = A232 & ~A200;
  assign \new_[77494]_  = \new_[77493]_  & \new_[77490]_ ;
  assign \new_[77495]_  = \new_[77494]_  & \new_[77487]_ ;
  assign \new_[77499]_  = A235 & A234;
  assign \new_[77500]_  = ~A233 & \new_[77499]_ ;
  assign \new_[77503]_  = ~A266 & A265;
  assign \new_[77506]_  = A269 & A267;
  assign \new_[77507]_  = \new_[77506]_  & \new_[77503]_ ;
  assign \new_[77508]_  = \new_[77507]_  & \new_[77500]_ ;
  assign \new_[77512]_  = ~A167 & A169;
  assign \new_[77513]_  = ~A170 & \new_[77512]_ ;
  assign \new_[77516]_  = ~A199 & ~A166;
  assign \new_[77519]_  = A232 & ~A200;
  assign \new_[77520]_  = \new_[77519]_  & \new_[77516]_ ;
  assign \new_[77521]_  = \new_[77520]_  & \new_[77513]_ ;
  assign \new_[77525]_  = A236 & A234;
  assign \new_[77526]_  = ~A233 & \new_[77525]_ ;
  assign \new_[77529]_  = ~A299 & A298;
  assign \new_[77532]_  = A301 & A300;
  assign \new_[77533]_  = \new_[77532]_  & \new_[77529]_ ;
  assign \new_[77534]_  = \new_[77533]_  & \new_[77526]_ ;
  assign \new_[77538]_  = ~A167 & A169;
  assign \new_[77539]_  = ~A170 & \new_[77538]_ ;
  assign \new_[77542]_  = ~A199 & ~A166;
  assign \new_[77545]_  = A232 & ~A200;
  assign \new_[77546]_  = \new_[77545]_  & \new_[77542]_ ;
  assign \new_[77547]_  = \new_[77546]_  & \new_[77539]_ ;
  assign \new_[77551]_  = A236 & A234;
  assign \new_[77552]_  = ~A233 & \new_[77551]_ ;
  assign \new_[77555]_  = ~A299 & A298;
  assign \new_[77558]_  = A302 & A300;
  assign \new_[77559]_  = \new_[77558]_  & \new_[77555]_ ;
  assign \new_[77560]_  = \new_[77559]_  & \new_[77552]_ ;
  assign \new_[77564]_  = ~A167 & A169;
  assign \new_[77565]_  = ~A170 & \new_[77564]_ ;
  assign \new_[77568]_  = ~A199 & ~A166;
  assign \new_[77571]_  = A232 & ~A200;
  assign \new_[77572]_  = \new_[77571]_  & \new_[77568]_ ;
  assign \new_[77573]_  = \new_[77572]_  & \new_[77565]_ ;
  assign \new_[77577]_  = A236 & A234;
  assign \new_[77578]_  = ~A233 & \new_[77577]_ ;
  assign \new_[77581]_  = ~A266 & A265;
  assign \new_[77584]_  = A268 & A267;
  assign \new_[77585]_  = \new_[77584]_  & \new_[77581]_ ;
  assign \new_[77586]_  = \new_[77585]_  & \new_[77578]_ ;
  assign \new_[77590]_  = ~A167 & A169;
  assign \new_[77591]_  = ~A170 & \new_[77590]_ ;
  assign \new_[77594]_  = ~A199 & ~A166;
  assign \new_[77597]_  = A232 & ~A200;
  assign \new_[77598]_  = \new_[77597]_  & \new_[77594]_ ;
  assign \new_[77599]_  = \new_[77598]_  & \new_[77591]_ ;
  assign \new_[77603]_  = A236 & A234;
  assign \new_[77604]_  = ~A233 & \new_[77603]_ ;
  assign \new_[77607]_  = ~A266 & A265;
  assign \new_[77610]_  = A269 & A267;
  assign \new_[77611]_  = \new_[77610]_  & \new_[77607]_ ;
  assign \new_[77612]_  = \new_[77611]_  & \new_[77604]_ ;
  assign \new_[77616]_  = ~A167 & A169;
  assign \new_[77617]_  = ~A170 & \new_[77616]_ ;
  assign \new_[77620]_  = ~A199 & ~A166;
  assign \new_[77623]_  = ~A232 & ~A200;
  assign \new_[77624]_  = \new_[77623]_  & \new_[77620]_ ;
  assign \new_[77625]_  = \new_[77624]_  & \new_[77617]_ ;
  assign \new_[77629]_  = ~A268 & ~A266;
  assign \new_[77630]_  = ~A233 & \new_[77629]_ ;
  assign \new_[77633]_  = A298 & ~A269;
  assign \new_[77636]_  = ~A302 & ~A301;
  assign \new_[77637]_  = \new_[77636]_  & \new_[77633]_ ;
  assign \new_[77638]_  = \new_[77637]_  & \new_[77630]_ ;
  assign \new_[77642]_  = ~A166 & ~A167;
  assign \new_[77643]_  = ~A169 & \new_[77642]_ ;
  assign \new_[77646]_  = A200 & ~A199;
  assign \new_[77649]_  = ~A235 & ~A233;
  assign \new_[77650]_  = \new_[77649]_  & \new_[77646]_ ;
  assign \new_[77651]_  = \new_[77650]_  & \new_[77643]_ ;
  assign \new_[77655]_  = ~A268 & ~A266;
  assign \new_[77656]_  = ~A236 & \new_[77655]_ ;
  assign \new_[77659]_  = A298 & ~A269;
  assign \new_[77662]_  = ~A302 & ~A301;
  assign \new_[77663]_  = \new_[77662]_  & \new_[77659]_ ;
  assign \new_[77664]_  = \new_[77663]_  & \new_[77656]_ ;
  assign \new_[77668]_  = ~A166 & ~A167;
  assign \new_[77669]_  = ~A169 & \new_[77668]_ ;
  assign \new_[77672]_  = ~A200 & A199;
  assign \new_[77675]_  = A202 & A201;
  assign \new_[77676]_  = \new_[77675]_  & \new_[77672]_ ;
  assign \new_[77677]_  = \new_[77676]_  & \new_[77669]_ ;
  assign \new_[77681]_  = A265 & A233;
  assign \new_[77682]_  = A232 & \new_[77681]_ ;
  assign \new_[77685]_  = ~A269 & ~A268;
  assign \new_[77688]_  = ~A300 & ~A299;
  assign \new_[77689]_  = \new_[77688]_  & \new_[77685]_ ;
  assign \new_[77690]_  = \new_[77689]_  & \new_[77682]_ ;
  assign \new_[77694]_  = ~A166 & ~A167;
  assign \new_[77695]_  = ~A169 & \new_[77694]_ ;
  assign \new_[77698]_  = ~A200 & A199;
  assign \new_[77701]_  = A202 & A201;
  assign \new_[77702]_  = \new_[77701]_  & \new_[77698]_ ;
  assign \new_[77703]_  = \new_[77702]_  & \new_[77695]_ ;
  assign \new_[77707]_  = A265 & A233;
  assign \new_[77708]_  = A232 & \new_[77707]_ ;
  assign \new_[77711]_  = ~A269 & ~A268;
  assign \new_[77714]_  = A299 & A298;
  assign \new_[77715]_  = \new_[77714]_  & \new_[77711]_ ;
  assign \new_[77716]_  = \new_[77715]_  & \new_[77708]_ ;
  assign \new_[77720]_  = ~A166 & ~A167;
  assign \new_[77721]_  = ~A169 & \new_[77720]_ ;
  assign \new_[77724]_  = ~A200 & A199;
  assign \new_[77727]_  = A202 & A201;
  assign \new_[77728]_  = \new_[77727]_  & \new_[77724]_ ;
  assign \new_[77729]_  = \new_[77728]_  & \new_[77721]_ ;
  assign \new_[77733]_  = A265 & A233;
  assign \new_[77734]_  = A232 & \new_[77733]_ ;
  assign \new_[77737]_  = ~A269 & ~A268;
  assign \new_[77740]_  = ~A299 & ~A298;
  assign \new_[77741]_  = \new_[77740]_  & \new_[77737]_ ;
  assign \new_[77742]_  = \new_[77741]_  & \new_[77734]_ ;
  assign \new_[77746]_  = ~A166 & ~A167;
  assign \new_[77747]_  = ~A169 & \new_[77746]_ ;
  assign \new_[77750]_  = ~A200 & A199;
  assign \new_[77753]_  = A202 & A201;
  assign \new_[77754]_  = \new_[77753]_  & \new_[77750]_ ;
  assign \new_[77755]_  = \new_[77754]_  & \new_[77747]_ ;
  assign \new_[77759]_  = A265 & A233;
  assign \new_[77760]_  = A232 & \new_[77759]_ ;
  assign \new_[77763]_  = ~A299 & ~A267;
  assign \new_[77766]_  = ~A302 & ~A301;
  assign \new_[77767]_  = \new_[77766]_  & \new_[77763]_ ;
  assign \new_[77768]_  = \new_[77767]_  & \new_[77760]_ ;
  assign \new_[77772]_  = ~A166 & ~A167;
  assign \new_[77773]_  = ~A169 & \new_[77772]_ ;
  assign \new_[77776]_  = ~A200 & A199;
  assign \new_[77779]_  = A202 & A201;
  assign \new_[77780]_  = \new_[77779]_  & \new_[77776]_ ;
  assign \new_[77781]_  = \new_[77780]_  & \new_[77773]_ ;
  assign \new_[77785]_  = A265 & A233;
  assign \new_[77786]_  = A232 & \new_[77785]_ ;
  assign \new_[77789]_  = ~A299 & A266;
  assign \new_[77792]_  = ~A302 & ~A301;
  assign \new_[77793]_  = \new_[77792]_  & \new_[77789]_ ;
  assign \new_[77794]_  = \new_[77793]_  & \new_[77786]_ ;
  assign \new_[77798]_  = ~A166 & ~A167;
  assign \new_[77799]_  = ~A169 & \new_[77798]_ ;
  assign \new_[77802]_  = ~A200 & A199;
  assign \new_[77805]_  = A202 & A201;
  assign \new_[77806]_  = \new_[77805]_  & \new_[77802]_ ;
  assign \new_[77807]_  = \new_[77806]_  & \new_[77799]_ ;
  assign \new_[77811]_  = ~A265 & A233;
  assign \new_[77812]_  = A232 & \new_[77811]_ ;
  assign \new_[77815]_  = ~A299 & ~A266;
  assign \new_[77818]_  = ~A302 & ~A301;
  assign \new_[77819]_  = \new_[77818]_  & \new_[77815]_ ;
  assign \new_[77820]_  = \new_[77819]_  & \new_[77812]_ ;
  assign \new_[77824]_  = ~A166 & ~A167;
  assign \new_[77825]_  = ~A169 & \new_[77824]_ ;
  assign \new_[77828]_  = ~A200 & A199;
  assign \new_[77831]_  = A202 & A201;
  assign \new_[77832]_  = \new_[77831]_  & \new_[77828]_ ;
  assign \new_[77833]_  = \new_[77832]_  & \new_[77825]_ ;
  assign \new_[77837]_  = ~A236 & ~A235;
  assign \new_[77838]_  = ~A233 & \new_[77837]_ ;
  assign \new_[77841]_  = A266 & A265;
  assign \new_[77844]_  = ~A300 & A298;
  assign \new_[77845]_  = \new_[77844]_  & \new_[77841]_ ;
  assign \new_[77846]_  = \new_[77845]_  & \new_[77838]_ ;
  assign \new_[77850]_  = ~A166 & ~A167;
  assign \new_[77851]_  = ~A169 & \new_[77850]_ ;
  assign \new_[77854]_  = ~A200 & A199;
  assign \new_[77857]_  = A202 & A201;
  assign \new_[77858]_  = \new_[77857]_  & \new_[77854]_ ;
  assign \new_[77859]_  = \new_[77858]_  & \new_[77851]_ ;
  assign \new_[77863]_  = ~A236 & ~A235;
  assign \new_[77864]_  = ~A233 & \new_[77863]_ ;
  assign \new_[77867]_  = A266 & A265;
  assign \new_[77870]_  = A299 & A298;
  assign \new_[77871]_  = \new_[77870]_  & \new_[77867]_ ;
  assign \new_[77872]_  = \new_[77871]_  & \new_[77864]_ ;
  assign \new_[77876]_  = ~A166 & ~A167;
  assign \new_[77877]_  = ~A169 & \new_[77876]_ ;
  assign \new_[77880]_  = ~A200 & A199;
  assign \new_[77883]_  = A202 & A201;
  assign \new_[77884]_  = \new_[77883]_  & \new_[77880]_ ;
  assign \new_[77885]_  = \new_[77884]_  & \new_[77877]_ ;
  assign \new_[77889]_  = ~A236 & ~A235;
  assign \new_[77890]_  = ~A233 & \new_[77889]_ ;
  assign \new_[77893]_  = A266 & A265;
  assign \new_[77896]_  = ~A299 & ~A298;
  assign \new_[77897]_  = \new_[77896]_  & \new_[77893]_ ;
  assign \new_[77898]_  = \new_[77897]_  & \new_[77890]_ ;
  assign \new_[77902]_  = ~A166 & ~A167;
  assign \new_[77903]_  = ~A169 & \new_[77902]_ ;
  assign \new_[77906]_  = ~A200 & A199;
  assign \new_[77909]_  = A202 & A201;
  assign \new_[77910]_  = \new_[77909]_  & \new_[77906]_ ;
  assign \new_[77911]_  = \new_[77910]_  & \new_[77903]_ ;
  assign \new_[77915]_  = ~A236 & ~A235;
  assign \new_[77916]_  = ~A233 & \new_[77915]_ ;
  assign \new_[77919]_  = ~A267 & ~A266;
  assign \new_[77922]_  = ~A300 & A298;
  assign \new_[77923]_  = \new_[77922]_  & \new_[77919]_ ;
  assign \new_[77924]_  = \new_[77923]_  & \new_[77916]_ ;
  assign \new_[77928]_  = ~A166 & ~A167;
  assign \new_[77929]_  = ~A169 & \new_[77928]_ ;
  assign \new_[77932]_  = ~A200 & A199;
  assign \new_[77935]_  = A202 & A201;
  assign \new_[77936]_  = \new_[77935]_  & \new_[77932]_ ;
  assign \new_[77937]_  = \new_[77936]_  & \new_[77929]_ ;
  assign \new_[77941]_  = ~A236 & ~A235;
  assign \new_[77942]_  = ~A233 & \new_[77941]_ ;
  assign \new_[77945]_  = ~A267 & ~A266;
  assign \new_[77948]_  = A299 & A298;
  assign \new_[77949]_  = \new_[77948]_  & \new_[77945]_ ;
  assign \new_[77950]_  = \new_[77949]_  & \new_[77942]_ ;
  assign \new_[77954]_  = ~A166 & ~A167;
  assign \new_[77955]_  = ~A169 & \new_[77954]_ ;
  assign \new_[77958]_  = ~A200 & A199;
  assign \new_[77961]_  = A202 & A201;
  assign \new_[77962]_  = \new_[77961]_  & \new_[77958]_ ;
  assign \new_[77963]_  = \new_[77962]_  & \new_[77955]_ ;
  assign \new_[77967]_  = ~A236 & ~A235;
  assign \new_[77968]_  = ~A233 & \new_[77967]_ ;
  assign \new_[77971]_  = ~A267 & ~A266;
  assign \new_[77974]_  = ~A299 & ~A298;
  assign \new_[77975]_  = \new_[77974]_  & \new_[77971]_ ;
  assign \new_[77976]_  = \new_[77975]_  & \new_[77968]_ ;
  assign \new_[77980]_  = ~A166 & ~A167;
  assign \new_[77981]_  = ~A169 & \new_[77980]_ ;
  assign \new_[77984]_  = ~A200 & A199;
  assign \new_[77987]_  = A202 & A201;
  assign \new_[77988]_  = \new_[77987]_  & \new_[77984]_ ;
  assign \new_[77989]_  = \new_[77988]_  & \new_[77981]_ ;
  assign \new_[77993]_  = ~A236 & ~A235;
  assign \new_[77994]_  = ~A233 & \new_[77993]_ ;
  assign \new_[77997]_  = ~A266 & ~A265;
  assign \new_[78000]_  = ~A300 & A298;
  assign \new_[78001]_  = \new_[78000]_  & \new_[77997]_ ;
  assign \new_[78002]_  = \new_[78001]_  & \new_[77994]_ ;
  assign \new_[78006]_  = ~A166 & ~A167;
  assign \new_[78007]_  = ~A169 & \new_[78006]_ ;
  assign \new_[78010]_  = ~A200 & A199;
  assign \new_[78013]_  = A202 & A201;
  assign \new_[78014]_  = \new_[78013]_  & \new_[78010]_ ;
  assign \new_[78015]_  = \new_[78014]_  & \new_[78007]_ ;
  assign \new_[78019]_  = ~A236 & ~A235;
  assign \new_[78020]_  = ~A233 & \new_[78019]_ ;
  assign \new_[78023]_  = ~A266 & ~A265;
  assign \new_[78026]_  = A299 & A298;
  assign \new_[78027]_  = \new_[78026]_  & \new_[78023]_ ;
  assign \new_[78028]_  = \new_[78027]_  & \new_[78020]_ ;
  assign \new_[78032]_  = ~A166 & ~A167;
  assign \new_[78033]_  = ~A169 & \new_[78032]_ ;
  assign \new_[78036]_  = ~A200 & A199;
  assign \new_[78039]_  = A202 & A201;
  assign \new_[78040]_  = \new_[78039]_  & \new_[78036]_ ;
  assign \new_[78041]_  = \new_[78040]_  & \new_[78033]_ ;
  assign \new_[78045]_  = ~A236 & ~A235;
  assign \new_[78046]_  = ~A233 & \new_[78045]_ ;
  assign \new_[78049]_  = ~A266 & ~A265;
  assign \new_[78052]_  = ~A299 & ~A298;
  assign \new_[78053]_  = \new_[78052]_  & \new_[78049]_ ;
  assign \new_[78054]_  = \new_[78053]_  & \new_[78046]_ ;
  assign \new_[78058]_  = ~A166 & ~A167;
  assign \new_[78059]_  = ~A169 & \new_[78058]_ ;
  assign \new_[78062]_  = ~A200 & A199;
  assign \new_[78065]_  = A202 & A201;
  assign \new_[78066]_  = \new_[78065]_  & \new_[78062]_ ;
  assign \new_[78067]_  = \new_[78066]_  & \new_[78059]_ ;
  assign \new_[78071]_  = A265 & ~A234;
  assign \new_[78072]_  = ~A233 & \new_[78071]_ ;
  assign \new_[78075]_  = A298 & A266;
  assign \new_[78078]_  = ~A302 & ~A301;
  assign \new_[78079]_  = \new_[78078]_  & \new_[78075]_ ;
  assign \new_[78080]_  = \new_[78079]_  & \new_[78072]_ ;
  assign \new_[78084]_  = ~A166 & ~A167;
  assign \new_[78085]_  = ~A169 & \new_[78084]_ ;
  assign \new_[78088]_  = ~A200 & A199;
  assign \new_[78091]_  = A202 & A201;
  assign \new_[78092]_  = \new_[78091]_  & \new_[78088]_ ;
  assign \new_[78093]_  = \new_[78092]_  & \new_[78085]_ ;
  assign \new_[78097]_  = ~A266 & ~A234;
  assign \new_[78098]_  = ~A233 & \new_[78097]_ ;
  assign \new_[78101]_  = ~A269 & ~A268;
  assign \new_[78104]_  = ~A300 & A298;
  assign \new_[78105]_  = \new_[78104]_  & \new_[78101]_ ;
  assign \new_[78106]_  = \new_[78105]_  & \new_[78098]_ ;
  assign \new_[78110]_  = ~A166 & ~A167;
  assign \new_[78111]_  = ~A169 & \new_[78110]_ ;
  assign \new_[78114]_  = ~A200 & A199;
  assign \new_[78117]_  = A202 & A201;
  assign \new_[78118]_  = \new_[78117]_  & \new_[78114]_ ;
  assign \new_[78119]_  = \new_[78118]_  & \new_[78111]_ ;
  assign \new_[78123]_  = ~A266 & ~A234;
  assign \new_[78124]_  = ~A233 & \new_[78123]_ ;
  assign \new_[78127]_  = ~A269 & ~A268;
  assign \new_[78130]_  = A299 & A298;
  assign \new_[78131]_  = \new_[78130]_  & \new_[78127]_ ;
  assign \new_[78132]_  = \new_[78131]_  & \new_[78124]_ ;
  assign \new_[78136]_  = ~A166 & ~A167;
  assign \new_[78137]_  = ~A169 & \new_[78136]_ ;
  assign \new_[78140]_  = ~A200 & A199;
  assign \new_[78143]_  = A202 & A201;
  assign \new_[78144]_  = \new_[78143]_  & \new_[78140]_ ;
  assign \new_[78145]_  = \new_[78144]_  & \new_[78137]_ ;
  assign \new_[78149]_  = ~A266 & ~A234;
  assign \new_[78150]_  = ~A233 & \new_[78149]_ ;
  assign \new_[78153]_  = ~A269 & ~A268;
  assign \new_[78156]_  = ~A299 & ~A298;
  assign \new_[78157]_  = \new_[78156]_  & \new_[78153]_ ;
  assign \new_[78158]_  = \new_[78157]_  & \new_[78150]_ ;
  assign \new_[78162]_  = ~A166 & ~A167;
  assign \new_[78163]_  = ~A169 & \new_[78162]_ ;
  assign \new_[78166]_  = ~A200 & A199;
  assign \new_[78169]_  = A202 & A201;
  assign \new_[78170]_  = \new_[78169]_  & \new_[78166]_ ;
  assign \new_[78171]_  = \new_[78170]_  & \new_[78163]_ ;
  assign \new_[78175]_  = ~A266 & ~A234;
  assign \new_[78176]_  = ~A233 & \new_[78175]_ ;
  assign \new_[78179]_  = A298 & ~A267;
  assign \new_[78182]_  = ~A302 & ~A301;
  assign \new_[78183]_  = \new_[78182]_  & \new_[78179]_ ;
  assign \new_[78184]_  = \new_[78183]_  & \new_[78176]_ ;
  assign \new_[78188]_  = ~A166 & ~A167;
  assign \new_[78189]_  = ~A169 & \new_[78188]_ ;
  assign \new_[78192]_  = ~A200 & A199;
  assign \new_[78195]_  = A202 & A201;
  assign \new_[78196]_  = \new_[78195]_  & \new_[78192]_ ;
  assign \new_[78197]_  = \new_[78196]_  & \new_[78189]_ ;
  assign \new_[78201]_  = ~A265 & ~A234;
  assign \new_[78202]_  = ~A233 & \new_[78201]_ ;
  assign \new_[78205]_  = A298 & ~A266;
  assign \new_[78208]_  = ~A302 & ~A301;
  assign \new_[78209]_  = \new_[78208]_  & \new_[78205]_ ;
  assign \new_[78210]_  = \new_[78209]_  & \new_[78202]_ ;
  assign \new_[78214]_  = ~A166 & ~A167;
  assign \new_[78215]_  = ~A169 & \new_[78214]_ ;
  assign \new_[78218]_  = ~A200 & A199;
  assign \new_[78221]_  = A202 & A201;
  assign \new_[78222]_  = \new_[78221]_  & \new_[78218]_ ;
  assign \new_[78223]_  = \new_[78222]_  & \new_[78215]_ ;
  assign \new_[78227]_  = A265 & ~A233;
  assign \new_[78228]_  = ~A232 & \new_[78227]_ ;
  assign \new_[78231]_  = A298 & A266;
  assign \new_[78234]_  = ~A302 & ~A301;
  assign \new_[78235]_  = \new_[78234]_  & \new_[78231]_ ;
  assign \new_[78236]_  = \new_[78235]_  & \new_[78228]_ ;
  assign \new_[78240]_  = ~A166 & ~A167;
  assign \new_[78241]_  = ~A169 & \new_[78240]_ ;
  assign \new_[78244]_  = ~A200 & A199;
  assign \new_[78247]_  = A202 & A201;
  assign \new_[78248]_  = \new_[78247]_  & \new_[78244]_ ;
  assign \new_[78249]_  = \new_[78248]_  & \new_[78241]_ ;
  assign \new_[78253]_  = ~A266 & ~A233;
  assign \new_[78254]_  = ~A232 & \new_[78253]_ ;
  assign \new_[78257]_  = ~A269 & ~A268;
  assign \new_[78260]_  = ~A300 & A298;
  assign \new_[78261]_  = \new_[78260]_  & \new_[78257]_ ;
  assign \new_[78262]_  = \new_[78261]_  & \new_[78254]_ ;
  assign \new_[78266]_  = ~A166 & ~A167;
  assign \new_[78267]_  = ~A169 & \new_[78266]_ ;
  assign \new_[78270]_  = ~A200 & A199;
  assign \new_[78273]_  = A202 & A201;
  assign \new_[78274]_  = \new_[78273]_  & \new_[78270]_ ;
  assign \new_[78275]_  = \new_[78274]_  & \new_[78267]_ ;
  assign \new_[78279]_  = ~A266 & ~A233;
  assign \new_[78280]_  = ~A232 & \new_[78279]_ ;
  assign \new_[78283]_  = ~A269 & ~A268;
  assign \new_[78286]_  = A299 & A298;
  assign \new_[78287]_  = \new_[78286]_  & \new_[78283]_ ;
  assign \new_[78288]_  = \new_[78287]_  & \new_[78280]_ ;
  assign \new_[78292]_  = ~A166 & ~A167;
  assign \new_[78293]_  = ~A169 & \new_[78292]_ ;
  assign \new_[78296]_  = ~A200 & A199;
  assign \new_[78299]_  = A202 & A201;
  assign \new_[78300]_  = \new_[78299]_  & \new_[78296]_ ;
  assign \new_[78301]_  = \new_[78300]_  & \new_[78293]_ ;
  assign \new_[78305]_  = ~A266 & ~A233;
  assign \new_[78306]_  = ~A232 & \new_[78305]_ ;
  assign \new_[78309]_  = ~A269 & ~A268;
  assign \new_[78312]_  = ~A299 & ~A298;
  assign \new_[78313]_  = \new_[78312]_  & \new_[78309]_ ;
  assign \new_[78314]_  = \new_[78313]_  & \new_[78306]_ ;
  assign \new_[78318]_  = ~A166 & ~A167;
  assign \new_[78319]_  = ~A169 & \new_[78318]_ ;
  assign \new_[78322]_  = ~A200 & A199;
  assign \new_[78325]_  = A202 & A201;
  assign \new_[78326]_  = \new_[78325]_  & \new_[78322]_ ;
  assign \new_[78327]_  = \new_[78326]_  & \new_[78319]_ ;
  assign \new_[78331]_  = ~A266 & ~A233;
  assign \new_[78332]_  = ~A232 & \new_[78331]_ ;
  assign \new_[78335]_  = A298 & ~A267;
  assign \new_[78338]_  = ~A302 & ~A301;
  assign \new_[78339]_  = \new_[78338]_  & \new_[78335]_ ;
  assign \new_[78340]_  = \new_[78339]_  & \new_[78332]_ ;
  assign \new_[78344]_  = ~A166 & ~A167;
  assign \new_[78345]_  = ~A169 & \new_[78344]_ ;
  assign \new_[78348]_  = ~A200 & A199;
  assign \new_[78351]_  = A202 & A201;
  assign \new_[78352]_  = \new_[78351]_  & \new_[78348]_ ;
  assign \new_[78353]_  = \new_[78352]_  & \new_[78345]_ ;
  assign \new_[78357]_  = ~A265 & ~A233;
  assign \new_[78358]_  = ~A232 & \new_[78357]_ ;
  assign \new_[78361]_  = A298 & ~A266;
  assign \new_[78364]_  = ~A302 & ~A301;
  assign \new_[78365]_  = \new_[78364]_  & \new_[78361]_ ;
  assign \new_[78366]_  = \new_[78365]_  & \new_[78358]_ ;
  assign \new_[78370]_  = ~A166 & ~A167;
  assign \new_[78371]_  = ~A169 & \new_[78370]_ ;
  assign \new_[78374]_  = ~A200 & A199;
  assign \new_[78377]_  = A203 & A201;
  assign \new_[78378]_  = \new_[78377]_  & \new_[78374]_ ;
  assign \new_[78379]_  = \new_[78378]_  & \new_[78371]_ ;
  assign \new_[78383]_  = A265 & A233;
  assign \new_[78384]_  = A232 & \new_[78383]_ ;
  assign \new_[78387]_  = ~A269 & ~A268;
  assign \new_[78390]_  = ~A300 & ~A299;
  assign \new_[78391]_  = \new_[78390]_  & \new_[78387]_ ;
  assign \new_[78392]_  = \new_[78391]_  & \new_[78384]_ ;
  assign \new_[78396]_  = ~A166 & ~A167;
  assign \new_[78397]_  = ~A169 & \new_[78396]_ ;
  assign \new_[78400]_  = ~A200 & A199;
  assign \new_[78403]_  = A203 & A201;
  assign \new_[78404]_  = \new_[78403]_  & \new_[78400]_ ;
  assign \new_[78405]_  = \new_[78404]_  & \new_[78397]_ ;
  assign \new_[78409]_  = A265 & A233;
  assign \new_[78410]_  = A232 & \new_[78409]_ ;
  assign \new_[78413]_  = ~A269 & ~A268;
  assign \new_[78416]_  = A299 & A298;
  assign \new_[78417]_  = \new_[78416]_  & \new_[78413]_ ;
  assign \new_[78418]_  = \new_[78417]_  & \new_[78410]_ ;
  assign \new_[78422]_  = ~A166 & ~A167;
  assign \new_[78423]_  = ~A169 & \new_[78422]_ ;
  assign \new_[78426]_  = ~A200 & A199;
  assign \new_[78429]_  = A203 & A201;
  assign \new_[78430]_  = \new_[78429]_  & \new_[78426]_ ;
  assign \new_[78431]_  = \new_[78430]_  & \new_[78423]_ ;
  assign \new_[78435]_  = A265 & A233;
  assign \new_[78436]_  = A232 & \new_[78435]_ ;
  assign \new_[78439]_  = ~A269 & ~A268;
  assign \new_[78442]_  = ~A299 & ~A298;
  assign \new_[78443]_  = \new_[78442]_  & \new_[78439]_ ;
  assign \new_[78444]_  = \new_[78443]_  & \new_[78436]_ ;
  assign \new_[78448]_  = ~A166 & ~A167;
  assign \new_[78449]_  = ~A169 & \new_[78448]_ ;
  assign \new_[78452]_  = ~A200 & A199;
  assign \new_[78455]_  = A203 & A201;
  assign \new_[78456]_  = \new_[78455]_  & \new_[78452]_ ;
  assign \new_[78457]_  = \new_[78456]_  & \new_[78449]_ ;
  assign \new_[78461]_  = A265 & A233;
  assign \new_[78462]_  = A232 & \new_[78461]_ ;
  assign \new_[78465]_  = ~A299 & ~A267;
  assign \new_[78468]_  = ~A302 & ~A301;
  assign \new_[78469]_  = \new_[78468]_  & \new_[78465]_ ;
  assign \new_[78470]_  = \new_[78469]_  & \new_[78462]_ ;
  assign \new_[78474]_  = ~A166 & ~A167;
  assign \new_[78475]_  = ~A169 & \new_[78474]_ ;
  assign \new_[78478]_  = ~A200 & A199;
  assign \new_[78481]_  = A203 & A201;
  assign \new_[78482]_  = \new_[78481]_  & \new_[78478]_ ;
  assign \new_[78483]_  = \new_[78482]_  & \new_[78475]_ ;
  assign \new_[78487]_  = A265 & A233;
  assign \new_[78488]_  = A232 & \new_[78487]_ ;
  assign \new_[78491]_  = ~A299 & A266;
  assign \new_[78494]_  = ~A302 & ~A301;
  assign \new_[78495]_  = \new_[78494]_  & \new_[78491]_ ;
  assign \new_[78496]_  = \new_[78495]_  & \new_[78488]_ ;
  assign \new_[78500]_  = ~A166 & ~A167;
  assign \new_[78501]_  = ~A169 & \new_[78500]_ ;
  assign \new_[78504]_  = ~A200 & A199;
  assign \new_[78507]_  = A203 & A201;
  assign \new_[78508]_  = \new_[78507]_  & \new_[78504]_ ;
  assign \new_[78509]_  = \new_[78508]_  & \new_[78501]_ ;
  assign \new_[78513]_  = ~A265 & A233;
  assign \new_[78514]_  = A232 & \new_[78513]_ ;
  assign \new_[78517]_  = ~A299 & ~A266;
  assign \new_[78520]_  = ~A302 & ~A301;
  assign \new_[78521]_  = \new_[78520]_  & \new_[78517]_ ;
  assign \new_[78522]_  = \new_[78521]_  & \new_[78514]_ ;
  assign \new_[78526]_  = ~A166 & ~A167;
  assign \new_[78527]_  = ~A169 & \new_[78526]_ ;
  assign \new_[78530]_  = ~A200 & A199;
  assign \new_[78533]_  = A203 & A201;
  assign \new_[78534]_  = \new_[78533]_  & \new_[78530]_ ;
  assign \new_[78535]_  = \new_[78534]_  & \new_[78527]_ ;
  assign \new_[78539]_  = ~A236 & ~A235;
  assign \new_[78540]_  = ~A233 & \new_[78539]_ ;
  assign \new_[78543]_  = A266 & A265;
  assign \new_[78546]_  = ~A300 & A298;
  assign \new_[78547]_  = \new_[78546]_  & \new_[78543]_ ;
  assign \new_[78548]_  = \new_[78547]_  & \new_[78540]_ ;
  assign \new_[78552]_  = ~A166 & ~A167;
  assign \new_[78553]_  = ~A169 & \new_[78552]_ ;
  assign \new_[78556]_  = ~A200 & A199;
  assign \new_[78559]_  = A203 & A201;
  assign \new_[78560]_  = \new_[78559]_  & \new_[78556]_ ;
  assign \new_[78561]_  = \new_[78560]_  & \new_[78553]_ ;
  assign \new_[78565]_  = ~A236 & ~A235;
  assign \new_[78566]_  = ~A233 & \new_[78565]_ ;
  assign \new_[78569]_  = A266 & A265;
  assign \new_[78572]_  = A299 & A298;
  assign \new_[78573]_  = \new_[78572]_  & \new_[78569]_ ;
  assign \new_[78574]_  = \new_[78573]_  & \new_[78566]_ ;
  assign \new_[78578]_  = ~A166 & ~A167;
  assign \new_[78579]_  = ~A169 & \new_[78578]_ ;
  assign \new_[78582]_  = ~A200 & A199;
  assign \new_[78585]_  = A203 & A201;
  assign \new_[78586]_  = \new_[78585]_  & \new_[78582]_ ;
  assign \new_[78587]_  = \new_[78586]_  & \new_[78579]_ ;
  assign \new_[78591]_  = ~A236 & ~A235;
  assign \new_[78592]_  = ~A233 & \new_[78591]_ ;
  assign \new_[78595]_  = A266 & A265;
  assign \new_[78598]_  = ~A299 & ~A298;
  assign \new_[78599]_  = \new_[78598]_  & \new_[78595]_ ;
  assign \new_[78600]_  = \new_[78599]_  & \new_[78592]_ ;
  assign \new_[78604]_  = ~A166 & ~A167;
  assign \new_[78605]_  = ~A169 & \new_[78604]_ ;
  assign \new_[78608]_  = ~A200 & A199;
  assign \new_[78611]_  = A203 & A201;
  assign \new_[78612]_  = \new_[78611]_  & \new_[78608]_ ;
  assign \new_[78613]_  = \new_[78612]_  & \new_[78605]_ ;
  assign \new_[78617]_  = ~A236 & ~A235;
  assign \new_[78618]_  = ~A233 & \new_[78617]_ ;
  assign \new_[78621]_  = ~A267 & ~A266;
  assign \new_[78624]_  = ~A300 & A298;
  assign \new_[78625]_  = \new_[78624]_  & \new_[78621]_ ;
  assign \new_[78626]_  = \new_[78625]_  & \new_[78618]_ ;
  assign \new_[78630]_  = ~A166 & ~A167;
  assign \new_[78631]_  = ~A169 & \new_[78630]_ ;
  assign \new_[78634]_  = ~A200 & A199;
  assign \new_[78637]_  = A203 & A201;
  assign \new_[78638]_  = \new_[78637]_  & \new_[78634]_ ;
  assign \new_[78639]_  = \new_[78638]_  & \new_[78631]_ ;
  assign \new_[78643]_  = ~A236 & ~A235;
  assign \new_[78644]_  = ~A233 & \new_[78643]_ ;
  assign \new_[78647]_  = ~A267 & ~A266;
  assign \new_[78650]_  = A299 & A298;
  assign \new_[78651]_  = \new_[78650]_  & \new_[78647]_ ;
  assign \new_[78652]_  = \new_[78651]_  & \new_[78644]_ ;
  assign \new_[78656]_  = ~A166 & ~A167;
  assign \new_[78657]_  = ~A169 & \new_[78656]_ ;
  assign \new_[78660]_  = ~A200 & A199;
  assign \new_[78663]_  = A203 & A201;
  assign \new_[78664]_  = \new_[78663]_  & \new_[78660]_ ;
  assign \new_[78665]_  = \new_[78664]_  & \new_[78657]_ ;
  assign \new_[78669]_  = ~A236 & ~A235;
  assign \new_[78670]_  = ~A233 & \new_[78669]_ ;
  assign \new_[78673]_  = ~A267 & ~A266;
  assign \new_[78676]_  = ~A299 & ~A298;
  assign \new_[78677]_  = \new_[78676]_  & \new_[78673]_ ;
  assign \new_[78678]_  = \new_[78677]_  & \new_[78670]_ ;
  assign \new_[78682]_  = ~A166 & ~A167;
  assign \new_[78683]_  = ~A169 & \new_[78682]_ ;
  assign \new_[78686]_  = ~A200 & A199;
  assign \new_[78689]_  = A203 & A201;
  assign \new_[78690]_  = \new_[78689]_  & \new_[78686]_ ;
  assign \new_[78691]_  = \new_[78690]_  & \new_[78683]_ ;
  assign \new_[78695]_  = ~A236 & ~A235;
  assign \new_[78696]_  = ~A233 & \new_[78695]_ ;
  assign \new_[78699]_  = ~A266 & ~A265;
  assign \new_[78702]_  = ~A300 & A298;
  assign \new_[78703]_  = \new_[78702]_  & \new_[78699]_ ;
  assign \new_[78704]_  = \new_[78703]_  & \new_[78696]_ ;
  assign \new_[78708]_  = ~A166 & ~A167;
  assign \new_[78709]_  = ~A169 & \new_[78708]_ ;
  assign \new_[78712]_  = ~A200 & A199;
  assign \new_[78715]_  = A203 & A201;
  assign \new_[78716]_  = \new_[78715]_  & \new_[78712]_ ;
  assign \new_[78717]_  = \new_[78716]_  & \new_[78709]_ ;
  assign \new_[78721]_  = ~A236 & ~A235;
  assign \new_[78722]_  = ~A233 & \new_[78721]_ ;
  assign \new_[78725]_  = ~A266 & ~A265;
  assign \new_[78728]_  = A299 & A298;
  assign \new_[78729]_  = \new_[78728]_  & \new_[78725]_ ;
  assign \new_[78730]_  = \new_[78729]_  & \new_[78722]_ ;
  assign \new_[78734]_  = ~A166 & ~A167;
  assign \new_[78735]_  = ~A169 & \new_[78734]_ ;
  assign \new_[78738]_  = ~A200 & A199;
  assign \new_[78741]_  = A203 & A201;
  assign \new_[78742]_  = \new_[78741]_  & \new_[78738]_ ;
  assign \new_[78743]_  = \new_[78742]_  & \new_[78735]_ ;
  assign \new_[78747]_  = ~A236 & ~A235;
  assign \new_[78748]_  = ~A233 & \new_[78747]_ ;
  assign \new_[78751]_  = ~A266 & ~A265;
  assign \new_[78754]_  = ~A299 & ~A298;
  assign \new_[78755]_  = \new_[78754]_  & \new_[78751]_ ;
  assign \new_[78756]_  = \new_[78755]_  & \new_[78748]_ ;
  assign \new_[78760]_  = ~A166 & ~A167;
  assign \new_[78761]_  = ~A169 & \new_[78760]_ ;
  assign \new_[78764]_  = ~A200 & A199;
  assign \new_[78767]_  = A203 & A201;
  assign \new_[78768]_  = \new_[78767]_  & \new_[78764]_ ;
  assign \new_[78769]_  = \new_[78768]_  & \new_[78761]_ ;
  assign \new_[78773]_  = A265 & ~A234;
  assign \new_[78774]_  = ~A233 & \new_[78773]_ ;
  assign \new_[78777]_  = A298 & A266;
  assign \new_[78780]_  = ~A302 & ~A301;
  assign \new_[78781]_  = \new_[78780]_  & \new_[78777]_ ;
  assign \new_[78782]_  = \new_[78781]_  & \new_[78774]_ ;
  assign \new_[78786]_  = ~A166 & ~A167;
  assign \new_[78787]_  = ~A169 & \new_[78786]_ ;
  assign \new_[78790]_  = ~A200 & A199;
  assign \new_[78793]_  = A203 & A201;
  assign \new_[78794]_  = \new_[78793]_  & \new_[78790]_ ;
  assign \new_[78795]_  = \new_[78794]_  & \new_[78787]_ ;
  assign \new_[78799]_  = ~A266 & ~A234;
  assign \new_[78800]_  = ~A233 & \new_[78799]_ ;
  assign \new_[78803]_  = ~A269 & ~A268;
  assign \new_[78806]_  = ~A300 & A298;
  assign \new_[78807]_  = \new_[78806]_  & \new_[78803]_ ;
  assign \new_[78808]_  = \new_[78807]_  & \new_[78800]_ ;
  assign \new_[78812]_  = ~A166 & ~A167;
  assign \new_[78813]_  = ~A169 & \new_[78812]_ ;
  assign \new_[78816]_  = ~A200 & A199;
  assign \new_[78819]_  = A203 & A201;
  assign \new_[78820]_  = \new_[78819]_  & \new_[78816]_ ;
  assign \new_[78821]_  = \new_[78820]_  & \new_[78813]_ ;
  assign \new_[78825]_  = ~A266 & ~A234;
  assign \new_[78826]_  = ~A233 & \new_[78825]_ ;
  assign \new_[78829]_  = ~A269 & ~A268;
  assign \new_[78832]_  = A299 & A298;
  assign \new_[78833]_  = \new_[78832]_  & \new_[78829]_ ;
  assign \new_[78834]_  = \new_[78833]_  & \new_[78826]_ ;
  assign \new_[78838]_  = ~A166 & ~A167;
  assign \new_[78839]_  = ~A169 & \new_[78838]_ ;
  assign \new_[78842]_  = ~A200 & A199;
  assign \new_[78845]_  = A203 & A201;
  assign \new_[78846]_  = \new_[78845]_  & \new_[78842]_ ;
  assign \new_[78847]_  = \new_[78846]_  & \new_[78839]_ ;
  assign \new_[78851]_  = ~A266 & ~A234;
  assign \new_[78852]_  = ~A233 & \new_[78851]_ ;
  assign \new_[78855]_  = ~A269 & ~A268;
  assign \new_[78858]_  = ~A299 & ~A298;
  assign \new_[78859]_  = \new_[78858]_  & \new_[78855]_ ;
  assign \new_[78860]_  = \new_[78859]_  & \new_[78852]_ ;
  assign \new_[78864]_  = ~A166 & ~A167;
  assign \new_[78865]_  = ~A169 & \new_[78864]_ ;
  assign \new_[78868]_  = ~A200 & A199;
  assign \new_[78871]_  = A203 & A201;
  assign \new_[78872]_  = \new_[78871]_  & \new_[78868]_ ;
  assign \new_[78873]_  = \new_[78872]_  & \new_[78865]_ ;
  assign \new_[78877]_  = ~A266 & ~A234;
  assign \new_[78878]_  = ~A233 & \new_[78877]_ ;
  assign \new_[78881]_  = A298 & ~A267;
  assign \new_[78884]_  = ~A302 & ~A301;
  assign \new_[78885]_  = \new_[78884]_  & \new_[78881]_ ;
  assign \new_[78886]_  = \new_[78885]_  & \new_[78878]_ ;
  assign \new_[78890]_  = ~A166 & ~A167;
  assign \new_[78891]_  = ~A169 & \new_[78890]_ ;
  assign \new_[78894]_  = ~A200 & A199;
  assign \new_[78897]_  = A203 & A201;
  assign \new_[78898]_  = \new_[78897]_  & \new_[78894]_ ;
  assign \new_[78899]_  = \new_[78898]_  & \new_[78891]_ ;
  assign \new_[78903]_  = ~A265 & ~A234;
  assign \new_[78904]_  = ~A233 & \new_[78903]_ ;
  assign \new_[78907]_  = A298 & ~A266;
  assign \new_[78910]_  = ~A302 & ~A301;
  assign \new_[78911]_  = \new_[78910]_  & \new_[78907]_ ;
  assign \new_[78912]_  = \new_[78911]_  & \new_[78904]_ ;
  assign \new_[78916]_  = ~A166 & ~A167;
  assign \new_[78917]_  = ~A169 & \new_[78916]_ ;
  assign \new_[78920]_  = ~A200 & A199;
  assign \new_[78923]_  = A203 & A201;
  assign \new_[78924]_  = \new_[78923]_  & \new_[78920]_ ;
  assign \new_[78925]_  = \new_[78924]_  & \new_[78917]_ ;
  assign \new_[78929]_  = A265 & ~A233;
  assign \new_[78930]_  = ~A232 & \new_[78929]_ ;
  assign \new_[78933]_  = A298 & A266;
  assign \new_[78936]_  = ~A302 & ~A301;
  assign \new_[78937]_  = \new_[78936]_  & \new_[78933]_ ;
  assign \new_[78938]_  = \new_[78937]_  & \new_[78930]_ ;
  assign \new_[78942]_  = ~A166 & ~A167;
  assign \new_[78943]_  = ~A169 & \new_[78942]_ ;
  assign \new_[78946]_  = ~A200 & A199;
  assign \new_[78949]_  = A203 & A201;
  assign \new_[78950]_  = \new_[78949]_  & \new_[78946]_ ;
  assign \new_[78951]_  = \new_[78950]_  & \new_[78943]_ ;
  assign \new_[78955]_  = ~A266 & ~A233;
  assign \new_[78956]_  = ~A232 & \new_[78955]_ ;
  assign \new_[78959]_  = ~A269 & ~A268;
  assign \new_[78962]_  = ~A300 & A298;
  assign \new_[78963]_  = \new_[78962]_  & \new_[78959]_ ;
  assign \new_[78964]_  = \new_[78963]_  & \new_[78956]_ ;
  assign \new_[78968]_  = ~A166 & ~A167;
  assign \new_[78969]_  = ~A169 & \new_[78968]_ ;
  assign \new_[78972]_  = ~A200 & A199;
  assign \new_[78975]_  = A203 & A201;
  assign \new_[78976]_  = \new_[78975]_  & \new_[78972]_ ;
  assign \new_[78977]_  = \new_[78976]_  & \new_[78969]_ ;
  assign \new_[78981]_  = ~A266 & ~A233;
  assign \new_[78982]_  = ~A232 & \new_[78981]_ ;
  assign \new_[78985]_  = ~A269 & ~A268;
  assign \new_[78988]_  = A299 & A298;
  assign \new_[78989]_  = \new_[78988]_  & \new_[78985]_ ;
  assign \new_[78990]_  = \new_[78989]_  & \new_[78982]_ ;
  assign \new_[78994]_  = ~A166 & ~A167;
  assign \new_[78995]_  = ~A169 & \new_[78994]_ ;
  assign \new_[78998]_  = ~A200 & A199;
  assign \new_[79001]_  = A203 & A201;
  assign \new_[79002]_  = \new_[79001]_  & \new_[78998]_ ;
  assign \new_[79003]_  = \new_[79002]_  & \new_[78995]_ ;
  assign \new_[79007]_  = ~A266 & ~A233;
  assign \new_[79008]_  = ~A232 & \new_[79007]_ ;
  assign \new_[79011]_  = ~A269 & ~A268;
  assign \new_[79014]_  = ~A299 & ~A298;
  assign \new_[79015]_  = \new_[79014]_  & \new_[79011]_ ;
  assign \new_[79016]_  = \new_[79015]_  & \new_[79008]_ ;
  assign \new_[79020]_  = ~A166 & ~A167;
  assign \new_[79021]_  = ~A169 & \new_[79020]_ ;
  assign \new_[79024]_  = ~A200 & A199;
  assign \new_[79027]_  = A203 & A201;
  assign \new_[79028]_  = \new_[79027]_  & \new_[79024]_ ;
  assign \new_[79029]_  = \new_[79028]_  & \new_[79021]_ ;
  assign \new_[79033]_  = ~A266 & ~A233;
  assign \new_[79034]_  = ~A232 & \new_[79033]_ ;
  assign \new_[79037]_  = A298 & ~A267;
  assign \new_[79040]_  = ~A302 & ~A301;
  assign \new_[79041]_  = \new_[79040]_  & \new_[79037]_ ;
  assign \new_[79042]_  = \new_[79041]_  & \new_[79034]_ ;
  assign \new_[79046]_  = ~A166 & ~A167;
  assign \new_[79047]_  = ~A169 & \new_[79046]_ ;
  assign \new_[79050]_  = ~A200 & A199;
  assign \new_[79053]_  = A203 & A201;
  assign \new_[79054]_  = \new_[79053]_  & \new_[79050]_ ;
  assign \new_[79055]_  = \new_[79054]_  & \new_[79047]_ ;
  assign \new_[79059]_  = ~A265 & ~A233;
  assign \new_[79060]_  = ~A232 & \new_[79059]_ ;
  assign \new_[79063]_  = A298 & ~A266;
  assign \new_[79066]_  = ~A302 & ~A301;
  assign \new_[79067]_  = \new_[79066]_  & \new_[79063]_ ;
  assign \new_[79068]_  = \new_[79067]_  & \new_[79060]_ ;
  assign \new_[79072]_  = A167 & ~A168;
  assign \new_[79073]_  = ~A169 & \new_[79072]_ ;
  assign \new_[79076]_  = ~A199 & A166;
  assign \new_[79079]_  = A232 & A200;
  assign \new_[79080]_  = \new_[79079]_  & \new_[79076]_ ;
  assign \new_[79081]_  = \new_[79080]_  & \new_[79073]_ ;
  assign \new_[79085]_  = ~A268 & A265;
  assign \new_[79086]_  = A233 & \new_[79085]_ ;
  assign \new_[79089]_  = ~A299 & ~A269;
  assign \new_[79092]_  = ~A302 & ~A301;
  assign \new_[79093]_  = \new_[79092]_  & \new_[79089]_ ;
  assign \new_[79094]_  = \new_[79093]_  & \new_[79086]_ ;
  assign \new_[79098]_  = A167 & ~A168;
  assign \new_[79099]_  = ~A169 & \new_[79098]_ ;
  assign \new_[79102]_  = ~A199 & A166;
  assign \new_[79105]_  = ~A233 & A200;
  assign \new_[79106]_  = \new_[79105]_  & \new_[79102]_ ;
  assign \new_[79107]_  = \new_[79106]_  & \new_[79099]_ ;
  assign \new_[79111]_  = A265 & ~A236;
  assign \new_[79112]_  = ~A235 & \new_[79111]_ ;
  assign \new_[79115]_  = A298 & A266;
  assign \new_[79118]_  = ~A302 & ~A301;
  assign \new_[79119]_  = \new_[79118]_  & \new_[79115]_ ;
  assign \new_[79120]_  = \new_[79119]_  & \new_[79112]_ ;
  assign \new_[79124]_  = A167 & ~A168;
  assign \new_[79125]_  = ~A169 & \new_[79124]_ ;
  assign \new_[79128]_  = ~A199 & A166;
  assign \new_[79131]_  = ~A233 & A200;
  assign \new_[79132]_  = \new_[79131]_  & \new_[79128]_ ;
  assign \new_[79133]_  = \new_[79132]_  & \new_[79125]_ ;
  assign \new_[79137]_  = ~A266 & ~A236;
  assign \new_[79138]_  = ~A235 & \new_[79137]_ ;
  assign \new_[79141]_  = ~A269 & ~A268;
  assign \new_[79144]_  = ~A300 & A298;
  assign \new_[79145]_  = \new_[79144]_  & \new_[79141]_ ;
  assign \new_[79146]_  = \new_[79145]_  & \new_[79138]_ ;
  assign \new_[79150]_  = A167 & ~A168;
  assign \new_[79151]_  = ~A169 & \new_[79150]_ ;
  assign \new_[79154]_  = ~A199 & A166;
  assign \new_[79157]_  = ~A233 & A200;
  assign \new_[79158]_  = \new_[79157]_  & \new_[79154]_ ;
  assign \new_[79159]_  = \new_[79158]_  & \new_[79151]_ ;
  assign \new_[79163]_  = ~A266 & ~A236;
  assign \new_[79164]_  = ~A235 & \new_[79163]_ ;
  assign \new_[79167]_  = ~A269 & ~A268;
  assign \new_[79170]_  = A299 & A298;
  assign \new_[79171]_  = \new_[79170]_  & \new_[79167]_ ;
  assign \new_[79172]_  = \new_[79171]_  & \new_[79164]_ ;
  assign \new_[79176]_  = A167 & ~A168;
  assign \new_[79177]_  = ~A169 & \new_[79176]_ ;
  assign \new_[79180]_  = ~A199 & A166;
  assign \new_[79183]_  = ~A233 & A200;
  assign \new_[79184]_  = \new_[79183]_  & \new_[79180]_ ;
  assign \new_[79185]_  = \new_[79184]_  & \new_[79177]_ ;
  assign \new_[79189]_  = ~A266 & ~A236;
  assign \new_[79190]_  = ~A235 & \new_[79189]_ ;
  assign \new_[79193]_  = ~A269 & ~A268;
  assign \new_[79196]_  = ~A299 & ~A298;
  assign \new_[79197]_  = \new_[79196]_  & \new_[79193]_ ;
  assign \new_[79198]_  = \new_[79197]_  & \new_[79190]_ ;
  assign \new_[79202]_  = A167 & ~A168;
  assign \new_[79203]_  = ~A169 & \new_[79202]_ ;
  assign \new_[79206]_  = ~A199 & A166;
  assign \new_[79209]_  = ~A233 & A200;
  assign \new_[79210]_  = \new_[79209]_  & \new_[79206]_ ;
  assign \new_[79211]_  = \new_[79210]_  & \new_[79203]_ ;
  assign \new_[79215]_  = ~A266 & ~A236;
  assign \new_[79216]_  = ~A235 & \new_[79215]_ ;
  assign \new_[79219]_  = A298 & ~A267;
  assign \new_[79222]_  = ~A302 & ~A301;
  assign \new_[79223]_  = \new_[79222]_  & \new_[79219]_ ;
  assign \new_[79224]_  = \new_[79223]_  & \new_[79216]_ ;
  assign \new_[79228]_  = A167 & ~A168;
  assign \new_[79229]_  = ~A169 & \new_[79228]_ ;
  assign \new_[79232]_  = ~A199 & A166;
  assign \new_[79235]_  = ~A233 & A200;
  assign \new_[79236]_  = \new_[79235]_  & \new_[79232]_ ;
  assign \new_[79237]_  = \new_[79236]_  & \new_[79229]_ ;
  assign \new_[79241]_  = ~A265 & ~A236;
  assign \new_[79242]_  = ~A235 & \new_[79241]_ ;
  assign \new_[79245]_  = A298 & ~A266;
  assign \new_[79248]_  = ~A302 & ~A301;
  assign \new_[79249]_  = \new_[79248]_  & \new_[79245]_ ;
  assign \new_[79250]_  = \new_[79249]_  & \new_[79242]_ ;
  assign \new_[79254]_  = A167 & ~A168;
  assign \new_[79255]_  = ~A169 & \new_[79254]_ ;
  assign \new_[79258]_  = ~A199 & A166;
  assign \new_[79261]_  = ~A233 & A200;
  assign \new_[79262]_  = \new_[79261]_  & \new_[79258]_ ;
  assign \new_[79263]_  = \new_[79262]_  & \new_[79255]_ ;
  assign \new_[79267]_  = ~A268 & ~A266;
  assign \new_[79268]_  = ~A234 & \new_[79267]_ ;
  assign \new_[79271]_  = A298 & ~A269;
  assign \new_[79274]_  = ~A302 & ~A301;
  assign \new_[79275]_  = \new_[79274]_  & \new_[79271]_ ;
  assign \new_[79276]_  = \new_[79275]_  & \new_[79268]_ ;
  assign \new_[79280]_  = A167 & ~A168;
  assign \new_[79281]_  = ~A169 & \new_[79280]_ ;
  assign \new_[79284]_  = ~A199 & A166;
  assign \new_[79287]_  = A232 & A200;
  assign \new_[79288]_  = \new_[79287]_  & \new_[79284]_ ;
  assign \new_[79289]_  = \new_[79288]_  & \new_[79281]_ ;
  assign \new_[79293]_  = A235 & A234;
  assign \new_[79294]_  = ~A233 & \new_[79293]_ ;
  assign \new_[79297]_  = ~A299 & A298;
  assign \new_[79300]_  = A301 & A300;
  assign \new_[79301]_  = \new_[79300]_  & \new_[79297]_ ;
  assign \new_[79302]_  = \new_[79301]_  & \new_[79294]_ ;
  assign \new_[79306]_  = A167 & ~A168;
  assign \new_[79307]_  = ~A169 & \new_[79306]_ ;
  assign \new_[79310]_  = ~A199 & A166;
  assign \new_[79313]_  = A232 & A200;
  assign \new_[79314]_  = \new_[79313]_  & \new_[79310]_ ;
  assign \new_[79315]_  = \new_[79314]_  & \new_[79307]_ ;
  assign \new_[79319]_  = A235 & A234;
  assign \new_[79320]_  = ~A233 & \new_[79319]_ ;
  assign \new_[79323]_  = ~A299 & A298;
  assign \new_[79326]_  = A302 & A300;
  assign \new_[79327]_  = \new_[79326]_  & \new_[79323]_ ;
  assign \new_[79328]_  = \new_[79327]_  & \new_[79320]_ ;
  assign \new_[79332]_  = A167 & ~A168;
  assign \new_[79333]_  = ~A169 & \new_[79332]_ ;
  assign \new_[79336]_  = ~A199 & A166;
  assign \new_[79339]_  = A232 & A200;
  assign \new_[79340]_  = \new_[79339]_  & \new_[79336]_ ;
  assign \new_[79341]_  = \new_[79340]_  & \new_[79333]_ ;
  assign \new_[79345]_  = A235 & A234;
  assign \new_[79346]_  = ~A233 & \new_[79345]_ ;
  assign \new_[79349]_  = ~A266 & A265;
  assign \new_[79352]_  = A268 & A267;
  assign \new_[79353]_  = \new_[79352]_  & \new_[79349]_ ;
  assign \new_[79354]_  = \new_[79353]_  & \new_[79346]_ ;
  assign \new_[79358]_  = A167 & ~A168;
  assign \new_[79359]_  = ~A169 & \new_[79358]_ ;
  assign \new_[79362]_  = ~A199 & A166;
  assign \new_[79365]_  = A232 & A200;
  assign \new_[79366]_  = \new_[79365]_  & \new_[79362]_ ;
  assign \new_[79367]_  = \new_[79366]_  & \new_[79359]_ ;
  assign \new_[79371]_  = A235 & A234;
  assign \new_[79372]_  = ~A233 & \new_[79371]_ ;
  assign \new_[79375]_  = ~A266 & A265;
  assign \new_[79378]_  = A269 & A267;
  assign \new_[79379]_  = \new_[79378]_  & \new_[79375]_ ;
  assign \new_[79380]_  = \new_[79379]_  & \new_[79372]_ ;
  assign \new_[79384]_  = A167 & ~A168;
  assign \new_[79385]_  = ~A169 & \new_[79384]_ ;
  assign \new_[79388]_  = ~A199 & A166;
  assign \new_[79391]_  = A232 & A200;
  assign \new_[79392]_  = \new_[79391]_  & \new_[79388]_ ;
  assign \new_[79393]_  = \new_[79392]_  & \new_[79385]_ ;
  assign \new_[79397]_  = A236 & A234;
  assign \new_[79398]_  = ~A233 & \new_[79397]_ ;
  assign \new_[79401]_  = ~A299 & A298;
  assign \new_[79404]_  = A301 & A300;
  assign \new_[79405]_  = \new_[79404]_  & \new_[79401]_ ;
  assign \new_[79406]_  = \new_[79405]_  & \new_[79398]_ ;
  assign \new_[79410]_  = A167 & ~A168;
  assign \new_[79411]_  = ~A169 & \new_[79410]_ ;
  assign \new_[79414]_  = ~A199 & A166;
  assign \new_[79417]_  = A232 & A200;
  assign \new_[79418]_  = \new_[79417]_  & \new_[79414]_ ;
  assign \new_[79419]_  = \new_[79418]_  & \new_[79411]_ ;
  assign \new_[79423]_  = A236 & A234;
  assign \new_[79424]_  = ~A233 & \new_[79423]_ ;
  assign \new_[79427]_  = ~A299 & A298;
  assign \new_[79430]_  = A302 & A300;
  assign \new_[79431]_  = \new_[79430]_  & \new_[79427]_ ;
  assign \new_[79432]_  = \new_[79431]_  & \new_[79424]_ ;
  assign \new_[79436]_  = A167 & ~A168;
  assign \new_[79437]_  = ~A169 & \new_[79436]_ ;
  assign \new_[79440]_  = ~A199 & A166;
  assign \new_[79443]_  = A232 & A200;
  assign \new_[79444]_  = \new_[79443]_  & \new_[79440]_ ;
  assign \new_[79445]_  = \new_[79444]_  & \new_[79437]_ ;
  assign \new_[79449]_  = A236 & A234;
  assign \new_[79450]_  = ~A233 & \new_[79449]_ ;
  assign \new_[79453]_  = ~A266 & A265;
  assign \new_[79456]_  = A268 & A267;
  assign \new_[79457]_  = \new_[79456]_  & \new_[79453]_ ;
  assign \new_[79458]_  = \new_[79457]_  & \new_[79450]_ ;
  assign \new_[79462]_  = A167 & ~A168;
  assign \new_[79463]_  = ~A169 & \new_[79462]_ ;
  assign \new_[79466]_  = ~A199 & A166;
  assign \new_[79469]_  = A232 & A200;
  assign \new_[79470]_  = \new_[79469]_  & \new_[79466]_ ;
  assign \new_[79471]_  = \new_[79470]_  & \new_[79463]_ ;
  assign \new_[79475]_  = A236 & A234;
  assign \new_[79476]_  = ~A233 & \new_[79475]_ ;
  assign \new_[79479]_  = ~A266 & A265;
  assign \new_[79482]_  = A269 & A267;
  assign \new_[79483]_  = \new_[79482]_  & \new_[79479]_ ;
  assign \new_[79484]_  = \new_[79483]_  & \new_[79476]_ ;
  assign \new_[79488]_  = A167 & ~A168;
  assign \new_[79489]_  = ~A169 & \new_[79488]_ ;
  assign \new_[79492]_  = ~A199 & A166;
  assign \new_[79495]_  = ~A232 & A200;
  assign \new_[79496]_  = \new_[79495]_  & \new_[79492]_ ;
  assign \new_[79497]_  = \new_[79496]_  & \new_[79489]_ ;
  assign \new_[79501]_  = ~A268 & ~A266;
  assign \new_[79502]_  = ~A233 & \new_[79501]_ ;
  assign \new_[79505]_  = A298 & ~A269;
  assign \new_[79508]_  = ~A302 & ~A301;
  assign \new_[79509]_  = \new_[79508]_  & \new_[79505]_ ;
  assign \new_[79510]_  = \new_[79509]_  & \new_[79502]_ ;
  assign \new_[79514]_  = A167 & ~A168;
  assign \new_[79515]_  = ~A169 & \new_[79514]_ ;
  assign \new_[79518]_  = A199 & A166;
  assign \new_[79521]_  = A201 & ~A200;
  assign \new_[79522]_  = \new_[79521]_  & \new_[79518]_ ;
  assign \new_[79523]_  = \new_[79522]_  & \new_[79515]_ ;
  assign \new_[79527]_  = A233 & A232;
  assign \new_[79528]_  = A202 & \new_[79527]_ ;
  assign \new_[79531]_  = ~A267 & A265;
  assign \new_[79534]_  = ~A300 & ~A299;
  assign \new_[79535]_  = \new_[79534]_  & \new_[79531]_ ;
  assign \new_[79536]_  = \new_[79535]_  & \new_[79528]_ ;
  assign \new_[79540]_  = A167 & ~A168;
  assign \new_[79541]_  = ~A169 & \new_[79540]_ ;
  assign \new_[79544]_  = A199 & A166;
  assign \new_[79547]_  = A201 & ~A200;
  assign \new_[79548]_  = \new_[79547]_  & \new_[79544]_ ;
  assign \new_[79549]_  = \new_[79548]_  & \new_[79541]_ ;
  assign \new_[79553]_  = A233 & A232;
  assign \new_[79554]_  = A202 & \new_[79553]_ ;
  assign \new_[79557]_  = ~A267 & A265;
  assign \new_[79560]_  = A299 & A298;
  assign \new_[79561]_  = \new_[79560]_  & \new_[79557]_ ;
  assign \new_[79562]_  = \new_[79561]_  & \new_[79554]_ ;
  assign \new_[79566]_  = A167 & ~A168;
  assign \new_[79567]_  = ~A169 & \new_[79566]_ ;
  assign \new_[79570]_  = A199 & A166;
  assign \new_[79573]_  = A201 & ~A200;
  assign \new_[79574]_  = \new_[79573]_  & \new_[79570]_ ;
  assign \new_[79575]_  = \new_[79574]_  & \new_[79567]_ ;
  assign \new_[79579]_  = A233 & A232;
  assign \new_[79580]_  = A202 & \new_[79579]_ ;
  assign \new_[79583]_  = ~A267 & A265;
  assign \new_[79586]_  = ~A299 & ~A298;
  assign \new_[79587]_  = \new_[79586]_  & \new_[79583]_ ;
  assign \new_[79588]_  = \new_[79587]_  & \new_[79580]_ ;
  assign \new_[79592]_  = A167 & ~A168;
  assign \new_[79593]_  = ~A169 & \new_[79592]_ ;
  assign \new_[79596]_  = A199 & A166;
  assign \new_[79599]_  = A201 & ~A200;
  assign \new_[79600]_  = \new_[79599]_  & \new_[79596]_ ;
  assign \new_[79601]_  = \new_[79600]_  & \new_[79593]_ ;
  assign \new_[79605]_  = A233 & A232;
  assign \new_[79606]_  = A202 & \new_[79605]_ ;
  assign \new_[79609]_  = A266 & A265;
  assign \new_[79612]_  = ~A300 & ~A299;
  assign \new_[79613]_  = \new_[79612]_  & \new_[79609]_ ;
  assign \new_[79614]_  = \new_[79613]_  & \new_[79606]_ ;
  assign \new_[79618]_  = A167 & ~A168;
  assign \new_[79619]_  = ~A169 & \new_[79618]_ ;
  assign \new_[79622]_  = A199 & A166;
  assign \new_[79625]_  = A201 & ~A200;
  assign \new_[79626]_  = \new_[79625]_  & \new_[79622]_ ;
  assign \new_[79627]_  = \new_[79626]_  & \new_[79619]_ ;
  assign \new_[79631]_  = A233 & A232;
  assign \new_[79632]_  = A202 & \new_[79631]_ ;
  assign \new_[79635]_  = A266 & A265;
  assign \new_[79638]_  = A299 & A298;
  assign \new_[79639]_  = \new_[79638]_  & \new_[79635]_ ;
  assign \new_[79640]_  = \new_[79639]_  & \new_[79632]_ ;
  assign \new_[79644]_  = A167 & ~A168;
  assign \new_[79645]_  = ~A169 & \new_[79644]_ ;
  assign \new_[79648]_  = A199 & A166;
  assign \new_[79651]_  = A201 & ~A200;
  assign \new_[79652]_  = \new_[79651]_  & \new_[79648]_ ;
  assign \new_[79653]_  = \new_[79652]_  & \new_[79645]_ ;
  assign \new_[79657]_  = A233 & A232;
  assign \new_[79658]_  = A202 & \new_[79657]_ ;
  assign \new_[79661]_  = A266 & A265;
  assign \new_[79664]_  = ~A299 & ~A298;
  assign \new_[79665]_  = \new_[79664]_  & \new_[79661]_ ;
  assign \new_[79666]_  = \new_[79665]_  & \new_[79658]_ ;
  assign \new_[79670]_  = A167 & ~A168;
  assign \new_[79671]_  = ~A169 & \new_[79670]_ ;
  assign \new_[79674]_  = A199 & A166;
  assign \new_[79677]_  = A201 & ~A200;
  assign \new_[79678]_  = \new_[79677]_  & \new_[79674]_ ;
  assign \new_[79679]_  = \new_[79678]_  & \new_[79671]_ ;
  assign \new_[79683]_  = A233 & A232;
  assign \new_[79684]_  = A202 & \new_[79683]_ ;
  assign \new_[79687]_  = ~A266 & ~A265;
  assign \new_[79690]_  = ~A300 & ~A299;
  assign \new_[79691]_  = \new_[79690]_  & \new_[79687]_ ;
  assign \new_[79692]_  = \new_[79691]_  & \new_[79684]_ ;
  assign \new_[79696]_  = A167 & ~A168;
  assign \new_[79697]_  = ~A169 & \new_[79696]_ ;
  assign \new_[79700]_  = A199 & A166;
  assign \new_[79703]_  = A201 & ~A200;
  assign \new_[79704]_  = \new_[79703]_  & \new_[79700]_ ;
  assign \new_[79705]_  = \new_[79704]_  & \new_[79697]_ ;
  assign \new_[79709]_  = A233 & A232;
  assign \new_[79710]_  = A202 & \new_[79709]_ ;
  assign \new_[79713]_  = ~A266 & ~A265;
  assign \new_[79716]_  = A299 & A298;
  assign \new_[79717]_  = \new_[79716]_  & \new_[79713]_ ;
  assign \new_[79718]_  = \new_[79717]_  & \new_[79710]_ ;
  assign \new_[79722]_  = A167 & ~A168;
  assign \new_[79723]_  = ~A169 & \new_[79722]_ ;
  assign \new_[79726]_  = A199 & A166;
  assign \new_[79729]_  = A201 & ~A200;
  assign \new_[79730]_  = \new_[79729]_  & \new_[79726]_ ;
  assign \new_[79731]_  = \new_[79730]_  & \new_[79723]_ ;
  assign \new_[79735]_  = A233 & A232;
  assign \new_[79736]_  = A202 & \new_[79735]_ ;
  assign \new_[79739]_  = ~A266 & ~A265;
  assign \new_[79742]_  = ~A299 & ~A298;
  assign \new_[79743]_  = \new_[79742]_  & \new_[79739]_ ;
  assign \new_[79744]_  = \new_[79743]_  & \new_[79736]_ ;
  assign \new_[79748]_  = A167 & ~A168;
  assign \new_[79749]_  = ~A169 & \new_[79748]_ ;
  assign \new_[79752]_  = A199 & A166;
  assign \new_[79755]_  = A201 & ~A200;
  assign \new_[79756]_  = \new_[79755]_  & \new_[79752]_ ;
  assign \new_[79757]_  = \new_[79756]_  & \new_[79749]_ ;
  assign \new_[79761]_  = A233 & ~A232;
  assign \new_[79762]_  = A202 & \new_[79761]_ ;
  assign \new_[79765]_  = ~A299 & A298;
  assign \new_[79768]_  = A301 & A300;
  assign \new_[79769]_  = \new_[79768]_  & \new_[79765]_ ;
  assign \new_[79770]_  = \new_[79769]_  & \new_[79762]_ ;
  assign \new_[79774]_  = A167 & ~A168;
  assign \new_[79775]_  = ~A169 & \new_[79774]_ ;
  assign \new_[79778]_  = A199 & A166;
  assign \new_[79781]_  = A201 & ~A200;
  assign \new_[79782]_  = \new_[79781]_  & \new_[79778]_ ;
  assign \new_[79783]_  = \new_[79782]_  & \new_[79775]_ ;
  assign \new_[79787]_  = A233 & ~A232;
  assign \new_[79788]_  = A202 & \new_[79787]_ ;
  assign \new_[79791]_  = ~A299 & A298;
  assign \new_[79794]_  = A302 & A300;
  assign \new_[79795]_  = \new_[79794]_  & \new_[79791]_ ;
  assign \new_[79796]_  = \new_[79795]_  & \new_[79788]_ ;
  assign \new_[79800]_  = A167 & ~A168;
  assign \new_[79801]_  = ~A169 & \new_[79800]_ ;
  assign \new_[79804]_  = A199 & A166;
  assign \new_[79807]_  = A201 & ~A200;
  assign \new_[79808]_  = \new_[79807]_  & \new_[79804]_ ;
  assign \new_[79809]_  = \new_[79808]_  & \new_[79801]_ ;
  assign \new_[79813]_  = A233 & ~A232;
  assign \new_[79814]_  = A202 & \new_[79813]_ ;
  assign \new_[79817]_  = ~A266 & A265;
  assign \new_[79820]_  = A268 & A267;
  assign \new_[79821]_  = \new_[79820]_  & \new_[79817]_ ;
  assign \new_[79822]_  = \new_[79821]_  & \new_[79814]_ ;
  assign \new_[79826]_  = A167 & ~A168;
  assign \new_[79827]_  = ~A169 & \new_[79826]_ ;
  assign \new_[79830]_  = A199 & A166;
  assign \new_[79833]_  = A201 & ~A200;
  assign \new_[79834]_  = \new_[79833]_  & \new_[79830]_ ;
  assign \new_[79835]_  = \new_[79834]_  & \new_[79827]_ ;
  assign \new_[79839]_  = A233 & ~A232;
  assign \new_[79840]_  = A202 & \new_[79839]_ ;
  assign \new_[79843]_  = ~A266 & A265;
  assign \new_[79846]_  = A269 & A267;
  assign \new_[79847]_  = \new_[79846]_  & \new_[79843]_ ;
  assign \new_[79848]_  = \new_[79847]_  & \new_[79840]_ ;
  assign \new_[79852]_  = A167 & ~A168;
  assign \new_[79853]_  = ~A169 & \new_[79852]_ ;
  assign \new_[79856]_  = A199 & A166;
  assign \new_[79859]_  = A201 & ~A200;
  assign \new_[79860]_  = \new_[79859]_  & \new_[79856]_ ;
  assign \new_[79861]_  = \new_[79860]_  & \new_[79853]_ ;
  assign \new_[79865]_  = ~A234 & ~A233;
  assign \new_[79866]_  = A202 & \new_[79865]_ ;
  assign \new_[79869]_  = A266 & A265;
  assign \new_[79872]_  = ~A300 & A298;
  assign \new_[79873]_  = \new_[79872]_  & \new_[79869]_ ;
  assign \new_[79874]_  = \new_[79873]_  & \new_[79866]_ ;
  assign \new_[79878]_  = A167 & ~A168;
  assign \new_[79879]_  = ~A169 & \new_[79878]_ ;
  assign \new_[79882]_  = A199 & A166;
  assign \new_[79885]_  = A201 & ~A200;
  assign \new_[79886]_  = \new_[79885]_  & \new_[79882]_ ;
  assign \new_[79887]_  = \new_[79886]_  & \new_[79879]_ ;
  assign \new_[79891]_  = ~A234 & ~A233;
  assign \new_[79892]_  = A202 & \new_[79891]_ ;
  assign \new_[79895]_  = A266 & A265;
  assign \new_[79898]_  = A299 & A298;
  assign \new_[79899]_  = \new_[79898]_  & \new_[79895]_ ;
  assign \new_[79900]_  = \new_[79899]_  & \new_[79892]_ ;
  assign \new_[79904]_  = A167 & ~A168;
  assign \new_[79905]_  = ~A169 & \new_[79904]_ ;
  assign \new_[79908]_  = A199 & A166;
  assign \new_[79911]_  = A201 & ~A200;
  assign \new_[79912]_  = \new_[79911]_  & \new_[79908]_ ;
  assign \new_[79913]_  = \new_[79912]_  & \new_[79905]_ ;
  assign \new_[79917]_  = ~A234 & ~A233;
  assign \new_[79918]_  = A202 & \new_[79917]_ ;
  assign \new_[79921]_  = A266 & A265;
  assign \new_[79924]_  = ~A299 & ~A298;
  assign \new_[79925]_  = \new_[79924]_  & \new_[79921]_ ;
  assign \new_[79926]_  = \new_[79925]_  & \new_[79918]_ ;
  assign \new_[79930]_  = A167 & ~A168;
  assign \new_[79931]_  = ~A169 & \new_[79930]_ ;
  assign \new_[79934]_  = A199 & A166;
  assign \new_[79937]_  = A201 & ~A200;
  assign \new_[79938]_  = \new_[79937]_  & \new_[79934]_ ;
  assign \new_[79939]_  = \new_[79938]_  & \new_[79931]_ ;
  assign \new_[79943]_  = ~A234 & ~A233;
  assign \new_[79944]_  = A202 & \new_[79943]_ ;
  assign \new_[79947]_  = ~A267 & ~A266;
  assign \new_[79950]_  = ~A300 & A298;
  assign \new_[79951]_  = \new_[79950]_  & \new_[79947]_ ;
  assign \new_[79952]_  = \new_[79951]_  & \new_[79944]_ ;
  assign \new_[79956]_  = A167 & ~A168;
  assign \new_[79957]_  = ~A169 & \new_[79956]_ ;
  assign \new_[79960]_  = A199 & A166;
  assign \new_[79963]_  = A201 & ~A200;
  assign \new_[79964]_  = \new_[79963]_  & \new_[79960]_ ;
  assign \new_[79965]_  = \new_[79964]_  & \new_[79957]_ ;
  assign \new_[79969]_  = ~A234 & ~A233;
  assign \new_[79970]_  = A202 & \new_[79969]_ ;
  assign \new_[79973]_  = ~A267 & ~A266;
  assign \new_[79976]_  = A299 & A298;
  assign \new_[79977]_  = \new_[79976]_  & \new_[79973]_ ;
  assign \new_[79978]_  = \new_[79977]_  & \new_[79970]_ ;
  assign \new_[79982]_  = A167 & ~A168;
  assign \new_[79983]_  = ~A169 & \new_[79982]_ ;
  assign \new_[79986]_  = A199 & A166;
  assign \new_[79989]_  = A201 & ~A200;
  assign \new_[79990]_  = \new_[79989]_  & \new_[79986]_ ;
  assign \new_[79991]_  = \new_[79990]_  & \new_[79983]_ ;
  assign \new_[79995]_  = ~A234 & ~A233;
  assign \new_[79996]_  = A202 & \new_[79995]_ ;
  assign \new_[79999]_  = ~A267 & ~A266;
  assign \new_[80002]_  = ~A299 & ~A298;
  assign \new_[80003]_  = \new_[80002]_  & \new_[79999]_ ;
  assign \new_[80004]_  = \new_[80003]_  & \new_[79996]_ ;
  assign \new_[80008]_  = A167 & ~A168;
  assign \new_[80009]_  = ~A169 & \new_[80008]_ ;
  assign \new_[80012]_  = A199 & A166;
  assign \new_[80015]_  = A201 & ~A200;
  assign \new_[80016]_  = \new_[80015]_  & \new_[80012]_ ;
  assign \new_[80017]_  = \new_[80016]_  & \new_[80009]_ ;
  assign \new_[80021]_  = ~A234 & ~A233;
  assign \new_[80022]_  = A202 & \new_[80021]_ ;
  assign \new_[80025]_  = ~A266 & ~A265;
  assign \new_[80028]_  = ~A300 & A298;
  assign \new_[80029]_  = \new_[80028]_  & \new_[80025]_ ;
  assign \new_[80030]_  = \new_[80029]_  & \new_[80022]_ ;
  assign \new_[80034]_  = A167 & ~A168;
  assign \new_[80035]_  = ~A169 & \new_[80034]_ ;
  assign \new_[80038]_  = A199 & A166;
  assign \new_[80041]_  = A201 & ~A200;
  assign \new_[80042]_  = \new_[80041]_  & \new_[80038]_ ;
  assign \new_[80043]_  = \new_[80042]_  & \new_[80035]_ ;
  assign \new_[80047]_  = ~A234 & ~A233;
  assign \new_[80048]_  = A202 & \new_[80047]_ ;
  assign \new_[80051]_  = ~A266 & ~A265;
  assign \new_[80054]_  = A299 & A298;
  assign \new_[80055]_  = \new_[80054]_  & \new_[80051]_ ;
  assign \new_[80056]_  = \new_[80055]_  & \new_[80048]_ ;
  assign \new_[80060]_  = A167 & ~A168;
  assign \new_[80061]_  = ~A169 & \new_[80060]_ ;
  assign \new_[80064]_  = A199 & A166;
  assign \new_[80067]_  = A201 & ~A200;
  assign \new_[80068]_  = \new_[80067]_  & \new_[80064]_ ;
  assign \new_[80069]_  = \new_[80068]_  & \new_[80061]_ ;
  assign \new_[80073]_  = ~A234 & ~A233;
  assign \new_[80074]_  = A202 & \new_[80073]_ ;
  assign \new_[80077]_  = ~A266 & ~A265;
  assign \new_[80080]_  = ~A299 & ~A298;
  assign \new_[80081]_  = \new_[80080]_  & \new_[80077]_ ;
  assign \new_[80082]_  = \new_[80081]_  & \new_[80074]_ ;
  assign \new_[80086]_  = A167 & ~A168;
  assign \new_[80087]_  = ~A169 & \new_[80086]_ ;
  assign \new_[80090]_  = A199 & A166;
  assign \new_[80093]_  = A201 & ~A200;
  assign \new_[80094]_  = \new_[80093]_  & \new_[80090]_ ;
  assign \new_[80095]_  = \new_[80094]_  & \new_[80087]_ ;
  assign \new_[80099]_  = ~A233 & A232;
  assign \new_[80100]_  = A202 & \new_[80099]_ ;
  assign \new_[80103]_  = A235 & A234;
  assign \new_[80106]_  = A299 & ~A298;
  assign \new_[80107]_  = \new_[80106]_  & \new_[80103]_ ;
  assign \new_[80108]_  = \new_[80107]_  & \new_[80100]_ ;
  assign \new_[80112]_  = A167 & ~A168;
  assign \new_[80113]_  = ~A169 & \new_[80112]_ ;
  assign \new_[80116]_  = A199 & A166;
  assign \new_[80119]_  = A201 & ~A200;
  assign \new_[80120]_  = \new_[80119]_  & \new_[80116]_ ;
  assign \new_[80121]_  = \new_[80120]_  & \new_[80113]_ ;
  assign \new_[80125]_  = ~A233 & A232;
  assign \new_[80126]_  = A202 & \new_[80125]_ ;
  assign \new_[80129]_  = A235 & A234;
  assign \new_[80132]_  = A266 & ~A265;
  assign \new_[80133]_  = \new_[80132]_  & \new_[80129]_ ;
  assign \new_[80134]_  = \new_[80133]_  & \new_[80126]_ ;
  assign \new_[80138]_  = A167 & ~A168;
  assign \new_[80139]_  = ~A169 & \new_[80138]_ ;
  assign \new_[80142]_  = A199 & A166;
  assign \new_[80145]_  = A201 & ~A200;
  assign \new_[80146]_  = \new_[80145]_  & \new_[80142]_ ;
  assign \new_[80147]_  = \new_[80146]_  & \new_[80139]_ ;
  assign \new_[80151]_  = ~A233 & A232;
  assign \new_[80152]_  = A202 & \new_[80151]_ ;
  assign \new_[80155]_  = A236 & A234;
  assign \new_[80158]_  = A299 & ~A298;
  assign \new_[80159]_  = \new_[80158]_  & \new_[80155]_ ;
  assign \new_[80160]_  = \new_[80159]_  & \new_[80152]_ ;
  assign \new_[80164]_  = A167 & ~A168;
  assign \new_[80165]_  = ~A169 & \new_[80164]_ ;
  assign \new_[80168]_  = A199 & A166;
  assign \new_[80171]_  = A201 & ~A200;
  assign \new_[80172]_  = \new_[80171]_  & \new_[80168]_ ;
  assign \new_[80173]_  = \new_[80172]_  & \new_[80165]_ ;
  assign \new_[80177]_  = ~A233 & A232;
  assign \new_[80178]_  = A202 & \new_[80177]_ ;
  assign \new_[80181]_  = A236 & A234;
  assign \new_[80184]_  = A266 & ~A265;
  assign \new_[80185]_  = \new_[80184]_  & \new_[80181]_ ;
  assign \new_[80186]_  = \new_[80185]_  & \new_[80178]_ ;
  assign \new_[80190]_  = A167 & ~A168;
  assign \new_[80191]_  = ~A169 & \new_[80190]_ ;
  assign \new_[80194]_  = A199 & A166;
  assign \new_[80197]_  = A201 & ~A200;
  assign \new_[80198]_  = \new_[80197]_  & \new_[80194]_ ;
  assign \new_[80199]_  = \new_[80198]_  & \new_[80191]_ ;
  assign \new_[80203]_  = ~A233 & ~A232;
  assign \new_[80204]_  = A202 & \new_[80203]_ ;
  assign \new_[80207]_  = A266 & A265;
  assign \new_[80210]_  = ~A300 & A298;
  assign \new_[80211]_  = \new_[80210]_  & \new_[80207]_ ;
  assign \new_[80212]_  = \new_[80211]_  & \new_[80204]_ ;
  assign \new_[80216]_  = A167 & ~A168;
  assign \new_[80217]_  = ~A169 & \new_[80216]_ ;
  assign \new_[80220]_  = A199 & A166;
  assign \new_[80223]_  = A201 & ~A200;
  assign \new_[80224]_  = \new_[80223]_  & \new_[80220]_ ;
  assign \new_[80225]_  = \new_[80224]_  & \new_[80217]_ ;
  assign \new_[80229]_  = ~A233 & ~A232;
  assign \new_[80230]_  = A202 & \new_[80229]_ ;
  assign \new_[80233]_  = A266 & A265;
  assign \new_[80236]_  = A299 & A298;
  assign \new_[80237]_  = \new_[80236]_  & \new_[80233]_ ;
  assign \new_[80238]_  = \new_[80237]_  & \new_[80230]_ ;
  assign \new_[80242]_  = A167 & ~A168;
  assign \new_[80243]_  = ~A169 & \new_[80242]_ ;
  assign \new_[80246]_  = A199 & A166;
  assign \new_[80249]_  = A201 & ~A200;
  assign \new_[80250]_  = \new_[80249]_  & \new_[80246]_ ;
  assign \new_[80251]_  = \new_[80250]_  & \new_[80243]_ ;
  assign \new_[80255]_  = ~A233 & ~A232;
  assign \new_[80256]_  = A202 & \new_[80255]_ ;
  assign \new_[80259]_  = A266 & A265;
  assign \new_[80262]_  = ~A299 & ~A298;
  assign \new_[80263]_  = \new_[80262]_  & \new_[80259]_ ;
  assign \new_[80264]_  = \new_[80263]_  & \new_[80256]_ ;
  assign \new_[80268]_  = A167 & ~A168;
  assign \new_[80269]_  = ~A169 & \new_[80268]_ ;
  assign \new_[80272]_  = A199 & A166;
  assign \new_[80275]_  = A201 & ~A200;
  assign \new_[80276]_  = \new_[80275]_  & \new_[80272]_ ;
  assign \new_[80277]_  = \new_[80276]_  & \new_[80269]_ ;
  assign \new_[80281]_  = ~A233 & ~A232;
  assign \new_[80282]_  = A202 & \new_[80281]_ ;
  assign \new_[80285]_  = ~A267 & ~A266;
  assign \new_[80288]_  = ~A300 & A298;
  assign \new_[80289]_  = \new_[80288]_  & \new_[80285]_ ;
  assign \new_[80290]_  = \new_[80289]_  & \new_[80282]_ ;
  assign \new_[80294]_  = A167 & ~A168;
  assign \new_[80295]_  = ~A169 & \new_[80294]_ ;
  assign \new_[80298]_  = A199 & A166;
  assign \new_[80301]_  = A201 & ~A200;
  assign \new_[80302]_  = \new_[80301]_  & \new_[80298]_ ;
  assign \new_[80303]_  = \new_[80302]_  & \new_[80295]_ ;
  assign \new_[80307]_  = ~A233 & ~A232;
  assign \new_[80308]_  = A202 & \new_[80307]_ ;
  assign \new_[80311]_  = ~A267 & ~A266;
  assign \new_[80314]_  = A299 & A298;
  assign \new_[80315]_  = \new_[80314]_  & \new_[80311]_ ;
  assign \new_[80316]_  = \new_[80315]_  & \new_[80308]_ ;
  assign \new_[80320]_  = A167 & ~A168;
  assign \new_[80321]_  = ~A169 & \new_[80320]_ ;
  assign \new_[80324]_  = A199 & A166;
  assign \new_[80327]_  = A201 & ~A200;
  assign \new_[80328]_  = \new_[80327]_  & \new_[80324]_ ;
  assign \new_[80329]_  = \new_[80328]_  & \new_[80321]_ ;
  assign \new_[80333]_  = ~A233 & ~A232;
  assign \new_[80334]_  = A202 & \new_[80333]_ ;
  assign \new_[80337]_  = ~A267 & ~A266;
  assign \new_[80340]_  = ~A299 & ~A298;
  assign \new_[80341]_  = \new_[80340]_  & \new_[80337]_ ;
  assign \new_[80342]_  = \new_[80341]_  & \new_[80334]_ ;
  assign \new_[80346]_  = A167 & ~A168;
  assign \new_[80347]_  = ~A169 & \new_[80346]_ ;
  assign \new_[80350]_  = A199 & A166;
  assign \new_[80353]_  = A201 & ~A200;
  assign \new_[80354]_  = \new_[80353]_  & \new_[80350]_ ;
  assign \new_[80355]_  = \new_[80354]_  & \new_[80347]_ ;
  assign \new_[80359]_  = ~A233 & ~A232;
  assign \new_[80360]_  = A202 & \new_[80359]_ ;
  assign \new_[80363]_  = ~A266 & ~A265;
  assign \new_[80366]_  = ~A300 & A298;
  assign \new_[80367]_  = \new_[80366]_  & \new_[80363]_ ;
  assign \new_[80368]_  = \new_[80367]_  & \new_[80360]_ ;
  assign \new_[80372]_  = A167 & ~A168;
  assign \new_[80373]_  = ~A169 & \new_[80372]_ ;
  assign \new_[80376]_  = A199 & A166;
  assign \new_[80379]_  = A201 & ~A200;
  assign \new_[80380]_  = \new_[80379]_  & \new_[80376]_ ;
  assign \new_[80381]_  = \new_[80380]_  & \new_[80373]_ ;
  assign \new_[80385]_  = ~A233 & ~A232;
  assign \new_[80386]_  = A202 & \new_[80385]_ ;
  assign \new_[80389]_  = ~A266 & ~A265;
  assign \new_[80392]_  = A299 & A298;
  assign \new_[80393]_  = \new_[80392]_  & \new_[80389]_ ;
  assign \new_[80394]_  = \new_[80393]_  & \new_[80386]_ ;
  assign \new_[80398]_  = A167 & ~A168;
  assign \new_[80399]_  = ~A169 & \new_[80398]_ ;
  assign \new_[80402]_  = A199 & A166;
  assign \new_[80405]_  = A201 & ~A200;
  assign \new_[80406]_  = \new_[80405]_  & \new_[80402]_ ;
  assign \new_[80407]_  = \new_[80406]_  & \new_[80399]_ ;
  assign \new_[80411]_  = ~A233 & ~A232;
  assign \new_[80412]_  = A202 & \new_[80411]_ ;
  assign \new_[80415]_  = ~A266 & ~A265;
  assign \new_[80418]_  = ~A299 & ~A298;
  assign \new_[80419]_  = \new_[80418]_  & \new_[80415]_ ;
  assign \new_[80420]_  = \new_[80419]_  & \new_[80412]_ ;
  assign \new_[80424]_  = A167 & ~A168;
  assign \new_[80425]_  = ~A169 & \new_[80424]_ ;
  assign \new_[80428]_  = A199 & A166;
  assign \new_[80431]_  = A201 & ~A200;
  assign \new_[80432]_  = \new_[80431]_  & \new_[80428]_ ;
  assign \new_[80433]_  = \new_[80432]_  & \new_[80425]_ ;
  assign \new_[80437]_  = A233 & A232;
  assign \new_[80438]_  = A203 & \new_[80437]_ ;
  assign \new_[80441]_  = ~A267 & A265;
  assign \new_[80444]_  = ~A300 & ~A299;
  assign \new_[80445]_  = \new_[80444]_  & \new_[80441]_ ;
  assign \new_[80446]_  = \new_[80445]_  & \new_[80438]_ ;
  assign \new_[80450]_  = A167 & ~A168;
  assign \new_[80451]_  = ~A169 & \new_[80450]_ ;
  assign \new_[80454]_  = A199 & A166;
  assign \new_[80457]_  = A201 & ~A200;
  assign \new_[80458]_  = \new_[80457]_  & \new_[80454]_ ;
  assign \new_[80459]_  = \new_[80458]_  & \new_[80451]_ ;
  assign \new_[80463]_  = A233 & A232;
  assign \new_[80464]_  = A203 & \new_[80463]_ ;
  assign \new_[80467]_  = ~A267 & A265;
  assign \new_[80470]_  = A299 & A298;
  assign \new_[80471]_  = \new_[80470]_  & \new_[80467]_ ;
  assign \new_[80472]_  = \new_[80471]_  & \new_[80464]_ ;
  assign \new_[80476]_  = A167 & ~A168;
  assign \new_[80477]_  = ~A169 & \new_[80476]_ ;
  assign \new_[80480]_  = A199 & A166;
  assign \new_[80483]_  = A201 & ~A200;
  assign \new_[80484]_  = \new_[80483]_  & \new_[80480]_ ;
  assign \new_[80485]_  = \new_[80484]_  & \new_[80477]_ ;
  assign \new_[80489]_  = A233 & A232;
  assign \new_[80490]_  = A203 & \new_[80489]_ ;
  assign \new_[80493]_  = ~A267 & A265;
  assign \new_[80496]_  = ~A299 & ~A298;
  assign \new_[80497]_  = \new_[80496]_  & \new_[80493]_ ;
  assign \new_[80498]_  = \new_[80497]_  & \new_[80490]_ ;
  assign \new_[80502]_  = A167 & ~A168;
  assign \new_[80503]_  = ~A169 & \new_[80502]_ ;
  assign \new_[80506]_  = A199 & A166;
  assign \new_[80509]_  = A201 & ~A200;
  assign \new_[80510]_  = \new_[80509]_  & \new_[80506]_ ;
  assign \new_[80511]_  = \new_[80510]_  & \new_[80503]_ ;
  assign \new_[80515]_  = A233 & A232;
  assign \new_[80516]_  = A203 & \new_[80515]_ ;
  assign \new_[80519]_  = A266 & A265;
  assign \new_[80522]_  = ~A300 & ~A299;
  assign \new_[80523]_  = \new_[80522]_  & \new_[80519]_ ;
  assign \new_[80524]_  = \new_[80523]_  & \new_[80516]_ ;
  assign \new_[80528]_  = A167 & ~A168;
  assign \new_[80529]_  = ~A169 & \new_[80528]_ ;
  assign \new_[80532]_  = A199 & A166;
  assign \new_[80535]_  = A201 & ~A200;
  assign \new_[80536]_  = \new_[80535]_  & \new_[80532]_ ;
  assign \new_[80537]_  = \new_[80536]_  & \new_[80529]_ ;
  assign \new_[80541]_  = A233 & A232;
  assign \new_[80542]_  = A203 & \new_[80541]_ ;
  assign \new_[80545]_  = A266 & A265;
  assign \new_[80548]_  = A299 & A298;
  assign \new_[80549]_  = \new_[80548]_  & \new_[80545]_ ;
  assign \new_[80550]_  = \new_[80549]_  & \new_[80542]_ ;
  assign \new_[80554]_  = A167 & ~A168;
  assign \new_[80555]_  = ~A169 & \new_[80554]_ ;
  assign \new_[80558]_  = A199 & A166;
  assign \new_[80561]_  = A201 & ~A200;
  assign \new_[80562]_  = \new_[80561]_  & \new_[80558]_ ;
  assign \new_[80563]_  = \new_[80562]_  & \new_[80555]_ ;
  assign \new_[80567]_  = A233 & A232;
  assign \new_[80568]_  = A203 & \new_[80567]_ ;
  assign \new_[80571]_  = A266 & A265;
  assign \new_[80574]_  = ~A299 & ~A298;
  assign \new_[80575]_  = \new_[80574]_  & \new_[80571]_ ;
  assign \new_[80576]_  = \new_[80575]_  & \new_[80568]_ ;
  assign \new_[80580]_  = A167 & ~A168;
  assign \new_[80581]_  = ~A169 & \new_[80580]_ ;
  assign \new_[80584]_  = A199 & A166;
  assign \new_[80587]_  = A201 & ~A200;
  assign \new_[80588]_  = \new_[80587]_  & \new_[80584]_ ;
  assign \new_[80589]_  = \new_[80588]_  & \new_[80581]_ ;
  assign \new_[80593]_  = A233 & A232;
  assign \new_[80594]_  = A203 & \new_[80593]_ ;
  assign \new_[80597]_  = ~A266 & ~A265;
  assign \new_[80600]_  = ~A300 & ~A299;
  assign \new_[80601]_  = \new_[80600]_  & \new_[80597]_ ;
  assign \new_[80602]_  = \new_[80601]_  & \new_[80594]_ ;
  assign \new_[80606]_  = A167 & ~A168;
  assign \new_[80607]_  = ~A169 & \new_[80606]_ ;
  assign \new_[80610]_  = A199 & A166;
  assign \new_[80613]_  = A201 & ~A200;
  assign \new_[80614]_  = \new_[80613]_  & \new_[80610]_ ;
  assign \new_[80615]_  = \new_[80614]_  & \new_[80607]_ ;
  assign \new_[80619]_  = A233 & A232;
  assign \new_[80620]_  = A203 & \new_[80619]_ ;
  assign \new_[80623]_  = ~A266 & ~A265;
  assign \new_[80626]_  = A299 & A298;
  assign \new_[80627]_  = \new_[80626]_  & \new_[80623]_ ;
  assign \new_[80628]_  = \new_[80627]_  & \new_[80620]_ ;
  assign \new_[80632]_  = A167 & ~A168;
  assign \new_[80633]_  = ~A169 & \new_[80632]_ ;
  assign \new_[80636]_  = A199 & A166;
  assign \new_[80639]_  = A201 & ~A200;
  assign \new_[80640]_  = \new_[80639]_  & \new_[80636]_ ;
  assign \new_[80641]_  = \new_[80640]_  & \new_[80633]_ ;
  assign \new_[80645]_  = A233 & A232;
  assign \new_[80646]_  = A203 & \new_[80645]_ ;
  assign \new_[80649]_  = ~A266 & ~A265;
  assign \new_[80652]_  = ~A299 & ~A298;
  assign \new_[80653]_  = \new_[80652]_  & \new_[80649]_ ;
  assign \new_[80654]_  = \new_[80653]_  & \new_[80646]_ ;
  assign \new_[80658]_  = A167 & ~A168;
  assign \new_[80659]_  = ~A169 & \new_[80658]_ ;
  assign \new_[80662]_  = A199 & A166;
  assign \new_[80665]_  = A201 & ~A200;
  assign \new_[80666]_  = \new_[80665]_  & \new_[80662]_ ;
  assign \new_[80667]_  = \new_[80666]_  & \new_[80659]_ ;
  assign \new_[80671]_  = A233 & ~A232;
  assign \new_[80672]_  = A203 & \new_[80671]_ ;
  assign \new_[80675]_  = ~A299 & A298;
  assign \new_[80678]_  = A301 & A300;
  assign \new_[80679]_  = \new_[80678]_  & \new_[80675]_ ;
  assign \new_[80680]_  = \new_[80679]_  & \new_[80672]_ ;
  assign \new_[80684]_  = A167 & ~A168;
  assign \new_[80685]_  = ~A169 & \new_[80684]_ ;
  assign \new_[80688]_  = A199 & A166;
  assign \new_[80691]_  = A201 & ~A200;
  assign \new_[80692]_  = \new_[80691]_  & \new_[80688]_ ;
  assign \new_[80693]_  = \new_[80692]_  & \new_[80685]_ ;
  assign \new_[80697]_  = A233 & ~A232;
  assign \new_[80698]_  = A203 & \new_[80697]_ ;
  assign \new_[80701]_  = ~A299 & A298;
  assign \new_[80704]_  = A302 & A300;
  assign \new_[80705]_  = \new_[80704]_  & \new_[80701]_ ;
  assign \new_[80706]_  = \new_[80705]_  & \new_[80698]_ ;
  assign \new_[80710]_  = A167 & ~A168;
  assign \new_[80711]_  = ~A169 & \new_[80710]_ ;
  assign \new_[80714]_  = A199 & A166;
  assign \new_[80717]_  = A201 & ~A200;
  assign \new_[80718]_  = \new_[80717]_  & \new_[80714]_ ;
  assign \new_[80719]_  = \new_[80718]_  & \new_[80711]_ ;
  assign \new_[80723]_  = A233 & ~A232;
  assign \new_[80724]_  = A203 & \new_[80723]_ ;
  assign \new_[80727]_  = ~A266 & A265;
  assign \new_[80730]_  = A268 & A267;
  assign \new_[80731]_  = \new_[80730]_  & \new_[80727]_ ;
  assign \new_[80732]_  = \new_[80731]_  & \new_[80724]_ ;
  assign \new_[80736]_  = A167 & ~A168;
  assign \new_[80737]_  = ~A169 & \new_[80736]_ ;
  assign \new_[80740]_  = A199 & A166;
  assign \new_[80743]_  = A201 & ~A200;
  assign \new_[80744]_  = \new_[80743]_  & \new_[80740]_ ;
  assign \new_[80745]_  = \new_[80744]_  & \new_[80737]_ ;
  assign \new_[80749]_  = A233 & ~A232;
  assign \new_[80750]_  = A203 & \new_[80749]_ ;
  assign \new_[80753]_  = ~A266 & A265;
  assign \new_[80756]_  = A269 & A267;
  assign \new_[80757]_  = \new_[80756]_  & \new_[80753]_ ;
  assign \new_[80758]_  = \new_[80757]_  & \new_[80750]_ ;
  assign \new_[80762]_  = A167 & ~A168;
  assign \new_[80763]_  = ~A169 & \new_[80762]_ ;
  assign \new_[80766]_  = A199 & A166;
  assign \new_[80769]_  = A201 & ~A200;
  assign \new_[80770]_  = \new_[80769]_  & \new_[80766]_ ;
  assign \new_[80771]_  = \new_[80770]_  & \new_[80763]_ ;
  assign \new_[80775]_  = ~A234 & ~A233;
  assign \new_[80776]_  = A203 & \new_[80775]_ ;
  assign \new_[80779]_  = A266 & A265;
  assign \new_[80782]_  = ~A300 & A298;
  assign \new_[80783]_  = \new_[80782]_  & \new_[80779]_ ;
  assign \new_[80784]_  = \new_[80783]_  & \new_[80776]_ ;
  assign \new_[80788]_  = A167 & ~A168;
  assign \new_[80789]_  = ~A169 & \new_[80788]_ ;
  assign \new_[80792]_  = A199 & A166;
  assign \new_[80795]_  = A201 & ~A200;
  assign \new_[80796]_  = \new_[80795]_  & \new_[80792]_ ;
  assign \new_[80797]_  = \new_[80796]_  & \new_[80789]_ ;
  assign \new_[80801]_  = ~A234 & ~A233;
  assign \new_[80802]_  = A203 & \new_[80801]_ ;
  assign \new_[80805]_  = A266 & A265;
  assign \new_[80808]_  = A299 & A298;
  assign \new_[80809]_  = \new_[80808]_  & \new_[80805]_ ;
  assign \new_[80810]_  = \new_[80809]_  & \new_[80802]_ ;
  assign \new_[80814]_  = A167 & ~A168;
  assign \new_[80815]_  = ~A169 & \new_[80814]_ ;
  assign \new_[80818]_  = A199 & A166;
  assign \new_[80821]_  = A201 & ~A200;
  assign \new_[80822]_  = \new_[80821]_  & \new_[80818]_ ;
  assign \new_[80823]_  = \new_[80822]_  & \new_[80815]_ ;
  assign \new_[80827]_  = ~A234 & ~A233;
  assign \new_[80828]_  = A203 & \new_[80827]_ ;
  assign \new_[80831]_  = A266 & A265;
  assign \new_[80834]_  = ~A299 & ~A298;
  assign \new_[80835]_  = \new_[80834]_  & \new_[80831]_ ;
  assign \new_[80836]_  = \new_[80835]_  & \new_[80828]_ ;
  assign \new_[80840]_  = A167 & ~A168;
  assign \new_[80841]_  = ~A169 & \new_[80840]_ ;
  assign \new_[80844]_  = A199 & A166;
  assign \new_[80847]_  = A201 & ~A200;
  assign \new_[80848]_  = \new_[80847]_  & \new_[80844]_ ;
  assign \new_[80849]_  = \new_[80848]_  & \new_[80841]_ ;
  assign \new_[80853]_  = ~A234 & ~A233;
  assign \new_[80854]_  = A203 & \new_[80853]_ ;
  assign \new_[80857]_  = ~A267 & ~A266;
  assign \new_[80860]_  = ~A300 & A298;
  assign \new_[80861]_  = \new_[80860]_  & \new_[80857]_ ;
  assign \new_[80862]_  = \new_[80861]_  & \new_[80854]_ ;
  assign \new_[80866]_  = A167 & ~A168;
  assign \new_[80867]_  = ~A169 & \new_[80866]_ ;
  assign \new_[80870]_  = A199 & A166;
  assign \new_[80873]_  = A201 & ~A200;
  assign \new_[80874]_  = \new_[80873]_  & \new_[80870]_ ;
  assign \new_[80875]_  = \new_[80874]_  & \new_[80867]_ ;
  assign \new_[80879]_  = ~A234 & ~A233;
  assign \new_[80880]_  = A203 & \new_[80879]_ ;
  assign \new_[80883]_  = ~A267 & ~A266;
  assign \new_[80886]_  = A299 & A298;
  assign \new_[80887]_  = \new_[80886]_  & \new_[80883]_ ;
  assign \new_[80888]_  = \new_[80887]_  & \new_[80880]_ ;
  assign \new_[80892]_  = A167 & ~A168;
  assign \new_[80893]_  = ~A169 & \new_[80892]_ ;
  assign \new_[80896]_  = A199 & A166;
  assign \new_[80899]_  = A201 & ~A200;
  assign \new_[80900]_  = \new_[80899]_  & \new_[80896]_ ;
  assign \new_[80901]_  = \new_[80900]_  & \new_[80893]_ ;
  assign \new_[80905]_  = ~A234 & ~A233;
  assign \new_[80906]_  = A203 & \new_[80905]_ ;
  assign \new_[80909]_  = ~A267 & ~A266;
  assign \new_[80912]_  = ~A299 & ~A298;
  assign \new_[80913]_  = \new_[80912]_  & \new_[80909]_ ;
  assign \new_[80914]_  = \new_[80913]_  & \new_[80906]_ ;
  assign \new_[80918]_  = A167 & ~A168;
  assign \new_[80919]_  = ~A169 & \new_[80918]_ ;
  assign \new_[80922]_  = A199 & A166;
  assign \new_[80925]_  = A201 & ~A200;
  assign \new_[80926]_  = \new_[80925]_  & \new_[80922]_ ;
  assign \new_[80927]_  = \new_[80926]_  & \new_[80919]_ ;
  assign \new_[80931]_  = ~A234 & ~A233;
  assign \new_[80932]_  = A203 & \new_[80931]_ ;
  assign \new_[80935]_  = ~A266 & ~A265;
  assign \new_[80938]_  = ~A300 & A298;
  assign \new_[80939]_  = \new_[80938]_  & \new_[80935]_ ;
  assign \new_[80940]_  = \new_[80939]_  & \new_[80932]_ ;
  assign \new_[80944]_  = A167 & ~A168;
  assign \new_[80945]_  = ~A169 & \new_[80944]_ ;
  assign \new_[80948]_  = A199 & A166;
  assign \new_[80951]_  = A201 & ~A200;
  assign \new_[80952]_  = \new_[80951]_  & \new_[80948]_ ;
  assign \new_[80953]_  = \new_[80952]_  & \new_[80945]_ ;
  assign \new_[80957]_  = ~A234 & ~A233;
  assign \new_[80958]_  = A203 & \new_[80957]_ ;
  assign \new_[80961]_  = ~A266 & ~A265;
  assign \new_[80964]_  = A299 & A298;
  assign \new_[80965]_  = \new_[80964]_  & \new_[80961]_ ;
  assign \new_[80966]_  = \new_[80965]_  & \new_[80958]_ ;
  assign \new_[80970]_  = A167 & ~A168;
  assign \new_[80971]_  = ~A169 & \new_[80970]_ ;
  assign \new_[80974]_  = A199 & A166;
  assign \new_[80977]_  = A201 & ~A200;
  assign \new_[80978]_  = \new_[80977]_  & \new_[80974]_ ;
  assign \new_[80979]_  = \new_[80978]_  & \new_[80971]_ ;
  assign \new_[80983]_  = ~A234 & ~A233;
  assign \new_[80984]_  = A203 & \new_[80983]_ ;
  assign \new_[80987]_  = ~A266 & ~A265;
  assign \new_[80990]_  = ~A299 & ~A298;
  assign \new_[80991]_  = \new_[80990]_  & \new_[80987]_ ;
  assign \new_[80992]_  = \new_[80991]_  & \new_[80984]_ ;
  assign \new_[80996]_  = A167 & ~A168;
  assign \new_[80997]_  = ~A169 & \new_[80996]_ ;
  assign \new_[81000]_  = A199 & A166;
  assign \new_[81003]_  = A201 & ~A200;
  assign \new_[81004]_  = \new_[81003]_  & \new_[81000]_ ;
  assign \new_[81005]_  = \new_[81004]_  & \new_[80997]_ ;
  assign \new_[81009]_  = ~A233 & A232;
  assign \new_[81010]_  = A203 & \new_[81009]_ ;
  assign \new_[81013]_  = A235 & A234;
  assign \new_[81016]_  = A299 & ~A298;
  assign \new_[81017]_  = \new_[81016]_  & \new_[81013]_ ;
  assign \new_[81018]_  = \new_[81017]_  & \new_[81010]_ ;
  assign \new_[81022]_  = A167 & ~A168;
  assign \new_[81023]_  = ~A169 & \new_[81022]_ ;
  assign \new_[81026]_  = A199 & A166;
  assign \new_[81029]_  = A201 & ~A200;
  assign \new_[81030]_  = \new_[81029]_  & \new_[81026]_ ;
  assign \new_[81031]_  = \new_[81030]_  & \new_[81023]_ ;
  assign \new_[81035]_  = ~A233 & A232;
  assign \new_[81036]_  = A203 & \new_[81035]_ ;
  assign \new_[81039]_  = A235 & A234;
  assign \new_[81042]_  = A266 & ~A265;
  assign \new_[81043]_  = \new_[81042]_  & \new_[81039]_ ;
  assign \new_[81044]_  = \new_[81043]_  & \new_[81036]_ ;
  assign \new_[81048]_  = A167 & ~A168;
  assign \new_[81049]_  = ~A169 & \new_[81048]_ ;
  assign \new_[81052]_  = A199 & A166;
  assign \new_[81055]_  = A201 & ~A200;
  assign \new_[81056]_  = \new_[81055]_  & \new_[81052]_ ;
  assign \new_[81057]_  = \new_[81056]_  & \new_[81049]_ ;
  assign \new_[81061]_  = ~A233 & A232;
  assign \new_[81062]_  = A203 & \new_[81061]_ ;
  assign \new_[81065]_  = A236 & A234;
  assign \new_[81068]_  = A299 & ~A298;
  assign \new_[81069]_  = \new_[81068]_  & \new_[81065]_ ;
  assign \new_[81070]_  = \new_[81069]_  & \new_[81062]_ ;
  assign \new_[81074]_  = A167 & ~A168;
  assign \new_[81075]_  = ~A169 & \new_[81074]_ ;
  assign \new_[81078]_  = A199 & A166;
  assign \new_[81081]_  = A201 & ~A200;
  assign \new_[81082]_  = \new_[81081]_  & \new_[81078]_ ;
  assign \new_[81083]_  = \new_[81082]_  & \new_[81075]_ ;
  assign \new_[81087]_  = ~A233 & A232;
  assign \new_[81088]_  = A203 & \new_[81087]_ ;
  assign \new_[81091]_  = A236 & A234;
  assign \new_[81094]_  = A266 & ~A265;
  assign \new_[81095]_  = \new_[81094]_  & \new_[81091]_ ;
  assign \new_[81096]_  = \new_[81095]_  & \new_[81088]_ ;
  assign \new_[81100]_  = A167 & ~A168;
  assign \new_[81101]_  = ~A169 & \new_[81100]_ ;
  assign \new_[81104]_  = A199 & A166;
  assign \new_[81107]_  = A201 & ~A200;
  assign \new_[81108]_  = \new_[81107]_  & \new_[81104]_ ;
  assign \new_[81109]_  = \new_[81108]_  & \new_[81101]_ ;
  assign \new_[81113]_  = ~A233 & ~A232;
  assign \new_[81114]_  = A203 & \new_[81113]_ ;
  assign \new_[81117]_  = A266 & A265;
  assign \new_[81120]_  = ~A300 & A298;
  assign \new_[81121]_  = \new_[81120]_  & \new_[81117]_ ;
  assign \new_[81122]_  = \new_[81121]_  & \new_[81114]_ ;
  assign \new_[81126]_  = A167 & ~A168;
  assign \new_[81127]_  = ~A169 & \new_[81126]_ ;
  assign \new_[81130]_  = A199 & A166;
  assign \new_[81133]_  = A201 & ~A200;
  assign \new_[81134]_  = \new_[81133]_  & \new_[81130]_ ;
  assign \new_[81135]_  = \new_[81134]_  & \new_[81127]_ ;
  assign \new_[81139]_  = ~A233 & ~A232;
  assign \new_[81140]_  = A203 & \new_[81139]_ ;
  assign \new_[81143]_  = A266 & A265;
  assign \new_[81146]_  = A299 & A298;
  assign \new_[81147]_  = \new_[81146]_  & \new_[81143]_ ;
  assign \new_[81148]_  = \new_[81147]_  & \new_[81140]_ ;
  assign \new_[81152]_  = A167 & ~A168;
  assign \new_[81153]_  = ~A169 & \new_[81152]_ ;
  assign \new_[81156]_  = A199 & A166;
  assign \new_[81159]_  = A201 & ~A200;
  assign \new_[81160]_  = \new_[81159]_  & \new_[81156]_ ;
  assign \new_[81161]_  = \new_[81160]_  & \new_[81153]_ ;
  assign \new_[81165]_  = ~A233 & ~A232;
  assign \new_[81166]_  = A203 & \new_[81165]_ ;
  assign \new_[81169]_  = A266 & A265;
  assign \new_[81172]_  = ~A299 & ~A298;
  assign \new_[81173]_  = \new_[81172]_  & \new_[81169]_ ;
  assign \new_[81174]_  = \new_[81173]_  & \new_[81166]_ ;
  assign \new_[81178]_  = A167 & ~A168;
  assign \new_[81179]_  = ~A169 & \new_[81178]_ ;
  assign \new_[81182]_  = A199 & A166;
  assign \new_[81185]_  = A201 & ~A200;
  assign \new_[81186]_  = \new_[81185]_  & \new_[81182]_ ;
  assign \new_[81187]_  = \new_[81186]_  & \new_[81179]_ ;
  assign \new_[81191]_  = ~A233 & ~A232;
  assign \new_[81192]_  = A203 & \new_[81191]_ ;
  assign \new_[81195]_  = ~A267 & ~A266;
  assign \new_[81198]_  = ~A300 & A298;
  assign \new_[81199]_  = \new_[81198]_  & \new_[81195]_ ;
  assign \new_[81200]_  = \new_[81199]_  & \new_[81192]_ ;
  assign \new_[81204]_  = A167 & ~A168;
  assign \new_[81205]_  = ~A169 & \new_[81204]_ ;
  assign \new_[81208]_  = A199 & A166;
  assign \new_[81211]_  = A201 & ~A200;
  assign \new_[81212]_  = \new_[81211]_  & \new_[81208]_ ;
  assign \new_[81213]_  = \new_[81212]_  & \new_[81205]_ ;
  assign \new_[81217]_  = ~A233 & ~A232;
  assign \new_[81218]_  = A203 & \new_[81217]_ ;
  assign \new_[81221]_  = ~A267 & ~A266;
  assign \new_[81224]_  = A299 & A298;
  assign \new_[81225]_  = \new_[81224]_  & \new_[81221]_ ;
  assign \new_[81226]_  = \new_[81225]_  & \new_[81218]_ ;
  assign \new_[81230]_  = A167 & ~A168;
  assign \new_[81231]_  = ~A169 & \new_[81230]_ ;
  assign \new_[81234]_  = A199 & A166;
  assign \new_[81237]_  = A201 & ~A200;
  assign \new_[81238]_  = \new_[81237]_  & \new_[81234]_ ;
  assign \new_[81239]_  = \new_[81238]_  & \new_[81231]_ ;
  assign \new_[81243]_  = ~A233 & ~A232;
  assign \new_[81244]_  = A203 & \new_[81243]_ ;
  assign \new_[81247]_  = ~A267 & ~A266;
  assign \new_[81250]_  = ~A299 & ~A298;
  assign \new_[81251]_  = \new_[81250]_  & \new_[81247]_ ;
  assign \new_[81252]_  = \new_[81251]_  & \new_[81244]_ ;
  assign \new_[81256]_  = A167 & ~A168;
  assign \new_[81257]_  = ~A169 & \new_[81256]_ ;
  assign \new_[81260]_  = A199 & A166;
  assign \new_[81263]_  = A201 & ~A200;
  assign \new_[81264]_  = \new_[81263]_  & \new_[81260]_ ;
  assign \new_[81265]_  = \new_[81264]_  & \new_[81257]_ ;
  assign \new_[81269]_  = ~A233 & ~A232;
  assign \new_[81270]_  = A203 & \new_[81269]_ ;
  assign \new_[81273]_  = ~A266 & ~A265;
  assign \new_[81276]_  = ~A300 & A298;
  assign \new_[81277]_  = \new_[81276]_  & \new_[81273]_ ;
  assign \new_[81278]_  = \new_[81277]_  & \new_[81270]_ ;
  assign \new_[81282]_  = A167 & ~A168;
  assign \new_[81283]_  = ~A169 & \new_[81282]_ ;
  assign \new_[81286]_  = A199 & A166;
  assign \new_[81289]_  = A201 & ~A200;
  assign \new_[81290]_  = \new_[81289]_  & \new_[81286]_ ;
  assign \new_[81291]_  = \new_[81290]_  & \new_[81283]_ ;
  assign \new_[81295]_  = ~A233 & ~A232;
  assign \new_[81296]_  = A203 & \new_[81295]_ ;
  assign \new_[81299]_  = ~A266 & ~A265;
  assign \new_[81302]_  = A299 & A298;
  assign \new_[81303]_  = \new_[81302]_  & \new_[81299]_ ;
  assign \new_[81304]_  = \new_[81303]_  & \new_[81296]_ ;
  assign \new_[81308]_  = A167 & ~A168;
  assign \new_[81309]_  = ~A169 & \new_[81308]_ ;
  assign \new_[81312]_  = A199 & A166;
  assign \new_[81315]_  = A201 & ~A200;
  assign \new_[81316]_  = \new_[81315]_  & \new_[81312]_ ;
  assign \new_[81317]_  = \new_[81316]_  & \new_[81309]_ ;
  assign \new_[81321]_  = ~A233 & ~A232;
  assign \new_[81322]_  = A203 & \new_[81321]_ ;
  assign \new_[81325]_  = ~A266 & ~A265;
  assign \new_[81328]_  = ~A299 & ~A298;
  assign \new_[81329]_  = \new_[81328]_  & \new_[81325]_ ;
  assign \new_[81330]_  = \new_[81329]_  & \new_[81322]_ ;
  assign \new_[81334]_  = A167 & ~A169;
  assign \new_[81335]_  = A170 & \new_[81334]_ ;
  assign \new_[81338]_  = A199 & ~A166;
  assign \new_[81341]_  = A232 & A200;
  assign \new_[81342]_  = \new_[81341]_  & \new_[81338]_ ;
  assign \new_[81343]_  = \new_[81342]_  & \new_[81335]_ ;
  assign \new_[81347]_  = ~A268 & A265;
  assign \new_[81348]_  = A233 & \new_[81347]_ ;
  assign \new_[81351]_  = ~A299 & ~A269;
  assign \new_[81354]_  = ~A302 & ~A301;
  assign \new_[81355]_  = \new_[81354]_  & \new_[81351]_ ;
  assign \new_[81356]_  = \new_[81355]_  & \new_[81348]_ ;
  assign \new_[81360]_  = A167 & ~A169;
  assign \new_[81361]_  = A170 & \new_[81360]_ ;
  assign \new_[81364]_  = A199 & ~A166;
  assign \new_[81367]_  = ~A233 & A200;
  assign \new_[81368]_  = \new_[81367]_  & \new_[81364]_ ;
  assign \new_[81369]_  = \new_[81368]_  & \new_[81361]_ ;
  assign \new_[81373]_  = A265 & ~A236;
  assign \new_[81374]_  = ~A235 & \new_[81373]_ ;
  assign \new_[81377]_  = A298 & A266;
  assign \new_[81380]_  = ~A302 & ~A301;
  assign \new_[81381]_  = \new_[81380]_  & \new_[81377]_ ;
  assign \new_[81382]_  = \new_[81381]_  & \new_[81374]_ ;
  assign \new_[81386]_  = A167 & ~A169;
  assign \new_[81387]_  = A170 & \new_[81386]_ ;
  assign \new_[81390]_  = A199 & ~A166;
  assign \new_[81393]_  = ~A233 & A200;
  assign \new_[81394]_  = \new_[81393]_  & \new_[81390]_ ;
  assign \new_[81395]_  = \new_[81394]_  & \new_[81387]_ ;
  assign \new_[81399]_  = ~A266 & ~A236;
  assign \new_[81400]_  = ~A235 & \new_[81399]_ ;
  assign \new_[81403]_  = ~A269 & ~A268;
  assign \new_[81406]_  = ~A300 & A298;
  assign \new_[81407]_  = \new_[81406]_  & \new_[81403]_ ;
  assign \new_[81408]_  = \new_[81407]_  & \new_[81400]_ ;
  assign \new_[81412]_  = A167 & ~A169;
  assign \new_[81413]_  = A170 & \new_[81412]_ ;
  assign \new_[81416]_  = A199 & ~A166;
  assign \new_[81419]_  = ~A233 & A200;
  assign \new_[81420]_  = \new_[81419]_  & \new_[81416]_ ;
  assign \new_[81421]_  = \new_[81420]_  & \new_[81413]_ ;
  assign \new_[81425]_  = ~A266 & ~A236;
  assign \new_[81426]_  = ~A235 & \new_[81425]_ ;
  assign \new_[81429]_  = ~A269 & ~A268;
  assign \new_[81432]_  = A299 & A298;
  assign \new_[81433]_  = \new_[81432]_  & \new_[81429]_ ;
  assign \new_[81434]_  = \new_[81433]_  & \new_[81426]_ ;
  assign \new_[81438]_  = A167 & ~A169;
  assign \new_[81439]_  = A170 & \new_[81438]_ ;
  assign \new_[81442]_  = A199 & ~A166;
  assign \new_[81445]_  = ~A233 & A200;
  assign \new_[81446]_  = \new_[81445]_  & \new_[81442]_ ;
  assign \new_[81447]_  = \new_[81446]_  & \new_[81439]_ ;
  assign \new_[81451]_  = ~A266 & ~A236;
  assign \new_[81452]_  = ~A235 & \new_[81451]_ ;
  assign \new_[81455]_  = ~A269 & ~A268;
  assign \new_[81458]_  = ~A299 & ~A298;
  assign \new_[81459]_  = \new_[81458]_  & \new_[81455]_ ;
  assign \new_[81460]_  = \new_[81459]_  & \new_[81452]_ ;
  assign \new_[81464]_  = A167 & ~A169;
  assign \new_[81465]_  = A170 & \new_[81464]_ ;
  assign \new_[81468]_  = A199 & ~A166;
  assign \new_[81471]_  = ~A233 & A200;
  assign \new_[81472]_  = \new_[81471]_  & \new_[81468]_ ;
  assign \new_[81473]_  = \new_[81472]_  & \new_[81465]_ ;
  assign \new_[81477]_  = ~A266 & ~A236;
  assign \new_[81478]_  = ~A235 & \new_[81477]_ ;
  assign \new_[81481]_  = A298 & ~A267;
  assign \new_[81484]_  = ~A302 & ~A301;
  assign \new_[81485]_  = \new_[81484]_  & \new_[81481]_ ;
  assign \new_[81486]_  = \new_[81485]_  & \new_[81478]_ ;
  assign \new_[81490]_  = A167 & ~A169;
  assign \new_[81491]_  = A170 & \new_[81490]_ ;
  assign \new_[81494]_  = A199 & ~A166;
  assign \new_[81497]_  = ~A233 & A200;
  assign \new_[81498]_  = \new_[81497]_  & \new_[81494]_ ;
  assign \new_[81499]_  = \new_[81498]_  & \new_[81491]_ ;
  assign \new_[81503]_  = ~A265 & ~A236;
  assign \new_[81504]_  = ~A235 & \new_[81503]_ ;
  assign \new_[81507]_  = A298 & ~A266;
  assign \new_[81510]_  = ~A302 & ~A301;
  assign \new_[81511]_  = \new_[81510]_  & \new_[81507]_ ;
  assign \new_[81512]_  = \new_[81511]_  & \new_[81504]_ ;
  assign \new_[81516]_  = A167 & ~A169;
  assign \new_[81517]_  = A170 & \new_[81516]_ ;
  assign \new_[81520]_  = A199 & ~A166;
  assign \new_[81523]_  = ~A233 & A200;
  assign \new_[81524]_  = \new_[81523]_  & \new_[81520]_ ;
  assign \new_[81525]_  = \new_[81524]_  & \new_[81517]_ ;
  assign \new_[81529]_  = ~A268 & ~A266;
  assign \new_[81530]_  = ~A234 & \new_[81529]_ ;
  assign \new_[81533]_  = A298 & ~A269;
  assign \new_[81536]_  = ~A302 & ~A301;
  assign \new_[81537]_  = \new_[81536]_  & \new_[81533]_ ;
  assign \new_[81538]_  = \new_[81537]_  & \new_[81530]_ ;
  assign \new_[81542]_  = A167 & ~A169;
  assign \new_[81543]_  = A170 & \new_[81542]_ ;
  assign \new_[81546]_  = A199 & ~A166;
  assign \new_[81549]_  = A232 & A200;
  assign \new_[81550]_  = \new_[81549]_  & \new_[81546]_ ;
  assign \new_[81551]_  = \new_[81550]_  & \new_[81543]_ ;
  assign \new_[81555]_  = A235 & A234;
  assign \new_[81556]_  = ~A233 & \new_[81555]_ ;
  assign \new_[81559]_  = ~A299 & A298;
  assign \new_[81562]_  = A301 & A300;
  assign \new_[81563]_  = \new_[81562]_  & \new_[81559]_ ;
  assign \new_[81564]_  = \new_[81563]_  & \new_[81556]_ ;
  assign \new_[81568]_  = A167 & ~A169;
  assign \new_[81569]_  = A170 & \new_[81568]_ ;
  assign \new_[81572]_  = A199 & ~A166;
  assign \new_[81575]_  = A232 & A200;
  assign \new_[81576]_  = \new_[81575]_  & \new_[81572]_ ;
  assign \new_[81577]_  = \new_[81576]_  & \new_[81569]_ ;
  assign \new_[81581]_  = A235 & A234;
  assign \new_[81582]_  = ~A233 & \new_[81581]_ ;
  assign \new_[81585]_  = ~A299 & A298;
  assign \new_[81588]_  = A302 & A300;
  assign \new_[81589]_  = \new_[81588]_  & \new_[81585]_ ;
  assign \new_[81590]_  = \new_[81589]_  & \new_[81582]_ ;
  assign \new_[81594]_  = A167 & ~A169;
  assign \new_[81595]_  = A170 & \new_[81594]_ ;
  assign \new_[81598]_  = A199 & ~A166;
  assign \new_[81601]_  = A232 & A200;
  assign \new_[81602]_  = \new_[81601]_  & \new_[81598]_ ;
  assign \new_[81603]_  = \new_[81602]_  & \new_[81595]_ ;
  assign \new_[81607]_  = A235 & A234;
  assign \new_[81608]_  = ~A233 & \new_[81607]_ ;
  assign \new_[81611]_  = ~A266 & A265;
  assign \new_[81614]_  = A268 & A267;
  assign \new_[81615]_  = \new_[81614]_  & \new_[81611]_ ;
  assign \new_[81616]_  = \new_[81615]_  & \new_[81608]_ ;
  assign \new_[81620]_  = A167 & ~A169;
  assign \new_[81621]_  = A170 & \new_[81620]_ ;
  assign \new_[81624]_  = A199 & ~A166;
  assign \new_[81627]_  = A232 & A200;
  assign \new_[81628]_  = \new_[81627]_  & \new_[81624]_ ;
  assign \new_[81629]_  = \new_[81628]_  & \new_[81621]_ ;
  assign \new_[81633]_  = A235 & A234;
  assign \new_[81634]_  = ~A233 & \new_[81633]_ ;
  assign \new_[81637]_  = ~A266 & A265;
  assign \new_[81640]_  = A269 & A267;
  assign \new_[81641]_  = \new_[81640]_  & \new_[81637]_ ;
  assign \new_[81642]_  = \new_[81641]_  & \new_[81634]_ ;
  assign \new_[81646]_  = A167 & ~A169;
  assign \new_[81647]_  = A170 & \new_[81646]_ ;
  assign \new_[81650]_  = A199 & ~A166;
  assign \new_[81653]_  = A232 & A200;
  assign \new_[81654]_  = \new_[81653]_  & \new_[81650]_ ;
  assign \new_[81655]_  = \new_[81654]_  & \new_[81647]_ ;
  assign \new_[81659]_  = A236 & A234;
  assign \new_[81660]_  = ~A233 & \new_[81659]_ ;
  assign \new_[81663]_  = ~A299 & A298;
  assign \new_[81666]_  = A301 & A300;
  assign \new_[81667]_  = \new_[81666]_  & \new_[81663]_ ;
  assign \new_[81668]_  = \new_[81667]_  & \new_[81660]_ ;
  assign \new_[81672]_  = A167 & ~A169;
  assign \new_[81673]_  = A170 & \new_[81672]_ ;
  assign \new_[81676]_  = A199 & ~A166;
  assign \new_[81679]_  = A232 & A200;
  assign \new_[81680]_  = \new_[81679]_  & \new_[81676]_ ;
  assign \new_[81681]_  = \new_[81680]_  & \new_[81673]_ ;
  assign \new_[81685]_  = A236 & A234;
  assign \new_[81686]_  = ~A233 & \new_[81685]_ ;
  assign \new_[81689]_  = ~A299 & A298;
  assign \new_[81692]_  = A302 & A300;
  assign \new_[81693]_  = \new_[81692]_  & \new_[81689]_ ;
  assign \new_[81694]_  = \new_[81693]_  & \new_[81686]_ ;
  assign \new_[81698]_  = A167 & ~A169;
  assign \new_[81699]_  = A170 & \new_[81698]_ ;
  assign \new_[81702]_  = A199 & ~A166;
  assign \new_[81705]_  = A232 & A200;
  assign \new_[81706]_  = \new_[81705]_  & \new_[81702]_ ;
  assign \new_[81707]_  = \new_[81706]_  & \new_[81699]_ ;
  assign \new_[81711]_  = A236 & A234;
  assign \new_[81712]_  = ~A233 & \new_[81711]_ ;
  assign \new_[81715]_  = ~A266 & A265;
  assign \new_[81718]_  = A268 & A267;
  assign \new_[81719]_  = \new_[81718]_  & \new_[81715]_ ;
  assign \new_[81720]_  = \new_[81719]_  & \new_[81712]_ ;
  assign \new_[81724]_  = A167 & ~A169;
  assign \new_[81725]_  = A170 & \new_[81724]_ ;
  assign \new_[81728]_  = A199 & ~A166;
  assign \new_[81731]_  = A232 & A200;
  assign \new_[81732]_  = \new_[81731]_  & \new_[81728]_ ;
  assign \new_[81733]_  = \new_[81732]_  & \new_[81725]_ ;
  assign \new_[81737]_  = A236 & A234;
  assign \new_[81738]_  = ~A233 & \new_[81737]_ ;
  assign \new_[81741]_  = ~A266 & A265;
  assign \new_[81744]_  = A269 & A267;
  assign \new_[81745]_  = \new_[81744]_  & \new_[81741]_ ;
  assign \new_[81746]_  = \new_[81745]_  & \new_[81738]_ ;
  assign \new_[81750]_  = A167 & ~A169;
  assign \new_[81751]_  = A170 & \new_[81750]_ ;
  assign \new_[81754]_  = A199 & ~A166;
  assign \new_[81757]_  = ~A232 & A200;
  assign \new_[81758]_  = \new_[81757]_  & \new_[81754]_ ;
  assign \new_[81759]_  = \new_[81758]_  & \new_[81751]_ ;
  assign \new_[81763]_  = ~A268 & ~A266;
  assign \new_[81764]_  = ~A233 & \new_[81763]_ ;
  assign \new_[81767]_  = A298 & ~A269;
  assign \new_[81770]_  = ~A302 & ~A301;
  assign \new_[81771]_  = \new_[81770]_  & \new_[81767]_ ;
  assign \new_[81772]_  = \new_[81771]_  & \new_[81764]_ ;
  assign \new_[81776]_  = A167 & ~A169;
  assign \new_[81777]_  = A170 & \new_[81776]_ ;
  assign \new_[81780]_  = ~A200 & ~A166;
  assign \new_[81783]_  = ~A203 & ~A202;
  assign \new_[81784]_  = \new_[81783]_  & \new_[81780]_ ;
  assign \new_[81785]_  = \new_[81784]_  & \new_[81777]_ ;
  assign \new_[81789]_  = A265 & A233;
  assign \new_[81790]_  = A232 & \new_[81789]_ ;
  assign \new_[81793]_  = ~A269 & ~A268;
  assign \new_[81796]_  = ~A300 & ~A299;
  assign \new_[81797]_  = \new_[81796]_  & \new_[81793]_ ;
  assign \new_[81798]_  = \new_[81797]_  & \new_[81790]_ ;
  assign \new_[81802]_  = A167 & ~A169;
  assign \new_[81803]_  = A170 & \new_[81802]_ ;
  assign \new_[81806]_  = ~A200 & ~A166;
  assign \new_[81809]_  = ~A203 & ~A202;
  assign \new_[81810]_  = \new_[81809]_  & \new_[81806]_ ;
  assign \new_[81811]_  = \new_[81810]_  & \new_[81803]_ ;
  assign \new_[81815]_  = A265 & A233;
  assign \new_[81816]_  = A232 & \new_[81815]_ ;
  assign \new_[81819]_  = ~A269 & ~A268;
  assign \new_[81822]_  = A299 & A298;
  assign \new_[81823]_  = \new_[81822]_  & \new_[81819]_ ;
  assign \new_[81824]_  = \new_[81823]_  & \new_[81816]_ ;
  assign \new_[81828]_  = A167 & ~A169;
  assign \new_[81829]_  = A170 & \new_[81828]_ ;
  assign \new_[81832]_  = ~A200 & ~A166;
  assign \new_[81835]_  = ~A203 & ~A202;
  assign \new_[81836]_  = \new_[81835]_  & \new_[81832]_ ;
  assign \new_[81837]_  = \new_[81836]_  & \new_[81829]_ ;
  assign \new_[81841]_  = A265 & A233;
  assign \new_[81842]_  = A232 & \new_[81841]_ ;
  assign \new_[81845]_  = ~A269 & ~A268;
  assign \new_[81848]_  = ~A299 & ~A298;
  assign \new_[81849]_  = \new_[81848]_  & \new_[81845]_ ;
  assign \new_[81850]_  = \new_[81849]_  & \new_[81842]_ ;
  assign \new_[81854]_  = A167 & ~A169;
  assign \new_[81855]_  = A170 & \new_[81854]_ ;
  assign \new_[81858]_  = ~A200 & ~A166;
  assign \new_[81861]_  = ~A203 & ~A202;
  assign \new_[81862]_  = \new_[81861]_  & \new_[81858]_ ;
  assign \new_[81863]_  = \new_[81862]_  & \new_[81855]_ ;
  assign \new_[81867]_  = A265 & A233;
  assign \new_[81868]_  = A232 & \new_[81867]_ ;
  assign \new_[81871]_  = ~A299 & ~A267;
  assign \new_[81874]_  = ~A302 & ~A301;
  assign \new_[81875]_  = \new_[81874]_  & \new_[81871]_ ;
  assign \new_[81876]_  = \new_[81875]_  & \new_[81868]_ ;
  assign \new_[81880]_  = A167 & ~A169;
  assign \new_[81881]_  = A170 & \new_[81880]_ ;
  assign \new_[81884]_  = ~A200 & ~A166;
  assign \new_[81887]_  = ~A203 & ~A202;
  assign \new_[81888]_  = \new_[81887]_  & \new_[81884]_ ;
  assign \new_[81889]_  = \new_[81888]_  & \new_[81881]_ ;
  assign \new_[81893]_  = A265 & A233;
  assign \new_[81894]_  = A232 & \new_[81893]_ ;
  assign \new_[81897]_  = ~A299 & A266;
  assign \new_[81900]_  = ~A302 & ~A301;
  assign \new_[81901]_  = \new_[81900]_  & \new_[81897]_ ;
  assign \new_[81902]_  = \new_[81901]_  & \new_[81894]_ ;
  assign \new_[81906]_  = A167 & ~A169;
  assign \new_[81907]_  = A170 & \new_[81906]_ ;
  assign \new_[81910]_  = ~A200 & ~A166;
  assign \new_[81913]_  = ~A203 & ~A202;
  assign \new_[81914]_  = \new_[81913]_  & \new_[81910]_ ;
  assign \new_[81915]_  = \new_[81914]_  & \new_[81907]_ ;
  assign \new_[81919]_  = ~A265 & A233;
  assign \new_[81920]_  = A232 & \new_[81919]_ ;
  assign \new_[81923]_  = ~A299 & ~A266;
  assign \new_[81926]_  = ~A302 & ~A301;
  assign \new_[81927]_  = \new_[81926]_  & \new_[81923]_ ;
  assign \new_[81928]_  = \new_[81927]_  & \new_[81920]_ ;
  assign \new_[81932]_  = A167 & ~A169;
  assign \new_[81933]_  = A170 & \new_[81932]_ ;
  assign \new_[81936]_  = ~A200 & ~A166;
  assign \new_[81939]_  = ~A203 & ~A202;
  assign \new_[81940]_  = \new_[81939]_  & \new_[81936]_ ;
  assign \new_[81941]_  = \new_[81940]_  & \new_[81933]_ ;
  assign \new_[81945]_  = ~A236 & ~A235;
  assign \new_[81946]_  = ~A233 & \new_[81945]_ ;
  assign \new_[81949]_  = A266 & A265;
  assign \new_[81952]_  = ~A300 & A298;
  assign \new_[81953]_  = \new_[81952]_  & \new_[81949]_ ;
  assign \new_[81954]_  = \new_[81953]_  & \new_[81946]_ ;
  assign \new_[81958]_  = A167 & ~A169;
  assign \new_[81959]_  = A170 & \new_[81958]_ ;
  assign \new_[81962]_  = ~A200 & ~A166;
  assign \new_[81965]_  = ~A203 & ~A202;
  assign \new_[81966]_  = \new_[81965]_  & \new_[81962]_ ;
  assign \new_[81967]_  = \new_[81966]_  & \new_[81959]_ ;
  assign \new_[81971]_  = ~A236 & ~A235;
  assign \new_[81972]_  = ~A233 & \new_[81971]_ ;
  assign \new_[81975]_  = A266 & A265;
  assign \new_[81978]_  = A299 & A298;
  assign \new_[81979]_  = \new_[81978]_  & \new_[81975]_ ;
  assign \new_[81980]_  = \new_[81979]_  & \new_[81972]_ ;
  assign \new_[81984]_  = A167 & ~A169;
  assign \new_[81985]_  = A170 & \new_[81984]_ ;
  assign \new_[81988]_  = ~A200 & ~A166;
  assign \new_[81991]_  = ~A203 & ~A202;
  assign \new_[81992]_  = \new_[81991]_  & \new_[81988]_ ;
  assign \new_[81993]_  = \new_[81992]_  & \new_[81985]_ ;
  assign \new_[81997]_  = ~A236 & ~A235;
  assign \new_[81998]_  = ~A233 & \new_[81997]_ ;
  assign \new_[82001]_  = A266 & A265;
  assign \new_[82004]_  = ~A299 & ~A298;
  assign \new_[82005]_  = \new_[82004]_  & \new_[82001]_ ;
  assign \new_[82006]_  = \new_[82005]_  & \new_[81998]_ ;
  assign \new_[82010]_  = A167 & ~A169;
  assign \new_[82011]_  = A170 & \new_[82010]_ ;
  assign \new_[82014]_  = ~A200 & ~A166;
  assign \new_[82017]_  = ~A203 & ~A202;
  assign \new_[82018]_  = \new_[82017]_  & \new_[82014]_ ;
  assign \new_[82019]_  = \new_[82018]_  & \new_[82011]_ ;
  assign \new_[82023]_  = ~A236 & ~A235;
  assign \new_[82024]_  = ~A233 & \new_[82023]_ ;
  assign \new_[82027]_  = ~A267 & ~A266;
  assign \new_[82030]_  = ~A300 & A298;
  assign \new_[82031]_  = \new_[82030]_  & \new_[82027]_ ;
  assign \new_[82032]_  = \new_[82031]_  & \new_[82024]_ ;
  assign \new_[82036]_  = A167 & ~A169;
  assign \new_[82037]_  = A170 & \new_[82036]_ ;
  assign \new_[82040]_  = ~A200 & ~A166;
  assign \new_[82043]_  = ~A203 & ~A202;
  assign \new_[82044]_  = \new_[82043]_  & \new_[82040]_ ;
  assign \new_[82045]_  = \new_[82044]_  & \new_[82037]_ ;
  assign \new_[82049]_  = ~A236 & ~A235;
  assign \new_[82050]_  = ~A233 & \new_[82049]_ ;
  assign \new_[82053]_  = ~A267 & ~A266;
  assign \new_[82056]_  = A299 & A298;
  assign \new_[82057]_  = \new_[82056]_  & \new_[82053]_ ;
  assign \new_[82058]_  = \new_[82057]_  & \new_[82050]_ ;
  assign \new_[82062]_  = A167 & ~A169;
  assign \new_[82063]_  = A170 & \new_[82062]_ ;
  assign \new_[82066]_  = ~A200 & ~A166;
  assign \new_[82069]_  = ~A203 & ~A202;
  assign \new_[82070]_  = \new_[82069]_  & \new_[82066]_ ;
  assign \new_[82071]_  = \new_[82070]_  & \new_[82063]_ ;
  assign \new_[82075]_  = ~A236 & ~A235;
  assign \new_[82076]_  = ~A233 & \new_[82075]_ ;
  assign \new_[82079]_  = ~A267 & ~A266;
  assign \new_[82082]_  = ~A299 & ~A298;
  assign \new_[82083]_  = \new_[82082]_  & \new_[82079]_ ;
  assign \new_[82084]_  = \new_[82083]_  & \new_[82076]_ ;
  assign \new_[82088]_  = A167 & ~A169;
  assign \new_[82089]_  = A170 & \new_[82088]_ ;
  assign \new_[82092]_  = ~A200 & ~A166;
  assign \new_[82095]_  = ~A203 & ~A202;
  assign \new_[82096]_  = \new_[82095]_  & \new_[82092]_ ;
  assign \new_[82097]_  = \new_[82096]_  & \new_[82089]_ ;
  assign \new_[82101]_  = ~A236 & ~A235;
  assign \new_[82102]_  = ~A233 & \new_[82101]_ ;
  assign \new_[82105]_  = ~A266 & ~A265;
  assign \new_[82108]_  = ~A300 & A298;
  assign \new_[82109]_  = \new_[82108]_  & \new_[82105]_ ;
  assign \new_[82110]_  = \new_[82109]_  & \new_[82102]_ ;
  assign \new_[82114]_  = A167 & ~A169;
  assign \new_[82115]_  = A170 & \new_[82114]_ ;
  assign \new_[82118]_  = ~A200 & ~A166;
  assign \new_[82121]_  = ~A203 & ~A202;
  assign \new_[82122]_  = \new_[82121]_  & \new_[82118]_ ;
  assign \new_[82123]_  = \new_[82122]_  & \new_[82115]_ ;
  assign \new_[82127]_  = ~A236 & ~A235;
  assign \new_[82128]_  = ~A233 & \new_[82127]_ ;
  assign \new_[82131]_  = ~A266 & ~A265;
  assign \new_[82134]_  = A299 & A298;
  assign \new_[82135]_  = \new_[82134]_  & \new_[82131]_ ;
  assign \new_[82136]_  = \new_[82135]_  & \new_[82128]_ ;
  assign \new_[82140]_  = A167 & ~A169;
  assign \new_[82141]_  = A170 & \new_[82140]_ ;
  assign \new_[82144]_  = ~A200 & ~A166;
  assign \new_[82147]_  = ~A203 & ~A202;
  assign \new_[82148]_  = \new_[82147]_  & \new_[82144]_ ;
  assign \new_[82149]_  = \new_[82148]_  & \new_[82141]_ ;
  assign \new_[82153]_  = ~A236 & ~A235;
  assign \new_[82154]_  = ~A233 & \new_[82153]_ ;
  assign \new_[82157]_  = ~A266 & ~A265;
  assign \new_[82160]_  = ~A299 & ~A298;
  assign \new_[82161]_  = \new_[82160]_  & \new_[82157]_ ;
  assign \new_[82162]_  = \new_[82161]_  & \new_[82154]_ ;
  assign \new_[82166]_  = A167 & ~A169;
  assign \new_[82167]_  = A170 & \new_[82166]_ ;
  assign \new_[82170]_  = ~A200 & ~A166;
  assign \new_[82173]_  = ~A203 & ~A202;
  assign \new_[82174]_  = \new_[82173]_  & \new_[82170]_ ;
  assign \new_[82175]_  = \new_[82174]_  & \new_[82167]_ ;
  assign \new_[82179]_  = A265 & ~A234;
  assign \new_[82180]_  = ~A233 & \new_[82179]_ ;
  assign \new_[82183]_  = A298 & A266;
  assign \new_[82186]_  = ~A302 & ~A301;
  assign \new_[82187]_  = \new_[82186]_  & \new_[82183]_ ;
  assign \new_[82188]_  = \new_[82187]_  & \new_[82180]_ ;
  assign \new_[82192]_  = A167 & ~A169;
  assign \new_[82193]_  = A170 & \new_[82192]_ ;
  assign \new_[82196]_  = ~A200 & ~A166;
  assign \new_[82199]_  = ~A203 & ~A202;
  assign \new_[82200]_  = \new_[82199]_  & \new_[82196]_ ;
  assign \new_[82201]_  = \new_[82200]_  & \new_[82193]_ ;
  assign \new_[82205]_  = ~A266 & ~A234;
  assign \new_[82206]_  = ~A233 & \new_[82205]_ ;
  assign \new_[82209]_  = ~A269 & ~A268;
  assign \new_[82212]_  = ~A300 & A298;
  assign \new_[82213]_  = \new_[82212]_  & \new_[82209]_ ;
  assign \new_[82214]_  = \new_[82213]_  & \new_[82206]_ ;
  assign \new_[82218]_  = A167 & ~A169;
  assign \new_[82219]_  = A170 & \new_[82218]_ ;
  assign \new_[82222]_  = ~A200 & ~A166;
  assign \new_[82225]_  = ~A203 & ~A202;
  assign \new_[82226]_  = \new_[82225]_  & \new_[82222]_ ;
  assign \new_[82227]_  = \new_[82226]_  & \new_[82219]_ ;
  assign \new_[82231]_  = ~A266 & ~A234;
  assign \new_[82232]_  = ~A233 & \new_[82231]_ ;
  assign \new_[82235]_  = ~A269 & ~A268;
  assign \new_[82238]_  = A299 & A298;
  assign \new_[82239]_  = \new_[82238]_  & \new_[82235]_ ;
  assign \new_[82240]_  = \new_[82239]_  & \new_[82232]_ ;
  assign \new_[82244]_  = A167 & ~A169;
  assign \new_[82245]_  = A170 & \new_[82244]_ ;
  assign \new_[82248]_  = ~A200 & ~A166;
  assign \new_[82251]_  = ~A203 & ~A202;
  assign \new_[82252]_  = \new_[82251]_  & \new_[82248]_ ;
  assign \new_[82253]_  = \new_[82252]_  & \new_[82245]_ ;
  assign \new_[82257]_  = ~A266 & ~A234;
  assign \new_[82258]_  = ~A233 & \new_[82257]_ ;
  assign \new_[82261]_  = ~A269 & ~A268;
  assign \new_[82264]_  = ~A299 & ~A298;
  assign \new_[82265]_  = \new_[82264]_  & \new_[82261]_ ;
  assign \new_[82266]_  = \new_[82265]_  & \new_[82258]_ ;
  assign \new_[82270]_  = A167 & ~A169;
  assign \new_[82271]_  = A170 & \new_[82270]_ ;
  assign \new_[82274]_  = ~A200 & ~A166;
  assign \new_[82277]_  = ~A203 & ~A202;
  assign \new_[82278]_  = \new_[82277]_  & \new_[82274]_ ;
  assign \new_[82279]_  = \new_[82278]_  & \new_[82271]_ ;
  assign \new_[82283]_  = ~A266 & ~A234;
  assign \new_[82284]_  = ~A233 & \new_[82283]_ ;
  assign \new_[82287]_  = A298 & ~A267;
  assign \new_[82290]_  = ~A302 & ~A301;
  assign \new_[82291]_  = \new_[82290]_  & \new_[82287]_ ;
  assign \new_[82292]_  = \new_[82291]_  & \new_[82284]_ ;
  assign \new_[82296]_  = A167 & ~A169;
  assign \new_[82297]_  = A170 & \new_[82296]_ ;
  assign \new_[82300]_  = ~A200 & ~A166;
  assign \new_[82303]_  = ~A203 & ~A202;
  assign \new_[82304]_  = \new_[82303]_  & \new_[82300]_ ;
  assign \new_[82305]_  = \new_[82304]_  & \new_[82297]_ ;
  assign \new_[82309]_  = ~A265 & ~A234;
  assign \new_[82310]_  = ~A233 & \new_[82309]_ ;
  assign \new_[82313]_  = A298 & ~A266;
  assign \new_[82316]_  = ~A302 & ~A301;
  assign \new_[82317]_  = \new_[82316]_  & \new_[82313]_ ;
  assign \new_[82318]_  = \new_[82317]_  & \new_[82310]_ ;
  assign \new_[82322]_  = A167 & ~A169;
  assign \new_[82323]_  = A170 & \new_[82322]_ ;
  assign \new_[82326]_  = ~A200 & ~A166;
  assign \new_[82329]_  = ~A203 & ~A202;
  assign \new_[82330]_  = \new_[82329]_  & \new_[82326]_ ;
  assign \new_[82331]_  = \new_[82330]_  & \new_[82323]_ ;
  assign \new_[82335]_  = A265 & ~A233;
  assign \new_[82336]_  = ~A232 & \new_[82335]_ ;
  assign \new_[82339]_  = A298 & A266;
  assign \new_[82342]_  = ~A302 & ~A301;
  assign \new_[82343]_  = \new_[82342]_  & \new_[82339]_ ;
  assign \new_[82344]_  = \new_[82343]_  & \new_[82336]_ ;
  assign \new_[82348]_  = A167 & ~A169;
  assign \new_[82349]_  = A170 & \new_[82348]_ ;
  assign \new_[82352]_  = ~A200 & ~A166;
  assign \new_[82355]_  = ~A203 & ~A202;
  assign \new_[82356]_  = \new_[82355]_  & \new_[82352]_ ;
  assign \new_[82357]_  = \new_[82356]_  & \new_[82349]_ ;
  assign \new_[82361]_  = ~A266 & ~A233;
  assign \new_[82362]_  = ~A232 & \new_[82361]_ ;
  assign \new_[82365]_  = ~A269 & ~A268;
  assign \new_[82368]_  = ~A300 & A298;
  assign \new_[82369]_  = \new_[82368]_  & \new_[82365]_ ;
  assign \new_[82370]_  = \new_[82369]_  & \new_[82362]_ ;
  assign \new_[82374]_  = A167 & ~A169;
  assign \new_[82375]_  = A170 & \new_[82374]_ ;
  assign \new_[82378]_  = ~A200 & ~A166;
  assign \new_[82381]_  = ~A203 & ~A202;
  assign \new_[82382]_  = \new_[82381]_  & \new_[82378]_ ;
  assign \new_[82383]_  = \new_[82382]_  & \new_[82375]_ ;
  assign \new_[82387]_  = ~A266 & ~A233;
  assign \new_[82388]_  = ~A232 & \new_[82387]_ ;
  assign \new_[82391]_  = ~A269 & ~A268;
  assign \new_[82394]_  = A299 & A298;
  assign \new_[82395]_  = \new_[82394]_  & \new_[82391]_ ;
  assign \new_[82396]_  = \new_[82395]_  & \new_[82388]_ ;
  assign \new_[82400]_  = A167 & ~A169;
  assign \new_[82401]_  = A170 & \new_[82400]_ ;
  assign \new_[82404]_  = ~A200 & ~A166;
  assign \new_[82407]_  = ~A203 & ~A202;
  assign \new_[82408]_  = \new_[82407]_  & \new_[82404]_ ;
  assign \new_[82409]_  = \new_[82408]_  & \new_[82401]_ ;
  assign \new_[82413]_  = ~A266 & ~A233;
  assign \new_[82414]_  = ~A232 & \new_[82413]_ ;
  assign \new_[82417]_  = ~A269 & ~A268;
  assign \new_[82420]_  = ~A299 & ~A298;
  assign \new_[82421]_  = \new_[82420]_  & \new_[82417]_ ;
  assign \new_[82422]_  = \new_[82421]_  & \new_[82414]_ ;
  assign \new_[82426]_  = A167 & ~A169;
  assign \new_[82427]_  = A170 & \new_[82426]_ ;
  assign \new_[82430]_  = ~A200 & ~A166;
  assign \new_[82433]_  = ~A203 & ~A202;
  assign \new_[82434]_  = \new_[82433]_  & \new_[82430]_ ;
  assign \new_[82435]_  = \new_[82434]_  & \new_[82427]_ ;
  assign \new_[82439]_  = ~A266 & ~A233;
  assign \new_[82440]_  = ~A232 & \new_[82439]_ ;
  assign \new_[82443]_  = A298 & ~A267;
  assign \new_[82446]_  = ~A302 & ~A301;
  assign \new_[82447]_  = \new_[82446]_  & \new_[82443]_ ;
  assign \new_[82448]_  = \new_[82447]_  & \new_[82440]_ ;
  assign \new_[82452]_  = A167 & ~A169;
  assign \new_[82453]_  = A170 & \new_[82452]_ ;
  assign \new_[82456]_  = ~A200 & ~A166;
  assign \new_[82459]_  = ~A203 & ~A202;
  assign \new_[82460]_  = \new_[82459]_  & \new_[82456]_ ;
  assign \new_[82461]_  = \new_[82460]_  & \new_[82453]_ ;
  assign \new_[82465]_  = ~A265 & ~A233;
  assign \new_[82466]_  = ~A232 & \new_[82465]_ ;
  assign \new_[82469]_  = A298 & ~A266;
  assign \new_[82472]_  = ~A302 & ~A301;
  assign \new_[82473]_  = \new_[82472]_  & \new_[82469]_ ;
  assign \new_[82474]_  = \new_[82473]_  & \new_[82466]_ ;
  assign \new_[82478]_  = A167 & ~A169;
  assign \new_[82479]_  = A170 & \new_[82478]_ ;
  assign \new_[82482]_  = ~A200 & ~A166;
  assign \new_[82485]_  = A232 & ~A201;
  assign \new_[82486]_  = \new_[82485]_  & \new_[82482]_ ;
  assign \new_[82487]_  = \new_[82486]_  & \new_[82479]_ ;
  assign \new_[82491]_  = ~A268 & A265;
  assign \new_[82492]_  = A233 & \new_[82491]_ ;
  assign \new_[82495]_  = ~A299 & ~A269;
  assign \new_[82498]_  = ~A302 & ~A301;
  assign \new_[82499]_  = \new_[82498]_  & \new_[82495]_ ;
  assign \new_[82500]_  = \new_[82499]_  & \new_[82492]_ ;
  assign \new_[82504]_  = A167 & ~A169;
  assign \new_[82505]_  = A170 & \new_[82504]_ ;
  assign \new_[82508]_  = ~A200 & ~A166;
  assign \new_[82511]_  = ~A233 & ~A201;
  assign \new_[82512]_  = \new_[82511]_  & \new_[82508]_ ;
  assign \new_[82513]_  = \new_[82512]_  & \new_[82505]_ ;
  assign \new_[82517]_  = A265 & ~A236;
  assign \new_[82518]_  = ~A235 & \new_[82517]_ ;
  assign \new_[82521]_  = A298 & A266;
  assign \new_[82524]_  = ~A302 & ~A301;
  assign \new_[82525]_  = \new_[82524]_  & \new_[82521]_ ;
  assign \new_[82526]_  = \new_[82525]_  & \new_[82518]_ ;
  assign \new_[82530]_  = A167 & ~A169;
  assign \new_[82531]_  = A170 & \new_[82530]_ ;
  assign \new_[82534]_  = ~A200 & ~A166;
  assign \new_[82537]_  = ~A233 & ~A201;
  assign \new_[82538]_  = \new_[82537]_  & \new_[82534]_ ;
  assign \new_[82539]_  = \new_[82538]_  & \new_[82531]_ ;
  assign \new_[82543]_  = ~A266 & ~A236;
  assign \new_[82544]_  = ~A235 & \new_[82543]_ ;
  assign \new_[82547]_  = ~A269 & ~A268;
  assign \new_[82550]_  = ~A300 & A298;
  assign \new_[82551]_  = \new_[82550]_  & \new_[82547]_ ;
  assign \new_[82552]_  = \new_[82551]_  & \new_[82544]_ ;
  assign \new_[82556]_  = A167 & ~A169;
  assign \new_[82557]_  = A170 & \new_[82556]_ ;
  assign \new_[82560]_  = ~A200 & ~A166;
  assign \new_[82563]_  = ~A233 & ~A201;
  assign \new_[82564]_  = \new_[82563]_  & \new_[82560]_ ;
  assign \new_[82565]_  = \new_[82564]_  & \new_[82557]_ ;
  assign \new_[82569]_  = ~A266 & ~A236;
  assign \new_[82570]_  = ~A235 & \new_[82569]_ ;
  assign \new_[82573]_  = ~A269 & ~A268;
  assign \new_[82576]_  = A299 & A298;
  assign \new_[82577]_  = \new_[82576]_  & \new_[82573]_ ;
  assign \new_[82578]_  = \new_[82577]_  & \new_[82570]_ ;
  assign \new_[82582]_  = A167 & ~A169;
  assign \new_[82583]_  = A170 & \new_[82582]_ ;
  assign \new_[82586]_  = ~A200 & ~A166;
  assign \new_[82589]_  = ~A233 & ~A201;
  assign \new_[82590]_  = \new_[82589]_  & \new_[82586]_ ;
  assign \new_[82591]_  = \new_[82590]_  & \new_[82583]_ ;
  assign \new_[82595]_  = ~A266 & ~A236;
  assign \new_[82596]_  = ~A235 & \new_[82595]_ ;
  assign \new_[82599]_  = ~A269 & ~A268;
  assign \new_[82602]_  = ~A299 & ~A298;
  assign \new_[82603]_  = \new_[82602]_  & \new_[82599]_ ;
  assign \new_[82604]_  = \new_[82603]_  & \new_[82596]_ ;
  assign \new_[82608]_  = A167 & ~A169;
  assign \new_[82609]_  = A170 & \new_[82608]_ ;
  assign \new_[82612]_  = ~A200 & ~A166;
  assign \new_[82615]_  = ~A233 & ~A201;
  assign \new_[82616]_  = \new_[82615]_  & \new_[82612]_ ;
  assign \new_[82617]_  = \new_[82616]_  & \new_[82609]_ ;
  assign \new_[82621]_  = ~A266 & ~A236;
  assign \new_[82622]_  = ~A235 & \new_[82621]_ ;
  assign \new_[82625]_  = A298 & ~A267;
  assign \new_[82628]_  = ~A302 & ~A301;
  assign \new_[82629]_  = \new_[82628]_  & \new_[82625]_ ;
  assign \new_[82630]_  = \new_[82629]_  & \new_[82622]_ ;
  assign \new_[82634]_  = A167 & ~A169;
  assign \new_[82635]_  = A170 & \new_[82634]_ ;
  assign \new_[82638]_  = ~A200 & ~A166;
  assign \new_[82641]_  = ~A233 & ~A201;
  assign \new_[82642]_  = \new_[82641]_  & \new_[82638]_ ;
  assign \new_[82643]_  = \new_[82642]_  & \new_[82635]_ ;
  assign \new_[82647]_  = ~A265 & ~A236;
  assign \new_[82648]_  = ~A235 & \new_[82647]_ ;
  assign \new_[82651]_  = A298 & ~A266;
  assign \new_[82654]_  = ~A302 & ~A301;
  assign \new_[82655]_  = \new_[82654]_  & \new_[82651]_ ;
  assign \new_[82656]_  = \new_[82655]_  & \new_[82648]_ ;
  assign \new_[82660]_  = A167 & ~A169;
  assign \new_[82661]_  = A170 & \new_[82660]_ ;
  assign \new_[82664]_  = ~A200 & ~A166;
  assign \new_[82667]_  = ~A233 & ~A201;
  assign \new_[82668]_  = \new_[82667]_  & \new_[82664]_ ;
  assign \new_[82669]_  = \new_[82668]_  & \new_[82661]_ ;
  assign \new_[82673]_  = ~A268 & ~A266;
  assign \new_[82674]_  = ~A234 & \new_[82673]_ ;
  assign \new_[82677]_  = A298 & ~A269;
  assign \new_[82680]_  = ~A302 & ~A301;
  assign \new_[82681]_  = \new_[82680]_  & \new_[82677]_ ;
  assign \new_[82682]_  = \new_[82681]_  & \new_[82674]_ ;
  assign \new_[82686]_  = A167 & ~A169;
  assign \new_[82687]_  = A170 & \new_[82686]_ ;
  assign \new_[82690]_  = ~A200 & ~A166;
  assign \new_[82693]_  = A232 & ~A201;
  assign \new_[82694]_  = \new_[82693]_  & \new_[82690]_ ;
  assign \new_[82695]_  = \new_[82694]_  & \new_[82687]_ ;
  assign \new_[82699]_  = A235 & A234;
  assign \new_[82700]_  = ~A233 & \new_[82699]_ ;
  assign \new_[82703]_  = ~A299 & A298;
  assign \new_[82706]_  = A301 & A300;
  assign \new_[82707]_  = \new_[82706]_  & \new_[82703]_ ;
  assign \new_[82708]_  = \new_[82707]_  & \new_[82700]_ ;
  assign \new_[82712]_  = A167 & ~A169;
  assign \new_[82713]_  = A170 & \new_[82712]_ ;
  assign \new_[82716]_  = ~A200 & ~A166;
  assign \new_[82719]_  = A232 & ~A201;
  assign \new_[82720]_  = \new_[82719]_  & \new_[82716]_ ;
  assign \new_[82721]_  = \new_[82720]_  & \new_[82713]_ ;
  assign \new_[82725]_  = A235 & A234;
  assign \new_[82726]_  = ~A233 & \new_[82725]_ ;
  assign \new_[82729]_  = ~A299 & A298;
  assign \new_[82732]_  = A302 & A300;
  assign \new_[82733]_  = \new_[82732]_  & \new_[82729]_ ;
  assign \new_[82734]_  = \new_[82733]_  & \new_[82726]_ ;
  assign \new_[82738]_  = A167 & ~A169;
  assign \new_[82739]_  = A170 & \new_[82738]_ ;
  assign \new_[82742]_  = ~A200 & ~A166;
  assign \new_[82745]_  = A232 & ~A201;
  assign \new_[82746]_  = \new_[82745]_  & \new_[82742]_ ;
  assign \new_[82747]_  = \new_[82746]_  & \new_[82739]_ ;
  assign \new_[82751]_  = A235 & A234;
  assign \new_[82752]_  = ~A233 & \new_[82751]_ ;
  assign \new_[82755]_  = ~A266 & A265;
  assign \new_[82758]_  = A268 & A267;
  assign \new_[82759]_  = \new_[82758]_  & \new_[82755]_ ;
  assign \new_[82760]_  = \new_[82759]_  & \new_[82752]_ ;
  assign \new_[82764]_  = A167 & ~A169;
  assign \new_[82765]_  = A170 & \new_[82764]_ ;
  assign \new_[82768]_  = ~A200 & ~A166;
  assign \new_[82771]_  = A232 & ~A201;
  assign \new_[82772]_  = \new_[82771]_  & \new_[82768]_ ;
  assign \new_[82773]_  = \new_[82772]_  & \new_[82765]_ ;
  assign \new_[82777]_  = A235 & A234;
  assign \new_[82778]_  = ~A233 & \new_[82777]_ ;
  assign \new_[82781]_  = ~A266 & A265;
  assign \new_[82784]_  = A269 & A267;
  assign \new_[82785]_  = \new_[82784]_  & \new_[82781]_ ;
  assign \new_[82786]_  = \new_[82785]_  & \new_[82778]_ ;
  assign \new_[82790]_  = A167 & ~A169;
  assign \new_[82791]_  = A170 & \new_[82790]_ ;
  assign \new_[82794]_  = ~A200 & ~A166;
  assign \new_[82797]_  = A232 & ~A201;
  assign \new_[82798]_  = \new_[82797]_  & \new_[82794]_ ;
  assign \new_[82799]_  = \new_[82798]_  & \new_[82791]_ ;
  assign \new_[82803]_  = A236 & A234;
  assign \new_[82804]_  = ~A233 & \new_[82803]_ ;
  assign \new_[82807]_  = ~A299 & A298;
  assign \new_[82810]_  = A301 & A300;
  assign \new_[82811]_  = \new_[82810]_  & \new_[82807]_ ;
  assign \new_[82812]_  = \new_[82811]_  & \new_[82804]_ ;
  assign \new_[82816]_  = A167 & ~A169;
  assign \new_[82817]_  = A170 & \new_[82816]_ ;
  assign \new_[82820]_  = ~A200 & ~A166;
  assign \new_[82823]_  = A232 & ~A201;
  assign \new_[82824]_  = \new_[82823]_  & \new_[82820]_ ;
  assign \new_[82825]_  = \new_[82824]_  & \new_[82817]_ ;
  assign \new_[82829]_  = A236 & A234;
  assign \new_[82830]_  = ~A233 & \new_[82829]_ ;
  assign \new_[82833]_  = ~A299 & A298;
  assign \new_[82836]_  = A302 & A300;
  assign \new_[82837]_  = \new_[82836]_  & \new_[82833]_ ;
  assign \new_[82838]_  = \new_[82837]_  & \new_[82830]_ ;
  assign \new_[82842]_  = A167 & ~A169;
  assign \new_[82843]_  = A170 & \new_[82842]_ ;
  assign \new_[82846]_  = ~A200 & ~A166;
  assign \new_[82849]_  = A232 & ~A201;
  assign \new_[82850]_  = \new_[82849]_  & \new_[82846]_ ;
  assign \new_[82851]_  = \new_[82850]_  & \new_[82843]_ ;
  assign \new_[82855]_  = A236 & A234;
  assign \new_[82856]_  = ~A233 & \new_[82855]_ ;
  assign \new_[82859]_  = ~A266 & A265;
  assign \new_[82862]_  = A268 & A267;
  assign \new_[82863]_  = \new_[82862]_  & \new_[82859]_ ;
  assign \new_[82864]_  = \new_[82863]_  & \new_[82856]_ ;
  assign \new_[82868]_  = A167 & ~A169;
  assign \new_[82869]_  = A170 & \new_[82868]_ ;
  assign \new_[82872]_  = ~A200 & ~A166;
  assign \new_[82875]_  = A232 & ~A201;
  assign \new_[82876]_  = \new_[82875]_  & \new_[82872]_ ;
  assign \new_[82877]_  = \new_[82876]_  & \new_[82869]_ ;
  assign \new_[82881]_  = A236 & A234;
  assign \new_[82882]_  = ~A233 & \new_[82881]_ ;
  assign \new_[82885]_  = ~A266 & A265;
  assign \new_[82888]_  = A269 & A267;
  assign \new_[82889]_  = \new_[82888]_  & \new_[82885]_ ;
  assign \new_[82890]_  = \new_[82889]_  & \new_[82882]_ ;
  assign \new_[82894]_  = A167 & ~A169;
  assign \new_[82895]_  = A170 & \new_[82894]_ ;
  assign \new_[82898]_  = ~A200 & ~A166;
  assign \new_[82901]_  = ~A232 & ~A201;
  assign \new_[82902]_  = \new_[82901]_  & \new_[82898]_ ;
  assign \new_[82903]_  = \new_[82902]_  & \new_[82895]_ ;
  assign \new_[82907]_  = ~A268 & ~A266;
  assign \new_[82908]_  = ~A233 & \new_[82907]_ ;
  assign \new_[82911]_  = A298 & ~A269;
  assign \new_[82914]_  = ~A302 & ~A301;
  assign \new_[82915]_  = \new_[82914]_  & \new_[82911]_ ;
  assign \new_[82916]_  = \new_[82915]_  & \new_[82908]_ ;
  assign \new_[82920]_  = A167 & ~A169;
  assign \new_[82921]_  = A170 & \new_[82920]_ ;
  assign \new_[82924]_  = ~A199 & ~A166;
  assign \new_[82927]_  = A232 & ~A200;
  assign \new_[82928]_  = \new_[82927]_  & \new_[82924]_ ;
  assign \new_[82929]_  = \new_[82928]_  & \new_[82921]_ ;
  assign \new_[82933]_  = ~A268 & A265;
  assign \new_[82934]_  = A233 & \new_[82933]_ ;
  assign \new_[82937]_  = ~A299 & ~A269;
  assign \new_[82940]_  = ~A302 & ~A301;
  assign \new_[82941]_  = \new_[82940]_  & \new_[82937]_ ;
  assign \new_[82942]_  = \new_[82941]_  & \new_[82934]_ ;
  assign \new_[82946]_  = A167 & ~A169;
  assign \new_[82947]_  = A170 & \new_[82946]_ ;
  assign \new_[82950]_  = ~A199 & ~A166;
  assign \new_[82953]_  = ~A233 & ~A200;
  assign \new_[82954]_  = \new_[82953]_  & \new_[82950]_ ;
  assign \new_[82955]_  = \new_[82954]_  & \new_[82947]_ ;
  assign \new_[82959]_  = A265 & ~A236;
  assign \new_[82960]_  = ~A235 & \new_[82959]_ ;
  assign \new_[82963]_  = A298 & A266;
  assign \new_[82966]_  = ~A302 & ~A301;
  assign \new_[82967]_  = \new_[82966]_  & \new_[82963]_ ;
  assign \new_[82968]_  = \new_[82967]_  & \new_[82960]_ ;
  assign \new_[82972]_  = A167 & ~A169;
  assign \new_[82973]_  = A170 & \new_[82972]_ ;
  assign \new_[82976]_  = ~A199 & ~A166;
  assign \new_[82979]_  = ~A233 & ~A200;
  assign \new_[82980]_  = \new_[82979]_  & \new_[82976]_ ;
  assign \new_[82981]_  = \new_[82980]_  & \new_[82973]_ ;
  assign \new_[82985]_  = ~A266 & ~A236;
  assign \new_[82986]_  = ~A235 & \new_[82985]_ ;
  assign \new_[82989]_  = ~A269 & ~A268;
  assign \new_[82992]_  = ~A300 & A298;
  assign \new_[82993]_  = \new_[82992]_  & \new_[82989]_ ;
  assign \new_[82994]_  = \new_[82993]_  & \new_[82986]_ ;
  assign \new_[82998]_  = A167 & ~A169;
  assign \new_[82999]_  = A170 & \new_[82998]_ ;
  assign \new_[83002]_  = ~A199 & ~A166;
  assign \new_[83005]_  = ~A233 & ~A200;
  assign \new_[83006]_  = \new_[83005]_  & \new_[83002]_ ;
  assign \new_[83007]_  = \new_[83006]_  & \new_[82999]_ ;
  assign \new_[83011]_  = ~A266 & ~A236;
  assign \new_[83012]_  = ~A235 & \new_[83011]_ ;
  assign \new_[83015]_  = ~A269 & ~A268;
  assign \new_[83018]_  = A299 & A298;
  assign \new_[83019]_  = \new_[83018]_  & \new_[83015]_ ;
  assign \new_[83020]_  = \new_[83019]_  & \new_[83012]_ ;
  assign \new_[83024]_  = A167 & ~A169;
  assign \new_[83025]_  = A170 & \new_[83024]_ ;
  assign \new_[83028]_  = ~A199 & ~A166;
  assign \new_[83031]_  = ~A233 & ~A200;
  assign \new_[83032]_  = \new_[83031]_  & \new_[83028]_ ;
  assign \new_[83033]_  = \new_[83032]_  & \new_[83025]_ ;
  assign \new_[83037]_  = ~A266 & ~A236;
  assign \new_[83038]_  = ~A235 & \new_[83037]_ ;
  assign \new_[83041]_  = ~A269 & ~A268;
  assign \new_[83044]_  = ~A299 & ~A298;
  assign \new_[83045]_  = \new_[83044]_  & \new_[83041]_ ;
  assign \new_[83046]_  = \new_[83045]_  & \new_[83038]_ ;
  assign \new_[83050]_  = A167 & ~A169;
  assign \new_[83051]_  = A170 & \new_[83050]_ ;
  assign \new_[83054]_  = ~A199 & ~A166;
  assign \new_[83057]_  = ~A233 & ~A200;
  assign \new_[83058]_  = \new_[83057]_  & \new_[83054]_ ;
  assign \new_[83059]_  = \new_[83058]_  & \new_[83051]_ ;
  assign \new_[83063]_  = ~A266 & ~A236;
  assign \new_[83064]_  = ~A235 & \new_[83063]_ ;
  assign \new_[83067]_  = A298 & ~A267;
  assign \new_[83070]_  = ~A302 & ~A301;
  assign \new_[83071]_  = \new_[83070]_  & \new_[83067]_ ;
  assign \new_[83072]_  = \new_[83071]_  & \new_[83064]_ ;
  assign \new_[83076]_  = A167 & ~A169;
  assign \new_[83077]_  = A170 & \new_[83076]_ ;
  assign \new_[83080]_  = ~A199 & ~A166;
  assign \new_[83083]_  = ~A233 & ~A200;
  assign \new_[83084]_  = \new_[83083]_  & \new_[83080]_ ;
  assign \new_[83085]_  = \new_[83084]_  & \new_[83077]_ ;
  assign \new_[83089]_  = ~A265 & ~A236;
  assign \new_[83090]_  = ~A235 & \new_[83089]_ ;
  assign \new_[83093]_  = A298 & ~A266;
  assign \new_[83096]_  = ~A302 & ~A301;
  assign \new_[83097]_  = \new_[83096]_  & \new_[83093]_ ;
  assign \new_[83098]_  = \new_[83097]_  & \new_[83090]_ ;
  assign \new_[83102]_  = A167 & ~A169;
  assign \new_[83103]_  = A170 & \new_[83102]_ ;
  assign \new_[83106]_  = ~A199 & ~A166;
  assign \new_[83109]_  = ~A233 & ~A200;
  assign \new_[83110]_  = \new_[83109]_  & \new_[83106]_ ;
  assign \new_[83111]_  = \new_[83110]_  & \new_[83103]_ ;
  assign \new_[83115]_  = ~A268 & ~A266;
  assign \new_[83116]_  = ~A234 & \new_[83115]_ ;
  assign \new_[83119]_  = A298 & ~A269;
  assign \new_[83122]_  = ~A302 & ~A301;
  assign \new_[83123]_  = \new_[83122]_  & \new_[83119]_ ;
  assign \new_[83124]_  = \new_[83123]_  & \new_[83116]_ ;
  assign \new_[83128]_  = A167 & ~A169;
  assign \new_[83129]_  = A170 & \new_[83128]_ ;
  assign \new_[83132]_  = ~A199 & ~A166;
  assign \new_[83135]_  = A232 & ~A200;
  assign \new_[83136]_  = \new_[83135]_  & \new_[83132]_ ;
  assign \new_[83137]_  = \new_[83136]_  & \new_[83129]_ ;
  assign \new_[83141]_  = A235 & A234;
  assign \new_[83142]_  = ~A233 & \new_[83141]_ ;
  assign \new_[83145]_  = ~A299 & A298;
  assign \new_[83148]_  = A301 & A300;
  assign \new_[83149]_  = \new_[83148]_  & \new_[83145]_ ;
  assign \new_[83150]_  = \new_[83149]_  & \new_[83142]_ ;
  assign \new_[83154]_  = A167 & ~A169;
  assign \new_[83155]_  = A170 & \new_[83154]_ ;
  assign \new_[83158]_  = ~A199 & ~A166;
  assign \new_[83161]_  = A232 & ~A200;
  assign \new_[83162]_  = \new_[83161]_  & \new_[83158]_ ;
  assign \new_[83163]_  = \new_[83162]_  & \new_[83155]_ ;
  assign \new_[83167]_  = A235 & A234;
  assign \new_[83168]_  = ~A233 & \new_[83167]_ ;
  assign \new_[83171]_  = ~A299 & A298;
  assign \new_[83174]_  = A302 & A300;
  assign \new_[83175]_  = \new_[83174]_  & \new_[83171]_ ;
  assign \new_[83176]_  = \new_[83175]_  & \new_[83168]_ ;
  assign \new_[83180]_  = A167 & ~A169;
  assign \new_[83181]_  = A170 & \new_[83180]_ ;
  assign \new_[83184]_  = ~A199 & ~A166;
  assign \new_[83187]_  = A232 & ~A200;
  assign \new_[83188]_  = \new_[83187]_  & \new_[83184]_ ;
  assign \new_[83189]_  = \new_[83188]_  & \new_[83181]_ ;
  assign \new_[83193]_  = A235 & A234;
  assign \new_[83194]_  = ~A233 & \new_[83193]_ ;
  assign \new_[83197]_  = ~A266 & A265;
  assign \new_[83200]_  = A268 & A267;
  assign \new_[83201]_  = \new_[83200]_  & \new_[83197]_ ;
  assign \new_[83202]_  = \new_[83201]_  & \new_[83194]_ ;
  assign \new_[83206]_  = A167 & ~A169;
  assign \new_[83207]_  = A170 & \new_[83206]_ ;
  assign \new_[83210]_  = ~A199 & ~A166;
  assign \new_[83213]_  = A232 & ~A200;
  assign \new_[83214]_  = \new_[83213]_  & \new_[83210]_ ;
  assign \new_[83215]_  = \new_[83214]_  & \new_[83207]_ ;
  assign \new_[83219]_  = A235 & A234;
  assign \new_[83220]_  = ~A233 & \new_[83219]_ ;
  assign \new_[83223]_  = ~A266 & A265;
  assign \new_[83226]_  = A269 & A267;
  assign \new_[83227]_  = \new_[83226]_  & \new_[83223]_ ;
  assign \new_[83228]_  = \new_[83227]_  & \new_[83220]_ ;
  assign \new_[83232]_  = A167 & ~A169;
  assign \new_[83233]_  = A170 & \new_[83232]_ ;
  assign \new_[83236]_  = ~A199 & ~A166;
  assign \new_[83239]_  = A232 & ~A200;
  assign \new_[83240]_  = \new_[83239]_  & \new_[83236]_ ;
  assign \new_[83241]_  = \new_[83240]_  & \new_[83233]_ ;
  assign \new_[83245]_  = A236 & A234;
  assign \new_[83246]_  = ~A233 & \new_[83245]_ ;
  assign \new_[83249]_  = ~A299 & A298;
  assign \new_[83252]_  = A301 & A300;
  assign \new_[83253]_  = \new_[83252]_  & \new_[83249]_ ;
  assign \new_[83254]_  = \new_[83253]_  & \new_[83246]_ ;
  assign \new_[83258]_  = A167 & ~A169;
  assign \new_[83259]_  = A170 & \new_[83258]_ ;
  assign \new_[83262]_  = ~A199 & ~A166;
  assign \new_[83265]_  = A232 & ~A200;
  assign \new_[83266]_  = \new_[83265]_  & \new_[83262]_ ;
  assign \new_[83267]_  = \new_[83266]_  & \new_[83259]_ ;
  assign \new_[83271]_  = A236 & A234;
  assign \new_[83272]_  = ~A233 & \new_[83271]_ ;
  assign \new_[83275]_  = ~A299 & A298;
  assign \new_[83278]_  = A302 & A300;
  assign \new_[83279]_  = \new_[83278]_  & \new_[83275]_ ;
  assign \new_[83280]_  = \new_[83279]_  & \new_[83272]_ ;
  assign \new_[83284]_  = A167 & ~A169;
  assign \new_[83285]_  = A170 & \new_[83284]_ ;
  assign \new_[83288]_  = ~A199 & ~A166;
  assign \new_[83291]_  = A232 & ~A200;
  assign \new_[83292]_  = \new_[83291]_  & \new_[83288]_ ;
  assign \new_[83293]_  = \new_[83292]_  & \new_[83285]_ ;
  assign \new_[83297]_  = A236 & A234;
  assign \new_[83298]_  = ~A233 & \new_[83297]_ ;
  assign \new_[83301]_  = ~A266 & A265;
  assign \new_[83304]_  = A268 & A267;
  assign \new_[83305]_  = \new_[83304]_  & \new_[83301]_ ;
  assign \new_[83306]_  = \new_[83305]_  & \new_[83298]_ ;
  assign \new_[83310]_  = A167 & ~A169;
  assign \new_[83311]_  = A170 & \new_[83310]_ ;
  assign \new_[83314]_  = ~A199 & ~A166;
  assign \new_[83317]_  = A232 & ~A200;
  assign \new_[83318]_  = \new_[83317]_  & \new_[83314]_ ;
  assign \new_[83319]_  = \new_[83318]_  & \new_[83311]_ ;
  assign \new_[83323]_  = A236 & A234;
  assign \new_[83324]_  = ~A233 & \new_[83323]_ ;
  assign \new_[83327]_  = ~A266 & A265;
  assign \new_[83330]_  = A269 & A267;
  assign \new_[83331]_  = \new_[83330]_  & \new_[83327]_ ;
  assign \new_[83332]_  = \new_[83331]_  & \new_[83324]_ ;
  assign \new_[83336]_  = A167 & ~A169;
  assign \new_[83337]_  = A170 & \new_[83336]_ ;
  assign \new_[83340]_  = ~A199 & ~A166;
  assign \new_[83343]_  = ~A232 & ~A200;
  assign \new_[83344]_  = \new_[83343]_  & \new_[83340]_ ;
  assign \new_[83345]_  = \new_[83344]_  & \new_[83337]_ ;
  assign \new_[83349]_  = ~A268 & ~A266;
  assign \new_[83350]_  = ~A233 & \new_[83349]_ ;
  assign \new_[83353]_  = A298 & ~A269;
  assign \new_[83356]_  = ~A302 & ~A301;
  assign \new_[83357]_  = \new_[83356]_  & \new_[83353]_ ;
  assign \new_[83358]_  = \new_[83357]_  & \new_[83350]_ ;
  assign \new_[83362]_  = ~A167 & ~A169;
  assign \new_[83363]_  = A170 & \new_[83362]_ ;
  assign \new_[83366]_  = A199 & A166;
  assign \new_[83369]_  = A232 & A200;
  assign \new_[83370]_  = \new_[83369]_  & \new_[83366]_ ;
  assign \new_[83371]_  = \new_[83370]_  & \new_[83363]_ ;
  assign \new_[83375]_  = ~A268 & A265;
  assign \new_[83376]_  = A233 & \new_[83375]_ ;
  assign \new_[83379]_  = ~A299 & ~A269;
  assign \new_[83382]_  = ~A302 & ~A301;
  assign \new_[83383]_  = \new_[83382]_  & \new_[83379]_ ;
  assign \new_[83384]_  = \new_[83383]_  & \new_[83376]_ ;
  assign \new_[83388]_  = ~A167 & ~A169;
  assign \new_[83389]_  = A170 & \new_[83388]_ ;
  assign \new_[83392]_  = A199 & A166;
  assign \new_[83395]_  = ~A233 & A200;
  assign \new_[83396]_  = \new_[83395]_  & \new_[83392]_ ;
  assign \new_[83397]_  = \new_[83396]_  & \new_[83389]_ ;
  assign \new_[83401]_  = A265 & ~A236;
  assign \new_[83402]_  = ~A235 & \new_[83401]_ ;
  assign \new_[83405]_  = A298 & A266;
  assign \new_[83408]_  = ~A302 & ~A301;
  assign \new_[83409]_  = \new_[83408]_  & \new_[83405]_ ;
  assign \new_[83410]_  = \new_[83409]_  & \new_[83402]_ ;
  assign \new_[83414]_  = ~A167 & ~A169;
  assign \new_[83415]_  = A170 & \new_[83414]_ ;
  assign \new_[83418]_  = A199 & A166;
  assign \new_[83421]_  = ~A233 & A200;
  assign \new_[83422]_  = \new_[83421]_  & \new_[83418]_ ;
  assign \new_[83423]_  = \new_[83422]_  & \new_[83415]_ ;
  assign \new_[83427]_  = ~A266 & ~A236;
  assign \new_[83428]_  = ~A235 & \new_[83427]_ ;
  assign \new_[83431]_  = ~A269 & ~A268;
  assign \new_[83434]_  = ~A300 & A298;
  assign \new_[83435]_  = \new_[83434]_  & \new_[83431]_ ;
  assign \new_[83436]_  = \new_[83435]_  & \new_[83428]_ ;
  assign \new_[83440]_  = ~A167 & ~A169;
  assign \new_[83441]_  = A170 & \new_[83440]_ ;
  assign \new_[83444]_  = A199 & A166;
  assign \new_[83447]_  = ~A233 & A200;
  assign \new_[83448]_  = \new_[83447]_  & \new_[83444]_ ;
  assign \new_[83449]_  = \new_[83448]_  & \new_[83441]_ ;
  assign \new_[83453]_  = ~A266 & ~A236;
  assign \new_[83454]_  = ~A235 & \new_[83453]_ ;
  assign \new_[83457]_  = ~A269 & ~A268;
  assign \new_[83460]_  = A299 & A298;
  assign \new_[83461]_  = \new_[83460]_  & \new_[83457]_ ;
  assign \new_[83462]_  = \new_[83461]_  & \new_[83454]_ ;
  assign \new_[83466]_  = ~A167 & ~A169;
  assign \new_[83467]_  = A170 & \new_[83466]_ ;
  assign \new_[83470]_  = A199 & A166;
  assign \new_[83473]_  = ~A233 & A200;
  assign \new_[83474]_  = \new_[83473]_  & \new_[83470]_ ;
  assign \new_[83475]_  = \new_[83474]_  & \new_[83467]_ ;
  assign \new_[83479]_  = ~A266 & ~A236;
  assign \new_[83480]_  = ~A235 & \new_[83479]_ ;
  assign \new_[83483]_  = ~A269 & ~A268;
  assign \new_[83486]_  = ~A299 & ~A298;
  assign \new_[83487]_  = \new_[83486]_  & \new_[83483]_ ;
  assign \new_[83488]_  = \new_[83487]_  & \new_[83480]_ ;
  assign \new_[83492]_  = ~A167 & ~A169;
  assign \new_[83493]_  = A170 & \new_[83492]_ ;
  assign \new_[83496]_  = A199 & A166;
  assign \new_[83499]_  = ~A233 & A200;
  assign \new_[83500]_  = \new_[83499]_  & \new_[83496]_ ;
  assign \new_[83501]_  = \new_[83500]_  & \new_[83493]_ ;
  assign \new_[83505]_  = ~A266 & ~A236;
  assign \new_[83506]_  = ~A235 & \new_[83505]_ ;
  assign \new_[83509]_  = A298 & ~A267;
  assign \new_[83512]_  = ~A302 & ~A301;
  assign \new_[83513]_  = \new_[83512]_  & \new_[83509]_ ;
  assign \new_[83514]_  = \new_[83513]_  & \new_[83506]_ ;
  assign \new_[83518]_  = ~A167 & ~A169;
  assign \new_[83519]_  = A170 & \new_[83518]_ ;
  assign \new_[83522]_  = A199 & A166;
  assign \new_[83525]_  = ~A233 & A200;
  assign \new_[83526]_  = \new_[83525]_  & \new_[83522]_ ;
  assign \new_[83527]_  = \new_[83526]_  & \new_[83519]_ ;
  assign \new_[83531]_  = ~A265 & ~A236;
  assign \new_[83532]_  = ~A235 & \new_[83531]_ ;
  assign \new_[83535]_  = A298 & ~A266;
  assign \new_[83538]_  = ~A302 & ~A301;
  assign \new_[83539]_  = \new_[83538]_  & \new_[83535]_ ;
  assign \new_[83540]_  = \new_[83539]_  & \new_[83532]_ ;
  assign \new_[83544]_  = ~A167 & ~A169;
  assign \new_[83545]_  = A170 & \new_[83544]_ ;
  assign \new_[83548]_  = A199 & A166;
  assign \new_[83551]_  = ~A233 & A200;
  assign \new_[83552]_  = \new_[83551]_  & \new_[83548]_ ;
  assign \new_[83553]_  = \new_[83552]_  & \new_[83545]_ ;
  assign \new_[83557]_  = ~A268 & ~A266;
  assign \new_[83558]_  = ~A234 & \new_[83557]_ ;
  assign \new_[83561]_  = A298 & ~A269;
  assign \new_[83564]_  = ~A302 & ~A301;
  assign \new_[83565]_  = \new_[83564]_  & \new_[83561]_ ;
  assign \new_[83566]_  = \new_[83565]_  & \new_[83558]_ ;
  assign \new_[83570]_  = ~A167 & ~A169;
  assign \new_[83571]_  = A170 & \new_[83570]_ ;
  assign \new_[83574]_  = A199 & A166;
  assign \new_[83577]_  = A232 & A200;
  assign \new_[83578]_  = \new_[83577]_  & \new_[83574]_ ;
  assign \new_[83579]_  = \new_[83578]_  & \new_[83571]_ ;
  assign \new_[83583]_  = A235 & A234;
  assign \new_[83584]_  = ~A233 & \new_[83583]_ ;
  assign \new_[83587]_  = ~A299 & A298;
  assign \new_[83590]_  = A301 & A300;
  assign \new_[83591]_  = \new_[83590]_  & \new_[83587]_ ;
  assign \new_[83592]_  = \new_[83591]_  & \new_[83584]_ ;
  assign \new_[83596]_  = ~A167 & ~A169;
  assign \new_[83597]_  = A170 & \new_[83596]_ ;
  assign \new_[83600]_  = A199 & A166;
  assign \new_[83603]_  = A232 & A200;
  assign \new_[83604]_  = \new_[83603]_  & \new_[83600]_ ;
  assign \new_[83605]_  = \new_[83604]_  & \new_[83597]_ ;
  assign \new_[83609]_  = A235 & A234;
  assign \new_[83610]_  = ~A233 & \new_[83609]_ ;
  assign \new_[83613]_  = ~A299 & A298;
  assign \new_[83616]_  = A302 & A300;
  assign \new_[83617]_  = \new_[83616]_  & \new_[83613]_ ;
  assign \new_[83618]_  = \new_[83617]_  & \new_[83610]_ ;
  assign \new_[83622]_  = ~A167 & ~A169;
  assign \new_[83623]_  = A170 & \new_[83622]_ ;
  assign \new_[83626]_  = A199 & A166;
  assign \new_[83629]_  = A232 & A200;
  assign \new_[83630]_  = \new_[83629]_  & \new_[83626]_ ;
  assign \new_[83631]_  = \new_[83630]_  & \new_[83623]_ ;
  assign \new_[83635]_  = A235 & A234;
  assign \new_[83636]_  = ~A233 & \new_[83635]_ ;
  assign \new_[83639]_  = ~A266 & A265;
  assign \new_[83642]_  = A268 & A267;
  assign \new_[83643]_  = \new_[83642]_  & \new_[83639]_ ;
  assign \new_[83644]_  = \new_[83643]_  & \new_[83636]_ ;
  assign \new_[83648]_  = ~A167 & ~A169;
  assign \new_[83649]_  = A170 & \new_[83648]_ ;
  assign \new_[83652]_  = A199 & A166;
  assign \new_[83655]_  = A232 & A200;
  assign \new_[83656]_  = \new_[83655]_  & \new_[83652]_ ;
  assign \new_[83657]_  = \new_[83656]_  & \new_[83649]_ ;
  assign \new_[83661]_  = A235 & A234;
  assign \new_[83662]_  = ~A233 & \new_[83661]_ ;
  assign \new_[83665]_  = ~A266 & A265;
  assign \new_[83668]_  = A269 & A267;
  assign \new_[83669]_  = \new_[83668]_  & \new_[83665]_ ;
  assign \new_[83670]_  = \new_[83669]_  & \new_[83662]_ ;
  assign \new_[83674]_  = ~A167 & ~A169;
  assign \new_[83675]_  = A170 & \new_[83674]_ ;
  assign \new_[83678]_  = A199 & A166;
  assign \new_[83681]_  = A232 & A200;
  assign \new_[83682]_  = \new_[83681]_  & \new_[83678]_ ;
  assign \new_[83683]_  = \new_[83682]_  & \new_[83675]_ ;
  assign \new_[83687]_  = A236 & A234;
  assign \new_[83688]_  = ~A233 & \new_[83687]_ ;
  assign \new_[83691]_  = ~A299 & A298;
  assign \new_[83694]_  = A301 & A300;
  assign \new_[83695]_  = \new_[83694]_  & \new_[83691]_ ;
  assign \new_[83696]_  = \new_[83695]_  & \new_[83688]_ ;
  assign \new_[83700]_  = ~A167 & ~A169;
  assign \new_[83701]_  = A170 & \new_[83700]_ ;
  assign \new_[83704]_  = A199 & A166;
  assign \new_[83707]_  = A232 & A200;
  assign \new_[83708]_  = \new_[83707]_  & \new_[83704]_ ;
  assign \new_[83709]_  = \new_[83708]_  & \new_[83701]_ ;
  assign \new_[83713]_  = A236 & A234;
  assign \new_[83714]_  = ~A233 & \new_[83713]_ ;
  assign \new_[83717]_  = ~A299 & A298;
  assign \new_[83720]_  = A302 & A300;
  assign \new_[83721]_  = \new_[83720]_  & \new_[83717]_ ;
  assign \new_[83722]_  = \new_[83721]_  & \new_[83714]_ ;
  assign \new_[83726]_  = ~A167 & ~A169;
  assign \new_[83727]_  = A170 & \new_[83726]_ ;
  assign \new_[83730]_  = A199 & A166;
  assign \new_[83733]_  = A232 & A200;
  assign \new_[83734]_  = \new_[83733]_  & \new_[83730]_ ;
  assign \new_[83735]_  = \new_[83734]_  & \new_[83727]_ ;
  assign \new_[83739]_  = A236 & A234;
  assign \new_[83740]_  = ~A233 & \new_[83739]_ ;
  assign \new_[83743]_  = ~A266 & A265;
  assign \new_[83746]_  = A268 & A267;
  assign \new_[83747]_  = \new_[83746]_  & \new_[83743]_ ;
  assign \new_[83748]_  = \new_[83747]_  & \new_[83740]_ ;
  assign \new_[83752]_  = ~A167 & ~A169;
  assign \new_[83753]_  = A170 & \new_[83752]_ ;
  assign \new_[83756]_  = A199 & A166;
  assign \new_[83759]_  = A232 & A200;
  assign \new_[83760]_  = \new_[83759]_  & \new_[83756]_ ;
  assign \new_[83761]_  = \new_[83760]_  & \new_[83753]_ ;
  assign \new_[83765]_  = A236 & A234;
  assign \new_[83766]_  = ~A233 & \new_[83765]_ ;
  assign \new_[83769]_  = ~A266 & A265;
  assign \new_[83772]_  = A269 & A267;
  assign \new_[83773]_  = \new_[83772]_  & \new_[83769]_ ;
  assign \new_[83774]_  = \new_[83773]_  & \new_[83766]_ ;
  assign \new_[83778]_  = ~A167 & ~A169;
  assign \new_[83779]_  = A170 & \new_[83778]_ ;
  assign \new_[83782]_  = A199 & A166;
  assign \new_[83785]_  = ~A232 & A200;
  assign \new_[83786]_  = \new_[83785]_  & \new_[83782]_ ;
  assign \new_[83787]_  = \new_[83786]_  & \new_[83779]_ ;
  assign \new_[83791]_  = ~A268 & ~A266;
  assign \new_[83792]_  = ~A233 & \new_[83791]_ ;
  assign \new_[83795]_  = A298 & ~A269;
  assign \new_[83798]_  = ~A302 & ~A301;
  assign \new_[83799]_  = \new_[83798]_  & \new_[83795]_ ;
  assign \new_[83800]_  = \new_[83799]_  & \new_[83792]_ ;
  assign \new_[83804]_  = ~A167 & ~A169;
  assign \new_[83805]_  = A170 & \new_[83804]_ ;
  assign \new_[83808]_  = ~A200 & A166;
  assign \new_[83811]_  = ~A203 & ~A202;
  assign \new_[83812]_  = \new_[83811]_  & \new_[83808]_ ;
  assign \new_[83813]_  = \new_[83812]_  & \new_[83805]_ ;
  assign \new_[83817]_  = A265 & A233;
  assign \new_[83818]_  = A232 & \new_[83817]_ ;
  assign \new_[83821]_  = ~A269 & ~A268;
  assign \new_[83824]_  = ~A300 & ~A299;
  assign \new_[83825]_  = \new_[83824]_  & \new_[83821]_ ;
  assign \new_[83826]_  = \new_[83825]_  & \new_[83818]_ ;
  assign \new_[83830]_  = ~A167 & ~A169;
  assign \new_[83831]_  = A170 & \new_[83830]_ ;
  assign \new_[83834]_  = ~A200 & A166;
  assign \new_[83837]_  = ~A203 & ~A202;
  assign \new_[83838]_  = \new_[83837]_  & \new_[83834]_ ;
  assign \new_[83839]_  = \new_[83838]_  & \new_[83831]_ ;
  assign \new_[83843]_  = A265 & A233;
  assign \new_[83844]_  = A232 & \new_[83843]_ ;
  assign \new_[83847]_  = ~A269 & ~A268;
  assign \new_[83850]_  = A299 & A298;
  assign \new_[83851]_  = \new_[83850]_  & \new_[83847]_ ;
  assign \new_[83852]_  = \new_[83851]_  & \new_[83844]_ ;
  assign \new_[83856]_  = ~A167 & ~A169;
  assign \new_[83857]_  = A170 & \new_[83856]_ ;
  assign \new_[83860]_  = ~A200 & A166;
  assign \new_[83863]_  = ~A203 & ~A202;
  assign \new_[83864]_  = \new_[83863]_  & \new_[83860]_ ;
  assign \new_[83865]_  = \new_[83864]_  & \new_[83857]_ ;
  assign \new_[83869]_  = A265 & A233;
  assign \new_[83870]_  = A232 & \new_[83869]_ ;
  assign \new_[83873]_  = ~A269 & ~A268;
  assign \new_[83876]_  = ~A299 & ~A298;
  assign \new_[83877]_  = \new_[83876]_  & \new_[83873]_ ;
  assign \new_[83878]_  = \new_[83877]_  & \new_[83870]_ ;
  assign \new_[83882]_  = ~A167 & ~A169;
  assign \new_[83883]_  = A170 & \new_[83882]_ ;
  assign \new_[83886]_  = ~A200 & A166;
  assign \new_[83889]_  = ~A203 & ~A202;
  assign \new_[83890]_  = \new_[83889]_  & \new_[83886]_ ;
  assign \new_[83891]_  = \new_[83890]_  & \new_[83883]_ ;
  assign \new_[83895]_  = A265 & A233;
  assign \new_[83896]_  = A232 & \new_[83895]_ ;
  assign \new_[83899]_  = ~A299 & ~A267;
  assign \new_[83902]_  = ~A302 & ~A301;
  assign \new_[83903]_  = \new_[83902]_  & \new_[83899]_ ;
  assign \new_[83904]_  = \new_[83903]_  & \new_[83896]_ ;
  assign \new_[83908]_  = ~A167 & ~A169;
  assign \new_[83909]_  = A170 & \new_[83908]_ ;
  assign \new_[83912]_  = ~A200 & A166;
  assign \new_[83915]_  = ~A203 & ~A202;
  assign \new_[83916]_  = \new_[83915]_  & \new_[83912]_ ;
  assign \new_[83917]_  = \new_[83916]_  & \new_[83909]_ ;
  assign \new_[83921]_  = A265 & A233;
  assign \new_[83922]_  = A232 & \new_[83921]_ ;
  assign \new_[83925]_  = ~A299 & A266;
  assign \new_[83928]_  = ~A302 & ~A301;
  assign \new_[83929]_  = \new_[83928]_  & \new_[83925]_ ;
  assign \new_[83930]_  = \new_[83929]_  & \new_[83922]_ ;
  assign \new_[83934]_  = ~A167 & ~A169;
  assign \new_[83935]_  = A170 & \new_[83934]_ ;
  assign \new_[83938]_  = ~A200 & A166;
  assign \new_[83941]_  = ~A203 & ~A202;
  assign \new_[83942]_  = \new_[83941]_  & \new_[83938]_ ;
  assign \new_[83943]_  = \new_[83942]_  & \new_[83935]_ ;
  assign \new_[83947]_  = ~A265 & A233;
  assign \new_[83948]_  = A232 & \new_[83947]_ ;
  assign \new_[83951]_  = ~A299 & ~A266;
  assign \new_[83954]_  = ~A302 & ~A301;
  assign \new_[83955]_  = \new_[83954]_  & \new_[83951]_ ;
  assign \new_[83956]_  = \new_[83955]_  & \new_[83948]_ ;
  assign \new_[83960]_  = ~A167 & ~A169;
  assign \new_[83961]_  = A170 & \new_[83960]_ ;
  assign \new_[83964]_  = ~A200 & A166;
  assign \new_[83967]_  = ~A203 & ~A202;
  assign \new_[83968]_  = \new_[83967]_  & \new_[83964]_ ;
  assign \new_[83969]_  = \new_[83968]_  & \new_[83961]_ ;
  assign \new_[83973]_  = ~A236 & ~A235;
  assign \new_[83974]_  = ~A233 & \new_[83973]_ ;
  assign \new_[83977]_  = A266 & A265;
  assign \new_[83980]_  = ~A300 & A298;
  assign \new_[83981]_  = \new_[83980]_  & \new_[83977]_ ;
  assign \new_[83982]_  = \new_[83981]_  & \new_[83974]_ ;
  assign \new_[83986]_  = ~A167 & ~A169;
  assign \new_[83987]_  = A170 & \new_[83986]_ ;
  assign \new_[83990]_  = ~A200 & A166;
  assign \new_[83993]_  = ~A203 & ~A202;
  assign \new_[83994]_  = \new_[83993]_  & \new_[83990]_ ;
  assign \new_[83995]_  = \new_[83994]_  & \new_[83987]_ ;
  assign \new_[83999]_  = ~A236 & ~A235;
  assign \new_[84000]_  = ~A233 & \new_[83999]_ ;
  assign \new_[84003]_  = A266 & A265;
  assign \new_[84006]_  = A299 & A298;
  assign \new_[84007]_  = \new_[84006]_  & \new_[84003]_ ;
  assign \new_[84008]_  = \new_[84007]_  & \new_[84000]_ ;
  assign \new_[84012]_  = ~A167 & ~A169;
  assign \new_[84013]_  = A170 & \new_[84012]_ ;
  assign \new_[84016]_  = ~A200 & A166;
  assign \new_[84019]_  = ~A203 & ~A202;
  assign \new_[84020]_  = \new_[84019]_  & \new_[84016]_ ;
  assign \new_[84021]_  = \new_[84020]_  & \new_[84013]_ ;
  assign \new_[84025]_  = ~A236 & ~A235;
  assign \new_[84026]_  = ~A233 & \new_[84025]_ ;
  assign \new_[84029]_  = A266 & A265;
  assign \new_[84032]_  = ~A299 & ~A298;
  assign \new_[84033]_  = \new_[84032]_  & \new_[84029]_ ;
  assign \new_[84034]_  = \new_[84033]_  & \new_[84026]_ ;
  assign \new_[84038]_  = ~A167 & ~A169;
  assign \new_[84039]_  = A170 & \new_[84038]_ ;
  assign \new_[84042]_  = ~A200 & A166;
  assign \new_[84045]_  = ~A203 & ~A202;
  assign \new_[84046]_  = \new_[84045]_  & \new_[84042]_ ;
  assign \new_[84047]_  = \new_[84046]_  & \new_[84039]_ ;
  assign \new_[84051]_  = ~A236 & ~A235;
  assign \new_[84052]_  = ~A233 & \new_[84051]_ ;
  assign \new_[84055]_  = ~A267 & ~A266;
  assign \new_[84058]_  = ~A300 & A298;
  assign \new_[84059]_  = \new_[84058]_  & \new_[84055]_ ;
  assign \new_[84060]_  = \new_[84059]_  & \new_[84052]_ ;
  assign \new_[84064]_  = ~A167 & ~A169;
  assign \new_[84065]_  = A170 & \new_[84064]_ ;
  assign \new_[84068]_  = ~A200 & A166;
  assign \new_[84071]_  = ~A203 & ~A202;
  assign \new_[84072]_  = \new_[84071]_  & \new_[84068]_ ;
  assign \new_[84073]_  = \new_[84072]_  & \new_[84065]_ ;
  assign \new_[84077]_  = ~A236 & ~A235;
  assign \new_[84078]_  = ~A233 & \new_[84077]_ ;
  assign \new_[84081]_  = ~A267 & ~A266;
  assign \new_[84084]_  = A299 & A298;
  assign \new_[84085]_  = \new_[84084]_  & \new_[84081]_ ;
  assign \new_[84086]_  = \new_[84085]_  & \new_[84078]_ ;
  assign \new_[84090]_  = ~A167 & ~A169;
  assign \new_[84091]_  = A170 & \new_[84090]_ ;
  assign \new_[84094]_  = ~A200 & A166;
  assign \new_[84097]_  = ~A203 & ~A202;
  assign \new_[84098]_  = \new_[84097]_  & \new_[84094]_ ;
  assign \new_[84099]_  = \new_[84098]_  & \new_[84091]_ ;
  assign \new_[84103]_  = ~A236 & ~A235;
  assign \new_[84104]_  = ~A233 & \new_[84103]_ ;
  assign \new_[84107]_  = ~A267 & ~A266;
  assign \new_[84110]_  = ~A299 & ~A298;
  assign \new_[84111]_  = \new_[84110]_  & \new_[84107]_ ;
  assign \new_[84112]_  = \new_[84111]_  & \new_[84104]_ ;
  assign \new_[84116]_  = ~A167 & ~A169;
  assign \new_[84117]_  = A170 & \new_[84116]_ ;
  assign \new_[84120]_  = ~A200 & A166;
  assign \new_[84123]_  = ~A203 & ~A202;
  assign \new_[84124]_  = \new_[84123]_  & \new_[84120]_ ;
  assign \new_[84125]_  = \new_[84124]_  & \new_[84117]_ ;
  assign \new_[84129]_  = ~A236 & ~A235;
  assign \new_[84130]_  = ~A233 & \new_[84129]_ ;
  assign \new_[84133]_  = ~A266 & ~A265;
  assign \new_[84136]_  = ~A300 & A298;
  assign \new_[84137]_  = \new_[84136]_  & \new_[84133]_ ;
  assign \new_[84138]_  = \new_[84137]_  & \new_[84130]_ ;
  assign \new_[84142]_  = ~A167 & ~A169;
  assign \new_[84143]_  = A170 & \new_[84142]_ ;
  assign \new_[84146]_  = ~A200 & A166;
  assign \new_[84149]_  = ~A203 & ~A202;
  assign \new_[84150]_  = \new_[84149]_  & \new_[84146]_ ;
  assign \new_[84151]_  = \new_[84150]_  & \new_[84143]_ ;
  assign \new_[84155]_  = ~A236 & ~A235;
  assign \new_[84156]_  = ~A233 & \new_[84155]_ ;
  assign \new_[84159]_  = ~A266 & ~A265;
  assign \new_[84162]_  = A299 & A298;
  assign \new_[84163]_  = \new_[84162]_  & \new_[84159]_ ;
  assign \new_[84164]_  = \new_[84163]_  & \new_[84156]_ ;
  assign \new_[84168]_  = ~A167 & ~A169;
  assign \new_[84169]_  = A170 & \new_[84168]_ ;
  assign \new_[84172]_  = ~A200 & A166;
  assign \new_[84175]_  = ~A203 & ~A202;
  assign \new_[84176]_  = \new_[84175]_  & \new_[84172]_ ;
  assign \new_[84177]_  = \new_[84176]_  & \new_[84169]_ ;
  assign \new_[84181]_  = ~A236 & ~A235;
  assign \new_[84182]_  = ~A233 & \new_[84181]_ ;
  assign \new_[84185]_  = ~A266 & ~A265;
  assign \new_[84188]_  = ~A299 & ~A298;
  assign \new_[84189]_  = \new_[84188]_  & \new_[84185]_ ;
  assign \new_[84190]_  = \new_[84189]_  & \new_[84182]_ ;
  assign \new_[84194]_  = ~A167 & ~A169;
  assign \new_[84195]_  = A170 & \new_[84194]_ ;
  assign \new_[84198]_  = ~A200 & A166;
  assign \new_[84201]_  = ~A203 & ~A202;
  assign \new_[84202]_  = \new_[84201]_  & \new_[84198]_ ;
  assign \new_[84203]_  = \new_[84202]_  & \new_[84195]_ ;
  assign \new_[84207]_  = A265 & ~A234;
  assign \new_[84208]_  = ~A233 & \new_[84207]_ ;
  assign \new_[84211]_  = A298 & A266;
  assign \new_[84214]_  = ~A302 & ~A301;
  assign \new_[84215]_  = \new_[84214]_  & \new_[84211]_ ;
  assign \new_[84216]_  = \new_[84215]_  & \new_[84208]_ ;
  assign \new_[84220]_  = ~A167 & ~A169;
  assign \new_[84221]_  = A170 & \new_[84220]_ ;
  assign \new_[84224]_  = ~A200 & A166;
  assign \new_[84227]_  = ~A203 & ~A202;
  assign \new_[84228]_  = \new_[84227]_  & \new_[84224]_ ;
  assign \new_[84229]_  = \new_[84228]_  & \new_[84221]_ ;
  assign \new_[84233]_  = ~A266 & ~A234;
  assign \new_[84234]_  = ~A233 & \new_[84233]_ ;
  assign \new_[84237]_  = ~A269 & ~A268;
  assign \new_[84240]_  = ~A300 & A298;
  assign \new_[84241]_  = \new_[84240]_  & \new_[84237]_ ;
  assign \new_[84242]_  = \new_[84241]_  & \new_[84234]_ ;
  assign \new_[84246]_  = ~A167 & ~A169;
  assign \new_[84247]_  = A170 & \new_[84246]_ ;
  assign \new_[84250]_  = ~A200 & A166;
  assign \new_[84253]_  = ~A203 & ~A202;
  assign \new_[84254]_  = \new_[84253]_  & \new_[84250]_ ;
  assign \new_[84255]_  = \new_[84254]_  & \new_[84247]_ ;
  assign \new_[84259]_  = ~A266 & ~A234;
  assign \new_[84260]_  = ~A233 & \new_[84259]_ ;
  assign \new_[84263]_  = ~A269 & ~A268;
  assign \new_[84266]_  = A299 & A298;
  assign \new_[84267]_  = \new_[84266]_  & \new_[84263]_ ;
  assign \new_[84268]_  = \new_[84267]_  & \new_[84260]_ ;
  assign \new_[84272]_  = ~A167 & ~A169;
  assign \new_[84273]_  = A170 & \new_[84272]_ ;
  assign \new_[84276]_  = ~A200 & A166;
  assign \new_[84279]_  = ~A203 & ~A202;
  assign \new_[84280]_  = \new_[84279]_  & \new_[84276]_ ;
  assign \new_[84281]_  = \new_[84280]_  & \new_[84273]_ ;
  assign \new_[84285]_  = ~A266 & ~A234;
  assign \new_[84286]_  = ~A233 & \new_[84285]_ ;
  assign \new_[84289]_  = ~A269 & ~A268;
  assign \new_[84292]_  = ~A299 & ~A298;
  assign \new_[84293]_  = \new_[84292]_  & \new_[84289]_ ;
  assign \new_[84294]_  = \new_[84293]_  & \new_[84286]_ ;
  assign \new_[84298]_  = ~A167 & ~A169;
  assign \new_[84299]_  = A170 & \new_[84298]_ ;
  assign \new_[84302]_  = ~A200 & A166;
  assign \new_[84305]_  = ~A203 & ~A202;
  assign \new_[84306]_  = \new_[84305]_  & \new_[84302]_ ;
  assign \new_[84307]_  = \new_[84306]_  & \new_[84299]_ ;
  assign \new_[84311]_  = ~A266 & ~A234;
  assign \new_[84312]_  = ~A233 & \new_[84311]_ ;
  assign \new_[84315]_  = A298 & ~A267;
  assign \new_[84318]_  = ~A302 & ~A301;
  assign \new_[84319]_  = \new_[84318]_  & \new_[84315]_ ;
  assign \new_[84320]_  = \new_[84319]_  & \new_[84312]_ ;
  assign \new_[84324]_  = ~A167 & ~A169;
  assign \new_[84325]_  = A170 & \new_[84324]_ ;
  assign \new_[84328]_  = ~A200 & A166;
  assign \new_[84331]_  = ~A203 & ~A202;
  assign \new_[84332]_  = \new_[84331]_  & \new_[84328]_ ;
  assign \new_[84333]_  = \new_[84332]_  & \new_[84325]_ ;
  assign \new_[84337]_  = ~A265 & ~A234;
  assign \new_[84338]_  = ~A233 & \new_[84337]_ ;
  assign \new_[84341]_  = A298 & ~A266;
  assign \new_[84344]_  = ~A302 & ~A301;
  assign \new_[84345]_  = \new_[84344]_  & \new_[84341]_ ;
  assign \new_[84346]_  = \new_[84345]_  & \new_[84338]_ ;
  assign \new_[84350]_  = ~A167 & ~A169;
  assign \new_[84351]_  = A170 & \new_[84350]_ ;
  assign \new_[84354]_  = ~A200 & A166;
  assign \new_[84357]_  = ~A203 & ~A202;
  assign \new_[84358]_  = \new_[84357]_  & \new_[84354]_ ;
  assign \new_[84359]_  = \new_[84358]_  & \new_[84351]_ ;
  assign \new_[84363]_  = A265 & ~A233;
  assign \new_[84364]_  = ~A232 & \new_[84363]_ ;
  assign \new_[84367]_  = A298 & A266;
  assign \new_[84370]_  = ~A302 & ~A301;
  assign \new_[84371]_  = \new_[84370]_  & \new_[84367]_ ;
  assign \new_[84372]_  = \new_[84371]_  & \new_[84364]_ ;
  assign \new_[84376]_  = ~A167 & ~A169;
  assign \new_[84377]_  = A170 & \new_[84376]_ ;
  assign \new_[84380]_  = ~A200 & A166;
  assign \new_[84383]_  = ~A203 & ~A202;
  assign \new_[84384]_  = \new_[84383]_  & \new_[84380]_ ;
  assign \new_[84385]_  = \new_[84384]_  & \new_[84377]_ ;
  assign \new_[84389]_  = ~A266 & ~A233;
  assign \new_[84390]_  = ~A232 & \new_[84389]_ ;
  assign \new_[84393]_  = ~A269 & ~A268;
  assign \new_[84396]_  = ~A300 & A298;
  assign \new_[84397]_  = \new_[84396]_  & \new_[84393]_ ;
  assign \new_[84398]_  = \new_[84397]_  & \new_[84390]_ ;
  assign \new_[84402]_  = ~A167 & ~A169;
  assign \new_[84403]_  = A170 & \new_[84402]_ ;
  assign \new_[84406]_  = ~A200 & A166;
  assign \new_[84409]_  = ~A203 & ~A202;
  assign \new_[84410]_  = \new_[84409]_  & \new_[84406]_ ;
  assign \new_[84411]_  = \new_[84410]_  & \new_[84403]_ ;
  assign \new_[84415]_  = ~A266 & ~A233;
  assign \new_[84416]_  = ~A232 & \new_[84415]_ ;
  assign \new_[84419]_  = ~A269 & ~A268;
  assign \new_[84422]_  = A299 & A298;
  assign \new_[84423]_  = \new_[84422]_  & \new_[84419]_ ;
  assign \new_[84424]_  = \new_[84423]_  & \new_[84416]_ ;
  assign \new_[84428]_  = ~A167 & ~A169;
  assign \new_[84429]_  = A170 & \new_[84428]_ ;
  assign \new_[84432]_  = ~A200 & A166;
  assign \new_[84435]_  = ~A203 & ~A202;
  assign \new_[84436]_  = \new_[84435]_  & \new_[84432]_ ;
  assign \new_[84437]_  = \new_[84436]_  & \new_[84429]_ ;
  assign \new_[84441]_  = ~A266 & ~A233;
  assign \new_[84442]_  = ~A232 & \new_[84441]_ ;
  assign \new_[84445]_  = ~A269 & ~A268;
  assign \new_[84448]_  = ~A299 & ~A298;
  assign \new_[84449]_  = \new_[84448]_  & \new_[84445]_ ;
  assign \new_[84450]_  = \new_[84449]_  & \new_[84442]_ ;
  assign \new_[84454]_  = ~A167 & ~A169;
  assign \new_[84455]_  = A170 & \new_[84454]_ ;
  assign \new_[84458]_  = ~A200 & A166;
  assign \new_[84461]_  = ~A203 & ~A202;
  assign \new_[84462]_  = \new_[84461]_  & \new_[84458]_ ;
  assign \new_[84463]_  = \new_[84462]_  & \new_[84455]_ ;
  assign \new_[84467]_  = ~A266 & ~A233;
  assign \new_[84468]_  = ~A232 & \new_[84467]_ ;
  assign \new_[84471]_  = A298 & ~A267;
  assign \new_[84474]_  = ~A302 & ~A301;
  assign \new_[84475]_  = \new_[84474]_  & \new_[84471]_ ;
  assign \new_[84476]_  = \new_[84475]_  & \new_[84468]_ ;
  assign \new_[84480]_  = ~A167 & ~A169;
  assign \new_[84481]_  = A170 & \new_[84480]_ ;
  assign \new_[84484]_  = ~A200 & A166;
  assign \new_[84487]_  = ~A203 & ~A202;
  assign \new_[84488]_  = \new_[84487]_  & \new_[84484]_ ;
  assign \new_[84489]_  = \new_[84488]_  & \new_[84481]_ ;
  assign \new_[84493]_  = ~A265 & ~A233;
  assign \new_[84494]_  = ~A232 & \new_[84493]_ ;
  assign \new_[84497]_  = A298 & ~A266;
  assign \new_[84500]_  = ~A302 & ~A301;
  assign \new_[84501]_  = \new_[84500]_  & \new_[84497]_ ;
  assign \new_[84502]_  = \new_[84501]_  & \new_[84494]_ ;
  assign \new_[84506]_  = ~A167 & ~A169;
  assign \new_[84507]_  = A170 & \new_[84506]_ ;
  assign \new_[84510]_  = ~A200 & A166;
  assign \new_[84513]_  = A232 & ~A201;
  assign \new_[84514]_  = \new_[84513]_  & \new_[84510]_ ;
  assign \new_[84515]_  = \new_[84514]_  & \new_[84507]_ ;
  assign \new_[84519]_  = ~A268 & A265;
  assign \new_[84520]_  = A233 & \new_[84519]_ ;
  assign \new_[84523]_  = ~A299 & ~A269;
  assign \new_[84526]_  = ~A302 & ~A301;
  assign \new_[84527]_  = \new_[84526]_  & \new_[84523]_ ;
  assign \new_[84528]_  = \new_[84527]_  & \new_[84520]_ ;
  assign \new_[84532]_  = ~A167 & ~A169;
  assign \new_[84533]_  = A170 & \new_[84532]_ ;
  assign \new_[84536]_  = ~A200 & A166;
  assign \new_[84539]_  = ~A233 & ~A201;
  assign \new_[84540]_  = \new_[84539]_  & \new_[84536]_ ;
  assign \new_[84541]_  = \new_[84540]_  & \new_[84533]_ ;
  assign \new_[84545]_  = A265 & ~A236;
  assign \new_[84546]_  = ~A235 & \new_[84545]_ ;
  assign \new_[84549]_  = A298 & A266;
  assign \new_[84552]_  = ~A302 & ~A301;
  assign \new_[84553]_  = \new_[84552]_  & \new_[84549]_ ;
  assign \new_[84554]_  = \new_[84553]_  & \new_[84546]_ ;
  assign \new_[84558]_  = ~A167 & ~A169;
  assign \new_[84559]_  = A170 & \new_[84558]_ ;
  assign \new_[84562]_  = ~A200 & A166;
  assign \new_[84565]_  = ~A233 & ~A201;
  assign \new_[84566]_  = \new_[84565]_  & \new_[84562]_ ;
  assign \new_[84567]_  = \new_[84566]_  & \new_[84559]_ ;
  assign \new_[84571]_  = ~A266 & ~A236;
  assign \new_[84572]_  = ~A235 & \new_[84571]_ ;
  assign \new_[84575]_  = ~A269 & ~A268;
  assign \new_[84578]_  = ~A300 & A298;
  assign \new_[84579]_  = \new_[84578]_  & \new_[84575]_ ;
  assign \new_[84580]_  = \new_[84579]_  & \new_[84572]_ ;
  assign \new_[84584]_  = ~A167 & ~A169;
  assign \new_[84585]_  = A170 & \new_[84584]_ ;
  assign \new_[84588]_  = ~A200 & A166;
  assign \new_[84591]_  = ~A233 & ~A201;
  assign \new_[84592]_  = \new_[84591]_  & \new_[84588]_ ;
  assign \new_[84593]_  = \new_[84592]_  & \new_[84585]_ ;
  assign \new_[84597]_  = ~A266 & ~A236;
  assign \new_[84598]_  = ~A235 & \new_[84597]_ ;
  assign \new_[84601]_  = ~A269 & ~A268;
  assign \new_[84604]_  = A299 & A298;
  assign \new_[84605]_  = \new_[84604]_  & \new_[84601]_ ;
  assign \new_[84606]_  = \new_[84605]_  & \new_[84598]_ ;
  assign \new_[84610]_  = ~A167 & ~A169;
  assign \new_[84611]_  = A170 & \new_[84610]_ ;
  assign \new_[84614]_  = ~A200 & A166;
  assign \new_[84617]_  = ~A233 & ~A201;
  assign \new_[84618]_  = \new_[84617]_  & \new_[84614]_ ;
  assign \new_[84619]_  = \new_[84618]_  & \new_[84611]_ ;
  assign \new_[84623]_  = ~A266 & ~A236;
  assign \new_[84624]_  = ~A235 & \new_[84623]_ ;
  assign \new_[84627]_  = ~A269 & ~A268;
  assign \new_[84630]_  = ~A299 & ~A298;
  assign \new_[84631]_  = \new_[84630]_  & \new_[84627]_ ;
  assign \new_[84632]_  = \new_[84631]_  & \new_[84624]_ ;
  assign \new_[84636]_  = ~A167 & ~A169;
  assign \new_[84637]_  = A170 & \new_[84636]_ ;
  assign \new_[84640]_  = ~A200 & A166;
  assign \new_[84643]_  = ~A233 & ~A201;
  assign \new_[84644]_  = \new_[84643]_  & \new_[84640]_ ;
  assign \new_[84645]_  = \new_[84644]_  & \new_[84637]_ ;
  assign \new_[84649]_  = ~A266 & ~A236;
  assign \new_[84650]_  = ~A235 & \new_[84649]_ ;
  assign \new_[84653]_  = A298 & ~A267;
  assign \new_[84656]_  = ~A302 & ~A301;
  assign \new_[84657]_  = \new_[84656]_  & \new_[84653]_ ;
  assign \new_[84658]_  = \new_[84657]_  & \new_[84650]_ ;
  assign \new_[84662]_  = ~A167 & ~A169;
  assign \new_[84663]_  = A170 & \new_[84662]_ ;
  assign \new_[84666]_  = ~A200 & A166;
  assign \new_[84669]_  = ~A233 & ~A201;
  assign \new_[84670]_  = \new_[84669]_  & \new_[84666]_ ;
  assign \new_[84671]_  = \new_[84670]_  & \new_[84663]_ ;
  assign \new_[84675]_  = ~A265 & ~A236;
  assign \new_[84676]_  = ~A235 & \new_[84675]_ ;
  assign \new_[84679]_  = A298 & ~A266;
  assign \new_[84682]_  = ~A302 & ~A301;
  assign \new_[84683]_  = \new_[84682]_  & \new_[84679]_ ;
  assign \new_[84684]_  = \new_[84683]_  & \new_[84676]_ ;
  assign \new_[84688]_  = ~A167 & ~A169;
  assign \new_[84689]_  = A170 & \new_[84688]_ ;
  assign \new_[84692]_  = ~A200 & A166;
  assign \new_[84695]_  = ~A233 & ~A201;
  assign \new_[84696]_  = \new_[84695]_  & \new_[84692]_ ;
  assign \new_[84697]_  = \new_[84696]_  & \new_[84689]_ ;
  assign \new_[84701]_  = ~A268 & ~A266;
  assign \new_[84702]_  = ~A234 & \new_[84701]_ ;
  assign \new_[84705]_  = A298 & ~A269;
  assign \new_[84708]_  = ~A302 & ~A301;
  assign \new_[84709]_  = \new_[84708]_  & \new_[84705]_ ;
  assign \new_[84710]_  = \new_[84709]_  & \new_[84702]_ ;
  assign \new_[84714]_  = ~A167 & ~A169;
  assign \new_[84715]_  = A170 & \new_[84714]_ ;
  assign \new_[84718]_  = ~A200 & A166;
  assign \new_[84721]_  = A232 & ~A201;
  assign \new_[84722]_  = \new_[84721]_  & \new_[84718]_ ;
  assign \new_[84723]_  = \new_[84722]_  & \new_[84715]_ ;
  assign \new_[84727]_  = A235 & A234;
  assign \new_[84728]_  = ~A233 & \new_[84727]_ ;
  assign \new_[84731]_  = ~A299 & A298;
  assign \new_[84734]_  = A301 & A300;
  assign \new_[84735]_  = \new_[84734]_  & \new_[84731]_ ;
  assign \new_[84736]_  = \new_[84735]_  & \new_[84728]_ ;
  assign \new_[84740]_  = ~A167 & ~A169;
  assign \new_[84741]_  = A170 & \new_[84740]_ ;
  assign \new_[84744]_  = ~A200 & A166;
  assign \new_[84747]_  = A232 & ~A201;
  assign \new_[84748]_  = \new_[84747]_  & \new_[84744]_ ;
  assign \new_[84749]_  = \new_[84748]_  & \new_[84741]_ ;
  assign \new_[84753]_  = A235 & A234;
  assign \new_[84754]_  = ~A233 & \new_[84753]_ ;
  assign \new_[84757]_  = ~A299 & A298;
  assign \new_[84760]_  = A302 & A300;
  assign \new_[84761]_  = \new_[84760]_  & \new_[84757]_ ;
  assign \new_[84762]_  = \new_[84761]_  & \new_[84754]_ ;
  assign \new_[84766]_  = ~A167 & ~A169;
  assign \new_[84767]_  = A170 & \new_[84766]_ ;
  assign \new_[84770]_  = ~A200 & A166;
  assign \new_[84773]_  = A232 & ~A201;
  assign \new_[84774]_  = \new_[84773]_  & \new_[84770]_ ;
  assign \new_[84775]_  = \new_[84774]_  & \new_[84767]_ ;
  assign \new_[84779]_  = A235 & A234;
  assign \new_[84780]_  = ~A233 & \new_[84779]_ ;
  assign \new_[84783]_  = ~A266 & A265;
  assign \new_[84786]_  = A268 & A267;
  assign \new_[84787]_  = \new_[84786]_  & \new_[84783]_ ;
  assign \new_[84788]_  = \new_[84787]_  & \new_[84780]_ ;
  assign \new_[84792]_  = ~A167 & ~A169;
  assign \new_[84793]_  = A170 & \new_[84792]_ ;
  assign \new_[84796]_  = ~A200 & A166;
  assign \new_[84799]_  = A232 & ~A201;
  assign \new_[84800]_  = \new_[84799]_  & \new_[84796]_ ;
  assign \new_[84801]_  = \new_[84800]_  & \new_[84793]_ ;
  assign \new_[84805]_  = A235 & A234;
  assign \new_[84806]_  = ~A233 & \new_[84805]_ ;
  assign \new_[84809]_  = ~A266 & A265;
  assign \new_[84812]_  = A269 & A267;
  assign \new_[84813]_  = \new_[84812]_  & \new_[84809]_ ;
  assign \new_[84814]_  = \new_[84813]_  & \new_[84806]_ ;
  assign \new_[84818]_  = ~A167 & ~A169;
  assign \new_[84819]_  = A170 & \new_[84818]_ ;
  assign \new_[84822]_  = ~A200 & A166;
  assign \new_[84825]_  = A232 & ~A201;
  assign \new_[84826]_  = \new_[84825]_  & \new_[84822]_ ;
  assign \new_[84827]_  = \new_[84826]_  & \new_[84819]_ ;
  assign \new_[84831]_  = A236 & A234;
  assign \new_[84832]_  = ~A233 & \new_[84831]_ ;
  assign \new_[84835]_  = ~A299 & A298;
  assign \new_[84838]_  = A301 & A300;
  assign \new_[84839]_  = \new_[84838]_  & \new_[84835]_ ;
  assign \new_[84840]_  = \new_[84839]_  & \new_[84832]_ ;
  assign \new_[84844]_  = ~A167 & ~A169;
  assign \new_[84845]_  = A170 & \new_[84844]_ ;
  assign \new_[84848]_  = ~A200 & A166;
  assign \new_[84851]_  = A232 & ~A201;
  assign \new_[84852]_  = \new_[84851]_  & \new_[84848]_ ;
  assign \new_[84853]_  = \new_[84852]_  & \new_[84845]_ ;
  assign \new_[84857]_  = A236 & A234;
  assign \new_[84858]_  = ~A233 & \new_[84857]_ ;
  assign \new_[84861]_  = ~A299 & A298;
  assign \new_[84864]_  = A302 & A300;
  assign \new_[84865]_  = \new_[84864]_  & \new_[84861]_ ;
  assign \new_[84866]_  = \new_[84865]_  & \new_[84858]_ ;
  assign \new_[84870]_  = ~A167 & ~A169;
  assign \new_[84871]_  = A170 & \new_[84870]_ ;
  assign \new_[84874]_  = ~A200 & A166;
  assign \new_[84877]_  = A232 & ~A201;
  assign \new_[84878]_  = \new_[84877]_  & \new_[84874]_ ;
  assign \new_[84879]_  = \new_[84878]_  & \new_[84871]_ ;
  assign \new_[84883]_  = A236 & A234;
  assign \new_[84884]_  = ~A233 & \new_[84883]_ ;
  assign \new_[84887]_  = ~A266 & A265;
  assign \new_[84890]_  = A268 & A267;
  assign \new_[84891]_  = \new_[84890]_  & \new_[84887]_ ;
  assign \new_[84892]_  = \new_[84891]_  & \new_[84884]_ ;
  assign \new_[84896]_  = ~A167 & ~A169;
  assign \new_[84897]_  = A170 & \new_[84896]_ ;
  assign \new_[84900]_  = ~A200 & A166;
  assign \new_[84903]_  = A232 & ~A201;
  assign \new_[84904]_  = \new_[84903]_  & \new_[84900]_ ;
  assign \new_[84905]_  = \new_[84904]_  & \new_[84897]_ ;
  assign \new_[84909]_  = A236 & A234;
  assign \new_[84910]_  = ~A233 & \new_[84909]_ ;
  assign \new_[84913]_  = ~A266 & A265;
  assign \new_[84916]_  = A269 & A267;
  assign \new_[84917]_  = \new_[84916]_  & \new_[84913]_ ;
  assign \new_[84918]_  = \new_[84917]_  & \new_[84910]_ ;
  assign \new_[84922]_  = ~A167 & ~A169;
  assign \new_[84923]_  = A170 & \new_[84922]_ ;
  assign \new_[84926]_  = ~A200 & A166;
  assign \new_[84929]_  = ~A232 & ~A201;
  assign \new_[84930]_  = \new_[84929]_  & \new_[84926]_ ;
  assign \new_[84931]_  = \new_[84930]_  & \new_[84923]_ ;
  assign \new_[84935]_  = ~A268 & ~A266;
  assign \new_[84936]_  = ~A233 & \new_[84935]_ ;
  assign \new_[84939]_  = A298 & ~A269;
  assign \new_[84942]_  = ~A302 & ~A301;
  assign \new_[84943]_  = \new_[84942]_  & \new_[84939]_ ;
  assign \new_[84944]_  = \new_[84943]_  & \new_[84936]_ ;
  assign \new_[84948]_  = ~A167 & ~A169;
  assign \new_[84949]_  = A170 & \new_[84948]_ ;
  assign \new_[84952]_  = ~A199 & A166;
  assign \new_[84955]_  = A232 & ~A200;
  assign \new_[84956]_  = \new_[84955]_  & \new_[84952]_ ;
  assign \new_[84957]_  = \new_[84956]_  & \new_[84949]_ ;
  assign \new_[84961]_  = ~A268 & A265;
  assign \new_[84962]_  = A233 & \new_[84961]_ ;
  assign \new_[84965]_  = ~A299 & ~A269;
  assign \new_[84968]_  = ~A302 & ~A301;
  assign \new_[84969]_  = \new_[84968]_  & \new_[84965]_ ;
  assign \new_[84970]_  = \new_[84969]_  & \new_[84962]_ ;
  assign \new_[84974]_  = ~A167 & ~A169;
  assign \new_[84975]_  = A170 & \new_[84974]_ ;
  assign \new_[84978]_  = ~A199 & A166;
  assign \new_[84981]_  = ~A233 & ~A200;
  assign \new_[84982]_  = \new_[84981]_  & \new_[84978]_ ;
  assign \new_[84983]_  = \new_[84982]_  & \new_[84975]_ ;
  assign \new_[84987]_  = A265 & ~A236;
  assign \new_[84988]_  = ~A235 & \new_[84987]_ ;
  assign \new_[84991]_  = A298 & A266;
  assign \new_[84994]_  = ~A302 & ~A301;
  assign \new_[84995]_  = \new_[84994]_  & \new_[84991]_ ;
  assign \new_[84996]_  = \new_[84995]_  & \new_[84988]_ ;
  assign \new_[85000]_  = ~A167 & ~A169;
  assign \new_[85001]_  = A170 & \new_[85000]_ ;
  assign \new_[85004]_  = ~A199 & A166;
  assign \new_[85007]_  = ~A233 & ~A200;
  assign \new_[85008]_  = \new_[85007]_  & \new_[85004]_ ;
  assign \new_[85009]_  = \new_[85008]_  & \new_[85001]_ ;
  assign \new_[85013]_  = ~A266 & ~A236;
  assign \new_[85014]_  = ~A235 & \new_[85013]_ ;
  assign \new_[85017]_  = ~A269 & ~A268;
  assign \new_[85020]_  = ~A300 & A298;
  assign \new_[85021]_  = \new_[85020]_  & \new_[85017]_ ;
  assign \new_[85022]_  = \new_[85021]_  & \new_[85014]_ ;
  assign \new_[85026]_  = ~A167 & ~A169;
  assign \new_[85027]_  = A170 & \new_[85026]_ ;
  assign \new_[85030]_  = ~A199 & A166;
  assign \new_[85033]_  = ~A233 & ~A200;
  assign \new_[85034]_  = \new_[85033]_  & \new_[85030]_ ;
  assign \new_[85035]_  = \new_[85034]_  & \new_[85027]_ ;
  assign \new_[85039]_  = ~A266 & ~A236;
  assign \new_[85040]_  = ~A235 & \new_[85039]_ ;
  assign \new_[85043]_  = ~A269 & ~A268;
  assign \new_[85046]_  = A299 & A298;
  assign \new_[85047]_  = \new_[85046]_  & \new_[85043]_ ;
  assign \new_[85048]_  = \new_[85047]_  & \new_[85040]_ ;
  assign \new_[85052]_  = ~A167 & ~A169;
  assign \new_[85053]_  = A170 & \new_[85052]_ ;
  assign \new_[85056]_  = ~A199 & A166;
  assign \new_[85059]_  = ~A233 & ~A200;
  assign \new_[85060]_  = \new_[85059]_  & \new_[85056]_ ;
  assign \new_[85061]_  = \new_[85060]_  & \new_[85053]_ ;
  assign \new_[85065]_  = ~A266 & ~A236;
  assign \new_[85066]_  = ~A235 & \new_[85065]_ ;
  assign \new_[85069]_  = ~A269 & ~A268;
  assign \new_[85072]_  = ~A299 & ~A298;
  assign \new_[85073]_  = \new_[85072]_  & \new_[85069]_ ;
  assign \new_[85074]_  = \new_[85073]_  & \new_[85066]_ ;
  assign \new_[85078]_  = ~A167 & ~A169;
  assign \new_[85079]_  = A170 & \new_[85078]_ ;
  assign \new_[85082]_  = ~A199 & A166;
  assign \new_[85085]_  = ~A233 & ~A200;
  assign \new_[85086]_  = \new_[85085]_  & \new_[85082]_ ;
  assign \new_[85087]_  = \new_[85086]_  & \new_[85079]_ ;
  assign \new_[85091]_  = ~A266 & ~A236;
  assign \new_[85092]_  = ~A235 & \new_[85091]_ ;
  assign \new_[85095]_  = A298 & ~A267;
  assign \new_[85098]_  = ~A302 & ~A301;
  assign \new_[85099]_  = \new_[85098]_  & \new_[85095]_ ;
  assign \new_[85100]_  = \new_[85099]_  & \new_[85092]_ ;
  assign \new_[85104]_  = ~A167 & ~A169;
  assign \new_[85105]_  = A170 & \new_[85104]_ ;
  assign \new_[85108]_  = ~A199 & A166;
  assign \new_[85111]_  = ~A233 & ~A200;
  assign \new_[85112]_  = \new_[85111]_  & \new_[85108]_ ;
  assign \new_[85113]_  = \new_[85112]_  & \new_[85105]_ ;
  assign \new_[85117]_  = ~A265 & ~A236;
  assign \new_[85118]_  = ~A235 & \new_[85117]_ ;
  assign \new_[85121]_  = A298 & ~A266;
  assign \new_[85124]_  = ~A302 & ~A301;
  assign \new_[85125]_  = \new_[85124]_  & \new_[85121]_ ;
  assign \new_[85126]_  = \new_[85125]_  & \new_[85118]_ ;
  assign \new_[85130]_  = ~A167 & ~A169;
  assign \new_[85131]_  = A170 & \new_[85130]_ ;
  assign \new_[85134]_  = ~A199 & A166;
  assign \new_[85137]_  = ~A233 & ~A200;
  assign \new_[85138]_  = \new_[85137]_  & \new_[85134]_ ;
  assign \new_[85139]_  = \new_[85138]_  & \new_[85131]_ ;
  assign \new_[85143]_  = ~A268 & ~A266;
  assign \new_[85144]_  = ~A234 & \new_[85143]_ ;
  assign \new_[85147]_  = A298 & ~A269;
  assign \new_[85150]_  = ~A302 & ~A301;
  assign \new_[85151]_  = \new_[85150]_  & \new_[85147]_ ;
  assign \new_[85152]_  = \new_[85151]_  & \new_[85144]_ ;
  assign \new_[85156]_  = ~A167 & ~A169;
  assign \new_[85157]_  = A170 & \new_[85156]_ ;
  assign \new_[85160]_  = ~A199 & A166;
  assign \new_[85163]_  = A232 & ~A200;
  assign \new_[85164]_  = \new_[85163]_  & \new_[85160]_ ;
  assign \new_[85165]_  = \new_[85164]_  & \new_[85157]_ ;
  assign \new_[85169]_  = A235 & A234;
  assign \new_[85170]_  = ~A233 & \new_[85169]_ ;
  assign \new_[85173]_  = ~A299 & A298;
  assign \new_[85176]_  = A301 & A300;
  assign \new_[85177]_  = \new_[85176]_  & \new_[85173]_ ;
  assign \new_[85178]_  = \new_[85177]_  & \new_[85170]_ ;
  assign \new_[85182]_  = ~A167 & ~A169;
  assign \new_[85183]_  = A170 & \new_[85182]_ ;
  assign \new_[85186]_  = ~A199 & A166;
  assign \new_[85189]_  = A232 & ~A200;
  assign \new_[85190]_  = \new_[85189]_  & \new_[85186]_ ;
  assign \new_[85191]_  = \new_[85190]_  & \new_[85183]_ ;
  assign \new_[85195]_  = A235 & A234;
  assign \new_[85196]_  = ~A233 & \new_[85195]_ ;
  assign \new_[85199]_  = ~A299 & A298;
  assign \new_[85202]_  = A302 & A300;
  assign \new_[85203]_  = \new_[85202]_  & \new_[85199]_ ;
  assign \new_[85204]_  = \new_[85203]_  & \new_[85196]_ ;
  assign \new_[85208]_  = ~A167 & ~A169;
  assign \new_[85209]_  = A170 & \new_[85208]_ ;
  assign \new_[85212]_  = ~A199 & A166;
  assign \new_[85215]_  = A232 & ~A200;
  assign \new_[85216]_  = \new_[85215]_  & \new_[85212]_ ;
  assign \new_[85217]_  = \new_[85216]_  & \new_[85209]_ ;
  assign \new_[85221]_  = A235 & A234;
  assign \new_[85222]_  = ~A233 & \new_[85221]_ ;
  assign \new_[85225]_  = ~A266 & A265;
  assign \new_[85228]_  = A268 & A267;
  assign \new_[85229]_  = \new_[85228]_  & \new_[85225]_ ;
  assign \new_[85230]_  = \new_[85229]_  & \new_[85222]_ ;
  assign \new_[85234]_  = ~A167 & ~A169;
  assign \new_[85235]_  = A170 & \new_[85234]_ ;
  assign \new_[85238]_  = ~A199 & A166;
  assign \new_[85241]_  = A232 & ~A200;
  assign \new_[85242]_  = \new_[85241]_  & \new_[85238]_ ;
  assign \new_[85243]_  = \new_[85242]_  & \new_[85235]_ ;
  assign \new_[85247]_  = A235 & A234;
  assign \new_[85248]_  = ~A233 & \new_[85247]_ ;
  assign \new_[85251]_  = ~A266 & A265;
  assign \new_[85254]_  = A269 & A267;
  assign \new_[85255]_  = \new_[85254]_  & \new_[85251]_ ;
  assign \new_[85256]_  = \new_[85255]_  & \new_[85248]_ ;
  assign \new_[85260]_  = ~A167 & ~A169;
  assign \new_[85261]_  = A170 & \new_[85260]_ ;
  assign \new_[85264]_  = ~A199 & A166;
  assign \new_[85267]_  = A232 & ~A200;
  assign \new_[85268]_  = \new_[85267]_  & \new_[85264]_ ;
  assign \new_[85269]_  = \new_[85268]_  & \new_[85261]_ ;
  assign \new_[85273]_  = A236 & A234;
  assign \new_[85274]_  = ~A233 & \new_[85273]_ ;
  assign \new_[85277]_  = ~A299 & A298;
  assign \new_[85280]_  = A301 & A300;
  assign \new_[85281]_  = \new_[85280]_  & \new_[85277]_ ;
  assign \new_[85282]_  = \new_[85281]_  & \new_[85274]_ ;
  assign \new_[85286]_  = ~A167 & ~A169;
  assign \new_[85287]_  = A170 & \new_[85286]_ ;
  assign \new_[85290]_  = ~A199 & A166;
  assign \new_[85293]_  = A232 & ~A200;
  assign \new_[85294]_  = \new_[85293]_  & \new_[85290]_ ;
  assign \new_[85295]_  = \new_[85294]_  & \new_[85287]_ ;
  assign \new_[85299]_  = A236 & A234;
  assign \new_[85300]_  = ~A233 & \new_[85299]_ ;
  assign \new_[85303]_  = ~A299 & A298;
  assign \new_[85306]_  = A302 & A300;
  assign \new_[85307]_  = \new_[85306]_  & \new_[85303]_ ;
  assign \new_[85308]_  = \new_[85307]_  & \new_[85300]_ ;
  assign \new_[85312]_  = ~A167 & ~A169;
  assign \new_[85313]_  = A170 & \new_[85312]_ ;
  assign \new_[85316]_  = ~A199 & A166;
  assign \new_[85319]_  = A232 & ~A200;
  assign \new_[85320]_  = \new_[85319]_  & \new_[85316]_ ;
  assign \new_[85321]_  = \new_[85320]_  & \new_[85313]_ ;
  assign \new_[85325]_  = A236 & A234;
  assign \new_[85326]_  = ~A233 & \new_[85325]_ ;
  assign \new_[85329]_  = ~A266 & A265;
  assign \new_[85332]_  = A268 & A267;
  assign \new_[85333]_  = \new_[85332]_  & \new_[85329]_ ;
  assign \new_[85334]_  = \new_[85333]_  & \new_[85326]_ ;
  assign \new_[85338]_  = ~A167 & ~A169;
  assign \new_[85339]_  = A170 & \new_[85338]_ ;
  assign \new_[85342]_  = ~A199 & A166;
  assign \new_[85345]_  = A232 & ~A200;
  assign \new_[85346]_  = \new_[85345]_  & \new_[85342]_ ;
  assign \new_[85347]_  = \new_[85346]_  & \new_[85339]_ ;
  assign \new_[85351]_  = A236 & A234;
  assign \new_[85352]_  = ~A233 & \new_[85351]_ ;
  assign \new_[85355]_  = ~A266 & A265;
  assign \new_[85358]_  = A269 & A267;
  assign \new_[85359]_  = \new_[85358]_  & \new_[85355]_ ;
  assign \new_[85360]_  = \new_[85359]_  & \new_[85352]_ ;
  assign \new_[85364]_  = ~A167 & ~A169;
  assign \new_[85365]_  = A170 & \new_[85364]_ ;
  assign \new_[85368]_  = ~A199 & A166;
  assign \new_[85371]_  = ~A232 & ~A200;
  assign \new_[85372]_  = \new_[85371]_  & \new_[85368]_ ;
  assign \new_[85373]_  = \new_[85372]_  & \new_[85365]_ ;
  assign \new_[85377]_  = ~A268 & ~A266;
  assign \new_[85378]_  = ~A233 & \new_[85377]_ ;
  assign \new_[85381]_  = A298 & ~A269;
  assign \new_[85384]_  = ~A302 & ~A301;
  assign \new_[85385]_  = \new_[85384]_  & \new_[85381]_ ;
  assign \new_[85386]_  = \new_[85385]_  & \new_[85378]_ ;
  assign \new_[85390]_  = ~A168 & ~A169;
  assign \new_[85391]_  = ~A170 & \new_[85390]_ ;
  assign \new_[85394]_  = ~A200 & A199;
  assign \new_[85397]_  = A202 & A201;
  assign \new_[85398]_  = \new_[85397]_  & \new_[85394]_ ;
  assign \new_[85399]_  = \new_[85398]_  & \new_[85391]_ ;
  assign \new_[85403]_  = A265 & A233;
  assign \new_[85404]_  = A232 & \new_[85403]_ ;
  assign \new_[85407]_  = ~A269 & ~A268;
  assign \new_[85410]_  = ~A300 & ~A299;
  assign \new_[85411]_  = \new_[85410]_  & \new_[85407]_ ;
  assign \new_[85412]_  = \new_[85411]_  & \new_[85404]_ ;
  assign \new_[85416]_  = ~A168 & ~A169;
  assign \new_[85417]_  = ~A170 & \new_[85416]_ ;
  assign \new_[85420]_  = ~A200 & A199;
  assign \new_[85423]_  = A202 & A201;
  assign \new_[85424]_  = \new_[85423]_  & \new_[85420]_ ;
  assign \new_[85425]_  = \new_[85424]_  & \new_[85417]_ ;
  assign \new_[85429]_  = A265 & A233;
  assign \new_[85430]_  = A232 & \new_[85429]_ ;
  assign \new_[85433]_  = ~A269 & ~A268;
  assign \new_[85436]_  = A299 & A298;
  assign \new_[85437]_  = \new_[85436]_  & \new_[85433]_ ;
  assign \new_[85438]_  = \new_[85437]_  & \new_[85430]_ ;
  assign \new_[85442]_  = ~A168 & ~A169;
  assign \new_[85443]_  = ~A170 & \new_[85442]_ ;
  assign \new_[85446]_  = ~A200 & A199;
  assign \new_[85449]_  = A202 & A201;
  assign \new_[85450]_  = \new_[85449]_  & \new_[85446]_ ;
  assign \new_[85451]_  = \new_[85450]_  & \new_[85443]_ ;
  assign \new_[85455]_  = A265 & A233;
  assign \new_[85456]_  = A232 & \new_[85455]_ ;
  assign \new_[85459]_  = ~A269 & ~A268;
  assign \new_[85462]_  = ~A299 & ~A298;
  assign \new_[85463]_  = \new_[85462]_  & \new_[85459]_ ;
  assign \new_[85464]_  = \new_[85463]_  & \new_[85456]_ ;
  assign \new_[85468]_  = ~A168 & ~A169;
  assign \new_[85469]_  = ~A170 & \new_[85468]_ ;
  assign \new_[85472]_  = ~A200 & A199;
  assign \new_[85475]_  = A202 & A201;
  assign \new_[85476]_  = \new_[85475]_  & \new_[85472]_ ;
  assign \new_[85477]_  = \new_[85476]_  & \new_[85469]_ ;
  assign \new_[85481]_  = A265 & A233;
  assign \new_[85482]_  = A232 & \new_[85481]_ ;
  assign \new_[85485]_  = ~A299 & ~A267;
  assign \new_[85488]_  = ~A302 & ~A301;
  assign \new_[85489]_  = \new_[85488]_  & \new_[85485]_ ;
  assign \new_[85490]_  = \new_[85489]_  & \new_[85482]_ ;
  assign \new_[85494]_  = ~A168 & ~A169;
  assign \new_[85495]_  = ~A170 & \new_[85494]_ ;
  assign \new_[85498]_  = ~A200 & A199;
  assign \new_[85501]_  = A202 & A201;
  assign \new_[85502]_  = \new_[85501]_  & \new_[85498]_ ;
  assign \new_[85503]_  = \new_[85502]_  & \new_[85495]_ ;
  assign \new_[85507]_  = A265 & A233;
  assign \new_[85508]_  = A232 & \new_[85507]_ ;
  assign \new_[85511]_  = ~A299 & A266;
  assign \new_[85514]_  = ~A302 & ~A301;
  assign \new_[85515]_  = \new_[85514]_  & \new_[85511]_ ;
  assign \new_[85516]_  = \new_[85515]_  & \new_[85508]_ ;
  assign \new_[85520]_  = ~A168 & ~A169;
  assign \new_[85521]_  = ~A170 & \new_[85520]_ ;
  assign \new_[85524]_  = ~A200 & A199;
  assign \new_[85527]_  = A202 & A201;
  assign \new_[85528]_  = \new_[85527]_  & \new_[85524]_ ;
  assign \new_[85529]_  = \new_[85528]_  & \new_[85521]_ ;
  assign \new_[85533]_  = ~A265 & A233;
  assign \new_[85534]_  = A232 & \new_[85533]_ ;
  assign \new_[85537]_  = ~A299 & ~A266;
  assign \new_[85540]_  = ~A302 & ~A301;
  assign \new_[85541]_  = \new_[85540]_  & \new_[85537]_ ;
  assign \new_[85542]_  = \new_[85541]_  & \new_[85534]_ ;
  assign \new_[85546]_  = ~A168 & ~A169;
  assign \new_[85547]_  = ~A170 & \new_[85546]_ ;
  assign \new_[85550]_  = ~A200 & A199;
  assign \new_[85553]_  = A202 & A201;
  assign \new_[85554]_  = \new_[85553]_  & \new_[85550]_ ;
  assign \new_[85555]_  = \new_[85554]_  & \new_[85547]_ ;
  assign \new_[85559]_  = ~A236 & ~A235;
  assign \new_[85560]_  = ~A233 & \new_[85559]_ ;
  assign \new_[85563]_  = A266 & A265;
  assign \new_[85566]_  = ~A300 & A298;
  assign \new_[85567]_  = \new_[85566]_  & \new_[85563]_ ;
  assign \new_[85568]_  = \new_[85567]_  & \new_[85560]_ ;
  assign \new_[85572]_  = ~A168 & ~A169;
  assign \new_[85573]_  = ~A170 & \new_[85572]_ ;
  assign \new_[85576]_  = ~A200 & A199;
  assign \new_[85579]_  = A202 & A201;
  assign \new_[85580]_  = \new_[85579]_  & \new_[85576]_ ;
  assign \new_[85581]_  = \new_[85580]_  & \new_[85573]_ ;
  assign \new_[85585]_  = ~A236 & ~A235;
  assign \new_[85586]_  = ~A233 & \new_[85585]_ ;
  assign \new_[85589]_  = A266 & A265;
  assign \new_[85592]_  = A299 & A298;
  assign \new_[85593]_  = \new_[85592]_  & \new_[85589]_ ;
  assign \new_[85594]_  = \new_[85593]_  & \new_[85586]_ ;
  assign \new_[85598]_  = ~A168 & ~A169;
  assign \new_[85599]_  = ~A170 & \new_[85598]_ ;
  assign \new_[85602]_  = ~A200 & A199;
  assign \new_[85605]_  = A202 & A201;
  assign \new_[85606]_  = \new_[85605]_  & \new_[85602]_ ;
  assign \new_[85607]_  = \new_[85606]_  & \new_[85599]_ ;
  assign \new_[85611]_  = ~A236 & ~A235;
  assign \new_[85612]_  = ~A233 & \new_[85611]_ ;
  assign \new_[85615]_  = A266 & A265;
  assign \new_[85618]_  = ~A299 & ~A298;
  assign \new_[85619]_  = \new_[85618]_  & \new_[85615]_ ;
  assign \new_[85620]_  = \new_[85619]_  & \new_[85612]_ ;
  assign \new_[85624]_  = ~A168 & ~A169;
  assign \new_[85625]_  = ~A170 & \new_[85624]_ ;
  assign \new_[85628]_  = ~A200 & A199;
  assign \new_[85631]_  = A202 & A201;
  assign \new_[85632]_  = \new_[85631]_  & \new_[85628]_ ;
  assign \new_[85633]_  = \new_[85632]_  & \new_[85625]_ ;
  assign \new_[85637]_  = ~A236 & ~A235;
  assign \new_[85638]_  = ~A233 & \new_[85637]_ ;
  assign \new_[85641]_  = ~A267 & ~A266;
  assign \new_[85644]_  = ~A300 & A298;
  assign \new_[85645]_  = \new_[85644]_  & \new_[85641]_ ;
  assign \new_[85646]_  = \new_[85645]_  & \new_[85638]_ ;
  assign \new_[85650]_  = ~A168 & ~A169;
  assign \new_[85651]_  = ~A170 & \new_[85650]_ ;
  assign \new_[85654]_  = ~A200 & A199;
  assign \new_[85657]_  = A202 & A201;
  assign \new_[85658]_  = \new_[85657]_  & \new_[85654]_ ;
  assign \new_[85659]_  = \new_[85658]_  & \new_[85651]_ ;
  assign \new_[85663]_  = ~A236 & ~A235;
  assign \new_[85664]_  = ~A233 & \new_[85663]_ ;
  assign \new_[85667]_  = ~A267 & ~A266;
  assign \new_[85670]_  = A299 & A298;
  assign \new_[85671]_  = \new_[85670]_  & \new_[85667]_ ;
  assign \new_[85672]_  = \new_[85671]_  & \new_[85664]_ ;
  assign \new_[85676]_  = ~A168 & ~A169;
  assign \new_[85677]_  = ~A170 & \new_[85676]_ ;
  assign \new_[85680]_  = ~A200 & A199;
  assign \new_[85683]_  = A202 & A201;
  assign \new_[85684]_  = \new_[85683]_  & \new_[85680]_ ;
  assign \new_[85685]_  = \new_[85684]_  & \new_[85677]_ ;
  assign \new_[85689]_  = ~A236 & ~A235;
  assign \new_[85690]_  = ~A233 & \new_[85689]_ ;
  assign \new_[85693]_  = ~A267 & ~A266;
  assign \new_[85696]_  = ~A299 & ~A298;
  assign \new_[85697]_  = \new_[85696]_  & \new_[85693]_ ;
  assign \new_[85698]_  = \new_[85697]_  & \new_[85690]_ ;
  assign \new_[85702]_  = ~A168 & ~A169;
  assign \new_[85703]_  = ~A170 & \new_[85702]_ ;
  assign \new_[85706]_  = ~A200 & A199;
  assign \new_[85709]_  = A202 & A201;
  assign \new_[85710]_  = \new_[85709]_  & \new_[85706]_ ;
  assign \new_[85711]_  = \new_[85710]_  & \new_[85703]_ ;
  assign \new_[85715]_  = ~A236 & ~A235;
  assign \new_[85716]_  = ~A233 & \new_[85715]_ ;
  assign \new_[85719]_  = ~A266 & ~A265;
  assign \new_[85722]_  = ~A300 & A298;
  assign \new_[85723]_  = \new_[85722]_  & \new_[85719]_ ;
  assign \new_[85724]_  = \new_[85723]_  & \new_[85716]_ ;
  assign \new_[85728]_  = ~A168 & ~A169;
  assign \new_[85729]_  = ~A170 & \new_[85728]_ ;
  assign \new_[85732]_  = ~A200 & A199;
  assign \new_[85735]_  = A202 & A201;
  assign \new_[85736]_  = \new_[85735]_  & \new_[85732]_ ;
  assign \new_[85737]_  = \new_[85736]_  & \new_[85729]_ ;
  assign \new_[85741]_  = ~A236 & ~A235;
  assign \new_[85742]_  = ~A233 & \new_[85741]_ ;
  assign \new_[85745]_  = ~A266 & ~A265;
  assign \new_[85748]_  = A299 & A298;
  assign \new_[85749]_  = \new_[85748]_  & \new_[85745]_ ;
  assign \new_[85750]_  = \new_[85749]_  & \new_[85742]_ ;
  assign \new_[85754]_  = ~A168 & ~A169;
  assign \new_[85755]_  = ~A170 & \new_[85754]_ ;
  assign \new_[85758]_  = ~A200 & A199;
  assign \new_[85761]_  = A202 & A201;
  assign \new_[85762]_  = \new_[85761]_  & \new_[85758]_ ;
  assign \new_[85763]_  = \new_[85762]_  & \new_[85755]_ ;
  assign \new_[85767]_  = ~A236 & ~A235;
  assign \new_[85768]_  = ~A233 & \new_[85767]_ ;
  assign \new_[85771]_  = ~A266 & ~A265;
  assign \new_[85774]_  = ~A299 & ~A298;
  assign \new_[85775]_  = \new_[85774]_  & \new_[85771]_ ;
  assign \new_[85776]_  = \new_[85775]_  & \new_[85768]_ ;
  assign \new_[85780]_  = ~A168 & ~A169;
  assign \new_[85781]_  = ~A170 & \new_[85780]_ ;
  assign \new_[85784]_  = ~A200 & A199;
  assign \new_[85787]_  = A202 & A201;
  assign \new_[85788]_  = \new_[85787]_  & \new_[85784]_ ;
  assign \new_[85789]_  = \new_[85788]_  & \new_[85781]_ ;
  assign \new_[85793]_  = A265 & ~A234;
  assign \new_[85794]_  = ~A233 & \new_[85793]_ ;
  assign \new_[85797]_  = A298 & A266;
  assign \new_[85800]_  = ~A302 & ~A301;
  assign \new_[85801]_  = \new_[85800]_  & \new_[85797]_ ;
  assign \new_[85802]_  = \new_[85801]_  & \new_[85794]_ ;
  assign \new_[85806]_  = ~A168 & ~A169;
  assign \new_[85807]_  = ~A170 & \new_[85806]_ ;
  assign \new_[85810]_  = ~A200 & A199;
  assign \new_[85813]_  = A202 & A201;
  assign \new_[85814]_  = \new_[85813]_  & \new_[85810]_ ;
  assign \new_[85815]_  = \new_[85814]_  & \new_[85807]_ ;
  assign \new_[85819]_  = ~A266 & ~A234;
  assign \new_[85820]_  = ~A233 & \new_[85819]_ ;
  assign \new_[85823]_  = ~A269 & ~A268;
  assign \new_[85826]_  = ~A300 & A298;
  assign \new_[85827]_  = \new_[85826]_  & \new_[85823]_ ;
  assign \new_[85828]_  = \new_[85827]_  & \new_[85820]_ ;
  assign \new_[85832]_  = ~A168 & ~A169;
  assign \new_[85833]_  = ~A170 & \new_[85832]_ ;
  assign \new_[85836]_  = ~A200 & A199;
  assign \new_[85839]_  = A202 & A201;
  assign \new_[85840]_  = \new_[85839]_  & \new_[85836]_ ;
  assign \new_[85841]_  = \new_[85840]_  & \new_[85833]_ ;
  assign \new_[85845]_  = ~A266 & ~A234;
  assign \new_[85846]_  = ~A233 & \new_[85845]_ ;
  assign \new_[85849]_  = ~A269 & ~A268;
  assign \new_[85852]_  = A299 & A298;
  assign \new_[85853]_  = \new_[85852]_  & \new_[85849]_ ;
  assign \new_[85854]_  = \new_[85853]_  & \new_[85846]_ ;
  assign \new_[85858]_  = ~A168 & ~A169;
  assign \new_[85859]_  = ~A170 & \new_[85858]_ ;
  assign \new_[85862]_  = ~A200 & A199;
  assign \new_[85865]_  = A202 & A201;
  assign \new_[85866]_  = \new_[85865]_  & \new_[85862]_ ;
  assign \new_[85867]_  = \new_[85866]_  & \new_[85859]_ ;
  assign \new_[85871]_  = ~A266 & ~A234;
  assign \new_[85872]_  = ~A233 & \new_[85871]_ ;
  assign \new_[85875]_  = ~A269 & ~A268;
  assign \new_[85878]_  = ~A299 & ~A298;
  assign \new_[85879]_  = \new_[85878]_  & \new_[85875]_ ;
  assign \new_[85880]_  = \new_[85879]_  & \new_[85872]_ ;
  assign \new_[85884]_  = ~A168 & ~A169;
  assign \new_[85885]_  = ~A170 & \new_[85884]_ ;
  assign \new_[85888]_  = ~A200 & A199;
  assign \new_[85891]_  = A202 & A201;
  assign \new_[85892]_  = \new_[85891]_  & \new_[85888]_ ;
  assign \new_[85893]_  = \new_[85892]_  & \new_[85885]_ ;
  assign \new_[85897]_  = ~A266 & ~A234;
  assign \new_[85898]_  = ~A233 & \new_[85897]_ ;
  assign \new_[85901]_  = A298 & ~A267;
  assign \new_[85904]_  = ~A302 & ~A301;
  assign \new_[85905]_  = \new_[85904]_  & \new_[85901]_ ;
  assign \new_[85906]_  = \new_[85905]_  & \new_[85898]_ ;
  assign \new_[85910]_  = ~A168 & ~A169;
  assign \new_[85911]_  = ~A170 & \new_[85910]_ ;
  assign \new_[85914]_  = ~A200 & A199;
  assign \new_[85917]_  = A202 & A201;
  assign \new_[85918]_  = \new_[85917]_  & \new_[85914]_ ;
  assign \new_[85919]_  = \new_[85918]_  & \new_[85911]_ ;
  assign \new_[85923]_  = ~A265 & ~A234;
  assign \new_[85924]_  = ~A233 & \new_[85923]_ ;
  assign \new_[85927]_  = A298 & ~A266;
  assign \new_[85930]_  = ~A302 & ~A301;
  assign \new_[85931]_  = \new_[85930]_  & \new_[85927]_ ;
  assign \new_[85932]_  = \new_[85931]_  & \new_[85924]_ ;
  assign \new_[85936]_  = ~A168 & ~A169;
  assign \new_[85937]_  = ~A170 & \new_[85936]_ ;
  assign \new_[85940]_  = ~A200 & A199;
  assign \new_[85943]_  = A202 & A201;
  assign \new_[85944]_  = \new_[85943]_  & \new_[85940]_ ;
  assign \new_[85945]_  = \new_[85944]_  & \new_[85937]_ ;
  assign \new_[85949]_  = A265 & ~A233;
  assign \new_[85950]_  = ~A232 & \new_[85949]_ ;
  assign \new_[85953]_  = A298 & A266;
  assign \new_[85956]_  = ~A302 & ~A301;
  assign \new_[85957]_  = \new_[85956]_  & \new_[85953]_ ;
  assign \new_[85958]_  = \new_[85957]_  & \new_[85950]_ ;
  assign \new_[85962]_  = ~A168 & ~A169;
  assign \new_[85963]_  = ~A170 & \new_[85962]_ ;
  assign \new_[85966]_  = ~A200 & A199;
  assign \new_[85969]_  = A202 & A201;
  assign \new_[85970]_  = \new_[85969]_  & \new_[85966]_ ;
  assign \new_[85971]_  = \new_[85970]_  & \new_[85963]_ ;
  assign \new_[85975]_  = ~A266 & ~A233;
  assign \new_[85976]_  = ~A232 & \new_[85975]_ ;
  assign \new_[85979]_  = ~A269 & ~A268;
  assign \new_[85982]_  = ~A300 & A298;
  assign \new_[85983]_  = \new_[85982]_  & \new_[85979]_ ;
  assign \new_[85984]_  = \new_[85983]_  & \new_[85976]_ ;
  assign \new_[85988]_  = ~A168 & ~A169;
  assign \new_[85989]_  = ~A170 & \new_[85988]_ ;
  assign \new_[85992]_  = ~A200 & A199;
  assign \new_[85995]_  = A202 & A201;
  assign \new_[85996]_  = \new_[85995]_  & \new_[85992]_ ;
  assign \new_[85997]_  = \new_[85996]_  & \new_[85989]_ ;
  assign \new_[86001]_  = ~A266 & ~A233;
  assign \new_[86002]_  = ~A232 & \new_[86001]_ ;
  assign \new_[86005]_  = ~A269 & ~A268;
  assign \new_[86008]_  = A299 & A298;
  assign \new_[86009]_  = \new_[86008]_  & \new_[86005]_ ;
  assign \new_[86010]_  = \new_[86009]_  & \new_[86002]_ ;
  assign \new_[86014]_  = ~A168 & ~A169;
  assign \new_[86015]_  = ~A170 & \new_[86014]_ ;
  assign \new_[86018]_  = ~A200 & A199;
  assign \new_[86021]_  = A202 & A201;
  assign \new_[86022]_  = \new_[86021]_  & \new_[86018]_ ;
  assign \new_[86023]_  = \new_[86022]_  & \new_[86015]_ ;
  assign \new_[86027]_  = ~A266 & ~A233;
  assign \new_[86028]_  = ~A232 & \new_[86027]_ ;
  assign \new_[86031]_  = ~A269 & ~A268;
  assign \new_[86034]_  = ~A299 & ~A298;
  assign \new_[86035]_  = \new_[86034]_  & \new_[86031]_ ;
  assign \new_[86036]_  = \new_[86035]_  & \new_[86028]_ ;
  assign \new_[86040]_  = ~A168 & ~A169;
  assign \new_[86041]_  = ~A170 & \new_[86040]_ ;
  assign \new_[86044]_  = ~A200 & A199;
  assign \new_[86047]_  = A202 & A201;
  assign \new_[86048]_  = \new_[86047]_  & \new_[86044]_ ;
  assign \new_[86049]_  = \new_[86048]_  & \new_[86041]_ ;
  assign \new_[86053]_  = ~A266 & ~A233;
  assign \new_[86054]_  = ~A232 & \new_[86053]_ ;
  assign \new_[86057]_  = A298 & ~A267;
  assign \new_[86060]_  = ~A302 & ~A301;
  assign \new_[86061]_  = \new_[86060]_  & \new_[86057]_ ;
  assign \new_[86062]_  = \new_[86061]_  & \new_[86054]_ ;
  assign \new_[86066]_  = ~A168 & ~A169;
  assign \new_[86067]_  = ~A170 & \new_[86066]_ ;
  assign \new_[86070]_  = ~A200 & A199;
  assign \new_[86073]_  = A202 & A201;
  assign \new_[86074]_  = \new_[86073]_  & \new_[86070]_ ;
  assign \new_[86075]_  = \new_[86074]_  & \new_[86067]_ ;
  assign \new_[86079]_  = ~A265 & ~A233;
  assign \new_[86080]_  = ~A232 & \new_[86079]_ ;
  assign \new_[86083]_  = A298 & ~A266;
  assign \new_[86086]_  = ~A302 & ~A301;
  assign \new_[86087]_  = \new_[86086]_  & \new_[86083]_ ;
  assign \new_[86088]_  = \new_[86087]_  & \new_[86080]_ ;
  assign \new_[86092]_  = ~A168 & ~A169;
  assign \new_[86093]_  = ~A170 & \new_[86092]_ ;
  assign \new_[86096]_  = ~A200 & A199;
  assign \new_[86099]_  = A203 & A201;
  assign \new_[86100]_  = \new_[86099]_  & \new_[86096]_ ;
  assign \new_[86101]_  = \new_[86100]_  & \new_[86093]_ ;
  assign \new_[86105]_  = A265 & A233;
  assign \new_[86106]_  = A232 & \new_[86105]_ ;
  assign \new_[86109]_  = ~A269 & ~A268;
  assign \new_[86112]_  = ~A300 & ~A299;
  assign \new_[86113]_  = \new_[86112]_  & \new_[86109]_ ;
  assign \new_[86114]_  = \new_[86113]_  & \new_[86106]_ ;
  assign \new_[86118]_  = ~A168 & ~A169;
  assign \new_[86119]_  = ~A170 & \new_[86118]_ ;
  assign \new_[86122]_  = ~A200 & A199;
  assign \new_[86125]_  = A203 & A201;
  assign \new_[86126]_  = \new_[86125]_  & \new_[86122]_ ;
  assign \new_[86127]_  = \new_[86126]_  & \new_[86119]_ ;
  assign \new_[86131]_  = A265 & A233;
  assign \new_[86132]_  = A232 & \new_[86131]_ ;
  assign \new_[86135]_  = ~A269 & ~A268;
  assign \new_[86138]_  = A299 & A298;
  assign \new_[86139]_  = \new_[86138]_  & \new_[86135]_ ;
  assign \new_[86140]_  = \new_[86139]_  & \new_[86132]_ ;
  assign \new_[86144]_  = ~A168 & ~A169;
  assign \new_[86145]_  = ~A170 & \new_[86144]_ ;
  assign \new_[86148]_  = ~A200 & A199;
  assign \new_[86151]_  = A203 & A201;
  assign \new_[86152]_  = \new_[86151]_  & \new_[86148]_ ;
  assign \new_[86153]_  = \new_[86152]_  & \new_[86145]_ ;
  assign \new_[86157]_  = A265 & A233;
  assign \new_[86158]_  = A232 & \new_[86157]_ ;
  assign \new_[86161]_  = ~A269 & ~A268;
  assign \new_[86164]_  = ~A299 & ~A298;
  assign \new_[86165]_  = \new_[86164]_  & \new_[86161]_ ;
  assign \new_[86166]_  = \new_[86165]_  & \new_[86158]_ ;
  assign \new_[86170]_  = ~A168 & ~A169;
  assign \new_[86171]_  = ~A170 & \new_[86170]_ ;
  assign \new_[86174]_  = ~A200 & A199;
  assign \new_[86177]_  = A203 & A201;
  assign \new_[86178]_  = \new_[86177]_  & \new_[86174]_ ;
  assign \new_[86179]_  = \new_[86178]_  & \new_[86171]_ ;
  assign \new_[86183]_  = A265 & A233;
  assign \new_[86184]_  = A232 & \new_[86183]_ ;
  assign \new_[86187]_  = ~A299 & ~A267;
  assign \new_[86190]_  = ~A302 & ~A301;
  assign \new_[86191]_  = \new_[86190]_  & \new_[86187]_ ;
  assign \new_[86192]_  = \new_[86191]_  & \new_[86184]_ ;
  assign \new_[86196]_  = ~A168 & ~A169;
  assign \new_[86197]_  = ~A170 & \new_[86196]_ ;
  assign \new_[86200]_  = ~A200 & A199;
  assign \new_[86203]_  = A203 & A201;
  assign \new_[86204]_  = \new_[86203]_  & \new_[86200]_ ;
  assign \new_[86205]_  = \new_[86204]_  & \new_[86197]_ ;
  assign \new_[86209]_  = A265 & A233;
  assign \new_[86210]_  = A232 & \new_[86209]_ ;
  assign \new_[86213]_  = ~A299 & A266;
  assign \new_[86216]_  = ~A302 & ~A301;
  assign \new_[86217]_  = \new_[86216]_  & \new_[86213]_ ;
  assign \new_[86218]_  = \new_[86217]_  & \new_[86210]_ ;
  assign \new_[86222]_  = ~A168 & ~A169;
  assign \new_[86223]_  = ~A170 & \new_[86222]_ ;
  assign \new_[86226]_  = ~A200 & A199;
  assign \new_[86229]_  = A203 & A201;
  assign \new_[86230]_  = \new_[86229]_  & \new_[86226]_ ;
  assign \new_[86231]_  = \new_[86230]_  & \new_[86223]_ ;
  assign \new_[86235]_  = ~A265 & A233;
  assign \new_[86236]_  = A232 & \new_[86235]_ ;
  assign \new_[86239]_  = ~A299 & ~A266;
  assign \new_[86242]_  = ~A302 & ~A301;
  assign \new_[86243]_  = \new_[86242]_  & \new_[86239]_ ;
  assign \new_[86244]_  = \new_[86243]_  & \new_[86236]_ ;
  assign \new_[86248]_  = ~A168 & ~A169;
  assign \new_[86249]_  = ~A170 & \new_[86248]_ ;
  assign \new_[86252]_  = ~A200 & A199;
  assign \new_[86255]_  = A203 & A201;
  assign \new_[86256]_  = \new_[86255]_  & \new_[86252]_ ;
  assign \new_[86257]_  = \new_[86256]_  & \new_[86249]_ ;
  assign \new_[86261]_  = ~A236 & ~A235;
  assign \new_[86262]_  = ~A233 & \new_[86261]_ ;
  assign \new_[86265]_  = A266 & A265;
  assign \new_[86268]_  = ~A300 & A298;
  assign \new_[86269]_  = \new_[86268]_  & \new_[86265]_ ;
  assign \new_[86270]_  = \new_[86269]_  & \new_[86262]_ ;
  assign \new_[86274]_  = ~A168 & ~A169;
  assign \new_[86275]_  = ~A170 & \new_[86274]_ ;
  assign \new_[86278]_  = ~A200 & A199;
  assign \new_[86281]_  = A203 & A201;
  assign \new_[86282]_  = \new_[86281]_  & \new_[86278]_ ;
  assign \new_[86283]_  = \new_[86282]_  & \new_[86275]_ ;
  assign \new_[86287]_  = ~A236 & ~A235;
  assign \new_[86288]_  = ~A233 & \new_[86287]_ ;
  assign \new_[86291]_  = A266 & A265;
  assign \new_[86294]_  = A299 & A298;
  assign \new_[86295]_  = \new_[86294]_  & \new_[86291]_ ;
  assign \new_[86296]_  = \new_[86295]_  & \new_[86288]_ ;
  assign \new_[86300]_  = ~A168 & ~A169;
  assign \new_[86301]_  = ~A170 & \new_[86300]_ ;
  assign \new_[86304]_  = ~A200 & A199;
  assign \new_[86307]_  = A203 & A201;
  assign \new_[86308]_  = \new_[86307]_  & \new_[86304]_ ;
  assign \new_[86309]_  = \new_[86308]_  & \new_[86301]_ ;
  assign \new_[86313]_  = ~A236 & ~A235;
  assign \new_[86314]_  = ~A233 & \new_[86313]_ ;
  assign \new_[86317]_  = A266 & A265;
  assign \new_[86320]_  = ~A299 & ~A298;
  assign \new_[86321]_  = \new_[86320]_  & \new_[86317]_ ;
  assign \new_[86322]_  = \new_[86321]_  & \new_[86314]_ ;
  assign \new_[86326]_  = ~A168 & ~A169;
  assign \new_[86327]_  = ~A170 & \new_[86326]_ ;
  assign \new_[86330]_  = ~A200 & A199;
  assign \new_[86333]_  = A203 & A201;
  assign \new_[86334]_  = \new_[86333]_  & \new_[86330]_ ;
  assign \new_[86335]_  = \new_[86334]_  & \new_[86327]_ ;
  assign \new_[86339]_  = ~A236 & ~A235;
  assign \new_[86340]_  = ~A233 & \new_[86339]_ ;
  assign \new_[86343]_  = ~A267 & ~A266;
  assign \new_[86346]_  = ~A300 & A298;
  assign \new_[86347]_  = \new_[86346]_  & \new_[86343]_ ;
  assign \new_[86348]_  = \new_[86347]_  & \new_[86340]_ ;
  assign \new_[86352]_  = ~A168 & ~A169;
  assign \new_[86353]_  = ~A170 & \new_[86352]_ ;
  assign \new_[86356]_  = ~A200 & A199;
  assign \new_[86359]_  = A203 & A201;
  assign \new_[86360]_  = \new_[86359]_  & \new_[86356]_ ;
  assign \new_[86361]_  = \new_[86360]_  & \new_[86353]_ ;
  assign \new_[86365]_  = ~A236 & ~A235;
  assign \new_[86366]_  = ~A233 & \new_[86365]_ ;
  assign \new_[86369]_  = ~A267 & ~A266;
  assign \new_[86372]_  = A299 & A298;
  assign \new_[86373]_  = \new_[86372]_  & \new_[86369]_ ;
  assign \new_[86374]_  = \new_[86373]_  & \new_[86366]_ ;
  assign \new_[86378]_  = ~A168 & ~A169;
  assign \new_[86379]_  = ~A170 & \new_[86378]_ ;
  assign \new_[86382]_  = ~A200 & A199;
  assign \new_[86385]_  = A203 & A201;
  assign \new_[86386]_  = \new_[86385]_  & \new_[86382]_ ;
  assign \new_[86387]_  = \new_[86386]_  & \new_[86379]_ ;
  assign \new_[86391]_  = ~A236 & ~A235;
  assign \new_[86392]_  = ~A233 & \new_[86391]_ ;
  assign \new_[86395]_  = ~A267 & ~A266;
  assign \new_[86398]_  = ~A299 & ~A298;
  assign \new_[86399]_  = \new_[86398]_  & \new_[86395]_ ;
  assign \new_[86400]_  = \new_[86399]_  & \new_[86392]_ ;
  assign \new_[86404]_  = ~A168 & ~A169;
  assign \new_[86405]_  = ~A170 & \new_[86404]_ ;
  assign \new_[86408]_  = ~A200 & A199;
  assign \new_[86411]_  = A203 & A201;
  assign \new_[86412]_  = \new_[86411]_  & \new_[86408]_ ;
  assign \new_[86413]_  = \new_[86412]_  & \new_[86405]_ ;
  assign \new_[86417]_  = ~A236 & ~A235;
  assign \new_[86418]_  = ~A233 & \new_[86417]_ ;
  assign \new_[86421]_  = ~A266 & ~A265;
  assign \new_[86424]_  = ~A300 & A298;
  assign \new_[86425]_  = \new_[86424]_  & \new_[86421]_ ;
  assign \new_[86426]_  = \new_[86425]_  & \new_[86418]_ ;
  assign \new_[86430]_  = ~A168 & ~A169;
  assign \new_[86431]_  = ~A170 & \new_[86430]_ ;
  assign \new_[86434]_  = ~A200 & A199;
  assign \new_[86437]_  = A203 & A201;
  assign \new_[86438]_  = \new_[86437]_  & \new_[86434]_ ;
  assign \new_[86439]_  = \new_[86438]_  & \new_[86431]_ ;
  assign \new_[86443]_  = ~A236 & ~A235;
  assign \new_[86444]_  = ~A233 & \new_[86443]_ ;
  assign \new_[86447]_  = ~A266 & ~A265;
  assign \new_[86450]_  = A299 & A298;
  assign \new_[86451]_  = \new_[86450]_  & \new_[86447]_ ;
  assign \new_[86452]_  = \new_[86451]_  & \new_[86444]_ ;
  assign \new_[86456]_  = ~A168 & ~A169;
  assign \new_[86457]_  = ~A170 & \new_[86456]_ ;
  assign \new_[86460]_  = ~A200 & A199;
  assign \new_[86463]_  = A203 & A201;
  assign \new_[86464]_  = \new_[86463]_  & \new_[86460]_ ;
  assign \new_[86465]_  = \new_[86464]_  & \new_[86457]_ ;
  assign \new_[86469]_  = ~A236 & ~A235;
  assign \new_[86470]_  = ~A233 & \new_[86469]_ ;
  assign \new_[86473]_  = ~A266 & ~A265;
  assign \new_[86476]_  = ~A299 & ~A298;
  assign \new_[86477]_  = \new_[86476]_  & \new_[86473]_ ;
  assign \new_[86478]_  = \new_[86477]_  & \new_[86470]_ ;
  assign \new_[86482]_  = ~A168 & ~A169;
  assign \new_[86483]_  = ~A170 & \new_[86482]_ ;
  assign \new_[86486]_  = ~A200 & A199;
  assign \new_[86489]_  = A203 & A201;
  assign \new_[86490]_  = \new_[86489]_  & \new_[86486]_ ;
  assign \new_[86491]_  = \new_[86490]_  & \new_[86483]_ ;
  assign \new_[86495]_  = A265 & ~A234;
  assign \new_[86496]_  = ~A233 & \new_[86495]_ ;
  assign \new_[86499]_  = A298 & A266;
  assign \new_[86502]_  = ~A302 & ~A301;
  assign \new_[86503]_  = \new_[86502]_  & \new_[86499]_ ;
  assign \new_[86504]_  = \new_[86503]_  & \new_[86496]_ ;
  assign \new_[86508]_  = ~A168 & ~A169;
  assign \new_[86509]_  = ~A170 & \new_[86508]_ ;
  assign \new_[86512]_  = ~A200 & A199;
  assign \new_[86515]_  = A203 & A201;
  assign \new_[86516]_  = \new_[86515]_  & \new_[86512]_ ;
  assign \new_[86517]_  = \new_[86516]_  & \new_[86509]_ ;
  assign \new_[86521]_  = ~A266 & ~A234;
  assign \new_[86522]_  = ~A233 & \new_[86521]_ ;
  assign \new_[86525]_  = ~A269 & ~A268;
  assign \new_[86528]_  = ~A300 & A298;
  assign \new_[86529]_  = \new_[86528]_  & \new_[86525]_ ;
  assign \new_[86530]_  = \new_[86529]_  & \new_[86522]_ ;
  assign \new_[86534]_  = ~A168 & ~A169;
  assign \new_[86535]_  = ~A170 & \new_[86534]_ ;
  assign \new_[86538]_  = ~A200 & A199;
  assign \new_[86541]_  = A203 & A201;
  assign \new_[86542]_  = \new_[86541]_  & \new_[86538]_ ;
  assign \new_[86543]_  = \new_[86542]_  & \new_[86535]_ ;
  assign \new_[86547]_  = ~A266 & ~A234;
  assign \new_[86548]_  = ~A233 & \new_[86547]_ ;
  assign \new_[86551]_  = ~A269 & ~A268;
  assign \new_[86554]_  = A299 & A298;
  assign \new_[86555]_  = \new_[86554]_  & \new_[86551]_ ;
  assign \new_[86556]_  = \new_[86555]_  & \new_[86548]_ ;
  assign \new_[86560]_  = ~A168 & ~A169;
  assign \new_[86561]_  = ~A170 & \new_[86560]_ ;
  assign \new_[86564]_  = ~A200 & A199;
  assign \new_[86567]_  = A203 & A201;
  assign \new_[86568]_  = \new_[86567]_  & \new_[86564]_ ;
  assign \new_[86569]_  = \new_[86568]_  & \new_[86561]_ ;
  assign \new_[86573]_  = ~A266 & ~A234;
  assign \new_[86574]_  = ~A233 & \new_[86573]_ ;
  assign \new_[86577]_  = ~A269 & ~A268;
  assign \new_[86580]_  = ~A299 & ~A298;
  assign \new_[86581]_  = \new_[86580]_  & \new_[86577]_ ;
  assign \new_[86582]_  = \new_[86581]_  & \new_[86574]_ ;
  assign \new_[86586]_  = ~A168 & ~A169;
  assign \new_[86587]_  = ~A170 & \new_[86586]_ ;
  assign \new_[86590]_  = ~A200 & A199;
  assign \new_[86593]_  = A203 & A201;
  assign \new_[86594]_  = \new_[86593]_  & \new_[86590]_ ;
  assign \new_[86595]_  = \new_[86594]_  & \new_[86587]_ ;
  assign \new_[86599]_  = ~A266 & ~A234;
  assign \new_[86600]_  = ~A233 & \new_[86599]_ ;
  assign \new_[86603]_  = A298 & ~A267;
  assign \new_[86606]_  = ~A302 & ~A301;
  assign \new_[86607]_  = \new_[86606]_  & \new_[86603]_ ;
  assign \new_[86608]_  = \new_[86607]_  & \new_[86600]_ ;
  assign \new_[86612]_  = ~A168 & ~A169;
  assign \new_[86613]_  = ~A170 & \new_[86612]_ ;
  assign \new_[86616]_  = ~A200 & A199;
  assign \new_[86619]_  = A203 & A201;
  assign \new_[86620]_  = \new_[86619]_  & \new_[86616]_ ;
  assign \new_[86621]_  = \new_[86620]_  & \new_[86613]_ ;
  assign \new_[86625]_  = ~A265 & ~A234;
  assign \new_[86626]_  = ~A233 & \new_[86625]_ ;
  assign \new_[86629]_  = A298 & ~A266;
  assign \new_[86632]_  = ~A302 & ~A301;
  assign \new_[86633]_  = \new_[86632]_  & \new_[86629]_ ;
  assign \new_[86634]_  = \new_[86633]_  & \new_[86626]_ ;
  assign \new_[86638]_  = ~A168 & ~A169;
  assign \new_[86639]_  = ~A170 & \new_[86638]_ ;
  assign \new_[86642]_  = ~A200 & A199;
  assign \new_[86645]_  = A203 & A201;
  assign \new_[86646]_  = \new_[86645]_  & \new_[86642]_ ;
  assign \new_[86647]_  = \new_[86646]_  & \new_[86639]_ ;
  assign \new_[86651]_  = A265 & ~A233;
  assign \new_[86652]_  = ~A232 & \new_[86651]_ ;
  assign \new_[86655]_  = A298 & A266;
  assign \new_[86658]_  = ~A302 & ~A301;
  assign \new_[86659]_  = \new_[86658]_  & \new_[86655]_ ;
  assign \new_[86660]_  = \new_[86659]_  & \new_[86652]_ ;
  assign \new_[86664]_  = ~A168 & ~A169;
  assign \new_[86665]_  = ~A170 & \new_[86664]_ ;
  assign \new_[86668]_  = ~A200 & A199;
  assign \new_[86671]_  = A203 & A201;
  assign \new_[86672]_  = \new_[86671]_  & \new_[86668]_ ;
  assign \new_[86673]_  = \new_[86672]_  & \new_[86665]_ ;
  assign \new_[86677]_  = ~A266 & ~A233;
  assign \new_[86678]_  = ~A232 & \new_[86677]_ ;
  assign \new_[86681]_  = ~A269 & ~A268;
  assign \new_[86684]_  = ~A300 & A298;
  assign \new_[86685]_  = \new_[86684]_  & \new_[86681]_ ;
  assign \new_[86686]_  = \new_[86685]_  & \new_[86678]_ ;
  assign \new_[86690]_  = ~A168 & ~A169;
  assign \new_[86691]_  = ~A170 & \new_[86690]_ ;
  assign \new_[86694]_  = ~A200 & A199;
  assign \new_[86697]_  = A203 & A201;
  assign \new_[86698]_  = \new_[86697]_  & \new_[86694]_ ;
  assign \new_[86699]_  = \new_[86698]_  & \new_[86691]_ ;
  assign \new_[86703]_  = ~A266 & ~A233;
  assign \new_[86704]_  = ~A232 & \new_[86703]_ ;
  assign \new_[86707]_  = ~A269 & ~A268;
  assign \new_[86710]_  = A299 & A298;
  assign \new_[86711]_  = \new_[86710]_  & \new_[86707]_ ;
  assign \new_[86712]_  = \new_[86711]_  & \new_[86704]_ ;
  assign \new_[86716]_  = ~A168 & ~A169;
  assign \new_[86717]_  = ~A170 & \new_[86716]_ ;
  assign \new_[86720]_  = ~A200 & A199;
  assign \new_[86723]_  = A203 & A201;
  assign \new_[86724]_  = \new_[86723]_  & \new_[86720]_ ;
  assign \new_[86725]_  = \new_[86724]_  & \new_[86717]_ ;
  assign \new_[86729]_  = ~A266 & ~A233;
  assign \new_[86730]_  = ~A232 & \new_[86729]_ ;
  assign \new_[86733]_  = ~A269 & ~A268;
  assign \new_[86736]_  = ~A299 & ~A298;
  assign \new_[86737]_  = \new_[86736]_  & \new_[86733]_ ;
  assign \new_[86738]_  = \new_[86737]_  & \new_[86730]_ ;
  assign \new_[86742]_  = ~A168 & ~A169;
  assign \new_[86743]_  = ~A170 & \new_[86742]_ ;
  assign \new_[86746]_  = ~A200 & A199;
  assign \new_[86749]_  = A203 & A201;
  assign \new_[86750]_  = \new_[86749]_  & \new_[86746]_ ;
  assign \new_[86751]_  = \new_[86750]_  & \new_[86743]_ ;
  assign \new_[86755]_  = ~A266 & ~A233;
  assign \new_[86756]_  = ~A232 & \new_[86755]_ ;
  assign \new_[86759]_  = A298 & ~A267;
  assign \new_[86762]_  = ~A302 & ~A301;
  assign \new_[86763]_  = \new_[86762]_  & \new_[86759]_ ;
  assign \new_[86764]_  = \new_[86763]_  & \new_[86756]_ ;
  assign \new_[86768]_  = ~A168 & ~A169;
  assign \new_[86769]_  = ~A170 & \new_[86768]_ ;
  assign \new_[86772]_  = ~A200 & A199;
  assign \new_[86775]_  = A203 & A201;
  assign \new_[86776]_  = \new_[86775]_  & \new_[86772]_ ;
  assign \new_[86777]_  = \new_[86776]_  & \new_[86769]_ ;
  assign \new_[86781]_  = ~A265 & ~A233;
  assign \new_[86782]_  = ~A232 & \new_[86781]_ ;
  assign \new_[86785]_  = A298 & ~A266;
  assign \new_[86788]_  = ~A302 & ~A301;
  assign \new_[86789]_  = \new_[86788]_  & \new_[86785]_ ;
  assign \new_[86790]_  = \new_[86789]_  & \new_[86782]_ ;
  assign \new_[86794]_  = ~A166 & ~A167;
  assign \new_[86795]_  = A170 & \new_[86794]_ ;
  assign \new_[86798]_  = ~A200 & A199;
  assign \new_[86801]_  = A202 & A201;
  assign \new_[86802]_  = \new_[86801]_  & \new_[86798]_ ;
  assign \new_[86803]_  = \new_[86802]_  & \new_[86795]_ ;
  assign \new_[86806]_  = A233 & A232;
  assign \new_[86809]_  = ~A268 & A265;
  assign \new_[86810]_  = \new_[86809]_  & \new_[86806]_ ;
  assign \new_[86813]_  = ~A299 & ~A269;
  assign \new_[86816]_  = ~A302 & ~A301;
  assign \new_[86817]_  = \new_[86816]_  & \new_[86813]_ ;
  assign \new_[86818]_  = \new_[86817]_  & \new_[86810]_ ;
  assign \new_[86822]_  = ~A166 & ~A167;
  assign \new_[86823]_  = A170 & \new_[86822]_ ;
  assign \new_[86826]_  = ~A200 & A199;
  assign \new_[86829]_  = A202 & A201;
  assign \new_[86830]_  = \new_[86829]_  & \new_[86826]_ ;
  assign \new_[86831]_  = \new_[86830]_  & \new_[86823]_ ;
  assign \new_[86834]_  = ~A235 & ~A233;
  assign \new_[86837]_  = A265 & ~A236;
  assign \new_[86838]_  = \new_[86837]_  & \new_[86834]_ ;
  assign \new_[86841]_  = A298 & A266;
  assign \new_[86844]_  = ~A302 & ~A301;
  assign \new_[86845]_  = \new_[86844]_  & \new_[86841]_ ;
  assign \new_[86846]_  = \new_[86845]_  & \new_[86838]_ ;
  assign \new_[86850]_  = ~A166 & ~A167;
  assign \new_[86851]_  = A170 & \new_[86850]_ ;
  assign \new_[86854]_  = ~A200 & A199;
  assign \new_[86857]_  = A202 & A201;
  assign \new_[86858]_  = \new_[86857]_  & \new_[86854]_ ;
  assign \new_[86859]_  = \new_[86858]_  & \new_[86851]_ ;
  assign \new_[86862]_  = ~A235 & ~A233;
  assign \new_[86865]_  = ~A266 & ~A236;
  assign \new_[86866]_  = \new_[86865]_  & \new_[86862]_ ;
  assign \new_[86869]_  = ~A269 & ~A268;
  assign \new_[86872]_  = ~A300 & A298;
  assign \new_[86873]_  = \new_[86872]_  & \new_[86869]_ ;
  assign \new_[86874]_  = \new_[86873]_  & \new_[86866]_ ;
  assign \new_[86878]_  = ~A166 & ~A167;
  assign \new_[86879]_  = A170 & \new_[86878]_ ;
  assign \new_[86882]_  = ~A200 & A199;
  assign \new_[86885]_  = A202 & A201;
  assign \new_[86886]_  = \new_[86885]_  & \new_[86882]_ ;
  assign \new_[86887]_  = \new_[86886]_  & \new_[86879]_ ;
  assign \new_[86890]_  = ~A235 & ~A233;
  assign \new_[86893]_  = ~A266 & ~A236;
  assign \new_[86894]_  = \new_[86893]_  & \new_[86890]_ ;
  assign \new_[86897]_  = ~A269 & ~A268;
  assign \new_[86900]_  = A299 & A298;
  assign \new_[86901]_  = \new_[86900]_  & \new_[86897]_ ;
  assign \new_[86902]_  = \new_[86901]_  & \new_[86894]_ ;
  assign \new_[86906]_  = ~A166 & ~A167;
  assign \new_[86907]_  = A170 & \new_[86906]_ ;
  assign \new_[86910]_  = ~A200 & A199;
  assign \new_[86913]_  = A202 & A201;
  assign \new_[86914]_  = \new_[86913]_  & \new_[86910]_ ;
  assign \new_[86915]_  = \new_[86914]_  & \new_[86907]_ ;
  assign \new_[86918]_  = ~A235 & ~A233;
  assign \new_[86921]_  = ~A266 & ~A236;
  assign \new_[86922]_  = \new_[86921]_  & \new_[86918]_ ;
  assign \new_[86925]_  = ~A269 & ~A268;
  assign \new_[86928]_  = ~A299 & ~A298;
  assign \new_[86929]_  = \new_[86928]_  & \new_[86925]_ ;
  assign \new_[86930]_  = \new_[86929]_  & \new_[86922]_ ;
  assign \new_[86934]_  = ~A166 & ~A167;
  assign \new_[86935]_  = A170 & \new_[86934]_ ;
  assign \new_[86938]_  = ~A200 & A199;
  assign \new_[86941]_  = A202 & A201;
  assign \new_[86942]_  = \new_[86941]_  & \new_[86938]_ ;
  assign \new_[86943]_  = \new_[86942]_  & \new_[86935]_ ;
  assign \new_[86946]_  = ~A235 & ~A233;
  assign \new_[86949]_  = ~A266 & ~A236;
  assign \new_[86950]_  = \new_[86949]_  & \new_[86946]_ ;
  assign \new_[86953]_  = A298 & ~A267;
  assign \new_[86956]_  = ~A302 & ~A301;
  assign \new_[86957]_  = \new_[86956]_  & \new_[86953]_ ;
  assign \new_[86958]_  = \new_[86957]_  & \new_[86950]_ ;
  assign \new_[86962]_  = ~A166 & ~A167;
  assign \new_[86963]_  = A170 & \new_[86962]_ ;
  assign \new_[86966]_  = ~A200 & A199;
  assign \new_[86969]_  = A202 & A201;
  assign \new_[86970]_  = \new_[86969]_  & \new_[86966]_ ;
  assign \new_[86971]_  = \new_[86970]_  & \new_[86963]_ ;
  assign \new_[86974]_  = ~A235 & ~A233;
  assign \new_[86977]_  = ~A265 & ~A236;
  assign \new_[86978]_  = \new_[86977]_  & \new_[86974]_ ;
  assign \new_[86981]_  = A298 & ~A266;
  assign \new_[86984]_  = ~A302 & ~A301;
  assign \new_[86985]_  = \new_[86984]_  & \new_[86981]_ ;
  assign \new_[86986]_  = \new_[86985]_  & \new_[86978]_ ;
  assign \new_[86990]_  = ~A166 & ~A167;
  assign \new_[86991]_  = A170 & \new_[86990]_ ;
  assign \new_[86994]_  = ~A200 & A199;
  assign \new_[86997]_  = A202 & A201;
  assign \new_[86998]_  = \new_[86997]_  & \new_[86994]_ ;
  assign \new_[86999]_  = \new_[86998]_  & \new_[86991]_ ;
  assign \new_[87002]_  = ~A234 & ~A233;
  assign \new_[87005]_  = ~A268 & ~A266;
  assign \new_[87006]_  = \new_[87005]_  & \new_[87002]_ ;
  assign \new_[87009]_  = A298 & ~A269;
  assign \new_[87012]_  = ~A302 & ~A301;
  assign \new_[87013]_  = \new_[87012]_  & \new_[87009]_ ;
  assign \new_[87014]_  = \new_[87013]_  & \new_[87006]_ ;
  assign \new_[87018]_  = ~A166 & ~A167;
  assign \new_[87019]_  = A170 & \new_[87018]_ ;
  assign \new_[87022]_  = ~A200 & A199;
  assign \new_[87025]_  = A202 & A201;
  assign \new_[87026]_  = \new_[87025]_  & \new_[87022]_ ;
  assign \new_[87027]_  = \new_[87026]_  & \new_[87019]_ ;
  assign \new_[87030]_  = ~A233 & A232;
  assign \new_[87033]_  = A235 & A234;
  assign \new_[87034]_  = \new_[87033]_  & \new_[87030]_ ;
  assign \new_[87037]_  = ~A299 & A298;
  assign \new_[87040]_  = A301 & A300;
  assign \new_[87041]_  = \new_[87040]_  & \new_[87037]_ ;
  assign \new_[87042]_  = \new_[87041]_  & \new_[87034]_ ;
  assign \new_[87046]_  = ~A166 & ~A167;
  assign \new_[87047]_  = A170 & \new_[87046]_ ;
  assign \new_[87050]_  = ~A200 & A199;
  assign \new_[87053]_  = A202 & A201;
  assign \new_[87054]_  = \new_[87053]_  & \new_[87050]_ ;
  assign \new_[87055]_  = \new_[87054]_  & \new_[87047]_ ;
  assign \new_[87058]_  = ~A233 & A232;
  assign \new_[87061]_  = A235 & A234;
  assign \new_[87062]_  = \new_[87061]_  & \new_[87058]_ ;
  assign \new_[87065]_  = ~A299 & A298;
  assign \new_[87068]_  = A302 & A300;
  assign \new_[87069]_  = \new_[87068]_  & \new_[87065]_ ;
  assign \new_[87070]_  = \new_[87069]_  & \new_[87062]_ ;
  assign \new_[87074]_  = ~A166 & ~A167;
  assign \new_[87075]_  = A170 & \new_[87074]_ ;
  assign \new_[87078]_  = ~A200 & A199;
  assign \new_[87081]_  = A202 & A201;
  assign \new_[87082]_  = \new_[87081]_  & \new_[87078]_ ;
  assign \new_[87083]_  = \new_[87082]_  & \new_[87075]_ ;
  assign \new_[87086]_  = ~A233 & A232;
  assign \new_[87089]_  = A235 & A234;
  assign \new_[87090]_  = \new_[87089]_  & \new_[87086]_ ;
  assign \new_[87093]_  = ~A266 & A265;
  assign \new_[87096]_  = A268 & A267;
  assign \new_[87097]_  = \new_[87096]_  & \new_[87093]_ ;
  assign \new_[87098]_  = \new_[87097]_  & \new_[87090]_ ;
  assign \new_[87102]_  = ~A166 & ~A167;
  assign \new_[87103]_  = A170 & \new_[87102]_ ;
  assign \new_[87106]_  = ~A200 & A199;
  assign \new_[87109]_  = A202 & A201;
  assign \new_[87110]_  = \new_[87109]_  & \new_[87106]_ ;
  assign \new_[87111]_  = \new_[87110]_  & \new_[87103]_ ;
  assign \new_[87114]_  = ~A233 & A232;
  assign \new_[87117]_  = A235 & A234;
  assign \new_[87118]_  = \new_[87117]_  & \new_[87114]_ ;
  assign \new_[87121]_  = ~A266 & A265;
  assign \new_[87124]_  = A269 & A267;
  assign \new_[87125]_  = \new_[87124]_  & \new_[87121]_ ;
  assign \new_[87126]_  = \new_[87125]_  & \new_[87118]_ ;
  assign \new_[87130]_  = ~A166 & ~A167;
  assign \new_[87131]_  = A170 & \new_[87130]_ ;
  assign \new_[87134]_  = ~A200 & A199;
  assign \new_[87137]_  = A202 & A201;
  assign \new_[87138]_  = \new_[87137]_  & \new_[87134]_ ;
  assign \new_[87139]_  = \new_[87138]_  & \new_[87131]_ ;
  assign \new_[87142]_  = ~A233 & A232;
  assign \new_[87145]_  = A236 & A234;
  assign \new_[87146]_  = \new_[87145]_  & \new_[87142]_ ;
  assign \new_[87149]_  = ~A299 & A298;
  assign \new_[87152]_  = A301 & A300;
  assign \new_[87153]_  = \new_[87152]_  & \new_[87149]_ ;
  assign \new_[87154]_  = \new_[87153]_  & \new_[87146]_ ;
  assign \new_[87158]_  = ~A166 & ~A167;
  assign \new_[87159]_  = A170 & \new_[87158]_ ;
  assign \new_[87162]_  = ~A200 & A199;
  assign \new_[87165]_  = A202 & A201;
  assign \new_[87166]_  = \new_[87165]_  & \new_[87162]_ ;
  assign \new_[87167]_  = \new_[87166]_  & \new_[87159]_ ;
  assign \new_[87170]_  = ~A233 & A232;
  assign \new_[87173]_  = A236 & A234;
  assign \new_[87174]_  = \new_[87173]_  & \new_[87170]_ ;
  assign \new_[87177]_  = ~A299 & A298;
  assign \new_[87180]_  = A302 & A300;
  assign \new_[87181]_  = \new_[87180]_  & \new_[87177]_ ;
  assign \new_[87182]_  = \new_[87181]_  & \new_[87174]_ ;
  assign \new_[87186]_  = ~A166 & ~A167;
  assign \new_[87187]_  = A170 & \new_[87186]_ ;
  assign \new_[87190]_  = ~A200 & A199;
  assign \new_[87193]_  = A202 & A201;
  assign \new_[87194]_  = \new_[87193]_  & \new_[87190]_ ;
  assign \new_[87195]_  = \new_[87194]_  & \new_[87187]_ ;
  assign \new_[87198]_  = ~A233 & A232;
  assign \new_[87201]_  = A236 & A234;
  assign \new_[87202]_  = \new_[87201]_  & \new_[87198]_ ;
  assign \new_[87205]_  = ~A266 & A265;
  assign \new_[87208]_  = A268 & A267;
  assign \new_[87209]_  = \new_[87208]_  & \new_[87205]_ ;
  assign \new_[87210]_  = \new_[87209]_  & \new_[87202]_ ;
  assign \new_[87214]_  = ~A166 & ~A167;
  assign \new_[87215]_  = A170 & \new_[87214]_ ;
  assign \new_[87218]_  = ~A200 & A199;
  assign \new_[87221]_  = A202 & A201;
  assign \new_[87222]_  = \new_[87221]_  & \new_[87218]_ ;
  assign \new_[87223]_  = \new_[87222]_  & \new_[87215]_ ;
  assign \new_[87226]_  = ~A233 & A232;
  assign \new_[87229]_  = A236 & A234;
  assign \new_[87230]_  = \new_[87229]_  & \new_[87226]_ ;
  assign \new_[87233]_  = ~A266 & A265;
  assign \new_[87236]_  = A269 & A267;
  assign \new_[87237]_  = \new_[87236]_  & \new_[87233]_ ;
  assign \new_[87238]_  = \new_[87237]_  & \new_[87230]_ ;
  assign \new_[87242]_  = ~A166 & ~A167;
  assign \new_[87243]_  = A170 & \new_[87242]_ ;
  assign \new_[87246]_  = ~A200 & A199;
  assign \new_[87249]_  = A202 & A201;
  assign \new_[87250]_  = \new_[87249]_  & \new_[87246]_ ;
  assign \new_[87251]_  = \new_[87250]_  & \new_[87243]_ ;
  assign \new_[87254]_  = ~A233 & ~A232;
  assign \new_[87257]_  = ~A268 & ~A266;
  assign \new_[87258]_  = \new_[87257]_  & \new_[87254]_ ;
  assign \new_[87261]_  = A298 & ~A269;
  assign \new_[87264]_  = ~A302 & ~A301;
  assign \new_[87265]_  = \new_[87264]_  & \new_[87261]_ ;
  assign \new_[87266]_  = \new_[87265]_  & \new_[87258]_ ;
  assign \new_[87270]_  = ~A166 & ~A167;
  assign \new_[87271]_  = A170 & \new_[87270]_ ;
  assign \new_[87274]_  = ~A200 & A199;
  assign \new_[87277]_  = A203 & A201;
  assign \new_[87278]_  = \new_[87277]_  & \new_[87274]_ ;
  assign \new_[87279]_  = \new_[87278]_  & \new_[87271]_ ;
  assign \new_[87282]_  = A233 & A232;
  assign \new_[87285]_  = ~A268 & A265;
  assign \new_[87286]_  = \new_[87285]_  & \new_[87282]_ ;
  assign \new_[87289]_  = ~A299 & ~A269;
  assign \new_[87292]_  = ~A302 & ~A301;
  assign \new_[87293]_  = \new_[87292]_  & \new_[87289]_ ;
  assign \new_[87294]_  = \new_[87293]_  & \new_[87286]_ ;
  assign \new_[87298]_  = ~A166 & ~A167;
  assign \new_[87299]_  = A170 & \new_[87298]_ ;
  assign \new_[87302]_  = ~A200 & A199;
  assign \new_[87305]_  = A203 & A201;
  assign \new_[87306]_  = \new_[87305]_  & \new_[87302]_ ;
  assign \new_[87307]_  = \new_[87306]_  & \new_[87299]_ ;
  assign \new_[87310]_  = ~A235 & ~A233;
  assign \new_[87313]_  = A265 & ~A236;
  assign \new_[87314]_  = \new_[87313]_  & \new_[87310]_ ;
  assign \new_[87317]_  = A298 & A266;
  assign \new_[87320]_  = ~A302 & ~A301;
  assign \new_[87321]_  = \new_[87320]_  & \new_[87317]_ ;
  assign \new_[87322]_  = \new_[87321]_  & \new_[87314]_ ;
  assign \new_[87326]_  = ~A166 & ~A167;
  assign \new_[87327]_  = A170 & \new_[87326]_ ;
  assign \new_[87330]_  = ~A200 & A199;
  assign \new_[87333]_  = A203 & A201;
  assign \new_[87334]_  = \new_[87333]_  & \new_[87330]_ ;
  assign \new_[87335]_  = \new_[87334]_  & \new_[87327]_ ;
  assign \new_[87338]_  = ~A235 & ~A233;
  assign \new_[87341]_  = ~A266 & ~A236;
  assign \new_[87342]_  = \new_[87341]_  & \new_[87338]_ ;
  assign \new_[87345]_  = ~A269 & ~A268;
  assign \new_[87348]_  = ~A300 & A298;
  assign \new_[87349]_  = \new_[87348]_  & \new_[87345]_ ;
  assign \new_[87350]_  = \new_[87349]_  & \new_[87342]_ ;
  assign \new_[87354]_  = ~A166 & ~A167;
  assign \new_[87355]_  = A170 & \new_[87354]_ ;
  assign \new_[87358]_  = ~A200 & A199;
  assign \new_[87361]_  = A203 & A201;
  assign \new_[87362]_  = \new_[87361]_  & \new_[87358]_ ;
  assign \new_[87363]_  = \new_[87362]_  & \new_[87355]_ ;
  assign \new_[87366]_  = ~A235 & ~A233;
  assign \new_[87369]_  = ~A266 & ~A236;
  assign \new_[87370]_  = \new_[87369]_  & \new_[87366]_ ;
  assign \new_[87373]_  = ~A269 & ~A268;
  assign \new_[87376]_  = A299 & A298;
  assign \new_[87377]_  = \new_[87376]_  & \new_[87373]_ ;
  assign \new_[87378]_  = \new_[87377]_  & \new_[87370]_ ;
  assign \new_[87382]_  = ~A166 & ~A167;
  assign \new_[87383]_  = A170 & \new_[87382]_ ;
  assign \new_[87386]_  = ~A200 & A199;
  assign \new_[87389]_  = A203 & A201;
  assign \new_[87390]_  = \new_[87389]_  & \new_[87386]_ ;
  assign \new_[87391]_  = \new_[87390]_  & \new_[87383]_ ;
  assign \new_[87394]_  = ~A235 & ~A233;
  assign \new_[87397]_  = ~A266 & ~A236;
  assign \new_[87398]_  = \new_[87397]_  & \new_[87394]_ ;
  assign \new_[87401]_  = ~A269 & ~A268;
  assign \new_[87404]_  = ~A299 & ~A298;
  assign \new_[87405]_  = \new_[87404]_  & \new_[87401]_ ;
  assign \new_[87406]_  = \new_[87405]_  & \new_[87398]_ ;
  assign \new_[87410]_  = ~A166 & ~A167;
  assign \new_[87411]_  = A170 & \new_[87410]_ ;
  assign \new_[87414]_  = ~A200 & A199;
  assign \new_[87417]_  = A203 & A201;
  assign \new_[87418]_  = \new_[87417]_  & \new_[87414]_ ;
  assign \new_[87419]_  = \new_[87418]_  & \new_[87411]_ ;
  assign \new_[87422]_  = ~A235 & ~A233;
  assign \new_[87425]_  = ~A266 & ~A236;
  assign \new_[87426]_  = \new_[87425]_  & \new_[87422]_ ;
  assign \new_[87429]_  = A298 & ~A267;
  assign \new_[87432]_  = ~A302 & ~A301;
  assign \new_[87433]_  = \new_[87432]_  & \new_[87429]_ ;
  assign \new_[87434]_  = \new_[87433]_  & \new_[87426]_ ;
  assign \new_[87438]_  = ~A166 & ~A167;
  assign \new_[87439]_  = A170 & \new_[87438]_ ;
  assign \new_[87442]_  = ~A200 & A199;
  assign \new_[87445]_  = A203 & A201;
  assign \new_[87446]_  = \new_[87445]_  & \new_[87442]_ ;
  assign \new_[87447]_  = \new_[87446]_  & \new_[87439]_ ;
  assign \new_[87450]_  = ~A235 & ~A233;
  assign \new_[87453]_  = ~A265 & ~A236;
  assign \new_[87454]_  = \new_[87453]_  & \new_[87450]_ ;
  assign \new_[87457]_  = A298 & ~A266;
  assign \new_[87460]_  = ~A302 & ~A301;
  assign \new_[87461]_  = \new_[87460]_  & \new_[87457]_ ;
  assign \new_[87462]_  = \new_[87461]_  & \new_[87454]_ ;
  assign \new_[87466]_  = ~A166 & ~A167;
  assign \new_[87467]_  = A170 & \new_[87466]_ ;
  assign \new_[87470]_  = ~A200 & A199;
  assign \new_[87473]_  = A203 & A201;
  assign \new_[87474]_  = \new_[87473]_  & \new_[87470]_ ;
  assign \new_[87475]_  = \new_[87474]_  & \new_[87467]_ ;
  assign \new_[87478]_  = ~A234 & ~A233;
  assign \new_[87481]_  = ~A268 & ~A266;
  assign \new_[87482]_  = \new_[87481]_  & \new_[87478]_ ;
  assign \new_[87485]_  = A298 & ~A269;
  assign \new_[87488]_  = ~A302 & ~A301;
  assign \new_[87489]_  = \new_[87488]_  & \new_[87485]_ ;
  assign \new_[87490]_  = \new_[87489]_  & \new_[87482]_ ;
  assign \new_[87494]_  = ~A166 & ~A167;
  assign \new_[87495]_  = A170 & \new_[87494]_ ;
  assign \new_[87498]_  = ~A200 & A199;
  assign \new_[87501]_  = A203 & A201;
  assign \new_[87502]_  = \new_[87501]_  & \new_[87498]_ ;
  assign \new_[87503]_  = \new_[87502]_  & \new_[87495]_ ;
  assign \new_[87506]_  = ~A233 & A232;
  assign \new_[87509]_  = A235 & A234;
  assign \new_[87510]_  = \new_[87509]_  & \new_[87506]_ ;
  assign \new_[87513]_  = ~A299 & A298;
  assign \new_[87516]_  = A301 & A300;
  assign \new_[87517]_  = \new_[87516]_  & \new_[87513]_ ;
  assign \new_[87518]_  = \new_[87517]_  & \new_[87510]_ ;
  assign \new_[87522]_  = ~A166 & ~A167;
  assign \new_[87523]_  = A170 & \new_[87522]_ ;
  assign \new_[87526]_  = ~A200 & A199;
  assign \new_[87529]_  = A203 & A201;
  assign \new_[87530]_  = \new_[87529]_  & \new_[87526]_ ;
  assign \new_[87531]_  = \new_[87530]_  & \new_[87523]_ ;
  assign \new_[87534]_  = ~A233 & A232;
  assign \new_[87537]_  = A235 & A234;
  assign \new_[87538]_  = \new_[87537]_  & \new_[87534]_ ;
  assign \new_[87541]_  = ~A299 & A298;
  assign \new_[87544]_  = A302 & A300;
  assign \new_[87545]_  = \new_[87544]_  & \new_[87541]_ ;
  assign \new_[87546]_  = \new_[87545]_  & \new_[87538]_ ;
  assign \new_[87550]_  = ~A166 & ~A167;
  assign \new_[87551]_  = A170 & \new_[87550]_ ;
  assign \new_[87554]_  = ~A200 & A199;
  assign \new_[87557]_  = A203 & A201;
  assign \new_[87558]_  = \new_[87557]_  & \new_[87554]_ ;
  assign \new_[87559]_  = \new_[87558]_  & \new_[87551]_ ;
  assign \new_[87562]_  = ~A233 & A232;
  assign \new_[87565]_  = A235 & A234;
  assign \new_[87566]_  = \new_[87565]_  & \new_[87562]_ ;
  assign \new_[87569]_  = ~A266 & A265;
  assign \new_[87572]_  = A268 & A267;
  assign \new_[87573]_  = \new_[87572]_  & \new_[87569]_ ;
  assign \new_[87574]_  = \new_[87573]_  & \new_[87566]_ ;
  assign \new_[87578]_  = ~A166 & ~A167;
  assign \new_[87579]_  = A170 & \new_[87578]_ ;
  assign \new_[87582]_  = ~A200 & A199;
  assign \new_[87585]_  = A203 & A201;
  assign \new_[87586]_  = \new_[87585]_  & \new_[87582]_ ;
  assign \new_[87587]_  = \new_[87586]_  & \new_[87579]_ ;
  assign \new_[87590]_  = ~A233 & A232;
  assign \new_[87593]_  = A235 & A234;
  assign \new_[87594]_  = \new_[87593]_  & \new_[87590]_ ;
  assign \new_[87597]_  = ~A266 & A265;
  assign \new_[87600]_  = A269 & A267;
  assign \new_[87601]_  = \new_[87600]_  & \new_[87597]_ ;
  assign \new_[87602]_  = \new_[87601]_  & \new_[87594]_ ;
  assign \new_[87606]_  = ~A166 & ~A167;
  assign \new_[87607]_  = A170 & \new_[87606]_ ;
  assign \new_[87610]_  = ~A200 & A199;
  assign \new_[87613]_  = A203 & A201;
  assign \new_[87614]_  = \new_[87613]_  & \new_[87610]_ ;
  assign \new_[87615]_  = \new_[87614]_  & \new_[87607]_ ;
  assign \new_[87618]_  = ~A233 & A232;
  assign \new_[87621]_  = A236 & A234;
  assign \new_[87622]_  = \new_[87621]_  & \new_[87618]_ ;
  assign \new_[87625]_  = ~A299 & A298;
  assign \new_[87628]_  = A301 & A300;
  assign \new_[87629]_  = \new_[87628]_  & \new_[87625]_ ;
  assign \new_[87630]_  = \new_[87629]_  & \new_[87622]_ ;
  assign \new_[87634]_  = ~A166 & ~A167;
  assign \new_[87635]_  = A170 & \new_[87634]_ ;
  assign \new_[87638]_  = ~A200 & A199;
  assign \new_[87641]_  = A203 & A201;
  assign \new_[87642]_  = \new_[87641]_  & \new_[87638]_ ;
  assign \new_[87643]_  = \new_[87642]_  & \new_[87635]_ ;
  assign \new_[87646]_  = ~A233 & A232;
  assign \new_[87649]_  = A236 & A234;
  assign \new_[87650]_  = \new_[87649]_  & \new_[87646]_ ;
  assign \new_[87653]_  = ~A299 & A298;
  assign \new_[87656]_  = A302 & A300;
  assign \new_[87657]_  = \new_[87656]_  & \new_[87653]_ ;
  assign \new_[87658]_  = \new_[87657]_  & \new_[87650]_ ;
  assign \new_[87662]_  = ~A166 & ~A167;
  assign \new_[87663]_  = A170 & \new_[87662]_ ;
  assign \new_[87666]_  = ~A200 & A199;
  assign \new_[87669]_  = A203 & A201;
  assign \new_[87670]_  = \new_[87669]_  & \new_[87666]_ ;
  assign \new_[87671]_  = \new_[87670]_  & \new_[87663]_ ;
  assign \new_[87674]_  = ~A233 & A232;
  assign \new_[87677]_  = A236 & A234;
  assign \new_[87678]_  = \new_[87677]_  & \new_[87674]_ ;
  assign \new_[87681]_  = ~A266 & A265;
  assign \new_[87684]_  = A268 & A267;
  assign \new_[87685]_  = \new_[87684]_  & \new_[87681]_ ;
  assign \new_[87686]_  = \new_[87685]_  & \new_[87678]_ ;
  assign \new_[87690]_  = ~A166 & ~A167;
  assign \new_[87691]_  = A170 & \new_[87690]_ ;
  assign \new_[87694]_  = ~A200 & A199;
  assign \new_[87697]_  = A203 & A201;
  assign \new_[87698]_  = \new_[87697]_  & \new_[87694]_ ;
  assign \new_[87699]_  = \new_[87698]_  & \new_[87691]_ ;
  assign \new_[87702]_  = ~A233 & A232;
  assign \new_[87705]_  = A236 & A234;
  assign \new_[87706]_  = \new_[87705]_  & \new_[87702]_ ;
  assign \new_[87709]_  = ~A266 & A265;
  assign \new_[87712]_  = A269 & A267;
  assign \new_[87713]_  = \new_[87712]_  & \new_[87709]_ ;
  assign \new_[87714]_  = \new_[87713]_  & \new_[87706]_ ;
  assign \new_[87718]_  = ~A166 & ~A167;
  assign \new_[87719]_  = A170 & \new_[87718]_ ;
  assign \new_[87722]_  = ~A200 & A199;
  assign \new_[87725]_  = A203 & A201;
  assign \new_[87726]_  = \new_[87725]_  & \new_[87722]_ ;
  assign \new_[87727]_  = \new_[87726]_  & \new_[87719]_ ;
  assign \new_[87730]_  = ~A233 & ~A232;
  assign \new_[87733]_  = ~A268 & ~A266;
  assign \new_[87734]_  = \new_[87733]_  & \new_[87730]_ ;
  assign \new_[87737]_  = A298 & ~A269;
  assign \new_[87740]_  = ~A302 & ~A301;
  assign \new_[87741]_  = \new_[87740]_  & \new_[87737]_ ;
  assign \new_[87742]_  = \new_[87741]_  & \new_[87734]_ ;
  assign \new_[87746]_  = A167 & ~A168;
  assign \new_[87747]_  = A170 & \new_[87746]_ ;
  assign \new_[87750]_  = ~A199 & A166;
  assign \new_[87753]_  = ~A233 & A200;
  assign \new_[87754]_  = \new_[87753]_  & \new_[87750]_ ;
  assign \new_[87755]_  = \new_[87754]_  & \new_[87747]_ ;
  assign \new_[87758]_  = ~A236 & ~A235;
  assign \new_[87761]_  = ~A268 & ~A266;
  assign \new_[87762]_  = \new_[87761]_  & \new_[87758]_ ;
  assign \new_[87765]_  = A298 & ~A269;
  assign \new_[87768]_  = ~A302 & ~A301;
  assign \new_[87769]_  = \new_[87768]_  & \new_[87765]_ ;
  assign \new_[87770]_  = \new_[87769]_  & \new_[87762]_ ;
  assign \new_[87774]_  = A167 & ~A168;
  assign \new_[87775]_  = ~A170 & \new_[87774]_ ;
  assign \new_[87778]_  = ~A199 & ~A166;
  assign \new_[87781]_  = ~A233 & A200;
  assign \new_[87782]_  = \new_[87781]_  & \new_[87778]_ ;
  assign \new_[87783]_  = \new_[87782]_  & \new_[87775]_ ;
  assign \new_[87786]_  = ~A236 & ~A235;
  assign \new_[87789]_  = ~A268 & ~A266;
  assign \new_[87790]_  = \new_[87789]_  & \new_[87786]_ ;
  assign \new_[87793]_  = A298 & ~A269;
  assign \new_[87796]_  = ~A302 & ~A301;
  assign \new_[87797]_  = \new_[87796]_  & \new_[87793]_ ;
  assign \new_[87798]_  = \new_[87797]_  & \new_[87790]_ ;
  assign \new_[87802]_  = ~A167 & ~A168;
  assign \new_[87803]_  = ~A170 & \new_[87802]_ ;
  assign \new_[87806]_  = ~A199 & A166;
  assign \new_[87809]_  = ~A233 & A200;
  assign \new_[87810]_  = \new_[87809]_  & \new_[87806]_ ;
  assign \new_[87811]_  = \new_[87810]_  & \new_[87803]_ ;
  assign \new_[87814]_  = ~A236 & ~A235;
  assign \new_[87817]_  = ~A268 & ~A266;
  assign \new_[87818]_  = \new_[87817]_  & \new_[87814]_ ;
  assign \new_[87821]_  = A298 & ~A269;
  assign \new_[87824]_  = ~A302 & ~A301;
  assign \new_[87825]_  = \new_[87824]_  & \new_[87821]_ ;
  assign \new_[87826]_  = \new_[87825]_  & \new_[87818]_ ;
  assign \new_[87830]_  = A167 & ~A168;
  assign \new_[87831]_  = A169 & \new_[87830]_ ;
  assign \new_[87834]_  = ~A199 & ~A166;
  assign \new_[87837]_  = ~A233 & A200;
  assign \new_[87838]_  = \new_[87837]_  & \new_[87834]_ ;
  assign \new_[87839]_  = \new_[87838]_  & \new_[87831]_ ;
  assign \new_[87842]_  = ~A236 & ~A235;
  assign \new_[87845]_  = ~A268 & ~A266;
  assign \new_[87846]_  = \new_[87845]_  & \new_[87842]_ ;
  assign \new_[87849]_  = A298 & ~A269;
  assign \new_[87852]_  = ~A302 & ~A301;
  assign \new_[87853]_  = \new_[87852]_  & \new_[87849]_ ;
  assign \new_[87854]_  = \new_[87853]_  & \new_[87846]_ ;
  assign \new_[87858]_  = A167 & ~A168;
  assign \new_[87859]_  = A169 & \new_[87858]_ ;
  assign \new_[87862]_  = A199 & ~A166;
  assign \new_[87865]_  = A201 & ~A200;
  assign \new_[87866]_  = \new_[87865]_  & \new_[87862]_ ;
  assign \new_[87867]_  = \new_[87866]_  & \new_[87859]_ ;
  assign \new_[87870]_  = A232 & A202;
  assign \new_[87873]_  = A265 & A233;
  assign \new_[87874]_  = \new_[87873]_  & \new_[87870]_ ;
  assign \new_[87877]_  = ~A269 & ~A268;
  assign \new_[87880]_  = ~A300 & ~A299;
  assign \new_[87881]_  = \new_[87880]_  & \new_[87877]_ ;
  assign \new_[87882]_  = \new_[87881]_  & \new_[87874]_ ;
  assign \new_[87886]_  = A167 & ~A168;
  assign \new_[87887]_  = A169 & \new_[87886]_ ;
  assign \new_[87890]_  = A199 & ~A166;
  assign \new_[87893]_  = A201 & ~A200;
  assign \new_[87894]_  = \new_[87893]_  & \new_[87890]_ ;
  assign \new_[87895]_  = \new_[87894]_  & \new_[87887]_ ;
  assign \new_[87898]_  = A232 & A202;
  assign \new_[87901]_  = A265 & A233;
  assign \new_[87902]_  = \new_[87901]_  & \new_[87898]_ ;
  assign \new_[87905]_  = ~A269 & ~A268;
  assign \new_[87908]_  = A299 & A298;
  assign \new_[87909]_  = \new_[87908]_  & \new_[87905]_ ;
  assign \new_[87910]_  = \new_[87909]_  & \new_[87902]_ ;
  assign \new_[87914]_  = A167 & ~A168;
  assign \new_[87915]_  = A169 & \new_[87914]_ ;
  assign \new_[87918]_  = A199 & ~A166;
  assign \new_[87921]_  = A201 & ~A200;
  assign \new_[87922]_  = \new_[87921]_  & \new_[87918]_ ;
  assign \new_[87923]_  = \new_[87922]_  & \new_[87915]_ ;
  assign \new_[87926]_  = A232 & A202;
  assign \new_[87929]_  = A265 & A233;
  assign \new_[87930]_  = \new_[87929]_  & \new_[87926]_ ;
  assign \new_[87933]_  = ~A269 & ~A268;
  assign \new_[87936]_  = ~A299 & ~A298;
  assign \new_[87937]_  = \new_[87936]_  & \new_[87933]_ ;
  assign \new_[87938]_  = \new_[87937]_  & \new_[87930]_ ;
  assign \new_[87942]_  = A167 & ~A168;
  assign \new_[87943]_  = A169 & \new_[87942]_ ;
  assign \new_[87946]_  = A199 & ~A166;
  assign \new_[87949]_  = A201 & ~A200;
  assign \new_[87950]_  = \new_[87949]_  & \new_[87946]_ ;
  assign \new_[87951]_  = \new_[87950]_  & \new_[87943]_ ;
  assign \new_[87954]_  = A232 & A202;
  assign \new_[87957]_  = A265 & A233;
  assign \new_[87958]_  = \new_[87957]_  & \new_[87954]_ ;
  assign \new_[87961]_  = ~A299 & ~A267;
  assign \new_[87964]_  = ~A302 & ~A301;
  assign \new_[87965]_  = \new_[87964]_  & \new_[87961]_ ;
  assign \new_[87966]_  = \new_[87965]_  & \new_[87958]_ ;
  assign \new_[87970]_  = A167 & ~A168;
  assign \new_[87971]_  = A169 & \new_[87970]_ ;
  assign \new_[87974]_  = A199 & ~A166;
  assign \new_[87977]_  = A201 & ~A200;
  assign \new_[87978]_  = \new_[87977]_  & \new_[87974]_ ;
  assign \new_[87979]_  = \new_[87978]_  & \new_[87971]_ ;
  assign \new_[87982]_  = A232 & A202;
  assign \new_[87985]_  = A265 & A233;
  assign \new_[87986]_  = \new_[87985]_  & \new_[87982]_ ;
  assign \new_[87989]_  = ~A299 & A266;
  assign \new_[87992]_  = ~A302 & ~A301;
  assign \new_[87993]_  = \new_[87992]_  & \new_[87989]_ ;
  assign \new_[87994]_  = \new_[87993]_  & \new_[87986]_ ;
  assign \new_[87998]_  = A167 & ~A168;
  assign \new_[87999]_  = A169 & \new_[87998]_ ;
  assign \new_[88002]_  = A199 & ~A166;
  assign \new_[88005]_  = A201 & ~A200;
  assign \new_[88006]_  = \new_[88005]_  & \new_[88002]_ ;
  assign \new_[88007]_  = \new_[88006]_  & \new_[87999]_ ;
  assign \new_[88010]_  = A232 & A202;
  assign \new_[88013]_  = ~A265 & A233;
  assign \new_[88014]_  = \new_[88013]_  & \new_[88010]_ ;
  assign \new_[88017]_  = ~A299 & ~A266;
  assign \new_[88020]_  = ~A302 & ~A301;
  assign \new_[88021]_  = \new_[88020]_  & \new_[88017]_ ;
  assign \new_[88022]_  = \new_[88021]_  & \new_[88014]_ ;
  assign \new_[88026]_  = A167 & ~A168;
  assign \new_[88027]_  = A169 & \new_[88026]_ ;
  assign \new_[88030]_  = A199 & ~A166;
  assign \new_[88033]_  = A201 & ~A200;
  assign \new_[88034]_  = \new_[88033]_  & \new_[88030]_ ;
  assign \new_[88035]_  = \new_[88034]_  & \new_[88027]_ ;
  assign \new_[88038]_  = ~A233 & A202;
  assign \new_[88041]_  = ~A236 & ~A235;
  assign \new_[88042]_  = \new_[88041]_  & \new_[88038]_ ;
  assign \new_[88045]_  = A266 & A265;
  assign \new_[88048]_  = ~A300 & A298;
  assign \new_[88049]_  = \new_[88048]_  & \new_[88045]_ ;
  assign \new_[88050]_  = \new_[88049]_  & \new_[88042]_ ;
  assign \new_[88054]_  = A167 & ~A168;
  assign \new_[88055]_  = A169 & \new_[88054]_ ;
  assign \new_[88058]_  = A199 & ~A166;
  assign \new_[88061]_  = A201 & ~A200;
  assign \new_[88062]_  = \new_[88061]_  & \new_[88058]_ ;
  assign \new_[88063]_  = \new_[88062]_  & \new_[88055]_ ;
  assign \new_[88066]_  = ~A233 & A202;
  assign \new_[88069]_  = ~A236 & ~A235;
  assign \new_[88070]_  = \new_[88069]_  & \new_[88066]_ ;
  assign \new_[88073]_  = A266 & A265;
  assign \new_[88076]_  = A299 & A298;
  assign \new_[88077]_  = \new_[88076]_  & \new_[88073]_ ;
  assign \new_[88078]_  = \new_[88077]_  & \new_[88070]_ ;
  assign \new_[88082]_  = A167 & ~A168;
  assign \new_[88083]_  = A169 & \new_[88082]_ ;
  assign \new_[88086]_  = A199 & ~A166;
  assign \new_[88089]_  = A201 & ~A200;
  assign \new_[88090]_  = \new_[88089]_  & \new_[88086]_ ;
  assign \new_[88091]_  = \new_[88090]_  & \new_[88083]_ ;
  assign \new_[88094]_  = ~A233 & A202;
  assign \new_[88097]_  = ~A236 & ~A235;
  assign \new_[88098]_  = \new_[88097]_  & \new_[88094]_ ;
  assign \new_[88101]_  = A266 & A265;
  assign \new_[88104]_  = ~A299 & ~A298;
  assign \new_[88105]_  = \new_[88104]_  & \new_[88101]_ ;
  assign \new_[88106]_  = \new_[88105]_  & \new_[88098]_ ;
  assign \new_[88110]_  = A167 & ~A168;
  assign \new_[88111]_  = A169 & \new_[88110]_ ;
  assign \new_[88114]_  = A199 & ~A166;
  assign \new_[88117]_  = A201 & ~A200;
  assign \new_[88118]_  = \new_[88117]_  & \new_[88114]_ ;
  assign \new_[88119]_  = \new_[88118]_  & \new_[88111]_ ;
  assign \new_[88122]_  = ~A233 & A202;
  assign \new_[88125]_  = ~A236 & ~A235;
  assign \new_[88126]_  = \new_[88125]_  & \new_[88122]_ ;
  assign \new_[88129]_  = ~A267 & ~A266;
  assign \new_[88132]_  = ~A300 & A298;
  assign \new_[88133]_  = \new_[88132]_  & \new_[88129]_ ;
  assign \new_[88134]_  = \new_[88133]_  & \new_[88126]_ ;
  assign \new_[88138]_  = A167 & ~A168;
  assign \new_[88139]_  = A169 & \new_[88138]_ ;
  assign \new_[88142]_  = A199 & ~A166;
  assign \new_[88145]_  = A201 & ~A200;
  assign \new_[88146]_  = \new_[88145]_  & \new_[88142]_ ;
  assign \new_[88147]_  = \new_[88146]_  & \new_[88139]_ ;
  assign \new_[88150]_  = ~A233 & A202;
  assign \new_[88153]_  = ~A236 & ~A235;
  assign \new_[88154]_  = \new_[88153]_  & \new_[88150]_ ;
  assign \new_[88157]_  = ~A267 & ~A266;
  assign \new_[88160]_  = A299 & A298;
  assign \new_[88161]_  = \new_[88160]_  & \new_[88157]_ ;
  assign \new_[88162]_  = \new_[88161]_  & \new_[88154]_ ;
  assign \new_[88166]_  = A167 & ~A168;
  assign \new_[88167]_  = A169 & \new_[88166]_ ;
  assign \new_[88170]_  = A199 & ~A166;
  assign \new_[88173]_  = A201 & ~A200;
  assign \new_[88174]_  = \new_[88173]_  & \new_[88170]_ ;
  assign \new_[88175]_  = \new_[88174]_  & \new_[88167]_ ;
  assign \new_[88178]_  = ~A233 & A202;
  assign \new_[88181]_  = ~A236 & ~A235;
  assign \new_[88182]_  = \new_[88181]_  & \new_[88178]_ ;
  assign \new_[88185]_  = ~A267 & ~A266;
  assign \new_[88188]_  = ~A299 & ~A298;
  assign \new_[88189]_  = \new_[88188]_  & \new_[88185]_ ;
  assign \new_[88190]_  = \new_[88189]_  & \new_[88182]_ ;
  assign \new_[88194]_  = A167 & ~A168;
  assign \new_[88195]_  = A169 & \new_[88194]_ ;
  assign \new_[88198]_  = A199 & ~A166;
  assign \new_[88201]_  = A201 & ~A200;
  assign \new_[88202]_  = \new_[88201]_  & \new_[88198]_ ;
  assign \new_[88203]_  = \new_[88202]_  & \new_[88195]_ ;
  assign \new_[88206]_  = ~A233 & A202;
  assign \new_[88209]_  = ~A236 & ~A235;
  assign \new_[88210]_  = \new_[88209]_  & \new_[88206]_ ;
  assign \new_[88213]_  = ~A266 & ~A265;
  assign \new_[88216]_  = ~A300 & A298;
  assign \new_[88217]_  = \new_[88216]_  & \new_[88213]_ ;
  assign \new_[88218]_  = \new_[88217]_  & \new_[88210]_ ;
  assign \new_[88222]_  = A167 & ~A168;
  assign \new_[88223]_  = A169 & \new_[88222]_ ;
  assign \new_[88226]_  = A199 & ~A166;
  assign \new_[88229]_  = A201 & ~A200;
  assign \new_[88230]_  = \new_[88229]_  & \new_[88226]_ ;
  assign \new_[88231]_  = \new_[88230]_  & \new_[88223]_ ;
  assign \new_[88234]_  = ~A233 & A202;
  assign \new_[88237]_  = ~A236 & ~A235;
  assign \new_[88238]_  = \new_[88237]_  & \new_[88234]_ ;
  assign \new_[88241]_  = ~A266 & ~A265;
  assign \new_[88244]_  = A299 & A298;
  assign \new_[88245]_  = \new_[88244]_  & \new_[88241]_ ;
  assign \new_[88246]_  = \new_[88245]_  & \new_[88238]_ ;
  assign \new_[88250]_  = A167 & ~A168;
  assign \new_[88251]_  = A169 & \new_[88250]_ ;
  assign \new_[88254]_  = A199 & ~A166;
  assign \new_[88257]_  = A201 & ~A200;
  assign \new_[88258]_  = \new_[88257]_  & \new_[88254]_ ;
  assign \new_[88259]_  = \new_[88258]_  & \new_[88251]_ ;
  assign \new_[88262]_  = ~A233 & A202;
  assign \new_[88265]_  = ~A236 & ~A235;
  assign \new_[88266]_  = \new_[88265]_  & \new_[88262]_ ;
  assign \new_[88269]_  = ~A266 & ~A265;
  assign \new_[88272]_  = ~A299 & ~A298;
  assign \new_[88273]_  = \new_[88272]_  & \new_[88269]_ ;
  assign \new_[88274]_  = \new_[88273]_  & \new_[88266]_ ;
  assign \new_[88278]_  = A167 & ~A168;
  assign \new_[88279]_  = A169 & \new_[88278]_ ;
  assign \new_[88282]_  = A199 & ~A166;
  assign \new_[88285]_  = A201 & ~A200;
  assign \new_[88286]_  = \new_[88285]_  & \new_[88282]_ ;
  assign \new_[88287]_  = \new_[88286]_  & \new_[88279]_ ;
  assign \new_[88290]_  = ~A233 & A202;
  assign \new_[88293]_  = A265 & ~A234;
  assign \new_[88294]_  = \new_[88293]_  & \new_[88290]_ ;
  assign \new_[88297]_  = A298 & A266;
  assign \new_[88300]_  = ~A302 & ~A301;
  assign \new_[88301]_  = \new_[88300]_  & \new_[88297]_ ;
  assign \new_[88302]_  = \new_[88301]_  & \new_[88294]_ ;
  assign \new_[88306]_  = A167 & ~A168;
  assign \new_[88307]_  = A169 & \new_[88306]_ ;
  assign \new_[88310]_  = A199 & ~A166;
  assign \new_[88313]_  = A201 & ~A200;
  assign \new_[88314]_  = \new_[88313]_  & \new_[88310]_ ;
  assign \new_[88315]_  = \new_[88314]_  & \new_[88307]_ ;
  assign \new_[88318]_  = ~A233 & A202;
  assign \new_[88321]_  = ~A266 & ~A234;
  assign \new_[88322]_  = \new_[88321]_  & \new_[88318]_ ;
  assign \new_[88325]_  = ~A269 & ~A268;
  assign \new_[88328]_  = ~A300 & A298;
  assign \new_[88329]_  = \new_[88328]_  & \new_[88325]_ ;
  assign \new_[88330]_  = \new_[88329]_  & \new_[88322]_ ;
  assign \new_[88334]_  = A167 & ~A168;
  assign \new_[88335]_  = A169 & \new_[88334]_ ;
  assign \new_[88338]_  = A199 & ~A166;
  assign \new_[88341]_  = A201 & ~A200;
  assign \new_[88342]_  = \new_[88341]_  & \new_[88338]_ ;
  assign \new_[88343]_  = \new_[88342]_  & \new_[88335]_ ;
  assign \new_[88346]_  = ~A233 & A202;
  assign \new_[88349]_  = ~A266 & ~A234;
  assign \new_[88350]_  = \new_[88349]_  & \new_[88346]_ ;
  assign \new_[88353]_  = ~A269 & ~A268;
  assign \new_[88356]_  = A299 & A298;
  assign \new_[88357]_  = \new_[88356]_  & \new_[88353]_ ;
  assign \new_[88358]_  = \new_[88357]_  & \new_[88350]_ ;
  assign \new_[88362]_  = A167 & ~A168;
  assign \new_[88363]_  = A169 & \new_[88362]_ ;
  assign \new_[88366]_  = A199 & ~A166;
  assign \new_[88369]_  = A201 & ~A200;
  assign \new_[88370]_  = \new_[88369]_  & \new_[88366]_ ;
  assign \new_[88371]_  = \new_[88370]_  & \new_[88363]_ ;
  assign \new_[88374]_  = ~A233 & A202;
  assign \new_[88377]_  = ~A266 & ~A234;
  assign \new_[88378]_  = \new_[88377]_  & \new_[88374]_ ;
  assign \new_[88381]_  = ~A269 & ~A268;
  assign \new_[88384]_  = ~A299 & ~A298;
  assign \new_[88385]_  = \new_[88384]_  & \new_[88381]_ ;
  assign \new_[88386]_  = \new_[88385]_  & \new_[88378]_ ;
  assign \new_[88390]_  = A167 & ~A168;
  assign \new_[88391]_  = A169 & \new_[88390]_ ;
  assign \new_[88394]_  = A199 & ~A166;
  assign \new_[88397]_  = A201 & ~A200;
  assign \new_[88398]_  = \new_[88397]_  & \new_[88394]_ ;
  assign \new_[88399]_  = \new_[88398]_  & \new_[88391]_ ;
  assign \new_[88402]_  = ~A233 & A202;
  assign \new_[88405]_  = ~A266 & ~A234;
  assign \new_[88406]_  = \new_[88405]_  & \new_[88402]_ ;
  assign \new_[88409]_  = A298 & ~A267;
  assign \new_[88412]_  = ~A302 & ~A301;
  assign \new_[88413]_  = \new_[88412]_  & \new_[88409]_ ;
  assign \new_[88414]_  = \new_[88413]_  & \new_[88406]_ ;
  assign \new_[88418]_  = A167 & ~A168;
  assign \new_[88419]_  = A169 & \new_[88418]_ ;
  assign \new_[88422]_  = A199 & ~A166;
  assign \new_[88425]_  = A201 & ~A200;
  assign \new_[88426]_  = \new_[88425]_  & \new_[88422]_ ;
  assign \new_[88427]_  = \new_[88426]_  & \new_[88419]_ ;
  assign \new_[88430]_  = ~A233 & A202;
  assign \new_[88433]_  = ~A265 & ~A234;
  assign \new_[88434]_  = \new_[88433]_  & \new_[88430]_ ;
  assign \new_[88437]_  = A298 & ~A266;
  assign \new_[88440]_  = ~A302 & ~A301;
  assign \new_[88441]_  = \new_[88440]_  & \new_[88437]_ ;
  assign \new_[88442]_  = \new_[88441]_  & \new_[88434]_ ;
  assign \new_[88446]_  = A167 & ~A168;
  assign \new_[88447]_  = A169 & \new_[88446]_ ;
  assign \new_[88450]_  = A199 & ~A166;
  assign \new_[88453]_  = A201 & ~A200;
  assign \new_[88454]_  = \new_[88453]_  & \new_[88450]_ ;
  assign \new_[88455]_  = \new_[88454]_  & \new_[88447]_ ;
  assign \new_[88458]_  = ~A232 & A202;
  assign \new_[88461]_  = A265 & ~A233;
  assign \new_[88462]_  = \new_[88461]_  & \new_[88458]_ ;
  assign \new_[88465]_  = A298 & A266;
  assign \new_[88468]_  = ~A302 & ~A301;
  assign \new_[88469]_  = \new_[88468]_  & \new_[88465]_ ;
  assign \new_[88470]_  = \new_[88469]_  & \new_[88462]_ ;
  assign \new_[88474]_  = A167 & ~A168;
  assign \new_[88475]_  = A169 & \new_[88474]_ ;
  assign \new_[88478]_  = A199 & ~A166;
  assign \new_[88481]_  = A201 & ~A200;
  assign \new_[88482]_  = \new_[88481]_  & \new_[88478]_ ;
  assign \new_[88483]_  = \new_[88482]_  & \new_[88475]_ ;
  assign \new_[88486]_  = ~A232 & A202;
  assign \new_[88489]_  = ~A266 & ~A233;
  assign \new_[88490]_  = \new_[88489]_  & \new_[88486]_ ;
  assign \new_[88493]_  = ~A269 & ~A268;
  assign \new_[88496]_  = ~A300 & A298;
  assign \new_[88497]_  = \new_[88496]_  & \new_[88493]_ ;
  assign \new_[88498]_  = \new_[88497]_  & \new_[88490]_ ;
  assign \new_[88502]_  = A167 & ~A168;
  assign \new_[88503]_  = A169 & \new_[88502]_ ;
  assign \new_[88506]_  = A199 & ~A166;
  assign \new_[88509]_  = A201 & ~A200;
  assign \new_[88510]_  = \new_[88509]_  & \new_[88506]_ ;
  assign \new_[88511]_  = \new_[88510]_  & \new_[88503]_ ;
  assign \new_[88514]_  = ~A232 & A202;
  assign \new_[88517]_  = ~A266 & ~A233;
  assign \new_[88518]_  = \new_[88517]_  & \new_[88514]_ ;
  assign \new_[88521]_  = ~A269 & ~A268;
  assign \new_[88524]_  = A299 & A298;
  assign \new_[88525]_  = \new_[88524]_  & \new_[88521]_ ;
  assign \new_[88526]_  = \new_[88525]_  & \new_[88518]_ ;
  assign \new_[88530]_  = A167 & ~A168;
  assign \new_[88531]_  = A169 & \new_[88530]_ ;
  assign \new_[88534]_  = A199 & ~A166;
  assign \new_[88537]_  = A201 & ~A200;
  assign \new_[88538]_  = \new_[88537]_  & \new_[88534]_ ;
  assign \new_[88539]_  = \new_[88538]_  & \new_[88531]_ ;
  assign \new_[88542]_  = ~A232 & A202;
  assign \new_[88545]_  = ~A266 & ~A233;
  assign \new_[88546]_  = \new_[88545]_  & \new_[88542]_ ;
  assign \new_[88549]_  = ~A269 & ~A268;
  assign \new_[88552]_  = ~A299 & ~A298;
  assign \new_[88553]_  = \new_[88552]_  & \new_[88549]_ ;
  assign \new_[88554]_  = \new_[88553]_  & \new_[88546]_ ;
  assign \new_[88558]_  = A167 & ~A168;
  assign \new_[88559]_  = A169 & \new_[88558]_ ;
  assign \new_[88562]_  = A199 & ~A166;
  assign \new_[88565]_  = A201 & ~A200;
  assign \new_[88566]_  = \new_[88565]_  & \new_[88562]_ ;
  assign \new_[88567]_  = \new_[88566]_  & \new_[88559]_ ;
  assign \new_[88570]_  = ~A232 & A202;
  assign \new_[88573]_  = ~A266 & ~A233;
  assign \new_[88574]_  = \new_[88573]_  & \new_[88570]_ ;
  assign \new_[88577]_  = A298 & ~A267;
  assign \new_[88580]_  = ~A302 & ~A301;
  assign \new_[88581]_  = \new_[88580]_  & \new_[88577]_ ;
  assign \new_[88582]_  = \new_[88581]_  & \new_[88574]_ ;
  assign \new_[88586]_  = A167 & ~A168;
  assign \new_[88587]_  = A169 & \new_[88586]_ ;
  assign \new_[88590]_  = A199 & ~A166;
  assign \new_[88593]_  = A201 & ~A200;
  assign \new_[88594]_  = \new_[88593]_  & \new_[88590]_ ;
  assign \new_[88595]_  = \new_[88594]_  & \new_[88587]_ ;
  assign \new_[88598]_  = ~A232 & A202;
  assign \new_[88601]_  = ~A265 & ~A233;
  assign \new_[88602]_  = \new_[88601]_  & \new_[88598]_ ;
  assign \new_[88605]_  = A298 & ~A266;
  assign \new_[88608]_  = ~A302 & ~A301;
  assign \new_[88609]_  = \new_[88608]_  & \new_[88605]_ ;
  assign \new_[88610]_  = \new_[88609]_  & \new_[88602]_ ;
  assign \new_[88614]_  = A167 & ~A168;
  assign \new_[88615]_  = A169 & \new_[88614]_ ;
  assign \new_[88618]_  = A199 & ~A166;
  assign \new_[88621]_  = A201 & ~A200;
  assign \new_[88622]_  = \new_[88621]_  & \new_[88618]_ ;
  assign \new_[88623]_  = \new_[88622]_  & \new_[88615]_ ;
  assign \new_[88626]_  = A232 & A203;
  assign \new_[88629]_  = A265 & A233;
  assign \new_[88630]_  = \new_[88629]_  & \new_[88626]_ ;
  assign \new_[88633]_  = ~A269 & ~A268;
  assign \new_[88636]_  = ~A300 & ~A299;
  assign \new_[88637]_  = \new_[88636]_  & \new_[88633]_ ;
  assign \new_[88638]_  = \new_[88637]_  & \new_[88630]_ ;
  assign \new_[88642]_  = A167 & ~A168;
  assign \new_[88643]_  = A169 & \new_[88642]_ ;
  assign \new_[88646]_  = A199 & ~A166;
  assign \new_[88649]_  = A201 & ~A200;
  assign \new_[88650]_  = \new_[88649]_  & \new_[88646]_ ;
  assign \new_[88651]_  = \new_[88650]_  & \new_[88643]_ ;
  assign \new_[88654]_  = A232 & A203;
  assign \new_[88657]_  = A265 & A233;
  assign \new_[88658]_  = \new_[88657]_  & \new_[88654]_ ;
  assign \new_[88661]_  = ~A269 & ~A268;
  assign \new_[88664]_  = A299 & A298;
  assign \new_[88665]_  = \new_[88664]_  & \new_[88661]_ ;
  assign \new_[88666]_  = \new_[88665]_  & \new_[88658]_ ;
  assign \new_[88670]_  = A167 & ~A168;
  assign \new_[88671]_  = A169 & \new_[88670]_ ;
  assign \new_[88674]_  = A199 & ~A166;
  assign \new_[88677]_  = A201 & ~A200;
  assign \new_[88678]_  = \new_[88677]_  & \new_[88674]_ ;
  assign \new_[88679]_  = \new_[88678]_  & \new_[88671]_ ;
  assign \new_[88682]_  = A232 & A203;
  assign \new_[88685]_  = A265 & A233;
  assign \new_[88686]_  = \new_[88685]_  & \new_[88682]_ ;
  assign \new_[88689]_  = ~A269 & ~A268;
  assign \new_[88692]_  = ~A299 & ~A298;
  assign \new_[88693]_  = \new_[88692]_  & \new_[88689]_ ;
  assign \new_[88694]_  = \new_[88693]_  & \new_[88686]_ ;
  assign \new_[88698]_  = A167 & ~A168;
  assign \new_[88699]_  = A169 & \new_[88698]_ ;
  assign \new_[88702]_  = A199 & ~A166;
  assign \new_[88705]_  = A201 & ~A200;
  assign \new_[88706]_  = \new_[88705]_  & \new_[88702]_ ;
  assign \new_[88707]_  = \new_[88706]_  & \new_[88699]_ ;
  assign \new_[88710]_  = A232 & A203;
  assign \new_[88713]_  = A265 & A233;
  assign \new_[88714]_  = \new_[88713]_  & \new_[88710]_ ;
  assign \new_[88717]_  = ~A299 & ~A267;
  assign \new_[88720]_  = ~A302 & ~A301;
  assign \new_[88721]_  = \new_[88720]_  & \new_[88717]_ ;
  assign \new_[88722]_  = \new_[88721]_  & \new_[88714]_ ;
  assign \new_[88726]_  = A167 & ~A168;
  assign \new_[88727]_  = A169 & \new_[88726]_ ;
  assign \new_[88730]_  = A199 & ~A166;
  assign \new_[88733]_  = A201 & ~A200;
  assign \new_[88734]_  = \new_[88733]_  & \new_[88730]_ ;
  assign \new_[88735]_  = \new_[88734]_  & \new_[88727]_ ;
  assign \new_[88738]_  = A232 & A203;
  assign \new_[88741]_  = A265 & A233;
  assign \new_[88742]_  = \new_[88741]_  & \new_[88738]_ ;
  assign \new_[88745]_  = ~A299 & A266;
  assign \new_[88748]_  = ~A302 & ~A301;
  assign \new_[88749]_  = \new_[88748]_  & \new_[88745]_ ;
  assign \new_[88750]_  = \new_[88749]_  & \new_[88742]_ ;
  assign \new_[88754]_  = A167 & ~A168;
  assign \new_[88755]_  = A169 & \new_[88754]_ ;
  assign \new_[88758]_  = A199 & ~A166;
  assign \new_[88761]_  = A201 & ~A200;
  assign \new_[88762]_  = \new_[88761]_  & \new_[88758]_ ;
  assign \new_[88763]_  = \new_[88762]_  & \new_[88755]_ ;
  assign \new_[88766]_  = A232 & A203;
  assign \new_[88769]_  = ~A265 & A233;
  assign \new_[88770]_  = \new_[88769]_  & \new_[88766]_ ;
  assign \new_[88773]_  = ~A299 & ~A266;
  assign \new_[88776]_  = ~A302 & ~A301;
  assign \new_[88777]_  = \new_[88776]_  & \new_[88773]_ ;
  assign \new_[88778]_  = \new_[88777]_  & \new_[88770]_ ;
  assign \new_[88782]_  = A167 & ~A168;
  assign \new_[88783]_  = A169 & \new_[88782]_ ;
  assign \new_[88786]_  = A199 & ~A166;
  assign \new_[88789]_  = A201 & ~A200;
  assign \new_[88790]_  = \new_[88789]_  & \new_[88786]_ ;
  assign \new_[88791]_  = \new_[88790]_  & \new_[88783]_ ;
  assign \new_[88794]_  = ~A233 & A203;
  assign \new_[88797]_  = ~A236 & ~A235;
  assign \new_[88798]_  = \new_[88797]_  & \new_[88794]_ ;
  assign \new_[88801]_  = A266 & A265;
  assign \new_[88804]_  = ~A300 & A298;
  assign \new_[88805]_  = \new_[88804]_  & \new_[88801]_ ;
  assign \new_[88806]_  = \new_[88805]_  & \new_[88798]_ ;
  assign \new_[88810]_  = A167 & ~A168;
  assign \new_[88811]_  = A169 & \new_[88810]_ ;
  assign \new_[88814]_  = A199 & ~A166;
  assign \new_[88817]_  = A201 & ~A200;
  assign \new_[88818]_  = \new_[88817]_  & \new_[88814]_ ;
  assign \new_[88819]_  = \new_[88818]_  & \new_[88811]_ ;
  assign \new_[88822]_  = ~A233 & A203;
  assign \new_[88825]_  = ~A236 & ~A235;
  assign \new_[88826]_  = \new_[88825]_  & \new_[88822]_ ;
  assign \new_[88829]_  = A266 & A265;
  assign \new_[88832]_  = A299 & A298;
  assign \new_[88833]_  = \new_[88832]_  & \new_[88829]_ ;
  assign \new_[88834]_  = \new_[88833]_  & \new_[88826]_ ;
  assign \new_[88838]_  = A167 & ~A168;
  assign \new_[88839]_  = A169 & \new_[88838]_ ;
  assign \new_[88842]_  = A199 & ~A166;
  assign \new_[88845]_  = A201 & ~A200;
  assign \new_[88846]_  = \new_[88845]_  & \new_[88842]_ ;
  assign \new_[88847]_  = \new_[88846]_  & \new_[88839]_ ;
  assign \new_[88850]_  = ~A233 & A203;
  assign \new_[88853]_  = ~A236 & ~A235;
  assign \new_[88854]_  = \new_[88853]_  & \new_[88850]_ ;
  assign \new_[88857]_  = A266 & A265;
  assign \new_[88860]_  = ~A299 & ~A298;
  assign \new_[88861]_  = \new_[88860]_  & \new_[88857]_ ;
  assign \new_[88862]_  = \new_[88861]_  & \new_[88854]_ ;
  assign \new_[88866]_  = A167 & ~A168;
  assign \new_[88867]_  = A169 & \new_[88866]_ ;
  assign \new_[88870]_  = A199 & ~A166;
  assign \new_[88873]_  = A201 & ~A200;
  assign \new_[88874]_  = \new_[88873]_  & \new_[88870]_ ;
  assign \new_[88875]_  = \new_[88874]_  & \new_[88867]_ ;
  assign \new_[88878]_  = ~A233 & A203;
  assign \new_[88881]_  = ~A236 & ~A235;
  assign \new_[88882]_  = \new_[88881]_  & \new_[88878]_ ;
  assign \new_[88885]_  = ~A267 & ~A266;
  assign \new_[88888]_  = ~A300 & A298;
  assign \new_[88889]_  = \new_[88888]_  & \new_[88885]_ ;
  assign \new_[88890]_  = \new_[88889]_  & \new_[88882]_ ;
  assign \new_[88894]_  = A167 & ~A168;
  assign \new_[88895]_  = A169 & \new_[88894]_ ;
  assign \new_[88898]_  = A199 & ~A166;
  assign \new_[88901]_  = A201 & ~A200;
  assign \new_[88902]_  = \new_[88901]_  & \new_[88898]_ ;
  assign \new_[88903]_  = \new_[88902]_  & \new_[88895]_ ;
  assign \new_[88906]_  = ~A233 & A203;
  assign \new_[88909]_  = ~A236 & ~A235;
  assign \new_[88910]_  = \new_[88909]_  & \new_[88906]_ ;
  assign \new_[88913]_  = ~A267 & ~A266;
  assign \new_[88916]_  = A299 & A298;
  assign \new_[88917]_  = \new_[88916]_  & \new_[88913]_ ;
  assign \new_[88918]_  = \new_[88917]_  & \new_[88910]_ ;
  assign \new_[88922]_  = A167 & ~A168;
  assign \new_[88923]_  = A169 & \new_[88922]_ ;
  assign \new_[88926]_  = A199 & ~A166;
  assign \new_[88929]_  = A201 & ~A200;
  assign \new_[88930]_  = \new_[88929]_  & \new_[88926]_ ;
  assign \new_[88931]_  = \new_[88930]_  & \new_[88923]_ ;
  assign \new_[88934]_  = ~A233 & A203;
  assign \new_[88937]_  = ~A236 & ~A235;
  assign \new_[88938]_  = \new_[88937]_  & \new_[88934]_ ;
  assign \new_[88941]_  = ~A267 & ~A266;
  assign \new_[88944]_  = ~A299 & ~A298;
  assign \new_[88945]_  = \new_[88944]_  & \new_[88941]_ ;
  assign \new_[88946]_  = \new_[88945]_  & \new_[88938]_ ;
  assign \new_[88950]_  = A167 & ~A168;
  assign \new_[88951]_  = A169 & \new_[88950]_ ;
  assign \new_[88954]_  = A199 & ~A166;
  assign \new_[88957]_  = A201 & ~A200;
  assign \new_[88958]_  = \new_[88957]_  & \new_[88954]_ ;
  assign \new_[88959]_  = \new_[88958]_  & \new_[88951]_ ;
  assign \new_[88962]_  = ~A233 & A203;
  assign \new_[88965]_  = ~A236 & ~A235;
  assign \new_[88966]_  = \new_[88965]_  & \new_[88962]_ ;
  assign \new_[88969]_  = ~A266 & ~A265;
  assign \new_[88972]_  = ~A300 & A298;
  assign \new_[88973]_  = \new_[88972]_  & \new_[88969]_ ;
  assign \new_[88974]_  = \new_[88973]_  & \new_[88966]_ ;
  assign \new_[88978]_  = A167 & ~A168;
  assign \new_[88979]_  = A169 & \new_[88978]_ ;
  assign \new_[88982]_  = A199 & ~A166;
  assign \new_[88985]_  = A201 & ~A200;
  assign \new_[88986]_  = \new_[88985]_  & \new_[88982]_ ;
  assign \new_[88987]_  = \new_[88986]_  & \new_[88979]_ ;
  assign \new_[88990]_  = ~A233 & A203;
  assign \new_[88993]_  = ~A236 & ~A235;
  assign \new_[88994]_  = \new_[88993]_  & \new_[88990]_ ;
  assign \new_[88997]_  = ~A266 & ~A265;
  assign \new_[89000]_  = A299 & A298;
  assign \new_[89001]_  = \new_[89000]_  & \new_[88997]_ ;
  assign \new_[89002]_  = \new_[89001]_  & \new_[88994]_ ;
  assign \new_[89006]_  = A167 & ~A168;
  assign \new_[89007]_  = A169 & \new_[89006]_ ;
  assign \new_[89010]_  = A199 & ~A166;
  assign \new_[89013]_  = A201 & ~A200;
  assign \new_[89014]_  = \new_[89013]_  & \new_[89010]_ ;
  assign \new_[89015]_  = \new_[89014]_  & \new_[89007]_ ;
  assign \new_[89018]_  = ~A233 & A203;
  assign \new_[89021]_  = ~A236 & ~A235;
  assign \new_[89022]_  = \new_[89021]_  & \new_[89018]_ ;
  assign \new_[89025]_  = ~A266 & ~A265;
  assign \new_[89028]_  = ~A299 & ~A298;
  assign \new_[89029]_  = \new_[89028]_  & \new_[89025]_ ;
  assign \new_[89030]_  = \new_[89029]_  & \new_[89022]_ ;
  assign \new_[89034]_  = A167 & ~A168;
  assign \new_[89035]_  = A169 & \new_[89034]_ ;
  assign \new_[89038]_  = A199 & ~A166;
  assign \new_[89041]_  = A201 & ~A200;
  assign \new_[89042]_  = \new_[89041]_  & \new_[89038]_ ;
  assign \new_[89043]_  = \new_[89042]_  & \new_[89035]_ ;
  assign \new_[89046]_  = ~A233 & A203;
  assign \new_[89049]_  = A265 & ~A234;
  assign \new_[89050]_  = \new_[89049]_  & \new_[89046]_ ;
  assign \new_[89053]_  = A298 & A266;
  assign \new_[89056]_  = ~A302 & ~A301;
  assign \new_[89057]_  = \new_[89056]_  & \new_[89053]_ ;
  assign \new_[89058]_  = \new_[89057]_  & \new_[89050]_ ;
  assign \new_[89062]_  = A167 & ~A168;
  assign \new_[89063]_  = A169 & \new_[89062]_ ;
  assign \new_[89066]_  = A199 & ~A166;
  assign \new_[89069]_  = A201 & ~A200;
  assign \new_[89070]_  = \new_[89069]_  & \new_[89066]_ ;
  assign \new_[89071]_  = \new_[89070]_  & \new_[89063]_ ;
  assign \new_[89074]_  = ~A233 & A203;
  assign \new_[89077]_  = ~A266 & ~A234;
  assign \new_[89078]_  = \new_[89077]_  & \new_[89074]_ ;
  assign \new_[89081]_  = ~A269 & ~A268;
  assign \new_[89084]_  = ~A300 & A298;
  assign \new_[89085]_  = \new_[89084]_  & \new_[89081]_ ;
  assign \new_[89086]_  = \new_[89085]_  & \new_[89078]_ ;
  assign \new_[89090]_  = A167 & ~A168;
  assign \new_[89091]_  = A169 & \new_[89090]_ ;
  assign \new_[89094]_  = A199 & ~A166;
  assign \new_[89097]_  = A201 & ~A200;
  assign \new_[89098]_  = \new_[89097]_  & \new_[89094]_ ;
  assign \new_[89099]_  = \new_[89098]_  & \new_[89091]_ ;
  assign \new_[89102]_  = ~A233 & A203;
  assign \new_[89105]_  = ~A266 & ~A234;
  assign \new_[89106]_  = \new_[89105]_  & \new_[89102]_ ;
  assign \new_[89109]_  = ~A269 & ~A268;
  assign \new_[89112]_  = A299 & A298;
  assign \new_[89113]_  = \new_[89112]_  & \new_[89109]_ ;
  assign \new_[89114]_  = \new_[89113]_  & \new_[89106]_ ;
  assign \new_[89118]_  = A167 & ~A168;
  assign \new_[89119]_  = A169 & \new_[89118]_ ;
  assign \new_[89122]_  = A199 & ~A166;
  assign \new_[89125]_  = A201 & ~A200;
  assign \new_[89126]_  = \new_[89125]_  & \new_[89122]_ ;
  assign \new_[89127]_  = \new_[89126]_  & \new_[89119]_ ;
  assign \new_[89130]_  = ~A233 & A203;
  assign \new_[89133]_  = ~A266 & ~A234;
  assign \new_[89134]_  = \new_[89133]_  & \new_[89130]_ ;
  assign \new_[89137]_  = ~A269 & ~A268;
  assign \new_[89140]_  = ~A299 & ~A298;
  assign \new_[89141]_  = \new_[89140]_  & \new_[89137]_ ;
  assign \new_[89142]_  = \new_[89141]_  & \new_[89134]_ ;
  assign \new_[89146]_  = A167 & ~A168;
  assign \new_[89147]_  = A169 & \new_[89146]_ ;
  assign \new_[89150]_  = A199 & ~A166;
  assign \new_[89153]_  = A201 & ~A200;
  assign \new_[89154]_  = \new_[89153]_  & \new_[89150]_ ;
  assign \new_[89155]_  = \new_[89154]_  & \new_[89147]_ ;
  assign \new_[89158]_  = ~A233 & A203;
  assign \new_[89161]_  = ~A266 & ~A234;
  assign \new_[89162]_  = \new_[89161]_  & \new_[89158]_ ;
  assign \new_[89165]_  = A298 & ~A267;
  assign \new_[89168]_  = ~A302 & ~A301;
  assign \new_[89169]_  = \new_[89168]_  & \new_[89165]_ ;
  assign \new_[89170]_  = \new_[89169]_  & \new_[89162]_ ;
  assign \new_[89174]_  = A167 & ~A168;
  assign \new_[89175]_  = A169 & \new_[89174]_ ;
  assign \new_[89178]_  = A199 & ~A166;
  assign \new_[89181]_  = A201 & ~A200;
  assign \new_[89182]_  = \new_[89181]_  & \new_[89178]_ ;
  assign \new_[89183]_  = \new_[89182]_  & \new_[89175]_ ;
  assign \new_[89186]_  = ~A233 & A203;
  assign \new_[89189]_  = ~A265 & ~A234;
  assign \new_[89190]_  = \new_[89189]_  & \new_[89186]_ ;
  assign \new_[89193]_  = A298 & ~A266;
  assign \new_[89196]_  = ~A302 & ~A301;
  assign \new_[89197]_  = \new_[89196]_  & \new_[89193]_ ;
  assign \new_[89198]_  = \new_[89197]_  & \new_[89190]_ ;
  assign \new_[89202]_  = A167 & ~A168;
  assign \new_[89203]_  = A169 & \new_[89202]_ ;
  assign \new_[89206]_  = A199 & ~A166;
  assign \new_[89209]_  = A201 & ~A200;
  assign \new_[89210]_  = \new_[89209]_  & \new_[89206]_ ;
  assign \new_[89211]_  = \new_[89210]_  & \new_[89203]_ ;
  assign \new_[89214]_  = ~A232 & A203;
  assign \new_[89217]_  = A265 & ~A233;
  assign \new_[89218]_  = \new_[89217]_  & \new_[89214]_ ;
  assign \new_[89221]_  = A298 & A266;
  assign \new_[89224]_  = ~A302 & ~A301;
  assign \new_[89225]_  = \new_[89224]_  & \new_[89221]_ ;
  assign \new_[89226]_  = \new_[89225]_  & \new_[89218]_ ;
  assign \new_[89230]_  = A167 & ~A168;
  assign \new_[89231]_  = A169 & \new_[89230]_ ;
  assign \new_[89234]_  = A199 & ~A166;
  assign \new_[89237]_  = A201 & ~A200;
  assign \new_[89238]_  = \new_[89237]_  & \new_[89234]_ ;
  assign \new_[89239]_  = \new_[89238]_  & \new_[89231]_ ;
  assign \new_[89242]_  = ~A232 & A203;
  assign \new_[89245]_  = ~A266 & ~A233;
  assign \new_[89246]_  = \new_[89245]_  & \new_[89242]_ ;
  assign \new_[89249]_  = ~A269 & ~A268;
  assign \new_[89252]_  = ~A300 & A298;
  assign \new_[89253]_  = \new_[89252]_  & \new_[89249]_ ;
  assign \new_[89254]_  = \new_[89253]_  & \new_[89246]_ ;
  assign \new_[89258]_  = A167 & ~A168;
  assign \new_[89259]_  = A169 & \new_[89258]_ ;
  assign \new_[89262]_  = A199 & ~A166;
  assign \new_[89265]_  = A201 & ~A200;
  assign \new_[89266]_  = \new_[89265]_  & \new_[89262]_ ;
  assign \new_[89267]_  = \new_[89266]_  & \new_[89259]_ ;
  assign \new_[89270]_  = ~A232 & A203;
  assign \new_[89273]_  = ~A266 & ~A233;
  assign \new_[89274]_  = \new_[89273]_  & \new_[89270]_ ;
  assign \new_[89277]_  = ~A269 & ~A268;
  assign \new_[89280]_  = A299 & A298;
  assign \new_[89281]_  = \new_[89280]_  & \new_[89277]_ ;
  assign \new_[89282]_  = \new_[89281]_  & \new_[89274]_ ;
  assign \new_[89286]_  = A167 & ~A168;
  assign \new_[89287]_  = A169 & \new_[89286]_ ;
  assign \new_[89290]_  = A199 & ~A166;
  assign \new_[89293]_  = A201 & ~A200;
  assign \new_[89294]_  = \new_[89293]_  & \new_[89290]_ ;
  assign \new_[89295]_  = \new_[89294]_  & \new_[89287]_ ;
  assign \new_[89298]_  = ~A232 & A203;
  assign \new_[89301]_  = ~A266 & ~A233;
  assign \new_[89302]_  = \new_[89301]_  & \new_[89298]_ ;
  assign \new_[89305]_  = ~A269 & ~A268;
  assign \new_[89308]_  = ~A299 & ~A298;
  assign \new_[89309]_  = \new_[89308]_  & \new_[89305]_ ;
  assign \new_[89310]_  = \new_[89309]_  & \new_[89302]_ ;
  assign \new_[89314]_  = A167 & ~A168;
  assign \new_[89315]_  = A169 & \new_[89314]_ ;
  assign \new_[89318]_  = A199 & ~A166;
  assign \new_[89321]_  = A201 & ~A200;
  assign \new_[89322]_  = \new_[89321]_  & \new_[89318]_ ;
  assign \new_[89323]_  = \new_[89322]_  & \new_[89315]_ ;
  assign \new_[89326]_  = ~A232 & A203;
  assign \new_[89329]_  = ~A266 & ~A233;
  assign \new_[89330]_  = \new_[89329]_  & \new_[89326]_ ;
  assign \new_[89333]_  = A298 & ~A267;
  assign \new_[89336]_  = ~A302 & ~A301;
  assign \new_[89337]_  = \new_[89336]_  & \new_[89333]_ ;
  assign \new_[89338]_  = \new_[89337]_  & \new_[89330]_ ;
  assign \new_[89342]_  = A167 & ~A168;
  assign \new_[89343]_  = A169 & \new_[89342]_ ;
  assign \new_[89346]_  = A199 & ~A166;
  assign \new_[89349]_  = A201 & ~A200;
  assign \new_[89350]_  = \new_[89349]_  & \new_[89346]_ ;
  assign \new_[89351]_  = \new_[89350]_  & \new_[89343]_ ;
  assign \new_[89354]_  = ~A232 & A203;
  assign \new_[89357]_  = ~A265 & ~A233;
  assign \new_[89358]_  = \new_[89357]_  & \new_[89354]_ ;
  assign \new_[89361]_  = A298 & ~A266;
  assign \new_[89364]_  = ~A302 & ~A301;
  assign \new_[89365]_  = \new_[89364]_  & \new_[89361]_ ;
  assign \new_[89366]_  = \new_[89365]_  & \new_[89358]_ ;
  assign \new_[89370]_  = ~A167 & ~A168;
  assign \new_[89371]_  = A169 & \new_[89370]_ ;
  assign \new_[89374]_  = ~A199 & A166;
  assign \new_[89377]_  = ~A233 & A200;
  assign \new_[89378]_  = \new_[89377]_  & \new_[89374]_ ;
  assign \new_[89379]_  = \new_[89378]_  & \new_[89371]_ ;
  assign \new_[89382]_  = ~A236 & ~A235;
  assign \new_[89385]_  = ~A268 & ~A266;
  assign \new_[89386]_  = \new_[89385]_  & \new_[89382]_ ;
  assign \new_[89389]_  = A298 & ~A269;
  assign \new_[89392]_  = ~A302 & ~A301;
  assign \new_[89393]_  = \new_[89392]_  & \new_[89389]_ ;
  assign \new_[89394]_  = \new_[89393]_  & \new_[89386]_ ;
  assign \new_[89398]_  = ~A167 & ~A168;
  assign \new_[89399]_  = A169 & \new_[89398]_ ;
  assign \new_[89402]_  = A199 & A166;
  assign \new_[89405]_  = A201 & ~A200;
  assign \new_[89406]_  = \new_[89405]_  & \new_[89402]_ ;
  assign \new_[89407]_  = \new_[89406]_  & \new_[89399]_ ;
  assign \new_[89410]_  = A232 & A202;
  assign \new_[89413]_  = A265 & A233;
  assign \new_[89414]_  = \new_[89413]_  & \new_[89410]_ ;
  assign \new_[89417]_  = ~A269 & ~A268;
  assign \new_[89420]_  = ~A300 & ~A299;
  assign \new_[89421]_  = \new_[89420]_  & \new_[89417]_ ;
  assign \new_[89422]_  = \new_[89421]_  & \new_[89414]_ ;
  assign \new_[89426]_  = ~A167 & ~A168;
  assign \new_[89427]_  = A169 & \new_[89426]_ ;
  assign \new_[89430]_  = A199 & A166;
  assign \new_[89433]_  = A201 & ~A200;
  assign \new_[89434]_  = \new_[89433]_  & \new_[89430]_ ;
  assign \new_[89435]_  = \new_[89434]_  & \new_[89427]_ ;
  assign \new_[89438]_  = A232 & A202;
  assign \new_[89441]_  = A265 & A233;
  assign \new_[89442]_  = \new_[89441]_  & \new_[89438]_ ;
  assign \new_[89445]_  = ~A269 & ~A268;
  assign \new_[89448]_  = A299 & A298;
  assign \new_[89449]_  = \new_[89448]_  & \new_[89445]_ ;
  assign \new_[89450]_  = \new_[89449]_  & \new_[89442]_ ;
  assign \new_[89454]_  = ~A167 & ~A168;
  assign \new_[89455]_  = A169 & \new_[89454]_ ;
  assign \new_[89458]_  = A199 & A166;
  assign \new_[89461]_  = A201 & ~A200;
  assign \new_[89462]_  = \new_[89461]_  & \new_[89458]_ ;
  assign \new_[89463]_  = \new_[89462]_  & \new_[89455]_ ;
  assign \new_[89466]_  = A232 & A202;
  assign \new_[89469]_  = A265 & A233;
  assign \new_[89470]_  = \new_[89469]_  & \new_[89466]_ ;
  assign \new_[89473]_  = ~A269 & ~A268;
  assign \new_[89476]_  = ~A299 & ~A298;
  assign \new_[89477]_  = \new_[89476]_  & \new_[89473]_ ;
  assign \new_[89478]_  = \new_[89477]_  & \new_[89470]_ ;
  assign \new_[89482]_  = ~A167 & ~A168;
  assign \new_[89483]_  = A169 & \new_[89482]_ ;
  assign \new_[89486]_  = A199 & A166;
  assign \new_[89489]_  = A201 & ~A200;
  assign \new_[89490]_  = \new_[89489]_  & \new_[89486]_ ;
  assign \new_[89491]_  = \new_[89490]_  & \new_[89483]_ ;
  assign \new_[89494]_  = A232 & A202;
  assign \new_[89497]_  = A265 & A233;
  assign \new_[89498]_  = \new_[89497]_  & \new_[89494]_ ;
  assign \new_[89501]_  = ~A299 & ~A267;
  assign \new_[89504]_  = ~A302 & ~A301;
  assign \new_[89505]_  = \new_[89504]_  & \new_[89501]_ ;
  assign \new_[89506]_  = \new_[89505]_  & \new_[89498]_ ;
  assign \new_[89510]_  = ~A167 & ~A168;
  assign \new_[89511]_  = A169 & \new_[89510]_ ;
  assign \new_[89514]_  = A199 & A166;
  assign \new_[89517]_  = A201 & ~A200;
  assign \new_[89518]_  = \new_[89517]_  & \new_[89514]_ ;
  assign \new_[89519]_  = \new_[89518]_  & \new_[89511]_ ;
  assign \new_[89522]_  = A232 & A202;
  assign \new_[89525]_  = A265 & A233;
  assign \new_[89526]_  = \new_[89525]_  & \new_[89522]_ ;
  assign \new_[89529]_  = ~A299 & A266;
  assign \new_[89532]_  = ~A302 & ~A301;
  assign \new_[89533]_  = \new_[89532]_  & \new_[89529]_ ;
  assign \new_[89534]_  = \new_[89533]_  & \new_[89526]_ ;
  assign \new_[89538]_  = ~A167 & ~A168;
  assign \new_[89539]_  = A169 & \new_[89538]_ ;
  assign \new_[89542]_  = A199 & A166;
  assign \new_[89545]_  = A201 & ~A200;
  assign \new_[89546]_  = \new_[89545]_  & \new_[89542]_ ;
  assign \new_[89547]_  = \new_[89546]_  & \new_[89539]_ ;
  assign \new_[89550]_  = A232 & A202;
  assign \new_[89553]_  = ~A265 & A233;
  assign \new_[89554]_  = \new_[89553]_  & \new_[89550]_ ;
  assign \new_[89557]_  = ~A299 & ~A266;
  assign \new_[89560]_  = ~A302 & ~A301;
  assign \new_[89561]_  = \new_[89560]_  & \new_[89557]_ ;
  assign \new_[89562]_  = \new_[89561]_  & \new_[89554]_ ;
  assign \new_[89566]_  = ~A167 & ~A168;
  assign \new_[89567]_  = A169 & \new_[89566]_ ;
  assign \new_[89570]_  = A199 & A166;
  assign \new_[89573]_  = A201 & ~A200;
  assign \new_[89574]_  = \new_[89573]_  & \new_[89570]_ ;
  assign \new_[89575]_  = \new_[89574]_  & \new_[89567]_ ;
  assign \new_[89578]_  = ~A233 & A202;
  assign \new_[89581]_  = ~A236 & ~A235;
  assign \new_[89582]_  = \new_[89581]_  & \new_[89578]_ ;
  assign \new_[89585]_  = A266 & A265;
  assign \new_[89588]_  = ~A300 & A298;
  assign \new_[89589]_  = \new_[89588]_  & \new_[89585]_ ;
  assign \new_[89590]_  = \new_[89589]_  & \new_[89582]_ ;
  assign \new_[89594]_  = ~A167 & ~A168;
  assign \new_[89595]_  = A169 & \new_[89594]_ ;
  assign \new_[89598]_  = A199 & A166;
  assign \new_[89601]_  = A201 & ~A200;
  assign \new_[89602]_  = \new_[89601]_  & \new_[89598]_ ;
  assign \new_[89603]_  = \new_[89602]_  & \new_[89595]_ ;
  assign \new_[89606]_  = ~A233 & A202;
  assign \new_[89609]_  = ~A236 & ~A235;
  assign \new_[89610]_  = \new_[89609]_  & \new_[89606]_ ;
  assign \new_[89613]_  = A266 & A265;
  assign \new_[89616]_  = A299 & A298;
  assign \new_[89617]_  = \new_[89616]_  & \new_[89613]_ ;
  assign \new_[89618]_  = \new_[89617]_  & \new_[89610]_ ;
  assign \new_[89622]_  = ~A167 & ~A168;
  assign \new_[89623]_  = A169 & \new_[89622]_ ;
  assign \new_[89626]_  = A199 & A166;
  assign \new_[89629]_  = A201 & ~A200;
  assign \new_[89630]_  = \new_[89629]_  & \new_[89626]_ ;
  assign \new_[89631]_  = \new_[89630]_  & \new_[89623]_ ;
  assign \new_[89634]_  = ~A233 & A202;
  assign \new_[89637]_  = ~A236 & ~A235;
  assign \new_[89638]_  = \new_[89637]_  & \new_[89634]_ ;
  assign \new_[89641]_  = A266 & A265;
  assign \new_[89644]_  = ~A299 & ~A298;
  assign \new_[89645]_  = \new_[89644]_  & \new_[89641]_ ;
  assign \new_[89646]_  = \new_[89645]_  & \new_[89638]_ ;
  assign \new_[89650]_  = ~A167 & ~A168;
  assign \new_[89651]_  = A169 & \new_[89650]_ ;
  assign \new_[89654]_  = A199 & A166;
  assign \new_[89657]_  = A201 & ~A200;
  assign \new_[89658]_  = \new_[89657]_  & \new_[89654]_ ;
  assign \new_[89659]_  = \new_[89658]_  & \new_[89651]_ ;
  assign \new_[89662]_  = ~A233 & A202;
  assign \new_[89665]_  = ~A236 & ~A235;
  assign \new_[89666]_  = \new_[89665]_  & \new_[89662]_ ;
  assign \new_[89669]_  = ~A267 & ~A266;
  assign \new_[89672]_  = ~A300 & A298;
  assign \new_[89673]_  = \new_[89672]_  & \new_[89669]_ ;
  assign \new_[89674]_  = \new_[89673]_  & \new_[89666]_ ;
  assign \new_[89678]_  = ~A167 & ~A168;
  assign \new_[89679]_  = A169 & \new_[89678]_ ;
  assign \new_[89682]_  = A199 & A166;
  assign \new_[89685]_  = A201 & ~A200;
  assign \new_[89686]_  = \new_[89685]_  & \new_[89682]_ ;
  assign \new_[89687]_  = \new_[89686]_  & \new_[89679]_ ;
  assign \new_[89690]_  = ~A233 & A202;
  assign \new_[89693]_  = ~A236 & ~A235;
  assign \new_[89694]_  = \new_[89693]_  & \new_[89690]_ ;
  assign \new_[89697]_  = ~A267 & ~A266;
  assign \new_[89700]_  = A299 & A298;
  assign \new_[89701]_  = \new_[89700]_  & \new_[89697]_ ;
  assign \new_[89702]_  = \new_[89701]_  & \new_[89694]_ ;
  assign \new_[89706]_  = ~A167 & ~A168;
  assign \new_[89707]_  = A169 & \new_[89706]_ ;
  assign \new_[89710]_  = A199 & A166;
  assign \new_[89713]_  = A201 & ~A200;
  assign \new_[89714]_  = \new_[89713]_  & \new_[89710]_ ;
  assign \new_[89715]_  = \new_[89714]_  & \new_[89707]_ ;
  assign \new_[89718]_  = ~A233 & A202;
  assign \new_[89721]_  = ~A236 & ~A235;
  assign \new_[89722]_  = \new_[89721]_  & \new_[89718]_ ;
  assign \new_[89725]_  = ~A267 & ~A266;
  assign \new_[89728]_  = ~A299 & ~A298;
  assign \new_[89729]_  = \new_[89728]_  & \new_[89725]_ ;
  assign \new_[89730]_  = \new_[89729]_  & \new_[89722]_ ;
  assign \new_[89734]_  = ~A167 & ~A168;
  assign \new_[89735]_  = A169 & \new_[89734]_ ;
  assign \new_[89738]_  = A199 & A166;
  assign \new_[89741]_  = A201 & ~A200;
  assign \new_[89742]_  = \new_[89741]_  & \new_[89738]_ ;
  assign \new_[89743]_  = \new_[89742]_  & \new_[89735]_ ;
  assign \new_[89746]_  = ~A233 & A202;
  assign \new_[89749]_  = ~A236 & ~A235;
  assign \new_[89750]_  = \new_[89749]_  & \new_[89746]_ ;
  assign \new_[89753]_  = ~A266 & ~A265;
  assign \new_[89756]_  = ~A300 & A298;
  assign \new_[89757]_  = \new_[89756]_  & \new_[89753]_ ;
  assign \new_[89758]_  = \new_[89757]_  & \new_[89750]_ ;
  assign \new_[89762]_  = ~A167 & ~A168;
  assign \new_[89763]_  = A169 & \new_[89762]_ ;
  assign \new_[89766]_  = A199 & A166;
  assign \new_[89769]_  = A201 & ~A200;
  assign \new_[89770]_  = \new_[89769]_  & \new_[89766]_ ;
  assign \new_[89771]_  = \new_[89770]_  & \new_[89763]_ ;
  assign \new_[89774]_  = ~A233 & A202;
  assign \new_[89777]_  = ~A236 & ~A235;
  assign \new_[89778]_  = \new_[89777]_  & \new_[89774]_ ;
  assign \new_[89781]_  = ~A266 & ~A265;
  assign \new_[89784]_  = A299 & A298;
  assign \new_[89785]_  = \new_[89784]_  & \new_[89781]_ ;
  assign \new_[89786]_  = \new_[89785]_  & \new_[89778]_ ;
  assign \new_[89790]_  = ~A167 & ~A168;
  assign \new_[89791]_  = A169 & \new_[89790]_ ;
  assign \new_[89794]_  = A199 & A166;
  assign \new_[89797]_  = A201 & ~A200;
  assign \new_[89798]_  = \new_[89797]_  & \new_[89794]_ ;
  assign \new_[89799]_  = \new_[89798]_  & \new_[89791]_ ;
  assign \new_[89802]_  = ~A233 & A202;
  assign \new_[89805]_  = ~A236 & ~A235;
  assign \new_[89806]_  = \new_[89805]_  & \new_[89802]_ ;
  assign \new_[89809]_  = ~A266 & ~A265;
  assign \new_[89812]_  = ~A299 & ~A298;
  assign \new_[89813]_  = \new_[89812]_  & \new_[89809]_ ;
  assign \new_[89814]_  = \new_[89813]_  & \new_[89806]_ ;
  assign \new_[89818]_  = ~A167 & ~A168;
  assign \new_[89819]_  = A169 & \new_[89818]_ ;
  assign \new_[89822]_  = A199 & A166;
  assign \new_[89825]_  = A201 & ~A200;
  assign \new_[89826]_  = \new_[89825]_  & \new_[89822]_ ;
  assign \new_[89827]_  = \new_[89826]_  & \new_[89819]_ ;
  assign \new_[89830]_  = ~A233 & A202;
  assign \new_[89833]_  = A265 & ~A234;
  assign \new_[89834]_  = \new_[89833]_  & \new_[89830]_ ;
  assign \new_[89837]_  = A298 & A266;
  assign \new_[89840]_  = ~A302 & ~A301;
  assign \new_[89841]_  = \new_[89840]_  & \new_[89837]_ ;
  assign \new_[89842]_  = \new_[89841]_  & \new_[89834]_ ;
  assign \new_[89846]_  = ~A167 & ~A168;
  assign \new_[89847]_  = A169 & \new_[89846]_ ;
  assign \new_[89850]_  = A199 & A166;
  assign \new_[89853]_  = A201 & ~A200;
  assign \new_[89854]_  = \new_[89853]_  & \new_[89850]_ ;
  assign \new_[89855]_  = \new_[89854]_  & \new_[89847]_ ;
  assign \new_[89858]_  = ~A233 & A202;
  assign \new_[89861]_  = ~A266 & ~A234;
  assign \new_[89862]_  = \new_[89861]_  & \new_[89858]_ ;
  assign \new_[89865]_  = ~A269 & ~A268;
  assign \new_[89868]_  = ~A300 & A298;
  assign \new_[89869]_  = \new_[89868]_  & \new_[89865]_ ;
  assign \new_[89870]_  = \new_[89869]_  & \new_[89862]_ ;
  assign \new_[89874]_  = ~A167 & ~A168;
  assign \new_[89875]_  = A169 & \new_[89874]_ ;
  assign \new_[89878]_  = A199 & A166;
  assign \new_[89881]_  = A201 & ~A200;
  assign \new_[89882]_  = \new_[89881]_  & \new_[89878]_ ;
  assign \new_[89883]_  = \new_[89882]_  & \new_[89875]_ ;
  assign \new_[89886]_  = ~A233 & A202;
  assign \new_[89889]_  = ~A266 & ~A234;
  assign \new_[89890]_  = \new_[89889]_  & \new_[89886]_ ;
  assign \new_[89893]_  = ~A269 & ~A268;
  assign \new_[89896]_  = A299 & A298;
  assign \new_[89897]_  = \new_[89896]_  & \new_[89893]_ ;
  assign \new_[89898]_  = \new_[89897]_  & \new_[89890]_ ;
  assign \new_[89902]_  = ~A167 & ~A168;
  assign \new_[89903]_  = A169 & \new_[89902]_ ;
  assign \new_[89906]_  = A199 & A166;
  assign \new_[89909]_  = A201 & ~A200;
  assign \new_[89910]_  = \new_[89909]_  & \new_[89906]_ ;
  assign \new_[89911]_  = \new_[89910]_  & \new_[89903]_ ;
  assign \new_[89914]_  = ~A233 & A202;
  assign \new_[89917]_  = ~A266 & ~A234;
  assign \new_[89918]_  = \new_[89917]_  & \new_[89914]_ ;
  assign \new_[89921]_  = ~A269 & ~A268;
  assign \new_[89924]_  = ~A299 & ~A298;
  assign \new_[89925]_  = \new_[89924]_  & \new_[89921]_ ;
  assign \new_[89926]_  = \new_[89925]_  & \new_[89918]_ ;
  assign \new_[89930]_  = ~A167 & ~A168;
  assign \new_[89931]_  = A169 & \new_[89930]_ ;
  assign \new_[89934]_  = A199 & A166;
  assign \new_[89937]_  = A201 & ~A200;
  assign \new_[89938]_  = \new_[89937]_  & \new_[89934]_ ;
  assign \new_[89939]_  = \new_[89938]_  & \new_[89931]_ ;
  assign \new_[89942]_  = ~A233 & A202;
  assign \new_[89945]_  = ~A266 & ~A234;
  assign \new_[89946]_  = \new_[89945]_  & \new_[89942]_ ;
  assign \new_[89949]_  = A298 & ~A267;
  assign \new_[89952]_  = ~A302 & ~A301;
  assign \new_[89953]_  = \new_[89952]_  & \new_[89949]_ ;
  assign \new_[89954]_  = \new_[89953]_  & \new_[89946]_ ;
  assign \new_[89958]_  = ~A167 & ~A168;
  assign \new_[89959]_  = A169 & \new_[89958]_ ;
  assign \new_[89962]_  = A199 & A166;
  assign \new_[89965]_  = A201 & ~A200;
  assign \new_[89966]_  = \new_[89965]_  & \new_[89962]_ ;
  assign \new_[89967]_  = \new_[89966]_  & \new_[89959]_ ;
  assign \new_[89970]_  = ~A233 & A202;
  assign \new_[89973]_  = ~A265 & ~A234;
  assign \new_[89974]_  = \new_[89973]_  & \new_[89970]_ ;
  assign \new_[89977]_  = A298 & ~A266;
  assign \new_[89980]_  = ~A302 & ~A301;
  assign \new_[89981]_  = \new_[89980]_  & \new_[89977]_ ;
  assign \new_[89982]_  = \new_[89981]_  & \new_[89974]_ ;
  assign \new_[89986]_  = ~A167 & ~A168;
  assign \new_[89987]_  = A169 & \new_[89986]_ ;
  assign \new_[89990]_  = A199 & A166;
  assign \new_[89993]_  = A201 & ~A200;
  assign \new_[89994]_  = \new_[89993]_  & \new_[89990]_ ;
  assign \new_[89995]_  = \new_[89994]_  & \new_[89987]_ ;
  assign \new_[89998]_  = ~A232 & A202;
  assign \new_[90001]_  = A265 & ~A233;
  assign \new_[90002]_  = \new_[90001]_  & \new_[89998]_ ;
  assign \new_[90005]_  = A298 & A266;
  assign \new_[90008]_  = ~A302 & ~A301;
  assign \new_[90009]_  = \new_[90008]_  & \new_[90005]_ ;
  assign \new_[90010]_  = \new_[90009]_  & \new_[90002]_ ;
  assign \new_[90014]_  = ~A167 & ~A168;
  assign \new_[90015]_  = A169 & \new_[90014]_ ;
  assign \new_[90018]_  = A199 & A166;
  assign \new_[90021]_  = A201 & ~A200;
  assign \new_[90022]_  = \new_[90021]_  & \new_[90018]_ ;
  assign \new_[90023]_  = \new_[90022]_  & \new_[90015]_ ;
  assign \new_[90026]_  = ~A232 & A202;
  assign \new_[90029]_  = ~A266 & ~A233;
  assign \new_[90030]_  = \new_[90029]_  & \new_[90026]_ ;
  assign \new_[90033]_  = ~A269 & ~A268;
  assign \new_[90036]_  = ~A300 & A298;
  assign \new_[90037]_  = \new_[90036]_  & \new_[90033]_ ;
  assign \new_[90038]_  = \new_[90037]_  & \new_[90030]_ ;
  assign \new_[90042]_  = ~A167 & ~A168;
  assign \new_[90043]_  = A169 & \new_[90042]_ ;
  assign \new_[90046]_  = A199 & A166;
  assign \new_[90049]_  = A201 & ~A200;
  assign \new_[90050]_  = \new_[90049]_  & \new_[90046]_ ;
  assign \new_[90051]_  = \new_[90050]_  & \new_[90043]_ ;
  assign \new_[90054]_  = ~A232 & A202;
  assign \new_[90057]_  = ~A266 & ~A233;
  assign \new_[90058]_  = \new_[90057]_  & \new_[90054]_ ;
  assign \new_[90061]_  = ~A269 & ~A268;
  assign \new_[90064]_  = A299 & A298;
  assign \new_[90065]_  = \new_[90064]_  & \new_[90061]_ ;
  assign \new_[90066]_  = \new_[90065]_  & \new_[90058]_ ;
  assign \new_[90070]_  = ~A167 & ~A168;
  assign \new_[90071]_  = A169 & \new_[90070]_ ;
  assign \new_[90074]_  = A199 & A166;
  assign \new_[90077]_  = A201 & ~A200;
  assign \new_[90078]_  = \new_[90077]_  & \new_[90074]_ ;
  assign \new_[90079]_  = \new_[90078]_  & \new_[90071]_ ;
  assign \new_[90082]_  = ~A232 & A202;
  assign \new_[90085]_  = ~A266 & ~A233;
  assign \new_[90086]_  = \new_[90085]_  & \new_[90082]_ ;
  assign \new_[90089]_  = ~A269 & ~A268;
  assign \new_[90092]_  = ~A299 & ~A298;
  assign \new_[90093]_  = \new_[90092]_  & \new_[90089]_ ;
  assign \new_[90094]_  = \new_[90093]_  & \new_[90086]_ ;
  assign \new_[90098]_  = ~A167 & ~A168;
  assign \new_[90099]_  = A169 & \new_[90098]_ ;
  assign \new_[90102]_  = A199 & A166;
  assign \new_[90105]_  = A201 & ~A200;
  assign \new_[90106]_  = \new_[90105]_  & \new_[90102]_ ;
  assign \new_[90107]_  = \new_[90106]_  & \new_[90099]_ ;
  assign \new_[90110]_  = ~A232 & A202;
  assign \new_[90113]_  = ~A266 & ~A233;
  assign \new_[90114]_  = \new_[90113]_  & \new_[90110]_ ;
  assign \new_[90117]_  = A298 & ~A267;
  assign \new_[90120]_  = ~A302 & ~A301;
  assign \new_[90121]_  = \new_[90120]_  & \new_[90117]_ ;
  assign \new_[90122]_  = \new_[90121]_  & \new_[90114]_ ;
  assign \new_[90126]_  = ~A167 & ~A168;
  assign \new_[90127]_  = A169 & \new_[90126]_ ;
  assign \new_[90130]_  = A199 & A166;
  assign \new_[90133]_  = A201 & ~A200;
  assign \new_[90134]_  = \new_[90133]_  & \new_[90130]_ ;
  assign \new_[90135]_  = \new_[90134]_  & \new_[90127]_ ;
  assign \new_[90138]_  = ~A232 & A202;
  assign \new_[90141]_  = ~A265 & ~A233;
  assign \new_[90142]_  = \new_[90141]_  & \new_[90138]_ ;
  assign \new_[90145]_  = A298 & ~A266;
  assign \new_[90148]_  = ~A302 & ~A301;
  assign \new_[90149]_  = \new_[90148]_  & \new_[90145]_ ;
  assign \new_[90150]_  = \new_[90149]_  & \new_[90142]_ ;
  assign \new_[90154]_  = ~A167 & ~A168;
  assign \new_[90155]_  = A169 & \new_[90154]_ ;
  assign \new_[90158]_  = A199 & A166;
  assign \new_[90161]_  = A201 & ~A200;
  assign \new_[90162]_  = \new_[90161]_  & \new_[90158]_ ;
  assign \new_[90163]_  = \new_[90162]_  & \new_[90155]_ ;
  assign \new_[90166]_  = A232 & A203;
  assign \new_[90169]_  = A265 & A233;
  assign \new_[90170]_  = \new_[90169]_  & \new_[90166]_ ;
  assign \new_[90173]_  = ~A269 & ~A268;
  assign \new_[90176]_  = ~A300 & ~A299;
  assign \new_[90177]_  = \new_[90176]_  & \new_[90173]_ ;
  assign \new_[90178]_  = \new_[90177]_  & \new_[90170]_ ;
  assign \new_[90182]_  = ~A167 & ~A168;
  assign \new_[90183]_  = A169 & \new_[90182]_ ;
  assign \new_[90186]_  = A199 & A166;
  assign \new_[90189]_  = A201 & ~A200;
  assign \new_[90190]_  = \new_[90189]_  & \new_[90186]_ ;
  assign \new_[90191]_  = \new_[90190]_  & \new_[90183]_ ;
  assign \new_[90194]_  = A232 & A203;
  assign \new_[90197]_  = A265 & A233;
  assign \new_[90198]_  = \new_[90197]_  & \new_[90194]_ ;
  assign \new_[90201]_  = ~A269 & ~A268;
  assign \new_[90204]_  = A299 & A298;
  assign \new_[90205]_  = \new_[90204]_  & \new_[90201]_ ;
  assign \new_[90206]_  = \new_[90205]_  & \new_[90198]_ ;
  assign \new_[90210]_  = ~A167 & ~A168;
  assign \new_[90211]_  = A169 & \new_[90210]_ ;
  assign \new_[90214]_  = A199 & A166;
  assign \new_[90217]_  = A201 & ~A200;
  assign \new_[90218]_  = \new_[90217]_  & \new_[90214]_ ;
  assign \new_[90219]_  = \new_[90218]_  & \new_[90211]_ ;
  assign \new_[90222]_  = A232 & A203;
  assign \new_[90225]_  = A265 & A233;
  assign \new_[90226]_  = \new_[90225]_  & \new_[90222]_ ;
  assign \new_[90229]_  = ~A269 & ~A268;
  assign \new_[90232]_  = ~A299 & ~A298;
  assign \new_[90233]_  = \new_[90232]_  & \new_[90229]_ ;
  assign \new_[90234]_  = \new_[90233]_  & \new_[90226]_ ;
  assign \new_[90238]_  = ~A167 & ~A168;
  assign \new_[90239]_  = A169 & \new_[90238]_ ;
  assign \new_[90242]_  = A199 & A166;
  assign \new_[90245]_  = A201 & ~A200;
  assign \new_[90246]_  = \new_[90245]_  & \new_[90242]_ ;
  assign \new_[90247]_  = \new_[90246]_  & \new_[90239]_ ;
  assign \new_[90250]_  = A232 & A203;
  assign \new_[90253]_  = A265 & A233;
  assign \new_[90254]_  = \new_[90253]_  & \new_[90250]_ ;
  assign \new_[90257]_  = ~A299 & ~A267;
  assign \new_[90260]_  = ~A302 & ~A301;
  assign \new_[90261]_  = \new_[90260]_  & \new_[90257]_ ;
  assign \new_[90262]_  = \new_[90261]_  & \new_[90254]_ ;
  assign \new_[90266]_  = ~A167 & ~A168;
  assign \new_[90267]_  = A169 & \new_[90266]_ ;
  assign \new_[90270]_  = A199 & A166;
  assign \new_[90273]_  = A201 & ~A200;
  assign \new_[90274]_  = \new_[90273]_  & \new_[90270]_ ;
  assign \new_[90275]_  = \new_[90274]_  & \new_[90267]_ ;
  assign \new_[90278]_  = A232 & A203;
  assign \new_[90281]_  = A265 & A233;
  assign \new_[90282]_  = \new_[90281]_  & \new_[90278]_ ;
  assign \new_[90285]_  = ~A299 & A266;
  assign \new_[90288]_  = ~A302 & ~A301;
  assign \new_[90289]_  = \new_[90288]_  & \new_[90285]_ ;
  assign \new_[90290]_  = \new_[90289]_  & \new_[90282]_ ;
  assign \new_[90294]_  = ~A167 & ~A168;
  assign \new_[90295]_  = A169 & \new_[90294]_ ;
  assign \new_[90298]_  = A199 & A166;
  assign \new_[90301]_  = A201 & ~A200;
  assign \new_[90302]_  = \new_[90301]_  & \new_[90298]_ ;
  assign \new_[90303]_  = \new_[90302]_  & \new_[90295]_ ;
  assign \new_[90306]_  = A232 & A203;
  assign \new_[90309]_  = ~A265 & A233;
  assign \new_[90310]_  = \new_[90309]_  & \new_[90306]_ ;
  assign \new_[90313]_  = ~A299 & ~A266;
  assign \new_[90316]_  = ~A302 & ~A301;
  assign \new_[90317]_  = \new_[90316]_  & \new_[90313]_ ;
  assign \new_[90318]_  = \new_[90317]_  & \new_[90310]_ ;
  assign \new_[90322]_  = ~A167 & ~A168;
  assign \new_[90323]_  = A169 & \new_[90322]_ ;
  assign \new_[90326]_  = A199 & A166;
  assign \new_[90329]_  = A201 & ~A200;
  assign \new_[90330]_  = \new_[90329]_  & \new_[90326]_ ;
  assign \new_[90331]_  = \new_[90330]_  & \new_[90323]_ ;
  assign \new_[90334]_  = ~A233 & A203;
  assign \new_[90337]_  = ~A236 & ~A235;
  assign \new_[90338]_  = \new_[90337]_  & \new_[90334]_ ;
  assign \new_[90341]_  = A266 & A265;
  assign \new_[90344]_  = ~A300 & A298;
  assign \new_[90345]_  = \new_[90344]_  & \new_[90341]_ ;
  assign \new_[90346]_  = \new_[90345]_  & \new_[90338]_ ;
  assign \new_[90350]_  = ~A167 & ~A168;
  assign \new_[90351]_  = A169 & \new_[90350]_ ;
  assign \new_[90354]_  = A199 & A166;
  assign \new_[90357]_  = A201 & ~A200;
  assign \new_[90358]_  = \new_[90357]_  & \new_[90354]_ ;
  assign \new_[90359]_  = \new_[90358]_  & \new_[90351]_ ;
  assign \new_[90362]_  = ~A233 & A203;
  assign \new_[90365]_  = ~A236 & ~A235;
  assign \new_[90366]_  = \new_[90365]_  & \new_[90362]_ ;
  assign \new_[90369]_  = A266 & A265;
  assign \new_[90372]_  = A299 & A298;
  assign \new_[90373]_  = \new_[90372]_  & \new_[90369]_ ;
  assign \new_[90374]_  = \new_[90373]_  & \new_[90366]_ ;
  assign \new_[90378]_  = ~A167 & ~A168;
  assign \new_[90379]_  = A169 & \new_[90378]_ ;
  assign \new_[90382]_  = A199 & A166;
  assign \new_[90385]_  = A201 & ~A200;
  assign \new_[90386]_  = \new_[90385]_  & \new_[90382]_ ;
  assign \new_[90387]_  = \new_[90386]_  & \new_[90379]_ ;
  assign \new_[90390]_  = ~A233 & A203;
  assign \new_[90393]_  = ~A236 & ~A235;
  assign \new_[90394]_  = \new_[90393]_  & \new_[90390]_ ;
  assign \new_[90397]_  = A266 & A265;
  assign \new_[90400]_  = ~A299 & ~A298;
  assign \new_[90401]_  = \new_[90400]_  & \new_[90397]_ ;
  assign \new_[90402]_  = \new_[90401]_  & \new_[90394]_ ;
  assign \new_[90406]_  = ~A167 & ~A168;
  assign \new_[90407]_  = A169 & \new_[90406]_ ;
  assign \new_[90410]_  = A199 & A166;
  assign \new_[90413]_  = A201 & ~A200;
  assign \new_[90414]_  = \new_[90413]_  & \new_[90410]_ ;
  assign \new_[90415]_  = \new_[90414]_  & \new_[90407]_ ;
  assign \new_[90418]_  = ~A233 & A203;
  assign \new_[90421]_  = ~A236 & ~A235;
  assign \new_[90422]_  = \new_[90421]_  & \new_[90418]_ ;
  assign \new_[90425]_  = ~A267 & ~A266;
  assign \new_[90428]_  = ~A300 & A298;
  assign \new_[90429]_  = \new_[90428]_  & \new_[90425]_ ;
  assign \new_[90430]_  = \new_[90429]_  & \new_[90422]_ ;
  assign \new_[90434]_  = ~A167 & ~A168;
  assign \new_[90435]_  = A169 & \new_[90434]_ ;
  assign \new_[90438]_  = A199 & A166;
  assign \new_[90441]_  = A201 & ~A200;
  assign \new_[90442]_  = \new_[90441]_  & \new_[90438]_ ;
  assign \new_[90443]_  = \new_[90442]_  & \new_[90435]_ ;
  assign \new_[90446]_  = ~A233 & A203;
  assign \new_[90449]_  = ~A236 & ~A235;
  assign \new_[90450]_  = \new_[90449]_  & \new_[90446]_ ;
  assign \new_[90453]_  = ~A267 & ~A266;
  assign \new_[90456]_  = A299 & A298;
  assign \new_[90457]_  = \new_[90456]_  & \new_[90453]_ ;
  assign \new_[90458]_  = \new_[90457]_  & \new_[90450]_ ;
  assign \new_[90462]_  = ~A167 & ~A168;
  assign \new_[90463]_  = A169 & \new_[90462]_ ;
  assign \new_[90466]_  = A199 & A166;
  assign \new_[90469]_  = A201 & ~A200;
  assign \new_[90470]_  = \new_[90469]_  & \new_[90466]_ ;
  assign \new_[90471]_  = \new_[90470]_  & \new_[90463]_ ;
  assign \new_[90474]_  = ~A233 & A203;
  assign \new_[90477]_  = ~A236 & ~A235;
  assign \new_[90478]_  = \new_[90477]_  & \new_[90474]_ ;
  assign \new_[90481]_  = ~A267 & ~A266;
  assign \new_[90484]_  = ~A299 & ~A298;
  assign \new_[90485]_  = \new_[90484]_  & \new_[90481]_ ;
  assign \new_[90486]_  = \new_[90485]_  & \new_[90478]_ ;
  assign \new_[90490]_  = ~A167 & ~A168;
  assign \new_[90491]_  = A169 & \new_[90490]_ ;
  assign \new_[90494]_  = A199 & A166;
  assign \new_[90497]_  = A201 & ~A200;
  assign \new_[90498]_  = \new_[90497]_  & \new_[90494]_ ;
  assign \new_[90499]_  = \new_[90498]_  & \new_[90491]_ ;
  assign \new_[90502]_  = ~A233 & A203;
  assign \new_[90505]_  = ~A236 & ~A235;
  assign \new_[90506]_  = \new_[90505]_  & \new_[90502]_ ;
  assign \new_[90509]_  = ~A266 & ~A265;
  assign \new_[90512]_  = ~A300 & A298;
  assign \new_[90513]_  = \new_[90512]_  & \new_[90509]_ ;
  assign \new_[90514]_  = \new_[90513]_  & \new_[90506]_ ;
  assign \new_[90518]_  = ~A167 & ~A168;
  assign \new_[90519]_  = A169 & \new_[90518]_ ;
  assign \new_[90522]_  = A199 & A166;
  assign \new_[90525]_  = A201 & ~A200;
  assign \new_[90526]_  = \new_[90525]_  & \new_[90522]_ ;
  assign \new_[90527]_  = \new_[90526]_  & \new_[90519]_ ;
  assign \new_[90530]_  = ~A233 & A203;
  assign \new_[90533]_  = ~A236 & ~A235;
  assign \new_[90534]_  = \new_[90533]_  & \new_[90530]_ ;
  assign \new_[90537]_  = ~A266 & ~A265;
  assign \new_[90540]_  = A299 & A298;
  assign \new_[90541]_  = \new_[90540]_  & \new_[90537]_ ;
  assign \new_[90542]_  = \new_[90541]_  & \new_[90534]_ ;
  assign \new_[90546]_  = ~A167 & ~A168;
  assign \new_[90547]_  = A169 & \new_[90546]_ ;
  assign \new_[90550]_  = A199 & A166;
  assign \new_[90553]_  = A201 & ~A200;
  assign \new_[90554]_  = \new_[90553]_  & \new_[90550]_ ;
  assign \new_[90555]_  = \new_[90554]_  & \new_[90547]_ ;
  assign \new_[90558]_  = ~A233 & A203;
  assign \new_[90561]_  = ~A236 & ~A235;
  assign \new_[90562]_  = \new_[90561]_  & \new_[90558]_ ;
  assign \new_[90565]_  = ~A266 & ~A265;
  assign \new_[90568]_  = ~A299 & ~A298;
  assign \new_[90569]_  = \new_[90568]_  & \new_[90565]_ ;
  assign \new_[90570]_  = \new_[90569]_  & \new_[90562]_ ;
  assign \new_[90574]_  = ~A167 & ~A168;
  assign \new_[90575]_  = A169 & \new_[90574]_ ;
  assign \new_[90578]_  = A199 & A166;
  assign \new_[90581]_  = A201 & ~A200;
  assign \new_[90582]_  = \new_[90581]_  & \new_[90578]_ ;
  assign \new_[90583]_  = \new_[90582]_  & \new_[90575]_ ;
  assign \new_[90586]_  = ~A233 & A203;
  assign \new_[90589]_  = A265 & ~A234;
  assign \new_[90590]_  = \new_[90589]_  & \new_[90586]_ ;
  assign \new_[90593]_  = A298 & A266;
  assign \new_[90596]_  = ~A302 & ~A301;
  assign \new_[90597]_  = \new_[90596]_  & \new_[90593]_ ;
  assign \new_[90598]_  = \new_[90597]_  & \new_[90590]_ ;
  assign \new_[90602]_  = ~A167 & ~A168;
  assign \new_[90603]_  = A169 & \new_[90602]_ ;
  assign \new_[90606]_  = A199 & A166;
  assign \new_[90609]_  = A201 & ~A200;
  assign \new_[90610]_  = \new_[90609]_  & \new_[90606]_ ;
  assign \new_[90611]_  = \new_[90610]_  & \new_[90603]_ ;
  assign \new_[90614]_  = ~A233 & A203;
  assign \new_[90617]_  = ~A266 & ~A234;
  assign \new_[90618]_  = \new_[90617]_  & \new_[90614]_ ;
  assign \new_[90621]_  = ~A269 & ~A268;
  assign \new_[90624]_  = ~A300 & A298;
  assign \new_[90625]_  = \new_[90624]_  & \new_[90621]_ ;
  assign \new_[90626]_  = \new_[90625]_  & \new_[90618]_ ;
  assign \new_[90630]_  = ~A167 & ~A168;
  assign \new_[90631]_  = A169 & \new_[90630]_ ;
  assign \new_[90634]_  = A199 & A166;
  assign \new_[90637]_  = A201 & ~A200;
  assign \new_[90638]_  = \new_[90637]_  & \new_[90634]_ ;
  assign \new_[90639]_  = \new_[90638]_  & \new_[90631]_ ;
  assign \new_[90642]_  = ~A233 & A203;
  assign \new_[90645]_  = ~A266 & ~A234;
  assign \new_[90646]_  = \new_[90645]_  & \new_[90642]_ ;
  assign \new_[90649]_  = ~A269 & ~A268;
  assign \new_[90652]_  = A299 & A298;
  assign \new_[90653]_  = \new_[90652]_  & \new_[90649]_ ;
  assign \new_[90654]_  = \new_[90653]_  & \new_[90646]_ ;
  assign \new_[90658]_  = ~A167 & ~A168;
  assign \new_[90659]_  = A169 & \new_[90658]_ ;
  assign \new_[90662]_  = A199 & A166;
  assign \new_[90665]_  = A201 & ~A200;
  assign \new_[90666]_  = \new_[90665]_  & \new_[90662]_ ;
  assign \new_[90667]_  = \new_[90666]_  & \new_[90659]_ ;
  assign \new_[90670]_  = ~A233 & A203;
  assign \new_[90673]_  = ~A266 & ~A234;
  assign \new_[90674]_  = \new_[90673]_  & \new_[90670]_ ;
  assign \new_[90677]_  = ~A269 & ~A268;
  assign \new_[90680]_  = ~A299 & ~A298;
  assign \new_[90681]_  = \new_[90680]_  & \new_[90677]_ ;
  assign \new_[90682]_  = \new_[90681]_  & \new_[90674]_ ;
  assign \new_[90686]_  = ~A167 & ~A168;
  assign \new_[90687]_  = A169 & \new_[90686]_ ;
  assign \new_[90690]_  = A199 & A166;
  assign \new_[90693]_  = A201 & ~A200;
  assign \new_[90694]_  = \new_[90693]_  & \new_[90690]_ ;
  assign \new_[90695]_  = \new_[90694]_  & \new_[90687]_ ;
  assign \new_[90698]_  = ~A233 & A203;
  assign \new_[90701]_  = ~A266 & ~A234;
  assign \new_[90702]_  = \new_[90701]_  & \new_[90698]_ ;
  assign \new_[90705]_  = A298 & ~A267;
  assign \new_[90708]_  = ~A302 & ~A301;
  assign \new_[90709]_  = \new_[90708]_  & \new_[90705]_ ;
  assign \new_[90710]_  = \new_[90709]_  & \new_[90702]_ ;
  assign \new_[90714]_  = ~A167 & ~A168;
  assign \new_[90715]_  = A169 & \new_[90714]_ ;
  assign \new_[90718]_  = A199 & A166;
  assign \new_[90721]_  = A201 & ~A200;
  assign \new_[90722]_  = \new_[90721]_  & \new_[90718]_ ;
  assign \new_[90723]_  = \new_[90722]_  & \new_[90715]_ ;
  assign \new_[90726]_  = ~A233 & A203;
  assign \new_[90729]_  = ~A265 & ~A234;
  assign \new_[90730]_  = \new_[90729]_  & \new_[90726]_ ;
  assign \new_[90733]_  = A298 & ~A266;
  assign \new_[90736]_  = ~A302 & ~A301;
  assign \new_[90737]_  = \new_[90736]_  & \new_[90733]_ ;
  assign \new_[90738]_  = \new_[90737]_  & \new_[90730]_ ;
  assign \new_[90742]_  = ~A167 & ~A168;
  assign \new_[90743]_  = A169 & \new_[90742]_ ;
  assign \new_[90746]_  = A199 & A166;
  assign \new_[90749]_  = A201 & ~A200;
  assign \new_[90750]_  = \new_[90749]_  & \new_[90746]_ ;
  assign \new_[90751]_  = \new_[90750]_  & \new_[90743]_ ;
  assign \new_[90754]_  = ~A232 & A203;
  assign \new_[90757]_  = A265 & ~A233;
  assign \new_[90758]_  = \new_[90757]_  & \new_[90754]_ ;
  assign \new_[90761]_  = A298 & A266;
  assign \new_[90764]_  = ~A302 & ~A301;
  assign \new_[90765]_  = \new_[90764]_  & \new_[90761]_ ;
  assign \new_[90766]_  = \new_[90765]_  & \new_[90758]_ ;
  assign \new_[90770]_  = ~A167 & ~A168;
  assign \new_[90771]_  = A169 & \new_[90770]_ ;
  assign \new_[90774]_  = A199 & A166;
  assign \new_[90777]_  = A201 & ~A200;
  assign \new_[90778]_  = \new_[90777]_  & \new_[90774]_ ;
  assign \new_[90779]_  = \new_[90778]_  & \new_[90771]_ ;
  assign \new_[90782]_  = ~A232 & A203;
  assign \new_[90785]_  = ~A266 & ~A233;
  assign \new_[90786]_  = \new_[90785]_  & \new_[90782]_ ;
  assign \new_[90789]_  = ~A269 & ~A268;
  assign \new_[90792]_  = ~A300 & A298;
  assign \new_[90793]_  = \new_[90792]_  & \new_[90789]_ ;
  assign \new_[90794]_  = \new_[90793]_  & \new_[90786]_ ;
  assign \new_[90798]_  = ~A167 & ~A168;
  assign \new_[90799]_  = A169 & \new_[90798]_ ;
  assign \new_[90802]_  = A199 & A166;
  assign \new_[90805]_  = A201 & ~A200;
  assign \new_[90806]_  = \new_[90805]_  & \new_[90802]_ ;
  assign \new_[90807]_  = \new_[90806]_  & \new_[90799]_ ;
  assign \new_[90810]_  = ~A232 & A203;
  assign \new_[90813]_  = ~A266 & ~A233;
  assign \new_[90814]_  = \new_[90813]_  & \new_[90810]_ ;
  assign \new_[90817]_  = ~A269 & ~A268;
  assign \new_[90820]_  = A299 & A298;
  assign \new_[90821]_  = \new_[90820]_  & \new_[90817]_ ;
  assign \new_[90822]_  = \new_[90821]_  & \new_[90814]_ ;
  assign \new_[90826]_  = ~A167 & ~A168;
  assign \new_[90827]_  = A169 & \new_[90826]_ ;
  assign \new_[90830]_  = A199 & A166;
  assign \new_[90833]_  = A201 & ~A200;
  assign \new_[90834]_  = \new_[90833]_  & \new_[90830]_ ;
  assign \new_[90835]_  = \new_[90834]_  & \new_[90827]_ ;
  assign \new_[90838]_  = ~A232 & A203;
  assign \new_[90841]_  = ~A266 & ~A233;
  assign \new_[90842]_  = \new_[90841]_  & \new_[90838]_ ;
  assign \new_[90845]_  = ~A269 & ~A268;
  assign \new_[90848]_  = ~A299 & ~A298;
  assign \new_[90849]_  = \new_[90848]_  & \new_[90845]_ ;
  assign \new_[90850]_  = \new_[90849]_  & \new_[90842]_ ;
  assign \new_[90854]_  = ~A167 & ~A168;
  assign \new_[90855]_  = A169 & \new_[90854]_ ;
  assign \new_[90858]_  = A199 & A166;
  assign \new_[90861]_  = A201 & ~A200;
  assign \new_[90862]_  = \new_[90861]_  & \new_[90858]_ ;
  assign \new_[90863]_  = \new_[90862]_  & \new_[90855]_ ;
  assign \new_[90866]_  = ~A232 & A203;
  assign \new_[90869]_  = ~A266 & ~A233;
  assign \new_[90870]_  = \new_[90869]_  & \new_[90866]_ ;
  assign \new_[90873]_  = A298 & ~A267;
  assign \new_[90876]_  = ~A302 & ~A301;
  assign \new_[90877]_  = \new_[90876]_  & \new_[90873]_ ;
  assign \new_[90878]_  = \new_[90877]_  & \new_[90870]_ ;
  assign \new_[90882]_  = ~A167 & ~A168;
  assign \new_[90883]_  = A169 & \new_[90882]_ ;
  assign \new_[90886]_  = A199 & A166;
  assign \new_[90889]_  = A201 & ~A200;
  assign \new_[90890]_  = \new_[90889]_  & \new_[90886]_ ;
  assign \new_[90891]_  = \new_[90890]_  & \new_[90883]_ ;
  assign \new_[90894]_  = ~A232 & A203;
  assign \new_[90897]_  = ~A265 & ~A233;
  assign \new_[90898]_  = \new_[90897]_  & \new_[90894]_ ;
  assign \new_[90901]_  = A298 & ~A266;
  assign \new_[90904]_  = ~A302 & ~A301;
  assign \new_[90905]_  = \new_[90904]_  & \new_[90901]_ ;
  assign \new_[90906]_  = \new_[90905]_  & \new_[90898]_ ;
  assign \new_[90910]_  = ~A168 & A169;
  assign \new_[90911]_  = A170 & \new_[90910]_ ;
  assign \new_[90914]_  = ~A200 & A199;
  assign \new_[90917]_  = A202 & A201;
  assign \new_[90918]_  = \new_[90917]_  & \new_[90914]_ ;
  assign \new_[90919]_  = \new_[90918]_  & \new_[90911]_ ;
  assign \new_[90922]_  = A233 & A232;
  assign \new_[90925]_  = ~A268 & A265;
  assign \new_[90926]_  = \new_[90925]_  & \new_[90922]_ ;
  assign \new_[90929]_  = ~A299 & ~A269;
  assign \new_[90932]_  = ~A302 & ~A301;
  assign \new_[90933]_  = \new_[90932]_  & \new_[90929]_ ;
  assign \new_[90934]_  = \new_[90933]_  & \new_[90926]_ ;
  assign \new_[90938]_  = ~A168 & A169;
  assign \new_[90939]_  = A170 & \new_[90938]_ ;
  assign \new_[90942]_  = ~A200 & A199;
  assign \new_[90945]_  = A202 & A201;
  assign \new_[90946]_  = \new_[90945]_  & \new_[90942]_ ;
  assign \new_[90947]_  = \new_[90946]_  & \new_[90939]_ ;
  assign \new_[90950]_  = ~A235 & ~A233;
  assign \new_[90953]_  = A265 & ~A236;
  assign \new_[90954]_  = \new_[90953]_  & \new_[90950]_ ;
  assign \new_[90957]_  = A298 & A266;
  assign \new_[90960]_  = ~A302 & ~A301;
  assign \new_[90961]_  = \new_[90960]_  & \new_[90957]_ ;
  assign \new_[90962]_  = \new_[90961]_  & \new_[90954]_ ;
  assign \new_[90966]_  = ~A168 & A169;
  assign \new_[90967]_  = A170 & \new_[90966]_ ;
  assign \new_[90970]_  = ~A200 & A199;
  assign \new_[90973]_  = A202 & A201;
  assign \new_[90974]_  = \new_[90973]_  & \new_[90970]_ ;
  assign \new_[90975]_  = \new_[90974]_  & \new_[90967]_ ;
  assign \new_[90978]_  = ~A235 & ~A233;
  assign \new_[90981]_  = ~A266 & ~A236;
  assign \new_[90982]_  = \new_[90981]_  & \new_[90978]_ ;
  assign \new_[90985]_  = ~A269 & ~A268;
  assign \new_[90988]_  = ~A300 & A298;
  assign \new_[90989]_  = \new_[90988]_  & \new_[90985]_ ;
  assign \new_[90990]_  = \new_[90989]_  & \new_[90982]_ ;
  assign \new_[90994]_  = ~A168 & A169;
  assign \new_[90995]_  = A170 & \new_[90994]_ ;
  assign \new_[90998]_  = ~A200 & A199;
  assign \new_[91001]_  = A202 & A201;
  assign \new_[91002]_  = \new_[91001]_  & \new_[90998]_ ;
  assign \new_[91003]_  = \new_[91002]_  & \new_[90995]_ ;
  assign \new_[91006]_  = ~A235 & ~A233;
  assign \new_[91009]_  = ~A266 & ~A236;
  assign \new_[91010]_  = \new_[91009]_  & \new_[91006]_ ;
  assign \new_[91013]_  = ~A269 & ~A268;
  assign \new_[91016]_  = A299 & A298;
  assign \new_[91017]_  = \new_[91016]_  & \new_[91013]_ ;
  assign \new_[91018]_  = \new_[91017]_  & \new_[91010]_ ;
  assign \new_[91022]_  = ~A168 & A169;
  assign \new_[91023]_  = A170 & \new_[91022]_ ;
  assign \new_[91026]_  = ~A200 & A199;
  assign \new_[91029]_  = A202 & A201;
  assign \new_[91030]_  = \new_[91029]_  & \new_[91026]_ ;
  assign \new_[91031]_  = \new_[91030]_  & \new_[91023]_ ;
  assign \new_[91034]_  = ~A235 & ~A233;
  assign \new_[91037]_  = ~A266 & ~A236;
  assign \new_[91038]_  = \new_[91037]_  & \new_[91034]_ ;
  assign \new_[91041]_  = ~A269 & ~A268;
  assign \new_[91044]_  = ~A299 & ~A298;
  assign \new_[91045]_  = \new_[91044]_  & \new_[91041]_ ;
  assign \new_[91046]_  = \new_[91045]_  & \new_[91038]_ ;
  assign \new_[91050]_  = ~A168 & A169;
  assign \new_[91051]_  = A170 & \new_[91050]_ ;
  assign \new_[91054]_  = ~A200 & A199;
  assign \new_[91057]_  = A202 & A201;
  assign \new_[91058]_  = \new_[91057]_  & \new_[91054]_ ;
  assign \new_[91059]_  = \new_[91058]_  & \new_[91051]_ ;
  assign \new_[91062]_  = ~A235 & ~A233;
  assign \new_[91065]_  = ~A266 & ~A236;
  assign \new_[91066]_  = \new_[91065]_  & \new_[91062]_ ;
  assign \new_[91069]_  = A298 & ~A267;
  assign \new_[91072]_  = ~A302 & ~A301;
  assign \new_[91073]_  = \new_[91072]_  & \new_[91069]_ ;
  assign \new_[91074]_  = \new_[91073]_  & \new_[91066]_ ;
  assign \new_[91078]_  = ~A168 & A169;
  assign \new_[91079]_  = A170 & \new_[91078]_ ;
  assign \new_[91082]_  = ~A200 & A199;
  assign \new_[91085]_  = A202 & A201;
  assign \new_[91086]_  = \new_[91085]_  & \new_[91082]_ ;
  assign \new_[91087]_  = \new_[91086]_  & \new_[91079]_ ;
  assign \new_[91090]_  = ~A235 & ~A233;
  assign \new_[91093]_  = ~A265 & ~A236;
  assign \new_[91094]_  = \new_[91093]_  & \new_[91090]_ ;
  assign \new_[91097]_  = A298 & ~A266;
  assign \new_[91100]_  = ~A302 & ~A301;
  assign \new_[91101]_  = \new_[91100]_  & \new_[91097]_ ;
  assign \new_[91102]_  = \new_[91101]_  & \new_[91094]_ ;
  assign \new_[91106]_  = ~A168 & A169;
  assign \new_[91107]_  = A170 & \new_[91106]_ ;
  assign \new_[91110]_  = ~A200 & A199;
  assign \new_[91113]_  = A202 & A201;
  assign \new_[91114]_  = \new_[91113]_  & \new_[91110]_ ;
  assign \new_[91115]_  = \new_[91114]_  & \new_[91107]_ ;
  assign \new_[91118]_  = ~A234 & ~A233;
  assign \new_[91121]_  = ~A268 & ~A266;
  assign \new_[91122]_  = \new_[91121]_  & \new_[91118]_ ;
  assign \new_[91125]_  = A298 & ~A269;
  assign \new_[91128]_  = ~A302 & ~A301;
  assign \new_[91129]_  = \new_[91128]_  & \new_[91125]_ ;
  assign \new_[91130]_  = \new_[91129]_  & \new_[91122]_ ;
  assign \new_[91134]_  = ~A168 & A169;
  assign \new_[91135]_  = A170 & \new_[91134]_ ;
  assign \new_[91138]_  = ~A200 & A199;
  assign \new_[91141]_  = A202 & A201;
  assign \new_[91142]_  = \new_[91141]_  & \new_[91138]_ ;
  assign \new_[91143]_  = \new_[91142]_  & \new_[91135]_ ;
  assign \new_[91146]_  = ~A233 & A232;
  assign \new_[91149]_  = A235 & A234;
  assign \new_[91150]_  = \new_[91149]_  & \new_[91146]_ ;
  assign \new_[91153]_  = ~A299 & A298;
  assign \new_[91156]_  = A301 & A300;
  assign \new_[91157]_  = \new_[91156]_  & \new_[91153]_ ;
  assign \new_[91158]_  = \new_[91157]_  & \new_[91150]_ ;
  assign \new_[91162]_  = ~A168 & A169;
  assign \new_[91163]_  = A170 & \new_[91162]_ ;
  assign \new_[91166]_  = ~A200 & A199;
  assign \new_[91169]_  = A202 & A201;
  assign \new_[91170]_  = \new_[91169]_  & \new_[91166]_ ;
  assign \new_[91171]_  = \new_[91170]_  & \new_[91163]_ ;
  assign \new_[91174]_  = ~A233 & A232;
  assign \new_[91177]_  = A235 & A234;
  assign \new_[91178]_  = \new_[91177]_  & \new_[91174]_ ;
  assign \new_[91181]_  = ~A299 & A298;
  assign \new_[91184]_  = A302 & A300;
  assign \new_[91185]_  = \new_[91184]_  & \new_[91181]_ ;
  assign \new_[91186]_  = \new_[91185]_  & \new_[91178]_ ;
  assign \new_[91190]_  = ~A168 & A169;
  assign \new_[91191]_  = A170 & \new_[91190]_ ;
  assign \new_[91194]_  = ~A200 & A199;
  assign \new_[91197]_  = A202 & A201;
  assign \new_[91198]_  = \new_[91197]_  & \new_[91194]_ ;
  assign \new_[91199]_  = \new_[91198]_  & \new_[91191]_ ;
  assign \new_[91202]_  = ~A233 & A232;
  assign \new_[91205]_  = A235 & A234;
  assign \new_[91206]_  = \new_[91205]_  & \new_[91202]_ ;
  assign \new_[91209]_  = ~A266 & A265;
  assign \new_[91212]_  = A268 & A267;
  assign \new_[91213]_  = \new_[91212]_  & \new_[91209]_ ;
  assign \new_[91214]_  = \new_[91213]_  & \new_[91206]_ ;
  assign \new_[91218]_  = ~A168 & A169;
  assign \new_[91219]_  = A170 & \new_[91218]_ ;
  assign \new_[91222]_  = ~A200 & A199;
  assign \new_[91225]_  = A202 & A201;
  assign \new_[91226]_  = \new_[91225]_  & \new_[91222]_ ;
  assign \new_[91227]_  = \new_[91226]_  & \new_[91219]_ ;
  assign \new_[91230]_  = ~A233 & A232;
  assign \new_[91233]_  = A235 & A234;
  assign \new_[91234]_  = \new_[91233]_  & \new_[91230]_ ;
  assign \new_[91237]_  = ~A266 & A265;
  assign \new_[91240]_  = A269 & A267;
  assign \new_[91241]_  = \new_[91240]_  & \new_[91237]_ ;
  assign \new_[91242]_  = \new_[91241]_  & \new_[91234]_ ;
  assign \new_[91246]_  = ~A168 & A169;
  assign \new_[91247]_  = A170 & \new_[91246]_ ;
  assign \new_[91250]_  = ~A200 & A199;
  assign \new_[91253]_  = A202 & A201;
  assign \new_[91254]_  = \new_[91253]_  & \new_[91250]_ ;
  assign \new_[91255]_  = \new_[91254]_  & \new_[91247]_ ;
  assign \new_[91258]_  = ~A233 & A232;
  assign \new_[91261]_  = A236 & A234;
  assign \new_[91262]_  = \new_[91261]_  & \new_[91258]_ ;
  assign \new_[91265]_  = ~A299 & A298;
  assign \new_[91268]_  = A301 & A300;
  assign \new_[91269]_  = \new_[91268]_  & \new_[91265]_ ;
  assign \new_[91270]_  = \new_[91269]_  & \new_[91262]_ ;
  assign \new_[91274]_  = ~A168 & A169;
  assign \new_[91275]_  = A170 & \new_[91274]_ ;
  assign \new_[91278]_  = ~A200 & A199;
  assign \new_[91281]_  = A202 & A201;
  assign \new_[91282]_  = \new_[91281]_  & \new_[91278]_ ;
  assign \new_[91283]_  = \new_[91282]_  & \new_[91275]_ ;
  assign \new_[91286]_  = ~A233 & A232;
  assign \new_[91289]_  = A236 & A234;
  assign \new_[91290]_  = \new_[91289]_  & \new_[91286]_ ;
  assign \new_[91293]_  = ~A299 & A298;
  assign \new_[91296]_  = A302 & A300;
  assign \new_[91297]_  = \new_[91296]_  & \new_[91293]_ ;
  assign \new_[91298]_  = \new_[91297]_  & \new_[91290]_ ;
  assign \new_[91302]_  = ~A168 & A169;
  assign \new_[91303]_  = A170 & \new_[91302]_ ;
  assign \new_[91306]_  = ~A200 & A199;
  assign \new_[91309]_  = A202 & A201;
  assign \new_[91310]_  = \new_[91309]_  & \new_[91306]_ ;
  assign \new_[91311]_  = \new_[91310]_  & \new_[91303]_ ;
  assign \new_[91314]_  = ~A233 & A232;
  assign \new_[91317]_  = A236 & A234;
  assign \new_[91318]_  = \new_[91317]_  & \new_[91314]_ ;
  assign \new_[91321]_  = ~A266 & A265;
  assign \new_[91324]_  = A268 & A267;
  assign \new_[91325]_  = \new_[91324]_  & \new_[91321]_ ;
  assign \new_[91326]_  = \new_[91325]_  & \new_[91318]_ ;
  assign \new_[91330]_  = ~A168 & A169;
  assign \new_[91331]_  = A170 & \new_[91330]_ ;
  assign \new_[91334]_  = ~A200 & A199;
  assign \new_[91337]_  = A202 & A201;
  assign \new_[91338]_  = \new_[91337]_  & \new_[91334]_ ;
  assign \new_[91339]_  = \new_[91338]_  & \new_[91331]_ ;
  assign \new_[91342]_  = ~A233 & A232;
  assign \new_[91345]_  = A236 & A234;
  assign \new_[91346]_  = \new_[91345]_  & \new_[91342]_ ;
  assign \new_[91349]_  = ~A266 & A265;
  assign \new_[91352]_  = A269 & A267;
  assign \new_[91353]_  = \new_[91352]_  & \new_[91349]_ ;
  assign \new_[91354]_  = \new_[91353]_  & \new_[91346]_ ;
  assign \new_[91358]_  = ~A168 & A169;
  assign \new_[91359]_  = A170 & \new_[91358]_ ;
  assign \new_[91362]_  = ~A200 & A199;
  assign \new_[91365]_  = A202 & A201;
  assign \new_[91366]_  = \new_[91365]_  & \new_[91362]_ ;
  assign \new_[91367]_  = \new_[91366]_  & \new_[91359]_ ;
  assign \new_[91370]_  = ~A233 & ~A232;
  assign \new_[91373]_  = ~A268 & ~A266;
  assign \new_[91374]_  = \new_[91373]_  & \new_[91370]_ ;
  assign \new_[91377]_  = A298 & ~A269;
  assign \new_[91380]_  = ~A302 & ~A301;
  assign \new_[91381]_  = \new_[91380]_  & \new_[91377]_ ;
  assign \new_[91382]_  = \new_[91381]_  & \new_[91374]_ ;
  assign \new_[91386]_  = ~A168 & A169;
  assign \new_[91387]_  = A170 & \new_[91386]_ ;
  assign \new_[91390]_  = ~A200 & A199;
  assign \new_[91393]_  = A203 & A201;
  assign \new_[91394]_  = \new_[91393]_  & \new_[91390]_ ;
  assign \new_[91395]_  = \new_[91394]_  & \new_[91387]_ ;
  assign \new_[91398]_  = A233 & A232;
  assign \new_[91401]_  = ~A268 & A265;
  assign \new_[91402]_  = \new_[91401]_  & \new_[91398]_ ;
  assign \new_[91405]_  = ~A299 & ~A269;
  assign \new_[91408]_  = ~A302 & ~A301;
  assign \new_[91409]_  = \new_[91408]_  & \new_[91405]_ ;
  assign \new_[91410]_  = \new_[91409]_  & \new_[91402]_ ;
  assign \new_[91414]_  = ~A168 & A169;
  assign \new_[91415]_  = A170 & \new_[91414]_ ;
  assign \new_[91418]_  = ~A200 & A199;
  assign \new_[91421]_  = A203 & A201;
  assign \new_[91422]_  = \new_[91421]_  & \new_[91418]_ ;
  assign \new_[91423]_  = \new_[91422]_  & \new_[91415]_ ;
  assign \new_[91426]_  = ~A235 & ~A233;
  assign \new_[91429]_  = A265 & ~A236;
  assign \new_[91430]_  = \new_[91429]_  & \new_[91426]_ ;
  assign \new_[91433]_  = A298 & A266;
  assign \new_[91436]_  = ~A302 & ~A301;
  assign \new_[91437]_  = \new_[91436]_  & \new_[91433]_ ;
  assign \new_[91438]_  = \new_[91437]_  & \new_[91430]_ ;
  assign \new_[91442]_  = ~A168 & A169;
  assign \new_[91443]_  = A170 & \new_[91442]_ ;
  assign \new_[91446]_  = ~A200 & A199;
  assign \new_[91449]_  = A203 & A201;
  assign \new_[91450]_  = \new_[91449]_  & \new_[91446]_ ;
  assign \new_[91451]_  = \new_[91450]_  & \new_[91443]_ ;
  assign \new_[91454]_  = ~A235 & ~A233;
  assign \new_[91457]_  = ~A266 & ~A236;
  assign \new_[91458]_  = \new_[91457]_  & \new_[91454]_ ;
  assign \new_[91461]_  = ~A269 & ~A268;
  assign \new_[91464]_  = ~A300 & A298;
  assign \new_[91465]_  = \new_[91464]_  & \new_[91461]_ ;
  assign \new_[91466]_  = \new_[91465]_  & \new_[91458]_ ;
  assign \new_[91470]_  = ~A168 & A169;
  assign \new_[91471]_  = A170 & \new_[91470]_ ;
  assign \new_[91474]_  = ~A200 & A199;
  assign \new_[91477]_  = A203 & A201;
  assign \new_[91478]_  = \new_[91477]_  & \new_[91474]_ ;
  assign \new_[91479]_  = \new_[91478]_  & \new_[91471]_ ;
  assign \new_[91482]_  = ~A235 & ~A233;
  assign \new_[91485]_  = ~A266 & ~A236;
  assign \new_[91486]_  = \new_[91485]_  & \new_[91482]_ ;
  assign \new_[91489]_  = ~A269 & ~A268;
  assign \new_[91492]_  = A299 & A298;
  assign \new_[91493]_  = \new_[91492]_  & \new_[91489]_ ;
  assign \new_[91494]_  = \new_[91493]_  & \new_[91486]_ ;
  assign \new_[91498]_  = ~A168 & A169;
  assign \new_[91499]_  = A170 & \new_[91498]_ ;
  assign \new_[91502]_  = ~A200 & A199;
  assign \new_[91505]_  = A203 & A201;
  assign \new_[91506]_  = \new_[91505]_  & \new_[91502]_ ;
  assign \new_[91507]_  = \new_[91506]_  & \new_[91499]_ ;
  assign \new_[91510]_  = ~A235 & ~A233;
  assign \new_[91513]_  = ~A266 & ~A236;
  assign \new_[91514]_  = \new_[91513]_  & \new_[91510]_ ;
  assign \new_[91517]_  = ~A269 & ~A268;
  assign \new_[91520]_  = ~A299 & ~A298;
  assign \new_[91521]_  = \new_[91520]_  & \new_[91517]_ ;
  assign \new_[91522]_  = \new_[91521]_  & \new_[91514]_ ;
  assign \new_[91526]_  = ~A168 & A169;
  assign \new_[91527]_  = A170 & \new_[91526]_ ;
  assign \new_[91530]_  = ~A200 & A199;
  assign \new_[91533]_  = A203 & A201;
  assign \new_[91534]_  = \new_[91533]_  & \new_[91530]_ ;
  assign \new_[91535]_  = \new_[91534]_  & \new_[91527]_ ;
  assign \new_[91538]_  = ~A235 & ~A233;
  assign \new_[91541]_  = ~A266 & ~A236;
  assign \new_[91542]_  = \new_[91541]_  & \new_[91538]_ ;
  assign \new_[91545]_  = A298 & ~A267;
  assign \new_[91548]_  = ~A302 & ~A301;
  assign \new_[91549]_  = \new_[91548]_  & \new_[91545]_ ;
  assign \new_[91550]_  = \new_[91549]_  & \new_[91542]_ ;
  assign \new_[91554]_  = ~A168 & A169;
  assign \new_[91555]_  = A170 & \new_[91554]_ ;
  assign \new_[91558]_  = ~A200 & A199;
  assign \new_[91561]_  = A203 & A201;
  assign \new_[91562]_  = \new_[91561]_  & \new_[91558]_ ;
  assign \new_[91563]_  = \new_[91562]_  & \new_[91555]_ ;
  assign \new_[91566]_  = ~A235 & ~A233;
  assign \new_[91569]_  = ~A265 & ~A236;
  assign \new_[91570]_  = \new_[91569]_  & \new_[91566]_ ;
  assign \new_[91573]_  = A298 & ~A266;
  assign \new_[91576]_  = ~A302 & ~A301;
  assign \new_[91577]_  = \new_[91576]_  & \new_[91573]_ ;
  assign \new_[91578]_  = \new_[91577]_  & \new_[91570]_ ;
  assign \new_[91582]_  = ~A168 & A169;
  assign \new_[91583]_  = A170 & \new_[91582]_ ;
  assign \new_[91586]_  = ~A200 & A199;
  assign \new_[91589]_  = A203 & A201;
  assign \new_[91590]_  = \new_[91589]_  & \new_[91586]_ ;
  assign \new_[91591]_  = \new_[91590]_  & \new_[91583]_ ;
  assign \new_[91594]_  = ~A234 & ~A233;
  assign \new_[91597]_  = ~A268 & ~A266;
  assign \new_[91598]_  = \new_[91597]_  & \new_[91594]_ ;
  assign \new_[91601]_  = A298 & ~A269;
  assign \new_[91604]_  = ~A302 & ~A301;
  assign \new_[91605]_  = \new_[91604]_  & \new_[91601]_ ;
  assign \new_[91606]_  = \new_[91605]_  & \new_[91598]_ ;
  assign \new_[91610]_  = ~A168 & A169;
  assign \new_[91611]_  = A170 & \new_[91610]_ ;
  assign \new_[91614]_  = ~A200 & A199;
  assign \new_[91617]_  = A203 & A201;
  assign \new_[91618]_  = \new_[91617]_  & \new_[91614]_ ;
  assign \new_[91619]_  = \new_[91618]_  & \new_[91611]_ ;
  assign \new_[91622]_  = ~A233 & A232;
  assign \new_[91625]_  = A235 & A234;
  assign \new_[91626]_  = \new_[91625]_  & \new_[91622]_ ;
  assign \new_[91629]_  = ~A299 & A298;
  assign \new_[91632]_  = A301 & A300;
  assign \new_[91633]_  = \new_[91632]_  & \new_[91629]_ ;
  assign \new_[91634]_  = \new_[91633]_  & \new_[91626]_ ;
  assign \new_[91638]_  = ~A168 & A169;
  assign \new_[91639]_  = A170 & \new_[91638]_ ;
  assign \new_[91642]_  = ~A200 & A199;
  assign \new_[91645]_  = A203 & A201;
  assign \new_[91646]_  = \new_[91645]_  & \new_[91642]_ ;
  assign \new_[91647]_  = \new_[91646]_  & \new_[91639]_ ;
  assign \new_[91650]_  = ~A233 & A232;
  assign \new_[91653]_  = A235 & A234;
  assign \new_[91654]_  = \new_[91653]_  & \new_[91650]_ ;
  assign \new_[91657]_  = ~A299 & A298;
  assign \new_[91660]_  = A302 & A300;
  assign \new_[91661]_  = \new_[91660]_  & \new_[91657]_ ;
  assign \new_[91662]_  = \new_[91661]_  & \new_[91654]_ ;
  assign \new_[91666]_  = ~A168 & A169;
  assign \new_[91667]_  = A170 & \new_[91666]_ ;
  assign \new_[91670]_  = ~A200 & A199;
  assign \new_[91673]_  = A203 & A201;
  assign \new_[91674]_  = \new_[91673]_  & \new_[91670]_ ;
  assign \new_[91675]_  = \new_[91674]_  & \new_[91667]_ ;
  assign \new_[91678]_  = ~A233 & A232;
  assign \new_[91681]_  = A235 & A234;
  assign \new_[91682]_  = \new_[91681]_  & \new_[91678]_ ;
  assign \new_[91685]_  = ~A266 & A265;
  assign \new_[91688]_  = A268 & A267;
  assign \new_[91689]_  = \new_[91688]_  & \new_[91685]_ ;
  assign \new_[91690]_  = \new_[91689]_  & \new_[91682]_ ;
  assign \new_[91694]_  = ~A168 & A169;
  assign \new_[91695]_  = A170 & \new_[91694]_ ;
  assign \new_[91698]_  = ~A200 & A199;
  assign \new_[91701]_  = A203 & A201;
  assign \new_[91702]_  = \new_[91701]_  & \new_[91698]_ ;
  assign \new_[91703]_  = \new_[91702]_  & \new_[91695]_ ;
  assign \new_[91706]_  = ~A233 & A232;
  assign \new_[91709]_  = A235 & A234;
  assign \new_[91710]_  = \new_[91709]_  & \new_[91706]_ ;
  assign \new_[91713]_  = ~A266 & A265;
  assign \new_[91716]_  = A269 & A267;
  assign \new_[91717]_  = \new_[91716]_  & \new_[91713]_ ;
  assign \new_[91718]_  = \new_[91717]_  & \new_[91710]_ ;
  assign \new_[91722]_  = ~A168 & A169;
  assign \new_[91723]_  = A170 & \new_[91722]_ ;
  assign \new_[91726]_  = ~A200 & A199;
  assign \new_[91729]_  = A203 & A201;
  assign \new_[91730]_  = \new_[91729]_  & \new_[91726]_ ;
  assign \new_[91731]_  = \new_[91730]_  & \new_[91723]_ ;
  assign \new_[91734]_  = ~A233 & A232;
  assign \new_[91737]_  = A236 & A234;
  assign \new_[91738]_  = \new_[91737]_  & \new_[91734]_ ;
  assign \new_[91741]_  = ~A299 & A298;
  assign \new_[91744]_  = A301 & A300;
  assign \new_[91745]_  = \new_[91744]_  & \new_[91741]_ ;
  assign \new_[91746]_  = \new_[91745]_  & \new_[91738]_ ;
  assign \new_[91750]_  = ~A168 & A169;
  assign \new_[91751]_  = A170 & \new_[91750]_ ;
  assign \new_[91754]_  = ~A200 & A199;
  assign \new_[91757]_  = A203 & A201;
  assign \new_[91758]_  = \new_[91757]_  & \new_[91754]_ ;
  assign \new_[91759]_  = \new_[91758]_  & \new_[91751]_ ;
  assign \new_[91762]_  = ~A233 & A232;
  assign \new_[91765]_  = A236 & A234;
  assign \new_[91766]_  = \new_[91765]_  & \new_[91762]_ ;
  assign \new_[91769]_  = ~A299 & A298;
  assign \new_[91772]_  = A302 & A300;
  assign \new_[91773]_  = \new_[91772]_  & \new_[91769]_ ;
  assign \new_[91774]_  = \new_[91773]_  & \new_[91766]_ ;
  assign \new_[91778]_  = ~A168 & A169;
  assign \new_[91779]_  = A170 & \new_[91778]_ ;
  assign \new_[91782]_  = ~A200 & A199;
  assign \new_[91785]_  = A203 & A201;
  assign \new_[91786]_  = \new_[91785]_  & \new_[91782]_ ;
  assign \new_[91787]_  = \new_[91786]_  & \new_[91779]_ ;
  assign \new_[91790]_  = ~A233 & A232;
  assign \new_[91793]_  = A236 & A234;
  assign \new_[91794]_  = \new_[91793]_  & \new_[91790]_ ;
  assign \new_[91797]_  = ~A266 & A265;
  assign \new_[91800]_  = A268 & A267;
  assign \new_[91801]_  = \new_[91800]_  & \new_[91797]_ ;
  assign \new_[91802]_  = \new_[91801]_  & \new_[91794]_ ;
  assign \new_[91806]_  = ~A168 & A169;
  assign \new_[91807]_  = A170 & \new_[91806]_ ;
  assign \new_[91810]_  = ~A200 & A199;
  assign \new_[91813]_  = A203 & A201;
  assign \new_[91814]_  = \new_[91813]_  & \new_[91810]_ ;
  assign \new_[91815]_  = \new_[91814]_  & \new_[91807]_ ;
  assign \new_[91818]_  = ~A233 & A232;
  assign \new_[91821]_  = A236 & A234;
  assign \new_[91822]_  = \new_[91821]_  & \new_[91818]_ ;
  assign \new_[91825]_  = ~A266 & A265;
  assign \new_[91828]_  = A269 & A267;
  assign \new_[91829]_  = \new_[91828]_  & \new_[91825]_ ;
  assign \new_[91830]_  = \new_[91829]_  & \new_[91822]_ ;
  assign \new_[91834]_  = ~A168 & A169;
  assign \new_[91835]_  = A170 & \new_[91834]_ ;
  assign \new_[91838]_  = ~A200 & A199;
  assign \new_[91841]_  = A203 & A201;
  assign \new_[91842]_  = \new_[91841]_  & \new_[91838]_ ;
  assign \new_[91843]_  = \new_[91842]_  & \new_[91835]_ ;
  assign \new_[91846]_  = ~A233 & ~A232;
  assign \new_[91849]_  = ~A268 & ~A266;
  assign \new_[91850]_  = \new_[91849]_  & \new_[91846]_ ;
  assign \new_[91853]_  = A298 & ~A269;
  assign \new_[91856]_  = ~A302 & ~A301;
  assign \new_[91857]_  = \new_[91856]_  & \new_[91853]_ ;
  assign \new_[91858]_  = \new_[91857]_  & \new_[91850]_ ;
  assign \new_[91862]_  = A167 & A169;
  assign \new_[91863]_  = ~A170 & \new_[91862]_ ;
  assign \new_[91866]_  = A199 & A166;
  assign \new_[91869]_  = ~A233 & A200;
  assign \new_[91870]_  = \new_[91869]_  & \new_[91866]_ ;
  assign \new_[91871]_  = \new_[91870]_  & \new_[91863]_ ;
  assign \new_[91874]_  = ~A236 & ~A235;
  assign \new_[91877]_  = ~A268 & ~A266;
  assign \new_[91878]_  = \new_[91877]_  & \new_[91874]_ ;
  assign \new_[91881]_  = A298 & ~A269;
  assign \new_[91884]_  = ~A302 & ~A301;
  assign \new_[91885]_  = \new_[91884]_  & \new_[91881]_ ;
  assign \new_[91886]_  = \new_[91885]_  & \new_[91878]_ ;
  assign \new_[91890]_  = A167 & A169;
  assign \new_[91891]_  = ~A170 & \new_[91890]_ ;
  assign \new_[91894]_  = ~A200 & A166;
  assign \new_[91897]_  = ~A203 & ~A202;
  assign \new_[91898]_  = \new_[91897]_  & \new_[91894]_ ;
  assign \new_[91899]_  = \new_[91898]_  & \new_[91891]_ ;
  assign \new_[91902]_  = A233 & A232;
  assign \new_[91905]_  = ~A268 & A265;
  assign \new_[91906]_  = \new_[91905]_  & \new_[91902]_ ;
  assign \new_[91909]_  = ~A299 & ~A269;
  assign \new_[91912]_  = ~A302 & ~A301;
  assign \new_[91913]_  = \new_[91912]_  & \new_[91909]_ ;
  assign \new_[91914]_  = \new_[91913]_  & \new_[91906]_ ;
  assign \new_[91918]_  = A167 & A169;
  assign \new_[91919]_  = ~A170 & \new_[91918]_ ;
  assign \new_[91922]_  = ~A200 & A166;
  assign \new_[91925]_  = ~A203 & ~A202;
  assign \new_[91926]_  = \new_[91925]_  & \new_[91922]_ ;
  assign \new_[91927]_  = \new_[91926]_  & \new_[91919]_ ;
  assign \new_[91930]_  = ~A235 & ~A233;
  assign \new_[91933]_  = A265 & ~A236;
  assign \new_[91934]_  = \new_[91933]_  & \new_[91930]_ ;
  assign \new_[91937]_  = A298 & A266;
  assign \new_[91940]_  = ~A302 & ~A301;
  assign \new_[91941]_  = \new_[91940]_  & \new_[91937]_ ;
  assign \new_[91942]_  = \new_[91941]_  & \new_[91934]_ ;
  assign \new_[91946]_  = A167 & A169;
  assign \new_[91947]_  = ~A170 & \new_[91946]_ ;
  assign \new_[91950]_  = ~A200 & A166;
  assign \new_[91953]_  = ~A203 & ~A202;
  assign \new_[91954]_  = \new_[91953]_  & \new_[91950]_ ;
  assign \new_[91955]_  = \new_[91954]_  & \new_[91947]_ ;
  assign \new_[91958]_  = ~A235 & ~A233;
  assign \new_[91961]_  = ~A266 & ~A236;
  assign \new_[91962]_  = \new_[91961]_  & \new_[91958]_ ;
  assign \new_[91965]_  = ~A269 & ~A268;
  assign \new_[91968]_  = ~A300 & A298;
  assign \new_[91969]_  = \new_[91968]_  & \new_[91965]_ ;
  assign \new_[91970]_  = \new_[91969]_  & \new_[91962]_ ;
  assign \new_[91974]_  = A167 & A169;
  assign \new_[91975]_  = ~A170 & \new_[91974]_ ;
  assign \new_[91978]_  = ~A200 & A166;
  assign \new_[91981]_  = ~A203 & ~A202;
  assign \new_[91982]_  = \new_[91981]_  & \new_[91978]_ ;
  assign \new_[91983]_  = \new_[91982]_  & \new_[91975]_ ;
  assign \new_[91986]_  = ~A235 & ~A233;
  assign \new_[91989]_  = ~A266 & ~A236;
  assign \new_[91990]_  = \new_[91989]_  & \new_[91986]_ ;
  assign \new_[91993]_  = ~A269 & ~A268;
  assign \new_[91996]_  = A299 & A298;
  assign \new_[91997]_  = \new_[91996]_  & \new_[91993]_ ;
  assign \new_[91998]_  = \new_[91997]_  & \new_[91990]_ ;
  assign \new_[92002]_  = A167 & A169;
  assign \new_[92003]_  = ~A170 & \new_[92002]_ ;
  assign \new_[92006]_  = ~A200 & A166;
  assign \new_[92009]_  = ~A203 & ~A202;
  assign \new_[92010]_  = \new_[92009]_  & \new_[92006]_ ;
  assign \new_[92011]_  = \new_[92010]_  & \new_[92003]_ ;
  assign \new_[92014]_  = ~A235 & ~A233;
  assign \new_[92017]_  = ~A266 & ~A236;
  assign \new_[92018]_  = \new_[92017]_  & \new_[92014]_ ;
  assign \new_[92021]_  = ~A269 & ~A268;
  assign \new_[92024]_  = ~A299 & ~A298;
  assign \new_[92025]_  = \new_[92024]_  & \new_[92021]_ ;
  assign \new_[92026]_  = \new_[92025]_  & \new_[92018]_ ;
  assign \new_[92030]_  = A167 & A169;
  assign \new_[92031]_  = ~A170 & \new_[92030]_ ;
  assign \new_[92034]_  = ~A200 & A166;
  assign \new_[92037]_  = ~A203 & ~A202;
  assign \new_[92038]_  = \new_[92037]_  & \new_[92034]_ ;
  assign \new_[92039]_  = \new_[92038]_  & \new_[92031]_ ;
  assign \new_[92042]_  = ~A235 & ~A233;
  assign \new_[92045]_  = ~A266 & ~A236;
  assign \new_[92046]_  = \new_[92045]_  & \new_[92042]_ ;
  assign \new_[92049]_  = A298 & ~A267;
  assign \new_[92052]_  = ~A302 & ~A301;
  assign \new_[92053]_  = \new_[92052]_  & \new_[92049]_ ;
  assign \new_[92054]_  = \new_[92053]_  & \new_[92046]_ ;
  assign \new_[92058]_  = A167 & A169;
  assign \new_[92059]_  = ~A170 & \new_[92058]_ ;
  assign \new_[92062]_  = ~A200 & A166;
  assign \new_[92065]_  = ~A203 & ~A202;
  assign \new_[92066]_  = \new_[92065]_  & \new_[92062]_ ;
  assign \new_[92067]_  = \new_[92066]_  & \new_[92059]_ ;
  assign \new_[92070]_  = ~A235 & ~A233;
  assign \new_[92073]_  = ~A265 & ~A236;
  assign \new_[92074]_  = \new_[92073]_  & \new_[92070]_ ;
  assign \new_[92077]_  = A298 & ~A266;
  assign \new_[92080]_  = ~A302 & ~A301;
  assign \new_[92081]_  = \new_[92080]_  & \new_[92077]_ ;
  assign \new_[92082]_  = \new_[92081]_  & \new_[92074]_ ;
  assign \new_[92086]_  = A167 & A169;
  assign \new_[92087]_  = ~A170 & \new_[92086]_ ;
  assign \new_[92090]_  = ~A200 & A166;
  assign \new_[92093]_  = ~A203 & ~A202;
  assign \new_[92094]_  = \new_[92093]_  & \new_[92090]_ ;
  assign \new_[92095]_  = \new_[92094]_  & \new_[92087]_ ;
  assign \new_[92098]_  = ~A234 & ~A233;
  assign \new_[92101]_  = ~A268 & ~A266;
  assign \new_[92102]_  = \new_[92101]_  & \new_[92098]_ ;
  assign \new_[92105]_  = A298 & ~A269;
  assign \new_[92108]_  = ~A302 & ~A301;
  assign \new_[92109]_  = \new_[92108]_  & \new_[92105]_ ;
  assign \new_[92110]_  = \new_[92109]_  & \new_[92102]_ ;
  assign \new_[92114]_  = A167 & A169;
  assign \new_[92115]_  = ~A170 & \new_[92114]_ ;
  assign \new_[92118]_  = ~A200 & A166;
  assign \new_[92121]_  = ~A203 & ~A202;
  assign \new_[92122]_  = \new_[92121]_  & \new_[92118]_ ;
  assign \new_[92123]_  = \new_[92122]_  & \new_[92115]_ ;
  assign \new_[92126]_  = ~A233 & A232;
  assign \new_[92129]_  = A235 & A234;
  assign \new_[92130]_  = \new_[92129]_  & \new_[92126]_ ;
  assign \new_[92133]_  = ~A299 & A298;
  assign \new_[92136]_  = A301 & A300;
  assign \new_[92137]_  = \new_[92136]_  & \new_[92133]_ ;
  assign \new_[92138]_  = \new_[92137]_  & \new_[92130]_ ;
  assign \new_[92142]_  = A167 & A169;
  assign \new_[92143]_  = ~A170 & \new_[92142]_ ;
  assign \new_[92146]_  = ~A200 & A166;
  assign \new_[92149]_  = ~A203 & ~A202;
  assign \new_[92150]_  = \new_[92149]_  & \new_[92146]_ ;
  assign \new_[92151]_  = \new_[92150]_  & \new_[92143]_ ;
  assign \new_[92154]_  = ~A233 & A232;
  assign \new_[92157]_  = A235 & A234;
  assign \new_[92158]_  = \new_[92157]_  & \new_[92154]_ ;
  assign \new_[92161]_  = ~A299 & A298;
  assign \new_[92164]_  = A302 & A300;
  assign \new_[92165]_  = \new_[92164]_  & \new_[92161]_ ;
  assign \new_[92166]_  = \new_[92165]_  & \new_[92158]_ ;
  assign \new_[92170]_  = A167 & A169;
  assign \new_[92171]_  = ~A170 & \new_[92170]_ ;
  assign \new_[92174]_  = ~A200 & A166;
  assign \new_[92177]_  = ~A203 & ~A202;
  assign \new_[92178]_  = \new_[92177]_  & \new_[92174]_ ;
  assign \new_[92179]_  = \new_[92178]_  & \new_[92171]_ ;
  assign \new_[92182]_  = ~A233 & A232;
  assign \new_[92185]_  = A235 & A234;
  assign \new_[92186]_  = \new_[92185]_  & \new_[92182]_ ;
  assign \new_[92189]_  = ~A266 & A265;
  assign \new_[92192]_  = A268 & A267;
  assign \new_[92193]_  = \new_[92192]_  & \new_[92189]_ ;
  assign \new_[92194]_  = \new_[92193]_  & \new_[92186]_ ;
  assign \new_[92198]_  = A167 & A169;
  assign \new_[92199]_  = ~A170 & \new_[92198]_ ;
  assign \new_[92202]_  = ~A200 & A166;
  assign \new_[92205]_  = ~A203 & ~A202;
  assign \new_[92206]_  = \new_[92205]_  & \new_[92202]_ ;
  assign \new_[92207]_  = \new_[92206]_  & \new_[92199]_ ;
  assign \new_[92210]_  = ~A233 & A232;
  assign \new_[92213]_  = A235 & A234;
  assign \new_[92214]_  = \new_[92213]_  & \new_[92210]_ ;
  assign \new_[92217]_  = ~A266 & A265;
  assign \new_[92220]_  = A269 & A267;
  assign \new_[92221]_  = \new_[92220]_  & \new_[92217]_ ;
  assign \new_[92222]_  = \new_[92221]_  & \new_[92214]_ ;
  assign \new_[92226]_  = A167 & A169;
  assign \new_[92227]_  = ~A170 & \new_[92226]_ ;
  assign \new_[92230]_  = ~A200 & A166;
  assign \new_[92233]_  = ~A203 & ~A202;
  assign \new_[92234]_  = \new_[92233]_  & \new_[92230]_ ;
  assign \new_[92235]_  = \new_[92234]_  & \new_[92227]_ ;
  assign \new_[92238]_  = ~A233 & A232;
  assign \new_[92241]_  = A236 & A234;
  assign \new_[92242]_  = \new_[92241]_  & \new_[92238]_ ;
  assign \new_[92245]_  = ~A299 & A298;
  assign \new_[92248]_  = A301 & A300;
  assign \new_[92249]_  = \new_[92248]_  & \new_[92245]_ ;
  assign \new_[92250]_  = \new_[92249]_  & \new_[92242]_ ;
  assign \new_[92254]_  = A167 & A169;
  assign \new_[92255]_  = ~A170 & \new_[92254]_ ;
  assign \new_[92258]_  = ~A200 & A166;
  assign \new_[92261]_  = ~A203 & ~A202;
  assign \new_[92262]_  = \new_[92261]_  & \new_[92258]_ ;
  assign \new_[92263]_  = \new_[92262]_  & \new_[92255]_ ;
  assign \new_[92266]_  = ~A233 & A232;
  assign \new_[92269]_  = A236 & A234;
  assign \new_[92270]_  = \new_[92269]_  & \new_[92266]_ ;
  assign \new_[92273]_  = ~A299 & A298;
  assign \new_[92276]_  = A302 & A300;
  assign \new_[92277]_  = \new_[92276]_  & \new_[92273]_ ;
  assign \new_[92278]_  = \new_[92277]_  & \new_[92270]_ ;
  assign \new_[92282]_  = A167 & A169;
  assign \new_[92283]_  = ~A170 & \new_[92282]_ ;
  assign \new_[92286]_  = ~A200 & A166;
  assign \new_[92289]_  = ~A203 & ~A202;
  assign \new_[92290]_  = \new_[92289]_  & \new_[92286]_ ;
  assign \new_[92291]_  = \new_[92290]_  & \new_[92283]_ ;
  assign \new_[92294]_  = ~A233 & A232;
  assign \new_[92297]_  = A236 & A234;
  assign \new_[92298]_  = \new_[92297]_  & \new_[92294]_ ;
  assign \new_[92301]_  = ~A266 & A265;
  assign \new_[92304]_  = A268 & A267;
  assign \new_[92305]_  = \new_[92304]_  & \new_[92301]_ ;
  assign \new_[92306]_  = \new_[92305]_  & \new_[92298]_ ;
  assign \new_[92310]_  = A167 & A169;
  assign \new_[92311]_  = ~A170 & \new_[92310]_ ;
  assign \new_[92314]_  = ~A200 & A166;
  assign \new_[92317]_  = ~A203 & ~A202;
  assign \new_[92318]_  = \new_[92317]_  & \new_[92314]_ ;
  assign \new_[92319]_  = \new_[92318]_  & \new_[92311]_ ;
  assign \new_[92322]_  = ~A233 & A232;
  assign \new_[92325]_  = A236 & A234;
  assign \new_[92326]_  = \new_[92325]_  & \new_[92322]_ ;
  assign \new_[92329]_  = ~A266 & A265;
  assign \new_[92332]_  = A269 & A267;
  assign \new_[92333]_  = \new_[92332]_  & \new_[92329]_ ;
  assign \new_[92334]_  = \new_[92333]_  & \new_[92326]_ ;
  assign \new_[92338]_  = A167 & A169;
  assign \new_[92339]_  = ~A170 & \new_[92338]_ ;
  assign \new_[92342]_  = ~A200 & A166;
  assign \new_[92345]_  = ~A203 & ~A202;
  assign \new_[92346]_  = \new_[92345]_  & \new_[92342]_ ;
  assign \new_[92347]_  = \new_[92346]_  & \new_[92339]_ ;
  assign \new_[92350]_  = ~A233 & ~A232;
  assign \new_[92353]_  = ~A268 & ~A266;
  assign \new_[92354]_  = \new_[92353]_  & \new_[92350]_ ;
  assign \new_[92357]_  = A298 & ~A269;
  assign \new_[92360]_  = ~A302 & ~A301;
  assign \new_[92361]_  = \new_[92360]_  & \new_[92357]_ ;
  assign \new_[92362]_  = \new_[92361]_  & \new_[92354]_ ;
  assign \new_[92366]_  = A167 & A169;
  assign \new_[92367]_  = ~A170 & \new_[92366]_ ;
  assign \new_[92370]_  = ~A200 & A166;
  assign \new_[92373]_  = ~A233 & ~A201;
  assign \new_[92374]_  = \new_[92373]_  & \new_[92370]_ ;
  assign \new_[92375]_  = \new_[92374]_  & \new_[92367]_ ;
  assign \new_[92378]_  = ~A236 & ~A235;
  assign \new_[92381]_  = ~A268 & ~A266;
  assign \new_[92382]_  = \new_[92381]_  & \new_[92378]_ ;
  assign \new_[92385]_  = A298 & ~A269;
  assign \new_[92388]_  = ~A302 & ~A301;
  assign \new_[92389]_  = \new_[92388]_  & \new_[92385]_ ;
  assign \new_[92390]_  = \new_[92389]_  & \new_[92382]_ ;
  assign \new_[92394]_  = A167 & A169;
  assign \new_[92395]_  = ~A170 & \new_[92394]_ ;
  assign \new_[92398]_  = ~A199 & A166;
  assign \new_[92401]_  = ~A233 & ~A200;
  assign \new_[92402]_  = \new_[92401]_  & \new_[92398]_ ;
  assign \new_[92403]_  = \new_[92402]_  & \new_[92395]_ ;
  assign \new_[92406]_  = ~A236 & ~A235;
  assign \new_[92409]_  = ~A268 & ~A266;
  assign \new_[92410]_  = \new_[92409]_  & \new_[92406]_ ;
  assign \new_[92413]_  = A298 & ~A269;
  assign \new_[92416]_  = ~A302 & ~A301;
  assign \new_[92417]_  = \new_[92416]_  & \new_[92413]_ ;
  assign \new_[92418]_  = \new_[92417]_  & \new_[92410]_ ;
  assign \new_[92422]_  = ~A167 & A169;
  assign \new_[92423]_  = ~A170 & \new_[92422]_ ;
  assign \new_[92426]_  = A199 & ~A166;
  assign \new_[92429]_  = ~A233 & A200;
  assign \new_[92430]_  = \new_[92429]_  & \new_[92426]_ ;
  assign \new_[92431]_  = \new_[92430]_  & \new_[92423]_ ;
  assign \new_[92434]_  = ~A236 & ~A235;
  assign \new_[92437]_  = ~A268 & ~A266;
  assign \new_[92438]_  = \new_[92437]_  & \new_[92434]_ ;
  assign \new_[92441]_  = A298 & ~A269;
  assign \new_[92444]_  = ~A302 & ~A301;
  assign \new_[92445]_  = \new_[92444]_  & \new_[92441]_ ;
  assign \new_[92446]_  = \new_[92445]_  & \new_[92438]_ ;
  assign \new_[92450]_  = ~A167 & A169;
  assign \new_[92451]_  = ~A170 & \new_[92450]_ ;
  assign \new_[92454]_  = ~A200 & ~A166;
  assign \new_[92457]_  = ~A203 & ~A202;
  assign \new_[92458]_  = \new_[92457]_  & \new_[92454]_ ;
  assign \new_[92459]_  = \new_[92458]_  & \new_[92451]_ ;
  assign \new_[92462]_  = A233 & A232;
  assign \new_[92465]_  = ~A268 & A265;
  assign \new_[92466]_  = \new_[92465]_  & \new_[92462]_ ;
  assign \new_[92469]_  = ~A299 & ~A269;
  assign \new_[92472]_  = ~A302 & ~A301;
  assign \new_[92473]_  = \new_[92472]_  & \new_[92469]_ ;
  assign \new_[92474]_  = \new_[92473]_  & \new_[92466]_ ;
  assign \new_[92478]_  = ~A167 & A169;
  assign \new_[92479]_  = ~A170 & \new_[92478]_ ;
  assign \new_[92482]_  = ~A200 & ~A166;
  assign \new_[92485]_  = ~A203 & ~A202;
  assign \new_[92486]_  = \new_[92485]_  & \new_[92482]_ ;
  assign \new_[92487]_  = \new_[92486]_  & \new_[92479]_ ;
  assign \new_[92490]_  = ~A235 & ~A233;
  assign \new_[92493]_  = A265 & ~A236;
  assign \new_[92494]_  = \new_[92493]_  & \new_[92490]_ ;
  assign \new_[92497]_  = A298 & A266;
  assign \new_[92500]_  = ~A302 & ~A301;
  assign \new_[92501]_  = \new_[92500]_  & \new_[92497]_ ;
  assign \new_[92502]_  = \new_[92501]_  & \new_[92494]_ ;
  assign \new_[92506]_  = ~A167 & A169;
  assign \new_[92507]_  = ~A170 & \new_[92506]_ ;
  assign \new_[92510]_  = ~A200 & ~A166;
  assign \new_[92513]_  = ~A203 & ~A202;
  assign \new_[92514]_  = \new_[92513]_  & \new_[92510]_ ;
  assign \new_[92515]_  = \new_[92514]_  & \new_[92507]_ ;
  assign \new_[92518]_  = ~A235 & ~A233;
  assign \new_[92521]_  = ~A266 & ~A236;
  assign \new_[92522]_  = \new_[92521]_  & \new_[92518]_ ;
  assign \new_[92525]_  = ~A269 & ~A268;
  assign \new_[92528]_  = ~A300 & A298;
  assign \new_[92529]_  = \new_[92528]_  & \new_[92525]_ ;
  assign \new_[92530]_  = \new_[92529]_  & \new_[92522]_ ;
  assign \new_[92534]_  = ~A167 & A169;
  assign \new_[92535]_  = ~A170 & \new_[92534]_ ;
  assign \new_[92538]_  = ~A200 & ~A166;
  assign \new_[92541]_  = ~A203 & ~A202;
  assign \new_[92542]_  = \new_[92541]_  & \new_[92538]_ ;
  assign \new_[92543]_  = \new_[92542]_  & \new_[92535]_ ;
  assign \new_[92546]_  = ~A235 & ~A233;
  assign \new_[92549]_  = ~A266 & ~A236;
  assign \new_[92550]_  = \new_[92549]_  & \new_[92546]_ ;
  assign \new_[92553]_  = ~A269 & ~A268;
  assign \new_[92556]_  = A299 & A298;
  assign \new_[92557]_  = \new_[92556]_  & \new_[92553]_ ;
  assign \new_[92558]_  = \new_[92557]_  & \new_[92550]_ ;
  assign \new_[92562]_  = ~A167 & A169;
  assign \new_[92563]_  = ~A170 & \new_[92562]_ ;
  assign \new_[92566]_  = ~A200 & ~A166;
  assign \new_[92569]_  = ~A203 & ~A202;
  assign \new_[92570]_  = \new_[92569]_  & \new_[92566]_ ;
  assign \new_[92571]_  = \new_[92570]_  & \new_[92563]_ ;
  assign \new_[92574]_  = ~A235 & ~A233;
  assign \new_[92577]_  = ~A266 & ~A236;
  assign \new_[92578]_  = \new_[92577]_  & \new_[92574]_ ;
  assign \new_[92581]_  = ~A269 & ~A268;
  assign \new_[92584]_  = ~A299 & ~A298;
  assign \new_[92585]_  = \new_[92584]_  & \new_[92581]_ ;
  assign \new_[92586]_  = \new_[92585]_  & \new_[92578]_ ;
  assign \new_[92590]_  = ~A167 & A169;
  assign \new_[92591]_  = ~A170 & \new_[92590]_ ;
  assign \new_[92594]_  = ~A200 & ~A166;
  assign \new_[92597]_  = ~A203 & ~A202;
  assign \new_[92598]_  = \new_[92597]_  & \new_[92594]_ ;
  assign \new_[92599]_  = \new_[92598]_  & \new_[92591]_ ;
  assign \new_[92602]_  = ~A235 & ~A233;
  assign \new_[92605]_  = ~A266 & ~A236;
  assign \new_[92606]_  = \new_[92605]_  & \new_[92602]_ ;
  assign \new_[92609]_  = A298 & ~A267;
  assign \new_[92612]_  = ~A302 & ~A301;
  assign \new_[92613]_  = \new_[92612]_  & \new_[92609]_ ;
  assign \new_[92614]_  = \new_[92613]_  & \new_[92606]_ ;
  assign \new_[92618]_  = ~A167 & A169;
  assign \new_[92619]_  = ~A170 & \new_[92618]_ ;
  assign \new_[92622]_  = ~A200 & ~A166;
  assign \new_[92625]_  = ~A203 & ~A202;
  assign \new_[92626]_  = \new_[92625]_  & \new_[92622]_ ;
  assign \new_[92627]_  = \new_[92626]_  & \new_[92619]_ ;
  assign \new_[92630]_  = ~A235 & ~A233;
  assign \new_[92633]_  = ~A265 & ~A236;
  assign \new_[92634]_  = \new_[92633]_  & \new_[92630]_ ;
  assign \new_[92637]_  = A298 & ~A266;
  assign \new_[92640]_  = ~A302 & ~A301;
  assign \new_[92641]_  = \new_[92640]_  & \new_[92637]_ ;
  assign \new_[92642]_  = \new_[92641]_  & \new_[92634]_ ;
  assign \new_[92646]_  = ~A167 & A169;
  assign \new_[92647]_  = ~A170 & \new_[92646]_ ;
  assign \new_[92650]_  = ~A200 & ~A166;
  assign \new_[92653]_  = ~A203 & ~A202;
  assign \new_[92654]_  = \new_[92653]_  & \new_[92650]_ ;
  assign \new_[92655]_  = \new_[92654]_  & \new_[92647]_ ;
  assign \new_[92658]_  = ~A234 & ~A233;
  assign \new_[92661]_  = ~A268 & ~A266;
  assign \new_[92662]_  = \new_[92661]_  & \new_[92658]_ ;
  assign \new_[92665]_  = A298 & ~A269;
  assign \new_[92668]_  = ~A302 & ~A301;
  assign \new_[92669]_  = \new_[92668]_  & \new_[92665]_ ;
  assign \new_[92670]_  = \new_[92669]_  & \new_[92662]_ ;
  assign \new_[92674]_  = ~A167 & A169;
  assign \new_[92675]_  = ~A170 & \new_[92674]_ ;
  assign \new_[92678]_  = ~A200 & ~A166;
  assign \new_[92681]_  = ~A203 & ~A202;
  assign \new_[92682]_  = \new_[92681]_  & \new_[92678]_ ;
  assign \new_[92683]_  = \new_[92682]_  & \new_[92675]_ ;
  assign \new_[92686]_  = ~A233 & A232;
  assign \new_[92689]_  = A235 & A234;
  assign \new_[92690]_  = \new_[92689]_  & \new_[92686]_ ;
  assign \new_[92693]_  = ~A299 & A298;
  assign \new_[92696]_  = A301 & A300;
  assign \new_[92697]_  = \new_[92696]_  & \new_[92693]_ ;
  assign \new_[92698]_  = \new_[92697]_  & \new_[92690]_ ;
  assign \new_[92702]_  = ~A167 & A169;
  assign \new_[92703]_  = ~A170 & \new_[92702]_ ;
  assign \new_[92706]_  = ~A200 & ~A166;
  assign \new_[92709]_  = ~A203 & ~A202;
  assign \new_[92710]_  = \new_[92709]_  & \new_[92706]_ ;
  assign \new_[92711]_  = \new_[92710]_  & \new_[92703]_ ;
  assign \new_[92714]_  = ~A233 & A232;
  assign \new_[92717]_  = A235 & A234;
  assign \new_[92718]_  = \new_[92717]_  & \new_[92714]_ ;
  assign \new_[92721]_  = ~A299 & A298;
  assign \new_[92724]_  = A302 & A300;
  assign \new_[92725]_  = \new_[92724]_  & \new_[92721]_ ;
  assign \new_[92726]_  = \new_[92725]_  & \new_[92718]_ ;
  assign \new_[92730]_  = ~A167 & A169;
  assign \new_[92731]_  = ~A170 & \new_[92730]_ ;
  assign \new_[92734]_  = ~A200 & ~A166;
  assign \new_[92737]_  = ~A203 & ~A202;
  assign \new_[92738]_  = \new_[92737]_  & \new_[92734]_ ;
  assign \new_[92739]_  = \new_[92738]_  & \new_[92731]_ ;
  assign \new_[92742]_  = ~A233 & A232;
  assign \new_[92745]_  = A235 & A234;
  assign \new_[92746]_  = \new_[92745]_  & \new_[92742]_ ;
  assign \new_[92749]_  = ~A266 & A265;
  assign \new_[92752]_  = A268 & A267;
  assign \new_[92753]_  = \new_[92752]_  & \new_[92749]_ ;
  assign \new_[92754]_  = \new_[92753]_  & \new_[92746]_ ;
  assign \new_[92758]_  = ~A167 & A169;
  assign \new_[92759]_  = ~A170 & \new_[92758]_ ;
  assign \new_[92762]_  = ~A200 & ~A166;
  assign \new_[92765]_  = ~A203 & ~A202;
  assign \new_[92766]_  = \new_[92765]_  & \new_[92762]_ ;
  assign \new_[92767]_  = \new_[92766]_  & \new_[92759]_ ;
  assign \new_[92770]_  = ~A233 & A232;
  assign \new_[92773]_  = A235 & A234;
  assign \new_[92774]_  = \new_[92773]_  & \new_[92770]_ ;
  assign \new_[92777]_  = ~A266 & A265;
  assign \new_[92780]_  = A269 & A267;
  assign \new_[92781]_  = \new_[92780]_  & \new_[92777]_ ;
  assign \new_[92782]_  = \new_[92781]_  & \new_[92774]_ ;
  assign \new_[92786]_  = ~A167 & A169;
  assign \new_[92787]_  = ~A170 & \new_[92786]_ ;
  assign \new_[92790]_  = ~A200 & ~A166;
  assign \new_[92793]_  = ~A203 & ~A202;
  assign \new_[92794]_  = \new_[92793]_  & \new_[92790]_ ;
  assign \new_[92795]_  = \new_[92794]_  & \new_[92787]_ ;
  assign \new_[92798]_  = ~A233 & A232;
  assign \new_[92801]_  = A236 & A234;
  assign \new_[92802]_  = \new_[92801]_  & \new_[92798]_ ;
  assign \new_[92805]_  = ~A299 & A298;
  assign \new_[92808]_  = A301 & A300;
  assign \new_[92809]_  = \new_[92808]_  & \new_[92805]_ ;
  assign \new_[92810]_  = \new_[92809]_  & \new_[92802]_ ;
  assign \new_[92814]_  = ~A167 & A169;
  assign \new_[92815]_  = ~A170 & \new_[92814]_ ;
  assign \new_[92818]_  = ~A200 & ~A166;
  assign \new_[92821]_  = ~A203 & ~A202;
  assign \new_[92822]_  = \new_[92821]_  & \new_[92818]_ ;
  assign \new_[92823]_  = \new_[92822]_  & \new_[92815]_ ;
  assign \new_[92826]_  = ~A233 & A232;
  assign \new_[92829]_  = A236 & A234;
  assign \new_[92830]_  = \new_[92829]_  & \new_[92826]_ ;
  assign \new_[92833]_  = ~A299 & A298;
  assign \new_[92836]_  = A302 & A300;
  assign \new_[92837]_  = \new_[92836]_  & \new_[92833]_ ;
  assign \new_[92838]_  = \new_[92837]_  & \new_[92830]_ ;
  assign \new_[92842]_  = ~A167 & A169;
  assign \new_[92843]_  = ~A170 & \new_[92842]_ ;
  assign \new_[92846]_  = ~A200 & ~A166;
  assign \new_[92849]_  = ~A203 & ~A202;
  assign \new_[92850]_  = \new_[92849]_  & \new_[92846]_ ;
  assign \new_[92851]_  = \new_[92850]_  & \new_[92843]_ ;
  assign \new_[92854]_  = ~A233 & A232;
  assign \new_[92857]_  = A236 & A234;
  assign \new_[92858]_  = \new_[92857]_  & \new_[92854]_ ;
  assign \new_[92861]_  = ~A266 & A265;
  assign \new_[92864]_  = A268 & A267;
  assign \new_[92865]_  = \new_[92864]_  & \new_[92861]_ ;
  assign \new_[92866]_  = \new_[92865]_  & \new_[92858]_ ;
  assign \new_[92870]_  = ~A167 & A169;
  assign \new_[92871]_  = ~A170 & \new_[92870]_ ;
  assign \new_[92874]_  = ~A200 & ~A166;
  assign \new_[92877]_  = ~A203 & ~A202;
  assign \new_[92878]_  = \new_[92877]_  & \new_[92874]_ ;
  assign \new_[92879]_  = \new_[92878]_  & \new_[92871]_ ;
  assign \new_[92882]_  = ~A233 & A232;
  assign \new_[92885]_  = A236 & A234;
  assign \new_[92886]_  = \new_[92885]_  & \new_[92882]_ ;
  assign \new_[92889]_  = ~A266 & A265;
  assign \new_[92892]_  = A269 & A267;
  assign \new_[92893]_  = \new_[92892]_  & \new_[92889]_ ;
  assign \new_[92894]_  = \new_[92893]_  & \new_[92886]_ ;
  assign \new_[92898]_  = ~A167 & A169;
  assign \new_[92899]_  = ~A170 & \new_[92898]_ ;
  assign \new_[92902]_  = ~A200 & ~A166;
  assign \new_[92905]_  = ~A203 & ~A202;
  assign \new_[92906]_  = \new_[92905]_  & \new_[92902]_ ;
  assign \new_[92907]_  = \new_[92906]_  & \new_[92899]_ ;
  assign \new_[92910]_  = ~A233 & ~A232;
  assign \new_[92913]_  = ~A268 & ~A266;
  assign \new_[92914]_  = \new_[92913]_  & \new_[92910]_ ;
  assign \new_[92917]_  = A298 & ~A269;
  assign \new_[92920]_  = ~A302 & ~A301;
  assign \new_[92921]_  = \new_[92920]_  & \new_[92917]_ ;
  assign \new_[92922]_  = \new_[92921]_  & \new_[92914]_ ;
  assign \new_[92926]_  = ~A167 & A169;
  assign \new_[92927]_  = ~A170 & \new_[92926]_ ;
  assign \new_[92930]_  = ~A200 & ~A166;
  assign \new_[92933]_  = ~A233 & ~A201;
  assign \new_[92934]_  = \new_[92933]_  & \new_[92930]_ ;
  assign \new_[92935]_  = \new_[92934]_  & \new_[92927]_ ;
  assign \new_[92938]_  = ~A236 & ~A235;
  assign \new_[92941]_  = ~A268 & ~A266;
  assign \new_[92942]_  = \new_[92941]_  & \new_[92938]_ ;
  assign \new_[92945]_  = A298 & ~A269;
  assign \new_[92948]_  = ~A302 & ~A301;
  assign \new_[92949]_  = \new_[92948]_  & \new_[92945]_ ;
  assign \new_[92950]_  = \new_[92949]_  & \new_[92942]_ ;
  assign \new_[92954]_  = ~A167 & A169;
  assign \new_[92955]_  = ~A170 & \new_[92954]_ ;
  assign \new_[92958]_  = ~A199 & ~A166;
  assign \new_[92961]_  = ~A233 & ~A200;
  assign \new_[92962]_  = \new_[92961]_  & \new_[92958]_ ;
  assign \new_[92963]_  = \new_[92962]_  & \new_[92955]_ ;
  assign \new_[92966]_  = ~A236 & ~A235;
  assign \new_[92969]_  = ~A268 & ~A266;
  assign \new_[92970]_  = \new_[92969]_  & \new_[92966]_ ;
  assign \new_[92973]_  = A298 & ~A269;
  assign \new_[92976]_  = ~A302 & ~A301;
  assign \new_[92977]_  = \new_[92976]_  & \new_[92973]_ ;
  assign \new_[92978]_  = \new_[92977]_  & \new_[92970]_ ;
  assign \new_[92982]_  = ~A166 & ~A167;
  assign \new_[92983]_  = ~A169 & \new_[92982]_ ;
  assign \new_[92986]_  = ~A200 & A199;
  assign \new_[92989]_  = A202 & A201;
  assign \new_[92990]_  = \new_[92989]_  & \new_[92986]_ ;
  assign \new_[92991]_  = \new_[92990]_  & \new_[92983]_ ;
  assign \new_[92994]_  = A233 & A232;
  assign \new_[92997]_  = ~A268 & A265;
  assign \new_[92998]_  = \new_[92997]_  & \new_[92994]_ ;
  assign \new_[93001]_  = ~A299 & ~A269;
  assign \new_[93004]_  = ~A302 & ~A301;
  assign \new_[93005]_  = \new_[93004]_  & \new_[93001]_ ;
  assign \new_[93006]_  = \new_[93005]_  & \new_[92998]_ ;
  assign \new_[93010]_  = ~A166 & ~A167;
  assign \new_[93011]_  = ~A169 & \new_[93010]_ ;
  assign \new_[93014]_  = ~A200 & A199;
  assign \new_[93017]_  = A202 & A201;
  assign \new_[93018]_  = \new_[93017]_  & \new_[93014]_ ;
  assign \new_[93019]_  = \new_[93018]_  & \new_[93011]_ ;
  assign \new_[93022]_  = ~A235 & ~A233;
  assign \new_[93025]_  = A265 & ~A236;
  assign \new_[93026]_  = \new_[93025]_  & \new_[93022]_ ;
  assign \new_[93029]_  = A298 & A266;
  assign \new_[93032]_  = ~A302 & ~A301;
  assign \new_[93033]_  = \new_[93032]_  & \new_[93029]_ ;
  assign \new_[93034]_  = \new_[93033]_  & \new_[93026]_ ;
  assign \new_[93038]_  = ~A166 & ~A167;
  assign \new_[93039]_  = ~A169 & \new_[93038]_ ;
  assign \new_[93042]_  = ~A200 & A199;
  assign \new_[93045]_  = A202 & A201;
  assign \new_[93046]_  = \new_[93045]_  & \new_[93042]_ ;
  assign \new_[93047]_  = \new_[93046]_  & \new_[93039]_ ;
  assign \new_[93050]_  = ~A235 & ~A233;
  assign \new_[93053]_  = ~A266 & ~A236;
  assign \new_[93054]_  = \new_[93053]_  & \new_[93050]_ ;
  assign \new_[93057]_  = ~A269 & ~A268;
  assign \new_[93060]_  = ~A300 & A298;
  assign \new_[93061]_  = \new_[93060]_  & \new_[93057]_ ;
  assign \new_[93062]_  = \new_[93061]_  & \new_[93054]_ ;
  assign \new_[93066]_  = ~A166 & ~A167;
  assign \new_[93067]_  = ~A169 & \new_[93066]_ ;
  assign \new_[93070]_  = ~A200 & A199;
  assign \new_[93073]_  = A202 & A201;
  assign \new_[93074]_  = \new_[93073]_  & \new_[93070]_ ;
  assign \new_[93075]_  = \new_[93074]_  & \new_[93067]_ ;
  assign \new_[93078]_  = ~A235 & ~A233;
  assign \new_[93081]_  = ~A266 & ~A236;
  assign \new_[93082]_  = \new_[93081]_  & \new_[93078]_ ;
  assign \new_[93085]_  = ~A269 & ~A268;
  assign \new_[93088]_  = A299 & A298;
  assign \new_[93089]_  = \new_[93088]_  & \new_[93085]_ ;
  assign \new_[93090]_  = \new_[93089]_  & \new_[93082]_ ;
  assign \new_[93094]_  = ~A166 & ~A167;
  assign \new_[93095]_  = ~A169 & \new_[93094]_ ;
  assign \new_[93098]_  = ~A200 & A199;
  assign \new_[93101]_  = A202 & A201;
  assign \new_[93102]_  = \new_[93101]_  & \new_[93098]_ ;
  assign \new_[93103]_  = \new_[93102]_  & \new_[93095]_ ;
  assign \new_[93106]_  = ~A235 & ~A233;
  assign \new_[93109]_  = ~A266 & ~A236;
  assign \new_[93110]_  = \new_[93109]_  & \new_[93106]_ ;
  assign \new_[93113]_  = ~A269 & ~A268;
  assign \new_[93116]_  = ~A299 & ~A298;
  assign \new_[93117]_  = \new_[93116]_  & \new_[93113]_ ;
  assign \new_[93118]_  = \new_[93117]_  & \new_[93110]_ ;
  assign \new_[93122]_  = ~A166 & ~A167;
  assign \new_[93123]_  = ~A169 & \new_[93122]_ ;
  assign \new_[93126]_  = ~A200 & A199;
  assign \new_[93129]_  = A202 & A201;
  assign \new_[93130]_  = \new_[93129]_  & \new_[93126]_ ;
  assign \new_[93131]_  = \new_[93130]_  & \new_[93123]_ ;
  assign \new_[93134]_  = ~A235 & ~A233;
  assign \new_[93137]_  = ~A266 & ~A236;
  assign \new_[93138]_  = \new_[93137]_  & \new_[93134]_ ;
  assign \new_[93141]_  = A298 & ~A267;
  assign \new_[93144]_  = ~A302 & ~A301;
  assign \new_[93145]_  = \new_[93144]_  & \new_[93141]_ ;
  assign \new_[93146]_  = \new_[93145]_  & \new_[93138]_ ;
  assign \new_[93150]_  = ~A166 & ~A167;
  assign \new_[93151]_  = ~A169 & \new_[93150]_ ;
  assign \new_[93154]_  = ~A200 & A199;
  assign \new_[93157]_  = A202 & A201;
  assign \new_[93158]_  = \new_[93157]_  & \new_[93154]_ ;
  assign \new_[93159]_  = \new_[93158]_  & \new_[93151]_ ;
  assign \new_[93162]_  = ~A235 & ~A233;
  assign \new_[93165]_  = ~A265 & ~A236;
  assign \new_[93166]_  = \new_[93165]_  & \new_[93162]_ ;
  assign \new_[93169]_  = A298 & ~A266;
  assign \new_[93172]_  = ~A302 & ~A301;
  assign \new_[93173]_  = \new_[93172]_  & \new_[93169]_ ;
  assign \new_[93174]_  = \new_[93173]_  & \new_[93166]_ ;
  assign \new_[93178]_  = ~A166 & ~A167;
  assign \new_[93179]_  = ~A169 & \new_[93178]_ ;
  assign \new_[93182]_  = ~A200 & A199;
  assign \new_[93185]_  = A202 & A201;
  assign \new_[93186]_  = \new_[93185]_  & \new_[93182]_ ;
  assign \new_[93187]_  = \new_[93186]_  & \new_[93179]_ ;
  assign \new_[93190]_  = ~A234 & ~A233;
  assign \new_[93193]_  = ~A268 & ~A266;
  assign \new_[93194]_  = \new_[93193]_  & \new_[93190]_ ;
  assign \new_[93197]_  = A298 & ~A269;
  assign \new_[93200]_  = ~A302 & ~A301;
  assign \new_[93201]_  = \new_[93200]_  & \new_[93197]_ ;
  assign \new_[93202]_  = \new_[93201]_  & \new_[93194]_ ;
  assign \new_[93206]_  = ~A166 & ~A167;
  assign \new_[93207]_  = ~A169 & \new_[93206]_ ;
  assign \new_[93210]_  = ~A200 & A199;
  assign \new_[93213]_  = A202 & A201;
  assign \new_[93214]_  = \new_[93213]_  & \new_[93210]_ ;
  assign \new_[93215]_  = \new_[93214]_  & \new_[93207]_ ;
  assign \new_[93218]_  = ~A233 & A232;
  assign \new_[93221]_  = A235 & A234;
  assign \new_[93222]_  = \new_[93221]_  & \new_[93218]_ ;
  assign \new_[93225]_  = ~A299 & A298;
  assign \new_[93228]_  = A301 & A300;
  assign \new_[93229]_  = \new_[93228]_  & \new_[93225]_ ;
  assign \new_[93230]_  = \new_[93229]_  & \new_[93222]_ ;
  assign \new_[93234]_  = ~A166 & ~A167;
  assign \new_[93235]_  = ~A169 & \new_[93234]_ ;
  assign \new_[93238]_  = ~A200 & A199;
  assign \new_[93241]_  = A202 & A201;
  assign \new_[93242]_  = \new_[93241]_  & \new_[93238]_ ;
  assign \new_[93243]_  = \new_[93242]_  & \new_[93235]_ ;
  assign \new_[93246]_  = ~A233 & A232;
  assign \new_[93249]_  = A235 & A234;
  assign \new_[93250]_  = \new_[93249]_  & \new_[93246]_ ;
  assign \new_[93253]_  = ~A299 & A298;
  assign \new_[93256]_  = A302 & A300;
  assign \new_[93257]_  = \new_[93256]_  & \new_[93253]_ ;
  assign \new_[93258]_  = \new_[93257]_  & \new_[93250]_ ;
  assign \new_[93262]_  = ~A166 & ~A167;
  assign \new_[93263]_  = ~A169 & \new_[93262]_ ;
  assign \new_[93266]_  = ~A200 & A199;
  assign \new_[93269]_  = A202 & A201;
  assign \new_[93270]_  = \new_[93269]_  & \new_[93266]_ ;
  assign \new_[93271]_  = \new_[93270]_  & \new_[93263]_ ;
  assign \new_[93274]_  = ~A233 & A232;
  assign \new_[93277]_  = A235 & A234;
  assign \new_[93278]_  = \new_[93277]_  & \new_[93274]_ ;
  assign \new_[93281]_  = ~A266 & A265;
  assign \new_[93284]_  = A268 & A267;
  assign \new_[93285]_  = \new_[93284]_  & \new_[93281]_ ;
  assign \new_[93286]_  = \new_[93285]_  & \new_[93278]_ ;
  assign \new_[93290]_  = ~A166 & ~A167;
  assign \new_[93291]_  = ~A169 & \new_[93290]_ ;
  assign \new_[93294]_  = ~A200 & A199;
  assign \new_[93297]_  = A202 & A201;
  assign \new_[93298]_  = \new_[93297]_  & \new_[93294]_ ;
  assign \new_[93299]_  = \new_[93298]_  & \new_[93291]_ ;
  assign \new_[93302]_  = ~A233 & A232;
  assign \new_[93305]_  = A235 & A234;
  assign \new_[93306]_  = \new_[93305]_  & \new_[93302]_ ;
  assign \new_[93309]_  = ~A266 & A265;
  assign \new_[93312]_  = A269 & A267;
  assign \new_[93313]_  = \new_[93312]_  & \new_[93309]_ ;
  assign \new_[93314]_  = \new_[93313]_  & \new_[93306]_ ;
  assign \new_[93318]_  = ~A166 & ~A167;
  assign \new_[93319]_  = ~A169 & \new_[93318]_ ;
  assign \new_[93322]_  = ~A200 & A199;
  assign \new_[93325]_  = A202 & A201;
  assign \new_[93326]_  = \new_[93325]_  & \new_[93322]_ ;
  assign \new_[93327]_  = \new_[93326]_  & \new_[93319]_ ;
  assign \new_[93330]_  = ~A233 & A232;
  assign \new_[93333]_  = A236 & A234;
  assign \new_[93334]_  = \new_[93333]_  & \new_[93330]_ ;
  assign \new_[93337]_  = ~A299 & A298;
  assign \new_[93340]_  = A301 & A300;
  assign \new_[93341]_  = \new_[93340]_  & \new_[93337]_ ;
  assign \new_[93342]_  = \new_[93341]_  & \new_[93334]_ ;
  assign \new_[93346]_  = ~A166 & ~A167;
  assign \new_[93347]_  = ~A169 & \new_[93346]_ ;
  assign \new_[93350]_  = ~A200 & A199;
  assign \new_[93353]_  = A202 & A201;
  assign \new_[93354]_  = \new_[93353]_  & \new_[93350]_ ;
  assign \new_[93355]_  = \new_[93354]_  & \new_[93347]_ ;
  assign \new_[93358]_  = ~A233 & A232;
  assign \new_[93361]_  = A236 & A234;
  assign \new_[93362]_  = \new_[93361]_  & \new_[93358]_ ;
  assign \new_[93365]_  = ~A299 & A298;
  assign \new_[93368]_  = A302 & A300;
  assign \new_[93369]_  = \new_[93368]_  & \new_[93365]_ ;
  assign \new_[93370]_  = \new_[93369]_  & \new_[93362]_ ;
  assign \new_[93374]_  = ~A166 & ~A167;
  assign \new_[93375]_  = ~A169 & \new_[93374]_ ;
  assign \new_[93378]_  = ~A200 & A199;
  assign \new_[93381]_  = A202 & A201;
  assign \new_[93382]_  = \new_[93381]_  & \new_[93378]_ ;
  assign \new_[93383]_  = \new_[93382]_  & \new_[93375]_ ;
  assign \new_[93386]_  = ~A233 & A232;
  assign \new_[93389]_  = A236 & A234;
  assign \new_[93390]_  = \new_[93389]_  & \new_[93386]_ ;
  assign \new_[93393]_  = ~A266 & A265;
  assign \new_[93396]_  = A268 & A267;
  assign \new_[93397]_  = \new_[93396]_  & \new_[93393]_ ;
  assign \new_[93398]_  = \new_[93397]_  & \new_[93390]_ ;
  assign \new_[93402]_  = ~A166 & ~A167;
  assign \new_[93403]_  = ~A169 & \new_[93402]_ ;
  assign \new_[93406]_  = ~A200 & A199;
  assign \new_[93409]_  = A202 & A201;
  assign \new_[93410]_  = \new_[93409]_  & \new_[93406]_ ;
  assign \new_[93411]_  = \new_[93410]_  & \new_[93403]_ ;
  assign \new_[93414]_  = ~A233 & A232;
  assign \new_[93417]_  = A236 & A234;
  assign \new_[93418]_  = \new_[93417]_  & \new_[93414]_ ;
  assign \new_[93421]_  = ~A266 & A265;
  assign \new_[93424]_  = A269 & A267;
  assign \new_[93425]_  = \new_[93424]_  & \new_[93421]_ ;
  assign \new_[93426]_  = \new_[93425]_  & \new_[93418]_ ;
  assign \new_[93430]_  = ~A166 & ~A167;
  assign \new_[93431]_  = ~A169 & \new_[93430]_ ;
  assign \new_[93434]_  = ~A200 & A199;
  assign \new_[93437]_  = A202 & A201;
  assign \new_[93438]_  = \new_[93437]_  & \new_[93434]_ ;
  assign \new_[93439]_  = \new_[93438]_  & \new_[93431]_ ;
  assign \new_[93442]_  = ~A233 & ~A232;
  assign \new_[93445]_  = ~A268 & ~A266;
  assign \new_[93446]_  = \new_[93445]_  & \new_[93442]_ ;
  assign \new_[93449]_  = A298 & ~A269;
  assign \new_[93452]_  = ~A302 & ~A301;
  assign \new_[93453]_  = \new_[93452]_  & \new_[93449]_ ;
  assign \new_[93454]_  = \new_[93453]_  & \new_[93446]_ ;
  assign \new_[93458]_  = ~A166 & ~A167;
  assign \new_[93459]_  = ~A169 & \new_[93458]_ ;
  assign \new_[93462]_  = ~A200 & A199;
  assign \new_[93465]_  = A203 & A201;
  assign \new_[93466]_  = \new_[93465]_  & \new_[93462]_ ;
  assign \new_[93467]_  = \new_[93466]_  & \new_[93459]_ ;
  assign \new_[93470]_  = A233 & A232;
  assign \new_[93473]_  = ~A268 & A265;
  assign \new_[93474]_  = \new_[93473]_  & \new_[93470]_ ;
  assign \new_[93477]_  = ~A299 & ~A269;
  assign \new_[93480]_  = ~A302 & ~A301;
  assign \new_[93481]_  = \new_[93480]_  & \new_[93477]_ ;
  assign \new_[93482]_  = \new_[93481]_  & \new_[93474]_ ;
  assign \new_[93486]_  = ~A166 & ~A167;
  assign \new_[93487]_  = ~A169 & \new_[93486]_ ;
  assign \new_[93490]_  = ~A200 & A199;
  assign \new_[93493]_  = A203 & A201;
  assign \new_[93494]_  = \new_[93493]_  & \new_[93490]_ ;
  assign \new_[93495]_  = \new_[93494]_  & \new_[93487]_ ;
  assign \new_[93498]_  = ~A235 & ~A233;
  assign \new_[93501]_  = A265 & ~A236;
  assign \new_[93502]_  = \new_[93501]_  & \new_[93498]_ ;
  assign \new_[93505]_  = A298 & A266;
  assign \new_[93508]_  = ~A302 & ~A301;
  assign \new_[93509]_  = \new_[93508]_  & \new_[93505]_ ;
  assign \new_[93510]_  = \new_[93509]_  & \new_[93502]_ ;
  assign \new_[93514]_  = ~A166 & ~A167;
  assign \new_[93515]_  = ~A169 & \new_[93514]_ ;
  assign \new_[93518]_  = ~A200 & A199;
  assign \new_[93521]_  = A203 & A201;
  assign \new_[93522]_  = \new_[93521]_  & \new_[93518]_ ;
  assign \new_[93523]_  = \new_[93522]_  & \new_[93515]_ ;
  assign \new_[93526]_  = ~A235 & ~A233;
  assign \new_[93529]_  = ~A266 & ~A236;
  assign \new_[93530]_  = \new_[93529]_  & \new_[93526]_ ;
  assign \new_[93533]_  = ~A269 & ~A268;
  assign \new_[93536]_  = ~A300 & A298;
  assign \new_[93537]_  = \new_[93536]_  & \new_[93533]_ ;
  assign \new_[93538]_  = \new_[93537]_  & \new_[93530]_ ;
  assign \new_[93542]_  = ~A166 & ~A167;
  assign \new_[93543]_  = ~A169 & \new_[93542]_ ;
  assign \new_[93546]_  = ~A200 & A199;
  assign \new_[93549]_  = A203 & A201;
  assign \new_[93550]_  = \new_[93549]_  & \new_[93546]_ ;
  assign \new_[93551]_  = \new_[93550]_  & \new_[93543]_ ;
  assign \new_[93554]_  = ~A235 & ~A233;
  assign \new_[93557]_  = ~A266 & ~A236;
  assign \new_[93558]_  = \new_[93557]_  & \new_[93554]_ ;
  assign \new_[93561]_  = ~A269 & ~A268;
  assign \new_[93564]_  = A299 & A298;
  assign \new_[93565]_  = \new_[93564]_  & \new_[93561]_ ;
  assign \new_[93566]_  = \new_[93565]_  & \new_[93558]_ ;
  assign \new_[93570]_  = ~A166 & ~A167;
  assign \new_[93571]_  = ~A169 & \new_[93570]_ ;
  assign \new_[93574]_  = ~A200 & A199;
  assign \new_[93577]_  = A203 & A201;
  assign \new_[93578]_  = \new_[93577]_  & \new_[93574]_ ;
  assign \new_[93579]_  = \new_[93578]_  & \new_[93571]_ ;
  assign \new_[93582]_  = ~A235 & ~A233;
  assign \new_[93585]_  = ~A266 & ~A236;
  assign \new_[93586]_  = \new_[93585]_  & \new_[93582]_ ;
  assign \new_[93589]_  = ~A269 & ~A268;
  assign \new_[93592]_  = ~A299 & ~A298;
  assign \new_[93593]_  = \new_[93592]_  & \new_[93589]_ ;
  assign \new_[93594]_  = \new_[93593]_  & \new_[93586]_ ;
  assign \new_[93598]_  = ~A166 & ~A167;
  assign \new_[93599]_  = ~A169 & \new_[93598]_ ;
  assign \new_[93602]_  = ~A200 & A199;
  assign \new_[93605]_  = A203 & A201;
  assign \new_[93606]_  = \new_[93605]_  & \new_[93602]_ ;
  assign \new_[93607]_  = \new_[93606]_  & \new_[93599]_ ;
  assign \new_[93610]_  = ~A235 & ~A233;
  assign \new_[93613]_  = ~A266 & ~A236;
  assign \new_[93614]_  = \new_[93613]_  & \new_[93610]_ ;
  assign \new_[93617]_  = A298 & ~A267;
  assign \new_[93620]_  = ~A302 & ~A301;
  assign \new_[93621]_  = \new_[93620]_  & \new_[93617]_ ;
  assign \new_[93622]_  = \new_[93621]_  & \new_[93614]_ ;
  assign \new_[93626]_  = ~A166 & ~A167;
  assign \new_[93627]_  = ~A169 & \new_[93626]_ ;
  assign \new_[93630]_  = ~A200 & A199;
  assign \new_[93633]_  = A203 & A201;
  assign \new_[93634]_  = \new_[93633]_  & \new_[93630]_ ;
  assign \new_[93635]_  = \new_[93634]_  & \new_[93627]_ ;
  assign \new_[93638]_  = ~A235 & ~A233;
  assign \new_[93641]_  = ~A265 & ~A236;
  assign \new_[93642]_  = \new_[93641]_  & \new_[93638]_ ;
  assign \new_[93645]_  = A298 & ~A266;
  assign \new_[93648]_  = ~A302 & ~A301;
  assign \new_[93649]_  = \new_[93648]_  & \new_[93645]_ ;
  assign \new_[93650]_  = \new_[93649]_  & \new_[93642]_ ;
  assign \new_[93654]_  = ~A166 & ~A167;
  assign \new_[93655]_  = ~A169 & \new_[93654]_ ;
  assign \new_[93658]_  = ~A200 & A199;
  assign \new_[93661]_  = A203 & A201;
  assign \new_[93662]_  = \new_[93661]_  & \new_[93658]_ ;
  assign \new_[93663]_  = \new_[93662]_  & \new_[93655]_ ;
  assign \new_[93666]_  = ~A234 & ~A233;
  assign \new_[93669]_  = ~A268 & ~A266;
  assign \new_[93670]_  = \new_[93669]_  & \new_[93666]_ ;
  assign \new_[93673]_  = A298 & ~A269;
  assign \new_[93676]_  = ~A302 & ~A301;
  assign \new_[93677]_  = \new_[93676]_  & \new_[93673]_ ;
  assign \new_[93678]_  = \new_[93677]_  & \new_[93670]_ ;
  assign \new_[93682]_  = ~A166 & ~A167;
  assign \new_[93683]_  = ~A169 & \new_[93682]_ ;
  assign \new_[93686]_  = ~A200 & A199;
  assign \new_[93689]_  = A203 & A201;
  assign \new_[93690]_  = \new_[93689]_  & \new_[93686]_ ;
  assign \new_[93691]_  = \new_[93690]_  & \new_[93683]_ ;
  assign \new_[93694]_  = ~A233 & A232;
  assign \new_[93697]_  = A235 & A234;
  assign \new_[93698]_  = \new_[93697]_  & \new_[93694]_ ;
  assign \new_[93701]_  = ~A299 & A298;
  assign \new_[93704]_  = A301 & A300;
  assign \new_[93705]_  = \new_[93704]_  & \new_[93701]_ ;
  assign \new_[93706]_  = \new_[93705]_  & \new_[93698]_ ;
  assign \new_[93710]_  = ~A166 & ~A167;
  assign \new_[93711]_  = ~A169 & \new_[93710]_ ;
  assign \new_[93714]_  = ~A200 & A199;
  assign \new_[93717]_  = A203 & A201;
  assign \new_[93718]_  = \new_[93717]_  & \new_[93714]_ ;
  assign \new_[93719]_  = \new_[93718]_  & \new_[93711]_ ;
  assign \new_[93722]_  = ~A233 & A232;
  assign \new_[93725]_  = A235 & A234;
  assign \new_[93726]_  = \new_[93725]_  & \new_[93722]_ ;
  assign \new_[93729]_  = ~A299 & A298;
  assign \new_[93732]_  = A302 & A300;
  assign \new_[93733]_  = \new_[93732]_  & \new_[93729]_ ;
  assign \new_[93734]_  = \new_[93733]_  & \new_[93726]_ ;
  assign \new_[93738]_  = ~A166 & ~A167;
  assign \new_[93739]_  = ~A169 & \new_[93738]_ ;
  assign \new_[93742]_  = ~A200 & A199;
  assign \new_[93745]_  = A203 & A201;
  assign \new_[93746]_  = \new_[93745]_  & \new_[93742]_ ;
  assign \new_[93747]_  = \new_[93746]_  & \new_[93739]_ ;
  assign \new_[93750]_  = ~A233 & A232;
  assign \new_[93753]_  = A235 & A234;
  assign \new_[93754]_  = \new_[93753]_  & \new_[93750]_ ;
  assign \new_[93757]_  = ~A266 & A265;
  assign \new_[93760]_  = A268 & A267;
  assign \new_[93761]_  = \new_[93760]_  & \new_[93757]_ ;
  assign \new_[93762]_  = \new_[93761]_  & \new_[93754]_ ;
  assign \new_[93766]_  = ~A166 & ~A167;
  assign \new_[93767]_  = ~A169 & \new_[93766]_ ;
  assign \new_[93770]_  = ~A200 & A199;
  assign \new_[93773]_  = A203 & A201;
  assign \new_[93774]_  = \new_[93773]_  & \new_[93770]_ ;
  assign \new_[93775]_  = \new_[93774]_  & \new_[93767]_ ;
  assign \new_[93778]_  = ~A233 & A232;
  assign \new_[93781]_  = A235 & A234;
  assign \new_[93782]_  = \new_[93781]_  & \new_[93778]_ ;
  assign \new_[93785]_  = ~A266 & A265;
  assign \new_[93788]_  = A269 & A267;
  assign \new_[93789]_  = \new_[93788]_  & \new_[93785]_ ;
  assign \new_[93790]_  = \new_[93789]_  & \new_[93782]_ ;
  assign \new_[93794]_  = ~A166 & ~A167;
  assign \new_[93795]_  = ~A169 & \new_[93794]_ ;
  assign \new_[93798]_  = ~A200 & A199;
  assign \new_[93801]_  = A203 & A201;
  assign \new_[93802]_  = \new_[93801]_  & \new_[93798]_ ;
  assign \new_[93803]_  = \new_[93802]_  & \new_[93795]_ ;
  assign \new_[93806]_  = ~A233 & A232;
  assign \new_[93809]_  = A236 & A234;
  assign \new_[93810]_  = \new_[93809]_  & \new_[93806]_ ;
  assign \new_[93813]_  = ~A299 & A298;
  assign \new_[93816]_  = A301 & A300;
  assign \new_[93817]_  = \new_[93816]_  & \new_[93813]_ ;
  assign \new_[93818]_  = \new_[93817]_  & \new_[93810]_ ;
  assign \new_[93822]_  = ~A166 & ~A167;
  assign \new_[93823]_  = ~A169 & \new_[93822]_ ;
  assign \new_[93826]_  = ~A200 & A199;
  assign \new_[93829]_  = A203 & A201;
  assign \new_[93830]_  = \new_[93829]_  & \new_[93826]_ ;
  assign \new_[93831]_  = \new_[93830]_  & \new_[93823]_ ;
  assign \new_[93834]_  = ~A233 & A232;
  assign \new_[93837]_  = A236 & A234;
  assign \new_[93838]_  = \new_[93837]_  & \new_[93834]_ ;
  assign \new_[93841]_  = ~A299 & A298;
  assign \new_[93844]_  = A302 & A300;
  assign \new_[93845]_  = \new_[93844]_  & \new_[93841]_ ;
  assign \new_[93846]_  = \new_[93845]_  & \new_[93838]_ ;
  assign \new_[93850]_  = ~A166 & ~A167;
  assign \new_[93851]_  = ~A169 & \new_[93850]_ ;
  assign \new_[93854]_  = ~A200 & A199;
  assign \new_[93857]_  = A203 & A201;
  assign \new_[93858]_  = \new_[93857]_  & \new_[93854]_ ;
  assign \new_[93859]_  = \new_[93858]_  & \new_[93851]_ ;
  assign \new_[93862]_  = ~A233 & A232;
  assign \new_[93865]_  = A236 & A234;
  assign \new_[93866]_  = \new_[93865]_  & \new_[93862]_ ;
  assign \new_[93869]_  = ~A266 & A265;
  assign \new_[93872]_  = A268 & A267;
  assign \new_[93873]_  = \new_[93872]_  & \new_[93869]_ ;
  assign \new_[93874]_  = \new_[93873]_  & \new_[93866]_ ;
  assign \new_[93878]_  = ~A166 & ~A167;
  assign \new_[93879]_  = ~A169 & \new_[93878]_ ;
  assign \new_[93882]_  = ~A200 & A199;
  assign \new_[93885]_  = A203 & A201;
  assign \new_[93886]_  = \new_[93885]_  & \new_[93882]_ ;
  assign \new_[93887]_  = \new_[93886]_  & \new_[93879]_ ;
  assign \new_[93890]_  = ~A233 & A232;
  assign \new_[93893]_  = A236 & A234;
  assign \new_[93894]_  = \new_[93893]_  & \new_[93890]_ ;
  assign \new_[93897]_  = ~A266 & A265;
  assign \new_[93900]_  = A269 & A267;
  assign \new_[93901]_  = \new_[93900]_  & \new_[93897]_ ;
  assign \new_[93902]_  = \new_[93901]_  & \new_[93894]_ ;
  assign \new_[93906]_  = ~A166 & ~A167;
  assign \new_[93907]_  = ~A169 & \new_[93906]_ ;
  assign \new_[93910]_  = ~A200 & A199;
  assign \new_[93913]_  = A203 & A201;
  assign \new_[93914]_  = \new_[93913]_  & \new_[93910]_ ;
  assign \new_[93915]_  = \new_[93914]_  & \new_[93907]_ ;
  assign \new_[93918]_  = ~A233 & ~A232;
  assign \new_[93921]_  = ~A268 & ~A266;
  assign \new_[93922]_  = \new_[93921]_  & \new_[93918]_ ;
  assign \new_[93925]_  = A298 & ~A269;
  assign \new_[93928]_  = ~A302 & ~A301;
  assign \new_[93929]_  = \new_[93928]_  & \new_[93925]_ ;
  assign \new_[93930]_  = \new_[93929]_  & \new_[93922]_ ;
  assign \new_[93934]_  = A167 & ~A168;
  assign \new_[93935]_  = ~A169 & \new_[93934]_ ;
  assign \new_[93938]_  = ~A199 & A166;
  assign \new_[93941]_  = ~A233 & A200;
  assign \new_[93942]_  = \new_[93941]_  & \new_[93938]_ ;
  assign \new_[93943]_  = \new_[93942]_  & \new_[93935]_ ;
  assign \new_[93946]_  = ~A236 & ~A235;
  assign \new_[93949]_  = ~A268 & ~A266;
  assign \new_[93950]_  = \new_[93949]_  & \new_[93946]_ ;
  assign \new_[93953]_  = A298 & ~A269;
  assign \new_[93956]_  = ~A302 & ~A301;
  assign \new_[93957]_  = \new_[93956]_  & \new_[93953]_ ;
  assign \new_[93958]_  = \new_[93957]_  & \new_[93950]_ ;
  assign \new_[93962]_  = A167 & ~A168;
  assign \new_[93963]_  = ~A169 & \new_[93962]_ ;
  assign \new_[93966]_  = A199 & A166;
  assign \new_[93969]_  = A201 & ~A200;
  assign \new_[93970]_  = \new_[93969]_  & \new_[93966]_ ;
  assign \new_[93971]_  = \new_[93970]_  & \new_[93963]_ ;
  assign \new_[93974]_  = A232 & A202;
  assign \new_[93977]_  = A265 & A233;
  assign \new_[93978]_  = \new_[93977]_  & \new_[93974]_ ;
  assign \new_[93981]_  = ~A269 & ~A268;
  assign \new_[93984]_  = ~A300 & ~A299;
  assign \new_[93985]_  = \new_[93984]_  & \new_[93981]_ ;
  assign \new_[93986]_  = \new_[93985]_  & \new_[93978]_ ;
  assign \new_[93990]_  = A167 & ~A168;
  assign \new_[93991]_  = ~A169 & \new_[93990]_ ;
  assign \new_[93994]_  = A199 & A166;
  assign \new_[93997]_  = A201 & ~A200;
  assign \new_[93998]_  = \new_[93997]_  & \new_[93994]_ ;
  assign \new_[93999]_  = \new_[93998]_  & \new_[93991]_ ;
  assign \new_[94002]_  = A232 & A202;
  assign \new_[94005]_  = A265 & A233;
  assign \new_[94006]_  = \new_[94005]_  & \new_[94002]_ ;
  assign \new_[94009]_  = ~A269 & ~A268;
  assign \new_[94012]_  = A299 & A298;
  assign \new_[94013]_  = \new_[94012]_  & \new_[94009]_ ;
  assign \new_[94014]_  = \new_[94013]_  & \new_[94006]_ ;
  assign \new_[94018]_  = A167 & ~A168;
  assign \new_[94019]_  = ~A169 & \new_[94018]_ ;
  assign \new_[94022]_  = A199 & A166;
  assign \new_[94025]_  = A201 & ~A200;
  assign \new_[94026]_  = \new_[94025]_  & \new_[94022]_ ;
  assign \new_[94027]_  = \new_[94026]_  & \new_[94019]_ ;
  assign \new_[94030]_  = A232 & A202;
  assign \new_[94033]_  = A265 & A233;
  assign \new_[94034]_  = \new_[94033]_  & \new_[94030]_ ;
  assign \new_[94037]_  = ~A269 & ~A268;
  assign \new_[94040]_  = ~A299 & ~A298;
  assign \new_[94041]_  = \new_[94040]_  & \new_[94037]_ ;
  assign \new_[94042]_  = \new_[94041]_  & \new_[94034]_ ;
  assign \new_[94046]_  = A167 & ~A168;
  assign \new_[94047]_  = ~A169 & \new_[94046]_ ;
  assign \new_[94050]_  = A199 & A166;
  assign \new_[94053]_  = A201 & ~A200;
  assign \new_[94054]_  = \new_[94053]_  & \new_[94050]_ ;
  assign \new_[94055]_  = \new_[94054]_  & \new_[94047]_ ;
  assign \new_[94058]_  = A232 & A202;
  assign \new_[94061]_  = A265 & A233;
  assign \new_[94062]_  = \new_[94061]_  & \new_[94058]_ ;
  assign \new_[94065]_  = ~A299 & ~A267;
  assign \new_[94068]_  = ~A302 & ~A301;
  assign \new_[94069]_  = \new_[94068]_  & \new_[94065]_ ;
  assign \new_[94070]_  = \new_[94069]_  & \new_[94062]_ ;
  assign \new_[94074]_  = A167 & ~A168;
  assign \new_[94075]_  = ~A169 & \new_[94074]_ ;
  assign \new_[94078]_  = A199 & A166;
  assign \new_[94081]_  = A201 & ~A200;
  assign \new_[94082]_  = \new_[94081]_  & \new_[94078]_ ;
  assign \new_[94083]_  = \new_[94082]_  & \new_[94075]_ ;
  assign \new_[94086]_  = A232 & A202;
  assign \new_[94089]_  = A265 & A233;
  assign \new_[94090]_  = \new_[94089]_  & \new_[94086]_ ;
  assign \new_[94093]_  = ~A299 & A266;
  assign \new_[94096]_  = ~A302 & ~A301;
  assign \new_[94097]_  = \new_[94096]_  & \new_[94093]_ ;
  assign \new_[94098]_  = \new_[94097]_  & \new_[94090]_ ;
  assign \new_[94102]_  = A167 & ~A168;
  assign \new_[94103]_  = ~A169 & \new_[94102]_ ;
  assign \new_[94106]_  = A199 & A166;
  assign \new_[94109]_  = A201 & ~A200;
  assign \new_[94110]_  = \new_[94109]_  & \new_[94106]_ ;
  assign \new_[94111]_  = \new_[94110]_  & \new_[94103]_ ;
  assign \new_[94114]_  = A232 & A202;
  assign \new_[94117]_  = ~A265 & A233;
  assign \new_[94118]_  = \new_[94117]_  & \new_[94114]_ ;
  assign \new_[94121]_  = ~A299 & ~A266;
  assign \new_[94124]_  = ~A302 & ~A301;
  assign \new_[94125]_  = \new_[94124]_  & \new_[94121]_ ;
  assign \new_[94126]_  = \new_[94125]_  & \new_[94118]_ ;
  assign \new_[94130]_  = A167 & ~A168;
  assign \new_[94131]_  = ~A169 & \new_[94130]_ ;
  assign \new_[94134]_  = A199 & A166;
  assign \new_[94137]_  = A201 & ~A200;
  assign \new_[94138]_  = \new_[94137]_  & \new_[94134]_ ;
  assign \new_[94139]_  = \new_[94138]_  & \new_[94131]_ ;
  assign \new_[94142]_  = ~A233 & A202;
  assign \new_[94145]_  = ~A236 & ~A235;
  assign \new_[94146]_  = \new_[94145]_  & \new_[94142]_ ;
  assign \new_[94149]_  = A266 & A265;
  assign \new_[94152]_  = ~A300 & A298;
  assign \new_[94153]_  = \new_[94152]_  & \new_[94149]_ ;
  assign \new_[94154]_  = \new_[94153]_  & \new_[94146]_ ;
  assign \new_[94158]_  = A167 & ~A168;
  assign \new_[94159]_  = ~A169 & \new_[94158]_ ;
  assign \new_[94162]_  = A199 & A166;
  assign \new_[94165]_  = A201 & ~A200;
  assign \new_[94166]_  = \new_[94165]_  & \new_[94162]_ ;
  assign \new_[94167]_  = \new_[94166]_  & \new_[94159]_ ;
  assign \new_[94170]_  = ~A233 & A202;
  assign \new_[94173]_  = ~A236 & ~A235;
  assign \new_[94174]_  = \new_[94173]_  & \new_[94170]_ ;
  assign \new_[94177]_  = A266 & A265;
  assign \new_[94180]_  = A299 & A298;
  assign \new_[94181]_  = \new_[94180]_  & \new_[94177]_ ;
  assign \new_[94182]_  = \new_[94181]_  & \new_[94174]_ ;
  assign \new_[94186]_  = A167 & ~A168;
  assign \new_[94187]_  = ~A169 & \new_[94186]_ ;
  assign \new_[94190]_  = A199 & A166;
  assign \new_[94193]_  = A201 & ~A200;
  assign \new_[94194]_  = \new_[94193]_  & \new_[94190]_ ;
  assign \new_[94195]_  = \new_[94194]_  & \new_[94187]_ ;
  assign \new_[94198]_  = ~A233 & A202;
  assign \new_[94201]_  = ~A236 & ~A235;
  assign \new_[94202]_  = \new_[94201]_  & \new_[94198]_ ;
  assign \new_[94205]_  = A266 & A265;
  assign \new_[94208]_  = ~A299 & ~A298;
  assign \new_[94209]_  = \new_[94208]_  & \new_[94205]_ ;
  assign \new_[94210]_  = \new_[94209]_  & \new_[94202]_ ;
  assign \new_[94214]_  = A167 & ~A168;
  assign \new_[94215]_  = ~A169 & \new_[94214]_ ;
  assign \new_[94218]_  = A199 & A166;
  assign \new_[94221]_  = A201 & ~A200;
  assign \new_[94222]_  = \new_[94221]_  & \new_[94218]_ ;
  assign \new_[94223]_  = \new_[94222]_  & \new_[94215]_ ;
  assign \new_[94226]_  = ~A233 & A202;
  assign \new_[94229]_  = ~A236 & ~A235;
  assign \new_[94230]_  = \new_[94229]_  & \new_[94226]_ ;
  assign \new_[94233]_  = ~A267 & ~A266;
  assign \new_[94236]_  = ~A300 & A298;
  assign \new_[94237]_  = \new_[94236]_  & \new_[94233]_ ;
  assign \new_[94238]_  = \new_[94237]_  & \new_[94230]_ ;
  assign \new_[94242]_  = A167 & ~A168;
  assign \new_[94243]_  = ~A169 & \new_[94242]_ ;
  assign \new_[94246]_  = A199 & A166;
  assign \new_[94249]_  = A201 & ~A200;
  assign \new_[94250]_  = \new_[94249]_  & \new_[94246]_ ;
  assign \new_[94251]_  = \new_[94250]_  & \new_[94243]_ ;
  assign \new_[94254]_  = ~A233 & A202;
  assign \new_[94257]_  = ~A236 & ~A235;
  assign \new_[94258]_  = \new_[94257]_  & \new_[94254]_ ;
  assign \new_[94261]_  = ~A267 & ~A266;
  assign \new_[94264]_  = A299 & A298;
  assign \new_[94265]_  = \new_[94264]_  & \new_[94261]_ ;
  assign \new_[94266]_  = \new_[94265]_  & \new_[94258]_ ;
  assign \new_[94270]_  = A167 & ~A168;
  assign \new_[94271]_  = ~A169 & \new_[94270]_ ;
  assign \new_[94274]_  = A199 & A166;
  assign \new_[94277]_  = A201 & ~A200;
  assign \new_[94278]_  = \new_[94277]_  & \new_[94274]_ ;
  assign \new_[94279]_  = \new_[94278]_  & \new_[94271]_ ;
  assign \new_[94282]_  = ~A233 & A202;
  assign \new_[94285]_  = ~A236 & ~A235;
  assign \new_[94286]_  = \new_[94285]_  & \new_[94282]_ ;
  assign \new_[94289]_  = ~A267 & ~A266;
  assign \new_[94292]_  = ~A299 & ~A298;
  assign \new_[94293]_  = \new_[94292]_  & \new_[94289]_ ;
  assign \new_[94294]_  = \new_[94293]_  & \new_[94286]_ ;
  assign \new_[94298]_  = A167 & ~A168;
  assign \new_[94299]_  = ~A169 & \new_[94298]_ ;
  assign \new_[94302]_  = A199 & A166;
  assign \new_[94305]_  = A201 & ~A200;
  assign \new_[94306]_  = \new_[94305]_  & \new_[94302]_ ;
  assign \new_[94307]_  = \new_[94306]_  & \new_[94299]_ ;
  assign \new_[94310]_  = ~A233 & A202;
  assign \new_[94313]_  = ~A236 & ~A235;
  assign \new_[94314]_  = \new_[94313]_  & \new_[94310]_ ;
  assign \new_[94317]_  = ~A266 & ~A265;
  assign \new_[94320]_  = ~A300 & A298;
  assign \new_[94321]_  = \new_[94320]_  & \new_[94317]_ ;
  assign \new_[94322]_  = \new_[94321]_  & \new_[94314]_ ;
  assign \new_[94326]_  = A167 & ~A168;
  assign \new_[94327]_  = ~A169 & \new_[94326]_ ;
  assign \new_[94330]_  = A199 & A166;
  assign \new_[94333]_  = A201 & ~A200;
  assign \new_[94334]_  = \new_[94333]_  & \new_[94330]_ ;
  assign \new_[94335]_  = \new_[94334]_  & \new_[94327]_ ;
  assign \new_[94338]_  = ~A233 & A202;
  assign \new_[94341]_  = ~A236 & ~A235;
  assign \new_[94342]_  = \new_[94341]_  & \new_[94338]_ ;
  assign \new_[94345]_  = ~A266 & ~A265;
  assign \new_[94348]_  = A299 & A298;
  assign \new_[94349]_  = \new_[94348]_  & \new_[94345]_ ;
  assign \new_[94350]_  = \new_[94349]_  & \new_[94342]_ ;
  assign \new_[94354]_  = A167 & ~A168;
  assign \new_[94355]_  = ~A169 & \new_[94354]_ ;
  assign \new_[94358]_  = A199 & A166;
  assign \new_[94361]_  = A201 & ~A200;
  assign \new_[94362]_  = \new_[94361]_  & \new_[94358]_ ;
  assign \new_[94363]_  = \new_[94362]_  & \new_[94355]_ ;
  assign \new_[94366]_  = ~A233 & A202;
  assign \new_[94369]_  = ~A236 & ~A235;
  assign \new_[94370]_  = \new_[94369]_  & \new_[94366]_ ;
  assign \new_[94373]_  = ~A266 & ~A265;
  assign \new_[94376]_  = ~A299 & ~A298;
  assign \new_[94377]_  = \new_[94376]_  & \new_[94373]_ ;
  assign \new_[94378]_  = \new_[94377]_  & \new_[94370]_ ;
  assign \new_[94382]_  = A167 & ~A168;
  assign \new_[94383]_  = ~A169 & \new_[94382]_ ;
  assign \new_[94386]_  = A199 & A166;
  assign \new_[94389]_  = A201 & ~A200;
  assign \new_[94390]_  = \new_[94389]_  & \new_[94386]_ ;
  assign \new_[94391]_  = \new_[94390]_  & \new_[94383]_ ;
  assign \new_[94394]_  = ~A233 & A202;
  assign \new_[94397]_  = A265 & ~A234;
  assign \new_[94398]_  = \new_[94397]_  & \new_[94394]_ ;
  assign \new_[94401]_  = A298 & A266;
  assign \new_[94404]_  = ~A302 & ~A301;
  assign \new_[94405]_  = \new_[94404]_  & \new_[94401]_ ;
  assign \new_[94406]_  = \new_[94405]_  & \new_[94398]_ ;
  assign \new_[94410]_  = A167 & ~A168;
  assign \new_[94411]_  = ~A169 & \new_[94410]_ ;
  assign \new_[94414]_  = A199 & A166;
  assign \new_[94417]_  = A201 & ~A200;
  assign \new_[94418]_  = \new_[94417]_  & \new_[94414]_ ;
  assign \new_[94419]_  = \new_[94418]_  & \new_[94411]_ ;
  assign \new_[94422]_  = ~A233 & A202;
  assign \new_[94425]_  = ~A266 & ~A234;
  assign \new_[94426]_  = \new_[94425]_  & \new_[94422]_ ;
  assign \new_[94429]_  = ~A269 & ~A268;
  assign \new_[94432]_  = ~A300 & A298;
  assign \new_[94433]_  = \new_[94432]_  & \new_[94429]_ ;
  assign \new_[94434]_  = \new_[94433]_  & \new_[94426]_ ;
  assign \new_[94438]_  = A167 & ~A168;
  assign \new_[94439]_  = ~A169 & \new_[94438]_ ;
  assign \new_[94442]_  = A199 & A166;
  assign \new_[94445]_  = A201 & ~A200;
  assign \new_[94446]_  = \new_[94445]_  & \new_[94442]_ ;
  assign \new_[94447]_  = \new_[94446]_  & \new_[94439]_ ;
  assign \new_[94450]_  = ~A233 & A202;
  assign \new_[94453]_  = ~A266 & ~A234;
  assign \new_[94454]_  = \new_[94453]_  & \new_[94450]_ ;
  assign \new_[94457]_  = ~A269 & ~A268;
  assign \new_[94460]_  = A299 & A298;
  assign \new_[94461]_  = \new_[94460]_  & \new_[94457]_ ;
  assign \new_[94462]_  = \new_[94461]_  & \new_[94454]_ ;
  assign \new_[94466]_  = A167 & ~A168;
  assign \new_[94467]_  = ~A169 & \new_[94466]_ ;
  assign \new_[94470]_  = A199 & A166;
  assign \new_[94473]_  = A201 & ~A200;
  assign \new_[94474]_  = \new_[94473]_  & \new_[94470]_ ;
  assign \new_[94475]_  = \new_[94474]_  & \new_[94467]_ ;
  assign \new_[94478]_  = ~A233 & A202;
  assign \new_[94481]_  = ~A266 & ~A234;
  assign \new_[94482]_  = \new_[94481]_  & \new_[94478]_ ;
  assign \new_[94485]_  = ~A269 & ~A268;
  assign \new_[94488]_  = ~A299 & ~A298;
  assign \new_[94489]_  = \new_[94488]_  & \new_[94485]_ ;
  assign \new_[94490]_  = \new_[94489]_  & \new_[94482]_ ;
  assign \new_[94494]_  = A167 & ~A168;
  assign \new_[94495]_  = ~A169 & \new_[94494]_ ;
  assign \new_[94498]_  = A199 & A166;
  assign \new_[94501]_  = A201 & ~A200;
  assign \new_[94502]_  = \new_[94501]_  & \new_[94498]_ ;
  assign \new_[94503]_  = \new_[94502]_  & \new_[94495]_ ;
  assign \new_[94506]_  = ~A233 & A202;
  assign \new_[94509]_  = ~A266 & ~A234;
  assign \new_[94510]_  = \new_[94509]_  & \new_[94506]_ ;
  assign \new_[94513]_  = A298 & ~A267;
  assign \new_[94516]_  = ~A302 & ~A301;
  assign \new_[94517]_  = \new_[94516]_  & \new_[94513]_ ;
  assign \new_[94518]_  = \new_[94517]_  & \new_[94510]_ ;
  assign \new_[94522]_  = A167 & ~A168;
  assign \new_[94523]_  = ~A169 & \new_[94522]_ ;
  assign \new_[94526]_  = A199 & A166;
  assign \new_[94529]_  = A201 & ~A200;
  assign \new_[94530]_  = \new_[94529]_  & \new_[94526]_ ;
  assign \new_[94531]_  = \new_[94530]_  & \new_[94523]_ ;
  assign \new_[94534]_  = ~A233 & A202;
  assign \new_[94537]_  = ~A265 & ~A234;
  assign \new_[94538]_  = \new_[94537]_  & \new_[94534]_ ;
  assign \new_[94541]_  = A298 & ~A266;
  assign \new_[94544]_  = ~A302 & ~A301;
  assign \new_[94545]_  = \new_[94544]_  & \new_[94541]_ ;
  assign \new_[94546]_  = \new_[94545]_  & \new_[94538]_ ;
  assign \new_[94550]_  = A167 & ~A168;
  assign \new_[94551]_  = ~A169 & \new_[94550]_ ;
  assign \new_[94554]_  = A199 & A166;
  assign \new_[94557]_  = A201 & ~A200;
  assign \new_[94558]_  = \new_[94557]_  & \new_[94554]_ ;
  assign \new_[94559]_  = \new_[94558]_  & \new_[94551]_ ;
  assign \new_[94562]_  = ~A232 & A202;
  assign \new_[94565]_  = A265 & ~A233;
  assign \new_[94566]_  = \new_[94565]_  & \new_[94562]_ ;
  assign \new_[94569]_  = A298 & A266;
  assign \new_[94572]_  = ~A302 & ~A301;
  assign \new_[94573]_  = \new_[94572]_  & \new_[94569]_ ;
  assign \new_[94574]_  = \new_[94573]_  & \new_[94566]_ ;
  assign \new_[94578]_  = A167 & ~A168;
  assign \new_[94579]_  = ~A169 & \new_[94578]_ ;
  assign \new_[94582]_  = A199 & A166;
  assign \new_[94585]_  = A201 & ~A200;
  assign \new_[94586]_  = \new_[94585]_  & \new_[94582]_ ;
  assign \new_[94587]_  = \new_[94586]_  & \new_[94579]_ ;
  assign \new_[94590]_  = ~A232 & A202;
  assign \new_[94593]_  = ~A266 & ~A233;
  assign \new_[94594]_  = \new_[94593]_  & \new_[94590]_ ;
  assign \new_[94597]_  = ~A269 & ~A268;
  assign \new_[94600]_  = ~A300 & A298;
  assign \new_[94601]_  = \new_[94600]_  & \new_[94597]_ ;
  assign \new_[94602]_  = \new_[94601]_  & \new_[94594]_ ;
  assign \new_[94606]_  = A167 & ~A168;
  assign \new_[94607]_  = ~A169 & \new_[94606]_ ;
  assign \new_[94610]_  = A199 & A166;
  assign \new_[94613]_  = A201 & ~A200;
  assign \new_[94614]_  = \new_[94613]_  & \new_[94610]_ ;
  assign \new_[94615]_  = \new_[94614]_  & \new_[94607]_ ;
  assign \new_[94618]_  = ~A232 & A202;
  assign \new_[94621]_  = ~A266 & ~A233;
  assign \new_[94622]_  = \new_[94621]_  & \new_[94618]_ ;
  assign \new_[94625]_  = ~A269 & ~A268;
  assign \new_[94628]_  = A299 & A298;
  assign \new_[94629]_  = \new_[94628]_  & \new_[94625]_ ;
  assign \new_[94630]_  = \new_[94629]_  & \new_[94622]_ ;
  assign \new_[94634]_  = A167 & ~A168;
  assign \new_[94635]_  = ~A169 & \new_[94634]_ ;
  assign \new_[94638]_  = A199 & A166;
  assign \new_[94641]_  = A201 & ~A200;
  assign \new_[94642]_  = \new_[94641]_  & \new_[94638]_ ;
  assign \new_[94643]_  = \new_[94642]_  & \new_[94635]_ ;
  assign \new_[94646]_  = ~A232 & A202;
  assign \new_[94649]_  = ~A266 & ~A233;
  assign \new_[94650]_  = \new_[94649]_  & \new_[94646]_ ;
  assign \new_[94653]_  = ~A269 & ~A268;
  assign \new_[94656]_  = ~A299 & ~A298;
  assign \new_[94657]_  = \new_[94656]_  & \new_[94653]_ ;
  assign \new_[94658]_  = \new_[94657]_  & \new_[94650]_ ;
  assign \new_[94662]_  = A167 & ~A168;
  assign \new_[94663]_  = ~A169 & \new_[94662]_ ;
  assign \new_[94666]_  = A199 & A166;
  assign \new_[94669]_  = A201 & ~A200;
  assign \new_[94670]_  = \new_[94669]_  & \new_[94666]_ ;
  assign \new_[94671]_  = \new_[94670]_  & \new_[94663]_ ;
  assign \new_[94674]_  = ~A232 & A202;
  assign \new_[94677]_  = ~A266 & ~A233;
  assign \new_[94678]_  = \new_[94677]_  & \new_[94674]_ ;
  assign \new_[94681]_  = A298 & ~A267;
  assign \new_[94684]_  = ~A302 & ~A301;
  assign \new_[94685]_  = \new_[94684]_  & \new_[94681]_ ;
  assign \new_[94686]_  = \new_[94685]_  & \new_[94678]_ ;
  assign \new_[94690]_  = A167 & ~A168;
  assign \new_[94691]_  = ~A169 & \new_[94690]_ ;
  assign \new_[94694]_  = A199 & A166;
  assign \new_[94697]_  = A201 & ~A200;
  assign \new_[94698]_  = \new_[94697]_  & \new_[94694]_ ;
  assign \new_[94699]_  = \new_[94698]_  & \new_[94691]_ ;
  assign \new_[94702]_  = ~A232 & A202;
  assign \new_[94705]_  = ~A265 & ~A233;
  assign \new_[94706]_  = \new_[94705]_  & \new_[94702]_ ;
  assign \new_[94709]_  = A298 & ~A266;
  assign \new_[94712]_  = ~A302 & ~A301;
  assign \new_[94713]_  = \new_[94712]_  & \new_[94709]_ ;
  assign \new_[94714]_  = \new_[94713]_  & \new_[94706]_ ;
  assign \new_[94718]_  = A167 & ~A168;
  assign \new_[94719]_  = ~A169 & \new_[94718]_ ;
  assign \new_[94722]_  = A199 & A166;
  assign \new_[94725]_  = A201 & ~A200;
  assign \new_[94726]_  = \new_[94725]_  & \new_[94722]_ ;
  assign \new_[94727]_  = \new_[94726]_  & \new_[94719]_ ;
  assign \new_[94730]_  = A232 & A203;
  assign \new_[94733]_  = A265 & A233;
  assign \new_[94734]_  = \new_[94733]_  & \new_[94730]_ ;
  assign \new_[94737]_  = ~A269 & ~A268;
  assign \new_[94740]_  = ~A300 & ~A299;
  assign \new_[94741]_  = \new_[94740]_  & \new_[94737]_ ;
  assign \new_[94742]_  = \new_[94741]_  & \new_[94734]_ ;
  assign \new_[94746]_  = A167 & ~A168;
  assign \new_[94747]_  = ~A169 & \new_[94746]_ ;
  assign \new_[94750]_  = A199 & A166;
  assign \new_[94753]_  = A201 & ~A200;
  assign \new_[94754]_  = \new_[94753]_  & \new_[94750]_ ;
  assign \new_[94755]_  = \new_[94754]_  & \new_[94747]_ ;
  assign \new_[94758]_  = A232 & A203;
  assign \new_[94761]_  = A265 & A233;
  assign \new_[94762]_  = \new_[94761]_  & \new_[94758]_ ;
  assign \new_[94765]_  = ~A269 & ~A268;
  assign \new_[94768]_  = A299 & A298;
  assign \new_[94769]_  = \new_[94768]_  & \new_[94765]_ ;
  assign \new_[94770]_  = \new_[94769]_  & \new_[94762]_ ;
  assign \new_[94774]_  = A167 & ~A168;
  assign \new_[94775]_  = ~A169 & \new_[94774]_ ;
  assign \new_[94778]_  = A199 & A166;
  assign \new_[94781]_  = A201 & ~A200;
  assign \new_[94782]_  = \new_[94781]_  & \new_[94778]_ ;
  assign \new_[94783]_  = \new_[94782]_  & \new_[94775]_ ;
  assign \new_[94786]_  = A232 & A203;
  assign \new_[94789]_  = A265 & A233;
  assign \new_[94790]_  = \new_[94789]_  & \new_[94786]_ ;
  assign \new_[94793]_  = ~A269 & ~A268;
  assign \new_[94796]_  = ~A299 & ~A298;
  assign \new_[94797]_  = \new_[94796]_  & \new_[94793]_ ;
  assign \new_[94798]_  = \new_[94797]_  & \new_[94790]_ ;
  assign \new_[94802]_  = A167 & ~A168;
  assign \new_[94803]_  = ~A169 & \new_[94802]_ ;
  assign \new_[94806]_  = A199 & A166;
  assign \new_[94809]_  = A201 & ~A200;
  assign \new_[94810]_  = \new_[94809]_  & \new_[94806]_ ;
  assign \new_[94811]_  = \new_[94810]_  & \new_[94803]_ ;
  assign \new_[94814]_  = A232 & A203;
  assign \new_[94817]_  = A265 & A233;
  assign \new_[94818]_  = \new_[94817]_  & \new_[94814]_ ;
  assign \new_[94821]_  = ~A299 & ~A267;
  assign \new_[94824]_  = ~A302 & ~A301;
  assign \new_[94825]_  = \new_[94824]_  & \new_[94821]_ ;
  assign \new_[94826]_  = \new_[94825]_  & \new_[94818]_ ;
  assign \new_[94830]_  = A167 & ~A168;
  assign \new_[94831]_  = ~A169 & \new_[94830]_ ;
  assign \new_[94834]_  = A199 & A166;
  assign \new_[94837]_  = A201 & ~A200;
  assign \new_[94838]_  = \new_[94837]_  & \new_[94834]_ ;
  assign \new_[94839]_  = \new_[94838]_  & \new_[94831]_ ;
  assign \new_[94842]_  = A232 & A203;
  assign \new_[94845]_  = A265 & A233;
  assign \new_[94846]_  = \new_[94845]_  & \new_[94842]_ ;
  assign \new_[94849]_  = ~A299 & A266;
  assign \new_[94852]_  = ~A302 & ~A301;
  assign \new_[94853]_  = \new_[94852]_  & \new_[94849]_ ;
  assign \new_[94854]_  = \new_[94853]_  & \new_[94846]_ ;
  assign \new_[94858]_  = A167 & ~A168;
  assign \new_[94859]_  = ~A169 & \new_[94858]_ ;
  assign \new_[94862]_  = A199 & A166;
  assign \new_[94865]_  = A201 & ~A200;
  assign \new_[94866]_  = \new_[94865]_  & \new_[94862]_ ;
  assign \new_[94867]_  = \new_[94866]_  & \new_[94859]_ ;
  assign \new_[94870]_  = A232 & A203;
  assign \new_[94873]_  = ~A265 & A233;
  assign \new_[94874]_  = \new_[94873]_  & \new_[94870]_ ;
  assign \new_[94877]_  = ~A299 & ~A266;
  assign \new_[94880]_  = ~A302 & ~A301;
  assign \new_[94881]_  = \new_[94880]_  & \new_[94877]_ ;
  assign \new_[94882]_  = \new_[94881]_  & \new_[94874]_ ;
  assign \new_[94886]_  = A167 & ~A168;
  assign \new_[94887]_  = ~A169 & \new_[94886]_ ;
  assign \new_[94890]_  = A199 & A166;
  assign \new_[94893]_  = A201 & ~A200;
  assign \new_[94894]_  = \new_[94893]_  & \new_[94890]_ ;
  assign \new_[94895]_  = \new_[94894]_  & \new_[94887]_ ;
  assign \new_[94898]_  = ~A233 & A203;
  assign \new_[94901]_  = ~A236 & ~A235;
  assign \new_[94902]_  = \new_[94901]_  & \new_[94898]_ ;
  assign \new_[94905]_  = A266 & A265;
  assign \new_[94908]_  = ~A300 & A298;
  assign \new_[94909]_  = \new_[94908]_  & \new_[94905]_ ;
  assign \new_[94910]_  = \new_[94909]_  & \new_[94902]_ ;
  assign \new_[94914]_  = A167 & ~A168;
  assign \new_[94915]_  = ~A169 & \new_[94914]_ ;
  assign \new_[94918]_  = A199 & A166;
  assign \new_[94921]_  = A201 & ~A200;
  assign \new_[94922]_  = \new_[94921]_  & \new_[94918]_ ;
  assign \new_[94923]_  = \new_[94922]_  & \new_[94915]_ ;
  assign \new_[94926]_  = ~A233 & A203;
  assign \new_[94929]_  = ~A236 & ~A235;
  assign \new_[94930]_  = \new_[94929]_  & \new_[94926]_ ;
  assign \new_[94933]_  = A266 & A265;
  assign \new_[94936]_  = A299 & A298;
  assign \new_[94937]_  = \new_[94936]_  & \new_[94933]_ ;
  assign \new_[94938]_  = \new_[94937]_  & \new_[94930]_ ;
  assign \new_[94942]_  = A167 & ~A168;
  assign \new_[94943]_  = ~A169 & \new_[94942]_ ;
  assign \new_[94946]_  = A199 & A166;
  assign \new_[94949]_  = A201 & ~A200;
  assign \new_[94950]_  = \new_[94949]_  & \new_[94946]_ ;
  assign \new_[94951]_  = \new_[94950]_  & \new_[94943]_ ;
  assign \new_[94954]_  = ~A233 & A203;
  assign \new_[94957]_  = ~A236 & ~A235;
  assign \new_[94958]_  = \new_[94957]_  & \new_[94954]_ ;
  assign \new_[94961]_  = A266 & A265;
  assign \new_[94964]_  = ~A299 & ~A298;
  assign \new_[94965]_  = \new_[94964]_  & \new_[94961]_ ;
  assign \new_[94966]_  = \new_[94965]_  & \new_[94958]_ ;
  assign \new_[94970]_  = A167 & ~A168;
  assign \new_[94971]_  = ~A169 & \new_[94970]_ ;
  assign \new_[94974]_  = A199 & A166;
  assign \new_[94977]_  = A201 & ~A200;
  assign \new_[94978]_  = \new_[94977]_  & \new_[94974]_ ;
  assign \new_[94979]_  = \new_[94978]_  & \new_[94971]_ ;
  assign \new_[94982]_  = ~A233 & A203;
  assign \new_[94985]_  = ~A236 & ~A235;
  assign \new_[94986]_  = \new_[94985]_  & \new_[94982]_ ;
  assign \new_[94989]_  = ~A267 & ~A266;
  assign \new_[94992]_  = ~A300 & A298;
  assign \new_[94993]_  = \new_[94992]_  & \new_[94989]_ ;
  assign \new_[94994]_  = \new_[94993]_  & \new_[94986]_ ;
  assign \new_[94998]_  = A167 & ~A168;
  assign \new_[94999]_  = ~A169 & \new_[94998]_ ;
  assign \new_[95002]_  = A199 & A166;
  assign \new_[95005]_  = A201 & ~A200;
  assign \new_[95006]_  = \new_[95005]_  & \new_[95002]_ ;
  assign \new_[95007]_  = \new_[95006]_  & \new_[94999]_ ;
  assign \new_[95010]_  = ~A233 & A203;
  assign \new_[95013]_  = ~A236 & ~A235;
  assign \new_[95014]_  = \new_[95013]_  & \new_[95010]_ ;
  assign \new_[95017]_  = ~A267 & ~A266;
  assign \new_[95020]_  = A299 & A298;
  assign \new_[95021]_  = \new_[95020]_  & \new_[95017]_ ;
  assign \new_[95022]_  = \new_[95021]_  & \new_[95014]_ ;
  assign \new_[95026]_  = A167 & ~A168;
  assign \new_[95027]_  = ~A169 & \new_[95026]_ ;
  assign \new_[95030]_  = A199 & A166;
  assign \new_[95033]_  = A201 & ~A200;
  assign \new_[95034]_  = \new_[95033]_  & \new_[95030]_ ;
  assign \new_[95035]_  = \new_[95034]_  & \new_[95027]_ ;
  assign \new_[95038]_  = ~A233 & A203;
  assign \new_[95041]_  = ~A236 & ~A235;
  assign \new_[95042]_  = \new_[95041]_  & \new_[95038]_ ;
  assign \new_[95045]_  = ~A267 & ~A266;
  assign \new_[95048]_  = ~A299 & ~A298;
  assign \new_[95049]_  = \new_[95048]_  & \new_[95045]_ ;
  assign \new_[95050]_  = \new_[95049]_  & \new_[95042]_ ;
  assign \new_[95054]_  = A167 & ~A168;
  assign \new_[95055]_  = ~A169 & \new_[95054]_ ;
  assign \new_[95058]_  = A199 & A166;
  assign \new_[95061]_  = A201 & ~A200;
  assign \new_[95062]_  = \new_[95061]_  & \new_[95058]_ ;
  assign \new_[95063]_  = \new_[95062]_  & \new_[95055]_ ;
  assign \new_[95066]_  = ~A233 & A203;
  assign \new_[95069]_  = ~A236 & ~A235;
  assign \new_[95070]_  = \new_[95069]_  & \new_[95066]_ ;
  assign \new_[95073]_  = ~A266 & ~A265;
  assign \new_[95076]_  = ~A300 & A298;
  assign \new_[95077]_  = \new_[95076]_  & \new_[95073]_ ;
  assign \new_[95078]_  = \new_[95077]_  & \new_[95070]_ ;
  assign \new_[95082]_  = A167 & ~A168;
  assign \new_[95083]_  = ~A169 & \new_[95082]_ ;
  assign \new_[95086]_  = A199 & A166;
  assign \new_[95089]_  = A201 & ~A200;
  assign \new_[95090]_  = \new_[95089]_  & \new_[95086]_ ;
  assign \new_[95091]_  = \new_[95090]_  & \new_[95083]_ ;
  assign \new_[95094]_  = ~A233 & A203;
  assign \new_[95097]_  = ~A236 & ~A235;
  assign \new_[95098]_  = \new_[95097]_  & \new_[95094]_ ;
  assign \new_[95101]_  = ~A266 & ~A265;
  assign \new_[95104]_  = A299 & A298;
  assign \new_[95105]_  = \new_[95104]_  & \new_[95101]_ ;
  assign \new_[95106]_  = \new_[95105]_  & \new_[95098]_ ;
  assign \new_[95110]_  = A167 & ~A168;
  assign \new_[95111]_  = ~A169 & \new_[95110]_ ;
  assign \new_[95114]_  = A199 & A166;
  assign \new_[95117]_  = A201 & ~A200;
  assign \new_[95118]_  = \new_[95117]_  & \new_[95114]_ ;
  assign \new_[95119]_  = \new_[95118]_  & \new_[95111]_ ;
  assign \new_[95122]_  = ~A233 & A203;
  assign \new_[95125]_  = ~A236 & ~A235;
  assign \new_[95126]_  = \new_[95125]_  & \new_[95122]_ ;
  assign \new_[95129]_  = ~A266 & ~A265;
  assign \new_[95132]_  = ~A299 & ~A298;
  assign \new_[95133]_  = \new_[95132]_  & \new_[95129]_ ;
  assign \new_[95134]_  = \new_[95133]_  & \new_[95126]_ ;
  assign \new_[95138]_  = A167 & ~A168;
  assign \new_[95139]_  = ~A169 & \new_[95138]_ ;
  assign \new_[95142]_  = A199 & A166;
  assign \new_[95145]_  = A201 & ~A200;
  assign \new_[95146]_  = \new_[95145]_  & \new_[95142]_ ;
  assign \new_[95147]_  = \new_[95146]_  & \new_[95139]_ ;
  assign \new_[95150]_  = ~A233 & A203;
  assign \new_[95153]_  = A265 & ~A234;
  assign \new_[95154]_  = \new_[95153]_  & \new_[95150]_ ;
  assign \new_[95157]_  = A298 & A266;
  assign \new_[95160]_  = ~A302 & ~A301;
  assign \new_[95161]_  = \new_[95160]_  & \new_[95157]_ ;
  assign \new_[95162]_  = \new_[95161]_  & \new_[95154]_ ;
  assign \new_[95166]_  = A167 & ~A168;
  assign \new_[95167]_  = ~A169 & \new_[95166]_ ;
  assign \new_[95170]_  = A199 & A166;
  assign \new_[95173]_  = A201 & ~A200;
  assign \new_[95174]_  = \new_[95173]_  & \new_[95170]_ ;
  assign \new_[95175]_  = \new_[95174]_  & \new_[95167]_ ;
  assign \new_[95178]_  = ~A233 & A203;
  assign \new_[95181]_  = ~A266 & ~A234;
  assign \new_[95182]_  = \new_[95181]_  & \new_[95178]_ ;
  assign \new_[95185]_  = ~A269 & ~A268;
  assign \new_[95188]_  = ~A300 & A298;
  assign \new_[95189]_  = \new_[95188]_  & \new_[95185]_ ;
  assign \new_[95190]_  = \new_[95189]_  & \new_[95182]_ ;
  assign \new_[95194]_  = A167 & ~A168;
  assign \new_[95195]_  = ~A169 & \new_[95194]_ ;
  assign \new_[95198]_  = A199 & A166;
  assign \new_[95201]_  = A201 & ~A200;
  assign \new_[95202]_  = \new_[95201]_  & \new_[95198]_ ;
  assign \new_[95203]_  = \new_[95202]_  & \new_[95195]_ ;
  assign \new_[95206]_  = ~A233 & A203;
  assign \new_[95209]_  = ~A266 & ~A234;
  assign \new_[95210]_  = \new_[95209]_  & \new_[95206]_ ;
  assign \new_[95213]_  = ~A269 & ~A268;
  assign \new_[95216]_  = A299 & A298;
  assign \new_[95217]_  = \new_[95216]_  & \new_[95213]_ ;
  assign \new_[95218]_  = \new_[95217]_  & \new_[95210]_ ;
  assign \new_[95222]_  = A167 & ~A168;
  assign \new_[95223]_  = ~A169 & \new_[95222]_ ;
  assign \new_[95226]_  = A199 & A166;
  assign \new_[95229]_  = A201 & ~A200;
  assign \new_[95230]_  = \new_[95229]_  & \new_[95226]_ ;
  assign \new_[95231]_  = \new_[95230]_  & \new_[95223]_ ;
  assign \new_[95234]_  = ~A233 & A203;
  assign \new_[95237]_  = ~A266 & ~A234;
  assign \new_[95238]_  = \new_[95237]_  & \new_[95234]_ ;
  assign \new_[95241]_  = ~A269 & ~A268;
  assign \new_[95244]_  = ~A299 & ~A298;
  assign \new_[95245]_  = \new_[95244]_  & \new_[95241]_ ;
  assign \new_[95246]_  = \new_[95245]_  & \new_[95238]_ ;
  assign \new_[95250]_  = A167 & ~A168;
  assign \new_[95251]_  = ~A169 & \new_[95250]_ ;
  assign \new_[95254]_  = A199 & A166;
  assign \new_[95257]_  = A201 & ~A200;
  assign \new_[95258]_  = \new_[95257]_  & \new_[95254]_ ;
  assign \new_[95259]_  = \new_[95258]_  & \new_[95251]_ ;
  assign \new_[95262]_  = ~A233 & A203;
  assign \new_[95265]_  = ~A266 & ~A234;
  assign \new_[95266]_  = \new_[95265]_  & \new_[95262]_ ;
  assign \new_[95269]_  = A298 & ~A267;
  assign \new_[95272]_  = ~A302 & ~A301;
  assign \new_[95273]_  = \new_[95272]_  & \new_[95269]_ ;
  assign \new_[95274]_  = \new_[95273]_  & \new_[95266]_ ;
  assign \new_[95278]_  = A167 & ~A168;
  assign \new_[95279]_  = ~A169 & \new_[95278]_ ;
  assign \new_[95282]_  = A199 & A166;
  assign \new_[95285]_  = A201 & ~A200;
  assign \new_[95286]_  = \new_[95285]_  & \new_[95282]_ ;
  assign \new_[95287]_  = \new_[95286]_  & \new_[95279]_ ;
  assign \new_[95290]_  = ~A233 & A203;
  assign \new_[95293]_  = ~A265 & ~A234;
  assign \new_[95294]_  = \new_[95293]_  & \new_[95290]_ ;
  assign \new_[95297]_  = A298 & ~A266;
  assign \new_[95300]_  = ~A302 & ~A301;
  assign \new_[95301]_  = \new_[95300]_  & \new_[95297]_ ;
  assign \new_[95302]_  = \new_[95301]_  & \new_[95294]_ ;
  assign \new_[95306]_  = A167 & ~A168;
  assign \new_[95307]_  = ~A169 & \new_[95306]_ ;
  assign \new_[95310]_  = A199 & A166;
  assign \new_[95313]_  = A201 & ~A200;
  assign \new_[95314]_  = \new_[95313]_  & \new_[95310]_ ;
  assign \new_[95315]_  = \new_[95314]_  & \new_[95307]_ ;
  assign \new_[95318]_  = ~A232 & A203;
  assign \new_[95321]_  = A265 & ~A233;
  assign \new_[95322]_  = \new_[95321]_  & \new_[95318]_ ;
  assign \new_[95325]_  = A298 & A266;
  assign \new_[95328]_  = ~A302 & ~A301;
  assign \new_[95329]_  = \new_[95328]_  & \new_[95325]_ ;
  assign \new_[95330]_  = \new_[95329]_  & \new_[95322]_ ;
  assign \new_[95334]_  = A167 & ~A168;
  assign \new_[95335]_  = ~A169 & \new_[95334]_ ;
  assign \new_[95338]_  = A199 & A166;
  assign \new_[95341]_  = A201 & ~A200;
  assign \new_[95342]_  = \new_[95341]_  & \new_[95338]_ ;
  assign \new_[95343]_  = \new_[95342]_  & \new_[95335]_ ;
  assign \new_[95346]_  = ~A232 & A203;
  assign \new_[95349]_  = ~A266 & ~A233;
  assign \new_[95350]_  = \new_[95349]_  & \new_[95346]_ ;
  assign \new_[95353]_  = ~A269 & ~A268;
  assign \new_[95356]_  = ~A300 & A298;
  assign \new_[95357]_  = \new_[95356]_  & \new_[95353]_ ;
  assign \new_[95358]_  = \new_[95357]_  & \new_[95350]_ ;
  assign \new_[95362]_  = A167 & ~A168;
  assign \new_[95363]_  = ~A169 & \new_[95362]_ ;
  assign \new_[95366]_  = A199 & A166;
  assign \new_[95369]_  = A201 & ~A200;
  assign \new_[95370]_  = \new_[95369]_  & \new_[95366]_ ;
  assign \new_[95371]_  = \new_[95370]_  & \new_[95363]_ ;
  assign \new_[95374]_  = ~A232 & A203;
  assign \new_[95377]_  = ~A266 & ~A233;
  assign \new_[95378]_  = \new_[95377]_  & \new_[95374]_ ;
  assign \new_[95381]_  = ~A269 & ~A268;
  assign \new_[95384]_  = A299 & A298;
  assign \new_[95385]_  = \new_[95384]_  & \new_[95381]_ ;
  assign \new_[95386]_  = \new_[95385]_  & \new_[95378]_ ;
  assign \new_[95390]_  = A167 & ~A168;
  assign \new_[95391]_  = ~A169 & \new_[95390]_ ;
  assign \new_[95394]_  = A199 & A166;
  assign \new_[95397]_  = A201 & ~A200;
  assign \new_[95398]_  = \new_[95397]_  & \new_[95394]_ ;
  assign \new_[95399]_  = \new_[95398]_  & \new_[95391]_ ;
  assign \new_[95402]_  = ~A232 & A203;
  assign \new_[95405]_  = ~A266 & ~A233;
  assign \new_[95406]_  = \new_[95405]_  & \new_[95402]_ ;
  assign \new_[95409]_  = ~A269 & ~A268;
  assign \new_[95412]_  = ~A299 & ~A298;
  assign \new_[95413]_  = \new_[95412]_  & \new_[95409]_ ;
  assign \new_[95414]_  = \new_[95413]_  & \new_[95406]_ ;
  assign \new_[95418]_  = A167 & ~A168;
  assign \new_[95419]_  = ~A169 & \new_[95418]_ ;
  assign \new_[95422]_  = A199 & A166;
  assign \new_[95425]_  = A201 & ~A200;
  assign \new_[95426]_  = \new_[95425]_  & \new_[95422]_ ;
  assign \new_[95427]_  = \new_[95426]_  & \new_[95419]_ ;
  assign \new_[95430]_  = ~A232 & A203;
  assign \new_[95433]_  = ~A266 & ~A233;
  assign \new_[95434]_  = \new_[95433]_  & \new_[95430]_ ;
  assign \new_[95437]_  = A298 & ~A267;
  assign \new_[95440]_  = ~A302 & ~A301;
  assign \new_[95441]_  = \new_[95440]_  & \new_[95437]_ ;
  assign \new_[95442]_  = \new_[95441]_  & \new_[95434]_ ;
  assign \new_[95446]_  = A167 & ~A168;
  assign \new_[95447]_  = ~A169 & \new_[95446]_ ;
  assign \new_[95450]_  = A199 & A166;
  assign \new_[95453]_  = A201 & ~A200;
  assign \new_[95454]_  = \new_[95453]_  & \new_[95450]_ ;
  assign \new_[95455]_  = \new_[95454]_  & \new_[95447]_ ;
  assign \new_[95458]_  = ~A232 & A203;
  assign \new_[95461]_  = ~A265 & ~A233;
  assign \new_[95462]_  = \new_[95461]_  & \new_[95458]_ ;
  assign \new_[95465]_  = A298 & ~A266;
  assign \new_[95468]_  = ~A302 & ~A301;
  assign \new_[95469]_  = \new_[95468]_  & \new_[95465]_ ;
  assign \new_[95470]_  = \new_[95469]_  & \new_[95462]_ ;
  assign \new_[95474]_  = A167 & ~A169;
  assign \new_[95475]_  = A170 & \new_[95474]_ ;
  assign \new_[95478]_  = A199 & ~A166;
  assign \new_[95481]_  = ~A233 & A200;
  assign \new_[95482]_  = \new_[95481]_  & \new_[95478]_ ;
  assign \new_[95483]_  = \new_[95482]_  & \new_[95475]_ ;
  assign \new_[95486]_  = ~A236 & ~A235;
  assign \new_[95489]_  = ~A268 & ~A266;
  assign \new_[95490]_  = \new_[95489]_  & \new_[95486]_ ;
  assign \new_[95493]_  = A298 & ~A269;
  assign \new_[95496]_  = ~A302 & ~A301;
  assign \new_[95497]_  = \new_[95496]_  & \new_[95493]_ ;
  assign \new_[95498]_  = \new_[95497]_  & \new_[95490]_ ;
  assign \new_[95502]_  = A167 & ~A169;
  assign \new_[95503]_  = A170 & \new_[95502]_ ;
  assign \new_[95506]_  = ~A200 & ~A166;
  assign \new_[95509]_  = ~A203 & ~A202;
  assign \new_[95510]_  = \new_[95509]_  & \new_[95506]_ ;
  assign \new_[95511]_  = \new_[95510]_  & \new_[95503]_ ;
  assign \new_[95514]_  = A233 & A232;
  assign \new_[95517]_  = ~A268 & A265;
  assign \new_[95518]_  = \new_[95517]_  & \new_[95514]_ ;
  assign \new_[95521]_  = ~A299 & ~A269;
  assign \new_[95524]_  = ~A302 & ~A301;
  assign \new_[95525]_  = \new_[95524]_  & \new_[95521]_ ;
  assign \new_[95526]_  = \new_[95525]_  & \new_[95518]_ ;
  assign \new_[95530]_  = A167 & ~A169;
  assign \new_[95531]_  = A170 & \new_[95530]_ ;
  assign \new_[95534]_  = ~A200 & ~A166;
  assign \new_[95537]_  = ~A203 & ~A202;
  assign \new_[95538]_  = \new_[95537]_  & \new_[95534]_ ;
  assign \new_[95539]_  = \new_[95538]_  & \new_[95531]_ ;
  assign \new_[95542]_  = ~A235 & ~A233;
  assign \new_[95545]_  = A265 & ~A236;
  assign \new_[95546]_  = \new_[95545]_  & \new_[95542]_ ;
  assign \new_[95549]_  = A298 & A266;
  assign \new_[95552]_  = ~A302 & ~A301;
  assign \new_[95553]_  = \new_[95552]_  & \new_[95549]_ ;
  assign \new_[95554]_  = \new_[95553]_  & \new_[95546]_ ;
  assign \new_[95558]_  = A167 & ~A169;
  assign \new_[95559]_  = A170 & \new_[95558]_ ;
  assign \new_[95562]_  = ~A200 & ~A166;
  assign \new_[95565]_  = ~A203 & ~A202;
  assign \new_[95566]_  = \new_[95565]_  & \new_[95562]_ ;
  assign \new_[95567]_  = \new_[95566]_  & \new_[95559]_ ;
  assign \new_[95570]_  = ~A235 & ~A233;
  assign \new_[95573]_  = ~A266 & ~A236;
  assign \new_[95574]_  = \new_[95573]_  & \new_[95570]_ ;
  assign \new_[95577]_  = ~A269 & ~A268;
  assign \new_[95580]_  = ~A300 & A298;
  assign \new_[95581]_  = \new_[95580]_  & \new_[95577]_ ;
  assign \new_[95582]_  = \new_[95581]_  & \new_[95574]_ ;
  assign \new_[95586]_  = A167 & ~A169;
  assign \new_[95587]_  = A170 & \new_[95586]_ ;
  assign \new_[95590]_  = ~A200 & ~A166;
  assign \new_[95593]_  = ~A203 & ~A202;
  assign \new_[95594]_  = \new_[95593]_  & \new_[95590]_ ;
  assign \new_[95595]_  = \new_[95594]_  & \new_[95587]_ ;
  assign \new_[95598]_  = ~A235 & ~A233;
  assign \new_[95601]_  = ~A266 & ~A236;
  assign \new_[95602]_  = \new_[95601]_  & \new_[95598]_ ;
  assign \new_[95605]_  = ~A269 & ~A268;
  assign \new_[95608]_  = A299 & A298;
  assign \new_[95609]_  = \new_[95608]_  & \new_[95605]_ ;
  assign \new_[95610]_  = \new_[95609]_  & \new_[95602]_ ;
  assign \new_[95614]_  = A167 & ~A169;
  assign \new_[95615]_  = A170 & \new_[95614]_ ;
  assign \new_[95618]_  = ~A200 & ~A166;
  assign \new_[95621]_  = ~A203 & ~A202;
  assign \new_[95622]_  = \new_[95621]_  & \new_[95618]_ ;
  assign \new_[95623]_  = \new_[95622]_  & \new_[95615]_ ;
  assign \new_[95626]_  = ~A235 & ~A233;
  assign \new_[95629]_  = ~A266 & ~A236;
  assign \new_[95630]_  = \new_[95629]_  & \new_[95626]_ ;
  assign \new_[95633]_  = ~A269 & ~A268;
  assign \new_[95636]_  = ~A299 & ~A298;
  assign \new_[95637]_  = \new_[95636]_  & \new_[95633]_ ;
  assign \new_[95638]_  = \new_[95637]_  & \new_[95630]_ ;
  assign \new_[95642]_  = A167 & ~A169;
  assign \new_[95643]_  = A170 & \new_[95642]_ ;
  assign \new_[95646]_  = ~A200 & ~A166;
  assign \new_[95649]_  = ~A203 & ~A202;
  assign \new_[95650]_  = \new_[95649]_  & \new_[95646]_ ;
  assign \new_[95651]_  = \new_[95650]_  & \new_[95643]_ ;
  assign \new_[95654]_  = ~A235 & ~A233;
  assign \new_[95657]_  = ~A266 & ~A236;
  assign \new_[95658]_  = \new_[95657]_  & \new_[95654]_ ;
  assign \new_[95661]_  = A298 & ~A267;
  assign \new_[95664]_  = ~A302 & ~A301;
  assign \new_[95665]_  = \new_[95664]_  & \new_[95661]_ ;
  assign \new_[95666]_  = \new_[95665]_  & \new_[95658]_ ;
  assign \new_[95670]_  = A167 & ~A169;
  assign \new_[95671]_  = A170 & \new_[95670]_ ;
  assign \new_[95674]_  = ~A200 & ~A166;
  assign \new_[95677]_  = ~A203 & ~A202;
  assign \new_[95678]_  = \new_[95677]_  & \new_[95674]_ ;
  assign \new_[95679]_  = \new_[95678]_  & \new_[95671]_ ;
  assign \new_[95682]_  = ~A235 & ~A233;
  assign \new_[95685]_  = ~A265 & ~A236;
  assign \new_[95686]_  = \new_[95685]_  & \new_[95682]_ ;
  assign \new_[95689]_  = A298 & ~A266;
  assign \new_[95692]_  = ~A302 & ~A301;
  assign \new_[95693]_  = \new_[95692]_  & \new_[95689]_ ;
  assign \new_[95694]_  = \new_[95693]_  & \new_[95686]_ ;
  assign \new_[95698]_  = A167 & ~A169;
  assign \new_[95699]_  = A170 & \new_[95698]_ ;
  assign \new_[95702]_  = ~A200 & ~A166;
  assign \new_[95705]_  = ~A203 & ~A202;
  assign \new_[95706]_  = \new_[95705]_  & \new_[95702]_ ;
  assign \new_[95707]_  = \new_[95706]_  & \new_[95699]_ ;
  assign \new_[95710]_  = ~A234 & ~A233;
  assign \new_[95713]_  = ~A268 & ~A266;
  assign \new_[95714]_  = \new_[95713]_  & \new_[95710]_ ;
  assign \new_[95717]_  = A298 & ~A269;
  assign \new_[95720]_  = ~A302 & ~A301;
  assign \new_[95721]_  = \new_[95720]_  & \new_[95717]_ ;
  assign \new_[95722]_  = \new_[95721]_  & \new_[95714]_ ;
  assign \new_[95726]_  = A167 & ~A169;
  assign \new_[95727]_  = A170 & \new_[95726]_ ;
  assign \new_[95730]_  = ~A200 & ~A166;
  assign \new_[95733]_  = ~A203 & ~A202;
  assign \new_[95734]_  = \new_[95733]_  & \new_[95730]_ ;
  assign \new_[95735]_  = \new_[95734]_  & \new_[95727]_ ;
  assign \new_[95738]_  = ~A233 & A232;
  assign \new_[95741]_  = A235 & A234;
  assign \new_[95742]_  = \new_[95741]_  & \new_[95738]_ ;
  assign \new_[95745]_  = ~A299 & A298;
  assign \new_[95748]_  = A301 & A300;
  assign \new_[95749]_  = \new_[95748]_  & \new_[95745]_ ;
  assign \new_[95750]_  = \new_[95749]_  & \new_[95742]_ ;
  assign \new_[95754]_  = A167 & ~A169;
  assign \new_[95755]_  = A170 & \new_[95754]_ ;
  assign \new_[95758]_  = ~A200 & ~A166;
  assign \new_[95761]_  = ~A203 & ~A202;
  assign \new_[95762]_  = \new_[95761]_  & \new_[95758]_ ;
  assign \new_[95763]_  = \new_[95762]_  & \new_[95755]_ ;
  assign \new_[95766]_  = ~A233 & A232;
  assign \new_[95769]_  = A235 & A234;
  assign \new_[95770]_  = \new_[95769]_  & \new_[95766]_ ;
  assign \new_[95773]_  = ~A299 & A298;
  assign \new_[95776]_  = A302 & A300;
  assign \new_[95777]_  = \new_[95776]_  & \new_[95773]_ ;
  assign \new_[95778]_  = \new_[95777]_  & \new_[95770]_ ;
  assign \new_[95782]_  = A167 & ~A169;
  assign \new_[95783]_  = A170 & \new_[95782]_ ;
  assign \new_[95786]_  = ~A200 & ~A166;
  assign \new_[95789]_  = ~A203 & ~A202;
  assign \new_[95790]_  = \new_[95789]_  & \new_[95786]_ ;
  assign \new_[95791]_  = \new_[95790]_  & \new_[95783]_ ;
  assign \new_[95794]_  = ~A233 & A232;
  assign \new_[95797]_  = A235 & A234;
  assign \new_[95798]_  = \new_[95797]_  & \new_[95794]_ ;
  assign \new_[95801]_  = ~A266 & A265;
  assign \new_[95804]_  = A268 & A267;
  assign \new_[95805]_  = \new_[95804]_  & \new_[95801]_ ;
  assign \new_[95806]_  = \new_[95805]_  & \new_[95798]_ ;
  assign \new_[95810]_  = A167 & ~A169;
  assign \new_[95811]_  = A170 & \new_[95810]_ ;
  assign \new_[95814]_  = ~A200 & ~A166;
  assign \new_[95817]_  = ~A203 & ~A202;
  assign \new_[95818]_  = \new_[95817]_  & \new_[95814]_ ;
  assign \new_[95819]_  = \new_[95818]_  & \new_[95811]_ ;
  assign \new_[95822]_  = ~A233 & A232;
  assign \new_[95825]_  = A235 & A234;
  assign \new_[95826]_  = \new_[95825]_  & \new_[95822]_ ;
  assign \new_[95829]_  = ~A266 & A265;
  assign \new_[95832]_  = A269 & A267;
  assign \new_[95833]_  = \new_[95832]_  & \new_[95829]_ ;
  assign \new_[95834]_  = \new_[95833]_  & \new_[95826]_ ;
  assign \new_[95838]_  = A167 & ~A169;
  assign \new_[95839]_  = A170 & \new_[95838]_ ;
  assign \new_[95842]_  = ~A200 & ~A166;
  assign \new_[95845]_  = ~A203 & ~A202;
  assign \new_[95846]_  = \new_[95845]_  & \new_[95842]_ ;
  assign \new_[95847]_  = \new_[95846]_  & \new_[95839]_ ;
  assign \new_[95850]_  = ~A233 & A232;
  assign \new_[95853]_  = A236 & A234;
  assign \new_[95854]_  = \new_[95853]_  & \new_[95850]_ ;
  assign \new_[95857]_  = ~A299 & A298;
  assign \new_[95860]_  = A301 & A300;
  assign \new_[95861]_  = \new_[95860]_  & \new_[95857]_ ;
  assign \new_[95862]_  = \new_[95861]_  & \new_[95854]_ ;
  assign \new_[95866]_  = A167 & ~A169;
  assign \new_[95867]_  = A170 & \new_[95866]_ ;
  assign \new_[95870]_  = ~A200 & ~A166;
  assign \new_[95873]_  = ~A203 & ~A202;
  assign \new_[95874]_  = \new_[95873]_  & \new_[95870]_ ;
  assign \new_[95875]_  = \new_[95874]_  & \new_[95867]_ ;
  assign \new_[95878]_  = ~A233 & A232;
  assign \new_[95881]_  = A236 & A234;
  assign \new_[95882]_  = \new_[95881]_  & \new_[95878]_ ;
  assign \new_[95885]_  = ~A299 & A298;
  assign \new_[95888]_  = A302 & A300;
  assign \new_[95889]_  = \new_[95888]_  & \new_[95885]_ ;
  assign \new_[95890]_  = \new_[95889]_  & \new_[95882]_ ;
  assign \new_[95894]_  = A167 & ~A169;
  assign \new_[95895]_  = A170 & \new_[95894]_ ;
  assign \new_[95898]_  = ~A200 & ~A166;
  assign \new_[95901]_  = ~A203 & ~A202;
  assign \new_[95902]_  = \new_[95901]_  & \new_[95898]_ ;
  assign \new_[95903]_  = \new_[95902]_  & \new_[95895]_ ;
  assign \new_[95906]_  = ~A233 & A232;
  assign \new_[95909]_  = A236 & A234;
  assign \new_[95910]_  = \new_[95909]_  & \new_[95906]_ ;
  assign \new_[95913]_  = ~A266 & A265;
  assign \new_[95916]_  = A268 & A267;
  assign \new_[95917]_  = \new_[95916]_  & \new_[95913]_ ;
  assign \new_[95918]_  = \new_[95917]_  & \new_[95910]_ ;
  assign \new_[95922]_  = A167 & ~A169;
  assign \new_[95923]_  = A170 & \new_[95922]_ ;
  assign \new_[95926]_  = ~A200 & ~A166;
  assign \new_[95929]_  = ~A203 & ~A202;
  assign \new_[95930]_  = \new_[95929]_  & \new_[95926]_ ;
  assign \new_[95931]_  = \new_[95930]_  & \new_[95923]_ ;
  assign \new_[95934]_  = ~A233 & A232;
  assign \new_[95937]_  = A236 & A234;
  assign \new_[95938]_  = \new_[95937]_  & \new_[95934]_ ;
  assign \new_[95941]_  = ~A266 & A265;
  assign \new_[95944]_  = A269 & A267;
  assign \new_[95945]_  = \new_[95944]_  & \new_[95941]_ ;
  assign \new_[95946]_  = \new_[95945]_  & \new_[95938]_ ;
  assign \new_[95950]_  = A167 & ~A169;
  assign \new_[95951]_  = A170 & \new_[95950]_ ;
  assign \new_[95954]_  = ~A200 & ~A166;
  assign \new_[95957]_  = ~A203 & ~A202;
  assign \new_[95958]_  = \new_[95957]_  & \new_[95954]_ ;
  assign \new_[95959]_  = \new_[95958]_  & \new_[95951]_ ;
  assign \new_[95962]_  = ~A233 & ~A232;
  assign \new_[95965]_  = ~A268 & ~A266;
  assign \new_[95966]_  = \new_[95965]_  & \new_[95962]_ ;
  assign \new_[95969]_  = A298 & ~A269;
  assign \new_[95972]_  = ~A302 & ~A301;
  assign \new_[95973]_  = \new_[95972]_  & \new_[95969]_ ;
  assign \new_[95974]_  = \new_[95973]_  & \new_[95966]_ ;
  assign \new_[95978]_  = A167 & ~A169;
  assign \new_[95979]_  = A170 & \new_[95978]_ ;
  assign \new_[95982]_  = ~A200 & ~A166;
  assign \new_[95985]_  = ~A233 & ~A201;
  assign \new_[95986]_  = \new_[95985]_  & \new_[95982]_ ;
  assign \new_[95987]_  = \new_[95986]_  & \new_[95979]_ ;
  assign \new_[95990]_  = ~A236 & ~A235;
  assign \new_[95993]_  = ~A268 & ~A266;
  assign \new_[95994]_  = \new_[95993]_  & \new_[95990]_ ;
  assign \new_[95997]_  = A298 & ~A269;
  assign \new_[96000]_  = ~A302 & ~A301;
  assign \new_[96001]_  = \new_[96000]_  & \new_[95997]_ ;
  assign \new_[96002]_  = \new_[96001]_  & \new_[95994]_ ;
  assign \new_[96006]_  = A167 & ~A169;
  assign \new_[96007]_  = A170 & \new_[96006]_ ;
  assign \new_[96010]_  = ~A199 & ~A166;
  assign \new_[96013]_  = ~A233 & ~A200;
  assign \new_[96014]_  = \new_[96013]_  & \new_[96010]_ ;
  assign \new_[96015]_  = \new_[96014]_  & \new_[96007]_ ;
  assign \new_[96018]_  = ~A236 & ~A235;
  assign \new_[96021]_  = ~A268 & ~A266;
  assign \new_[96022]_  = \new_[96021]_  & \new_[96018]_ ;
  assign \new_[96025]_  = A298 & ~A269;
  assign \new_[96028]_  = ~A302 & ~A301;
  assign \new_[96029]_  = \new_[96028]_  & \new_[96025]_ ;
  assign \new_[96030]_  = \new_[96029]_  & \new_[96022]_ ;
  assign \new_[96034]_  = ~A167 & ~A169;
  assign \new_[96035]_  = A170 & \new_[96034]_ ;
  assign \new_[96038]_  = A199 & A166;
  assign \new_[96041]_  = ~A233 & A200;
  assign \new_[96042]_  = \new_[96041]_  & \new_[96038]_ ;
  assign \new_[96043]_  = \new_[96042]_  & \new_[96035]_ ;
  assign \new_[96046]_  = ~A236 & ~A235;
  assign \new_[96049]_  = ~A268 & ~A266;
  assign \new_[96050]_  = \new_[96049]_  & \new_[96046]_ ;
  assign \new_[96053]_  = A298 & ~A269;
  assign \new_[96056]_  = ~A302 & ~A301;
  assign \new_[96057]_  = \new_[96056]_  & \new_[96053]_ ;
  assign \new_[96058]_  = \new_[96057]_  & \new_[96050]_ ;
  assign \new_[96062]_  = ~A167 & ~A169;
  assign \new_[96063]_  = A170 & \new_[96062]_ ;
  assign \new_[96066]_  = ~A200 & A166;
  assign \new_[96069]_  = ~A203 & ~A202;
  assign \new_[96070]_  = \new_[96069]_  & \new_[96066]_ ;
  assign \new_[96071]_  = \new_[96070]_  & \new_[96063]_ ;
  assign \new_[96074]_  = A233 & A232;
  assign \new_[96077]_  = ~A268 & A265;
  assign \new_[96078]_  = \new_[96077]_  & \new_[96074]_ ;
  assign \new_[96081]_  = ~A299 & ~A269;
  assign \new_[96084]_  = ~A302 & ~A301;
  assign \new_[96085]_  = \new_[96084]_  & \new_[96081]_ ;
  assign \new_[96086]_  = \new_[96085]_  & \new_[96078]_ ;
  assign \new_[96090]_  = ~A167 & ~A169;
  assign \new_[96091]_  = A170 & \new_[96090]_ ;
  assign \new_[96094]_  = ~A200 & A166;
  assign \new_[96097]_  = ~A203 & ~A202;
  assign \new_[96098]_  = \new_[96097]_  & \new_[96094]_ ;
  assign \new_[96099]_  = \new_[96098]_  & \new_[96091]_ ;
  assign \new_[96102]_  = ~A235 & ~A233;
  assign \new_[96105]_  = A265 & ~A236;
  assign \new_[96106]_  = \new_[96105]_  & \new_[96102]_ ;
  assign \new_[96109]_  = A298 & A266;
  assign \new_[96112]_  = ~A302 & ~A301;
  assign \new_[96113]_  = \new_[96112]_  & \new_[96109]_ ;
  assign \new_[96114]_  = \new_[96113]_  & \new_[96106]_ ;
  assign \new_[96118]_  = ~A167 & ~A169;
  assign \new_[96119]_  = A170 & \new_[96118]_ ;
  assign \new_[96122]_  = ~A200 & A166;
  assign \new_[96125]_  = ~A203 & ~A202;
  assign \new_[96126]_  = \new_[96125]_  & \new_[96122]_ ;
  assign \new_[96127]_  = \new_[96126]_  & \new_[96119]_ ;
  assign \new_[96130]_  = ~A235 & ~A233;
  assign \new_[96133]_  = ~A266 & ~A236;
  assign \new_[96134]_  = \new_[96133]_  & \new_[96130]_ ;
  assign \new_[96137]_  = ~A269 & ~A268;
  assign \new_[96140]_  = ~A300 & A298;
  assign \new_[96141]_  = \new_[96140]_  & \new_[96137]_ ;
  assign \new_[96142]_  = \new_[96141]_  & \new_[96134]_ ;
  assign \new_[96146]_  = ~A167 & ~A169;
  assign \new_[96147]_  = A170 & \new_[96146]_ ;
  assign \new_[96150]_  = ~A200 & A166;
  assign \new_[96153]_  = ~A203 & ~A202;
  assign \new_[96154]_  = \new_[96153]_  & \new_[96150]_ ;
  assign \new_[96155]_  = \new_[96154]_  & \new_[96147]_ ;
  assign \new_[96158]_  = ~A235 & ~A233;
  assign \new_[96161]_  = ~A266 & ~A236;
  assign \new_[96162]_  = \new_[96161]_  & \new_[96158]_ ;
  assign \new_[96165]_  = ~A269 & ~A268;
  assign \new_[96168]_  = A299 & A298;
  assign \new_[96169]_  = \new_[96168]_  & \new_[96165]_ ;
  assign \new_[96170]_  = \new_[96169]_  & \new_[96162]_ ;
  assign \new_[96174]_  = ~A167 & ~A169;
  assign \new_[96175]_  = A170 & \new_[96174]_ ;
  assign \new_[96178]_  = ~A200 & A166;
  assign \new_[96181]_  = ~A203 & ~A202;
  assign \new_[96182]_  = \new_[96181]_  & \new_[96178]_ ;
  assign \new_[96183]_  = \new_[96182]_  & \new_[96175]_ ;
  assign \new_[96186]_  = ~A235 & ~A233;
  assign \new_[96189]_  = ~A266 & ~A236;
  assign \new_[96190]_  = \new_[96189]_  & \new_[96186]_ ;
  assign \new_[96193]_  = ~A269 & ~A268;
  assign \new_[96196]_  = ~A299 & ~A298;
  assign \new_[96197]_  = \new_[96196]_  & \new_[96193]_ ;
  assign \new_[96198]_  = \new_[96197]_  & \new_[96190]_ ;
  assign \new_[96202]_  = ~A167 & ~A169;
  assign \new_[96203]_  = A170 & \new_[96202]_ ;
  assign \new_[96206]_  = ~A200 & A166;
  assign \new_[96209]_  = ~A203 & ~A202;
  assign \new_[96210]_  = \new_[96209]_  & \new_[96206]_ ;
  assign \new_[96211]_  = \new_[96210]_  & \new_[96203]_ ;
  assign \new_[96214]_  = ~A235 & ~A233;
  assign \new_[96217]_  = ~A266 & ~A236;
  assign \new_[96218]_  = \new_[96217]_  & \new_[96214]_ ;
  assign \new_[96221]_  = A298 & ~A267;
  assign \new_[96224]_  = ~A302 & ~A301;
  assign \new_[96225]_  = \new_[96224]_  & \new_[96221]_ ;
  assign \new_[96226]_  = \new_[96225]_  & \new_[96218]_ ;
  assign \new_[96230]_  = ~A167 & ~A169;
  assign \new_[96231]_  = A170 & \new_[96230]_ ;
  assign \new_[96234]_  = ~A200 & A166;
  assign \new_[96237]_  = ~A203 & ~A202;
  assign \new_[96238]_  = \new_[96237]_  & \new_[96234]_ ;
  assign \new_[96239]_  = \new_[96238]_  & \new_[96231]_ ;
  assign \new_[96242]_  = ~A235 & ~A233;
  assign \new_[96245]_  = ~A265 & ~A236;
  assign \new_[96246]_  = \new_[96245]_  & \new_[96242]_ ;
  assign \new_[96249]_  = A298 & ~A266;
  assign \new_[96252]_  = ~A302 & ~A301;
  assign \new_[96253]_  = \new_[96252]_  & \new_[96249]_ ;
  assign \new_[96254]_  = \new_[96253]_  & \new_[96246]_ ;
  assign \new_[96258]_  = ~A167 & ~A169;
  assign \new_[96259]_  = A170 & \new_[96258]_ ;
  assign \new_[96262]_  = ~A200 & A166;
  assign \new_[96265]_  = ~A203 & ~A202;
  assign \new_[96266]_  = \new_[96265]_  & \new_[96262]_ ;
  assign \new_[96267]_  = \new_[96266]_  & \new_[96259]_ ;
  assign \new_[96270]_  = ~A234 & ~A233;
  assign \new_[96273]_  = ~A268 & ~A266;
  assign \new_[96274]_  = \new_[96273]_  & \new_[96270]_ ;
  assign \new_[96277]_  = A298 & ~A269;
  assign \new_[96280]_  = ~A302 & ~A301;
  assign \new_[96281]_  = \new_[96280]_  & \new_[96277]_ ;
  assign \new_[96282]_  = \new_[96281]_  & \new_[96274]_ ;
  assign \new_[96286]_  = ~A167 & ~A169;
  assign \new_[96287]_  = A170 & \new_[96286]_ ;
  assign \new_[96290]_  = ~A200 & A166;
  assign \new_[96293]_  = ~A203 & ~A202;
  assign \new_[96294]_  = \new_[96293]_  & \new_[96290]_ ;
  assign \new_[96295]_  = \new_[96294]_  & \new_[96287]_ ;
  assign \new_[96298]_  = ~A233 & A232;
  assign \new_[96301]_  = A235 & A234;
  assign \new_[96302]_  = \new_[96301]_  & \new_[96298]_ ;
  assign \new_[96305]_  = ~A299 & A298;
  assign \new_[96308]_  = A301 & A300;
  assign \new_[96309]_  = \new_[96308]_  & \new_[96305]_ ;
  assign \new_[96310]_  = \new_[96309]_  & \new_[96302]_ ;
  assign \new_[96314]_  = ~A167 & ~A169;
  assign \new_[96315]_  = A170 & \new_[96314]_ ;
  assign \new_[96318]_  = ~A200 & A166;
  assign \new_[96321]_  = ~A203 & ~A202;
  assign \new_[96322]_  = \new_[96321]_  & \new_[96318]_ ;
  assign \new_[96323]_  = \new_[96322]_  & \new_[96315]_ ;
  assign \new_[96326]_  = ~A233 & A232;
  assign \new_[96329]_  = A235 & A234;
  assign \new_[96330]_  = \new_[96329]_  & \new_[96326]_ ;
  assign \new_[96333]_  = ~A299 & A298;
  assign \new_[96336]_  = A302 & A300;
  assign \new_[96337]_  = \new_[96336]_  & \new_[96333]_ ;
  assign \new_[96338]_  = \new_[96337]_  & \new_[96330]_ ;
  assign \new_[96342]_  = ~A167 & ~A169;
  assign \new_[96343]_  = A170 & \new_[96342]_ ;
  assign \new_[96346]_  = ~A200 & A166;
  assign \new_[96349]_  = ~A203 & ~A202;
  assign \new_[96350]_  = \new_[96349]_  & \new_[96346]_ ;
  assign \new_[96351]_  = \new_[96350]_  & \new_[96343]_ ;
  assign \new_[96354]_  = ~A233 & A232;
  assign \new_[96357]_  = A235 & A234;
  assign \new_[96358]_  = \new_[96357]_  & \new_[96354]_ ;
  assign \new_[96361]_  = ~A266 & A265;
  assign \new_[96364]_  = A268 & A267;
  assign \new_[96365]_  = \new_[96364]_  & \new_[96361]_ ;
  assign \new_[96366]_  = \new_[96365]_  & \new_[96358]_ ;
  assign \new_[96370]_  = ~A167 & ~A169;
  assign \new_[96371]_  = A170 & \new_[96370]_ ;
  assign \new_[96374]_  = ~A200 & A166;
  assign \new_[96377]_  = ~A203 & ~A202;
  assign \new_[96378]_  = \new_[96377]_  & \new_[96374]_ ;
  assign \new_[96379]_  = \new_[96378]_  & \new_[96371]_ ;
  assign \new_[96382]_  = ~A233 & A232;
  assign \new_[96385]_  = A235 & A234;
  assign \new_[96386]_  = \new_[96385]_  & \new_[96382]_ ;
  assign \new_[96389]_  = ~A266 & A265;
  assign \new_[96392]_  = A269 & A267;
  assign \new_[96393]_  = \new_[96392]_  & \new_[96389]_ ;
  assign \new_[96394]_  = \new_[96393]_  & \new_[96386]_ ;
  assign \new_[96398]_  = ~A167 & ~A169;
  assign \new_[96399]_  = A170 & \new_[96398]_ ;
  assign \new_[96402]_  = ~A200 & A166;
  assign \new_[96405]_  = ~A203 & ~A202;
  assign \new_[96406]_  = \new_[96405]_  & \new_[96402]_ ;
  assign \new_[96407]_  = \new_[96406]_  & \new_[96399]_ ;
  assign \new_[96410]_  = ~A233 & A232;
  assign \new_[96413]_  = A236 & A234;
  assign \new_[96414]_  = \new_[96413]_  & \new_[96410]_ ;
  assign \new_[96417]_  = ~A299 & A298;
  assign \new_[96420]_  = A301 & A300;
  assign \new_[96421]_  = \new_[96420]_  & \new_[96417]_ ;
  assign \new_[96422]_  = \new_[96421]_  & \new_[96414]_ ;
  assign \new_[96426]_  = ~A167 & ~A169;
  assign \new_[96427]_  = A170 & \new_[96426]_ ;
  assign \new_[96430]_  = ~A200 & A166;
  assign \new_[96433]_  = ~A203 & ~A202;
  assign \new_[96434]_  = \new_[96433]_  & \new_[96430]_ ;
  assign \new_[96435]_  = \new_[96434]_  & \new_[96427]_ ;
  assign \new_[96438]_  = ~A233 & A232;
  assign \new_[96441]_  = A236 & A234;
  assign \new_[96442]_  = \new_[96441]_  & \new_[96438]_ ;
  assign \new_[96445]_  = ~A299 & A298;
  assign \new_[96448]_  = A302 & A300;
  assign \new_[96449]_  = \new_[96448]_  & \new_[96445]_ ;
  assign \new_[96450]_  = \new_[96449]_  & \new_[96442]_ ;
  assign \new_[96454]_  = ~A167 & ~A169;
  assign \new_[96455]_  = A170 & \new_[96454]_ ;
  assign \new_[96458]_  = ~A200 & A166;
  assign \new_[96461]_  = ~A203 & ~A202;
  assign \new_[96462]_  = \new_[96461]_  & \new_[96458]_ ;
  assign \new_[96463]_  = \new_[96462]_  & \new_[96455]_ ;
  assign \new_[96466]_  = ~A233 & A232;
  assign \new_[96469]_  = A236 & A234;
  assign \new_[96470]_  = \new_[96469]_  & \new_[96466]_ ;
  assign \new_[96473]_  = ~A266 & A265;
  assign \new_[96476]_  = A268 & A267;
  assign \new_[96477]_  = \new_[96476]_  & \new_[96473]_ ;
  assign \new_[96478]_  = \new_[96477]_  & \new_[96470]_ ;
  assign \new_[96482]_  = ~A167 & ~A169;
  assign \new_[96483]_  = A170 & \new_[96482]_ ;
  assign \new_[96486]_  = ~A200 & A166;
  assign \new_[96489]_  = ~A203 & ~A202;
  assign \new_[96490]_  = \new_[96489]_  & \new_[96486]_ ;
  assign \new_[96491]_  = \new_[96490]_  & \new_[96483]_ ;
  assign \new_[96494]_  = ~A233 & A232;
  assign \new_[96497]_  = A236 & A234;
  assign \new_[96498]_  = \new_[96497]_  & \new_[96494]_ ;
  assign \new_[96501]_  = ~A266 & A265;
  assign \new_[96504]_  = A269 & A267;
  assign \new_[96505]_  = \new_[96504]_  & \new_[96501]_ ;
  assign \new_[96506]_  = \new_[96505]_  & \new_[96498]_ ;
  assign \new_[96510]_  = ~A167 & ~A169;
  assign \new_[96511]_  = A170 & \new_[96510]_ ;
  assign \new_[96514]_  = ~A200 & A166;
  assign \new_[96517]_  = ~A203 & ~A202;
  assign \new_[96518]_  = \new_[96517]_  & \new_[96514]_ ;
  assign \new_[96519]_  = \new_[96518]_  & \new_[96511]_ ;
  assign \new_[96522]_  = ~A233 & ~A232;
  assign \new_[96525]_  = ~A268 & ~A266;
  assign \new_[96526]_  = \new_[96525]_  & \new_[96522]_ ;
  assign \new_[96529]_  = A298 & ~A269;
  assign \new_[96532]_  = ~A302 & ~A301;
  assign \new_[96533]_  = \new_[96532]_  & \new_[96529]_ ;
  assign \new_[96534]_  = \new_[96533]_  & \new_[96526]_ ;
  assign \new_[96538]_  = ~A167 & ~A169;
  assign \new_[96539]_  = A170 & \new_[96538]_ ;
  assign \new_[96542]_  = ~A200 & A166;
  assign \new_[96545]_  = ~A233 & ~A201;
  assign \new_[96546]_  = \new_[96545]_  & \new_[96542]_ ;
  assign \new_[96547]_  = \new_[96546]_  & \new_[96539]_ ;
  assign \new_[96550]_  = ~A236 & ~A235;
  assign \new_[96553]_  = ~A268 & ~A266;
  assign \new_[96554]_  = \new_[96553]_  & \new_[96550]_ ;
  assign \new_[96557]_  = A298 & ~A269;
  assign \new_[96560]_  = ~A302 & ~A301;
  assign \new_[96561]_  = \new_[96560]_  & \new_[96557]_ ;
  assign \new_[96562]_  = \new_[96561]_  & \new_[96554]_ ;
  assign \new_[96566]_  = ~A167 & ~A169;
  assign \new_[96567]_  = A170 & \new_[96566]_ ;
  assign \new_[96570]_  = ~A199 & A166;
  assign \new_[96573]_  = ~A233 & ~A200;
  assign \new_[96574]_  = \new_[96573]_  & \new_[96570]_ ;
  assign \new_[96575]_  = \new_[96574]_  & \new_[96567]_ ;
  assign \new_[96578]_  = ~A236 & ~A235;
  assign \new_[96581]_  = ~A268 & ~A266;
  assign \new_[96582]_  = \new_[96581]_  & \new_[96578]_ ;
  assign \new_[96585]_  = A298 & ~A269;
  assign \new_[96588]_  = ~A302 & ~A301;
  assign \new_[96589]_  = \new_[96588]_  & \new_[96585]_ ;
  assign \new_[96590]_  = \new_[96589]_  & \new_[96582]_ ;
  assign \new_[96594]_  = ~A168 & ~A169;
  assign \new_[96595]_  = ~A170 & \new_[96594]_ ;
  assign \new_[96598]_  = ~A200 & A199;
  assign \new_[96601]_  = A202 & A201;
  assign \new_[96602]_  = \new_[96601]_  & \new_[96598]_ ;
  assign \new_[96603]_  = \new_[96602]_  & \new_[96595]_ ;
  assign \new_[96606]_  = A233 & A232;
  assign \new_[96609]_  = ~A268 & A265;
  assign \new_[96610]_  = \new_[96609]_  & \new_[96606]_ ;
  assign \new_[96613]_  = ~A299 & ~A269;
  assign \new_[96616]_  = ~A302 & ~A301;
  assign \new_[96617]_  = \new_[96616]_  & \new_[96613]_ ;
  assign \new_[96618]_  = \new_[96617]_  & \new_[96610]_ ;
  assign \new_[96622]_  = ~A168 & ~A169;
  assign \new_[96623]_  = ~A170 & \new_[96622]_ ;
  assign \new_[96626]_  = ~A200 & A199;
  assign \new_[96629]_  = A202 & A201;
  assign \new_[96630]_  = \new_[96629]_  & \new_[96626]_ ;
  assign \new_[96631]_  = \new_[96630]_  & \new_[96623]_ ;
  assign \new_[96634]_  = ~A235 & ~A233;
  assign \new_[96637]_  = A265 & ~A236;
  assign \new_[96638]_  = \new_[96637]_  & \new_[96634]_ ;
  assign \new_[96641]_  = A298 & A266;
  assign \new_[96644]_  = ~A302 & ~A301;
  assign \new_[96645]_  = \new_[96644]_  & \new_[96641]_ ;
  assign \new_[96646]_  = \new_[96645]_  & \new_[96638]_ ;
  assign \new_[96650]_  = ~A168 & ~A169;
  assign \new_[96651]_  = ~A170 & \new_[96650]_ ;
  assign \new_[96654]_  = ~A200 & A199;
  assign \new_[96657]_  = A202 & A201;
  assign \new_[96658]_  = \new_[96657]_  & \new_[96654]_ ;
  assign \new_[96659]_  = \new_[96658]_  & \new_[96651]_ ;
  assign \new_[96662]_  = ~A235 & ~A233;
  assign \new_[96665]_  = ~A266 & ~A236;
  assign \new_[96666]_  = \new_[96665]_  & \new_[96662]_ ;
  assign \new_[96669]_  = ~A269 & ~A268;
  assign \new_[96672]_  = ~A300 & A298;
  assign \new_[96673]_  = \new_[96672]_  & \new_[96669]_ ;
  assign \new_[96674]_  = \new_[96673]_  & \new_[96666]_ ;
  assign \new_[96678]_  = ~A168 & ~A169;
  assign \new_[96679]_  = ~A170 & \new_[96678]_ ;
  assign \new_[96682]_  = ~A200 & A199;
  assign \new_[96685]_  = A202 & A201;
  assign \new_[96686]_  = \new_[96685]_  & \new_[96682]_ ;
  assign \new_[96687]_  = \new_[96686]_  & \new_[96679]_ ;
  assign \new_[96690]_  = ~A235 & ~A233;
  assign \new_[96693]_  = ~A266 & ~A236;
  assign \new_[96694]_  = \new_[96693]_  & \new_[96690]_ ;
  assign \new_[96697]_  = ~A269 & ~A268;
  assign \new_[96700]_  = A299 & A298;
  assign \new_[96701]_  = \new_[96700]_  & \new_[96697]_ ;
  assign \new_[96702]_  = \new_[96701]_  & \new_[96694]_ ;
  assign \new_[96706]_  = ~A168 & ~A169;
  assign \new_[96707]_  = ~A170 & \new_[96706]_ ;
  assign \new_[96710]_  = ~A200 & A199;
  assign \new_[96713]_  = A202 & A201;
  assign \new_[96714]_  = \new_[96713]_  & \new_[96710]_ ;
  assign \new_[96715]_  = \new_[96714]_  & \new_[96707]_ ;
  assign \new_[96718]_  = ~A235 & ~A233;
  assign \new_[96721]_  = ~A266 & ~A236;
  assign \new_[96722]_  = \new_[96721]_  & \new_[96718]_ ;
  assign \new_[96725]_  = ~A269 & ~A268;
  assign \new_[96728]_  = ~A299 & ~A298;
  assign \new_[96729]_  = \new_[96728]_  & \new_[96725]_ ;
  assign \new_[96730]_  = \new_[96729]_  & \new_[96722]_ ;
  assign \new_[96734]_  = ~A168 & ~A169;
  assign \new_[96735]_  = ~A170 & \new_[96734]_ ;
  assign \new_[96738]_  = ~A200 & A199;
  assign \new_[96741]_  = A202 & A201;
  assign \new_[96742]_  = \new_[96741]_  & \new_[96738]_ ;
  assign \new_[96743]_  = \new_[96742]_  & \new_[96735]_ ;
  assign \new_[96746]_  = ~A235 & ~A233;
  assign \new_[96749]_  = ~A266 & ~A236;
  assign \new_[96750]_  = \new_[96749]_  & \new_[96746]_ ;
  assign \new_[96753]_  = A298 & ~A267;
  assign \new_[96756]_  = ~A302 & ~A301;
  assign \new_[96757]_  = \new_[96756]_  & \new_[96753]_ ;
  assign \new_[96758]_  = \new_[96757]_  & \new_[96750]_ ;
  assign \new_[96762]_  = ~A168 & ~A169;
  assign \new_[96763]_  = ~A170 & \new_[96762]_ ;
  assign \new_[96766]_  = ~A200 & A199;
  assign \new_[96769]_  = A202 & A201;
  assign \new_[96770]_  = \new_[96769]_  & \new_[96766]_ ;
  assign \new_[96771]_  = \new_[96770]_  & \new_[96763]_ ;
  assign \new_[96774]_  = ~A235 & ~A233;
  assign \new_[96777]_  = ~A265 & ~A236;
  assign \new_[96778]_  = \new_[96777]_  & \new_[96774]_ ;
  assign \new_[96781]_  = A298 & ~A266;
  assign \new_[96784]_  = ~A302 & ~A301;
  assign \new_[96785]_  = \new_[96784]_  & \new_[96781]_ ;
  assign \new_[96786]_  = \new_[96785]_  & \new_[96778]_ ;
  assign \new_[96790]_  = ~A168 & ~A169;
  assign \new_[96791]_  = ~A170 & \new_[96790]_ ;
  assign \new_[96794]_  = ~A200 & A199;
  assign \new_[96797]_  = A202 & A201;
  assign \new_[96798]_  = \new_[96797]_  & \new_[96794]_ ;
  assign \new_[96799]_  = \new_[96798]_  & \new_[96791]_ ;
  assign \new_[96802]_  = ~A234 & ~A233;
  assign \new_[96805]_  = ~A268 & ~A266;
  assign \new_[96806]_  = \new_[96805]_  & \new_[96802]_ ;
  assign \new_[96809]_  = A298 & ~A269;
  assign \new_[96812]_  = ~A302 & ~A301;
  assign \new_[96813]_  = \new_[96812]_  & \new_[96809]_ ;
  assign \new_[96814]_  = \new_[96813]_  & \new_[96806]_ ;
  assign \new_[96818]_  = ~A168 & ~A169;
  assign \new_[96819]_  = ~A170 & \new_[96818]_ ;
  assign \new_[96822]_  = ~A200 & A199;
  assign \new_[96825]_  = A202 & A201;
  assign \new_[96826]_  = \new_[96825]_  & \new_[96822]_ ;
  assign \new_[96827]_  = \new_[96826]_  & \new_[96819]_ ;
  assign \new_[96830]_  = ~A233 & A232;
  assign \new_[96833]_  = A235 & A234;
  assign \new_[96834]_  = \new_[96833]_  & \new_[96830]_ ;
  assign \new_[96837]_  = ~A299 & A298;
  assign \new_[96840]_  = A301 & A300;
  assign \new_[96841]_  = \new_[96840]_  & \new_[96837]_ ;
  assign \new_[96842]_  = \new_[96841]_  & \new_[96834]_ ;
  assign \new_[96846]_  = ~A168 & ~A169;
  assign \new_[96847]_  = ~A170 & \new_[96846]_ ;
  assign \new_[96850]_  = ~A200 & A199;
  assign \new_[96853]_  = A202 & A201;
  assign \new_[96854]_  = \new_[96853]_  & \new_[96850]_ ;
  assign \new_[96855]_  = \new_[96854]_  & \new_[96847]_ ;
  assign \new_[96858]_  = ~A233 & A232;
  assign \new_[96861]_  = A235 & A234;
  assign \new_[96862]_  = \new_[96861]_  & \new_[96858]_ ;
  assign \new_[96865]_  = ~A299 & A298;
  assign \new_[96868]_  = A302 & A300;
  assign \new_[96869]_  = \new_[96868]_  & \new_[96865]_ ;
  assign \new_[96870]_  = \new_[96869]_  & \new_[96862]_ ;
  assign \new_[96874]_  = ~A168 & ~A169;
  assign \new_[96875]_  = ~A170 & \new_[96874]_ ;
  assign \new_[96878]_  = ~A200 & A199;
  assign \new_[96881]_  = A202 & A201;
  assign \new_[96882]_  = \new_[96881]_  & \new_[96878]_ ;
  assign \new_[96883]_  = \new_[96882]_  & \new_[96875]_ ;
  assign \new_[96886]_  = ~A233 & A232;
  assign \new_[96889]_  = A235 & A234;
  assign \new_[96890]_  = \new_[96889]_  & \new_[96886]_ ;
  assign \new_[96893]_  = ~A266 & A265;
  assign \new_[96896]_  = A268 & A267;
  assign \new_[96897]_  = \new_[96896]_  & \new_[96893]_ ;
  assign \new_[96898]_  = \new_[96897]_  & \new_[96890]_ ;
  assign \new_[96902]_  = ~A168 & ~A169;
  assign \new_[96903]_  = ~A170 & \new_[96902]_ ;
  assign \new_[96906]_  = ~A200 & A199;
  assign \new_[96909]_  = A202 & A201;
  assign \new_[96910]_  = \new_[96909]_  & \new_[96906]_ ;
  assign \new_[96911]_  = \new_[96910]_  & \new_[96903]_ ;
  assign \new_[96914]_  = ~A233 & A232;
  assign \new_[96917]_  = A235 & A234;
  assign \new_[96918]_  = \new_[96917]_  & \new_[96914]_ ;
  assign \new_[96921]_  = ~A266 & A265;
  assign \new_[96924]_  = A269 & A267;
  assign \new_[96925]_  = \new_[96924]_  & \new_[96921]_ ;
  assign \new_[96926]_  = \new_[96925]_  & \new_[96918]_ ;
  assign \new_[96930]_  = ~A168 & ~A169;
  assign \new_[96931]_  = ~A170 & \new_[96930]_ ;
  assign \new_[96934]_  = ~A200 & A199;
  assign \new_[96937]_  = A202 & A201;
  assign \new_[96938]_  = \new_[96937]_  & \new_[96934]_ ;
  assign \new_[96939]_  = \new_[96938]_  & \new_[96931]_ ;
  assign \new_[96942]_  = ~A233 & A232;
  assign \new_[96945]_  = A236 & A234;
  assign \new_[96946]_  = \new_[96945]_  & \new_[96942]_ ;
  assign \new_[96949]_  = ~A299 & A298;
  assign \new_[96952]_  = A301 & A300;
  assign \new_[96953]_  = \new_[96952]_  & \new_[96949]_ ;
  assign \new_[96954]_  = \new_[96953]_  & \new_[96946]_ ;
  assign \new_[96958]_  = ~A168 & ~A169;
  assign \new_[96959]_  = ~A170 & \new_[96958]_ ;
  assign \new_[96962]_  = ~A200 & A199;
  assign \new_[96965]_  = A202 & A201;
  assign \new_[96966]_  = \new_[96965]_  & \new_[96962]_ ;
  assign \new_[96967]_  = \new_[96966]_  & \new_[96959]_ ;
  assign \new_[96970]_  = ~A233 & A232;
  assign \new_[96973]_  = A236 & A234;
  assign \new_[96974]_  = \new_[96973]_  & \new_[96970]_ ;
  assign \new_[96977]_  = ~A299 & A298;
  assign \new_[96980]_  = A302 & A300;
  assign \new_[96981]_  = \new_[96980]_  & \new_[96977]_ ;
  assign \new_[96982]_  = \new_[96981]_  & \new_[96974]_ ;
  assign \new_[96986]_  = ~A168 & ~A169;
  assign \new_[96987]_  = ~A170 & \new_[96986]_ ;
  assign \new_[96990]_  = ~A200 & A199;
  assign \new_[96993]_  = A202 & A201;
  assign \new_[96994]_  = \new_[96993]_  & \new_[96990]_ ;
  assign \new_[96995]_  = \new_[96994]_  & \new_[96987]_ ;
  assign \new_[96998]_  = ~A233 & A232;
  assign \new_[97001]_  = A236 & A234;
  assign \new_[97002]_  = \new_[97001]_  & \new_[96998]_ ;
  assign \new_[97005]_  = ~A266 & A265;
  assign \new_[97008]_  = A268 & A267;
  assign \new_[97009]_  = \new_[97008]_  & \new_[97005]_ ;
  assign \new_[97010]_  = \new_[97009]_  & \new_[97002]_ ;
  assign \new_[97014]_  = ~A168 & ~A169;
  assign \new_[97015]_  = ~A170 & \new_[97014]_ ;
  assign \new_[97018]_  = ~A200 & A199;
  assign \new_[97021]_  = A202 & A201;
  assign \new_[97022]_  = \new_[97021]_  & \new_[97018]_ ;
  assign \new_[97023]_  = \new_[97022]_  & \new_[97015]_ ;
  assign \new_[97026]_  = ~A233 & A232;
  assign \new_[97029]_  = A236 & A234;
  assign \new_[97030]_  = \new_[97029]_  & \new_[97026]_ ;
  assign \new_[97033]_  = ~A266 & A265;
  assign \new_[97036]_  = A269 & A267;
  assign \new_[97037]_  = \new_[97036]_  & \new_[97033]_ ;
  assign \new_[97038]_  = \new_[97037]_  & \new_[97030]_ ;
  assign \new_[97042]_  = ~A168 & ~A169;
  assign \new_[97043]_  = ~A170 & \new_[97042]_ ;
  assign \new_[97046]_  = ~A200 & A199;
  assign \new_[97049]_  = A202 & A201;
  assign \new_[97050]_  = \new_[97049]_  & \new_[97046]_ ;
  assign \new_[97051]_  = \new_[97050]_  & \new_[97043]_ ;
  assign \new_[97054]_  = ~A233 & ~A232;
  assign \new_[97057]_  = ~A268 & ~A266;
  assign \new_[97058]_  = \new_[97057]_  & \new_[97054]_ ;
  assign \new_[97061]_  = A298 & ~A269;
  assign \new_[97064]_  = ~A302 & ~A301;
  assign \new_[97065]_  = \new_[97064]_  & \new_[97061]_ ;
  assign \new_[97066]_  = \new_[97065]_  & \new_[97058]_ ;
  assign \new_[97070]_  = ~A168 & ~A169;
  assign \new_[97071]_  = ~A170 & \new_[97070]_ ;
  assign \new_[97074]_  = ~A200 & A199;
  assign \new_[97077]_  = A203 & A201;
  assign \new_[97078]_  = \new_[97077]_  & \new_[97074]_ ;
  assign \new_[97079]_  = \new_[97078]_  & \new_[97071]_ ;
  assign \new_[97082]_  = A233 & A232;
  assign \new_[97085]_  = ~A268 & A265;
  assign \new_[97086]_  = \new_[97085]_  & \new_[97082]_ ;
  assign \new_[97089]_  = ~A299 & ~A269;
  assign \new_[97092]_  = ~A302 & ~A301;
  assign \new_[97093]_  = \new_[97092]_  & \new_[97089]_ ;
  assign \new_[97094]_  = \new_[97093]_  & \new_[97086]_ ;
  assign \new_[97098]_  = ~A168 & ~A169;
  assign \new_[97099]_  = ~A170 & \new_[97098]_ ;
  assign \new_[97102]_  = ~A200 & A199;
  assign \new_[97105]_  = A203 & A201;
  assign \new_[97106]_  = \new_[97105]_  & \new_[97102]_ ;
  assign \new_[97107]_  = \new_[97106]_  & \new_[97099]_ ;
  assign \new_[97110]_  = ~A235 & ~A233;
  assign \new_[97113]_  = A265 & ~A236;
  assign \new_[97114]_  = \new_[97113]_  & \new_[97110]_ ;
  assign \new_[97117]_  = A298 & A266;
  assign \new_[97120]_  = ~A302 & ~A301;
  assign \new_[97121]_  = \new_[97120]_  & \new_[97117]_ ;
  assign \new_[97122]_  = \new_[97121]_  & \new_[97114]_ ;
  assign \new_[97126]_  = ~A168 & ~A169;
  assign \new_[97127]_  = ~A170 & \new_[97126]_ ;
  assign \new_[97130]_  = ~A200 & A199;
  assign \new_[97133]_  = A203 & A201;
  assign \new_[97134]_  = \new_[97133]_  & \new_[97130]_ ;
  assign \new_[97135]_  = \new_[97134]_  & \new_[97127]_ ;
  assign \new_[97138]_  = ~A235 & ~A233;
  assign \new_[97141]_  = ~A266 & ~A236;
  assign \new_[97142]_  = \new_[97141]_  & \new_[97138]_ ;
  assign \new_[97145]_  = ~A269 & ~A268;
  assign \new_[97148]_  = ~A300 & A298;
  assign \new_[97149]_  = \new_[97148]_  & \new_[97145]_ ;
  assign \new_[97150]_  = \new_[97149]_  & \new_[97142]_ ;
  assign \new_[97154]_  = ~A168 & ~A169;
  assign \new_[97155]_  = ~A170 & \new_[97154]_ ;
  assign \new_[97158]_  = ~A200 & A199;
  assign \new_[97161]_  = A203 & A201;
  assign \new_[97162]_  = \new_[97161]_  & \new_[97158]_ ;
  assign \new_[97163]_  = \new_[97162]_  & \new_[97155]_ ;
  assign \new_[97166]_  = ~A235 & ~A233;
  assign \new_[97169]_  = ~A266 & ~A236;
  assign \new_[97170]_  = \new_[97169]_  & \new_[97166]_ ;
  assign \new_[97173]_  = ~A269 & ~A268;
  assign \new_[97176]_  = A299 & A298;
  assign \new_[97177]_  = \new_[97176]_  & \new_[97173]_ ;
  assign \new_[97178]_  = \new_[97177]_  & \new_[97170]_ ;
  assign \new_[97182]_  = ~A168 & ~A169;
  assign \new_[97183]_  = ~A170 & \new_[97182]_ ;
  assign \new_[97186]_  = ~A200 & A199;
  assign \new_[97189]_  = A203 & A201;
  assign \new_[97190]_  = \new_[97189]_  & \new_[97186]_ ;
  assign \new_[97191]_  = \new_[97190]_  & \new_[97183]_ ;
  assign \new_[97194]_  = ~A235 & ~A233;
  assign \new_[97197]_  = ~A266 & ~A236;
  assign \new_[97198]_  = \new_[97197]_  & \new_[97194]_ ;
  assign \new_[97201]_  = ~A269 & ~A268;
  assign \new_[97204]_  = ~A299 & ~A298;
  assign \new_[97205]_  = \new_[97204]_  & \new_[97201]_ ;
  assign \new_[97206]_  = \new_[97205]_  & \new_[97198]_ ;
  assign \new_[97210]_  = ~A168 & ~A169;
  assign \new_[97211]_  = ~A170 & \new_[97210]_ ;
  assign \new_[97214]_  = ~A200 & A199;
  assign \new_[97217]_  = A203 & A201;
  assign \new_[97218]_  = \new_[97217]_  & \new_[97214]_ ;
  assign \new_[97219]_  = \new_[97218]_  & \new_[97211]_ ;
  assign \new_[97222]_  = ~A235 & ~A233;
  assign \new_[97225]_  = ~A266 & ~A236;
  assign \new_[97226]_  = \new_[97225]_  & \new_[97222]_ ;
  assign \new_[97229]_  = A298 & ~A267;
  assign \new_[97232]_  = ~A302 & ~A301;
  assign \new_[97233]_  = \new_[97232]_  & \new_[97229]_ ;
  assign \new_[97234]_  = \new_[97233]_  & \new_[97226]_ ;
  assign \new_[97238]_  = ~A168 & ~A169;
  assign \new_[97239]_  = ~A170 & \new_[97238]_ ;
  assign \new_[97242]_  = ~A200 & A199;
  assign \new_[97245]_  = A203 & A201;
  assign \new_[97246]_  = \new_[97245]_  & \new_[97242]_ ;
  assign \new_[97247]_  = \new_[97246]_  & \new_[97239]_ ;
  assign \new_[97250]_  = ~A235 & ~A233;
  assign \new_[97253]_  = ~A265 & ~A236;
  assign \new_[97254]_  = \new_[97253]_  & \new_[97250]_ ;
  assign \new_[97257]_  = A298 & ~A266;
  assign \new_[97260]_  = ~A302 & ~A301;
  assign \new_[97261]_  = \new_[97260]_  & \new_[97257]_ ;
  assign \new_[97262]_  = \new_[97261]_  & \new_[97254]_ ;
  assign \new_[97266]_  = ~A168 & ~A169;
  assign \new_[97267]_  = ~A170 & \new_[97266]_ ;
  assign \new_[97270]_  = ~A200 & A199;
  assign \new_[97273]_  = A203 & A201;
  assign \new_[97274]_  = \new_[97273]_  & \new_[97270]_ ;
  assign \new_[97275]_  = \new_[97274]_  & \new_[97267]_ ;
  assign \new_[97278]_  = ~A234 & ~A233;
  assign \new_[97281]_  = ~A268 & ~A266;
  assign \new_[97282]_  = \new_[97281]_  & \new_[97278]_ ;
  assign \new_[97285]_  = A298 & ~A269;
  assign \new_[97288]_  = ~A302 & ~A301;
  assign \new_[97289]_  = \new_[97288]_  & \new_[97285]_ ;
  assign \new_[97290]_  = \new_[97289]_  & \new_[97282]_ ;
  assign \new_[97294]_  = ~A168 & ~A169;
  assign \new_[97295]_  = ~A170 & \new_[97294]_ ;
  assign \new_[97298]_  = ~A200 & A199;
  assign \new_[97301]_  = A203 & A201;
  assign \new_[97302]_  = \new_[97301]_  & \new_[97298]_ ;
  assign \new_[97303]_  = \new_[97302]_  & \new_[97295]_ ;
  assign \new_[97306]_  = ~A233 & A232;
  assign \new_[97309]_  = A235 & A234;
  assign \new_[97310]_  = \new_[97309]_  & \new_[97306]_ ;
  assign \new_[97313]_  = ~A299 & A298;
  assign \new_[97316]_  = A301 & A300;
  assign \new_[97317]_  = \new_[97316]_  & \new_[97313]_ ;
  assign \new_[97318]_  = \new_[97317]_  & \new_[97310]_ ;
  assign \new_[97322]_  = ~A168 & ~A169;
  assign \new_[97323]_  = ~A170 & \new_[97322]_ ;
  assign \new_[97326]_  = ~A200 & A199;
  assign \new_[97329]_  = A203 & A201;
  assign \new_[97330]_  = \new_[97329]_  & \new_[97326]_ ;
  assign \new_[97331]_  = \new_[97330]_  & \new_[97323]_ ;
  assign \new_[97334]_  = ~A233 & A232;
  assign \new_[97337]_  = A235 & A234;
  assign \new_[97338]_  = \new_[97337]_  & \new_[97334]_ ;
  assign \new_[97341]_  = ~A299 & A298;
  assign \new_[97344]_  = A302 & A300;
  assign \new_[97345]_  = \new_[97344]_  & \new_[97341]_ ;
  assign \new_[97346]_  = \new_[97345]_  & \new_[97338]_ ;
  assign \new_[97350]_  = ~A168 & ~A169;
  assign \new_[97351]_  = ~A170 & \new_[97350]_ ;
  assign \new_[97354]_  = ~A200 & A199;
  assign \new_[97357]_  = A203 & A201;
  assign \new_[97358]_  = \new_[97357]_  & \new_[97354]_ ;
  assign \new_[97359]_  = \new_[97358]_  & \new_[97351]_ ;
  assign \new_[97362]_  = ~A233 & A232;
  assign \new_[97365]_  = A235 & A234;
  assign \new_[97366]_  = \new_[97365]_  & \new_[97362]_ ;
  assign \new_[97369]_  = ~A266 & A265;
  assign \new_[97372]_  = A268 & A267;
  assign \new_[97373]_  = \new_[97372]_  & \new_[97369]_ ;
  assign \new_[97374]_  = \new_[97373]_  & \new_[97366]_ ;
  assign \new_[97378]_  = ~A168 & ~A169;
  assign \new_[97379]_  = ~A170 & \new_[97378]_ ;
  assign \new_[97382]_  = ~A200 & A199;
  assign \new_[97385]_  = A203 & A201;
  assign \new_[97386]_  = \new_[97385]_  & \new_[97382]_ ;
  assign \new_[97387]_  = \new_[97386]_  & \new_[97379]_ ;
  assign \new_[97390]_  = ~A233 & A232;
  assign \new_[97393]_  = A235 & A234;
  assign \new_[97394]_  = \new_[97393]_  & \new_[97390]_ ;
  assign \new_[97397]_  = ~A266 & A265;
  assign \new_[97400]_  = A269 & A267;
  assign \new_[97401]_  = \new_[97400]_  & \new_[97397]_ ;
  assign \new_[97402]_  = \new_[97401]_  & \new_[97394]_ ;
  assign \new_[97406]_  = ~A168 & ~A169;
  assign \new_[97407]_  = ~A170 & \new_[97406]_ ;
  assign \new_[97410]_  = ~A200 & A199;
  assign \new_[97413]_  = A203 & A201;
  assign \new_[97414]_  = \new_[97413]_  & \new_[97410]_ ;
  assign \new_[97415]_  = \new_[97414]_  & \new_[97407]_ ;
  assign \new_[97418]_  = ~A233 & A232;
  assign \new_[97421]_  = A236 & A234;
  assign \new_[97422]_  = \new_[97421]_  & \new_[97418]_ ;
  assign \new_[97425]_  = ~A299 & A298;
  assign \new_[97428]_  = A301 & A300;
  assign \new_[97429]_  = \new_[97428]_  & \new_[97425]_ ;
  assign \new_[97430]_  = \new_[97429]_  & \new_[97422]_ ;
  assign \new_[97434]_  = ~A168 & ~A169;
  assign \new_[97435]_  = ~A170 & \new_[97434]_ ;
  assign \new_[97438]_  = ~A200 & A199;
  assign \new_[97441]_  = A203 & A201;
  assign \new_[97442]_  = \new_[97441]_  & \new_[97438]_ ;
  assign \new_[97443]_  = \new_[97442]_  & \new_[97435]_ ;
  assign \new_[97446]_  = ~A233 & A232;
  assign \new_[97449]_  = A236 & A234;
  assign \new_[97450]_  = \new_[97449]_  & \new_[97446]_ ;
  assign \new_[97453]_  = ~A299 & A298;
  assign \new_[97456]_  = A302 & A300;
  assign \new_[97457]_  = \new_[97456]_  & \new_[97453]_ ;
  assign \new_[97458]_  = \new_[97457]_  & \new_[97450]_ ;
  assign \new_[97462]_  = ~A168 & ~A169;
  assign \new_[97463]_  = ~A170 & \new_[97462]_ ;
  assign \new_[97466]_  = ~A200 & A199;
  assign \new_[97469]_  = A203 & A201;
  assign \new_[97470]_  = \new_[97469]_  & \new_[97466]_ ;
  assign \new_[97471]_  = \new_[97470]_  & \new_[97463]_ ;
  assign \new_[97474]_  = ~A233 & A232;
  assign \new_[97477]_  = A236 & A234;
  assign \new_[97478]_  = \new_[97477]_  & \new_[97474]_ ;
  assign \new_[97481]_  = ~A266 & A265;
  assign \new_[97484]_  = A268 & A267;
  assign \new_[97485]_  = \new_[97484]_  & \new_[97481]_ ;
  assign \new_[97486]_  = \new_[97485]_  & \new_[97478]_ ;
  assign \new_[97490]_  = ~A168 & ~A169;
  assign \new_[97491]_  = ~A170 & \new_[97490]_ ;
  assign \new_[97494]_  = ~A200 & A199;
  assign \new_[97497]_  = A203 & A201;
  assign \new_[97498]_  = \new_[97497]_  & \new_[97494]_ ;
  assign \new_[97499]_  = \new_[97498]_  & \new_[97491]_ ;
  assign \new_[97502]_  = ~A233 & A232;
  assign \new_[97505]_  = A236 & A234;
  assign \new_[97506]_  = \new_[97505]_  & \new_[97502]_ ;
  assign \new_[97509]_  = ~A266 & A265;
  assign \new_[97512]_  = A269 & A267;
  assign \new_[97513]_  = \new_[97512]_  & \new_[97509]_ ;
  assign \new_[97514]_  = \new_[97513]_  & \new_[97506]_ ;
  assign \new_[97518]_  = ~A168 & ~A169;
  assign \new_[97519]_  = ~A170 & \new_[97518]_ ;
  assign \new_[97522]_  = ~A200 & A199;
  assign \new_[97525]_  = A203 & A201;
  assign \new_[97526]_  = \new_[97525]_  & \new_[97522]_ ;
  assign \new_[97527]_  = \new_[97526]_  & \new_[97519]_ ;
  assign \new_[97530]_  = ~A233 & ~A232;
  assign \new_[97533]_  = ~A268 & ~A266;
  assign \new_[97534]_  = \new_[97533]_  & \new_[97530]_ ;
  assign \new_[97537]_  = A298 & ~A269;
  assign \new_[97540]_  = ~A302 & ~A301;
  assign \new_[97541]_  = \new_[97540]_  & \new_[97537]_ ;
  assign \new_[97542]_  = \new_[97541]_  & \new_[97534]_ ;
  assign \new_[97545]_  = ~A167 & A170;
  assign \new_[97548]_  = A199 & ~A166;
  assign \new_[97549]_  = \new_[97548]_  & \new_[97545]_ ;
  assign \new_[97552]_  = A201 & ~A200;
  assign \new_[97555]_  = ~A233 & A202;
  assign \new_[97556]_  = \new_[97555]_  & \new_[97552]_ ;
  assign \new_[97557]_  = \new_[97556]_  & \new_[97549]_ ;
  assign \new_[97560]_  = ~A236 & ~A235;
  assign \new_[97563]_  = ~A268 & ~A266;
  assign \new_[97564]_  = \new_[97563]_  & \new_[97560]_ ;
  assign \new_[97567]_  = A298 & ~A269;
  assign \new_[97570]_  = ~A302 & ~A301;
  assign \new_[97571]_  = \new_[97570]_  & \new_[97567]_ ;
  assign \new_[97572]_  = \new_[97571]_  & \new_[97564]_ ;
  assign \new_[97575]_  = ~A167 & A170;
  assign \new_[97578]_  = A199 & ~A166;
  assign \new_[97579]_  = \new_[97578]_  & \new_[97575]_ ;
  assign \new_[97582]_  = A201 & ~A200;
  assign \new_[97585]_  = ~A233 & A203;
  assign \new_[97586]_  = \new_[97585]_  & \new_[97582]_ ;
  assign \new_[97587]_  = \new_[97586]_  & \new_[97579]_ ;
  assign \new_[97590]_  = ~A236 & ~A235;
  assign \new_[97593]_  = ~A268 & ~A266;
  assign \new_[97594]_  = \new_[97593]_  & \new_[97590]_ ;
  assign \new_[97597]_  = A298 & ~A269;
  assign \new_[97600]_  = ~A302 & ~A301;
  assign \new_[97601]_  = \new_[97600]_  & \new_[97597]_ ;
  assign \new_[97602]_  = \new_[97601]_  & \new_[97594]_ ;
  assign \new_[97605]_  = ~A168 & A169;
  assign \new_[97608]_  = ~A166 & A167;
  assign \new_[97609]_  = \new_[97608]_  & \new_[97605]_ ;
  assign \new_[97612]_  = ~A200 & A199;
  assign \new_[97615]_  = A202 & A201;
  assign \new_[97616]_  = \new_[97615]_  & \new_[97612]_ ;
  assign \new_[97617]_  = \new_[97616]_  & \new_[97609]_ ;
  assign \new_[97620]_  = A233 & A232;
  assign \new_[97623]_  = ~A268 & A265;
  assign \new_[97624]_  = \new_[97623]_  & \new_[97620]_ ;
  assign \new_[97627]_  = ~A299 & ~A269;
  assign \new_[97630]_  = ~A302 & ~A301;
  assign \new_[97631]_  = \new_[97630]_  & \new_[97627]_ ;
  assign \new_[97632]_  = \new_[97631]_  & \new_[97624]_ ;
  assign \new_[97635]_  = ~A168 & A169;
  assign \new_[97638]_  = ~A166 & A167;
  assign \new_[97639]_  = \new_[97638]_  & \new_[97635]_ ;
  assign \new_[97642]_  = ~A200 & A199;
  assign \new_[97645]_  = A202 & A201;
  assign \new_[97646]_  = \new_[97645]_  & \new_[97642]_ ;
  assign \new_[97647]_  = \new_[97646]_  & \new_[97639]_ ;
  assign \new_[97650]_  = ~A235 & ~A233;
  assign \new_[97653]_  = A265 & ~A236;
  assign \new_[97654]_  = \new_[97653]_  & \new_[97650]_ ;
  assign \new_[97657]_  = A298 & A266;
  assign \new_[97660]_  = ~A302 & ~A301;
  assign \new_[97661]_  = \new_[97660]_  & \new_[97657]_ ;
  assign \new_[97662]_  = \new_[97661]_  & \new_[97654]_ ;
  assign \new_[97665]_  = ~A168 & A169;
  assign \new_[97668]_  = ~A166 & A167;
  assign \new_[97669]_  = \new_[97668]_  & \new_[97665]_ ;
  assign \new_[97672]_  = ~A200 & A199;
  assign \new_[97675]_  = A202 & A201;
  assign \new_[97676]_  = \new_[97675]_  & \new_[97672]_ ;
  assign \new_[97677]_  = \new_[97676]_  & \new_[97669]_ ;
  assign \new_[97680]_  = ~A235 & ~A233;
  assign \new_[97683]_  = ~A266 & ~A236;
  assign \new_[97684]_  = \new_[97683]_  & \new_[97680]_ ;
  assign \new_[97687]_  = ~A269 & ~A268;
  assign \new_[97690]_  = ~A300 & A298;
  assign \new_[97691]_  = \new_[97690]_  & \new_[97687]_ ;
  assign \new_[97692]_  = \new_[97691]_  & \new_[97684]_ ;
  assign \new_[97695]_  = ~A168 & A169;
  assign \new_[97698]_  = ~A166 & A167;
  assign \new_[97699]_  = \new_[97698]_  & \new_[97695]_ ;
  assign \new_[97702]_  = ~A200 & A199;
  assign \new_[97705]_  = A202 & A201;
  assign \new_[97706]_  = \new_[97705]_  & \new_[97702]_ ;
  assign \new_[97707]_  = \new_[97706]_  & \new_[97699]_ ;
  assign \new_[97710]_  = ~A235 & ~A233;
  assign \new_[97713]_  = ~A266 & ~A236;
  assign \new_[97714]_  = \new_[97713]_  & \new_[97710]_ ;
  assign \new_[97717]_  = ~A269 & ~A268;
  assign \new_[97720]_  = A299 & A298;
  assign \new_[97721]_  = \new_[97720]_  & \new_[97717]_ ;
  assign \new_[97722]_  = \new_[97721]_  & \new_[97714]_ ;
  assign \new_[97725]_  = ~A168 & A169;
  assign \new_[97728]_  = ~A166 & A167;
  assign \new_[97729]_  = \new_[97728]_  & \new_[97725]_ ;
  assign \new_[97732]_  = ~A200 & A199;
  assign \new_[97735]_  = A202 & A201;
  assign \new_[97736]_  = \new_[97735]_  & \new_[97732]_ ;
  assign \new_[97737]_  = \new_[97736]_  & \new_[97729]_ ;
  assign \new_[97740]_  = ~A235 & ~A233;
  assign \new_[97743]_  = ~A266 & ~A236;
  assign \new_[97744]_  = \new_[97743]_  & \new_[97740]_ ;
  assign \new_[97747]_  = ~A269 & ~A268;
  assign \new_[97750]_  = ~A299 & ~A298;
  assign \new_[97751]_  = \new_[97750]_  & \new_[97747]_ ;
  assign \new_[97752]_  = \new_[97751]_  & \new_[97744]_ ;
  assign \new_[97755]_  = ~A168 & A169;
  assign \new_[97758]_  = ~A166 & A167;
  assign \new_[97759]_  = \new_[97758]_  & \new_[97755]_ ;
  assign \new_[97762]_  = ~A200 & A199;
  assign \new_[97765]_  = A202 & A201;
  assign \new_[97766]_  = \new_[97765]_  & \new_[97762]_ ;
  assign \new_[97767]_  = \new_[97766]_  & \new_[97759]_ ;
  assign \new_[97770]_  = ~A235 & ~A233;
  assign \new_[97773]_  = ~A266 & ~A236;
  assign \new_[97774]_  = \new_[97773]_  & \new_[97770]_ ;
  assign \new_[97777]_  = A298 & ~A267;
  assign \new_[97780]_  = ~A302 & ~A301;
  assign \new_[97781]_  = \new_[97780]_  & \new_[97777]_ ;
  assign \new_[97782]_  = \new_[97781]_  & \new_[97774]_ ;
  assign \new_[97785]_  = ~A168 & A169;
  assign \new_[97788]_  = ~A166 & A167;
  assign \new_[97789]_  = \new_[97788]_  & \new_[97785]_ ;
  assign \new_[97792]_  = ~A200 & A199;
  assign \new_[97795]_  = A202 & A201;
  assign \new_[97796]_  = \new_[97795]_  & \new_[97792]_ ;
  assign \new_[97797]_  = \new_[97796]_  & \new_[97789]_ ;
  assign \new_[97800]_  = ~A235 & ~A233;
  assign \new_[97803]_  = ~A265 & ~A236;
  assign \new_[97804]_  = \new_[97803]_  & \new_[97800]_ ;
  assign \new_[97807]_  = A298 & ~A266;
  assign \new_[97810]_  = ~A302 & ~A301;
  assign \new_[97811]_  = \new_[97810]_  & \new_[97807]_ ;
  assign \new_[97812]_  = \new_[97811]_  & \new_[97804]_ ;
  assign \new_[97815]_  = ~A168 & A169;
  assign \new_[97818]_  = ~A166 & A167;
  assign \new_[97819]_  = \new_[97818]_  & \new_[97815]_ ;
  assign \new_[97822]_  = ~A200 & A199;
  assign \new_[97825]_  = A202 & A201;
  assign \new_[97826]_  = \new_[97825]_  & \new_[97822]_ ;
  assign \new_[97827]_  = \new_[97826]_  & \new_[97819]_ ;
  assign \new_[97830]_  = ~A234 & ~A233;
  assign \new_[97833]_  = ~A268 & ~A266;
  assign \new_[97834]_  = \new_[97833]_  & \new_[97830]_ ;
  assign \new_[97837]_  = A298 & ~A269;
  assign \new_[97840]_  = ~A302 & ~A301;
  assign \new_[97841]_  = \new_[97840]_  & \new_[97837]_ ;
  assign \new_[97842]_  = \new_[97841]_  & \new_[97834]_ ;
  assign \new_[97845]_  = ~A168 & A169;
  assign \new_[97848]_  = ~A166 & A167;
  assign \new_[97849]_  = \new_[97848]_  & \new_[97845]_ ;
  assign \new_[97852]_  = ~A200 & A199;
  assign \new_[97855]_  = A202 & A201;
  assign \new_[97856]_  = \new_[97855]_  & \new_[97852]_ ;
  assign \new_[97857]_  = \new_[97856]_  & \new_[97849]_ ;
  assign \new_[97860]_  = ~A233 & A232;
  assign \new_[97863]_  = A235 & A234;
  assign \new_[97864]_  = \new_[97863]_  & \new_[97860]_ ;
  assign \new_[97867]_  = ~A299 & A298;
  assign \new_[97870]_  = A301 & A300;
  assign \new_[97871]_  = \new_[97870]_  & \new_[97867]_ ;
  assign \new_[97872]_  = \new_[97871]_  & \new_[97864]_ ;
  assign \new_[97875]_  = ~A168 & A169;
  assign \new_[97878]_  = ~A166 & A167;
  assign \new_[97879]_  = \new_[97878]_  & \new_[97875]_ ;
  assign \new_[97882]_  = ~A200 & A199;
  assign \new_[97885]_  = A202 & A201;
  assign \new_[97886]_  = \new_[97885]_  & \new_[97882]_ ;
  assign \new_[97887]_  = \new_[97886]_  & \new_[97879]_ ;
  assign \new_[97890]_  = ~A233 & A232;
  assign \new_[97893]_  = A235 & A234;
  assign \new_[97894]_  = \new_[97893]_  & \new_[97890]_ ;
  assign \new_[97897]_  = ~A299 & A298;
  assign \new_[97900]_  = A302 & A300;
  assign \new_[97901]_  = \new_[97900]_  & \new_[97897]_ ;
  assign \new_[97902]_  = \new_[97901]_  & \new_[97894]_ ;
  assign \new_[97905]_  = ~A168 & A169;
  assign \new_[97908]_  = ~A166 & A167;
  assign \new_[97909]_  = \new_[97908]_  & \new_[97905]_ ;
  assign \new_[97912]_  = ~A200 & A199;
  assign \new_[97915]_  = A202 & A201;
  assign \new_[97916]_  = \new_[97915]_  & \new_[97912]_ ;
  assign \new_[97917]_  = \new_[97916]_  & \new_[97909]_ ;
  assign \new_[97920]_  = ~A233 & A232;
  assign \new_[97923]_  = A235 & A234;
  assign \new_[97924]_  = \new_[97923]_  & \new_[97920]_ ;
  assign \new_[97927]_  = ~A266 & A265;
  assign \new_[97930]_  = A268 & A267;
  assign \new_[97931]_  = \new_[97930]_  & \new_[97927]_ ;
  assign \new_[97932]_  = \new_[97931]_  & \new_[97924]_ ;
  assign \new_[97935]_  = ~A168 & A169;
  assign \new_[97938]_  = ~A166 & A167;
  assign \new_[97939]_  = \new_[97938]_  & \new_[97935]_ ;
  assign \new_[97942]_  = ~A200 & A199;
  assign \new_[97945]_  = A202 & A201;
  assign \new_[97946]_  = \new_[97945]_  & \new_[97942]_ ;
  assign \new_[97947]_  = \new_[97946]_  & \new_[97939]_ ;
  assign \new_[97950]_  = ~A233 & A232;
  assign \new_[97953]_  = A235 & A234;
  assign \new_[97954]_  = \new_[97953]_  & \new_[97950]_ ;
  assign \new_[97957]_  = ~A266 & A265;
  assign \new_[97960]_  = A269 & A267;
  assign \new_[97961]_  = \new_[97960]_  & \new_[97957]_ ;
  assign \new_[97962]_  = \new_[97961]_  & \new_[97954]_ ;
  assign \new_[97965]_  = ~A168 & A169;
  assign \new_[97968]_  = ~A166 & A167;
  assign \new_[97969]_  = \new_[97968]_  & \new_[97965]_ ;
  assign \new_[97972]_  = ~A200 & A199;
  assign \new_[97975]_  = A202 & A201;
  assign \new_[97976]_  = \new_[97975]_  & \new_[97972]_ ;
  assign \new_[97977]_  = \new_[97976]_  & \new_[97969]_ ;
  assign \new_[97980]_  = ~A233 & A232;
  assign \new_[97983]_  = A236 & A234;
  assign \new_[97984]_  = \new_[97983]_  & \new_[97980]_ ;
  assign \new_[97987]_  = ~A299 & A298;
  assign \new_[97990]_  = A301 & A300;
  assign \new_[97991]_  = \new_[97990]_  & \new_[97987]_ ;
  assign \new_[97992]_  = \new_[97991]_  & \new_[97984]_ ;
  assign \new_[97995]_  = ~A168 & A169;
  assign \new_[97998]_  = ~A166 & A167;
  assign \new_[97999]_  = \new_[97998]_  & \new_[97995]_ ;
  assign \new_[98002]_  = ~A200 & A199;
  assign \new_[98005]_  = A202 & A201;
  assign \new_[98006]_  = \new_[98005]_  & \new_[98002]_ ;
  assign \new_[98007]_  = \new_[98006]_  & \new_[97999]_ ;
  assign \new_[98010]_  = ~A233 & A232;
  assign \new_[98013]_  = A236 & A234;
  assign \new_[98014]_  = \new_[98013]_  & \new_[98010]_ ;
  assign \new_[98017]_  = ~A299 & A298;
  assign \new_[98020]_  = A302 & A300;
  assign \new_[98021]_  = \new_[98020]_  & \new_[98017]_ ;
  assign \new_[98022]_  = \new_[98021]_  & \new_[98014]_ ;
  assign \new_[98025]_  = ~A168 & A169;
  assign \new_[98028]_  = ~A166 & A167;
  assign \new_[98029]_  = \new_[98028]_  & \new_[98025]_ ;
  assign \new_[98032]_  = ~A200 & A199;
  assign \new_[98035]_  = A202 & A201;
  assign \new_[98036]_  = \new_[98035]_  & \new_[98032]_ ;
  assign \new_[98037]_  = \new_[98036]_  & \new_[98029]_ ;
  assign \new_[98040]_  = ~A233 & A232;
  assign \new_[98043]_  = A236 & A234;
  assign \new_[98044]_  = \new_[98043]_  & \new_[98040]_ ;
  assign \new_[98047]_  = ~A266 & A265;
  assign \new_[98050]_  = A268 & A267;
  assign \new_[98051]_  = \new_[98050]_  & \new_[98047]_ ;
  assign \new_[98052]_  = \new_[98051]_  & \new_[98044]_ ;
  assign \new_[98055]_  = ~A168 & A169;
  assign \new_[98058]_  = ~A166 & A167;
  assign \new_[98059]_  = \new_[98058]_  & \new_[98055]_ ;
  assign \new_[98062]_  = ~A200 & A199;
  assign \new_[98065]_  = A202 & A201;
  assign \new_[98066]_  = \new_[98065]_  & \new_[98062]_ ;
  assign \new_[98067]_  = \new_[98066]_  & \new_[98059]_ ;
  assign \new_[98070]_  = ~A233 & A232;
  assign \new_[98073]_  = A236 & A234;
  assign \new_[98074]_  = \new_[98073]_  & \new_[98070]_ ;
  assign \new_[98077]_  = ~A266 & A265;
  assign \new_[98080]_  = A269 & A267;
  assign \new_[98081]_  = \new_[98080]_  & \new_[98077]_ ;
  assign \new_[98082]_  = \new_[98081]_  & \new_[98074]_ ;
  assign \new_[98085]_  = ~A168 & A169;
  assign \new_[98088]_  = ~A166 & A167;
  assign \new_[98089]_  = \new_[98088]_  & \new_[98085]_ ;
  assign \new_[98092]_  = ~A200 & A199;
  assign \new_[98095]_  = A202 & A201;
  assign \new_[98096]_  = \new_[98095]_  & \new_[98092]_ ;
  assign \new_[98097]_  = \new_[98096]_  & \new_[98089]_ ;
  assign \new_[98100]_  = ~A233 & ~A232;
  assign \new_[98103]_  = ~A268 & ~A266;
  assign \new_[98104]_  = \new_[98103]_  & \new_[98100]_ ;
  assign \new_[98107]_  = A298 & ~A269;
  assign \new_[98110]_  = ~A302 & ~A301;
  assign \new_[98111]_  = \new_[98110]_  & \new_[98107]_ ;
  assign \new_[98112]_  = \new_[98111]_  & \new_[98104]_ ;
  assign \new_[98115]_  = ~A168 & A169;
  assign \new_[98118]_  = ~A166 & A167;
  assign \new_[98119]_  = \new_[98118]_  & \new_[98115]_ ;
  assign \new_[98122]_  = ~A200 & A199;
  assign \new_[98125]_  = A203 & A201;
  assign \new_[98126]_  = \new_[98125]_  & \new_[98122]_ ;
  assign \new_[98127]_  = \new_[98126]_  & \new_[98119]_ ;
  assign \new_[98130]_  = A233 & A232;
  assign \new_[98133]_  = ~A268 & A265;
  assign \new_[98134]_  = \new_[98133]_  & \new_[98130]_ ;
  assign \new_[98137]_  = ~A299 & ~A269;
  assign \new_[98140]_  = ~A302 & ~A301;
  assign \new_[98141]_  = \new_[98140]_  & \new_[98137]_ ;
  assign \new_[98142]_  = \new_[98141]_  & \new_[98134]_ ;
  assign \new_[98145]_  = ~A168 & A169;
  assign \new_[98148]_  = ~A166 & A167;
  assign \new_[98149]_  = \new_[98148]_  & \new_[98145]_ ;
  assign \new_[98152]_  = ~A200 & A199;
  assign \new_[98155]_  = A203 & A201;
  assign \new_[98156]_  = \new_[98155]_  & \new_[98152]_ ;
  assign \new_[98157]_  = \new_[98156]_  & \new_[98149]_ ;
  assign \new_[98160]_  = ~A235 & ~A233;
  assign \new_[98163]_  = A265 & ~A236;
  assign \new_[98164]_  = \new_[98163]_  & \new_[98160]_ ;
  assign \new_[98167]_  = A298 & A266;
  assign \new_[98170]_  = ~A302 & ~A301;
  assign \new_[98171]_  = \new_[98170]_  & \new_[98167]_ ;
  assign \new_[98172]_  = \new_[98171]_  & \new_[98164]_ ;
  assign \new_[98175]_  = ~A168 & A169;
  assign \new_[98178]_  = ~A166 & A167;
  assign \new_[98179]_  = \new_[98178]_  & \new_[98175]_ ;
  assign \new_[98182]_  = ~A200 & A199;
  assign \new_[98185]_  = A203 & A201;
  assign \new_[98186]_  = \new_[98185]_  & \new_[98182]_ ;
  assign \new_[98187]_  = \new_[98186]_  & \new_[98179]_ ;
  assign \new_[98190]_  = ~A235 & ~A233;
  assign \new_[98193]_  = ~A266 & ~A236;
  assign \new_[98194]_  = \new_[98193]_  & \new_[98190]_ ;
  assign \new_[98197]_  = ~A269 & ~A268;
  assign \new_[98200]_  = ~A300 & A298;
  assign \new_[98201]_  = \new_[98200]_  & \new_[98197]_ ;
  assign \new_[98202]_  = \new_[98201]_  & \new_[98194]_ ;
  assign \new_[98205]_  = ~A168 & A169;
  assign \new_[98208]_  = ~A166 & A167;
  assign \new_[98209]_  = \new_[98208]_  & \new_[98205]_ ;
  assign \new_[98212]_  = ~A200 & A199;
  assign \new_[98215]_  = A203 & A201;
  assign \new_[98216]_  = \new_[98215]_  & \new_[98212]_ ;
  assign \new_[98217]_  = \new_[98216]_  & \new_[98209]_ ;
  assign \new_[98220]_  = ~A235 & ~A233;
  assign \new_[98223]_  = ~A266 & ~A236;
  assign \new_[98224]_  = \new_[98223]_  & \new_[98220]_ ;
  assign \new_[98227]_  = ~A269 & ~A268;
  assign \new_[98230]_  = A299 & A298;
  assign \new_[98231]_  = \new_[98230]_  & \new_[98227]_ ;
  assign \new_[98232]_  = \new_[98231]_  & \new_[98224]_ ;
  assign \new_[98235]_  = ~A168 & A169;
  assign \new_[98238]_  = ~A166 & A167;
  assign \new_[98239]_  = \new_[98238]_  & \new_[98235]_ ;
  assign \new_[98242]_  = ~A200 & A199;
  assign \new_[98245]_  = A203 & A201;
  assign \new_[98246]_  = \new_[98245]_  & \new_[98242]_ ;
  assign \new_[98247]_  = \new_[98246]_  & \new_[98239]_ ;
  assign \new_[98250]_  = ~A235 & ~A233;
  assign \new_[98253]_  = ~A266 & ~A236;
  assign \new_[98254]_  = \new_[98253]_  & \new_[98250]_ ;
  assign \new_[98257]_  = ~A269 & ~A268;
  assign \new_[98260]_  = ~A299 & ~A298;
  assign \new_[98261]_  = \new_[98260]_  & \new_[98257]_ ;
  assign \new_[98262]_  = \new_[98261]_  & \new_[98254]_ ;
  assign \new_[98265]_  = ~A168 & A169;
  assign \new_[98268]_  = ~A166 & A167;
  assign \new_[98269]_  = \new_[98268]_  & \new_[98265]_ ;
  assign \new_[98272]_  = ~A200 & A199;
  assign \new_[98275]_  = A203 & A201;
  assign \new_[98276]_  = \new_[98275]_  & \new_[98272]_ ;
  assign \new_[98277]_  = \new_[98276]_  & \new_[98269]_ ;
  assign \new_[98280]_  = ~A235 & ~A233;
  assign \new_[98283]_  = ~A266 & ~A236;
  assign \new_[98284]_  = \new_[98283]_  & \new_[98280]_ ;
  assign \new_[98287]_  = A298 & ~A267;
  assign \new_[98290]_  = ~A302 & ~A301;
  assign \new_[98291]_  = \new_[98290]_  & \new_[98287]_ ;
  assign \new_[98292]_  = \new_[98291]_  & \new_[98284]_ ;
  assign \new_[98295]_  = ~A168 & A169;
  assign \new_[98298]_  = ~A166 & A167;
  assign \new_[98299]_  = \new_[98298]_  & \new_[98295]_ ;
  assign \new_[98302]_  = ~A200 & A199;
  assign \new_[98305]_  = A203 & A201;
  assign \new_[98306]_  = \new_[98305]_  & \new_[98302]_ ;
  assign \new_[98307]_  = \new_[98306]_  & \new_[98299]_ ;
  assign \new_[98310]_  = ~A235 & ~A233;
  assign \new_[98313]_  = ~A265 & ~A236;
  assign \new_[98314]_  = \new_[98313]_  & \new_[98310]_ ;
  assign \new_[98317]_  = A298 & ~A266;
  assign \new_[98320]_  = ~A302 & ~A301;
  assign \new_[98321]_  = \new_[98320]_  & \new_[98317]_ ;
  assign \new_[98322]_  = \new_[98321]_  & \new_[98314]_ ;
  assign \new_[98325]_  = ~A168 & A169;
  assign \new_[98328]_  = ~A166 & A167;
  assign \new_[98329]_  = \new_[98328]_  & \new_[98325]_ ;
  assign \new_[98332]_  = ~A200 & A199;
  assign \new_[98335]_  = A203 & A201;
  assign \new_[98336]_  = \new_[98335]_  & \new_[98332]_ ;
  assign \new_[98337]_  = \new_[98336]_  & \new_[98329]_ ;
  assign \new_[98340]_  = ~A234 & ~A233;
  assign \new_[98343]_  = ~A268 & ~A266;
  assign \new_[98344]_  = \new_[98343]_  & \new_[98340]_ ;
  assign \new_[98347]_  = A298 & ~A269;
  assign \new_[98350]_  = ~A302 & ~A301;
  assign \new_[98351]_  = \new_[98350]_  & \new_[98347]_ ;
  assign \new_[98352]_  = \new_[98351]_  & \new_[98344]_ ;
  assign \new_[98355]_  = ~A168 & A169;
  assign \new_[98358]_  = ~A166 & A167;
  assign \new_[98359]_  = \new_[98358]_  & \new_[98355]_ ;
  assign \new_[98362]_  = ~A200 & A199;
  assign \new_[98365]_  = A203 & A201;
  assign \new_[98366]_  = \new_[98365]_  & \new_[98362]_ ;
  assign \new_[98367]_  = \new_[98366]_  & \new_[98359]_ ;
  assign \new_[98370]_  = ~A233 & A232;
  assign \new_[98373]_  = A235 & A234;
  assign \new_[98374]_  = \new_[98373]_  & \new_[98370]_ ;
  assign \new_[98377]_  = ~A299 & A298;
  assign \new_[98380]_  = A301 & A300;
  assign \new_[98381]_  = \new_[98380]_  & \new_[98377]_ ;
  assign \new_[98382]_  = \new_[98381]_  & \new_[98374]_ ;
  assign \new_[98385]_  = ~A168 & A169;
  assign \new_[98388]_  = ~A166 & A167;
  assign \new_[98389]_  = \new_[98388]_  & \new_[98385]_ ;
  assign \new_[98392]_  = ~A200 & A199;
  assign \new_[98395]_  = A203 & A201;
  assign \new_[98396]_  = \new_[98395]_  & \new_[98392]_ ;
  assign \new_[98397]_  = \new_[98396]_  & \new_[98389]_ ;
  assign \new_[98400]_  = ~A233 & A232;
  assign \new_[98403]_  = A235 & A234;
  assign \new_[98404]_  = \new_[98403]_  & \new_[98400]_ ;
  assign \new_[98407]_  = ~A299 & A298;
  assign \new_[98410]_  = A302 & A300;
  assign \new_[98411]_  = \new_[98410]_  & \new_[98407]_ ;
  assign \new_[98412]_  = \new_[98411]_  & \new_[98404]_ ;
  assign \new_[98415]_  = ~A168 & A169;
  assign \new_[98418]_  = ~A166 & A167;
  assign \new_[98419]_  = \new_[98418]_  & \new_[98415]_ ;
  assign \new_[98422]_  = ~A200 & A199;
  assign \new_[98425]_  = A203 & A201;
  assign \new_[98426]_  = \new_[98425]_  & \new_[98422]_ ;
  assign \new_[98427]_  = \new_[98426]_  & \new_[98419]_ ;
  assign \new_[98430]_  = ~A233 & A232;
  assign \new_[98433]_  = A235 & A234;
  assign \new_[98434]_  = \new_[98433]_  & \new_[98430]_ ;
  assign \new_[98437]_  = ~A266 & A265;
  assign \new_[98440]_  = A268 & A267;
  assign \new_[98441]_  = \new_[98440]_  & \new_[98437]_ ;
  assign \new_[98442]_  = \new_[98441]_  & \new_[98434]_ ;
  assign \new_[98445]_  = ~A168 & A169;
  assign \new_[98448]_  = ~A166 & A167;
  assign \new_[98449]_  = \new_[98448]_  & \new_[98445]_ ;
  assign \new_[98452]_  = ~A200 & A199;
  assign \new_[98455]_  = A203 & A201;
  assign \new_[98456]_  = \new_[98455]_  & \new_[98452]_ ;
  assign \new_[98457]_  = \new_[98456]_  & \new_[98449]_ ;
  assign \new_[98460]_  = ~A233 & A232;
  assign \new_[98463]_  = A235 & A234;
  assign \new_[98464]_  = \new_[98463]_  & \new_[98460]_ ;
  assign \new_[98467]_  = ~A266 & A265;
  assign \new_[98470]_  = A269 & A267;
  assign \new_[98471]_  = \new_[98470]_  & \new_[98467]_ ;
  assign \new_[98472]_  = \new_[98471]_  & \new_[98464]_ ;
  assign \new_[98475]_  = ~A168 & A169;
  assign \new_[98478]_  = ~A166 & A167;
  assign \new_[98479]_  = \new_[98478]_  & \new_[98475]_ ;
  assign \new_[98482]_  = ~A200 & A199;
  assign \new_[98485]_  = A203 & A201;
  assign \new_[98486]_  = \new_[98485]_  & \new_[98482]_ ;
  assign \new_[98487]_  = \new_[98486]_  & \new_[98479]_ ;
  assign \new_[98490]_  = ~A233 & A232;
  assign \new_[98493]_  = A236 & A234;
  assign \new_[98494]_  = \new_[98493]_  & \new_[98490]_ ;
  assign \new_[98497]_  = ~A299 & A298;
  assign \new_[98500]_  = A301 & A300;
  assign \new_[98501]_  = \new_[98500]_  & \new_[98497]_ ;
  assign \new_[98502]_  = \new_[98501]_  & \new_[98494]_ ;
  assign \new_[98505]_  = ~A168 & A169;
  assign \new_[98508]_  = ~A166 & A167;
  assign \new_[98509]_  = \new_[98508]_  & \new_[98505]_ ;
  assign \new_[98512]_  = ~A200 & A199;
  assign \new_[98515]_  = A203 & A201;
  assign \new_[98516]_  = \new_[98515]_  & \new_[98512]_ ;
  assign \new_[98517]_  = \new_[98516]_  & \new_[98509]_ ;
  assign \new_[98520]_  = ~A233 & A232;
  assign \new_[98523]_  = A236 & A234;
  assign \new_[98524]_  = \new_[98523]_  & \new_[98520]_ ;
  assign \new_[98527]_  = ~A299 & A298;
  assign \new_[98530]_  = A302 & A300;
  assign \new_[98531]_  = \new_[98530]_  & \new_[98527]_ ;
  assign \new_[98532]_  = \new_[98531]_  & \new_[98524]_ ;
  assign \new_[98535]_  = ~A168 & A169;
  assign \new_[98538]_  = ~A166 & A167;
  assign \new_[98539]_  = \new_[98538]_  & \new_[98535]_ ;
  assign \new_[98542]_  = ~A200 & A199;
  assign \new_[98545]_  = A203 & A201;
  assign \new_[98546]_  = \new_[98545]_  & \new_[98542]_ ;
  assign \new_[98547]_  = \new_[98546]_  & \new_[98539]_ ;
  assign \new_[98550]_  = ~A233 & A232;
  assign \new_[98553]_  = A236 & A234;
  assign \new_[98554]_  = \new_[98553]_  & \new_[98550]_ ;
  assign \new_[98557]_  = ~A266 & A265;
  assign \new_[98560]_  = A268 & A267;
  assign \new_[98561]_  = \new_[98560]_  & \new_[98557]_ ;
  assign \new_[98562]_  = \new_[98561]_  & \new_[98554]_ ;
  assign \new_[98565]_  = ~A168 & A169;
  assign \new_[98568]_  = ~A166 & A167;
  assign \new_[98569]_  = \new_[98568]_  & \new_[98565]_ ;
  assign \new_[98572]_  = ~A200 & A199;
  assign \new_[98575]_  = A203 & A201;
  assign \new_[98576]_  = \new_[98575]_  & \new_[98572]_ ;
  assign \new_[98577]_  = \new_[98576]_  & \new_[98569]_ ;
  assign \new_[98580]_  = ~A233 & A232;
  assign \new_[98583]_  = A236 & A234;
  assign \new_[98584]_  = \new_[98583]_  & \new_[98580]_ ;
  assign \new_[98587]_  = ~A266 & A265;
  assign \new_[98590]_  = A269 & A267;
  assign \new_[98591]_  = \new_[98590]_  & \new_[98587]_ ;
  assign \new_[98592]_  = \new_[98591]_  & \new_[98584]_ ;
  assign \new_[98595]_  = ~A168 & A169;
  assign \new_[98598]_  = ~A166 & A167;
  assign \new_[98599]_  = \new_[98598]_  & \new_[98595]_ ;
  assign \new_[98602]_  = ~A200 & A199;
  assign \new_[98605]_  = A203 & A201;
  assign \new_[98606]_  = \new_[98605]_  & \new_[98602]_ ;
  assign \new_[98607]_  = \new_[98606]_  & \new_[98599]_ ;
  assign \new_[98610]_  = ~A233 & ~A232;
  assign \new_[98613]_  = ~A268 & ~A266;
  assign \new_[98614]_  = \new_[98613]_  & \new_[98610]_ ;
  assign \new_[98617]_  = A298 & ~A269;
  assign \new_[98620]_  = ~A302 & ~A301;
  assign \new_[98621]_  = \new_[98620]_  & \new_[98617]_ ;
  assign \new_[98622]_  = \new_[98621]_  & \new_[98614]_ ;
  assign \new_[98625]_  = ~A168 & A169;
  assign \new_[98628]_  = A166 & ~A167;
  assign \new_[98629]_  = \new_[98628]_  & \new_[98625]_ ;
  assign \new_[98632]_  = ~A200 & A199;
  assign \new_[98635]_  = A202 & A201;
  assign \new_[98636]_  = \new_[98635]_  & \new_[98632]_ ;
  assign \new_[98637]_  = \new_[98636]_  & \new_[98629]_ ;
  assign \new_[98640]_  = A233 & A232;
  assign \new_[98643]_  = ~A268 & A265;
  assign \new_[98644]_  = \new_[98643]_  & \new_[98640]_ ;
  assign \new_[98647]_  = ~A299 & ~A269;
  assign \new_[98650]_  = ~A302 & ~A301;
  assign \new_[98651]_  = \new_[98650]_  & \new_[98647]_ ;
  assign \new_[98652]_  = \new_[98651]_  & \new_[98644]_ ;
  assign \new_[98655]_  = ~A168 & A169;
  assign \new_[98658]_  = A166 & ~A167;
  assign \new_[98659]_  = \new_[98658]_  & \new_[98655]_ ;
  assign \new_[98662]_  = ~A200 & A199;
  assign \new_[98665]_  = A202 & A201;
  assign \new_[98666]_  = \new_[98665]_  & \new_[98662]_ ;
  assign \new_[98667]_  = \new_[98666]_  & \new_[98659]_ ;
  assign \new_[98670]_  = ~A235 & ~A233;
  assign \new_[98673]_  = A265 & ~A236;
  assign \new_[98674]_  = \new_[98673]_  & \new_[98670]_ ;
  assign \new_[98677]_  = A298 & A266;
  assign \new_[98680]_  = ~A302 & ~A301;
  assign \new_[98681]_  = \new_[98680]_  & \new_[98677]_ ;
  assign \new_[98682]_  = \new_[98681]_  & \new_[98674]_ ;
  assign \new_[98685]_  = ~A168 & A169;
  assign \new_[98688]_  = A166 & ~A167;
  assign \new_[98689]_  = \new_[98688]_  & \new_[98685]_ ;
  assign \new_[98692]_  = ~A200 & A199;
  assign \new_[98695]_  = A202 & A201;
  assign \new_[98696]_  = \new_[98695]_  & \new_[98692]_ ;
  assign \new_[98697]_  = \new_[98696]_  & \new_[98689]_ ;
  assign \new_[98700]_  = ~A235 & ~A233;
  assign \new_[98703]_  = ~A266 & ~A236;
  assign \new_[98704]_  = \new_[98703]_  & \new_[98700]_ ;
  assign \new_[98707]_  = ~A269 & ~A268;
  assign \new_[98710]_  = ~A300 & A298;
  assign \new_[98711]_  = \new_[98710]_  & \new_[98707]_ ;
  assign \new_[98712]_  = \new_[98711]_  & \new_[98704]_ ;
  assign \new_[98715]_  = ~A168 & A169;
  assign \new_[98718]_  = A166 & ~A167;
  assign \new_[98719]_  = \new_[98718]_  & \new_[98715]_ ;
  assign \new_[98722]_  = ~A200 & A199;
  assign \new_[98725]_  = A202 & A201;
  assign \new_[98726]_  = \new_[98725]_  & \new_[98722]_ ;
  assign \new_[98727]_  = \new_[98726]_  & \new_[98719]_ ;
  assign \new_[98730]_  = ~A235 & ~A233;
  assign \new_[98733]_  = ~A266 & ~A236;
  assign \new_[98734]_  = \new_[98733]_  & \new_[98730]_ ;
  assign \new_[98737]_  = ~A269 & ~A268;
  assign \new_[98740]_  = A299 & A298;
  assign \new_[98741]_  = \new_[98740]_  & \new_[98737]_ ;
  assign \new_[98742]_  = \new_[98741]_  & \new_[98734]_ ;
  assign \new_[98745]_  = ~A168 & A169;
  assign \new_[98748]_  = A166 & ~A167;
  assign \new_[98749]_  = \new_[98748]_  & \new_[98745]_ ;
  assign \new_[98752]_  = ~A200 & A199;
  assign \new_[98755]_  = A202 & A201;
  assign \new_[98756]_  = \new_[98755]_  & \new_[98752]_ ;
  assign \new_[98757]_  = \new_[98756]_  & \new_[98749]_ ;
  assign \new_[98760]_  = ~A235 & ~A233;
  assign \new_[98763]_  = ~A266 & ~A236;
  assign \new_[98764]_  = \new_[98763]_  & \new_[98760]_ ;
  assign \new_[98767]_  = ~A269 & ~A268;
  assign \new_[98770]_  = ~A299 & ~A298;
  assign \new_[98771]_  = \new_[98770]_  & \new_[98767]_ ;
  assign \new_[98772]_  = \new_[98771]_  & \new_[98764]_ ;
  assign \new_[98775]_  = ~A168 & A169;
  assign \new_[98778]_  = A166 & ~A167;
  assign \new_[98779]_  = \new_[98778]_  & \new_[98775]_ ;
  assign \new_[98782]_  = ~A200 & A199;
  assign \new_[98785]_  = A202 & A201;
  assign \new_[98786]_  = \new_[98785]_  & \new_[98782]_ ;
  assign \new_[98787]_  = \new_[98786]_  & \new_[98779]_ ;
  assign \new_[98790]_  = ~A235 & ~A233;
  assign \new_[98793]_  = ~A266 & ~A236;
  assign \new_[98794]_  = \new_[98793]_  & \new_[98790]_ ;
  assign \new_[98797]_  = A298 & ~A267;
  assign \new_[98800]_  = ~A302 & ~A301;
  assign \new_[98801]_  = \new_[98800]_  & \new_[98797]_ ;
  assign \new_[98802]_  = \new_[98801]_  & \new_[98794]_ ;
  assign \new_[98805]_  = ~A168 & A169;
  assign \new_[98808]_  = A166 & ~A167;
  assign \new_[98809]_  = \new_[98808]_  & \new_[98805]_ ;
  assign \new_[98812]_  = ~A200 & A199;
  assign \new_[98815]_  = A202 & A201;
  assign \new_[98816]_  = \new_[98815]_  & \new_[98812]_ ;
  assign \new_[98817]_  = \new_[98816]_  & \new_[98809]_ ;
  assign \new_[98820]_  = ~A235 & ~A233;
  assign \new_[98823]_  = ~A265 & ~A236;
  assign \new_[98824]_  = \new_[98823]_  & \new_[98820]_ ;
  assign \new_[98827]_  = A298 & ~A266;
  assign \new_[98830]_  = ~A302 & ~A301;
  assign \new_[98831]_  = \new_[98830]_  & \new_[98827]_ ;
  assign \new_[98832]_  = \new_[98831]_  & \new_[98824]_ ;
  assign \new_[98835]_  = ~A168 & A169;
  assign \new_[98838]_  = A166 & ~A167;
  assign \new_[98839]_  = \new_[98838]_  & \new_[98835]_ ;
  assign \new_[98842]_  = ~A200 & A199;
  assign \new_[98845]_  = A202 & A201;
  assign \new_[98846]_  = \new_[98845]_  & \new_[98842]_ ;
  assign \new_[98847]_  = \new_[98846]_  & \new_[98839]_ ;
  assign \new_[98850]_  = ~A234 & ~A233;
  assign \new_[98853]_  = ~A268 & ~A266;
  assign \new_[98854]_  = \new_[98853]_  & \new_[98850]_ ;
  assign \new_[98857]_  = A298 & ~A269;
  assign \new_[98860]_  = ~A302 & ~A301;
  assign \new_[98861]_  = \new_[98860]_  & \new_[98857]_ ;
  assign \new_[98862]_  = \new_[98861]_  & \new_[98854]_ ;
  assign \new_[98865]_  = ~A168 & A169;
  assign \new_[98868]_  = A166 & ~A167;
  assign \new_[98869]_  = \new_[98868]_  & \new_[98865]_ ;
  assign \new_[98872]_  = ~A200 & A199;
  assign \new_[98875]_  = A202 & A201;
  assign \new_[98876]_  = \new_[98875]_  & \new_[98872]_ ;
  assign \new_[98877]_  = \new_[98876]_  & \new_[98869]_ ;
  assign \new_[98880]_  = ~A233 & A232;
  assign \new_[98883]_  = A235 & A234;
  assign \new_[98884]_  = \new_[98883]_  & \new_[98880]_ ;
  assign \new_[98887]_  = ~A299 & A298;
  assign \new_[98890]_  = A301 & A300;
  assign \new_[98891]_  = \new_[98890]_  & \new_[98887]_ ;
  assign \new_[98892]_  = \new_[98891]_  & \new_[98884]_ ;
  assign \new_[98895]_  = ~A168 & A169;
  assign \new_[98898]_  = A166 & ~A167;
  assign \new_[98899]_  = \new_[98898]_  & \new_[98895]_ ;
  assign \new_[98902]_  = ~A200 & A199;
  assign \new_[98905]_  = A202 & A201;
  assign \new_[98906]_  = \new_[98905]_  & \new_[98902]_ ;
  assign \new_[98907]_  = \new_[98906]_  & \new_[98899]_ ;
  assign \new_[98910]_  = ~A233 & A232;
  assign \new_[98913]_  = A235 & A234;
  assign \new_[98914]_  = \new_[98913]_  & \new_[98910]_ ;
  assign \new_[98917]_  = ~A299 & A298;
  assign \new_[98920]_  = A302 & A300;
  assign \new_[98921]_  = \new_[98920]_  & \new_[98917]_ ;
  assign \new_[98922]_  = \new_[98921]_  & \new_[98914]_ ;
  assign \new_[98925]_  = ~A168 & A169;
  assign \new_[98928]_  = A166 & ~A167;
  assign \new_[98929]_  = \new_[98928]_  & \new_[98925]_ ;
  assign \new_[98932]_  = ~A200 & A199;
  assign \new_[98935]_  = A202 & A201;
  assign \new_[98936]_  = \new_[98935]_  & \new_[98932]_ ;
  assign \new_[98937]_  = \new_[98936]_  & \new_[98929]_ ;
  assign \new_[98940]_  = ~A233 & A232;
  assign \new_[98943]_  = A235 & A234;
  assign \new_[98944]_  = \new_[98943]_  & \new_[98940]_ ;
  assign \new_[98947]_  = ~A266 & A265;
  assign \new_[98950]_  = A268 & A267;
  assign \new_[98951]_  = \new_[98950]_  & \new_[98947]_ ;
  assign \new_[98952]_  = \new_[98951]_  & \new_[98944]_ ;
  assign \new_[98955]_  = ~A168 & A169;
  assign \new_[98958]_  = A166 & ~A167;
  assign \new_[98959]_  = \new_[98958]_  & \new_[98955]_ ;
  assign \new_[98962]_  = ~A200 & A199;
  assign \new_[98965]_  = A202 & A201;
  assign \new_[98966]_  = \new_[98965]_  & \new_[98962]_ ;
  assign \new_[98967]_  = \new_[98966]_  & \new_[98959]_ ;
  assign \new_[98970]_  = ~A233 & A232;
  assign \new_[98973]_  = A235 & A234;
  assign \new_[98974]_  = \new_[98973]_  & \new_[98970]_ ;
  assign \new_[98977]_  = ~A266 & A265;
  assign \new_[98980]_  = A269 & A267;
  assign \new_[98981]_  = \new_[98980]_  & \new_[98977]_ ;
  assign \new_[98982]_  = \new_[98981]_  & \new_[98974]_ ;
  assign \new_[98985]_  = ~A168 & A169;
  assign \new_[98988]_  = A166 & ~A167;
  assign \new_[98989]_  = \new_[98988]_  & \new_[98985]_ ;
  assign \new_[98992]_  = ~A200 & A199;
  assign \new_[98995]_  = A202 & A201;
  assign \new_[98996]_  = \new_[98995]_  & \new_[98992]_ ;
  assign \new_[98997]_  = \new_[98996]_  & \new_[98989]_ ;
  assign \new_[99000]_  = ~A233 & A232;
  assign \new_[99003]_  = A236 & A234;
  assign \new_[99004]_  = \new_[99003]_  & \new_[99000]_ ;
  assign \new_[99007]_  = ~A299 & A298;
  assign \new_[99010]_  = A301 & A300;
  assign \new_[99011]_  = \new_[99010]_  & \new_[99007]_ ;
  assign \new_[99012]_  = \new_[99011]_  & \new_[99004]_ ;
  assign \new_[99015]_  = ~A168 & A169;
  assign \new_[99018]_  = A166 & ~A167;
  assign \new_[99019]_  = \new_[99018]_  & \new_[99015]_ ;
  assign \new_[99022]_  = ~A200 & A199;
  assign \new_[99025]_  = A202 & A201;
  assign \new_[99026]_  = \new_[99025]_  & \new_[99022]_ ;
  assign \new_[99027]_  = \new_[99026]_  & \new_[99019]_ ;
  assign \new_[99030]_  = ~A233 & A232;
  assign \new_[99033]_  = A236 & A234;
  assign \new_[99034]_  = \new_[99033]_  & \new_[99030]_ ;
  assign \new_[99037]_  = ~A299 & A298;
  assign \new_[99040]_  = A302 & A300;
  assign \new_[99041]_  = \new_[99040]_  & \new_[99037]_ ;
  assign \new_[99042]_  = \new_[99041]_  & \new_[99034]_ ;
  assign \new_[99045]_  = ~A168 & A169;
  assign \new_[99048]_  = A166 & ~A167;
  assign \new_[99049]_  = \new_[99048]_  & \new_[99045]_ ;
  assign \new_[99052]_  = ~A200 & A199;
  assign \new_[99055]_  = A202 & A201;
  assign \new_[99056]_  = \new_[99055]_  & \new_[99052]_ ;
  assign \new_[99057]_  = \new_[99056]_  & \new_[99049]_ ;
  assign \new_[99060]_  = ~A233 & A232;
  assign \new_[99063]_  = A236 & A234;
  assign \new_[99064]_  = \new_[99063]_  & \new_[99060]_ ;
  assign \new_[99067]_  = ~A266 & A265;
  assign \new_[99070]_  = A268 & A267;
  assign \new_[99071]_  = \new_[99070]_  & \new_[99067]_ ;
  assign \new_[99072]_  = \new_[99071]_  & \new_[99064]_ ;
  assign \new_[99075]_  = ~A168 & A169;
  assign \new_[99078]_  = A166 & ~A167;
  assign \new_[99079]_  = \new_[99078]_  & \new_[99075]_ ;
  assign \new_[99082]_  = ~A200 & A199;
  assign \new_[99085]_  = A202 & A201;
  assign \new_[99086]_  = \new_[99085]_  & \new_[99082]_ ;
  assign \new_[99087]_  = \new_[99086]_  & \new_[99079]_ ;
  assign \new_[99090]_  = ~A233 & A232;
  assign \new_[99093]_  = A236 & A234;
  assign \new_[99094]_  = \new_[99093]_  & \new_[99090]_ ;
  assign \new_[99097]_  = ~A266 & A265;
  assign \new_[99100]_  = A269 & A267;
  assign \new_[99101]_  = \new_[99100]_  & \new_[99097]_ ;
  assign \new_[99102]_  = \new_[99101]_  & \new_[99094]_ ;
  assign \new_[99105]_  = ~A168 & A169;
  assign \new_[99108]_  = A166 & ~A167;
  assign \new_[99109]_  = \new_[99108]_  & \new_[99105]_ ;
  assign \new_[99112]_  = ~A200 & A199;
  assign \new_[99115]_  = A202 & A201;
  assign \new_[99116]_  = \new_[99115]_  & \new_[99112]_ ;
  assign \new_[99117]_  = \new_[99116]_  & \new_[99109]_ ;
  assign \new_[99120]_  = ~A233 & ~A232;
  assign \new_[99123]_  = ~A268 & ~A266;
  assign \new_[99124]_  = \new_[99123]_  & \new_[99120]_ ;
  assign \new_[99127]_  = A298 & ~A269;
  assign \new_[99130]_  = ~A302 & ~A301;
  assign \new_[99131]_  = \new_[99130]_  & \new_[99127]_ ;
  assign \new_[99132]_  = \new_[99131]_  & \new_[99124]_ ;
  assign \new_[99135]_  = ~A168 & A169;
  assign \new_[99138]_  = A166 & ~A167;
  assign \new_[99139]_  = \new_[99138]_  & \new_[99135]_ ;
  assign \new_[99142]_  = ~A200 & A199;
  assign \new_[99145]_  = A203 & A201;
  assign \new_[99146]_  = \new_[99145]_  & \new_[99142]_ ;
  assign \new_[99147]_  = \new_[99146]_  & \new_[99139]_ ;
  assign \new_[99150]_  = A233 & A232;
  assign \new_[99153]_  = ~A268 & A265;
  assign \new_[99154]_  = \new_[99153]_  & \new_[99150]_ ;
  assign \new_[99157]_  = ~A299 & ~A269;
  assign \new_[99160]_  = ~A302 & ~A301;
  assign \new_[99161]_  = \new_[99160]_  & \new_[99157]_ ;
  assign \new_[99162]_  = \new_[99161]_  & \new_[99154]_ ;
  assign \new_[99165]_  = ~A168 & A169;
  assign \new_[99168]_  = A166 & ~A167;
  assign \new_[99169]_  = \new_[99168]_  & \new_[99165]_ ;
  assign \new_[99172]_  = ~A200 & A199;
  assign \new_[99175]_  = A203 & A201;
  assign \new_[99176]_  = \new_[99175]_  & \new_[99172]_ ;
  assign \new_[99177]_  = \new_[99176]_  & \new_[99169]_ ;
  assign \new_[99180]_  = ~A235 & ~A233;
  assign \new_[99183]_  = A265 & ~A236;
  assign \new_[99184]_  = \new_[99183]_  & \new_[99180]_ ;
  assign \new_[99187]_  = A298 & A266;
  assign \new_[99190]_  = ~A302 & ~A301;
  assign \new_[99191]_  = \new_[99190]_  & \new_[99187]_ ;
  assign \new_[99192]_  = \new_[99191]_  & \new_[99184]_ ;
  assign \new_[99195]_  = ~A168 & A169;
  assign \new_[99198]_  = A166 & ~A167;
  assign \new_[99199]_  = \new_[99198]_  & \new_[99195]_ ;
  assign \new_[99202]_  = ~A200 & A199;
  assign \new_[99205]_  = A203 & A201;
  assign \new_[99206]_  = \new_[99205]_  & \new_[99202]_ ;
  assign \new_[99207]_  = \new_[99206]_  & \new_[99199]_ ;
  assign \new_[99210]_  = ~A235 & ~A233;
  assign \new_[99213]_  = ~A266 & ~A236;
  assign \new_[99214]_  = \new_[99213]_  & \new_[99210]_ ;
  assign \new_[99217]_  = ~A269 & ~A268;
  assign \new_[99220]_  = ~A300 & A298;
  assign \new_[99221]_  = \new_[99220]_  & \new_[99217]_ ;
  assign \new_[99222]_  = \new_[99221]_  & \new_[99214]_ ;
  assign \new_[99225]_  = ~A168 & A169;
  assign \new_[99228]_  = A166 & ~A167;
  assign \new_[99229]_  = \new_[99228]_  & \new_[99225]_ ;
  assign \new_[99232]_  = ~A200 & A199;
  assign \new_[99235]_  = A203 & A201;
  assign \new_[99236]_  = \new_[99235]_  & \new_[99232]_ ;
  assign \new_[99237]_  = \new_[99236]_  & \new_[99229]_ ;
  assign \new_[99240]_  = ~A235 & ~A233;
  assign \new_[99243]_  = ~A266 & ~A236;
  assign \new_[99244]_  = \new_[99243]_  & \new_[99240]_ ;
  assign \new_[99247]_  = ~A269 & ~A268;
  assign \new_[99250]_  = A299 & A298;
  assign \new_[99251]_  = \new_[99250]_  & \new_[99247]_ ;
  assign \new_[99252]_  = \new_[99251]_  & \new_[99244]_ ;
  assign \new_[99255]_  = ~A168 & A169;
  assign \new_[99258]_  = A166 & ~A167;
  assign \new_[99259]_  = \new_[99258]_  & \new_[99255]_ ;
  assign \new_[99262]_  = ~A200 & A199;
  assign \new_[99265]_  = A203 & A201;
  assign \new_[99266]_  = \new_[99265]_  & \new_[99262]_ ;
  assign \new_[99267]_  = \new_[99266]_  & \new_[99259]_ ;
  assign \new_[99270]_  = ~A235 & ~A233;
  assign \new_[99273]_  = ~A266 & ~A236;
  assign \new_[99274]_  = \new_[99273]_  & \new_[99270]_ ;
  assign \new_[99277]_  = ~A269 & ~A268;
  assign \new_[99280]_  = ~A299 & ~A298;
  assign \new_[99281]_  = \new_[99280]_  & \new_[99277]_ ;
  assign \new_[99282]_  = \new_[99281]_  & \new_[99274]_ ;
  assign \new_[99285]_  = ~A168 & A169;
  assign \new_[99288]_  = A166 & ~A167;
  assign \new_[99289]_  = \new_[99288]_  & \new_[99285]_ ;
  assign \new_[99292]_  = ~A200 & A199;
  assign \new_[99295]_  = A203 & A201;
  assign \new_[99296]_  = \new_[99295]_  & \new_[99292]_ ;
  assign \new_[99297]_  = \new_[99296]_  & \new_[99289]_ ;
  assign \new_[99300]_  = ~A235 & ~A233;
  assign \new_[99303]_  = ~A266 & ~A236;
  assign \new_[99304]_  = \new_[99303]_  & \new_[99300]_ ;
  assign \new_[99307]_  = A298 & ~A267;
  assign \new_[99310]_  = ~A302 & ~A301;
  assign \new_[99311]_  = \new_[99310]_  & \new_[99307]_ ;
  assign \new_[99312]_  = \new_[99311]_  & \new_[99304]_ ;
  assign \new_[99315]_  = ~A168 & A169;
  assign \new_[99318]_  = A166 & ~A167;
  assign \new_[99319]_  = \new_[99318]_  & \new_[99315]_ ;
  assign \new_[99322]_  = ~A200 & A199;
  assign \new_[99325]_  = A203 & A201;
  assign \new_[99326]_  = \new_[99325]_  & \new_[99322]_ ;
  assign \new_[99327]_  = \new_[99326]_  & \new_[99319]_ ;
  assign \new_[99330]_  = ~A235 & ~A233;
  assign \new_[99333]_  = ~A265 & ~A236;
  assign \new_[99334]_  = \new_[99333]_  & \new_[99330]_ ;
  assign \new_[99337]_  = A298 & ~A266;
  assign \new_[99340]_  = ~A302 & ~A301;
  assign \new_[99341]_  = \new_[99340]_  & \new_[99337]_ ;
  assign \new_[99342]_  = \new_[99341]_  & \new_[99334]_ ;
  assign \new_[99345]_  = ~A168 & A169;
  assign \new_[99348]_  = A166 & ~A167;
  assign \new_[99349]_  = \new_[99348]_  & \new_[99345]_ ;
  assign \new_[99352]_  = ~A200 & A199;
  assign \new_[99355]_  = A203 & A201;
  assign \new_[99356]_  = \new_[99355]_  & \new_[99352]_ ;
  assign \new_[99357]_  = \new_[99356]_  & \new_[99349]_ ;
  assign \new_[99360]_  = ~A234 & ~A233;
  assign \new_[99363]_  = ~A268 & ~A266;
  assign \new_[99364]_  = \new_[99363]_  & \new_[99360]_ ;
  assign \new_[99367]_  = A298 & ~A269;
  assign \new_[99370]_  = ~A302 & ~A301;
  assign \new_[99371]_  = \new_[99370]_  & \new_[99367]_ ;
  assign \new_[99372]_  = \new_[99371]_  & \new_[99364]_ ;
  assign \new_[99375]_  = ~A168 & A169;
  assign \new_[99378]_  = A166 & ~A167;
  assign \new_[99379]_  = \new_[99378]_  & \new_[99375]_ ;
  assign \new_[99382]_  = ~A200 & A199;
  assign \new_[99385]_  = A203 & A201;
  assign \new_[99386]_  = \new_[99385]_  & \new_[99382]_ ;
  assign \new_[99387]_  = \new_[99386]_  & \new_[99379]_ ;
  assign \new_[99390]_  = ~A233 & A232;
  assign \new_[99393]_  = A235 & A234;
  assign \new_[99394]_  = \new_[99393]_  & \new_[99390]_ ;
  assign \new_[99397]_  = ~A299 & A298;
  assign \new_[99400]_  = A301 & A300;
  assign \new_[99401]_  = \new_[99400]_  & \new_[99397]_ ;
  assign \new_[99402]_  = \new_[99401]_  & \new_[99394]_ ;
  assign \new_[99405]_  = ~A168 & A169;
  assign \new_[99408]_  = A166 & ~A167;
  assign \new_[99409]_  = \new_[99408]_  & \new_[99405]_ ;
  assign \new_[99412]_  = ~A200 & A199;
  assign \new_[99415]_  = A203 & A201;
  assign \new_[99416]_  = \new_[99415]_  & \new_[99412]_ ;
  assign \new_[99417]_  = \new_[99416]_  & \new_[99409]_ ;
  assign \new_[99420]_  = ~A233 & A232;
  assign \new_[99423]_  = A235 & A234;
  assign \new_[99424]_  = \new_[99423]_  & \new_[99420]_ ;
  assign \new_[99427]_  = ~A299 & A298;
  assign \new_[99430]_  = A302 & A300;
  assign \new_[99431]_  = \new_[99430]_  & \new_[99427]_ ;
  assign \new_[99432]_  = \new_[99431]_  & \new_[99424]_ ;
  assign \new_[99435]_  = ~A168 & A169;
  assign \new_[99438]_  = A166 & ~A167;
  assign \new_[99439]_  = \new_[99438]_  & \new_[99435]_ ;
  assign \new_[99442]_  = ~A200 & A199;
  assign \new_[99445]_  = A203 & A201;
  assign \new_[99446]_  = \new_[99445]_  & \new_[99442]_ ;
  assign \new_[99447]_  = \new_[99446]_  & \new_[99439]_ ;
  assign \new_[99450]_  = ~A233 & A232;
  assign \new_[99453]_  = A235 & A234;
  assign \new_[99454]_  = \new_[99453]_  & \new_[99450]_ ;
  assign \new_[99457]_  = ~A266 & A265;
  assign \new_[99460]_  = A268 & A267;
  assign \new_[99461]_  = \new_[99460]_  & \new_[99457]_ ;
  assign \new_[99462]_  = \new_[99461]_  & \new_[99454]_ ;
  assign \new_[99465]_  = ~A168 & A169;
  assign \new_[99468]_  = A166 & ~A167;
  assign \new_[99469]_  = \new_[99468]_  & \new_[99465]_ ;
  assign \new_[99472]_  = ~A200 & A199;
  assign \new_[99475]_  = A203 & A201;
  assign \new_[99476]_  = \new_[99475]_  & \new_[99472]_ ;
  assign \new_[99477]_  = \new_[99476]_  & \new_[99469]_ ;
  assign \new_[99480]_  = ~A233 & A232;
  assign \new_[99483]_  = A235 & A234;
  assign \new_[99484]_  = \new_[99483]_  & \new_[99480]_ ;
  assign \new_[99487]_  = ~A266 & A265;
  assign \new_[99490]_  = A269 & A267;
  assign \new_[99491]_  = \new_[99490]_  & \new_[99487]_ ;
  assign \new_[99492]_  = \new_[99491]_  & \new_[99484]_ ;
  assign \new_[99495]_  = ~A168 & A169;
  assign \new_[99498]_  = A166 & ~A167;
  assign \new_[99499]_  = \new_[99498]_  & \new_[99495]_ ;
  assign \new_[99502]_  = ~A200 & A199;
  assign \new_[99505]_  = A203 & A201;
  assign \new_[99506]_  = \new_[99505]_  & \new_[99502]_ ;
  assign \new_[99507]_  = \new_[99506]_  & \new_[99499]_ ;
  assign \new_[99510]_  = ~A233 & A232;
  assign \new_[99513]_  = A236 & A234;
  assign \new_[99514]_  = \new_[99513]_  & \new_[99510]_ ;
  assign \new_[99517]_  = ~A299 & A298;
  assign \new_[99520]_  = A301 & A300;
  assign \new_[99521]_  = \new_[99520]_  & \new_[99517]_ ;
  assign \new_[99522]_  = \new_[99521]_  & \new_[99514]_ ;
  assign \new_[99525]_  = ~A168 & A169;
  assign \new_[99528]_  = A166 & ~A167;
  assign \new_[99529]_  = \new_[99528]_  & \new_[99525]_ ;
  assign \new_[99532]_  = ~A200 & A199;
  assign \new_[99535]_  = A203 & A201;
  assign \new_[99536]_  = \new_[99535]_  & \new_[99532]_ ;
  assign \new_[99537]_  = \new_[99536]_  & \new_[99529]_ ;
  assign \new_[99540]_  = ~A233 & A232;
  assign \new_[99543]_  = A236 & A234;
  assign \new_[99544]_  = \new_[99543]_  & \new_[99540]_ ;
  assign \new_[99547]_  = ~A299 & A298;
  assign \new_[99550]_  = A302 & A300;
  assign \new_[99551]_  = \new_[99550]_  & \new_[99547]_ ;
  assign \new_[99552]_  = \new_[99551]_  & \new_[99544]_ ;
  assign \new_[99555]_  = ~A168 & A169;
  assign \new_[99558]_  = A166 & ~A167;
  assign \new_[99559]_  = \new_[99558]_  & \new_[99555]_ ;
  assign \new_[99562]_  = ~A200 & A199;
  assign \new_[99565]_  = A203 & A201;
  assign \new_[99566]_  = \new_[99565]_  & \new_[99562]_ ;
  assign \new_[99567]_  = \new_[99566]_  & \new_[99559]_ ;
  assign \new_[99570]_  = ~A233 & A232;
  assign \new_[99573]_  = A236 & A234;
  assign \new_[99574]_  = \new_[99573]_  & \new_[99570]_ ;
  assign \new_[99577]_  = ~A266 & A265;
  assign \new_[99580]_  = A268 & A267;
  assign \new_[99581]_  = \new_[99580]_  & \new_[99577]_ ;
  assign \new_[99582]_  = \new_[99581]_  & \new_[99574]_ ;
  assign \new_[99585]_  = ~A168 & A169;
  assign \new_[99588]_  = A166 & ~A167;
  assign \new_[99589]_  = \new_[99588]_  & \new_[99585]_ ;
  assign \new_[99592]_  = ~A200 & A199;
  assign \new_[99595]_  = A203 & A201;
  assign \new_[99596]_  = \new_[99595]_  & \new_[99592]_ ;
  assign \new_[99597]_  = \new_[99596]_  & \new_[99589]_ ;
  assign \new_[99600]_  = ~A233 & A232;
  assign \new_[99603]_  = A236 & A234;
  assign \new_[99604]_  = \new_[99603]_  & \new_[99600]_ ;
  assign \new_[99607]_  = ~A266 & A265;
  assign \new_[99610]_  = A269 & A267;
  assign \new_[99611]_  = \new_[99610]_  & \new_[99607]_ ;
  assign \new_[99612]_  = \new_[99611]_  & \new_[99604]_ ;
  assign \new_[99615]_  = ~A168 & A169;
  assign \new_[99618]_  = A166 & ~A167;
  assign \new_[99619]_  = \new_[99618]_  & \new_[99615]_ ;
  assign \new_[99622]_  = ~A200 & A199;
  assign \new_[99625]_  = A203 & A201;
  assign \new_[99626]_  = \new_[99625]_  & \new_[99622]_ ;
  assign \new_[99627]_  = \new_[99626]_  & \new_[99619]_ ;
  assign \new_[99630]_  = ~A233 & ~A232;
  assign \new_[99633]_  = ~A268 & ~A266;
  assign \new_[99634]_  = \new_[99633]_  & \new_[99630]_ ;
  assign \new_[99637]_  = A298 & ~A269;
  assign \new_[99640]_  = ~A302 & ~A301;
  assign \new_[99641]_  = \new_[99640]_  & \new_[99637]_ ;
  assign \new_[99642]_  = \new_[99641]_  & \new_[99634]_ ;
  assign \new_[99645]_  = A169 & A170;
  assign \new_[99648]_  = A199 & ~A168;
  assign \new_[99649]_  = \new_[99648]_  & \new_[99645]_ ;
  assign \new_[99652]_  = A201 & ~A200;
  assign \new_[99655]_  = ~A233 & A202;
  assign \new_[99656]_  = \new_[99655]_  & \new_[99652]_ ;
  assign \new_[99657]_  = \new_[99656]_  & \new_[99649]_ ;
  assign \new_[99660]_  = ~A236 & ~A235;
  assign \new_[99663]_  = ~A268 & ~A266;
  assign \new_[99664]_  = \new_[99663]_  & \new_[99660]_ ;
  assign \new_[99667]_  = A298 & ~A269;
  assign \new_[99670]_  = ~A302 & ~A301;
  assign \new_[99671]_  = \new_[99670]_  & \new_[99667]_ ;
  assign \new_[99672]_  = \new_[99671]_  & \new_[99664]_ ;
  assign \new_[99675]_  = A169 & A170;
  assign \new_[99678]_  = A199 & ~A168;
  assign \new_[99679]_  = \new_[99678]_  & \new_[99675]_ ;
  assign \new_[99682]_  = A201 & ~A200;
  assign \new_[99685]_  = ~A233 & A203;
  assign \new_[99686]_  = \new_[99685]_  & \new_[99682]_ ;
  assign \new_[99687]_  = \new_[99686]_  & \new_[99679]_ ;
  assign \new_[99690]_  = ~A236 & ~A235;
  assign \new_[99693]_  = ~A268 & ~A266;
  assign \new_[99694]_  = \new_[99693]_  & \new_[99690]_ ;
  assign \new_[99697]_  = A298 & ~A269;
  assign \new_[99700]_  = ~A302 & ~A301;
  assign \new_[99701]_  = \new_[99700]_  & \new_[99697]_ ;
  assign \new_[99702]_  = \new_[99701]_  & \new_[99694]_ ;
  assign \new_[99705]_  = A169 & ~A170;
  assign \new_[99708]_  = A166 & A167;
  assign \new_[99709]_  = \new_[99708]_  & \new_[99705]_ ;
  assign \new_[99712]_  = ~A202 & ~A200;
  assign \new_[99715]_  = ~A233 & ~A203;
  assign \new_[99716]_  = \new_[99715]_  & \new_[99712]_ ;
  assign \new_[99717]_  = \new_[99716]_  & \new_[99709]_ ;
  assign \new_[99720]_  = ~A236 & ~A235;
  assign \new_[99723]_  = ~A268 & ~A266;
  assign \new_[99724]_  = \new_[99723]_  & \new_[99720]_ ;
  assign \new_[99727]_  = A298 & ~A269;
  assign \new_[99730]_  = ~A302 & ~A301;
  assign \new_[99731]_  = \new_[99730]_  & \new_[99727]_ ;
  assign \new_[99732]_  = \new_[99731]_  & \new_[99724]_ ;
  assign \new_[99735]_  = A169 & ~A170;
  assign \new_[99738]_  = ~A166 & ~A167;
  assign \new_[99739]_  = \new_[99738]_  & \new_[99735]_ ;
  assign \new_[99742]_  = ~A202 & ~A200;
  assign \new_[99745]_  = ~A233 & ~A203;
  assign \new_[99746]_  = \new_[99745]_  & \new_[99742]_ ;
  assign \new_[99747]_  = \new_[99746]_  & \new_[99739]_ ;
  assign \new_[99750]_  = ~A236 & ~A235;
  assign \new_[99753]_  = ~A268 & ~A266;
  assign \new_[99754]_  = \new_[99753]_  & \new_[99750]_ ;
  assign \new_[99757]_  = A298 & ~A269;
  assign \new_[99760]_  = ~A302 & ~A301;
  assign \new_[99761]_  = \new_[99760]_  & \new_[99757]_ ;
  assign \new_[99762]_  = \new_[99761]_  & \new_[99754]_ ;
  assign \new_[99765]_  = ~A167 & ~A169;
  assign \new_[99768]_  = A199 & ~A166;
  assign \new_[99769]_  = \new_[99768]_  & \new_[99765]_ ;
  assign \new_[99772]_  = A201 & ~A200;
  assign \new_[99775]_  = ~A233 & A202;
  assign \new_[99776]_  = \new_[99775]_  & \new_[99772]_ ;
  assign \new_[99777]_  = \new_[99776]_  & \new_[99769]_ ;
  assign \new_[99780]_  = ~A236 & ~A235;
  assign \new_[99783]_  = ~A268 & ~A266;
  assign \new_[99784]_  = \new_[99783]_  & \new_[99780]_ ;
  assign \new_[99787]_  = A298 & ~A269;
  assign \new_[99790]_  = ~A302 & ~A301;
  assign \new_[99791]_  = \new_[99790]_  & \new_[99787]_ ;
  assign \new_[99792]_  = \new_[99791]_  & \new_[99784]_ ;
  assign \new_[99795]_  = ~A167 & ~A169;
  assign \new_[99798]_  = A199 & ~A166;
  assign \new_[99799]_  = \new_[99798]_  & \new_[99795]_ ;
  assign \new_[99802]_  = A201 & ~A200;
  assign \new_[99805]_  = ~A233 & A203;
  assign \new_[99806]_  = \new_[99805]_  & \new_[99802]_ ;
  assign \new_[99807]_  = \new_[99806]_  & \new_[99799]_ ;
  assign \new_[99810]_  = ~A236 & ~A235;
  assign \new_[99813]_  = ~A268 & ~A266;
  assign \new_[99814]_  = \new_[99813]_  & \new_[99810]_ ;
  assign \new_[99817]_  = A298 & ~A269;
  assign \new_[99820]_  = ~A302 & ~A301;
  assign \new_[99821]_  = \new_[99820]_  & \new_[99817]_ ;
  assign \new_[99822]_  = \new_[99821]_  & \new_[99814]_ ;
  assign \new_[99825]_  = ~A168 & ~A169;
  assign \new_[99828]_  = A166 & A167;
  assign \new_[99829]_  = \new_[99828]_  & \new_[99825]_ ;
  assign \new_[99832]_  = ~A200 & A199;
  assign \new_[99835]_  = A202 & A201;
  assign \new_[99836]_  = \new_[99835]_  & \new_[99832]_ ;
  assign \new_[99837]_  = \new_[99836]_  & \new_[99829]_ ;
  assign \new_[99840]_  = A233 & A232;
  assign \new_[99843]_  = ~A268 & A265;
  assign \new_[99844]_  = \new_[99843]_  & \new_[99840]_ ;
  assign \new_[99847]_  = ~A299 & ~A269;
  assign \new_[99850]_  = ~A302 & ~A301;
  assign \new_[99851]_  = \new_[99850]_  & \new_[99847]_ ;
  assign \new_[99852]_  = \new_[99851]_  & \new_[99844]_ ;
  assign \new_[99855]_  = ~A168 & ~A169;
  assign \new_[99858]_  = A166 & A167;
  assign \new_[99859]_  = \new_[99858]_  & \new_[99855]_ ;
  assign \new_[99862]_  = ~A200 & A199;
  assign \new_[99865]_  = A202 & A201;
  assign \new_[99866]_  = \new_[99865]_  & \new_[99862]_ ;
  assign \new_[99867]_  = \new_[99866]_  & \new_[99859]_ ;
  assign \new_[99870]_  = ~A235 & ~A233;
  assign \new_[99873]_  = A265 & ~A236;
  assign \new_[99874]_  = \new_[99873]_  & \new_[99870]_ ;
  assign \new_[99877]_  = A298 & A266;
  assign \new_[99880]_  = ~A302 & ~A301;
  assign \new_[99881]_  = \new_[99880]_  & \new_[99877]_ ;
  assign \new_[99882]_  = \new_[99881]_  & \new_[99874]_ ;
  assign \new_[99885]_  = ~A168 & ~A169;
  assign \new_[99888]_  = A166 & A167;
  assign \new_[99889]_  = \new_[99888]_  & \new_[99885]_ ;
  assign \new_[99892]_  = ~A200 & A199;
  assign \new_[99895]_  = A202 & A201;
  assign \new_[99896]_  = \new_[99895]_  & \new_[99892]_ ;
  assign \new_[99897]_  = \new_[99896]_  & \new_[99889]_ ;
  assign \new_[99900]_  = ~A235 & ~A233;
  assign \new_[99903]_  = ~A266 & ~A236;
  assign \new_[99904]_  = \new_[99903]_  & \new_[99900]_ ;
  assign \new_[99907]_  = ~A269 & ~A268;
  assign \new_[99910]_  = ~A300 & A298;
  assign \new_[99911]_  = \new_[99910]_  & \new_[99907]_ ;
  assign \new_[99912]_  = \new_[99911]_  & \new_[99904]_ ;
  assign \new_[99915]_  = ~A168 & ~A169;
  assign \new_[99918]_  = A166 & A167;
  assign \new_[99919]_  = \new_[99918]_  & \new_[99915]_ ;
  assign \new_[99922]_  = ~A200 & A199;
  assign \new_[99925]_  = A202 & A201;
  assign \new_[99926]_  = \new_[99925]_  & \new_[99922]_ ;
  assign \new_[99927]_  = \new_[99926]_  & \new_[99919]_ ;
  assign \new_[99930]_  = ~A235 & ~A233;
  assign \new_[99933]_  = ~A266 & ~A236;
  assign \new_[99934]_  = \new_[99933]_  & \new_[99930]_ ;
  assign \new_[99937]_  = ~A269 & ~A268;
  assign \new_[99940]_  = A299 & A298;
  assign \new_[99941]_  = \new_[99940]_  & \new_[99937]_ ;
  assign \new_[99942]_  = \new_[99941]_  & \new_[99934]_ ;
  assign \new_[99945]_  = ~A168 & ~A169;
  assign \new_[99948]_  = A166 & A167;
  assign \new_[99949]_  = \new_[99948]_  & \new_[99945]_ ;
  assign \new_[99952]_  = ~A200 & A199;
  assign \new_[99955]_  = A202 & A201;
  assign \new_[99956]_  = \new_[99955]_  & \new_[99952]_ ;
  assign \new_[99957]_  = \new_[99956]_  & \new_[99949]_ ;
  assign \new_[99960]_  = ~A235 & ~A233;
  assign \new_[99963]_  = ~A266 & ~A236;
  assign \new_[99964]_  = \new_[99963]_  & \new_[99960]_ ;
  assign \new_[99967]_  = ~A269 & ~A268;
  assign \new_[99970]_  = ~A299 & ~A298;
  assign \new_[99971]_  = \new_[99970]_  & \new_[99967]_ ;
  assign \new_[99972]_  = \new_[99971]_  & \new_[99964]_ ;
  assign \new_[99975]_  = ~A168 & ~A169;
  assign \new_[99978]_  = A166 & A167;
  assign \new_[99979]_  = \new_[99978]_  & \new_[99975]_ ;
  assign \new_[99982]_  = ~A200 & A199;
  assign \new_[99985]_  = A202 & A201;
  assign \new_[99986]_  = \new_[99985]_  & \new_[99982]_ ;
  assign \new_[99987]_  = \new_[99986]_  & \new_[99979]_ ;
  assign \new_[99990]_  = ~A235 & ~A233;
  assign \new_[99993]_  = ~A266 & ~A236;
  assign \new_[99994]_  = \new_[99993]_  & \new_[99990]_ ;
  assign \new_[99997]_  = A298 & ~A267;
  assign \new_[100000]_  = ~A302 & ~A301;
  assign \new_[100001]_  = \new_[100000]_  & \new_[99997]_ ;
  assign \new_[100002]_  = \new_[100001]_  & \new_[99994]_ ;
  assign \new_[100005]_  = ~A168 & ~A169;
  assign \new_[100008]_  = A166 & A167;
  assign \new_[100009]_  = \new_[100008]_  & \new_[100005]_ ;
  assign \new_[100012]_  = ~A200 & A199;
  assign \new_[100015]_  = A202 & A201;
  assign \new_[100016]_  = \new_[100015]_  & \new_[100012]_ ;
  assign \new_[100017]_  = \new_[100016]_  & \new_[100009]_ ;
  assign \new_[100020]_  = ~A235 & ~A233;
  assign \new_[100023]_  = ~A265 & ~A236;
  assign \new_[100024]_  = \new_[100023]_  & \new_[100020]_ ;
  assign \new_[100027]_  = A298 & ~A266;
  assign \new_[100030]_  = ~A302 & ~A301;
  assign \new_[100031]_  = \new_[100030]_  & \new_[100027]_ ;
  assign \new_[100032]_  = \new_[100031]_  & \new_[100024]_ ;
  assign \new_[100035]_  = ~A168 & ~A169;
  assign \new_[100038]_  = A166 & A167;
  assign \new_[100039]_  = \new_[100038]_  & \new_[100035]_ ;
  assign \new_[100042]_  = ~A200 & A199;
  assign \new_[100045]_  = A202 & A201;
  assign \new_[100046]_  = \new_[100045]_  & \new_[100042]_ ;
  assign \new_[100047]_  = \new_[100046]_  & \new_[100039]_ ;
  assign \new_[100050]_  = ~A234 & ~A233;
  assign \new_[100053]_  = ~A268 & ~A266;
  assign \new_[100054]_  = \new_[100053]_  & \new_[100050]_ ;
  assign \new_[100057]_  = A298 & ~A269;
  assign \new_[100060]_  = ~A302 & ~A301;
  assign \new_[100061]_  = \new_[100060]_  & \new_[100057]_ ;
  assign \new_[100062]_  = \new_[100061]_  & \new_[100054]_ ;
  assign \new_[100065]_  = ~A168 & ~A169;
  assign \new_[100068]_  = A166 & A167;
  assign \new_[100069]_  = \new_[100068]_  & \new_[100065]_ ;
  assign \new_[100072]_  = ~A200 & A199;
  assign \new_[100075]_  = A202 & A201;
  assign \new_[100076]_  = \new_[100075]_  & \new_[100072]_ ;
  assign \new_[100077]_  = \new_[100076]_  & \new_[100069]_ ;
  assign \new_[100080]_  = ~A233 & A232;
  assign \new_[100083]_  = A235 & A234;
  assign \new_[100084]_  = \new_[100083]_  & \new_[100080]_ ;
  assign \new_[100087]_  = ~A299 & A298;
  assign \new_[100090]_  = A301 & A300;
  assign \new_[100091]_  = \new_[100090]_  & \new_[100087]_ ;
  assign \new_[100092]_  = \new_[100091]_  & \new_[100084]_ ;
  assign \new_[100095]_  = ~A168 & ~A169;
  assign \new_[100098]_  = A166 & A167;
  assign \new_[100099]_  = \new_[100098]_  & \new_[100095]_ ;
  assign \new_[100102]_  = ~A200 & A199;
  assign \new_[100105]_  = A202 & A201;
  assign \new_[100106]_  = \new_[100105]_  & \new_[100102]_ ;
  assign \new_[100107]_  = \new_[100106]_  & \new_[100099]_ ;
  assign \new_[100110]_  = ~A233 & A232;
  assign \new_[100113]_  = A235 & A234;
  assign \new_[100114]_  = \new_[100113]_  & \new_[100110]_ ;
  assign \new_[100117]_  = ~A299 & A298;
  assign \new_[100120]_  = A302 & A300;
  assign \new_[100121]_  = \new_[100120]_  & \new_[100117]_ ;
  assign \new_[100122]_  = \new_[100121]_  & \new_[100114]_ ;
  assign \new_[100125]_  = ~A168 & ~A169;
  assign \new_[100128]_  = A166 & A167;
  assign \new_[100129]_  = \new_[100128]_  & \new_[100125]_ ;
  assign \new_[100132]_  = ~A200 & A199;
  assign \new_[100135]_  = A202 & A201;
  assign \new_[100136]_  = \new_[100135]_  & \new_[100132]_ ;
  assign \new_[100137]_  = \new_[100136]_  & \new_[100129]_ ;
  assign \new_[100140]_  = ~A233 & A232;
  assign \new_[100143]_  = A235 & A234;
  assign \new_[100144]_  = \new_[100143]_  & \new_[100140]_ ;
  assign \new_[100147]_  = ~A266 & A265;
  assign \new_[100150]_  = A268 & A267;
  assign \new_[100151]_  = \new_[100150]_  & \new_[100147]_ ;
  assign \new_[100152]_  = \new_[100151]_  & \new_[100144]_ ;
  assign \new_[100155]_  = ~A168 & ~A169;
  assign \new_[100158]_  = A166 & A167;
  assign \new_[100159]_  = \new_[100158]_  & \new_[100155]_ ;
  assign \new_[100162]_  = ~A200 & A199;
  assign \new_[100165]_  = A202 & A201;
  assign \new_[100166]_  = \new_[100165]_  & \new_[100162]_ ;
  assign \new_[100167]_  = \new_[100166]_  & \new_[100159]_ ;
  assign \new_[100170]_  = ~A233 & A232;
  assign \new_[100173]_  = A235 & A234;
  assign \new_[100174]_  = \new_[100173]_  & \new_[100170]_ ;
  assign \new_[100177]_  = ~A266 & A265;
  assign \new_[100180]_  = A269 & A267;
  assign \new_[100181]_  = \new_[100180]_  & \new_[100177]_ ;
  assign \new_[100182]_  = \new_[100181]_  & \new_[100174]_ ;
  assign \new_[100185]_  = ~A168 & ~A169;
  assign \new_[100188]_  = A166 & A167;
  assign \new_[100189]_  = \new_[100188]_  & \new_[100185]_ ;
  assign \new_[100192]_  = ~A200 & A199;
  assign \new_[100195]_  = A202 & A201;
  assign \new_[100196]_  = \new_[100195]_  & \new_[100192]_ ;
  assign \new_[100197]_  = \new_[100196]_  & \new_[100189]_ ;
  assign \new_[100200]_  = ~A233 & A232;
  assign \new_[100203]_  = A236 & A234;
  assign \new_[100204]_  = \new_[100203]_  & \new_[100200]_ ;
  assign \new_[100207]_  = ~A299 & A298;
  assign \new_[100210]_  = A301 & A300;
  assign \new_[100211]_  = \new_[100210]_  & \new_[100207]_ ;
  assign \new_[100212]_  = \new_[100211]_  & \new_[100204]_ ;
  assign \new_[100215]_  = ~A168 & ~A169;
  assign \new_[100218]_  = A166 & A167;
  assign \new_[100219]_  = \new_[100218]_  & \new_[100215]_ ;
  assign \new_[100222]_  = ~A200 & A199;
  assign \new_[100225]_  = A202 & A201;
  assign \new_[100226]_  = \new_[100225]_  & \new_[100222]_ ;
  assign \new_[100227]_  = \new_[100226]_  & \new_[100219]_ ;
  assign \new_[100230]_  = ~A233 & A232;
  assign \new_[100233]_  = A236 & A234;
  assign \new_[100234]_  = \new_[100233]_  & \new_[100230]_ ;
  assign \new_[100237]_  = ~A299 & A298;
  assign \new_[100240]_  = A302 & A300;
  assign \new_[100241]_  = \new_[100240]_  & \new_[100237]_ ;
  assign \new_[100242]_  = \new_[100241]_  & \new_[100234]_ ;
  assign \new_[100245]_  = ~A168 & ~A169;
  assign \new_[100248]_  = A166 & A167;
  assign \new_[100249]_  = \new_[100248]_  & \new_[100245]_ ;
  assign \new_[100252]_  = ~A200 & A199;
  assign \new_[100255]_  = A202 & A201;
  assign \new_[100256]_  = \new_[100255]_  & \new_[100252]_ ;
  assign \new_[100257]_  = \new_[100256]_  & \new_[100249]_ ;
  assign \new_[100260]_  = ~A233 & A232;
  assign \new_[100263]_  = A236 & A234;
  assign \new_[100264]_  = \new_[100263]_  & \new_[100260]_ ;
  assign \new_[100267]_  = ~A266 & A265;
  assign \new_[100270]_  = A268 & A267;
  assign \new_[100271]_  = \new_[100270]_  & \new_[100267]_ ;
  assign \new_[100272]_  = \new_[100271]_  & \new_[100264]_ ;
  assign \new_[100275]_  = ~A168 & ~A169;
  assign \new_[100278]_  = A166 & A167;
  assign \new_[100279]_  = \new_[100278]_  & \new_[100275]_ ;
  assign \new_[100282]_  = ~A200 & A199;
  assign \new_[100285]_  = A202 & A201;
  assign \new_[100286]_  = \new_[100285]_  & \new_[100282]_ ;
  assign \new_[100287]_  = \new_[100286]_  & \new_[100279]_ ;
  assign \new_[100290]_  = ~A233 & A232;
  assign \new_[100293]_  = A236 & A234;
  assign \new_[100294]_  = \new_[100293]_  & \new_[100290]_ ;
  assign \new_[100297]_  = ~A266 & A265;
  assign \new_[100300]_  = A269 & A267;
  assign \new_[100301]_  = \new_[100300]_  & \new_[100297]_ ;
  assign \new_[100302]_  = \new_[100301]_  & \new_[100294]_ ;
  assign \new_[100305]_  = ~A168 & ~A169;
  assign \new_[100308]_  = A166 & A167;
  assign \new_[100309]_  = \new_[100308]_  & \new_[100305]_ ;
  assign \new_[100312]_  = ~A200 & A199;
  assign \new_[100315]_  = A202 & A201;
  assign \new_[100316]_  = \new_[100315]_  & \new_[100312]_ ;
  assign \new_[100317]_  = \new_[100316]_  & \new_[100309]_ ;
  assign \new_[100320]_  = ~A233 & ~A232;
  assign \new_[100323]_  = ~A268 & ~A266;
  assign \new_[100324]_  = \new_[100323]_  & \new_[100320]_ ;
  assign \new_[100327]_  = A298 & ~A269;
  assign \new_[100330]_  = ~A302 & ~A301;
  assign \new_[100331]_  = \new_[100330]_  & \new_[100327]_ ;
  assign \new_[100332]_  = \new_[100331]_  & \new_[100324]_ ;
  assign \new_[100335]_  = ~A168 & ~A169;
  assign \new_[100338]_  = A166 & A167;
  assign \new_[100339]_  = \new_[100338]_  & \new_[100335]_ ;
  assign \new_[100342]_  = ~A200 & A199;
  assign \new_[100345]_  = A203 & A201;
  assign \new_[100346]_  = \new_[100345]_  & \new_[100342]_ ;
  assign \new_[100347]_  = \new_[100346]_  & \new_[100339]_ ;
  assign \new_[100350]_  = A233 & A232;
  assign \new_[100353]_  = ~A268 & A265;
  assign \new_[100354]_  = \new_[100353]_  & \new_[100350]_ ;
  assign \new_[100357]_  = ~A299 & ~A269;
  assign \new_[100360]_  = ~A302 & ~A301;
  assign \new_[100361]_  = \new_[100360]_  & \new_[100357]_ ;
  assign \new_[100362]_  = \new_[100361]_  & \new_[100354]_ ;
  assign \new_[100365]_  = ~A168 & ~A169;
  assign \new_[100368]_  = A166 & A167;
  assign \new_[100369]_  = \new_[100368]_  & \new_[100365]_ ;
  assign \new_[100372]_  = ~A200 & A199;
  assign \new_[100375]_  = A203 & A201;
  assign \new_[100376]_  = \new_[100375]_  & \new_[100372]_ ;
  assign \new_[100377]_  = \new_[100376]_  & \new_[100369]_ ;
  assign \new_[100380]_  = ~A235 & ~A233;
  assign \new_[100383]_  = A265 & ~A236;
  assign \new_[100384]_  = \new_[100383]_  & \new_[100380]_ ;
  assign \new_[100387]_  = A298 & A266;
  assign \new_[100390]_  = ~A302 & ~A301;
  assign \new_[100391]_  = \new_[100390]_  & \new_[100387]_ ;
  assign \new_[100392]_  = \new_[100391]_  & \new_[100384]_ ;
  assign \new_[100395]_  = ~A168 & ~A169;
  assign \new_[100398]_  = A166 & A167;
  assign \new_[100399]_  = \new_[100398]_  & \new_[100395]_ ;
  assign \new_[100402]_  = ~A200 & A199;
  assign \new_[100405]_  = A203 & A201;
  assign \new_[100406]_  = \new_[100405]_  & \new_[100402]_ ;
  assign \new_[100407]_  = \new_[100406]_  & \new_[100399]_ ;
  assign \new_[100410]_  = ~A235 & ~A233;
  assign \new_[100413]_  = ~A266 & ~A236;
  assign \new_[100414]_  = \new_[100413]_  & \new_[100410]_ ;
  assign \new_[100417]_  = ~A269 & ~A268;
  assign \new_[100420]_  = ~A300 & A298;
  assign \new_[100421]_  = \new_[100420]_  & \new_[100417]_ ;
  assign \new_[100422]_  = \new_[100421]_  & \new_[100414]_ ;
  assign \new_[100425]_  = ~A168 & ~A169;
  assign \new_[100428]_  = A166 & A167;
  assign \new_[100429]_  = \new_[100428]_  & \new_[100425]_ ;
  assign \new_[100432]_  = ~A200 & A199;
  assign \new_[100435]_  = A203 & A201;
  assign \new_[100436]_  = \new_[100435]_  & \new_[100432]_ ;
  assign \new_[100437]_  = \new_[100436]_  & \new_[100429]_ ;
  assign \new_[100440]_  = ~A235 & ~A233;
  assign \new_[100443]_  = ~A266 & ~A236;
  assign \new_[100444]_  = \new_[100443]_  & \new_[100440]_ ;
  assign \new_[100447]_  = ~A269 & ~A268;
  assign \new_[100450]_  = A299 & A298;
  assign \new_[100451]_  = \new_[100450]_  & \new_[100447]_ ;
  assign \new_[100452]_  = \new_[100451]_  & \new_[100444]_ ;
  assign \new_[100455]_  = ~A168 & ~A169;
  assign \new_[100458]_  = A166 & A167;
  assign \new_[100459]_  = \new_[100458]_  & \new_[100455]_ ;
  assign \new_[100462]_  = ~A200 & A199;
  assign \new_[100465]_  = A203 & A201;
  assign \new_[100466]_  = \new_[100465]_  & \new_[100462]_ ;
  assign \new_[100467]_  = \new_[100466]_  & \new_[100459]_ ;
  assign \new_[100470]_  = ~A235 & ~A233;
  assign \new_[100473]_  = ~A266 & ~A236;
  assign \new_[100474]_  = \new_[100473]_  & \new_[100470]_ ;
  assign \new_[100477]_  = ~A269 & ~A268;
  assign \new_[100480]_  = ~A299 & ~A298;
  assign \new_[100481]_  = \new_[100480]_  & \new_[100477]_ ;
  assign \new_[100482]_  = \new_[100481]_  & \new_[100474]_ ;
  assign \new_[100485]_  = ~A168 & ~A169;
  assign \new_[100488]_  = A166 & A167;
  assign \new_[100489]_  = \new_[100488]_  & \new_[100485]_ ;
  assign \new_[100492]_  = ~A200 & A199;
  assign \new_[100495]_  = A203 & A201;
  assign \new_[100496]_  = \new_[100495]_  & \new_[100492]_ ;
  assign \new_[100497]_  = \new_[100496]_  & \new_[100489]_ ;
  assign \new_[100500]_  = ~A235 & ~A233;
  assign \new_[100503]_  = ~A266 & ~A236;
  assign \new_[100504]_  = \new_[100503]_  & \new_[100500]_ ;
  assign \new_[100507]_  = A298 & ~A267;
  assign \new_[100510]_  = ~A302 & ~A301;
  assign \new_[100511]_  = \new_[100510]_  & \new_[100507]_ ;
  assign \new_[100512]_  = \new_[100511]_  & \new_[100504]_ ;
  assign \new_[100515]_  = ~A168 & ~A169;
  assign \new_[100518]_  = A166 & A167;
  assign \new_[100519]_  = \new_[100518]_  & \new_[100515]_ ;
  assign \new_[100522]_  = ~A200 & A199;
  assign \new_[100525]_  = A203 & A201;
  assign \new_[100526]_  = \new_[100525]_  & \new_[100522]_ ;
  assign \new_[100527]_  = \new_[100526]_  & \new_[100519]_ ;
  assign \new_[100530]_  = ~A235 & ~A233;
  assign \new_[100533]_  = ~A265 & ~A236;
  assign \new_[100534]_  = \new_[100533]_  & \new_[100530]_ ;
  assign \new_[100537]_  = A298 & ~A266;
  assign \new_[100540]_  = ~A302 & ~A301;
  assign \new_[100541]_  = \new_[100540]_  & \new_[100537]_ ;
  assign \new_[100542]_  = \new_[100541]_  & \new_[100534]_ ;
  assign \new_[100545]_  = ~A168 & ~A169;
  assign \new_[100548]_  = A166 & A167;
  assign \new_[100549]_  = \new_[100548]_  & \new_[100545]_ ;
  assign \new_[100552]_  = ~A200 & A199;
  assign \new_[100555]_  = A203 & A201;
  assign \new_[100556]_  = \new_[100555]_  & \new_[100552]_ ;
  assign \new_[100557]_  = \new_[100556]_  & \new_[100549]_ ;
  assign \new_[100560]_  = ~A234 & ~A233;
  assign \new_[100563]_  = ~A268 & ~A266;
  assign \new_[100564]_  = \new_[100563]_  & \new_[100560]_ ;
  assign \new_[100567]_  = A298 & ~A269;
  assign \new_[100570]_  = ~A302 & ~A301;
  assign \new_[100571]_  = \new_[100570]_  & \new_[100567]_ ;
  assign \new_[100572]_  = \new_[100571]_  & \new_[100564]_ ;
  assign \new_[100575]_  = ~A168 & ~A169;
  assign \new_[100578]_  = A166 & A167;
  assign \new_[100579]_  = \new_[100578]_  & \new_[100575]_ ;
  assign \new_[100582]_  = ~A200 & A199;
  assign \new_[100585]_  = A203 & A201;
  assign \new_[100586]_  = \new_[100585]_  & \new_[100582]_ ;
  assign \new_[100587]_  = \new_[100586]_  & \new_[100579]_ ;
  assign \new_[100590]_  = ~A233 & A232;
  assign \new_[100593]_  = A235 & A234;
  assign \new_[100594]_  = \new_[100593]_  & \new_[100590]_ ;
  assign \new_[100597]_  = ~A299 & A298;
  assign \new_[100600]_  = A301 & A300;
  assign \new_[100601]_  = \new_[100600]_  & \new_[100597]_ ;
  assign \new_[100602]_  = \new_[100601]_  & \new_[100594]_ ;
  assign \new_[100605]_  = ~A168 & ~A169;
  assign \new_[100608]_  = A166 & A167;
  assign \new_[100609]_  = \new_[100608]_  & \new_[100605]_ ;
  assign \new_[100612]_  = ~A200 & A199;
  assign \new_[100615]_  = A203 & A201;
  assign \new_[100616]_  = \new_[100615]_  & \new_[100612]_ ;
  assign \new_[100617]_  = \new_[100616]_  & \new_[100609]_ ;
  assign \new_[100620]_  = ~A233 & A232;
  assign \new_[100623]_  = A235 & A234;
  assign \new_[100624]_  = \new_[100623]_  & \new_[100620]_ ;
  assign \new_[100627]_  = ~A299 & A298;
  assign \new_[100630]_  = A302 & A300;
  assign \new_[100631]_  = \new_[100630]_  & \new_[100627]_ ;
  assign \new_[100632]_  = \new_[100631]_  & \new_[100624]_ ;
  assign \new_[100635]_  = ~A168 & ~A169;
  assign \new_[100638]_  = A166 & A167;
  assign \new_[100639]_  = \new_[100638]_  & \new_[100635]_ ;
  assign \new_[100642]_  = ~A200 & A199;
  assign \new_[100645]_  = A203 & A201;
  assign \new_[100646]_  = \new_[100645]_  & \new_[100642]_ ;
  assign \new_[100647]_  = \new_[100646]_  & \new_[100639]_ ;
  assign \new_[100650]_  = ~A233 & A232;
  assign \new_[100653]_  = A235 & A234;
  assign \new_[100654]_  = \new_[100653]_  & \new_[100650]_ ;
  assign \new_[100657]_  = ~A266 & A265;
  assign \new_[100660]_  = A268 & A267;
  assign \new_[100661]_  = \new_[100660]_  & \new_[100657]_ ;
  assign \new_[100662]_  = \new_[100661]_  & \new_[100654]_ ;
  assign \new_[100665]_  = ~A168 & ~A169;
  assign \new_[100668]_  = A166 & A167;
  assign \new_[100669]_  = \new_[100668]_  & \new_[100665]_ ;
  assign \new_[100672]_  = ~A200 & A199;
  assign \new_[100675]_  = A203 & A201;
  assign \new_[100676]_  = \new_[100675]_  & \new_[100672]_ ;
  assign \new_[100677]_  = \new_[100676]_  & \new_[100669]_ ;
  assign \new_[100680]_  = ~A233 & A232;
  assign \new_[100683]_  = A235 & A234;
  assign \new_[100684]_  = \new_[100683]_  & \new_[100680]_ ;
  assign \new_[100687]_  = ~A266 & A265;
  assign \new_[100690]_  = A269 & A267;
  assign \new_[100691]_  = \new_[100690]_  & \new_[100687]_ ;
  assign \new_[100692]_  = \new_[100691]_  & \new_[100684]_ ;
  assign \new_[100695]_  = ~A168 & ~A169;
  assign \new_[100698]_  = A166 & A167;
  assign \new_[100699]_  = \new_[100698]_  & \new_[100695]_ ;
  assign \new_[100702]_  = ~A200 & A199;
  assign \new_[100705]_  = A203 & A201;
  assign \new_[100706]_  = \new_[100705]_  & \new_[100702]_ ;
  assign \new_[100707]_  = \new_[100706]_  & \new_[100699]_ ;
  assign \new_[100710]_  = ~A233 & A232;
  assign \new_[100713]_  = A236 & A234;
  assign \new_[100714]_  = \new_[100713]_  & \new_[100710]_ ;
  assign \new_[100717]_  = ~A299 & A298;
  assign \new_[100720]_  = A301 & A300;
  assign \new_[100721]_  = \new_[100720]_  & \new_[100717]_ ;
  assign \new_[100722]_  = \new_[100721]_  & \new_[100714]_ ;
  assign \new_[100725]_  = ~A168 & ~A169;
  assign \new_[100728]_  = A166 & A167;
  assign \new_[100729]_  = \new_[100728]_  & \new_[100725]_ ;
  assign \new_[100732]_  = ~A200 & A199;
  assign \new_[100735]_  = A203 & A201;
  assign \new_[100736]_  = \new_[100735]_  & \new_[100732]_ ;
  assign \new_[100737]_  = \new_[100736]_  & \new_[100729]_ ;
  assign \new_[100740]_  = ~A233 & A232;
  assign \new_[100743]_  = A236 & A234;
  assign \new_[100744]_  = \new_[100743]_  & \new_[100740]_ ;
  assign \new_[100747]_  = ~A299 & A298;
  assign \new_[100750]_  = A302 & A300;
  assign \new_[100751]_  = \new_[100750]_  & \new_[100747]_ ;
  assign \new_[100752]_  = \new_[100751]_  & \new_[100744]_ ;
  assign \new_[100755]_  = ~A168 & ~A169;
  assign \new_[100758]_  = A166 & A167;
  assign \new_[100759]_  = \new_[100758]_  & \new_[100755]_ ;
  assign \new_[100762]_  = ~A200 & A199;
  assign \new_[100765]_  = A203 & A201;
  assign \new_[100766]_  = \new_[100765]_  & \new_[100762]_ ;
  assign \new_[100767]_  = \new_[100766]_  & \new_[100759]_ ;
  assign \new_[100770]_  = ~A233 & A232;
  assign \new_[100773]_  = A236 & A234;
  assign \new_[100774]_  = \new_[100773]_  & \new_[100770]_ ;
  assign \new_[100777]_  = ~A266 & A265;
  assign \new_[100780]_  = A268 & A267;
  assign \new_[100781]_  = \new_[100780]_  & \new_[100777]_ ;
  assign \new_[100782]_  = \new_[100781]_  & \new_[100774]_ ;
  assign \new_[100785]_  = ~A168 & ~A169;
  assign \new_[100788]_  = A166 & A167;
  assign \new_[100789]_  = \new_[100788]_  & \new_[100785]_ ;
  assign \new_[100792]_  = ~A200 & A199;
  assign \new_[100795]_  = A203 & A201;
  assign \new_[100796]_  = \new_[100795]_  & \new_[100792]_ ;
  assign \new_[100797]_  = \new_[100796]_  & \new_[100789]_ ;
  assign \new_[100800]_  = ~A233 & A232;
  assign \new_[100803]_  = A236 & A234;
  assign \new_[100804]_  = \new_[100803]_  & \new_[100800]_ ;
  assign \new_[100807]_  = ~A266 & A265;
  assign \new_[100810]_  = A269 & A267;
  assign \new_[100811]_  = \new_[100810]_  & \new_[100807]_ ;
  assign \new_[100812]_  = \new_[100811]_  & \new_[100804]_ ;
  assign \new_[100815]_  = ~A168 & ~A169;
  assign \new_[100818]_  = A166 & A167;
  assign \new_[100819]_  = \new_[100818]_  & \new_[100815]_ ;
  assign \new_[100822]_  = ~A200 & A199;
  assign \new_[100825]_  = A203 & A201;
  assign \new_[100826]_  = \new_[100825]_  & \new_[100822]_ ;
  assign \new_[100827]_  = \new_[100826]_  & \new_[100819]_ ;
  assign \new_[100830]_  = ~A233 & ~A232;
  assign \new_[100833]_  = ~A268 & ~A266;
  assign \new_[100834]_  = \new_[100833]_  & \new_[100830]_ ;
  assign \new_[100837]_  = A298 & ~A269;
  assign \new_[100840]_  = ~A302 & ~A301;
  assign \new_[100841]_  = \new_[100840]_  & \new_[100837]_ ;
  assign \new_[100842]_  = \new_[100841]_  & \new_[100834]_ ;
  assign \new_[100845]_  = ~A169 & A170;
  assign \new_[100848]_  = ~A166 & A167;
  assign \new_[100849]_  = \new_[100848]_  & \new_[100845]_ ;
  assign \new_[100852]_  = ~A202 & ~A200;
  assign \new_[100855]_  = ~A233 & ~A203;
  assign \new_[100856]_  = \new_[100855]_  & \new_[100852]_ ;
  assign \new_[100857]_  = \new_[100856]_  & \new_[100849]_ ;
  assign \new_[100860]_  = ~A236 & ~A235;
  assign \new_[100863]_  = ~A268 & ~A266;
  assign \new_[100864]_  = \new_[100863]_  & \new_[100860]_ ;
  assign \new_[100867]_  = A298 & ~A269;
  assign \new_[100870]_  = ~A302 & ~A301;
  assign \new_[100871]_  = \new_[100870]_  & \new_[100867]_ ;
  assign \new_[100872]_  = \new_[100871]_  & \new_[100864]_ ;
  assign \new_[100875]_  = ~A169 & A170;
  assign \new_[100878]_  = A166 & ~A167;
  assign \new_[100879]_  = \new_[100878]_  & \new_[100875]_ ;
  assign \new_[100882]_  = ~A202 & ~A200;
  assign \new_[100885]_  = ~A233 & ~A203;
  assign \new_[100886]_  = \new_[100885]_  & \new_[100882]_ ;
  assign \new_[100887]_  = \new_[100886]_  & \new_[100879]_ ;
  assign \new_[100890]_  = ~A236 & ~A235;
  assign \new_[100893]_  = ~A268 & ~A266;
  assign \new_[100894]_  = \new_[100893]_  & \new_[100890]_ ;
  assign \new_[100897]_  = A298 & ~A269;
  assign \new_[100900]_  = ~A302 & ~A301;
  assign \new_[100901]_  = \new_[100900]_  & \new_[100897]_ ;
  assign \new_[100902]_  = \new_[100901]_  & \new_[100894]_ ;
  assign \new_[100905]_  = ~A169 & ~A170;
  assign \new_[100908]_  = A199 & ~A168;
  assign \new_[100909]_  = \new_[100908]_  & \new_[100905]_ ;
  assign \new_[100912]_  = A201 & ~A200;
  assign \new_[100915]_  = ~A233 & A202;
  assign \new_[100916]_  = \new_[100915]_  & \new_[100912]_ ;
  assign \new_[100917]_  = \new_[100916]_  & \new_[100909]_ ;
  assign \new_[100920]_  = ~A236 & ~A235;
  assign \new_[100923]_  = ~A268 & ~A266;
  assign \new_[100924]_  = \new_[100923]_  & \new_[100920]_ ;
  assign \new_[100927]_  = A298 & ~A269;
  assign \new_[100930]_  = ~A302 & ~A301;
  assign \new_[100931]_  = \new_[100930]_  & \new_[100927]_ ;
  assign \new_[100932]_  = \new_[100931]_  & \new_[100924]_ ;
  assign \new_[100935]_  = ~A169 & ~A170;
  assign \new_[100938]_  = A199 & ~A168;
  assign \new_[100939]_  = \new_[100938]_  & \new_[100935]_ ;
  assign \new_[100942]_  = A201 & ~A200;
  assign \new_[100945]_  = ~A233 & A203;
  assign \new_[100946]_  = \new_[100945]_  & \new_[100942]_ ;
  assign \new_[100947]_  = \new_[100946]_  & \new_[100939]_ ;
  assign \new_[100950]_  = ~A236 & ~A235;
  assign \new_[100953]_  = ~A268 & ~A266;
  assign \new_[100954]_  = \new_[100953]_  & \new_[100950]_ ;
  assign \new_[100957]_  = A298 & ~A269;
  assign \new_[100960]_  = ~A302 & ~A301;
  assign \new_[100961]_  = \new_[100960]_  & \new_[100957]_ ;
  assign \new_[100962]_  = \new_[100961]_  & \new_[100954]_ ;
  assign \new_[100965]_  = ~A168 & A169;
  assign \new_[100968]_  = ~A166 & A167;
  assign \new_[100969]_  = \new_[100968]_  & \new_[100965]_ ;
  assign \new_[100972]_  = ~A200 & A199;
  assign \new_[100975]_  = A202 & A201;
  assign \new_[100976]_  = \new_[100975]_  & \new_[100972]_ ;
  assign \new_[100977]_  = \new_[100976]_  & \new_[100969]_ ;
  assign \new_[100980]_  = ~A235 & ~A233;
  assign \new_[100983]_  = ~A266 & ~A236;
  assign \new_[100984]_  = \new_[100983]_  & \new_[100980]_ ;
  assign \new_[100987]_  = ~A269 & ~A268;
  assign \new_[100991]_  = ~A302 & ~A301;
  assign \new_[100992]_  = A298 & \new_[100991]_ ;
  assign \new_[100993]_  = \new_[100992]_  & \new_[100987]_ ;
  assign \new_[100994]_  = \new_[100993]_  & \new_[100984]_ ;
  assign \new_[100997]_  = ~A168 & A169;
  assign \new_[101000]_  = ~A166 & A167;
  assign \new_[101001]_  = \new_[101000]_  & \new_[100997]_ ;
  assign \new_[101004]_  = ~A200 & A199;
  assign \new_[101007]_  = A203 & A201;
  assign \new_[101008]_  = \new_[101007]_  & \new_[101004]_ ;
  assign \new_[101009]_  = \new_[101008]_  & \new_[101001]_ ;
  assign \new_[101012]_  = ~A235 & ~A233;
  assign \new_[101015]_  = ~A266 & ~A236;
  assign \new_[101016]_  = \new_[101015]_  & \new_[101012]_ ;
  assign \new_[101019]_  = ~A269 & ~A268;
  assign \new_[101023]_  = ~A302 & ~A301;
  assign \new_[101024]_  = A298 & \new_[101023]_ ;
  assign \new_[101025]_  = \new_[101024]_  & \new_[101019]_ ;
  assign \new_[101026]_  = \new_[101025]_  & \new_[101016]_ ;
  assign \new_[101029]_  = ~A168 & A169;
  assign \new_[101032]_  = A166 & ~A167;
  assign \new_[101033]_  = \new_[101032]_  & \new_[101029]_ ;
  assign \new_[101036]_  = ~A200 & A199;
  assign \new_[101039]_  = A202 & A201;
  assign \new_[101040]_  = \new_[101039]_  & \new_[101036]_ ;
  assign \new_[101041]_  = \new_[101040]_  & \new_[101033]_ ;
  assign \new_[101044]_  = ~A235 & ~A233;
  assign \new_[101047]_  = ~A266 & ~A236;
  assign \new_[101048]_  = \new_[101047]_  & \new_[101044]_ ;
  assign \new_[101051]_  = ~A269 & ~A268;
  assign \new_[101055]_  = ~A302 & ~A301;
  assign \new_[101056]_  = A298 & \new_[101055]_ ;
  assign \new_[101057]_  = \new_[101056]_  & \new_[101051]_ ;
  assign \new_[101058]_  = \new_[101057]_  & \new_[101048]_ ;
  assign \new_[101061]_  = ~A168 & A169;
  assign \new_[101064]_  = A166 & ~A167;
  assign \new_[101065]_  = \new_[101064]_  & \new_[101061]_ ;
  assign \new_[101068]_  = ~A200 & A199;
  assign \new_[101071]_  = A203 & A201;
  assign \new_[101072]_  = \new_[101071]_  & \new_[101068]_ ;
  assign \new_[101073]_  = \new_[101072]_  & \new_[101065]_ ;
  assign \new_[101076]_  = ~A235 & ~A233;
  assign \new_[101079]_  = ~A266 & ~A236;
  assign \new_[101080]_  = \new_[101079]_  & \new_[101076]_ ;
  assign \new_[101083]_  = ~A269 & ~A268;
  assign \new_[101087]_  = ~A302 & ~A301;
  assign \new_[101088]_  = A298 & \new_[101087]_ ;
  assign \new_[101089]_  = \new_[101088]_  & \new_[101083]_ ;
  assign \new_[101090]_  = \new_[101089]_  & \new_[101080]_ ;
  assign \new_[101093]_  = ~A168 & ~A169;
  assign \new_[101096]_  = A166 & A167;
  assign \new_[101097]_  = \new_[101096]_  & \new_[101093]_ ;
  assign \new_[101100]_  = ~A200 & A199;
  assign \new_[101103]_  = A202 & A201;
  assign \new_[101104]_  = \new_[101103]_  & \new_[101100]_ ;
  assign \new_[101105]_  = \new_[101104]_  & \new_[101097]_ ;
  assign \new_[101108]_  = ~A235 & ~A233;
  assign \new_[101111]_  = ~A266 & ~A236;
  assign \new_[101112]_  = \new_[101111]_  & \new_[101108]_ ;
  assign \new_[101115]_  = ~A269 & ~A268;
  assign \new_[101119]_  = ~A302 & ~A301;
  assign \new_[101120]_  = A298 & \new_[101119]_ ;
  assign \new_[101121]_  = \new_[101120]_  & \new_[101115]_ ;
  assign \new_[101122]_  = \new_[101121]_  & \new_[101112]_ ;
  assign \new_[101125]_  = ~A168 & ~A169;
  assign \new_[101128]_  = A166 & A167;
  assign \new_[101129]_  = \new_[101128]_  & \new_[101125]_ ;
  assign \new_[101132]_  = ~A200 & A199;
  assign \new_[101135]_  = A203 & A201;
  assign \new_[101136]_  = \new_[101135]_  & \new_[101132]_ ;
  assign \new_[101137]_  = \new_[101136]_  & \new_[101129]_ ;
  assign \new_[101140]_  = ~A235 & ~A233;
  assign \new_[101143]_  = ~A266 & ~A236;
  assign \new_[101144]_  = \new_[101143]_  & \new_[101140]_ ;
  assign \new_[101147]_  = ~A269 & ~A268;
  assign \new_[101151]_  = ~A302 & ~A301;
  assign \new_[101152]_  = A298 & \new_[101151]_ ;
  assign \new_[101153]_  = \new_[101152]_  & \new_[101147]_ ;
  assign \new_[101154]_  = \new_[101153]_  & \new_[101144]_ ;
endmodule


