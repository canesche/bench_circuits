module top ( clock, 
    p_10, p_12, p_11, pclk, p_9, p_8, p_7, p_6, p_5, p_4, p_3, p_2, p_1,
    p_40, p_45, p_46, p_47, p_48, p_41, p_42, p_43, p_44  );
  input  clock;
  input  p_10, p_12, p_11, pclk, p_9, p_8, p_7, p_6, p_5, p_4, p_3, p_2,
    p_1;
  output p_40, p_45, p_46, p_47, p_48, p_41, p_42, p_43, p_44;
  reg n_22, n_18, n_19, n_20, n_21, n_14, n_15, n_16, n_17, n_13, n_23,
    n_34, n_24, n_33, n_25, n_36, n_26, n_35, n_27, n_38, n_28, n_37, n_29,
    n_30, n_39, n_31, n_32;
  wire new_n104_, new_n105_, new_n106_1_, new_n107_, new_n108_, new_n109_,
    new_n110_, new_n111_1_, new_n112_, new_n113_, new_n114_, new_n115_,
    new_n116_1_, new_n117_, new_n118_, new_n119_, new_n120_, new_n121_1_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_1_, new_n127_,
    new_n128_, new_n129_, new_n130_, new_n131_1_, new_n132_, new_n133_,
    new_n134_, new_n135_, new_n136_1_, new_n137_, new_n138_, new_n139_,
    new_n140_, new_n141_1_, new_n142_, new_n143_, new_n144_, new_n145_,
    new_n146_1_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_1_,
    new_n152_, new_n153_, new_n154_, new_n155_, new_n156_1_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_1_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_1_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_1_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_1_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n474_, new_n475_, new_n477_, new_n478_, new_n480_, new_n481_,
    new_n483_, new_n484_, new_n486_, new_n487_, new_n489_, new_n490_,
    new_n492_, new_n493_, new_n495_, new_n496_, new_n498_, new_n499_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n507_,
    new_n508_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n516_, new_n517_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n525_, new_n526_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n534_, new_n535_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n543_, new_n544_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n552_, new_n553_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n567_, new_n568_,
    new_n570_, new_n571_, new_n573_, new_n574_, n46, n51, n56, n61, n66,
    n71, n76, n81, n86, n91, n96, n101, n106, n111, n116, n121, n126, n131,
    n136, n141, n146, n151, n156, n161, n166, n171, n176;
  assign new_n104_ = ~p_3 & p_2;
  assign new_n105_ = ~p_1 & new_n104_;
  assign new_n106_1_ = ~p_4 & n_31;
  assign new_n107_ = p_4 & ~n_31;
  assign new_n108_ = ~new_n106_1_ & ~new_n107_;
  assign new_n109_ = p_4 & ~new_n108_;
  assign new_n110_ = ~p_5 & n_32;
  assign new_n111_1_ = p_5 & ~n_32;
  assign new_n112_ = ~new_n110_ & ~new_n111_1_;
  assign new_n113_ = new_n109_ & new_n112_;
  assign new_n114_ = p_5 & ~new_n112_;
  assign new_n115_ = ~new_n113_ & ~new_n114_;
  assign new_n116_1_ = ~p_6 & n_33;
  assign new_n117_ = p_6 & ~n_33;
  assign new_n118_ = ~new_n116_1_ & ~new_n117_;
  assign new_n119_ = ~new_n115_ & new_n118_;
  assign new_n120_ = p_6 & ~new_n118_;
  assign new_n121_1_ = ~new_n119_ & ~new_n120_;
  assign new_n122_ = ~p_7 & n_34;
  assign new_n123_ = p_7 & ~n_34;
  assign new_n124_ = ~new_n122_ & ~new_n123_;
  assign new_n125_ = ~new_n121_1_ & new_n124_;
  assign new_n126_1_ = p_7 & ~new_n124_;
  assign new_n127_ = ~new_n125_ & ~new_n126_1_;
  assign new_n128_ = ~p_8 & n_35;
  assign new_n129_ = p_8 & ~n_35;
  assign new_n130_ = ~new_n128_ & ~new_n129_;
  assign new_n131_1_ = ~new_n127_ & new_n130_;
  assign new_n132_ = p_8 & ~new_n130_;
  assign new_n133_ = ~new_n131_1_ & ~new_n132_;
  assign new_n134_ = ~p_9 & n_36;
  assign new_n135_ = p_9 & ~n_36;
  assign new_n136_1_ = ~new_n134_ & ~new_n135_;
  assign new_n137_ = ~new_n133_ & new_n136_1_;
  assign new_n138_ = p_9 & ~new_n136_1_;
  assign new_n139_ = ~new_n137_ & ~new_n138_;
  assign new_n140_ = ~p_10 & n_37;
  assign new_n141_1_ = p_10 & ~n_37;
  assign new_n142_ = ~new_n140_ & ~new_n141_1_;
  assign new_n143_ = ~new_n139_ & new_n142_;
  assign new_n144_ = p_10 & ~new_n142_;
  assign new_n145_ = ~new_n143_ & ~new_n144_;
  assign new_n146_1_ = ~p_11 & n_38;
  assign new_n147_ = p_11 & ~n_38;
  assign new_n148_ = ~new_n146_1_ & ~new_n147_;
  assign new_n149_ = ~new_n145_ & new_n148_;
  assign new_n150_ = p_11 & ~new_n148_;
  assign new_n151_1_ = ~new_n149_ & ~new_n150_;
  assign new_n152_ = ~p_12 & n_39;
  assign new_n153_ = p_12 & ~n_39;
  assign new_n154_ = ~new_n152_ & ~new_n153_;
  assign new_n155_ = ~new_n151_1_ & new_n154_;
  assign new_n156_1_ = p_12 & ~new_n154_;
  assign new_n157_ = ~new_n155_ & ~new_n156_1_;
  assign new_n158_ = new_n105_ & ~new_n157_;
  assign new_n159_ = n_32 & ~new_n158_;
  assign new_n160_ = p_5 & new_n158_;
  assign new_n161_1_ = ~new_n159_ & ~new_n160_;
  assign new_n162_ = new_n105_ & ~new_n161_1_;
  assign new_n163_ = ~p_4 & n_22;
  assign new_n164_ = p_4 & ~n_22;
  assign new_n165_ = ~new_n163_ & ~new_n164_;
  assign new_n166_1_ = p_4 & ~new_n165_;
  assign new_n167_ = ~p_5 & n_23;
  assign new_n168_ = p_5 & ~n_23;
  assign new_n169_ = ~new_n167_ & ~new_n168_;
  assign new_n170_ = new_n166_1_ & new_n169_;
  assign new_n171_1_ = p_5 & ~new_n169_;
  assign new_n172_ = ~new_n170_ & ~new_n171_1_;
  assign new_n173_ = ~p_6 & n_24;
  assign new_n174_ = p_6 & ~n_24;
  assign new_n175_ = ~new_n173_ & ~new_n174_;
  assign new_n176_1_ = ~new_n172_ & new_n175_;
  assign new_n177_ = p_6 & ~new_n175_;
  assign new_n178_ = ~new_n176_1_ & ~new_n177_;
  assign new_n179_ = ~p_7 & n_25;
  assign new_n180_ = p_7 & ~n_25;
  assign new_n181_ = ~new_n179_ & ~new_n180_;
  assign new_n182_ = ~new_n178_ & new_n181_;
  assign new_n183_ = p_7 & ~new_n181_;
  assign new_n184_ = ~new_n182_ & ~new_n183_;
  assign new_n185_ = ~p_8 & n_26;
  assign new_n186_ = p_8 & ~n_26;
  assign new_n187_ = ~new_n185_ & ~new_n186_;
  assign new_n188_ = ~new_n184_ & new_n187_;
  assign new_n189_ = p_8 & ~new_n187_;
  assign new_n190_ = ~new_n188_ & ~new_n189_;
  assign new_n191_ = ~p_9 & n_27;
  assign new_n192_ = p_9 & ~n_27;
  assign new_n193_ = ~new_n191_ & ~new_n192_;
  assign new_n194_ = ~new_n190_ & new_n193_;
  assign new_n195_ = p_9 & ~new_n193_;
  assign new_n196_ = ~new_n194_ & ~new_n195_;
  assign new_n197_ = ~p_10 & n_28;
  assign new_n198_ = p_10 & ~n_28;
  assign new_n199_ = ~new_n197_ & ~new_n198_;
  assign new_n200_ = ~new_n196_ & new_n199_;
  assign new_n201_ = p_10 & ~new_n199_;
  assign new_n202_ = ~new_n200_ & ~new_n201_;
  assign new_n203_ = ~p_11 & n_29;
  assign new_n204_ = p_11 & ~n_29;
  assign new_n205_ = ~new_n203_ & ~new_n204_;
  assign new_n206_ = ~new_n202_ & new_n205_;
  assign new_n207_ = p_11 & ~new_n205_;
  assign new_n208_ = ~new_n206_ & ~new_n207_;
  assign new_n209_ = ~p_12 & n_30;
  assign new_n210_ = p_12 & ~n_30;
  assign new_n211_ = ~new_n209_ & ~new_n210_;
  assign new_n212_ = ~new_n208_ & new_n211_;
  assign new_n213_ = p_12 & ~new_n211_;
  assign new_n214_ = ~new_n212_ & ~new_n213_;
  assign new_n215_ = new_n105_ & ~new_n214_;
  assign new_n216_ = n_23 & new_n215_;
  assign new_n217_ = p_5 & ~new_n215_;
  assign new_n218_ = ~new_n216_ & ~new_n217_;
  assign new_n219_ = new_n105_ & ~new_n218_;
  assign new_n220_ = n_22 & new_n215_;
  assign new_n221_ = p_4 & ~new_n215_;
  assign new_n222_ = ~new_n220_ & ~new_n221_;
  assign new_n223_ = new_n105_ & ~new_n222_;
  assign new_n224_ = n_31 & ~new_n158_;
  assign new_n225_ = p_4 & new_n158_;
  assign new_n226_ = ~new_n224_ & ~new_n225_;
  assign new_n227_ = new_n105_ & ~new_n226_;
  assign new_n228_ = new_n223_ & new_n227_;
  assign new_n229_ = new_n162_ & new_n219_;
  assign new_n230_ = new_n228_ & new_n229_;
  assign new_n231_ = ~new_n162_ & new_n219_;
  assign new_n232_ = ~new_n228_ & new_n231_;
  assign new_n233_ = new_n162_ & ~new_n219_;
  assign new_n234_ = ~new_n228_ & new_n233_;
  assign new_n235_ = ~new_n162_ & ~new_n219_;
  assign new_n236_ = new_n228_ & new_n235_;
  assign new_n237_ = ~new_n230_ & ~new_n232_;
  assign new_n238_ = ~new_n234_ & ~new_n236_;
  assign new_n239_ = new_n237_ & new_n238_;
  assign new_n240_ = ~p_3 & ~new_n239_;
  assign new_n241_ = p_4 & p_3;
  assign new_n242_ = ~new_n240_ & ~new_n241_;
  assign new_n243_ = p_2 & ~new_n242_;
  assign new_n244_ = ~p_2 & n_13;
  assign new_n245_ = ~new_n243_ & ~new_n244_;
  assign p_40 = ~p_1 & ~new_n245_;
  assign new_n247_ = n_37 & ~new_n158_;
  assign new_n248_ = p_10 & new_n158_;
  assign new_n249_ = ~new_n247_ & ~new_n248_;
  assign new_n250_ = new_n105_ & ~new_n249_;
  assign new_n251_ = n_28 & new_n215_;
  assign new_n252_ = p_10 & ~new_n215_;
  assign new_n253_ = ~new_n251_ & ~new_n252_;
  assign new_n254_ = new_n105_ & ~new_n253_;
  assign new_n255_ = n_27 & new_n215_;
  assign new_n256_ = p_9 & ~new_n215_;
  assign new_n257_ = ~new_n255_ & ~new_n256_;
  assign new_n258_ = new_n105_ & ~new_n257_;
  assign new_n259_ = n_36 & ~new_n158_;
  assign new_n260_ = p_9 & new_n158_;
  assign new_n261_ = ~new_n259_ & ~new_n260_;
  assign new_n262_ = new_n105_ & ~new_n261_;
  assign new_n263_ = new_n258_ & new_n262_;
  assign new_n264_ = n_26 & new_n215_;
  assign new_n265_ = p_8 & ~new_n215_;
  assign new_n266_ = ~new_n264_ & ~new_n265_;
  assign new_n267_ = new_n105_ & ~new_n266_;
  assign new_n268_ = n_35 & ~new_n158_;
  assign new_n269_ = p_8 & new_n158_;
  assign new_n270_ = ~new_n268_ & ~new_n269_;
  assign new_n271_ = new_n105_ & ~new_n270_;
  assign new_n272_ = new_n267_ & new_n271_;
  assign new_n273_ = n_25 & new_n215_;
  assign new_n274_ = p_7 & ~new_n215_;
  assign new_n275_ = ~new_n273_ & ~new_n274_;
  assign new_n276_ = new_n105_ & ~new_n275_;
  assign new_n277_ = n_34 & ~new_n158_;
  assign new_n278_ = p_7 & new_n158_;
  assign new_n279_ = ~new_n277_ & ~new_n278_;
  assign new_n280_ = new_n105_ & ~new_n279_;
  assign new_n281_ = new_n276_ & new_n280_;
  assign new_n282_ = n_24 & new_n215_;
  assign new_n283_ = p_6 & ~new_n215_;
  assign new_n284_ = ~new_n282_ & ~new_n283_;
  assign new_n285_ = new_n105_ & ~new_n284_;
  assign new_n286_ = n_33 & ~new_n158_;
  assign new_n287_ = p_6 & new_n158_;
  assign new_n288_ = ~new_n286_ & ~new_n287_;
  assign new_n289_ = new_n105_ & ~new_n288_;
  assign new_n290_ = new_n285_ & new_n289_;
  assign new_n291_ = new_n162_ & new_n228_;
  assign new_n292_ = new_n219_ & new_n228_;
  assign new_n293_ = ~new_n229_ & ~new_n291_;
  assign new_n294_ = ~new_n292_ & new_n293_;
  assign new_n295_ = new_n289_ & ~new_n294_;
  assign new_n296_ = new_n285_ & ~new_n294_;
  assign new_n297_ = ~new_n290_ & ~new_n295_;
  assign new_n298_ = ~new_n296_ & new_n297_;
  assign new_n299_ = new_n280_ & ~new_n298_;
  assign new_n300_ = new_n276_ & ~new_n298_;
  assign new_n301_ = ~new_n281_ & ~new_n299_;
  assign new_n302_ = ~new_n300_ & new_n301_;
  assign new_n303_ = new_n271_ & ~new_n302_;
  assign new_n304_ = new_n267_ & ~new_n302_;
  assign new_n305_ = ~new_n272_ & ~new_n303_;
  assign new_n306_ = ~new_n304_ & new_n305_;
  assign new_n307_ = new_n262_ & ~new_n306_;
  assign new_n308_ = new_n258_ & ~new_n306_;
  assign new_n309_ = ~new_n263_ & ~new_n307_;
  assign new_n310_ = ~new_n308_ & new_n309_;
  assign new_n311_ = new_n250_ & new_n254_;
  assign new_n312_ = ~new_n310_ & new_n311_;
  assign new_n313_ = ~new_n250_ & new_n254_;
  assign new_n314_ = new_n310_ & new_n313_;
  assign new_n315_ = new_n250_ & ~new_n254_;
  assign new_n316_ = new_n310_ & new_n315_;
  assign new_n317_ = ~new_n250_ & ~new_n254_;
  assign new_n318_ = ~new_n310_ & new_n317_;
  assign new_n319_ = ~new_n312_ & ~new_n314_;
  assign new_n320_ = ~new_n316_ & ~new_n318_;
  assign new_n321_ = new_n319_ & new_n320_;
  assign new_n322_ = ~p_3 & ~new_n321_;
  assign new_n323_ = p_9 & p_3;
  assign new_n324_ = ~new_n322_ & ~new_n323_;
  assign new_n325_ = p_2 & ~new_n324_;
  assign new_n326_ = ~p_2 & n_18;
  assign new_n327_ = ~new_n325_ & ~new_n326_;
  assign p_45 = ~p_1 & ~new_n327_;
  assign new_n329_ = n_38 & ~new_n158_;
  assign new_n330_ = p_11 & new_n158_;
  assign new_n331_ = ~new_n329_ & ~new_n330_;
  assign new_n332_ = new_n105_ & ~new_n331_;
  assign new_n333_ = n_29 & new_n215_;
  assign new_n334_ = p_11 & ~new_n215_;
  assign new_n335_ = ~new_n333_ & ~new_n334_;
  assign new_n336_ = new_n105_ & ~new_n335_;
  assign new_n337_ = new_n250_ & ~new_n310_;
  assign new_n338_ = new_n254_ & ~new_n310_;
  assign new_n339_ = ~new_n311_ & ~new_n337_;
  assign new_n340_ = ~new_n338_ & new_n339_;
  assign new_n341_ = new_n332_ & new_n336_;
  assign new_n342_ = ~new_n340_ & new_n341_;
  assign new_n343_ = ~new_n332_ & new_n336_;
  assign new_n344_ = new_n340_ & new_n343_;
  assign new_n345_ = new_n332_ & ~new_n336_;
  assign new_n346_ = new_n340_ & new_n345_;
  assign new_n347_ = ~new_n332_ & ~new_n336_;
  assign new_n348_ = ~new_n340_ & new_n347_;
  assign new_n349_ = ~new_n342_ & ~new_n344_;
  assign new_n350_ = ~new_n346_ & ~new_n348_;
  assign new_n351_ = new_n349_ & new_n350_;
  assign new_n352_ = ~p_3 & ~new_n351_;
  assign new_n353_ = p_10 & p_3;
  assign new_n354_ = ~new_n352_ & ~new_n353_;
  assign new_n355_ = p_2 & ~new_n354_;
  assign new_n356_ = ~p_2 & n_19;
  assign new_n357_ = ~new_n355_ & ~new_n356_;
  assign p_46 = ~p_1 & ~new_n357_;
  assign new_n359_ = n_39 & ~new_n158_;
  assign new_n360_ = p_12 & new_n158_;
  assign new_n361_ = ~new_n359_ & ~new_n360_;
  assign new_n362_ = new_n105_ & ~new_n361_;
  assign new_n363_ = n_30 & new_n215_;
  assign new_n364_ = p_12 & ~new_n215_;
  assign new_n365_ = ~new_n363_ & ~new_n364_;
  assign new_n366_ = new_n105_ & ~new_n365_;
  assign new_n367_ = new_n332_ & ~new_n340_;
  assign new_n368_ = new_n336_ & ~new_n340_;
  assign new_n369_ = ~new_n341_ & ~new_n367_;
  assign new_n370_ = ~new_n368_ & new_n369_;
  assign new_n371_ = new_n362_ & new_n366_;
  assign new_n372_ = ~new_n370_ & new_n371_;
  assign new_n373_ = ~new_n362_ & new_n366_;
  assign new_n374_ = new_n370_ & new_n373_;
  assign new_n375_ = new_n362_ & ~new_n366_;
  assign new_n376_ = new_n370_ & new_n375_;
  assign new_n377_ = ~new_n362_ & ~new_n366_;
  assign new_n378_ = ~new_n370_ & new_n377_;
  assign new_n379_ = ~new_n372_ & ~new_n374_;
  assign new_n380_ = ~new_n376_ & ~new_n378_;
  assign new_n381_ = new_n379_ & new_n380_;
  assign new_n382_ = ~p_3 & ~new_n381_;
  assign new_n383_ = p_11 & p_3;
  assign new_n384_ = ~new_n382_ & ~new_n383_;
  assign new_n385_ = p_2 & ~new_n384_;
  assign new_n386_ = ~p_2 & n_20;
  assign new_n387_ = ~new_n385_ & ~new_n386_;
  assign p_47 = ~p_1 & ~new_n387_;
  assign new_n389_ = new_n362_ & ~new_n370_;
  assign new_n390_ = new_n366_ & ~new_n370_;
  assign new_n391_ = ~new_n371_ & ~new_n389_;
  assign new_n392_ = ~new_n390_ & new_n391_;
  assign new_n393_ = ~p_3 & ~new_n392_;
  assign new_n394_ = p_12 & p_3;
  assign new_n395_ = ~new_n393_ & ~new_n394_;
  assign new_n396_ = p_2 & ~new_n395_;
  assign new_n397_ = ~p_2 & n_21;
  assign new_n398_ = ~new_n396_ & ~new_n397_;
  assign p_48 = ~p_1 & ~new_n398_;
  assign new_n400_ = new_n290_ & ~new_n294_;
  assign new_n401_ = new_n285_ & ~new_n289_;
  assign new_n402_ = new_n294_ & new_n401_;
  assign new_n403_ = ~new_n285_ & new_n289_;
  assign new_n404_ = new_n294_ & new_n403_;
  assign new_n405_ = ~new_n285_ & ~new_n289_;
  assign new_n406_ = ~new_n294_ & new_n405_;
  assign new_n407_ = ~new_n400_ & ~new_n402_;
  assign new_n408_ = ~new_n404_ & ~new_n406_;
  assign new_n409_ = new_n407_ & new_n408_;
  assign new_n410_ = ~p_3 & ~new_n409_;
  assign new_n411_ = p_5 & p_3;
  assign new_n412_ = ~new_n410_ & ~new_n411_;
  assign new_n413_ = p_2 & ~new_n412_;
  assign new_n414_ = ~p_2 & n_14;
  assign new_n415_ = ~new_n413_ & ~new_n414_;
  assign p_41 = ~p_1 & ~new_n415_;
  assign new_n417_ = new_n281_ & ~new_n298_;
  assign new_n418_ = new_n276_ & ~new_n280_;
  assign new_n419_ = new_n298_ & new_n418_;
  assign new_n420_ = ~new_n276_ & new_n280_;
  assign new_n421_ = new_n298_ & new_n420_;
  assign new_n422_ = ~new_n276_ & ~new_n280_;
  assign new_n423_ = ~new_n298_ & new_n422_;
  assign new_n424_ = ~new_n417_ & ~new_n419_;
  assign new_n425_ = ~new_n421_ & ~new_n423_;
  assign new_n426_ = new_n424_ & new_n425_;
  assign new_n427_ = ~p_3 & ~new_n426_;
  assign new_n428_ = p_6 & p_3;
  assign new_n429_ = ~new_n427_ & ~new_n428_;
  assign new_n430_ = p_2 & ~new_n429_;
  assign new_n431_ = ~p_2 & n_15;
  assign new_n432_ = ~new_n430_ & ~new_n431_;
  assign p_42 = ~p_1 & ~new_n432_;
  assign new_n434_ = new_n272_ & ~new_n302_;
  assign new_n435_ = new_n267_ & ~new_n271_;
  assign new_n436_ = new_n302_ & new_n435_;
  assign new_n437_ = ~new_n267_ & new_n271_;
  assign new_n438_ = new_n302_ & new_n437_;
  assign new_n439_ = ~new_n267_ & ~new_n271_;
  assign new_n440_ = ~new_n302_ & new_n439_;
  assign new_n441_ = ~new_n434_ & ~new_n436_;
  assign new_n442_ = ~new_n438_ & ~new_n440_;
  assign new_n443_ = new_n441_ & new_n442_;
  assign new_n444_ = ~p_3 & ~new_n443_;
  assign new_n445_ = p_7 & p_3;
  assign new_n446_ = ~new_n444_ & ~new_n445_;
  assign new_n447_ = p_2 & ~new_n446_;
  assign new_n448_ = ~p_2 & n_16;
  assign new_n449_ = ~new_n447_ & ~new_n448_;
  assign p_43 = ~p_1 & ~new_n449_;
  assign new_n451_ = new_n263_ & ~new_n306_;
  assign new_n452_ = new_n258_ & ~new_n262_;
  assign new_n453_ = new_n306_ & new_n452_;
  assign new_n454_ = ~new_n258_ & new_n262_;
  assign new_n455_ = new_n306_ & new_n454_;
  assign new_n456_ = ~new_n258_ & ~new_n262_;
  assign new_n457_ = ~new_n306_ & new_n456_;
  assign new_n458_ = ~new_n451_ & ~new_n453_;
  assign new_n459_ = ~new_n455_ & ~new_n457_;
  assign new_n460_ = new_n458_ & new_n459_;
  assign new_n461_ = ~p_3 & ~new_n460_;
  assign new_n462_ = p_8 & p_3;
  assign new_n463_ = ~new_n461_ & ~new_n462_;
  assign new_n464_ = p_2 & ~new_n463_;
  assign new_n465_ = ~p_2 & n_17;
  assign new_n466_ = ~new_n464_ & ~new_n465_;
  assign p_44 = ~p_1 & ~new_n466_;
  assign new_n468_ = ~p_3 & new_n223_;
  assign new_n469_ = ~p_3 & ~new_n468_;
  assign new_n470_ = p_2 & ~new_n469_;
  assign new_n471_ = p_2 & ~new_n470_;
  assign new_n472_ = ~p_1 & ~new_n471_;
  assign n46 = p_1 | new_n472_;
  assign new_n474_ = p_9 & p_2;
  assign new_n475_ = ~new_n326_ & ~new_n474_;
  assign n51 = ~p_1 & ~new_n475_;
  assign new_n477_ = p_10 & p_2;
  assign new_n478_ = ~new_n356_ & ~new_n477_;
  assign n56 = ~p_1 & ~new_n478_;
  assign new_n480_ = p_11 & p_2;
  assign new_n481_ = ~new_n386_ & ~new_n480_;
  assign n61 = ~p_1 & ~new_n481_;
  assign new_n483_ = p_12 & p_2;
  assign new_n484_ = ~new_n397_ & ~new_n483_;
  assign n66 = ~p_1 & ~new_n484_;
  assign new_n486_ = p_5 & p_2;
  assign new_n487_ = ~new_n414_ & ~new_n486_;
  assign n71 = ~p_1 & ~new_n487_;
  assign new_n489_ = p_6 & p_2;
  assign new_n490_ = ~new_n431_ & ~new_n489_;
  assign n76 = ~p_1 & ~new_n490_;
  assign new_n492_ = p_7 & p_2;
  assign new_n493_ = ~new_n448_ & ~new_n492_;
  assign n81 = ~p_1 & ~new_n493_;
  assign new_n495_ = p_8 & p_2;
  assign new_n496_ = ~new_n465_ & ~new_n495_;
  assign n86 = ~p_1 & ~new_n496_;
  assign new_n498_ = p_4 & p_2;
  assign new_n499_ = ~new_n244_ & ~new_n498_;
  assign n91 = ~p_1 & ~new_n499_;
  assign new_n501_ = ~p_3 & new_n219_;
  assign new_n502_ = ~p_3 & ~new_n501_;
  assign new_n503_ = p_2 & ~new_n502_;
  assign new_n504_ = p_2 & ~new_n503_;
  assign new_n505_ = ~p_1 & ~new_n504_;
  assign n96 = p_1 | new_n505_;
  assign new_n507_ = ~p_3 & new_n280_;
  assign new_n508_ = p_2 & new_n507_;
  assign n101 = ~p_1 & new_n508_;
  assign new_n510_ = ~p_3 & new_n285_;
  assign new_n511_ = ~p_3 & ~new_n510_;
  assign new_n512_ = p_2 & ~new_n511_;
  assign new_n513_ = p_2 & ~new_n512_;
  assign new_n514_ = ~p_1 & ~new_n513_;
  assign n106 = p_1 | new_n514_;
  assign new_n516_ = ~p_3 & new_n289_;
  assign new_n517_ = p_2 & new_n516_;
  assign n111 = ~p_1 & new_n517_;
  assign new_n519_ = ~p_3 & new_n276_;
  assign new_n520_ = ~p_3 & ~new_n519_;
  assign new_n521_ = p_2 & ~new_n520_;
  assign new_n522_ = p_2 & ~new_n521_;
  assign new_n523_ = ~p_1 & ~new_n522_;
  assign n116 = p_1 | new_n523_;
  assign new_n525_ = ~p_3 & new_n262_;
  assign new_n526_ = p_2 & new_n525_;
  assign n121 = ~p_1 & new_n526_;
  assign new_n528_ = ~p_3 & new_n267_;
  assign new_n529_ = ~p_3 & ~new_n528_;
  assign new_n530_ = p_2 & ~new_n529_;
  assign new_n531_ = p_2 & ~new_n530_;
  assign new_n532_ = ~p_1 & ~new_n531_;
  assign n126 = p_1 | new_n532_;
  assign new_n534_ = ~p_3 & new_n271_;
  assign new_n535_ = p_2 & new_n534_;
  assign n131 = ~p_1 & new_n535_;
  assign new_n537_ = ~p_3 & new_n258_;
  assign new_n538_ = ~p_3 & ~new_n537_;
  assign new_n539_ = p_2 & ~new_n538_;
  assign new_n540_ = p_2 & ~new_n539_;
  assign new_n541_ = ~p_1 & ~new_n540_;
  assign n136 = p_1 | new_n541_;
  assign new_n543_ = ~p_3 & new_n332_;
  assign new_n544_ = p_2 & new_n543_;
  assign n141 = ~p_1 & new_n544_;
  assign new_n546_ = ~p_3 & new_n254_;
  assign new_n547_ = ~p_3 & ~new_n546_;
  assign new_n548_ = p_2 & ~new_n547_;
  assign new_n549_ = p_2 & ~new_n548_;
  assign new_n550_ = ~p_1 & ~new_n549_;
  assign n146 = p_1 | new_n550_;
  assign new_n552_ = ~p_3 & new_n250_;
  assign new_n553_ = p_2 & new_n552_;
  assign n151 = ~p_1 & new_n553_;
  assign new_n555_ = ~p_3 & new_n336_;
  assign new_n556_ = ~p_3 & ~new_n555_;
  assign new_n557_ = p_2 & ~new_n556_;
  assign new_n558_ = p_2 & ~new_n557_;
  assign new_n559_ = ~p_1 & ~new_n558_;
  assign n156 = p_1 | new_n559_;
  assign new_n561_ = ~p_3 & new_n366_;
  assign new_n562_ = ~p_3 & ~new_n561_;
  assign new_n563_ = p_2 & ~new_n562_;
  assign new_n564_ = p_2 & ~new_n563_;
  assign new_n565_ = ~p_1 & ~new_n564_;
  assign n161 = p_1 | new_n565_;
  assign new_n567_ = ~p_3 & new_n362_;
  assign new_n568_ = p_2 & new_n567_;
  assign n166 = ~p_1 & new_n568_;
  assign new_n570_ = ~p_3 & new_n227_;
  assign new_n571_ = p_2 & new_n570_;
  assign n171 = ~p_1 & new_n571_;
  assign new_n573_ = ~p_3 & new_n162_;
  assign new_n574_ = p_2 & new_n573_;
  assign n176 = ~p_1 & new_n574_;
  always @ (posedge clock) begin
    n_22 <= n46;
    n_18 <= n51;
    n_19 <= n56;
    n_20 <= n61;
    n_21 <= n66;
    n_14 <= n71;
    n_15 <= n76;
    n_16 <= n81;
    n_17 <= n86;
    n_13 <= n91;
    n_23 <= n96;
    n_34 <= n101;
    n_24 <= n106;
    n_33 <= n111;
    n_25 <= n116;
    n_36 <= n121;
    n_26 <= n126;
    n_35 <= n131;
    n_27 <= n136;
    n_38 <= n141;
    n_28 <= n146;
    n_37 <= n151;
    n_29 <= n156;
    n_30 <= n161;
    n_39 <= n166;
    n_31 <= n171;
    n_32 <= n176;
  end
endmodule

