// Benchmark "des_area" written by ABC on Thu Oct  8 22:03:23 2020

module des_area ( clock, 
    \desIn[0] , \desIn[1] , \desIn[2] , \desIn[3] , \desIn[4] , \desIn[5] ,
    \desIn[6] , \desIn[7] , \desIn[8] , \desIn[9] , \desIn[10] ,
    \desIn[11] , \desIn[12] , \desIn[13] , \desIn[14] , \desIn[15] ,
    \desIn[16] , \desIn[17] , \desIn[18] , \desIn[19] , \desIn[20] ,
    \desIn[21] , \desIn[22] , \desIn[23] , \desIn[24] , \desIn[25] ,
    \desIn[26] , \desIn[27] , \desIn[28] , \desIn[29] , \desIn[30] ,
    \desIn[31] , \desIn[32] , \desIn[33] , \desIn[34] , \desIn[35] ,
    \desIn[36] , \desIn[37] , \desIn[38] , \desIn[39] , \desIn[40] ,
    \desIn[41] , \desIn[42] , \desIn[43] , \desIn[44] , \desIn[45] ,
    \desIn[46] , \desIn[47] , \desIn[48] , \desIn[49] , \desIn[50] ,
    \desIn[51] , \desIn[52] , \desIn[53] , \desIn[54] , \desIn[55] ,
    \desIn[56] , \desIn[57] , \desIn[58] , \desIn[59] , \desIn[60] ,
    \desIn[61] , \desIn[62] , \desIn[63] , \key1[0] , \key1[1] , \key1[2] ,
    \key1[3] , \key1[4] , \key1[5] , \key1[6] , \key1[7] , \key1[8] ,
    \key1[9] , \key1[10] , \key1[11] , \key1[12] , \key1[13] , \key1[14] ,
    \key1[15] , \key1[16] , \key1[17] , \key1[18] , \key1[19] , \key1[20] ,
    \key1[21] , \key1[22] , \key1[23] , \key1[24] , \key1[25] , \key1[26] ,
    \key1[27] , \key1[28] , \key1[29] , \key1[30] , \key1[31] , \key1[32] ,
    \key1[33] , \key1[34] , \key1[35] , \key1[36] , \key1[37] , \key1[38] ,
    \key1[39] , \key1[40] , \key1[41] , \key1[42] , \key1[43] , \key1[44] ,
    \key1[45] , \key1[46] , \key1[47] , \key1[48] , \key1[49] , \key1[50] ,
    \key1[51] , \key1[52] , \key1[53] , \key1[54] , \key1[55] , \key2[0] ,
    \key2[1] , \key2[2] , \key2[3] , \key2[4] , \key2[5] , \key2[6] ,
    \key2[7] , \key2[8] , \key2[9] , \key2[10] , \key2[11] , \key2[12] ,
    \key2[13] , \key2[14] , \key2[15] , \key2[16] , \key2[17] , \key2[18] ,
    \key2[19] , \key2[20] , \key2[21] , \key2[22] , \key2[23] , \key2[24] ,
    \key2[25] , \key2[26] , \key2[27] , \key2[28] , \key2[29] , \key2[30] ,
    \key2[31] , \key2[32] , \key2[33] , \key2[34] , \key2[35] , \key2[36] ,
    \key2[37] , \key2[38] , \key2[39] , \key2[40] , \key2[41] , \key2[42] ,
    \key2[43] , \key2[44] , \key2[45] , \key2[46] , \key2[47] , \key2[48] ,
    \key2[49] , \key2[50] , \key2[51] , \key2[52] , \key2[53] , \key2[54] ,
    \key2[55] , \key3[0] , \key3[1] , \key3[2] , \key3[3] , \key3[4] ,
    \key3[5] , \key3[6] , \key3[7] , \key3[8] , \key3[9] , \key3[10] ,
    \key3[11] , \key3[12] , \key3[13] , \key3[14] , \key3[15] , \key3[16] ,
    \key3[17] , \key3[18] , \key3[19] , \key3[20] , \key3[21] , \key3[22] ,
    \key3[23] , \key3[24] , \key3[25] , \key3[26] , \key3[27] , \key3[28] ,
    \key3[29] , \key3[30] , \key3[31] , \key3[32] , \key3[33] , \key3[34] ,
    \key3[35] , \key3[36] , \key3[37] , \key3[38] , \key3[39] , \key3[40] ,
    \key3[41] , \key3[42] , \key3[43] , \key3[44] , \key3[45] , \key3[46] ,
    \key3[47] , \key3[48] , \key3[49] , \key3[50] , \key3[51] , \key3[52] ,
    \key3[53] , \key3[54] , \key3[55] , decrypt, clk, \roundSel[0] ,
    \roundSel[1] , \roundSel[2] , \roundSel[3] , \roundSel[4] ,
    \roundSel[5] ,
    \desOut[0] , \desOut[1] , \desOut[2] , \desOut[3] , \desOut[4] ,
    \desOut[5] , \desOut[6] , \desOut[7] , \desOut[8] , \desOut[9] ,
    \desOut[10] , \desOut[11] , \desOut[12] , \desOut[13] , \desOut[14] ,
    \desOut[15] , \desOut[16] , \desOut[17] , \desOut[18] , \desOut[19] ,
    \desOut[20] , \desOut[21] , \desOut[22] , \desOut[23] , \desOut[24] ,
    \desOut[25] , \desOut[26] , \desOut[27] , \desOut[28] , \desOut[29] ,
    \desOut[30] , \desOut[31] , \desOut[32] , \desOut[33] , \desOut[34] ,
    \desOut[35] , \desOut[36] , \desOut[37] , \desOut[38] , \desOut[39] ,
    \desOut[40] , \desOut[41] , \desOut[42] , \desOut[43] , \desOut[44] ,
    \desOut[45] , \desOut[46] , \desOut[47] , \desOut[48] , \desOut[49] ,
    \desOut[50] , \desOut[51] , \desOut[52] , \desOut[53] , \desOut[54] ,
    \desOut[55] , \desOut[56] , \desOut[57] , \desOut[58] , \desOut[59] ,
    \desOut[60] , \desOut[61] , \desOut[62] , \desOut[63]   );
  input  clock;
  input  \desIn[0] , \desIn[1] , \desIn[2] , \desIn[3] , \desIn[4] ,
    \desIn[5] , \desIn[6] , \desIn[7] , \desIn[8] , \desIn[9] ,
    \desIn[10] , \desIn[11] , \desIn[12] , \desIn[13] , \desIn[14] ,
    \desIn[15] , \desIn[16] , \desIn[17] , \desIn[18] , \desIn[19] ,
    \desIn[20] , \desIn[21] , \desIn[22] , \desIn[23] , \desIn[24] ,
    \desIn[25] , \desIn[26] , \desIn[27] , \desIn[28] , \desIn[29] ,
    \desIn[30] , \desIn[31] , \desIn[32] , \desIn[33] , \desIn[34] ,
    \desIn[35] , \desIn[36] , \desIn[37] , \desIn[38] , \desIn[39] ,
    \desIn[40] , \desIn[41] , \desIn[42] , \desIn[43] , \desIn[44] ,
    \desIn[45] , \desIn[46] , \desIn[47] , \desIn[48] , \desIn[49] ,
    \desIn[50] , \desIn[51] , \desIn[52] , \desIn[53] , \desIn[54] ,
    \desIn[55] , \desIn[56] , \desIn[57] , \desIn[58] , \desIn[59] ,
    \desIn[60] , \desIn[61] , \desIn[62] , \desIn[63] , \key1[0] ,
    \key1[1] , \key1[2] , \key1[3] , \key1[4] , \key1[5] , \key1[6] ,
    \key1[7] , \key1[8] , \key1[9] , \key1[10] , \key1[11] , \key1[12] ,
    \key1[13] , \key1[14] , \key1[15] , \key1[16] , \key1[17] , \key1[18] ,
    \key1[19] , \key1[20] , \key1[21] , \key1[22] , \key1[23] , \key1[24] ,
    \key1[25] , \key1[26] , \key1[27] , \key1[28] , \key1[29] , \key1[30] ,
    \key1[31] , \key1[32] , \key1[33] , \key1[34] , \key1[35] , \key1[36] ,
    \key1[37] , \key1[38] , \key1[39] , \key1[40] , \key1[41] , \key1[42] ,
    \key1[43] , \key1[44] , \key1[45] , \key1[46] , \key1[47] , \key1[48] ,
    \key1[49] , \key1[50] , \key1[51] , \key1[52] , \key1[53] , \key1[54] ,
    \key1[55] , \key2[0] , \key2[1] , \key2[2] , \key2[3] , \key2[4] ,
    \key2[5] , \key2[6] , \key2[7] , \key2[8] , \key2[9] , \key2[10] ,
    \key2[11] , \key2[12] , \key2[13] , \key2[14] , \key2[15] , \key2[16] ,
    \key2[17] , \key2[18] , \key2[19] , \key2[20] , \key2[21] , \key2[22] ,
    \key2[23] , \key2[24] , \key2[25] , \key2[26] , \key2[27] , \key2[28] ,
    \key2[29] , \key2[30] , \key2[31] , \key2[32] , \key2[33] , \key2[34] ,
    \key2[35] , \key2[36] , \key2[37] , \key2[38] , \key2[39] , \key2[40] ,
    \key2[41] , \key2[42] , \key2[43] , \key2[44] , \key2[45] , \key2[46] ,
    \key2[47] , \key2[48] , \key2[49] , \key2[50] , \key2[51] , \key2[52] ,
    \key2[53] , \key2[54] , \key2[55] , \key3[0] , \key3[1] , \key3[2] ,
    \key3[3] , \key3[4] , \key3[5] , \key3[6] , \key3[7] , \key3[8] ,
    \key3[9] , \key3[10] , \key3[11] , \key3[12] , \key3[13] , \key3[14] ,
    \key3[15] , \key3[16] , \key3[17] , \key3[18] , \key3[19] , \key3[20] ,
    \key3[21] , \key3[22] , \key3[23] , \key3[24] , \key3[25] , \key3[26] ,
    \key3[27] , \key3[28] , \key3[29] , \key3[30] , \key3[31] , \key3[32] ,
    \key3[33] , \key3[34] , \key3[35] , \key3[36] , \key3[37] , \key3[38] ,
    \key3[39] , \key3[40] , \key3[41] , \key3[42] , \key3[43] , \key3[44] ,
    \key3[45] , \key3[46] , \key3[47] , \key3[48] , \key3[49] , \key3[50] ,
    \key3[51] , \key3[52] , \key3[53] , \key3[54] , \key3[55] , decrypt,
    clk, \roundSel[0] , \roundSel[1] , \roundSel[2] , \roundSel[3] ,
    \roundSel[4] , \roundSel[5] ;
  output \desOut[0] , \desOut[1] , \desOut[2] , \desOut[3] , \desOut[4] ,
    \desOut[5] , \desOut[6] , \desOut[7] , \desOut[8] , \desOut[9] ,
    \desOut[10] , \desOut[11] , \desOut[12] , \desOut[13] , \desOut[14] ,
    \desOut[15] , \desOut[16] , \desOut[17] , \desOut[18] , \desOut[19] ,
    \desOut[20] , \desOut[21] , \desOut[22] , \desOut[23] , \desOut[24] ,
    \desOut[25] , \desOut[26] , \desOut[27] , \desOut[28] , \desOut[29] ,
    \desOut[30] , \desOut[31] , \desOut[32] , \desOut[33] , \desOut[34] ,
    \desOut[35] , \desOut[36] , \desOut[37] , \desOut[38] , \desOut[39] ,
    \desOut[40] , \desOut[41] , \desOut[42] , \desOut[43] , \desOut[44] ,
    \desOut[45] , \desOut[46] , \desOut[47] , \desOut[48] , \desOut[49] ,
    \desOut[50] , \desOut[51] , \desOut[52] , \desOut[53] , \desOut[54] ,
    \desOut[55] , \desOut[56] , \desOut[57] , \desOut[58] , \desOut[59] ,
    \desOut[60] , \desOut[61] , \desOut[62] , \desOut[63] ;
  reg \\FP_R_reg[25] , \\R_reg[25] , \\FP_R_reg[11] , \\R_reg[11] ,
    \\FP_R_reg[3] , \\R_reg[7] , \\FP_R_reg[7] , \\R_reg[3] ,
    \\FP_R_reg[15] , \\R_reg[15] , \\FP_R_reg[4] , \\R_reg[4] ,
    \\FP_R_reg[29] , \\R_reg[29] , \\FP_R_reg[22] , \\R_reg[22] ,
    \\R_reg[14] , \\R_reg[2] , \\FP_R_reg[5] , \\R_reg[5] ,
    \\FP_R_reg[28] , \\FP_R_reg[14] , \\FP_R_reg[2] , \\R_reg[13] ,
    \\R_reg[28] , \\FP_R_reg[13] , \\FP_R_reg[31] , \\R_reg[26] ,
    \\FP_R_reg[8] , \\FP_R_reg[20] , \\R_reg[31] , \\R_reg[20] ,
    \\R_reg[8] , \\FP_R_reg[12] , \\R_reg[12] , \\FP_R_reg[26] ,
    \\FP_R_reg[27] , \\FP_R_reg[19] , \\FP_R_reg[10] , \\FP_R_reg[21] ,
    \\FP_R_reg[6] , \\R_reg[10] , \\R_reg[19] , \\R_reg[21] , \\R_reg[27] ,
    \\R_reg[6] , \\FP_R_reg[9] , \\R_reg[9] , \\FP_R_reg[18] ,
    \\R_reg[18] , \\FP_R_reg[30] , \\FP_R_reg[32] , \\R_reg[32] ,
    \\FP_R_reg[23] , \\R_reg[23] , \\FP_R_reg[1] , \\R_reg[1] ,
    \\R_reg[30] , \\FP_R_reg[17] , \\R_reg[17] , \\FP_R_reg[24] ,
    \\R_reg[24] , \\FP_R_reg[16] , \\R_reg[16] , \\L_reg[15] ,
    \\L_reg[23] , \\L_reg[30] , \\L_reg[19] , \\L_reg[11] , \\L_reg[27] ,
    \\L_reg[28] , \\L_reg[17] , \\L_reg[3] , \\L_reg[24] , \\L_reg[31] ,
    \\FP_R_reg[49] , \\FP_R_reg[35] , \\FP_R_reg[56] , \\FP_R_reg[55] ,
    \\FP_R_reg[62] , \\FP_R_reg[47] , \\FP_R_reg[60] , \\FP_R_reg[59] ,
    \\FP_R_reg[43] , \\FP_R_reg[51] , \\FP_R_reg[63] , \\FP_R_reg[64] ,
    \\L_reg[8] , \\L_reg[26] , \\L_reg[32] , \\L_reg[25] , \\L_reg[13] ,
    \\L_reg[6] , \\L_reg[5] , \\L_reg[21] , \\L_reg[16] , \\L_reg[22] ,
    \\L_reg[1] , \\L_reg[7] , \\FP_R_reg[58] , \\FP_R_reg[54] ,
    \\FP_R_reg[53] , \\FP_R_reg[40] , \\FP_R_reg[38] , \\FP_R_reg[37] ,
    \\FP_R_reg[45] , \\FP_R_reg[57] , \\FP_R_reg[48] , \\FP_R_reg[33] ,
    \\FP_R_reg[39] , \\L_reg[12] , \\FP_R_reg[52] , \\FP_R_reg[36] ,
    \\FP_R_reg[42] , \\FP_R_reg[34] , \\L_reg[10] , \\L_reg[20] ,
    \\L_reg[14] , \\L_reg[18] , \\FP_R_reg[50] , \\L_reg[2] ,
    \\FP_R_reg[44] , \\L_reg[4] , \\FP_R_reg[46] , \\FP_R_reg[61] ,
    \\FP_R_reg[41] , \\L_reg[29] , \\L_reg[9] ;
  wire \new_[434]_ , \new_[435]_ , \new_[436]_ , \new_[437]_ , \new_[438]_ ,
    \new_[439]_ , \new_[440]_ , \new_[441]_ , \new_[442]_ , \new_[443]_ ,
    \new_[444]_ , \new_[445]_ , \new_[446]_ , \new_[447]_ , \new_[448]_ ,
    \new_[449]_ , \new_[450]_ , \new_[451]_ , \new_[452]_ , \new_[453]_ ,
    \new_[454]_ , \new_[455]_ , \new_[456]_ , \new_[457]_ , \new_[458]_ ,
    \new_[459]_ , \new_[463]_ , \new_[464]_ , \new_[465]_ , \new_[466]_ ,
    \new_[467]_ , \new_[468]_ , \new_[469]_ , \new_[470]_ , \new_[471]_ ,
    \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ , \new_[476]_ ,
    \new_[477]_ , \new_[478]_ , \new_[479]_ , \new_[480]_ , \new_[481]_ ,
    \new_[482]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ , \new_[486]_ ,
    \new_[489]_ , \new_[490]_ , \new_[491]_ , \new_[492]_ , \new_[493]_ ,
    \new_[494]_ , \new_[495]_ , \new_[496]_ , \new_[497]_ , \new_[499]_ ,
    \new_[500]_ , \new_[501]_ , \new_[502]_ , \new_[503]_ , \new_[504]_ ,
    \new_[505]_ , \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ ,
    \new_[510]_ , \new_[511]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ ,
    \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ ,
    \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ ,
    \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ ,
    \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ ,
    \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ ,
    \new_[686]_ , \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ ,
    \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ ,
    \new_[696]_ , \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ ,
    \new_[701]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ ,
    \new_[706]_ , \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ ,
    \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ ,
    \new_[716]_ , \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[726]_ , \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ ,
    \new_[731]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ ,
    \new_[741]_ , \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[746]_ , \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ ,
    \new_[751]_ , \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ ,
    \new_[756]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ ,
    \new_[766]_ , \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ ,
    \new_[771]_ , \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ ,
    \new_[776]_ , \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ ,
    \new_[781]_ , \new_[782]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ ,
    \new_[786]_ , \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ ,
    \new_[791]_ , \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ ,
    \new_[796]_ , \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ ,
    \new_[801]_ , \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ ,
    \new_[806]_ , \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ ,
    \new_[811]_ , \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ ,
    \new_[816]_ , \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[824]_ , \new_[825]_ ,
    \new_[826]_ , \new_[827]_ , \new_[828]_ , \new_[829]_ , \new_[830]_ ,
    \new_[831]_ , \new_[832]_ , \new_[833]_ , \new_[834]_ , \new_[835]_ ,
    \new_[836]_ , \new_[837]_ , \new_[838]_ , \new_[839]_ , \new_[840]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[845]_ ,
    \new_[846]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ , \new_[850]_ ,
    \new_[851]_ , \new_[852]_ , \new_[853]_ , \new_[854]_ , \new_[855]_ ,
    \new_[856]_ , \new_[857]_ , \new_[858]_ , \new_[859]_ , \new_[860]_ ,
    \new_[861]_ , \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ ,
    \new_[866]_ , \new_[867]_ , \new_[868]_ , \new_[869]_ , \new_[870]_ ,
    \new_[871]_ , \new_[872]_ , \new_[873]_ , \new_[874]_ , \new_[875]_ ,
    \new_[876]_ , \new_[877]_ , \new_[878]_ , \new_[879]_ , \new_[880]_ ,
    \new_[881]_ , \new_[882]_ , \new_[883]_ , \new_[884]_ , \new_[885]_ ,
    \new_[886]_ , \new_[887]_ , \new_[888]_ , \new_[889]_ , \new_[890]_ ,
    \new_[891]_ , \new_[892]_ , \new_[893]_ , \new_[894]_ , \new_[895]_ ,
    \new_[896]_ , \new_[897]_ , \new_[898]_ , \new_[899]_ , \new_[900]_ ,
    \new_[901]_ , \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ ,
    \new_[906]_ , \new_[907]_ , \new_[908]_ , \new_[909]_ , \new_[910]_ ,
    \new_[911]_ , \new_[912]_ , \new_[913]_ , \new_[914]_ , \new_[915]_ ,
    \new_[916]_ , \new_[917]_ , \new_[918]_ , \new_[919]_ , \new_[920]_ ,
    \new_[921]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[925]_ ,
    \new_[926]_ , \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ ,
    \new_[931]_ , \new_[932]_ , \new_[933]_ , \new_[934]_ , \new_[935]_ ,
    \new_[936]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ , \new_[940]_ ,
    \new_[941]_ , \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ ,
    \new_[946]_ , \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ ,
    \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ ,
    \new_[956]_ , \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ ,
    \new_[961]_ , \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ ,
    \new_[966]_ , \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ ,
    \new_[971]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ ,
    \new_[976]_ , \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ ,
    \new_[986]_ , \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ ,
    \new_[996]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1002]_ , \new_[1003]_ , \new_[1004]_ ,
    \new_[1005]_ , \new_[1006]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1009]_ , \new_[1010]_ , \new_[1011]_ , \new_[1012]_ ,
    \new_[1013]_ , \new_[1014]_ , \new_[1015]_ , \new_[1016]_ ,
    \new_[1017]_ , \new_[1018]_ , \new_[1019]_ , \new_[1020]_ ,
    \new_[1021]_ , \new_[1022]_ , \new_[1023]_ , \new_[1024]_ ,
    \new_[1025]_ , \new_[1026]_ , \new_[1027]_ , \new_[1028]_ ,
    \new_[1029]_ , \new_[1030]_ , \new_[1031]_ , \new_[1032]_ ,
    \new_[1033]_ , \new_[1034]_ , \new_[1035]_ , \new_[1036]_ ,
    \new_[1037]_ , \new_[1038]_ , \new_[1039]_ , \new_[1040]_ ,
    \new_[1041]_ , \new_[1042]_ , \new_[1043]_ , \new_[1044]_ ,
    \new_[1045]_ , \new_[1046]_ , \new_[1047]_ , \new_[1048]_ ,
    \new_[1049]_ , \new_[1050]_ , \new_[1051]_ , \new_[1052]_ ,
    \new_[1053]_ , \new_[1054]_ , \new_[1055]_ , \new_[1056]_ ,
    \new_[1057]_ , \new_[1058]_ , \new_[1059]_ , \new_[1060]_ ,
    \new_[1061]_ , \new_[1062]_ , \new_[1063]_ , \new_[1064]_ ,
    \new_[1065]_ , \new_[1066]_ , \new_[1067]_ , \new_[1068]_ ,
    \new_[1069]_ , \new_[1070]_ , \new_[1071]_ , \new_[1072]_ ,
    \new_[1073]_ , \new_[1074]_ , \new_[1075]_ , \new_[1076]_ ,
    \new_[1077]_ , \new_[1078]_ , \new_[1079]_ , \new_[1080]_ ,
    \new_[1081]_ , \new_[1082]_ , \new_[1083]_ , \new_[1084]_ ,
    \new_[1085]_ , \new_[1086]_ , \new_[1087]_ , \new_[1088]_ ,
    \new_[1089]_ , \new_[1090]_ , \new_[1091]_ , \new_[1092]_ ,
    \new_[1093]_ , \new_[1094]_ , \new_[1095]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1098]_ , \new_[1099]_ , \new_[1100]_ ,
    \new_[1101]_ , \new_[1102]_ , \new_[1103]_ , \new_[1104]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1107]_ , \new_[1108]_ ,
    \new_[1109]_ , \new_[1110]_ , \new_[1111]_ , \new_[1112]_ ,
    \new_[1113]_ , \new_[1114]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1118]_ , \new_[1119]_ , \new_[1120]_ ,
    \new_[1121]_ , \new_[1122]_ , \new_[1123]_ , \new_[1124]_ ,
    \new_[1125]_ , \new_[1126]_ , \new_[1127]_ , \new_[1128]_ ,
    \new_[1129]_ , \new_[1130]_ , \new_[1131]_ , \new_[1132]_ ,
    \new_[1133]_ , \new_[1134]_ , \new_[1135]_ , \new_[1136]_ ,
    \new_[1137]_ , \new_[1138]_ , \new_[1139]_ , \new_[1140]_ ,
    \new_[1141]_ , \new_[1142]_ , \new_[1143]_ , \new_[1144]_ ,
    \new_[1145]_ , \new_[1146]_ , \new_[1147]_ , \new_[1148]_ ,
    \new_[1149]_ , \new_[1150]_ , \new_[1151]_ , \new_[1152]_ ,
    \new_[1153]_ , \new_[1154]_ , \new_[1155]_ , \new_[1156]_ ,
    \new_[1157]_ , \new_[1158]_ , \new_[1159]_ , \new_[1160]_ ,
    \new_[1161]_ , \new_[1162]_ , \new_[1163]_ , \new_[1164]_ ,
    \new_[1165]_ , \new_[1166]_ , \new_[1167]_ , \new_[1168]_ ,
    \new_[1169]_ , \new_[1170]_ , \new_[1171]_ , \new_[1172]_ ,
    \new_[1173]_ , \new_[1174]_ , \new_[1175]_ , \new_[1176]_ ,
    \new_[1177]_ , \new_[1178]_ , \new_[1179]_ , \new_[1180]_ ,
    \new_[1181]_ , \new_[1182]_ , \new_[1183]_ , \new_[1184]_ ,
    \new_[1185]_ , \new_[1186]_ , \new_[1187]_ , \new_[1188]_ ,
    \new_[1189]_ , \new_[1190]_ , \new_[1191]_ , \new_[1192]_ ,
    \new_[1193]_ , \new_[1194]_ , \new_[1195]_ , \new_[1196]_ ,
    \new_[1197]_ , \new_[1198]_ , \new_[1199]_ , \new_[1200]_ ,
    \new_[1201]_ , \new_[1202]_ , \new_[1203]_ , \new_[1204]_ ,
    \new_[1205]_ , \new_[1206]_ , \new_[1207]_ , \new_[1208]_ ,
    \new_[1209]_ , \new_[1210]_ , \new_[1211]_ , \new_[1212]_ ,
    \new_[1213]_ , \new_[1214]_ , \new_[1215]_ , \new_[1216]_ ,
    \new_[1217]_ , \new_[1218]_ , \new_[1219]_ , \new_[1220]_ ,
    \new_[1221]_ , \new_[1222]_ , \new_[1223]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1226]_ , \new_[1227]_ , \new_[1228]_ ,
    \new_[1229]_ , \new_[1230]_ , \new_[1231]_ , \new_[1232]_ ,
    \new_[1233]_ , \new_[1234]_ , \new_[1235]_ , \new_[1236]_ ,
    \new_[1237]_ , \new_[1238]_ , \new_[1239]_ , \new_[1240]_ ,
    \new_[1241]_ , \new_[1242]_ , \new_[1243]_ , \new_[1244]_ ,
    \new_[1245]_ , \new_[1246]_ , \new_[1247]_ , \new_[1248]_ ,
    \new_[1249]_ , \new_[1250]_ , \new_[1251]_ , \new_[1252]_ ,
    \new_[1253]_ , \new_[1254]_ , \new_[1255]_ , \new_[1256]_ ,
    \new_[1257]_ , \new_[1258]_ , \new_[1259]_ , \new_[1260]_ ,
    \new_[1261]_ , \new_[1262]_ , \new_[1263]_ , \new_[1264]_ ,
    \new_[1265]_ , \new_[1266]_ , \new_[1267]_ , \new_[1268]_ ,
    \new_[1269]_ , \new_[1270]_ , \new_[1271]_ , \new_[1272]_ ,
    \new_[1273]_ , \new_[1274]_ , \new_[1275]_ , \new_[1276]_ ,
    \new_[1277]_ , \new_[1278]_ , \new_[1279]_ , \new_[1280]_ ,
    \new_[1281]_ , \new_[1282]_ , \new_[1283]_ , \new_[1284]_ ,
    \new_[1285]_ , \new_[1286]_ , \new_[1287]_ , \new_[1288]_ ,
    \new_[1289]_ , \new_[1290]_ , \new_[1291]_ , \new_[1292]_ ,
    \new_[1293]_ , \new_[1294]_ , \new_[1295]_ , \new_[1296]_ ,
    \new_[1297]_ , \new_[1298]_ , \new_[1299]_ , \new_[1300]_ ,
    \new_[1301]_ , \new_[1302]_ , \new_[1303]_ , \new_[1304]_ ,
    \new_[1305]_ , \new_[1306]_ , \new_[1307]_ , \new_[1308]_ ,
    \new_[1309]_ , \new_[1310]_ , \new_[1311]_ , \new_[1312]_ ,
    \new_[1313]_ , \new_[1314]_ , \new_[1315]_ , \new_[1316]_ ,
    \new_[1317]_ , \new_[1318]_ , \new_[1319]_ , \new_[1320]_ ,
    \new_[1321]_ , \new_[1322]_ , \new_[1323]_ , \new_[1324]_ ,
    \new_[1325]_ , \new_[1326]_ , \new_[1327]_ , \new_[1328]_ ,
    \new_[1329]_ , \new_[1330]_ , \new_[1331]_ , \new_[1332]_ ,
    \new_[1333]_ , \new_[1334]_ , \new_[1335]_ , \new_[1336]_ ,
    \new_[1337]_ , \new_[1338]_ , \new_[1339]_ , \new_[1340]_ ,
    \new_[1341]_ , \new_[1342]_ , \new_[1343]_ , \new_[1344]_ ,
    \new_[1345]_ , \new_[1346]_ , \new_[1347]_ , \new_[1348]_ ,
    \new_[1349]_ , \new_[1350]_ , \new_[1351]_ , \new_[1352]_ ,
    \new_[1353]_ , \new_[1354]_ , \new_[1355]_ , \new_[1356]_ ,
    \new_[1357]_ , \new_[1358]_ , \new_[1359]_ , \new_[1360]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1363]_ , \new_[1364]_ ,
    \new_[1365]_ , \new_[1366]_ , \new_[1367]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1370]_ , \new_[1371]_ , \new_[1372]_ ,
    \new_[1373]_ , \new_[1374]_ , \new_[1375]_ , \new_[1376]_ ,
    \new_[1377]_ , \new_[1378]_ , \new_[1379]_ , \new_[1380]_ ,
    \new_[1381]_ , \new_[1382]_ , \new_[1383]_ , \new_[1384]_ ,
    \new_[1385]_ , \new_[1386]_ , \new_[1387]_ , \new_[1388]_ ,
    \new_[1389]_ , \new_[1390]_ , \new_[1391]_ , \new_[1392]_ ,
    \new_[1393]_ , \new_[1394]_ , \new_[1395]_ , \new_[1396]_ ,
    \new_[1397]_ , \new_[1398]_ , \new_[1399]_ , \new_[1400]_ ,
    \new_[1401]_ , \new_[1402]_ , \new_[1403]_ , \new_[1404]_ ,
    \new_[1405]_ , \new_[1406]_ , \new_[1407]_ , \new_[1408]_ ,
    \new_[1409]_ , \new_[1410]_ , \new_[1411]_ , \new_[1412]_ ,
    \new_[1413]_ , \new_[1414]_ , \new_[1415]_ , \new_[1416]_ ,
    \new_[1417]_ , \new_[1418]_ , \new_[1419]_ , \new_[1420]_ ,
    \new_[1421]_ , \new_[1422]_ , \new_[1423]_ , \new_[1424]_ ,
    \new_[1425]_ , \new_[1426]_ , \new_[1427]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1430]_ , \new_[1431]_ , \new_[1432]_ ,
    \new_[1433]_ , \new_[1434]_ , \new_[1435]_ , \new_[1436]_ ,
    \new_[1437]_ , \new_[1438]_ , \new_[1439]_ , \new_[1440]_ ,
    \new_[1441]_ , \new_[1442]_ , \new_[1443]_ , \new_[1444]_ ,
    \new_[1445]_ , \new_[1446]_ , \new_[1447]_ , \new_[1448]_ ,
    \new_[1449]_ , \new_[1450]_ , \new_[1451]_ , \new_[1452]_ ,
    \new_[1453]_ , \new_[1454]_ , \new_[1455]_ , \new_[1456]_ ,
    \new_[1457]_ , \new_[1458]_ , \new_[1459]_ , \new_[1460]_ ,
    \new_[1461]_ , \new_[1462]_ , \new_[1463]_ , \new_[1464]_ ,
    \new_[1465]_ , \new_[1466]_ , \new_[1467]_ , \new_[1468]_ ,
    \new_[1469]_ , \new_[1470]_ , \new_[1471]_ , \new_[1472]_ ,
    \new_[1473]_ , \new_[1474]_ , \new_[1475]_ , \new_[1476]_ ,
    \new_[1477]_ , \new_[1478]_ , \new_[1479]_ , \new_[1480]_ ,
    \new_[1481]_ , \new_[1482]_ , \new_[1483]_ , \new_[1484]_ ,
    \new_[1485]_ , \new_[1486]_ , \new_[1487]_ , \new_[1488]_ ,
    \new_[1489]_ , \new_[1490]_ , \new_[1491]_ , \new_[1492]_ ,
    \new_[1493]_ , \new_[1494]_ , \new_[1495]_ , \new_[1496]_ ,
    \new_[1497]_ , \new_[1498]_ , \new_[1499]_ , \new_[1500]_ ,
    \new_[1501]_ , \new_[1502]_ , \new_[1503]_ , \new_[1504]_ ,
    \new_[1505]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1514]_ , \new_[1515]_ , \new_[1516]_ ,
    \new_[1517]_ , \new_[1518]_ , \new_[1519]_ , \new_[1520]_ ,
    \new_[1521]_ , \new_[1522]_ , \new_[1523]_ , \new_[1524]_ ,
    \new_[1525]_ , \new_[1526]_ , \new_[1527]_ , \new_[1528]_ ,
    \new_[1529]_ , \new_[1530]_ , \new_[1531]_ , \new_[1532]_ ,
    \new_[1533]_ , \new_[1534]_ , \new_[1535]_ , \new_[1536]_ ,
    \new_[1537]_ , \new_[1538]_ , \new_[1539]_ , \new_[1540]_ ,
    \new_[1541]_ , \new_[1542]_ , \new_[1543]_ , \new_[1544]_ ,
    \new_[1545]_ , \new_[1546]_ , \new_[1547]_ , \new_[1548]_ ,
    \new_[1549]_ , \new_[1550]_ , \new_[1551]_ , \new_[1552]_ ,
    \new_[1553]_ , \new_[1554]_ , \new_[1555]_ , \new_[1556]_ ,
    \new_[1557]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1563]_ , \new_[1564]_ ,
    \new_[1565]_ , \new_[1566]_ , \new_[1567]_ , \new_[1568]_ ,
    \new_[1569]_ , \new_[1570]_ , \new_[1571]_ , \new_[1572]_ ,
    \new_[1573]_ , \new_[1574]_ , \new_[1575]_ , \new_[1576]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1579]_ , \new_[1580]_ ,
    \new_[1581]_ , \new_[1582]_ , \new_[1583]_ , \new_[1584]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1587]_ , \new_[1588]_ ,
    \new_[1589]_ , \new_[1590]_ , \new_[1591]_ , \new_[1592]_ ,
    \new_[1593]_ , \new_[1594]_ , \new_[1595]_ , \new_[1596]_ ,
    \new_[1597]_ , \new_[1598]_ , \new_[1599]_ , \new_[1600]_ ,
    \new_[1601]_ , \new_[1602]_ , \new_[1603]_ , \new_[1604]_ ,
    \new_[1605]_ , \new_[1606]_ , \new_[1607]_ , \new_[1608]_ ,
    \new_[1609]_ , \new_[1610]_ , \new_[1611]_ , \new_[1612]_ ,
    \new_[1613]_ , \new_[1614]_ , \new_[1615]_ , \new_[1616]_ ,
    \new_[1617]_ , \new_[1618]_ , \new_[1619]_ , \new_[1620]_ ,
    \new_[1621]_ , \new_[1622]_ , \new_[1623]_ , \new_[1624]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1627]_ , \new_[1628]_ ,
    \new_[1629]_ , \new_[1630]_ , \new_[1631]_ , \new_[1632]_ ,
    \new_[1633]_ , \new_[1634]_ , \new_[1635]_ , \new_[1636]_ ,
    \new_[1637]_ , \new_[1638]_ , \new_[1639]_ , \new_[1640]_ ,
    \new_[1641]_ , \new_[1642]_ , \new_[1643]_ , \new_[1644]_ ,
    \new_[1645]_ , \new_[1646]_ , \new_[1647]_ , \new_[1648]_ ,
    \new_[1649]_ , \new_[1650]_ , \new_[1651]_ , \new_[1652]_ ,
    \new_[1653]_ , \new_[1654]_ , \new_[1655]_ , \new_[1656]_ ,
    \new_[1657]_ , \new_[1658]_ , \new_[1659]_ , \new_[1660]_ ,
    \new_[1661]_ , \new_[1662]_ , \new_[1663]_ , \new_[1664]_ ,
    \new_[1665]_ , \new_[1666]_ , \new_[1667]_ , \new_[1668]_ ,
    \new_[1669]_ , \new_[1670]_ , \new_[1671]_ , \new_[1672]_ ,
    \new_[1673]_ , \new_[1674]_ , \new_[1675]_ , \new_[1676]_ ,
    \new_[1677]_ , \new_[1678]_ , \new_[1679]_ , \new_[1680]_ ,
    \new_[1681]_ , \new_[1682]_ , \new_[1683]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1686]_ , \new_[1687]_ , \new_[1688]_ ,
    \new_[1689]_ , \new_[1690]_ , \new_[1691]_ , \new_[1692]_ ,
    \new_[1693]_ , \new_[1694]_ , \new_[1695]_ , \new_[1696]_ ,
    \new_[1697]_ , \new_[1698]_ , \new_[1699]_ , \new_[1700]_ ,
    \new_[1701]_ , \new_[1702]_ , \new_[1703]_ , \new_[1704]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1707]_ , \new_[1708]_ ,
    \new_[1709]_ , \new_[1710]_ , \new_[1711]_ , \new_[1712]_ ,
    \new_[1713]_ , \new_[1714]_ , \new_[1715]_ , \new_[1716]_ ,
    \new_[1717]_ , \new_[1718]_ , \new_[1719]_ , \new_[1720]_ ,
    \new_[1721]_ , \new_[1722]_ , \new_[1723]_ , \new_[1724]_ ,
    \new_[1725]_ , \new_[1726]_ , \new_[1727]_ , \new_[1728]_ ,
    \new_[1729]_ , \new_[1730]_ , \new_[1731]_ , \new_[1732]_ ,
    \new_[1733]_ , \new_[1734]_ , \new_[1735]_ , \new_[1736]_ ,
    \new_[1737]_ , \new_[1738]_ , \new_[1739]_ , \new_[1740]_ ,
    \new_[1741]_ , \new_[1742]_ , \new_[1743]_ , \new_[1744]_ ,
    \new_[1745]_ , \new_[1746]_ , \new_[1747]_ , \new_[1748]_ ,
    \new_[1749]_ , \new_[1750]_ , \new_[1751]_ , \new_[1752]_ ,
    \new_[1753]_ , \new_[1754]_ , \new_[1755]_ , \new_[1756]_ ,
    \new_[1757]_ , \new_[1758]_ , \new_[1759]_ , \new_[1760]_ ,
    \new_[1761]_ , \new_[1762]_ , \new_[1763]_ , \new_[1764]_ ,
    \new_[1765]_ , \new_[1766]_ , \new_[1767]_ , \new_[1768]_ ,
    \new_[1769]_ , \new_[1770]_ , \new_[1771]_ , \new_[1772]_ ,
    \new_[1773]_ , \new_[1774]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1780]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1783]_ , \new_[1784]_ ,
    \new_[1785]_ , \new_[1786]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1792]_ ,
    \new_[1793]_ , \new_[1794]_ , \new_[1795]_ , \new_[1796]_ ,
    \new_[1797]_ , \new_[1798]_ , \new_[1799]_ , \new_[1800]_ ,
    \new_[1801]_ , \new_[1802]_ , \new_[1803]_ , \new_[1804]_ ,
    \new_[1805]_ , \new_[1806]_ , \new_[1807]_ , \new_[1808]_ ,
    \new_[1809]_ , \new_[1810]_ , \new_[1811]_ , \new_[1812]_ ,
    \new_[1813]_ , \new_[1814]_ , \new_[1815]_ , \new_[1816]_ ,
    \new_[1817]_ , \new_[1818]_ , \new_[1819]_ , \new_[1820]_ ,
    \new_[1821]_ , \new_[1822]_ , \new_[1823]_ , \new_[1824]_ ,
    \new_[1825]_ , \new_[1826]_ , \new_[1827]_ , \new_[1828]_ ,
    \new_[1829]_ , \new_[1830]_ , \new_[1831]_ , \new_[1832]_ ,
    \new_[1833]_ , \new_[1834]_ , \new_[1835]_ , \new_[1836]_ ,
    \new_[1837]_ , \new_[1838]_ , \new_[1839]_ , \new_[1840]_ ,
    \new_[1841]_ , \new_[1842]_ , \new_[1843]_ , \new_[1844]_ ,
    \new_[1845]_ , \new_[1846]_ , \new_[1847]_ , \new_[1848]_ ,
    \new_[1849]_ , \new_[1850]_ , \new_[1851]_ , \new_[1852]_ ,
    \new_[1853]_ , \new_[1854]_ , \new_[1855]_ , \new_[1856]_ ,
    \new_[1857]_ , \new_[1858]_ , \new_[1859]_ , \new_[1860]_ ,
    \new_[1861]_ , \new_[1862]_ , \new_[1863]_ , \new_[1864]_ ,
    \new_[1865]_ , \new_[1866]_ , \new_[1867]_ , \new_[1868]_ ,
    \new_[1869]_ , \new_[1870]_ , \new_[1871]_ , \new_[1872]_ ,
    \new_[1873]_ , \new_[1874]_ , \new_[1875]_ , \new_[1876]_ ,
    \new_[1877]_ , \new_[1878]_ , \new_[1879]_ , \new_[1880]_ ,
    \new_[1881]_ , \new_[1882]_ , \new_[1883]_ , \new_[1884]_ ,
    \new_[1885]_ , \new_[1886]_ , \new_[1887]_ , \new_[1888]_ ,
    \new_[1889]_ , \new_[1890]_ , \new_[1891]_ , \new_[1892]_ ,
    \new_[1893]_ , \new_[1894]_ , \new_[1895]_ , \new_[1896]_ ,
    \new_[1897]_ , \new_[1898]_ , \new_[1899]_ , \new_[1900]_ ,
    \new_[1901]_ , \new_[1902]_ , \new_[1903]_ , \new_[1904]_ ,
    \new_[1905]_ , \new_[1906]_ , \new_[1907]_ , \new_[1908]_ ,
    \new_[1909]_ , \new_[1910]_ , \new_[1911]_ , \new_[1912]_ ,
    \new_[1913]_ , \new_[1914]_ , \new_[1915]_ , \new_[1916]_ ,
    \new_[1917]_ , \new_[1918]_ , \new_[1919]_ , \new_[1920]_ ,
    \new_[1921]_ , \new_[1922]_ , \new_[1923]_ , \new_[1924]_ ,
    \new_[1925]_ , \new_[1926]_ , \new_[1927]_ , \new_[1928]_ ,
    \new_[1929]_ , \new_[1930]_ , \new_[1931]_ , \new_[1932]_ ,
    \new_[1933]_ , \new_[1934]_ , \new_[1935]_ , \new_[1936]_ ,
    \new_[1937]_ , \new_[1938]_ , \new_[1939]_ , \new_[1940]_ ,
    \new_[1941]_ , \new_[1942]_ , \new_[1943]_ , \new_[1944]_ ,
    \new_[1945]_ , \new_[1946]_ , \new_[1947]_ , \new_[1948]_ ,
    \new_[1949]_ , \new_[1950]_ , \new_[1951]_ , \new_[1952]_ ,
    \new_[1953]_ , \new_[1954]_ , \new_[1955]_ , \new_[1956]_ ,
    \new_[1957]_ , \new_[1958]_ , \new_[1959]_ , \new_[1960]_ ,
    \new_[1961]_ , \new_[1962]_ , \new_[1963]_ , \new_[1964]_ ,
    \new_[1965]_ , \new_[1966]_ , \new_[1967]_ , \new_[1968]_ ,
    \new_[1969]_ , \new_[1970]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1978]_ , \new_[1979]_ , \new_[1980]_ ,
    \new_[1981]_ , \new_[1982]_ , \new_[1983]_ , \new_[1984]_ ,
    \new_[1985]_ , \new_[1986]_ , \new_[1987]_ , \new_[1988]_ ,
    \new_[1989]_ , \new_[1990]_ , \new_[1991]_ , \new_[1992]_ ,
    \new_[1993]_ , \new_[1994]_ , \new_[1995]_ , \new_[1996]_ ,
    \new_[1997]_ , \new_[1998]_ , \new_[1999]_ , \new_[2000]_ ,
    \new_[2001]_ , \new_[2002]_ , \new_[2003]_ , \new_[2004]_ ,
    \new_[2005]_ , \new_[2006]_ , \new_[2007]_ , \new_[2008]_ ,
    \new_[2009]_ , \new_[2010]_ , \new_[2011]_ , \new_[2012]_ ,
    \new_[2013]_ , \new_[2014]_ , \new_[2015]_ , \new_[2016]_ ,
    \new_[2017]_ , \new_[2018]_ , \new_[2019]_ , \new_[2020]_ ,
    \new_[2021]_ , \new_[2022]_ , \new_[2023]_ , \new_[2024]_ ,
    \new_[2025]_ , \new_[2026]_ , \new_[2027]_ , \new_[2028]_ ,
    \new_[2029]_ , \new_[2030]_ , \new_[2031]_ , \new_[2032]_ ,
    \new_[2033]_ , \new_[2034]_ , \new_[2035]_ , \new_[2036]_ ,
    \new_[2037]_ , \new_[2038]_ , \new_[2039]_ , \new_[2040]_ ,
    \new_[2041]_ , \new_[2042]_ , \new_[2043]_ , \new_[2044]_ ,
    \new_[2045]_ , \new_[2046]_ , \new_[2047]_ , \new_[2048]_ ,
    \new_[2049]_ , \new_[2050]_ , \new_[2051]_ , \new_[2052]_ ,
    \new_[2053]_ , \new_[2054]_ , \new_[2055]_ , \new_[2056]_ ,
    \new_[2057]_ , \new_[2058]_ , \new_[2059]_ , \new_[2060]_ ,
    \new_[2061]_ , \new_[2062]_ , \new_[2063]_ , \new_[2064]_ ,
    \new_[2065]_ , \new_[2066]_ , \new_[2067]_ , \new_[2068]_ ,
    \new_[2069]_ , \new_[2070]_ , \new_[2071]_ , \new_[2072]_ ,
    \new_[2073]_ , \new_[2074]_ , \new_[2075]_ , \new_[2076]_ ,
    \new_[2077]_ , \new_[2078]_ , \new_[2079]_ , \new_[2080]_ ,
    \new_[2081]_ , \new_[2082]_ , \new_[2083]_ , \new_[2084]_ ,
    \new_[2085]_ , \new_[2086]_ , \new_[2087]_ , \new_[2088]_ ,
    \new_[2089]_ , \new_[2090]_ , \new_[2091]_ , \new_[2092]_ ,
    \new_[2093]_ , \new_[2094]_ , \new_[2095]_ , \new_[2096]_ ,
    \new_[2097]_ , \new_[2098]_ , \new_[2099]_ , \new_[2100]_ ,
    \new_[2101]_ , \new_[2102]_ , \new_[2103]_ , \new_[2104]_ ,
    \new_[2105]_ , \new_[2106]_ , \new_[2107]_ , \new_[2108]_ ,
    \new_[2109]_ , \new_[2110]_ , \new_[2111]_ , \new_[2112]_ ,
    \new_[2113]_ , \new_[2114]_ , \new_[2115]_ , \new_[2116]_ ,
    \new_[2117]_ , \new_[2118]_ , \new_[2119]_ , \new_[2120]_ ,
    \new_[2121]_ , \new_[2122]_ , \new_[2123]_ , \new_[2124]_ ,
    \new_[2125]_ , \new_[2126]_ , \new_[2127]_ , \new_[2128]_ ,
    \new_[2129]_ , \new_[2130]_ , \new_[2131]_ , \new_[2132]_ ,
    \new_[2133]_ , \new_[2134]_ , \new_[2135]_ , \new_[2136]_ ,
    \new_[2137]_ , \new_[2138]_ , \new_[2139]_ , \new_[2140]_ ,
    \new_[2141]_ , \new_[2142]_ , \new_[2143]_ , \new_[2144]_ ,
    \new_[2145]_ , \new_[2146]_ , \new_[2147]_ , \new_[2148]_ ,
    \new_[2149]_ , \new_[2150]_ , \new_[2151]_ , \new_[2152]_ ,
    \new_[2153]_ , \new_[2154]_ , \new_[2155]_ , \new_[2156]_ ,
    \new_[2157]_ , \new_[2158]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2162]_ , \new_[2163]_ , \new_[2164]_ ,
    \new_[2165]_ , \new_[2166]_ , \new_[2167]_ , \new_[2168]_ ,
    \new_[2169]_ , \new_[2170]_ , \new_[2171]_ , \new_[2172]_ ,
    \new_[2173]_ , \new_[2174]_ , \new_[2175]_ , \new_[2176]_ ,
    \new_[2177]_ , \new_[2178]_ , \new_[2179]_ , \new_[2180]_ ,
    \new_[2181]_ , \new_[2182]_ , \new_[2183]_ , \new_[2184]_ ,
    \new_[2185]_ , \new_[2186]_ , \new_[2187]_ , \new_[2188]_ ,
    \new_[2189]_ , \new_[2190]_ , \new_[2191]_ , \new_[2192]_ ,
    \new_[2193]_ , \new_[2194]_ , \new_[2195]_ , \new_[2196]_ ,
    \new_[2197]_ , \new_[2198]_ , \new_[2199]_ , \new_[2200]_ ,
    \new_[2201]_ , \new_[2202]_ , \new_[2203]_ , \new_[2204]_ ,
    \new_[2205]_ , \new_[2206]_ , \new_[2207]_ , \new_[2208]_ ,
    \new_[2209]_ , \new_[2210]_ , \new_[2211]_ , \new_[2212]_ ,
    \new_[2213]_ , \new_[2214]_ , \new_[2215]_ , \new_[2216]_ ,
    \new_[2217]_ , \new_[2218]_ , \new_[2219]_ , \new_[2220]_ ,
    \new_[2221]_ , \new_[2222]_ , \new_[2223]_ , \new_[2224]_ ,
    \new_[2225]_ , \new_[2226]_ , \new_[2227]_ , \new_[2228]_ ,
    \new_[2229]_ , \new_[2230]_ , \new_[2231]_ , \new_[2232]_ ,
    \new_[2233]_ , \new_[2234]_ , \new_[2235]_ , \new_[2236]_ ,
    \new_[2237]_ , \new_[2239]_ , \new_[2240]_ , \new_[2241]_ ,
    \new_[2242]_ , \new_[2243]_ , \new_[2244]_ , \new_[2245]_ ,
    \new_[2246]_ , \new_[2247]_ , \new_[2248]_ , \new_[2249]_ ,
    \new_[2250]_ , \new_[2251]_ , \new_[2252]_ , \new_[2253]_ ,
    \new_[2254]_ , \new_[2255]_ , \new_[2256]_ , \new_[2257]_ ,
    \new_[2258]_ , \new_[2259]_ , \new_[2260]_ , \new_[2261]_ ,
    \new_[2262]_ , \new_[2263]_ , \new_[2264]_ , \new_[2265]_ ,
    \new_[2266]_ , \new_[2267]_ , \new_[2268]_ , \new_[2269]_ ,
    \new_[2270]_ , \new_[2271]_ , \new_[2272]_ , \new_[2273]_ ,
    \new_[2274]_ , \new_[2275]_ , \new_[2276]_ , \new_[2277]_ ,
    \new_[2278]_ , \new_[2279]_ , \new_[2280]_ , \new_[2281]_ ,
    \new_[2282]_ , \new_[2283]_ , \new_[2284]_ , \new_[2285]_ ,
    \new_[2286]_ , \new_[2287]_ , \new_[2291]_ , \new_[2294]_ ,
    \new_[2295]_ , \new_[2296]_ , \new_[2298]_ , \new_[2299]_ ,
    \new_[2300]_ , \new_[2301]_ , \new_[2302]_ , \new_[2303]_ ,
    \new_[2304]_ , \new_[2305]_ , \new_[2306]_ , \new_[2307]_ ,
    \new_[2308]_ , \new_[2309]_ , \new_[2310]_ , \new_[2311]_ ,
    \new_[2312]_ , \new_[2313]_ , \new_[2314]_ , \new_[2315]_ ,
    \new_[2316]_ , \new_[2317]_ , \new_[2318]_ , \new_[2319]_ ,
    \new_[2320]_ , \new_[2321]_ , \new_[2322]_ , \new_[2323]_ ,
    \new_[2324]_ , \new_[2325]_ , \new_[2326]_ , \new_[2327]_ ,
    \new_[2328]_ , \new_[2329]_ , \new_[2330]_ , \new_[2331]_ ,
    \new_[2332]_ , \new_[2333]_ , \new_[2334]_ , \new_[2335]_ ,
    \new_[2336]_ , \new_[2337]_ , \new_[2338]_ , \new_[2339]_ ,
    \new_[2340]_ , \new_[2341]_ , \new_[2342]_ , \new_[2343]_ ,
    \new_[2344]_ , \new_[2345]_ , \new_[2346]_ , \new_[2347]_ ,
    \new_[2348]_ , \new_[2349]_ , \new_[2350]_ , \new_[2351]_ ,
    \new_[2352]_ , \new_[2353]_ , \new_[2354]_ , \new_[2355]_ ,
    \new_[2356]_ , \new_[2357]_ , \new_[2358]_ , \new_[2359]_ ,
    \new_[2360]_ , \new_[2361]_ , \new_[2362]_ , \new_[2363]_ ,
    \new_[2364]_ , \new_[2365]_ , \new_[2366]_ , \new_[2367]_ ,
    \new_[2368]_ , \new_[2369]_ , \new_[2370]_ , \new_[2371]_ ,
    \new_[2372]_ , \new_[2373]_ , \new_[2374]_ , \new_[2375]_ ,
    \new_[2376]_ , \new_[2377]_ , \new_[2378]_ , \new_[2379]_ ,
    \new_[2380]_ , \new_[2381]_ , \new_[2382]_ , \new_[2383]_ ,
    \new_[2384]_ , \new_[2385]_ , \new_[2386]_ , \new_[2387]_ ,
    \new_[2388]_ , \new_[2389]_ , \new_[2390]_ , \new_[2391]_ ,
    \new_[2392]_ , \new_[2393]_ , \new_[2394]_ , \new_[2395]_ ,
    \new_[2396]_ , \new_[2397]_ , \new_[2398]_ , \new_[2399]_ ,
    \new_[2400]_ , \new_[2401]_ , \new_[2402]_ , \new_[2403]_ ,
    \new_[2404]_ , \new_[2405]_ , \new_[2406]_ , \new_[2407]_ ,
    \new_[2408]_ , \new_[2409]_ , \new_[2410]_ , \new_[2411]_ ,
    \new_[2412]_ , \new_[2413]_ , \new_[2414]_ , \new_[2415]_ ,
    \new_[2416]_ , \new_[2417]_ , \new_[2418]_ , \new_[2420]_ ,
    \new_[2421]_ , \new_[2422]_ , \new_[2423]_ , \new_[2424]_ ,
    \new_[2425]_ , \new_[2426]_ , \new_[2427]_ , \new_[2428]_ ,
    \new_[2429]_ , \new_[2430]_ , \new_[2431]_ , \new_[2432]_ ,
    \new_[2433]_ , \new_[2434]_ , \new_[2435]_ , \new_[2436]_ ,
    \new_[2437]_ , \new_[2438]_ , \new_[2439]_ , \new_[2440]_ ,
    \new_[2441]_ , \new_[2442]_ , \new_[2443]_ , \new_[2444]_ ,
    \new_[2445]_ , \new_[2446]_ , \new_[2447]_ , \new_[2448]_ ,
    \new_[2449]_ , \new_[2450]_ , \new_[2451]_ , \new_[2452]_ ,
    \new_[2453]_ , \new_[2454]_ , \new_[2455]_ , \new_[2456]_ ,
    \new_[2457]_ , \new_[2458]_ , \new_[2459]_ , \new_[2460]_ ,
    \new_[2461]_ , \new_[2462]_ , \new_[2463]_ , \new_[2464]_ ,
    \new_[2465]_ , \new_[2466]_ , \new_[2467]_ , \new_[2468]_ ,
    \new_[2469]_ , \new_[2470]_ , \new_[2471]_ , \new_[2472]_ ,
    \new_[2473]_ , \new_[2474]_ , \new_[2475]_ , \new_[2476]_ ,
    \new_[2477]_ , \new_[2478]_ , \new_[2479]_ , \new_[2480]_ ,
    \new_[2481]_ , \new_[2482]_ , \new_[2483]_ , \new_[2484]_ ,
    \new_[2485]_ , \new_[2486]_ , \new_[2487]_ , \new_[2488]_ ,
    \new_[2490]_ , \new_[2491]_ , \new_[2492]_ , \new_[2493]_ ,
    \new_[2494]_ , \new_[2495]_ , \new_[2496]_ , \new_[2497]_ ,
    \new_[2498]_ , \new_[2499]_ , \new_[2500]_ , \new_[2501]_ ,
    \new_[2502]_ , \new_[2503]_ , \new_[2504]_ , \new_[2505]_ ,
    \new_[2506]_ , \new_[2507]_ , \new_[2508]_ , \new_[2509]_ ,
    \new_[2510]_ , \new_[2511]_ , \new_[2512]_ , \new_[2513]_ ,
    \new_[2514]_ , \new_[2515]_ , \new_[2516]_ , \new_[2517]_ ,
    \new_[2518]_ , \new_[2519]_ , \new_[2520]_ , \new_[2521]_ ,
    \new_[2522]_ , \new_[2523]_ , \new_[2524]_ , \new_[2525]_ ,
    \new_[2526]_ , \new_[2527]_ , \new_[2528]_ , \new_[2529]_ ,
    \new_[2530]_ , \new_[2531]_ , \new_[2532]_ , \new_[2533]_ ,
    \new_[2534]_ , \new_[2535]_ , \new_[2536]_ , \new_[2537]_ ,
    \new_[2538]_ , \new_[2539]_ , \new_[2540]_ , \new_[2541]_ ,
    \new_[2542]_ , \new_[2543]_ , \new_[2544]_ , \new_[2545]_ ,
    \new_[2546]_ , \new_[2547]_ , \new_[2548]_ , \new_[2549]_ ,
    \new_[2550]_ , \new_[2551]_ , \new_[2552]_ , \new_[2553]_ ,
    \new_[2554]_ , \new_[2555]_ , \new_[2556]_ , \new_[2557]_ ,
    \new_[2558]_ , \new_[2559]_ , \new_[2560]_ , \new_[2561]_ ,
    \new_[2562]_ , \new_[2563]_ , \new_[2564]_ , \new_[2565]_ ,
    \new_[2566]_ , \new_[2567]_ , \new_[2568]_ , \new_[2569]_ ,
    \new_[2570]_ , \new_[2571]_ , \new_[2572]_ , \new_[2573]_ ,
    \new_[2574]_ , \new_[2575]_ , \new_[2576]_ , \new_[2577]_ ,
    \new_[2578]_ , \new_[2579]_ , \new_[2580]_ , \new_[2581]_ ,
    \new_[2582]_ , \new_[2583]_ , \new_[2584]_ , \new_[2585]_ ,
    \new_[2586]_ , \new_[2587]_ , \new_[2588]_ , \new_[2589]_ ,
    \new_[2590]_ , \new_[2591]_ , \new_[2592]_ , \new_[2593]_ ,
    \new_[2595]_ , \new_[2596]_ , \new_[2597]_ , \new_[2599]_ ,
    \new_[2600]_ , \new_[2601]_ , \new_[2602]_ , \new_[2605]_ ,
    \new_[2606]_ , \new_[2607]_ , \new_[2608]_ , \new_[2609]_ ,
    \new_[2610]_ , \new_[2611]_ , \new_[2612]_ , \new_[2613]_ ,
    \new_[2614]_ , \new_[2615]_ , \new_[2616]_ , \new_[2617]_ ,
    \new_[2618]_ , \new_[2619]_ , \new_[2620]_ , \new_[2621]_ ,
    \new_[2622]_ , \new_[2623]_ , \new_[2624]_ , \new_[2625]_ ,
    \new_[2626]_ , \new_[2627]_ , \new_[2628]_ , \new_[2629]_ ,
    \new_[2630]_ , \new_[2631]_ , \new_[2632]_ , \new_[2633]_ ,
    \new_[2634]_ , \new_[2635]_ , \new_[2636]_ , \new_[2637]_ ,
    \new_[2638]_ , \new_[2639]_ , \new_[2640]_ , \new_[2641]_ ,
    \new_[2642]_ , \new_[2643]_ , \new_[2644]_ , \new_[2645]_ ,
    \new_[2646]_ , \new_[2647]_ , \new_[2648]_ , \new_[2649]_ ,
    \new_[2650]_ , \new_[2651]_ , \new_[2652]_ , \new_[2653]_ ,
    \new_[2654]_ , \new_[2655]_ , \new_[2656]_ , \new_[2657]_ ,
    \new_[2658]_ , \new_[2659]_ , \new_[2660]_ , \new_[2661]_ ,
    \new_[2662]_ , \new_[2663]_ , \new_[2664]_ , \new_[2665]_ ,
    \new_[2666]_ , \new_[2667]_ , \new_[2668]_ , \new_[2669]_ ,
    \new_[2670]_ , \new_[2671]_ , \new_[2672]_ , \new_[2673]_ ,
    \new_[2674]_ , \new_[2675]_ , \new_[2676]_ , \new_[2677]_ ,
    \new_[2678]_ , \new_[2679]_ , \new_[2680]_ , \new_[2681]_ ,
    \new_[2682]_ , \new_[2683]_ , \new_[2684]_ , \new_[2685]_ ,
    \new_[2686]_ , \new_[2687]_ , \new_[2688]_ , \new_[2689]_ ,
    \new_[2690]_ , \new_[2691]_ , \new_[2692]_ , \new_[2693]_ ,
    \new_[2694]_ , \new_[2695]_ , \new_[2696]_ , \new_[2697]_ ,
    \new_[2698]_ , \new_[2699]_ , \new_[2700]_ , \new_[2701]_ ,
    \new_[2702]_ , \new_[2703]_ , \new_[2704]_ , \new_[2705]_ ,
    \new_[2706]_ , \new_[2707]_ , \new_[2708]_ , \new_[2709]_ ,
    \new_[2710]_ , \new_[2711]_ , \new_[2712]_ , \new_[2713]_ ,
    \new_[2714]_ , \new_[2715]_ , \new_[2716]_ , \new_[2717]_ ,
    \new_[2718]_ , \new_[2719]_ , \new_[2720]_ , \new_[2721]_ ,
    \new_[2722]_ , \new_[2723]_ , \new_[2724]_ , \new_[2725]_ ,
    \new_[2726]_ , \new_[2727]_ , \new_[2728]_ , \new_[2729]_ ,
    \new_[2730]_ , \new_[2731]_ , \new_[2732]_ , \new_[2733]_ ,
    \new_[2734]_ , \new_[2735]_ , \new_[2736]_ , \new_[2737]_ ,
    \new_[2738]_ , \new_[2739]_ , \new_[2740]_ , \new_[2741]_ ,
    \new_[2742]_ , \new_[2743]_ , \new_[2744]_ , \new_[2745]_ ,
    \new_[2746]_ , \new_[2747]_ , \new_[2748]_ , \new_[2749]_ ,
    \new_[2750]_ , \new_[2751]_ , \new_[2752]_ , \new_[2753]_ ,
    \new_[2754]_ , \new_[2755]_ , \new_[2756]_ , \new_[2757]_ ,
    \new_[2758]_ , \new_[2759]_ , \new_[2760]_ , \new_[2761]_ ,
    \new_[2762]_ , \new_[2763]_ , \new_[2764]_ , \new_[2765]_ ,
    \new_[2766]_ , \new_[2767]_ , \new_[2768]_ , \new_[2769]_ ,
    \new_[2770]_ , \new_[2771]_ , \new_[2772]_ , \new_[2773]_ ,
    \new_[2774]_ , \new_[2775]_ , \new_[2776]_ , \new_[2777]_ ,
    \new_[2778]_ , \new_[2779]_ , \new_[2780]_ , \new_[2781]_ ,
    \new_[2782]_ , \new_[2783]_ , \new_[2784]_ , \new_[2785]_ ,
    \new_[2786]_ , \new_[2787]_ , \new_[2788]_ , \new_[2789]_ ,
    \new_[2790]_ , \new_[2791]_ , \new_[2792]_ , \new_[2793]_ ,
    \new_[2794]_ , \new_[2795]_ , \new_[2796]_ , \new_[2797]_ ,
    \new_[2798]_ , \new_[2799]_ , \new_[2800]_ , \new_[2801]_ ,
    \new_[2802]_ , \new_[2803]_ , \new_[2804]_ , \new_[2805]_ ,
    \new_[2806]_ , \new_[2807]_ , \new_[2808]_ , \new_[2809]_ ,
    \new_[2810]_ , \new_[2811]_ , \new_[2812]_ , \new_[2813]_ ,
    \new_[2814]_ , \new_[2815]_ , \new_[2816]_ , \new_[2817]_ ,
    \new_[2818]_ , \new_[2819]_ , \new_[2820]_ , \new_[2821]_ ,
    \new_[2822]_ , \new_[2823]_ , \new_[2824]_ , \new_[2825]_ ,
    \new_[2826]_ , \new_[2827]_ , \new_[2828]_ , \new_[2829]_ ,
    \new_[2830]_ , \new_[2831]_ , \new_[2832]_ , \new_[2833]_ ,
    \new_[2834]_ , \new_[2835]_ , \new_[2836]_ , \new_[2837]_ ,
    \new_[2838]_ , \new_[2839]_ , \new_[2840]_ , \new_[2841]_ ,
    \new_[2842]_ , \new_[2843]_ , \new_[2844]_ , \new_[2845]_ ,
    \new_[2846]_ , \new_[2847]_ , \new_[2848]_ , \new_[2851]_ ,
    \new_[2852]_ , \new_[2853]_ , \new_[2854]_ , \new_[2856]_ ,
    \new_[2858]_ , \new_[2859]_ , \new_[2860]_ , \new_[2861]_ ,
    \new_[2862]_ , \new_[2863]_ , \new_[2864]_ , \new_[2865]_ ,
    \new_[2866]_ , \new_[2867]_ , \new_[2868]_ , \new_[2869]_ ,
    \new_[2870]_ , \new_[2871]_ , \new_[2872]_ , \new_[2873]_ ,
    \new_[2874]_ , \new_[2875]_ , \new_[2876]_ , \new_[2877]_ ,
    \new_[2878]_ , \new_[2879]_ , \new_[2880]_ , \new_[2881]_ ,
    \new_[2882]_ , \new_[2883]_ , \new_[2884]_ , \new_[2885]_ ,
    \new_[2886]_ , \new_[2887]_ , \new_[2888]_ , \new_[2889]_ ,
    \new_[2890]_ , \new_[2891]_ , \new_[2892]_ , \new_[2893]_ ,
    \new_[2894]_ , \new_[2895]_ , \new_[2896]_ , \new_[2897]_ ,
    \new_[2898]_ , \new_[2899]_ , \new_[2900]_ , \new_[2901]_ ,
    \new_[2902]_ , \new_[2903]_ , \new_[2904]_ , \new_[2905]_ ,
    \new_[2906]_ , \new_[2907]_ , \new_[2908]_ , \new_[2909]_ ,
    \new_[2910]_ , \new_[2911]_ , \new_[2912]_ , \new_[2913]_ ,
    \new_[2914]_ , \new_[2915]_ , \new_[2916]_ , \new_[2917]_ ,
    \new_[2918]_ , \new_[2919]_ , \new_[2920]_ , \new_[2921]_ ,
    \new_[2922]_ , \new_[2923]_ , \new_[2924]_ , \new_[2925]_ ,
    \new_[2926]_ , \new_[2927]_ , \new_[2928]_ , \new_[2930]_ ,
    \new_[2932]_ , \new_[2933]_ , \new_[2934]_ , \new_[2935]_ ,
    \new_[2936]_ , \new_[2937]_ , \new_[2938]_ , \new_[2939]_ ,
    \new_[2940]_ , \new_[2941]_ , \new_[2942]_ , \new_[2943]_ ,
    \new_[2944]_ , \new_[2945]_ , \new_[2946]_ , \new_[2947]_ ,
    \new_[2948]_ , \new_[2949]_ , \new_[2950]_ , \new_[2951]_ ,
    \new_[2952]_ , \new_[2953]_ , \new_[2954]_ , \new_[2955]_ ,
    \new_[2956]_ , \new_[2957]_ , \new_[2958]_ , \new_[2959]_ ,
    \new_[2960]_ , \new_[2961]_ , \new_[2962]_ , \new_[2963]_ ,
    \new_[2964]_ , \new_[2965]_ , \new_[2966]_ , \new_[2967]_ ,
    \new_[2968]_ , \new_[2969]_ , \new_[2970]_ , \new_[2971]_ ,
    \new_[2972]_ , \new_[2974]_ , \new_[2975]_ , \new_[2976]_ ,
    \new_[2978]_ , \new_[2979]_ , \new_[2980]_ , \new_[2981]_ ,
    \new_[2982]_ , \new_[2983]_ , \new_[2984]_ , \new_[2985]_ ,
    \new_[2986]_ , \new_[2987]_ , \new_[2988]_ , \new_[2989]_ ,
    \new_[2990]_ , \new_[2991]_ , \new_[2992]_ , \new_[2993]_ ,
    \new_[2994]_ , \new_[2995]_ , \new_[2996]_ , \new_[2997]_ ,
    \new_[2998]_ , \new_[2999]_ , \new_[3000]_ , \new_[3001]_ ,
    \new_[3002]_ , \new_[3003]_ , \new_[3004]_ , \new_[3005]_ ,
    \new_[3006]_ , \new_[3007]_ , \new_[3008]_ , \new_[3009]_ ,
    \new_[3010]_ , \new_[3011]_ , \new_[3012]_ , \new_[3013]_ ,
    \new_[3014]_ , \new_[3015]_ , \new_[3016]_ , \new_[3017]_ ,
    \new_[3018]_ , \new_[3019]_ , \new_[3020]_ , \new_[3021]_ ,
    \new_[3022]_ , \new_[3023]_ , \new_[3024]_ , \new_[3025]_ ,
    \new_[3026]_ , \new_[3027]_ , \new_[3028]_ , \new_[3029]_ ,
    \new_[3030]_ , \new_[3031]_ , \new_[3032]_ , \new_[3033]_ ,
    \new_[3034]_ , \new_[3035]_ , \new_[3036]_ , \new_[3037]_ ,
    \new_[3038]_ , \new_[3039]_ , \new_[3040]_ , \new_[3041]_ ,
    \new_[3042]_ , \new_[3043]_ , \new_[3044]_ , \new_[3045]_ ,
    \new_[3046]_ , \new_[3047]_ , \new_[3048]_ , \new_[3049]_ ,
    \new_[3050]_ , \new_[3051]_ , \new_[3052]_ , \new_[3053]_ ,
    \new_[3054]_ , \new_[3055]_ , \new_[3056]_ , \new_[3057]_ ,
    \new_[3058]_ , \new_[3059]_ , \new_[3060]_ , \new_[3061]_ ,
    \new_[3062]_ , \new_[3063]_ , \new_[3064]_ , \new_[3065]_ ,
    \new_[3066]_ , \new_[3067]_ , \new_[3068]_ , \new_[3069]_ ,
    \new_[3070]_ , \new_[3071]_ , \new_[3072]_ , \new_[3073]_ ,
    \new_[3074]_ , \new_[3075]_ , \new_[3076]_ , \new_[3077]_ ,
    \new_[3078]_ , \new_[3079]_ , \new_[3080]_ , \new_[3081]_ ,
    \new_[3082]_ , \new_[3083]_ , \new_[3084]_ , \new_[3085]_ ,
    \new_[3086]_ , \new_[3087]_ , \new_[3088]_ , \new_[3089]_ ,
    \new_[3090]_ , \new_[3091]_ , \new_[3092]_ , \new_[3093]_ ,
    \new_[3094]_ , \new_[3095]_ , \new_[3096]_ , \new_[3097]_ ,
    \new_[3098]_ , \new_[3099]_ , \new_[3100]_ , \new_[3101]_ ,
    \new_[3102]_ , \new_[3103]_ , \new_[3104]_ , \new_[3105]_ ,
    \new_[3106]_ , \new_[3107]_ , \new_[3108]_ , \new_[3109]_ ,
    \new_[3110]_ , \new_[3111]_ , \new_[3112]_ , \new_[3113]_ ,
    \new_[3114]_ , \new_[3115]_ , \new_[3116]_ , \new_[3117]_ ,
    \new_[3118]_ , \new_[3119]_ , \new_[3120]_ , \new_[3121]_ ,
    \new_[3122]_ , \new_[3123]_ , \new_[3124]_ , \new_[3125]_ ,
    \new_[3126]_ , \new_[3127]_ , \new_[3128]_ , \new_[3129]_ ,
    \new_[3130]_ , \new_[3131]_ , \new_[3132]_ , \new_[3133]_ ,
    \new_[3134]_ , \new_[3135]_ , \new_[3136]_ , \new_[3137]_ ,
    \new_[3138]_ , \new_[3139]_ , \new_[3140]_ , \new_[3141]_ ,
    \new_[3142]_ , \new_[3143]_ , \new_[3144]_ , \new_[3145]_ ,
    \new_[3146]_ , \new_[3147]_ , \new_[3148]_ , \new_[3149]_ ,
    \new_[3150]_ , \new_[3151]_ , \new_[3152]_ , \new_[3153]_ ,
    \new_[3154]_ , \new_[3155]_ , \new_[3156]_ , \new_[3157]_ ,
    \new_[3158]_ , \new_[3159]_ , \new_[3160]_ , \new_[3161]_ ,
    \new_[3164]_ , \new_[3165]_ , \new_[3166]_ , \new_[3167]_ ,
    \new_[3168]_ , \new_[3169]_ , \new_[3170]_ , \new_[3171]_ ,
    \new_[3172]_ , \new_[3173]_ , \new_[3174]_ , \new_[3175]_ ,
    \new_[3176]_ , \new_[3177]_ , \new_[3178]_ , \new_[3179]_ ,
    \new_[3180]_ , \new_[3181]_ , \new_[3182]_ , \new_[3183]_ ,
    \new_[3184]_ , \new_[3185]_ , \new_[3186]_ , \new_[3187]_ ,
    \new_[3188]_ , \new_[3189]_ , \new_[3190]_ , \new_[3191]_ ,
    \new_[3192]_ , \new_[3193]_ , \new_[3194]_ , \new_[3195]_ ,
    \new_[3196]_ , \new_[3197]_ , \new_[3198]_ , \new_[3199]_ ,
    \new_[3200]_ , \new_[3201]_ , \new_[3202]_ , \new_[3203]_ ,
    \new_[3204]_ , \new_[3205]_ , \new_[3206]_ , \new_[3207]_ ,
    \new_[3208]_ , \new_[3209]_ , \new_[3210]_ , \new_[3211]_ ,
    \new_[3212]_ , \new_[3213]_ , \new_[3214]_ , \new_[3215]_ ,
    \new_[3216]_ , \new_[3217]_ , \new_[3218]_ , \new_[3219]_ ,
    \new_[3220]_ , \new_[3221]_ , \new_[3222]_ , \new_[3223]_ ,
    \new_[3224]_ , \new_[3225]_ , \new_[3226]_ , \new_[3227]_ ,
    \new_[3228]_ , \new_[3229]_ , \new_[3230]_ , \new_[3231]_ ,
    \new_[3232]_ , \new_[3233]_ , \new_[3234]_ , \new_[3235]_ ,
    \new_[3236]_ , \new_[3237]_ , \new_[3238]_ , \new_[3239]_ ,
    \new_[3240]_ , \new_[3241]_ , \new_[3242]_ , \new_[3243]_ ,
    \new_[3244]_ , \new_[3245]_ , \new_[3246]_ , \new_[3247]_ ,
    \new_[3248]_ , \new_[3249]_ , \new_[3250]_ , \new_[3251]_ ,
    \new_[3252]_ , \new_[3253]_ , \new_[3254]_ , \new_[3255]_ ,
    \new_[3256]_ , \new_[3257]_ , \new_[3258]_ , \new_[3259]_ ,
    \new_[3260]_ , \new_[3261]_ , \new_[3262]_ , \new_[3263]_ ,
    \new_[3264]_ , \new_[3265]_ , \new_[3266]_ , \new_[3267]_ ,
    \new_[3268]_ , \new_[3269]_ , \new_[3270]_ , \new_[3271]_ ,
    \new_[3272]_ , \new_[3273]_ , \new_[3274]_ , \new_[3275]_ ,
    \new_[3276]_ , \new_[3277]_ , \new_[3278]_ , \new_[3279]_ ,
    \new_[3280]_ , \new_[3281]_ , \new_[3283]_ , \new_[3284]_ ,
    \new_[3285]_ , \new_[3286]_ , \new_[3287]_ , \new_[3288]_ ,
    \new_[3289]_ , \new_[3290]_ , \new_[3291]_ , \new_[3292]_ ,
    \new_[3293]_ , \new_[3294]_ , \new_[3295]_ , \new_[3296]_ ,
    \new_[3297]_ , \new_[3298]_ , \new_[3299]_ , \new_[3300]_ ,
    \new_[3301]_ , \new_[3302]_ , \new_[3303]_ , \new_[3304]_ ,
    \new_[3305]_ , \new_[3306]_ , \new_[3307]_ , \new_[3308]_ ,
    \new_[3309]_ , \new_[3310]_ , \new_[3311]_ , \new_[3312]_ ,
    \new_[3313]_ , \new_[3314]_ , \new_[3315]_ , \new_[3316]_ ,
    \new_[3317]_ , \new_[3318]_ , \new_[3319]_ , \new_[3320]_ ,
    \new_[3321]_ , \new_[3322]_ , \new_[3323]_ , \new_[3324]_ ,
    \new_[3325]_ , \new_[3326]_ , \new_[3327]_ , \new_[3328]_ ,
    \new_[3329]_ , \new_[3330]_ , \new_[3331]_ , \new_[3332]_ ,
    \new_[3333]_ , \new_[3334]_ , \new_[3335]_ , \new_[3336]_ ,
    \new_[3337]_ , \new_[3338]_ , \new_[3339]_ , \new_[3340]_ ,
    \new_[3341]_ , \new_[3342]_ , \new_[3343]_ , \new_[3344]_ ,
    \new_[3345]_ , \new_[3346]_ , \new_[3347]_ , \new_[3348]_ ,
    \new_[3349]_ , \new_[3350]_ , \new_[3351]_ , \new_[3352]_ ,
    \new_[3353]_ , \new_[3354]_ , \new_[3355]_ , \new_[3356]_ ,
    \new_[3357]_ , \new_[3358]_ , \new_[3359]_ , \new_[3360]_ ,
    \new_[3361]_ , \new_[3362]_ , \new_[3363]_ , \new_[3364]_ ,
    \new_[3365]_ , \new_[3366]_ , \new_[3367]_ , \new_[3368]_ ,
    \new_[3369]_ , \new_[3370]_ , \new_[3371]_ , \new_[3372]_ ,
    \new_[3373]_ , \new_[3374]_ , \new_[3375]_ , \new_[3376]_ ,
    \new_[3377]_ , \new_[3378]_ , \new_[3379]_ , \new_[3380]_ ,
    \new_[3381]_ , \new_[3382]_ , \new_[3383]_ , \new_[3384]_ ,
    \new_[3385]_ , \new_[3386]_ , \new_[3387]_ , \new_[3388]_ ,
    \new_[3389]_ , \new_[3390]_ , \new_[3391]_ , \new_[3392]_ ,
    \new_[3393]_ , \new_[3394]_ , \new_[3395]_ , \new_[3396]_ ,
    \new_[3397]_ , \new_[3398]_ , \new_[3399]_ , \new_[3400]_ ,
    \new_[3401]_ , \new_[3402]_ , \new_[3403]_ , \new_[3404]_ ,
    \new_[3405]_ , \new_[3406]_ , \new_[3407]_ , \new_[3408]_ ,
    \new_[3409]_ , \new_[3410]_ , \new_[3411]_ , \new_[3412]_ ,
    \new_[3413]_ , \new_[3414]_ , \new_[3415]_ , \new_[3416]_ ,
    \new_[3417]_ , \new_[3418]_ , \new_[3419]_ , \new_[3420]_ ,
    \new_[3421]_ , \new_[3422]_ , \new_[3423]_ , \new_[3424]_ ,
    \new_[3425]_ , \new_[3426]_ , \new_[3427]_ , \new_[3428]_ ,
    \new_[3429]_ , \new_[3430]_ , \new_[3431]_ , \new_[3432]_ ,
    \new_[3433]_ , \new_[3434]_ , \new_[3435]_ , \new_[3436]_ ,
    \new_[3437]_ , \new_[3438]_ , \new_[3439]_ , \new_[3440]_ ,
    \new_[3441]_ , \new_[3442]_ , \new_[3443]_ , \new_[3444]_ ,
    \new_[3445]_ , \new_[3446]_ , \new_[3447]_ , \new_[3448]_ ,
    \new_[3449]_ , \new_[3450]_ , \new_[3451]_ , \new_[3452]_ ,
    \new_[3453]_ , \new_[3454]_ , \new_[3455]_ , \new_[3456]_ ,
    \new_[3457]_ , \new_[3458]_ , \new_[3459]_ , \new_[3460]_ ,
    \new_[3461]_ , \new_[3462]_ , \new_[3463]_ , \new_[3464]_ ,
    \new_[3465]_ , \new_[3466]_ , \new_[3467]_ , \new_[3468]_ ,
    \new_[3469]_ , \new_[3470]_ , \new_[3471]_ , \new_[3472]_ ,
    \new_[3473]_ , \new_[3474]_ , \new_[3475]_ , \new_[3476]_ ,
    \new_[3477]_ , \new_[3478]_ , \new_[3479]_ , \new_[3480]_ ,
    \new_[3481]_ , \new_[3482]_ , \new_[3483]_ , \new_[3484]_ ,
    \new_[3485]_ , \new_[3486]_ , \new_[3487]_ , \new_[3488]_ ,
    \new_[3489]_ , \new_[3490]_ , \new_[3491]_ , \new_[3492]_ ,
    \new_[3493]_ , \new_[3494]_ , \new_[3495]_ , \new_[3496]_ ,
    \new_[3497]_ , \new_[3498]_ , \new_[3499]_ , \new_[3500]_ ,
    \new_[3501]_ , \new_[3502]_ , \new_[3503]_ , \new_[3504]_ ,
    \new_[3505]_ , \new_[3506]_ , \new_[3507]_ , \new_[3508]_ ,
    \new_[3509]_ , \new_[3510]_ , \new_[3511]_ , \new_[3512]_ ,
    \new_[3513]_ , \new_[3514]_ , \new_[3515]_ , \new_[3516]_ ,
    \new_[3517]_ , \new_[3518]_ , \new_[3519]_ , \new_[3520]_ ,
    \new_[3521]_ , \new_[3522]_ , \new_[3523]_ , \new_[3524]_ ,
    \new_[3525]_ , \new_[3526]_ , \new_[3527]_ , \new_[3528]_ ,
    \new_[3529]_ , \new_[3530]_ , \new_[3531]_ , \new_[3532]_ ,
    \new_[3533]_ , \new_[3534]_ , \new_[3535]_ , \new_[3536]_ ,
    \new_[3537]_ , \new_[3538]_ , \new_[3539]_ , \new_[3540]_ ,
    \new_[3541]_ , \new_[3542]_ , \new_[3543]_ , \new_[3544]_ ,
    \new_[3545]_ , \new_[3546]_ , \new_[3547]_ , \new_[3548]_ ,
    \new_[3549]_ , \new_[3550]_ , \new_[3551]_ , \new_[3552]_ ,
    \new_[3553]_ , \new_[3554]_ , \new_[3555]_ , \new_[3556]_ ,
    \new_[3557]_ , \new_[3558]_ , \new_[3559]_ , \new_[3560]_ ,
    \new_[3561]_ , \new_[3562]_ , \new_[3563]_ , \new_[3564]_ ,
    \new_[3565]_ , \new_[3566]_ , \new_[3567]_ , \new_[3568]_ ,
    \new_[3569]_ , \new_[3570]_ , \new_[3571]_ , \new_[3572]_ ,
    \new_[3573]_ , \new_[3574]_ , \new_[3575]_ , \new_[3576]_ ,
    \new_[3577]_ , \new_[3578]_ , \new_[3579]_ , \new_[3580]_ ,
    \new_[3581]_ , \new_[3582]_ , \new_[3583]_ , \new_[3584]_ ,
    \new_[3585]_ , \new_[3586]_ , \new_[3587]_ , \new_[3588]_ ,
    \new_[3589]_ , \new_[3590]_ , \new_[3591]_ , \new_[3592]_ ,
    \new_[3593]_ , \new_[3594]_ , \new_[3595]_ , \new_[3596]_ ,
    \new_[3597]_ , \new_[3598]_ , \new_[3599]_ , \new_[3600]_ ,
    \new_[3601]_ , \new_[3602]_ , \new_[3603]_ , \new_[3604]_ ,
    \new_[3605]_ , \new_[3606]_ , \new_[3607]_ , \new_[3608]_ ,
    \new_[3609]_ , \new_[3610]_ , \new_[3611]_ , \new_[3612]_ ,
    \new_[3613]_ , \new_[3614]_ , \new_[3615]_ , \new_[3616]_ ,
    \new_[3617]_ , \new_[3618]_ , \new_[3619]_ , \new_[3620]_ ,
    \new_[3621]_ , \new_[3622]_ , \new_[3623]_ , \new_[3624]_ ,
    \new_[3625]_ , \new_[3626]_ , \new_[3627]_ , \new_[3628]_ ,
    \new_[3629]_ , \new_[3630]_ , \new_[3631]_ , \new_[3632]_ ,
    \new_[3633]_ , \new_[3634]_ , \new_[3635]_ , \new_[3636]_ ,
    \new_[3637]_ , \new_[3638]_ , \new_[3639]_ , \new_[3640]_ ,
    \new_[3641]_ , \new_[3642]_ , \new_[3643]_ , \new_[3644]_ ,
    \new_[3645]_ , \new_[3646]_ , \new_[3647]_ , \new_[3648]_ ,
    \new_[3649]_ , \new_[3650]_ , \new_[3651]_ , \new_[3652]_ ,
    \new_[3653]_ , \new_[3654]_ , \new_[3655]_ , \new_[3656]_ ,
    \new_[3657]_ , \new_[3658]_ , \new_[3659]_ , \new_[3660]_ ,
    \new_[3661]_ , \new_[3662]_ , \new_[3663]_ , \new_[3664]_ ,
    \new_[3665]_ , \new_[3666]_ , \new_[3667]_ , \new_[3668]_ ,
    \new_[3669]_ , \new_[3670]_ , \new_[3671]_ , \new_[3672]_ ,
    \new_[3673]_ , \new_[3674]_ , \new_[3675]_ , \new_[3676]_ ,
    \new_[3677]_ , \new_[3678]_ , \new_[3679]_ , \new_[3680]_ ,
    \new_[3681]_ , \new_[3682]_ , \new_[3683]_ , \new_[3684]_ ,
    \new_[3685]_ , \new_[3686]_ , \new_[3687]_ , \new_[3688]_ ,
    \new_[3689]_ , \new_[3690]_ , \new_[3691]_ , \new_[3692]_ ,
    \new_[3693]_ , \new_[3694]_ , \new_[3695]_ , \new_[3696]_ ,
    \new_[3697]_ , \new_[3698]_ , \new_[3699]_ , \new_[3700]_ ,
    \new_[3701]_ , \new_[3702]_ , \new_[3703]_ , \new_[3704]_ ,
    \new_[3705]_ , \new_[3706]_ , \new_[3707]_ , \new_[3708]_ ,
    \new_[3709]_ , \new_[3710]_ , \new_[3711]_ , \new_[3712]_ ,
    \new_[3713]_ , \new_[3714]_ , \new_[3715]_ , \new_[3716]_ ,
    \new_[3717]_ , \new_[3718]_ , \new_[3719]_ , \new_[3720]_ ,
    \new_[3721]_ , \new_[3722]_ , \new_[3723]_ , \new_[3724]_ ,
    \new_[3725]_ , \new_[3726]_ , \new_[3727]_ , \new_[3728]_ ,
    \new_[3729]_ , \new_[3730]_ , \new_[3731]_ , \new_[3732]_ ,
    \new_[3733]_ , \new_[3734]_ , \new_[3735]_ , \new_[3736]_ ,
    \new_[3737]_ , \new_[3738]_ , \new_[3739]_ , \new_[3740]_ ,
    \new_[3741]_ , \new_[3742]_ , \new_[3743]_ , \new_[3744]_ ,
    \new_[3745]_ , \new_[3746]_ , \new_[3747]_ , \new_[3748]_ ,
    \new_[3749]_ , \new_[3750]_ , \new_[3751]_ , \new_[3752]_ ,
    \new_[3753]_ , \new_[3754]_ , \new_[3755]_ , \new_[3756]_ ,
    \new_[3757]_ , \new_[3758]_ , \new_[3759]_ , \new_[3760]_ ,
    \new_[3761]_ , \new_[3762]_ , \new_[3763]_ , \new_[3764]_ ,
    \new_[3765]_ , \new_[3766]_ , \new_[3767]_ , \new_[3768]_ ,
    \new_[3769]_ , \new_[3770]_ , \new_[3771]_ , \new_[3772]_ ,
    \new_[3773]_ , \new_[3774]_ , \new_[3775]_ , \new_[3776]_ ,
    \new_[3777]_ , \new_[3778]_ , \new_[3779]_ , \new_[3780]_ ,
    \new_[3781]_ , \new_[3782]_ , \new_[3783]_ , \new_[3784]_ ,
    \new_[3785]_ , \new_[3786]_ , \new_[3787]_ , \new_[3788]_ ,
    \new_[3789]_ , \new_[3790]_ , \new_[3791]_ , \new_[3792]_ ,
    \new_[3793]_ , \new_[3794]_ , \new_[3795]_ , \new_[3796]_ ,
    \new_[3797]_ , \new_[3798]_ , \new_[3799]_ , \new_[3800]_ ,
    \new_[3801]_ , \new_[3802]_ , \new_[3803]_ , \new_[3804]_ ,
    \new_[3805]_ , \new_[3806]_ , \new_[3807]_ , \new_[3808]_ ,
    \new_[3809]_ , \new_[3810]_ , \new_[3811]_ , \new_[3812]_ ,
    \new_[3813]_ , \new_[3814]_ , \new_[3815]_ , \new_[3816]_ ,
    \new_[3817]_ , \new_[3818]_ , \new_[3819]_ , \new_[3820]_ ,
    \new_[3821]_ , \new_[3822]_ , \new_[3823]_ , \new_[3824]_ ,
    \new_[3825]_ , \new_[3826]_ , \new_[3827]_ , \new_[3828]_ ,
    \new_[3829]_ , \new_[3830]_ , \new_[3831]_ , \new_[3832]_ ,
    \new_[3833]_ , \new_[3834]_ , \new_[3835]_ , \new_[3836]_ ,
    \new_[3837]_ , \new_[3838]_ , \new_[3839]_ , \new_[3840]_ ,
    \new_[3841]_ , \new_[3842]_ , \new_[3843]_ , \new_[3844]_ ,
    \new_[3845]_ , \new_[3846]_ , \new_[3847]_ , \new_[3848]_ ,
    \new_[3849]_ , \new_[3850]_ , \new_[3851]_ , \new_[3852]_ ,
    \new_[3853]_ , \new_[3854]_ , \new_[3855]_ , \new_[3856]_ ,
    \new_[3857]_ , \new_[3858]_ , \new_[3859]_ , \new_[3860]_ ,
    \new_[3861]_ , \new_[3862]_ , \new_[3863]_ , \new_[3864]_ ,
    \new_[3865]_ , \new_[3866]_ , \new_[3867]_ , \new_[3868]_ ,
    \new_[3869]_ , \new_[3870]_ , \new_[3871]_ , \new_[3872]_ ,
    \new_[3873]_ , \new_[3874]_ , \new_[3875]_ , \new_[3876]_ ,
    \new_[3877]_ , \new_[3878]_ , \new_[3879]_ , \new_[3880]_ ,
    \new_[3881]_ , \new_[3882]_ , \new_[3883]_ , \new_[3884]_ ,
    \new_[3885]_ , \new_[3886]_ , \new_[3887]_ , \new_[3888]_ ,
    \new_[3889]_ , \new_[3890]_ , \new_[3891]_ , \new_[3892]_ ,
    \new_[3893]_ , \new_[3894]_ , \new_[3895]_ , \new_[3896]_ ,
    \new_[3897]_ , \new_[3898]_ , \new_[3899]_ , \new_[3900]_ ,
    \new_[3901]_ , \new_[3902]_ , \new_[3903]_ , \new_[3904]_ ,
    \new_[3905]_ , \new_[3906]_ , \new_[3907]_ , \new_[3908]_ ,
    \new_[3909]_ , \new_[3910]_ , \new_[3911]_ , \new_[3912]_ ,
    \new_[3913]_ , \new_[3914]_ , \new_[3915]_ , \new_[3916]_ ,
    \new_[3917]_ , \new_[3918]_ , \new_[3919]_ , \new_[3920]_ ,
    \new_[3921]_ , \new_[3922]_ , \new_[3923]_ , \new_[3924]_ ,
    \new_[3925]_ , \new_[3926]_ , \new_[3927]_ , \new_[3928]_ ,
    \new_[3929]_ , \new_[3930]_ , \new_[3931]_ , \new_[3932]_ ,
    \new_[3933]_ , \new_[3934]_ , \new_[3935]_ , \new_[3936]_ ,
    \new_[3937]_ , \new_[3938]_ , \new_[3939]_ , \new_[3940]_ ,
    \new_[3941]_ , \new_[3942]_ , \new_[3943]_ , \new_[3944]_ ,
    \new_[3945]_ , \new_[3946]_ , \new_[3947]_ , \new_[3948]_ ,
    \new_[3949]_ , \new_[3950]_ , \new_[3951]_ , \new_[3952]_ ,
    \new_[3953]_ , \new_[3954]_ , \new_[3955]_ , \new_[3956]_ ,
    \new_[3957]_ , \new_[3958]_ , \new_[3959]_ , \new_[3960]_ ,
    \new_[3961]_ , \new_[3962]_ , \new_[3963]_ , \new_[3964]_ ,
    \new_[3965]_ , \new_[3966]_ , \new_[3967]_ , \new_[3968]_ ,
    \new_[3969]_ , \new_[3970]_ , \new_[3971]_ , \new_[3972]_ ,
    \new_[3973]_ , \new_[3974]_ , \new_[3975]_ , \new_[3976]_ ,
    \new_[3977]_ , \new_[3978]_ , \new_[3979]_ , \new_[3980]_ ,
    \new_[3981]_ , \new_[3982]_ , \new_[3983]_ , \new_[3984]_ ,
    \new_[3985]_ , \new_[3986]_ , \new_[3987]_ , \new_[3988]_ ,
    \new_[3989]_ , \new_[3990]_ , \new_[3991]_ , \new_[3992]_ ,
    \new_[3993]_ , \new_[3994]_ , \new_[3995]_ , \new_[3996]_ ,
    \new_[3997]_ , \new_[3998]_ , \new_[3999]_ , \new_[4000]_ ,
    \new_[4001]_ , \new_[4002]_ , \new_[4003]_ , \new_[4004]_ ,
    \new_[4005]_ , \new_[4006]_ , \new_[4007]_ , \new_[4008]_ ,
    \new_[4009]_ , \new_[4010]_ , \new_[4011]_ , \new_[4012]_ ,
    \new_[4013]_ , \new_[4014]_ , \new_[4015]_ , \new_[4016]_ ,
    \new_[4017]_ , \new_[4018]_ , \new_[4019]_ , \new_[4020]_ ,
    \new_[4021]_ , \new_[4022]_ , \new_[4023]_ , \new_[4024]_ ,
    \new_[4025]_ , \new_[4026]_ , \new_[4027]_ , \new_[4028]_ ,
    \new_[4029]_ , \new_[4030]_ , \new_[4031]_ , \new_[4032]_ ,
    \new_[4033]_ , \new_[4034]_ , \new_[4035]_ , \new_[4036]_ ,
    \new_[4037]_ , \new_[4038]_ , \new_[4039]_ , \new_[4040]_ ,
    \new_[4041]_ , \new_[4042]_ , \new_[4043]_ , \new_[4044]_ ,
    \new_[4045]_ , \new_[4046]_ , \new_[4047]_ , \new_[4048]_ ,
    \new_[4049]_ , \new_[4050]_ , \new_[4051]_ , \new_[4052]_ ,
    \new_[4053]_ , \new_[4054]_ , \new_[4055]_ , \new_[4056]_ ,
    \new_[4057]_ , \new_[4058]_ , \new_[4059]_ , \new_[4060]_ ,
    \new_[4061]_ , \new_[4062]_ , \new_[4063]_ , \new_[4064]_ ,
    \new_[4065]_ , \new_[4066]_ , \new_[4067]_ , \new_[4068]_ ,
    \new_[4069]_ , \new_[4070]_ , \new_[4071]_ , \new_[4072]_ ,
    \new_[4073]_ , \new_[4074]_ , \new_[4075]_ , \new_[4076]_ ,
    \new_[4077]_ , \new_[4078]_ , \new_[4079]_ , \new_[4080]_ ,
    \new_[4081]_ , \new_[4082]_ , \new_[4083]_ , \new_[4084]_ ,
    \new_[4085]_ , \new_[4086]_ , \new_[4087]_ , \new_[4088]_ ,
    \new_[4089]_ , \new_[4090]_ , \new_[4091]_ , \new_[4092]_ ,
    \new_[4093]_ , \new_[4094]_ , \new_[4095]_ , \new_[4096]_ ,
    \new_[4097]_ , \new_[4098]_ , \new_[4099]_ , \new_[4100]_ ,
    \new_[4101]_ , \new_[4102]_ , \new_[4103]_ , \new_[4104]_ ,
    \new_[4105]_ , \new_[4106]_ , \new_[4107]_ , \new_[4108]_ ,
    \new_[4109]_ , \new_[4110]_ , \new_[4111]_ , \new_[4112]_ ,
    \new_[4113]_ , \new_[4114]_ , \new_[4115]_ , \new_[4116]_ ,
    \new_[4117]_ , \new_[4118]_ , \new_[4119]_ , \new_[4120]_ ,
    \new_[4121]_ , \new_[4122]_ , \new_[4123]_ , \new_[4124]_ ,
    \new_[4125]_ , \new_[4126]_ , \new_[4127]_ , \new_[4128]_ ,
    \new_[4129]_ , \new_[4130]_ , \new_[4131]_ , \new_[4132]_ ,
    \new_[4133]_ , \new_[4134]_ , \new_[4135]_ , \new_[4136]_ ,
    \new_[4137]_ , \new_[4138]_ , \new_[4139]_ , \new_[4140]_ ,
    \new_[4141]_ , \new_[4142]_ , \new_[4143]_ , \new_[4144]_ ,
    \new_[4145]_ , \new_[4146]_ , \new_[4147]_ , \new_[4148]_ ,
    \new_[4149]_ , \new_[4150]_ , \new_[4151]_ , \new_[4152]_ ,
    \new_[4153]_ , \new_[4154]_ , \new_[4155]_ , \new_[4156]_ ,
    \new_[4157]_ , \new_[4158]_ , \new_[4159]_ , \new_[4160]_ ,
    \new_[4161]_ , \new_[4162]_ , \new_[4163]_ , \new_[4164]_ ,
    \new_[4165]_ , \new_[4166]_ , \new_[4167]_ , \new_[4168]_ ,
    \new_[4169]_ , \new_[4170]_ , \new_[4171]_ , \new_[4172]_ ,
    \new_[4173]_ , \new_[4174]_ , \new_[4175]_ , \new_[4176]_ ,
    \new_[4177]_ , \new_[4178]_ , \new_[4179]_ , \new_[4180]_ ,
    \new_[4181]_ , \new_[4182]_ , \new_[4183]_ , \new_[4184]_ ,
    \new_[4185]_ , \new_[4186]_ , \new_[4187]_ , \new_[4188]_ ,
    \new_[4189]_ , \new_[4190]_ , \new_[4191]_ , \new_[4192]_ ,
    \new_[4193]_ , \new_[4194]_ , \new_[4195]_ , \new_[4196]_ ,
    \new_[4197]_ , \new_[4198]_ , \new_[4199]_ , \new_[4200]_ ,
    \new_[4201]_ , \new_[4202]_ , \new_[4203]_ , \new_[4204]_ ,
    \new_[4205]_ , \new_[4206]_ , \new_[4207]_ , \new_[4208]_ ,
    \new_[4209]_ , \new_[4210]_ , \new_[4211]_ , \new_[4212]_ ,
    \new_[4213]_ , \new_[4214]_ , \new_[4215]_ , \new_[4216]_ ,
    \new_[4217]_ , \new_[4218]_ , \new_[4219]_ , \new_[4220]_ ,
    \new_[4221]_ , \new_[4222]_ , \new_[4223]_ , \new_[4224]_ ,
    \new_[4225]_ , \new_[4226]_ , \new_[4227]_ , \new_[4228]_ ,
    \new_[4229]_ , \new_[4230]_ , \new_[4231]_ , \new_[4232]_ ,
    \new_[4233]_ , \new_[4234]_ , \new_[4235]_ , \new_[4236]_ ,
    \new_[4237]_ , \new_[4238]_ , \new_[4239]_ , \new_[4240]_ ,
    \new_[4241]_ , \new_[4242]_ , \new_[4243]_ , \new_[4244]_ ,
    \new_[4245]_ , \new_[4246]_ , \new_[4247]_ , \new_[4248]_ ,
    \new_[4249]_ , \new_[4250]_ , \new_[4251]_ , \new_[4252]_ ,
    \new_[4253]_ , \new_[4254]_ , \new_[4255]_ , \new_[4256]_ ,
    \new_[4257]_ , \new_[4258]_ , \new_[4259]_ , \new_[4260]_ ,
    \new_[4261]_ , \new_[4262]_ , \new_[4263]_ , \new_[4264]_ ,
    \new_[4265]_ , \new_[4266]_ , \new_[4267]_ , \new_[4268]_ ,
    \new_[4269]_ , \new_[4270]_ , \new_[4271]_ , \new_[4272]_ ,
    \new_[4273]_ , \new_[4274]_ , \new_[4275]_ , \new_[4276]_ ,
    \new_[4277]_ , \new_[4278]_ , \new_[4279]_ , \new_[4280]_ ,
    \new_[4281]_ , \new_[4282]_ , \new_[4283]_ , \new_[4284]_ ,
    \new_[4285]_ , \new_[4286]_ , \new_[4287]_ , \new_[4288]_ ,
    \new_[4289]_ , \new_[4290]_ , \new_[4291]_ , \new_[4292]_ ,
    \new_[4293]_ , \new_[4294]_ , \new_[4295]_ , \new_[4296]_ ,
    \new_[4297]_ , \new_[4298]_ , \new_[4299]_ , \new_[4300]_ ,
    \new_[4301]_ , \new_[4302]_ , \new_[4303]_ , \new_[4304]_ ,
    \new_[4305]_ , \new_[4306]_ , \new_[4307]_ , \new_[4308]_ ,
    \new_[4309]_ , \new_[4310]_ , \new_[4311]_ , \new_[4312]_ ,
    \new_[4313]_ , \new_[4314]_ , \new_[4315]_ , \new_[4316]_ ,
    \new_[4317]_ , \new_[4318]_ , \new_[4319]_ , \new_[4320]_ ,
    \new_[4321]_ , \new_[4322]_ , \new_[4323]_ , \new_[4324]_ ,
    \new_[4325]_ , \new_[4326]_ , \new_[4327]_ , \new_[4328]_ ,
    \new_[4329]_ , \new_[4330]_ , \new_[4331]_ , \new_[4332]_ ,
    \new_[4333]_ , \new_[4334]_ , \new_[4335]_ , \new_[4336]_ ,
    \new_[4337]_ , \new_[4338]_ , \new_[4339]_ , \new_[4340]_ ,
    \new_[4341]_ , \new_[4342]_ , \new_[4343]_ , \new_[4344]_ ,
    \new_[4345]_ , \new_[4346]_ , \new_[4347]_ , \new_[4348]_ ,
    \new_[4349]_ , \new_[4350]_ , \new_[4351]_ , \new_[4352]_ ,
    \new_[4353]_ , \new_[4354]_ , \new_[4355]_ , \new_[4356]_ ,
    \new_[4357]_ , \new_[4358]_ , \new_[4359]_ , \new_[4360]_ ,
    \new_[4361]_ , \new_[4362]_ , \new_[4363]_ , \new_[4364]_ ,
    \new_[4365]_ , \new_[4366]_ , \new_[4367]_ , \new_[4368]_ ,
    \new_[4369]_ , \new_[4370]_ , \new_[4371]_ , \new_[4372]_ ,
    \new_[4373]_ , \new_[4374]_ , \new_[4375]_ , \new_[4376]_ ,
    \new_[4377]_ , \new_[4378]_ , \new_[4379]_ , \new_[4380]_ ,
    \new_[4381]_ , \new_[4382]_ , \new_[4383]_ , \new_[4384]_ ,
    \new_[4385]_ , \new_[4386]_ , \new_[4387]_ , \new_[4388]_ ,
    \new_[4389]_ , \new_[4390]_ , \new_[4391]_ , \new_[4392]_ ,
    \new_[4393]_ , \new_[4394]_ , \new_[4395]_ , \new_[4396]_ ,
    \new_[4397]_ , \new_[4398]_ , \new_[4399]_ , \new_[4400]_ ,
    \new_[4401]_ , \new_[4402]_ , \new_[4403]_ , \new_[4404]_ ,
    \new_[4405]_ , \new_[4406]_ , \new_[4407]_ , \new_[4408]_ ,
    \new_[4410]_ , \new_[4411]_ , \new_[4412]_ , \new_[4413]_ ,
    \new_[4414]_ , \new_[4415]_ , \new_[4416]_ , \new_[4417]_ ,
    \new_[4418]_ , \new_[4419]_ , \new_[4420]_ , \new_[4422]_ ,
    \new_[4423]_ , \new_[4424]_ , \new_[4425]_ , \new_[4426]_ ,
    \new_[4427]_ , \new_[4428]_ , \new_[4430]_ , \new_[4431]_ ,
    \new_[4432]_ , \new_[4434]_ , \new_[4435]_ , \new_[4436]_ ,
    \new_[4437]_ , \new_[4438]_ , \new_[4439]_ , \new_[4440]_ ,
    \new_[4441]_ , \new_[4442]_ , \new_[4443]_ , \new_[4444]_ ,
    \new_[4445]_ , \new_[4447]_ , \new_[4448]_ , \new_[4449]_ ,
    \new_[4450]_ , \new_[4451]_ , \new_[4452]_ , \new_[4453]_ ,
    \new_[4454]_ , \new_[4455]_ , \new_[4456]_ , \new_[4457]_ ,
    \new_[4458]_ , \new_[4459]_ , \new_[4460]_ , \new_[4461]_ ,
    \new_[4462]_ , \new_[4463]_ , \new_[4464]_ , \new_[4466]_ ,
    \new_[4467]_ , \new_[4468]_ , \new_[4469]_ , \new_[4470]_ ,
    \new_[4471]_ , \new_[4472]_ , \new_[4473]_ , \new_[4474]_ ,
    \new_[4475]_ , \new_[4476]_ , \new_[4477]_ , \new_[4478]_ ,
    \new_[4480]_ , \new_[4481]_ , \new_[4482]_ , \new_[4483]_ ,
    \new_[4484]_ , \new_[4485]_ , \new_[4486]_ , \new_[4487]_ ,
    \new_[4488]_ , \new_[4489]_ , \new_[4490]_ , \new_[4491]_ ,
    \new_[4492]_ , \new_[4493]_ , \new_[4494]_ , \new_[4495]_ ,
    \new_[4496]_ , \new_[4497]_ , \new_[4498]_ , \new_[4499]_ ,
    \new_[4500]_ , \new_[4501]_ , \new_[4502]_ , \new_[4503]_ ,
    \new_[4504]_ , \new_[4505]_ , \new_[4506]_ , \new_[4507]_ ,
    \new_[4508]_ , \new_[4509]_ , \new_[4510]_ , \new_[4511]_ ,
    \new_[4513]_ , \new_[4514]_ , \new_[4515]_ , \new_[4516]_ ,
    \new_[4517]_ , \new_[4518]_ , \new_[4519]_ , \new_[4520]_ ,
    \new_[4521]_ , \new_[4522]_ , \new_[4523]_ , \new_[4524]_ ,
    \new_[4525]_ , \new_[4526]_ , \new_[4527]_ , \new_[4528]_ ,
    \new_[4529]_ , \new_[4530]_ , \new_[4531]_ , \new_[4532]_ ,
    \new_[4533]_ , \new_[4534]_ , \new_[4535]_ , \new_[4536]_ ,
    \new_[4537]_ , \new_[4538]_ , \new_[4539]_ , \new_[4540]_ ,
    \new_[4541]_ , \new_[4542]_ , \new_[4543]_ , \new_[4544]_ ,
    \new_[4545]_ , \new_[4546]_ , \new_[4547]_ , \new_[4548]_ ,
    \new_[4549]_ , \new_[4550]_ , \new_[4551]_ , \new_[4552]_ ,
    \new_[4553]_ , \new_[4554]_ , \new_[4555]_ , \new_[4556]_ ,
    \new_[4557]_ , \new_[4558]_ , \new_[4559]_ , \new_[4560]_ ,
    \new_[4561]_ , \new_[4562]_ , \new_[4563]_ , \new_[4564]_ ,
    \new_[4565]_ , \new_[4566]_ , \new_[4567]_ , \new_[4568]_ ,
    \new_[4569]_ , \new_[4570]_ , \new_[4571]_ , \new_[4572]_ ,
    \new_[4573]_ , \new_[4574]_ , \new_[4575]_ , \new_[4576]_ ,
    \new_[4577]_ , \new_[4578]_ , \new_[4579]_ , \new_[4580]_ ,
    \new_[4581]_ , \new_[4582]_ , \new_[4583]_ , \new_[4584]_ ,
    \new_[4585]_ , \new_[4587]_ , \new_[4588]_ , \new_[4589]_ ,
    \new_[4590]_ , \new_[4591]_ , \new_[4592]_ , \new_[4593]_ ,
    \new_[4594]_ , \new_[4595]_ , \new_[4596]_ , \new_[4597]_ ,
    \new_[4598]_ , \new_[4599]_ , \new_[4600]_ , \new_[4601]_ ,
    \new_[4602]_ , \new_[4603]_ , \new_[4604]_ , \new_[4605]_ ,
    \new_[4606]_ , \new_[4607]_ , \new_[4608]_ , \new_[4609]_ ,
    \new_[4610]_ , \new_[4611]_ , \new_[4612]_ , \new_[4613]_ ,
    \new_[4614]_ , \new_[4615]_ , \new_[4616]_ , \new_[4617]_ ,
    \new_[4618]_ , \new_[4619]_ , \new_[4620]_ , \new_[4622]_ ,
    \new_[4623]_ , \new_[4624]_ , \new_[4625]_ , \new_[4626]_ ,
    \new_[4627]_ , \new_[4628]_ , \new_[4629]_ , \new_[4630]_ ,
    \new_[4631]_ , \new_[4632]_ , \new_[4633]_ , \new_[4634]_ ,
    \new_[4635]_ , \new_[4636]_ , \new_[4637]_ , \new_[4638]_ ,
    \new_[4639]_ , \new_[4640]_ , \new_[4641]_ , \new_[4642]_ ,
    \new_[4643]_ , \new_[4644]_ , \new_[4645]_ , \new_[4646]_ ,
    \new_[4647]_ , \new_[4648]_ , \new_[4649]_ , \new_[4650]_ ,
    \new_[4651]_ , \new_[4652]_ , \new_[4653]_ , \new_[4654]_ ,
    \new_[4655]_ , \new_[4656]_ , \new_[4657]_ , \new_[4658]_ ,
    \new_[4659]_ , \new_[4660]_ , \new_[4661]_ , \new_[4662]_ ,
    \new_[4663]_ , \new_[4664]_ , \new_[4665]_ , \new_[4666]_ ,
    \new_[4667]_ , \new_[4668]_ , \new_[4669]_ , \new_[4670]_ ,
    \new_[4671]_ , \new_[4672]_ , \new_[4673]_ , \new_[4674]_ ,
    \new_[4675]_ , \new_[4676]_ , \new_[4677]_ , \new_[4678]_ ,
    \new_[4680]_ , \new_[4681]_ , \new_[4682]_ , \new_[4683]_ ,
    \new_[4684]_ , \new_[4685]_ , \new_[4686]_ , \new_[4687]_ ,
    \new_[4688]_ , \new_[4689]_ , \new_[4690]_ , \new_[4691]_ ,
    \new_[4692]_ , \new_[4693]_ , \new_[4694]_ , \new_[4695]_ ,
    \new_[4696]_ , \new_[4697]_ , \new_[4698]_ , \new_[4699]_ ,
    \new_[4700]_ , \new_[4701]_ , \new_[4702]_ , \new_[4703]_ ,
    \new_[4704]_ , \new_[4706]_ , \new_[4707]_ , \new_[4708]_ ,
    \new_[4709]_ , \new_[4710]_ , \new_[4711]_ , \new_[4712]_ ,
    \new_[4713]_ , \new_[4714]_ , \new_[4715]_ , \new_[4716]_ ,
    \new_[4717]_ , \new_[4718]_ , \new_[4719]_ , \new_[4720]_ ,
    \new_[4721]_ , \new_[4722]_ , \new_[4723]_ , \new_[4724]_ ,
    \new_[4725]_ , \new_[4726]_ , \new_[4727]_ , \new_[4728]_ ,
    \new_[4729]_ , \new_[4730]_ , \new_[4731]_ , \new_[4732]_ ,
    \new_[4733]_ , \new_[4734]_ , \new_[4735]_ , \new_[4736]_ ,
    \new_[4737]_ , \new_[4738]_ , \new_[4739]_ , \new_[4740]_ ,
    \new_[4741]_ , \new_[4742]_ , \new_[4743]_ , \new_[4744]_ ,
    \new_[4745]_ , \new_[4746]_ , \new_[4747]_ , \new_[4749]_ ,
    \new_[4750]_ , \new_[4751]_ , \new_[4752]_ , \new_[4753]_ ,
    \new_[4754]_ , \new_[4755]_ , \new_[4756]_ , \new_[4757]_ ,
    \new_[4758]_ , \new_[4759]_ , \new_[4760]_ , \new_[4761]_ ,
    \new_[4762]_ , \new_[4763]_ , \new_[4764]_ , \new_[4765]_ ,
    \new_[4766]_ , \new_[4767]_ , \new_[4768]_ , \new_[4769]_ ,
    \new_[4771]_ , \new_[4772]_ , \new_[4773]_ , \new_[4774]_ ,
    \new_[4775]_ , \new_[4776]_ , \new_[4777]_ , \new_[4778]_ ,
    \new_[4779]_ , \new_[4780]_ , \new_[4781]_ , \new_[4782]_ ,
    \new_[4783]_ , \new_[4784]_ , \new_[4785]_ , \new_[4786]_ ,
    \new_[4787]_ , \new_[4788]_ , \new_[4789]_ , \new_[4790]_ ,
    \new_[4791]_ , \new_[4792]_ , \new_[4793]_ , \new_[4794]_ ,
    \new_[4795]_ , \new_[4796]_ , \new_[4797]_ , \new_[4798]_ ,
    \new_[4799]_ , \new_[4800]_ , \new_[4801]_ , \new_[4802]_ ,
    \new_[4803]_ , \new_[4804]_ , \new_[4805]_ , \new_[4806]_ ,
    \new_[4807]_ , \new_[4808]_ , \new_[4809]_ , \new_[4810]_ ,
    \new_[4811]_ , \new_[4812]_ , \new_[4813]_ , \new_[4814]_ ,
    \new_[4815]_ , \new_[4816]_ , \new_[4817]_ , \new_[4818]_ ,
    \new_[4819]_ , \new_[4820]_ , \new_[4821]_ , \new_[4822]_ ,
    \new_[4823]_ , \new_[4824]_ , \new_[4825]_ , \new_[4826]_ ,
    \new_[4827]_ , \new_[4828]_ , \new_[4829]_ , \new_[4830]_ ,
    \new_[4831]_ , \new_[4832]_ , \new_[4833]_ , \new_[4836]_ ,
    \new_[4837]_ , \new_[4838]_ , \new_[4839]_ , \new_[4840]_ ,
    \new_[4841]_ , \new_[4842]_ , \new_[4843]_ , \new_[4844]_ ,
    \new_[4845]_ , \new_[4846]_ , \new_[4847]_ , \new_[4848]_ ,
    \new_[4849]_ , \new_[4850]_ , \new_[4851]_ , \new_[4852]_ ,
    \new_[4853]_ , \new_[4854]_ , \new_[4855]_ , \new_[4856]_ ,
    \new_[4857]_ , \new_[4858]_ , \new_[4859]_ , \new_[4860]_ ,
    \new_[4861]_ , \new_[4862]_ , \new_[4863]_ , \new_[4864]_ ,
    \new_[4865]_ , \new_[4866]_ , \new_[4867]_ , \new_[4868]_ ,
    \new_[4869]_ , \new_[4870]_ , \new_[4871]_ , \new_[4872]_ ,
    \new_[4873]_ , \new_[4874]_ , \new_[4875]_ , \new_[4877]_ ,
    \new_[4878]_ , \new_[4879]_ , \new_[4880]_ , \new_[4881]_ ,
    \new_[4882]_ , \new_[4883]_ , \new_[4884]_ , \new_[4885]_ ,
    \new_[4886]_ , \new_[4887]_ , \new_[4888]_ , \new_[4889]_ ,
    \new_[4890]_ , \new_[4891]_ , \new_[4892]_ , \new_[4893]_ ,
    \new_[4894]_ , \new_[4895]_ , \new_[4896]_ , \new_[4897]_ ,
    \new_[4898]_ , \new_[4899]_ , \new_[4901]_ , \new_[4902]_ ,
    \new_[4903]_ , \new_[4904]_ , \new_[4905]_ , \new_[4906]_ ,
    \new_[4907]_ , \new_[4908]_ , \new_[4909]_ , \new_[4910]_ ,
    \new_[4911]_ , \new_[4912]_ , \new_[4913]_ , \new_[4914]_ ,
    \new_[4916]_ , \new_[4917]_ , \new_[4918]_ , \new_[4919]_ ,
    \new_[4920]_ , \new_[4921]_ , \new_[4922]_ , \new_[4924]_ ,
    \new_[4925]_ , \new_[4926]_ , \new_[4927]_ , \new_[4928]_ ,
    \new_[4929]_ , \new_[4930]_ , \new_[4931]_ , \new_[4932]_ ,
    \new_[4933]_ , \new_[4934]_ , \new_[4935]_ , \new_[4936]_ ,
    \new_[4937]_ , \new_[4938]_ , \new_[4939]_ , \new_[4940]_ ,
    \new_[4942]_ , \new_[4943]_ , \new_[4944]_ , \new_[4945]_ ,
    \new_[4946]_ , \new_[4947]_ , \new_[4948]_ , \new_[4949]_ ,
    \new_[4950]_ , \new_[4951]_ , \new_[4952]_ , \new_[4953]_ ,
    \new_[4954]_ , \new_[4955]_ , \new_[4956]_ , \new_[4957]_ ,
    \new_[4958]_ , \new_[4959]_ , \new_[4960]_ , \new_[4961]_ ,
    \new_[4962]_ , \new_[4963]_ , \new_[4964]_ , \new_[4965]_ ,
    \new_[4966]_ , \new_[4967]_ , \new_[4968]_ , \new_[4969]_ ,
    \new_[4970]_ , \new_[4971]_ , \new_[4972]_ , \new_[4973]_ ,
    \new_[4974]_ , \new_[4975]_ , \new_[4976]_ , \new_[4977]_ ,
    \new_[4978]_ , \new_[4980]_ , \new_[4981]_ , \new_[4982]_ ,
    \new_[4983]_ , \new_[4984]_ , \new_[4985]_ , \new_[4986]_ ,
    \new_[4987]_ , \new_[4988]_ , \new_[4989]_ , \new_[4990]_ ,
    \new_[4992]_ , \new_[4993]_ , \new_[4994]_ , \new_[4995]_ ,
    \new_[4996]_ , \new_[4997]_ , \new_[4998]_ , \new_[4999]_ ,
    \new_[5000]_ , \new_[5001]_ , \new_[5002]_ , \new_[5003]_ ,
    \new_[5004]_ , \new_[5005]_ , \new_[5007]_ , \new_[5008]_ ,
    \new_[5009]_ , \new_[5010]_ , \new_[5011]_ , \new_[5012]_ ,
    \new_[5013]_ , \new_[5014]_ , \new_[5015]_ , \new_[5016]_ ,
    \new_[5017]_ , \new_[5018]_ , \new_[5019]_ , \new_[5020]_ ,
    \new_[5021]_ , \new_[5022]_ , \new_[5023]_ , \new_[5024]_ ,
    \new_[5025]_ , \new_[5026]_ , \new_[5027]_ , \new_[5028]_ ,
    \new_[5030]_ , \new_[5031]_ , \new_[5032]_ , \new_[5033]_ ,
    \new_[5034]_ , \new_[5035]_ , \new_[5036]_ , \new_[5037]_ ,
    \new_[5038]_ , \new_[5039]_ , \new_[5040]_ , \new_[5041]_ ,
    \new_[5042]_ , \new_[5043]_ , \new_[5044]_ , \new_[5045]_ ,
    \new_[5046]_ , \new_[5047]_ , \new_[5048]_ , \new_[5049]_ ,
    \new_[5050]_ , \new_[5051]_ , \new_[5052]_ , \new_[5053]_ ,
    \new_[5054]_ , \new_[5055]_ , \new_[5056]_ , \new_[5057]_ ,
    \new_[5058]_ , \new_[5059]_ , \new_[5060]_ , \new_[5061]_ ,
    \new_[5062]_ , \new_[5063]_ , \new_[5064]_ , \new_[5065]_ ,
    \new_[5066]_ , \new_[5067]_ , \new_[5068]_ , \new_[5069]_ ,
    \new_[5070]_ , \new_[5071]_ , \new_[5072]_ , \new_[5073]_ ,
    \new_[5075]_ , \new_[5076]_ , \new_[5077]_ , \new_[5078]_ ,
    \new_[5079]_ , \new_[5080]_ , \new_[5081]_ , \new_[5082]_ ,
    \new_[5083]_ , \new_[5084]_ , \new_[5085]_ , \new_[5086]_ ,
    \new_[5087]_ , \new_[5088]_ , \new_[5089]_ , \new_[5090]_ ,
    \new_[5091]_ , \new_[5092]_ , \new_[5093]_ , \new_[5094]_ ,
    \new_[5095]_ , \new_[5096]_ , \new_[5097]_ , \new_[5098]_ ,
    \new_[5099]_ , \new_[5100]_ , \new_[5101]_ , \new_[5102]_ ,
    \new_[5103]_ , \new_[5104]_ , \new_[5105]_ , \new_[5106]_ ,
    \new_[5107]_ , \new_[5108]_ , \new_[5109]_ , \new_[5110]_ ,
    \new_[5111]_ , \new_[5112]_ , \new_[5113]_ , \new_[5114]_ ,
    \new_[5115]_ , \new_[5116]_ , \new_[5117]_ , \new_[5118]_ ,
    \new_[5119]_ , \new_[5120]_ , \new_[5121]_ , \new_[5122]_ ,
    \new_[5123]_ , \new_[5124]_ , \new_[5125]_ , \new_[5126]_ ,
    \new_[5127]_ , \new_[5128]_ , \new_[5129]_ , \new_[5130]_ ,
    \new_[5131]_ , \new_[5132]_ , \new_[5133]_ , \new_[5134]_ ,
    \new_[5135]_ , \new_[5136]_ , \new_[5137]_ , \new_[5138]_ ,
    \new_[5139]_ , \new_[5140]_ , \new_[5141]_ , \new_[5142]_ ,
    \new_[5143]_ , \new_[5144]_ , \new_[5145]_ , \new_[5146]_ ,
    \new_[5147]_ , \new_[5148]_ , \new_[5149]_ , \new_[5150]_ ,
    \new_[5151]_ , \new_[5152]_ , \new_[5153]_ , \new_[5154]_ ,
    \new_[5155]_ , \new_[5156]_ , \new_[5157]_ , \new_[5158]_ ,
    \new_[5159]_ , \new_[5160]_ , \new_[5161]_ , \new_[5163]_ ,
    \new_[5164]_ , \new_[5165]_ , \new_[5166]_ , \new_[5167]_ ,
    \new_[5168]_ , \new_[5169]_ , \new_[5170]_ , \new_[5171]_ ,
    \new_[5172]_ , \new_[5173]_ , \new_[5174]_ , \new_[5175]_ ,
    \new_[5176]_ , \new_[5177]_ , \new_[5178]_ , \new_[5179]_ ,
    \new_[5180]_ , \new_[5181]_ , \new_[5182]_ , \new_[5183]_ ,
    \new_[5185]_ , \new_[5186]_ , \new_[5187]_ , \new_[5188]_ ,
    \new_[5189]_ , \new_[5190]_ , \new_[5191]_ , \new_[5192]_ ,
    \new_[5193]_ , \new_[5194]_ , \new_[5195]_ , \new_[5196]_ ,
    \new_[5197]_ , \new_[5198]_ , \new_[5199]_ , \new_[5200]_ ,
    \new_[5201]_ , \new_[5202]_ , \new_[5203]_ , \new_[5204]_ ,
    \new_[5205]_ , \new_[5207]_ , \new_[5208]_ , \new_[5209]_ ,
    \new_[5210]_ , \new_[5211]_ , \new_[5212]_ , \new_[5213]_ ,
    \new_[5214]_ , \new_[5215]_ , \new_[5216]_ , \new_[5217]_ ,
    \new_[5218]_ , \new_[5219]_ , \new_[5220]_ , \new_[5221]_ ,
    \new_[5222]_ , \new_[5223]_ , \new_[5224]_ , \new_[5225]_ ,
    \new_[5226]_ , \new_[5227]_ , \new_[5228]_ , \new_[5229]_ ,
    \new_[5230]_ , \new_[5231]_ , \new_[5232]_ , \new_[5233]_ ,
    \new_[5234]_ , \new_[5235]_ , \new_[5236]_ , \new_[5237]_ ,
    \new_[5240]_ , \new_[5241]_ , \new_[5242]_ , \new_[5243]_ ,
    \new_[5244]_ , \new_[5245]_ , \new_[5246]_ , \new_[5247]_ ,
    \new_[5248]_ , \new_[5249]_ , \new_[5250]_ , \new_[5255]_ ,
    \new_[5256]_ , \new_[5257]_ , \new_[5258]_ , \new_[5259]_ ,
    \new_[5260]_ , \new_[5261]_ , \new_[5262]_ , \new_[5263]_ ,
    \new_[5266]_ , \new_[5267]_ , \new_[5268]_ , \new_[5269]_ ,
    \new_[5270]_ , \new_[5271]_ , \new_[5272]_ , \new_[5273]_ ,
    \new_[5276]_ , \new_[5277]_ , \new_[5278]_ , \new_[5279]_ ,
    \new_[5280]_ , \new_[5281]_ , \new_[5282]_ , \new_[5283]_ ,
    \new_[5284]_ , \new_[5285]_ , \new_[5286]_ , \new_[5287]_ ,
    \new_[5288]_ , \new_[5289]_ , \new_[5290]_ , \new_[5291]_ ,
    \new_[5292]_ , \new_[5293]_ , \new_[5294]_ , \new_[5295]_ ,
    \new_[5296]_ , \new_[5297]_ , \new_[5298]_ , \new_[5299]_ ,
    \new_[5300]_ , \new_[5301]_ , \new_[5302]_ , \new_[5303]_ ,
    \new_[5304]_ , \new_[5305]_ , \new_[5306]_ , \new_[5307]_ ,
    \new_[5308]_ , \new_[5309]_ , \new_[5310]_ , \new_[5311]_ ,
    \new_[5312]_ , \new_[5313]_ , \new_[5314]_ , n610, n615, n620, n625,
    n630, n635, n640, n645, n650, n655, n660, n665, n670, n675, n680, n685,
    n690, n695, n700, n705, n710, n715, n720, n725, n730, n735, n740, n745,
    n750, n755, n760, n765, n770, n775, n780, n785, n790, n795, n800, n805,
    n810, n815, n820, n825, n830, n835, n840, n845, n850, n855, n860, n865,
    n870, n875, n880, n885, n890, n895, n900, n905, n910, n915, n920, n925,
    n930, n935, n940, n945, n950, n955, n960, n965, n970, n975, n980, n985,
    n990, n995, n1000, n1005, n1010, n1015, n1020, n1025, n1030, n1035,
    n1040, n1045, n1050, n1055, n1060, n1065, n1070, n1075, n1080, n1085,
    n1090, n1095, n1100, n1105, n1110, n1115, n1120, n1125, n1130, n1135,
    n1140, n1145, n1150, n1155, n1160, n1165, n1170, n1175, n1180, n1185,
    n1190, n1195, n1200, n1205, n1210, n1215, n1220, n1225, n1230, n1235,
    n1240, n1245;
  assign \new_[434]_  = \\FP_R_reg[25] ;
  assign \new_[435]_  = \\R_reg[25] ;
  assign \new_[436]_  = \\FP_R_reg[11] ;
  assign \new_[437]_  = \\R_reg[11] ;
  assign \new_[438]_  = \\FP_R_reg[3] ;
  assign \new_[439]_  = \\R_reg[7] ;
  assign \new_[440]_  = \\FP_R_reg[7] ;
  assign \new_[441]_  = \\R_reg[3] ;
  assign \new_[442]_  = \\FP_R_reg[15] ;
  assign \new_[443]_  = \\R_reg[15] ;
  assign \new_[444]_  = \\FP_R_reg[4] ;
  assign \new_[445]_  = \\R_reg[4] ;
  assign \new_[446]_  = \\FP_R_reg[29] ;
  assign \new_[447]_  = \\R_reg[29] ;
  assign \new_[448]_  = \\FP_R_reg[22] ;
  assign \new_[449]_  = \\R_reg[22] ;
  assign \new_[450]_  = \\R_reg[14] ;
  assign \new_[451]_  = \\R_reg[2] ;
  assign \new_[452]_  = \\FP_R_reg[5] ;
  assign \new_[453]_  = \\R_reg[5] ;
  assign \new_[454]_  = \\FP_R_reg[28] ;
  assign \new_[455]_  = \\FP_R_reg[14] ;
  assign \new_[456]_  = \\FP_R_reg[2] ;
  assign \new_[457]_  = \\R_reg[13] ;
  assign \new_[458]_  = \\R_reg[28] ;
  assign \new_[459]_  = \\FP_R_reg[13] ;
  assign n640 = ~\new_[514]_  | ~\new_[499]_ ;
  assign n645 = ~\new_[500]_  | ~\new_[516]_ ;
  assign n655 = ~\new_[507]_  | ~\new_[497]_ ;
  assign \new_[463]_  = \\FP_R_reg[31] ;
  assign \new_[464]_  = \\R_reg[26] ;
  assign \new_[465]_  = \\FP_R_reg[8] ;
  assign \new_[466]_  = \\FP_R_reg[20] ;
  assign \new_[467]_  = \\R_reg[31] ;
  assign \new_[468]_  = \\R_reg[20] ;
  assign \new_[469]_  = \\R_reg[8] ;
  assign \new_[470]_  = \\FP_R_reg[12] ;
  assign \new_[471]_  = \\R_reg[12] ;
  assign \new_[472]_  = \\FP_R_reg[26] ;
  assign \new_[473]_  = \\FP_R_reg[27] ;
  assign \new_[474]_  = \\FP_R_reg[19] ;
  assign \new_[475]_  = \\FP_R_reg[10] ;
  assign \new_[476]_  = \\FP_R_reg[21] ;
  assign \new_[477]_  = \\FP_R_reg[6] ;
  assign \new_[478]_  = \\R_reg[10] ;
  assign \new_[479]_  = \\R_reg[19] ;
  assign \new_[480]_  = \\R_reg[21] ;
  assign \new_[481]_  = \\R_reg[27] ;
  assign \new_[482]_  = \\R_reg[6] ;
  assign \new_[483]_  = \\FP_R_reg[9] ;
  assign \new_[484]_  = \\R_reg[9] ;
  assign \new_[485]_  = ~\\FP_R_reg[18] ;
  assign \new_[486]_  = \\R_reg[18] ;
  assign n730 = ~\new_[515]_  | ~\new_[509]_ ;
  assign n685 = ~\new_[518]_  | ~\new_[510]_ ;
  assign \new_[489]_  = ~\\FP_R_reg[30] ;
  assign \new_[490]_  = \\FP_R_reg[32] ;
  assign \new_[491]_  = \\R_reg[32] ;
  assign \new_[492]_  = \\FP_R_reg[23] ;
  assign \new_[493]_  = \\R_reg[23] ;
  assign \new_[494]_  = \\FP_R_reg[1] ;
  assign \new_[495]_  = \\R_reg[1] ;
  assign \new_[496]_  = \\R_reg[30] ;
  assign \new_[497]_  = ~\new_[513]_  | ~\new_[1695]_ ;
  assign n815 = ~\new_[522]_  | ~\new_[517]_ ;
  assign \new_[499]_  = ~\new_[5020]_  | ~\new_[1714]_ ;
  assign \new_[500]_  = ~\new_[4575]_  | ~\new_[1693]_ ;
  assign \new_[501]_  = ~\\FP_R_reg[17] ;
  assign \new_[502]_  = \\R_reg[17] ;
  assign \new_[503]_  = \\FP_R_reg[24] ;
  assign \new_[504]_  = \\R_reg[24] ;
  assign \new_[505]_  = \\FP_R_reg[16] ;
  assign \new_[506]_  = \\R_reg[16] ;
  assign \new_[507]_  = ~\new_[521]_  | ~\new_[1674]_ ;
  assign \new_[508]_  = ~\new_[520]_  | ~\new_[1696]_ ;
  assign \new_[509]_  = ~\new_[519]_  | ~\new_[1692]_ ;
  assign \new_[510]_  = ~\new_[524]_  | ~\new_[1713]_ ;
  assign \new_[511]_  = ~\new_[4524]_  | ~\new_[1710]_ ;
  assign n925 = ~\new_[526]_  | ~\new_[528]_ ;
  assign \new_[513]_  = ~\new_[521]_ ;
  assign \new_[514]_  = \new_[5027]_  | \new_[5028]_  | \new_[1714]_  | \new_[5022]_ ;
  assign \new_[515]_  = ~\new_[4560]_  | ~\new_[1673]_ ;
  assign \new_[516]_  = \new_[4582]_  | \new_[589]_  | \new_[1693]_  | \new_[4580]_ ;
  assign \new_[517]_  = ~\new_[525]_  | ~\new_[1728]_ ;
  assign \new_[518]_  = ~\new_[4531]_  | ~\new_[1698]_ ;
  assign \new_[519]_  = ~\new_[4560]_ ;
  assign \new_[520]_  = ~\new_[4524]_ ;
  assign \new_[521]_  = ~\new_[624]_  | ~\new_[540]_  | ~\new_[538]_  | ~\new_[603]_ ;
  assign \new_[522]_  = ~\new_[4774]_  | ~\new_[1709]_ ;
  assign \new_[523]_  = ~\new_[4989]_  | ~\new_[1694]_ ;
  assign \new_[524]_  = ~\new_[4531]_ ;
  assign \new_[525]_  = ~\new_[4774]_ ;
  assign \new_[526]_  = ~\new_[4845]_  | ~\new_[1697]_ ;
  assign \new_[527]_  = ~\new_[1177]_  | (~\new_[550]_  & ~\new_[732]_ );
  assign \new_[528]_  = ~\new_[4852]_  | ~\new_[4851]_  | ~\new_[1712]_  | ~\new_[4846]_ ;
  assign \new_[529]_  = ~\new_[539]_  | ~\new_[607]_ ;
  assign \new_[530]_  = (~\new_[4873]_  | ~\new_[562]_ ) & (~\new_[672]_  | ~\new_[5189]_ );
  assign \new_[531]_  = ~\new_[546]_  & (~\new_[578]_  | ~\new_[4782]_ );
  assign \new_[532]_  = ~\new_[549]_  | ~\new_[1318]_ ;
  assign \new_[533]_  = ~\new_[542]_  | ~\new_[1177]_ ;
  assign \new_[534]_  = (~\new_[4874]_  | ~\new_[558]_ ) & (~\new_[800]_  | ~\new_[5190]_ );
  assign \new_[535]_  = ~\new_[1308]_  | (~\new_[577]_  & ~\new_[997]_ );
  assign \new_[536]_  = ~\new_[583]_  & (~\new_[575]_  | ~\new_[1523]_ );
  assign \new_[537]_  = ~\new_[756]_  & ~\new_[561]_ ;
  assign \new_[538]_  = ~\new_[552]_  | ~\new_[1524]_ ;
  assign \new_[539]_  = ~\new_[4873]_  | (~\new_[573]_  & ~\new_[960]_ );
  assign \new_[540]_  = ~\new_[854]_  & ~\new_[551]_ ;
  assign \new_[541]_  = ~\new_[5149]_  | ~\new_[4535]_ ;
  assign \new_[542]_  = ~\new_[617]_  | (~\new_[598]_  & ~\new_[5004]_ );
  assign \new_[543]_  = ~\new_[553]_ ;
  assign \new_[544]_  = ~\new_[609]_  | ~\new_[615]_  | ~\new_[655]_  | ~\new_[599]_ ;
  assign \new_[545]_  = (~\new_[600]_  | ~\new_[1318]_ ) & (~\new_[1133]_  | ~\new_[696]_ );
  assign \new_[546]_  = ~\new_[675]_  | ~\new_[625]_  | ~\new_[618]_  | ~\new_[679]_ ;
  assign \new_[547]_  = ~\new_[568]_  | ~\new_[1319]_ ;
  assign \new_[548]_  = ~\new_[993]_  & ~\new_[570]_ ;
  assign \new_[549]_  = ~\new_[720]_  | ~\new_[593]_  | ~\new_[799]_ ;
  assign \new_[550]_  = ~\new_[620]_  | ~\new_[846]_  | ~\new_[649]_  | ~\new_[1033]_ ;
  assign \new_[551]_  = ~\new_[1524]_  & (~\new_[753]_  | ~\new_[4753]_ );
  assign \new_[552]_  = ~\new_[932]_  | ~\new_[1167]_  | ~\new_[666]_  | ~\new_[971]_ ;
  assign \new_[553]_  = ~\new_[627]_  | ~\new_[661]_  | ~\new_[900]_ ;
  assign \new_[554]_  = ~\new_[821]_  & ~\new_[590]_ ;
  assign \new_[555]_  = ~\new_[595]_  | ~\new_[5126]_ ;
  assign \new_[556]_  = ~\new_[596]_  | ~\new_[1178]_ ;
  assign \new_[557]_  = ~\new_[5121]_  | (~\new_[601]_  & ~\new_[885]_ );
  assign \new_[558]_  = ~\new_[832]_  | ~\new_[638]_  | ~\new_[622]_  | ~\new_[941]_ ;
  assign \new_[559]_  = ~\new_[822]_  | ~\new_[702]_  | ~\new_[635]_  | ~\new_[1049]_ ;
  assign \new_[560]_  = ~\new_[4462]_  | (~\new_[608]_  & ~\new_[904]_ );
  assign \new_[561]_  = ~\new_[1523]_  & (~\new_[882]_  | ~\new_[612]_ );
  assign \new_[562]_  = ~\new_[835]_  | ~\new_[652]_  | ~\new_[639]_  | ~\new_[726]_ ;
  assign \new_[563]_  = ~\new_[616]_  | ~\new_[613]_ ;
  assign \new_[564]_  = ~\new_[646]_  | ~\new_[752]_  | ~\new_[692]_ ;
  assign \new_[565]_  = ~\new_[614]_  & (~\new_[1087]_  | ~\new_[5039]_ );
  assign \new_[566]_  = ~\new_[605]_  | ~\new_[4975]_ ;
  assign \new_[567]_  = ~\new_[650]_  | ~\new_[657]_  | ~\new_[648]_ ;
  assign \new_[568]_  = ~\new_[884]_  | ~\new_[712]_  | ~\new_[761]_  | ~\new_[751]_ ;
  assign \new_[569]_  = ~\new_[768]_  | ~\new_[804]_  | ~\new_[602]_  | ~\new_[689]_ ;
  assign \new_[570]_  = ~\new_[4453]_  & (~\new_[660]_  | ~\new_[663]_ );
  assign \new_[571]_  = ~\new_[746]_  & ~\new_[606]_ ;
  assign \new_[572]_  = ~\new_[737]_  | ~\new_[668]_  | ~\new_[845]_ ;
  assign \new_[573]_  = ~\new_[1024]_  | ~\new_[619]_  | ~\new_[671]_ ;
  assign \new_[574]_  = ~\new_[658]_  | ~\new_[636]_  | ~\new_[893]_ ;
  assign \new_[575]_  = ~\new_[936]_  | ~\new_[986]_  | ~\new_[786]_  | ~\new_[710]_ ;
  assign \new_[576]_  = ~\new_[820]_  | ~\new_[797]_  | ~\new_[641]_ ;
  assign \new_[577]_  = ~\new_[1211]_  | ~\new_[834]_  | ~\new_[697]_  | ~\new_[1096]_ ;
  assign \new_[578]_  = ~\new_[977]_  | ~\new_[711]_  | ~\new_[688]_  | ~\new_[1182]_ ;
  assign \new_[579]_  = ~\new_[952]_  | ~\new_[805]_  | ~\new_[707]_  | ~\new_[731]_ ;
  assign \new_[580]_  = ~\new_[747]_  | ~\new_[631]_  | ~\new_[659]_ ;
  assign \new_[581]_  = ~\new_[811]_  | ~\new_[764]_  | ~\new_[623]_  | ~\new_[892]_ ;
  assign \new_[582]_  = ~\new_[695]_  | ~\new_[723]_  | ~\new_[1184]_ ;
  assign \new_[583]_  = ~\new_[1310]_  & (~\new_[701]_  | ~\new_[828]_ );
  assign \new_[584]_  = ~\new_[841]_  | ~\new_[670]_  | ~\new_[792]_ ;
  assign \new_[585]_  = ~\new_[644]_  & ~\new_[721]_ ;
  assign \new_[586]_  = ~\new_[766]_  | ~\new_[762]_  | ~\new_[735]_ ;
  assign \new_[587]_  = ~\new_[833]_  | ~\new_[653]_ ;
  assign \new_[588]_  = ~\new_[1317]_  & (~\new_[713]_  | ~\new_[5199]_ );
  assign \new_[589]_  = ~\new_[4581]_ ;
  assign \new_[590]_  = ~\new_[4880]_  | ~\new_[734]_  | ~\new_[859]_ ;
  assign \new_[591]_  = ~\new_[654]_  | ~\new_[716]_ ;
  assign \new_[592]_  = ~\new_[717]_  | ~\new_[839]_  | ~\new_[840]_ ;
  assign \new_[593]_  = ~\new_[1067]_  & ~\new_[642]_ ;
  assign \new_[594]_  = ~\new_[632]_  | ~\new_[5004]_ ;
  assign \new_[595]_  = ~\new_[4603]_  | ~\new_[690]_  | ~\new_[694]_ ;
  assign \new_[596]_  = ~\new_[634]_  | ~\new_[803]_ ;
  assign \new_[597]_  = ~\new_[1075]_  | (~\new_[693]_  & ~\new_[5209]_ );
  assign \new_[598]_  = ~\new_[948]_  & ~\new_[633]_ ;
  assign \new_[599]_  = ~\new_[640]_  | ~\new_[4417]_ ;
  assign \new_[600]_  = ~\new_[637]_  | ~\new_[1042]_ ;
  assign \new_[601]_  = ~\new_[741]_  | ~\new_[677]_ ;
  assign \new_[602]_  = ~\new_[1280]_  | ~\new_[685]_ ;
  assign \new_[603]_  = ~\new_[1310]_  | (~\new_[788]_  & ~\new_[975]_ );
  assign \new_[604]_  = ~\new_[787]_  & ~\new_[672]_ ;
  assign \new_[605]_  = ~\new_[703]_  | ~\new_[1037]_ ;
  assign \new_[606]_  = ~\new_[1187]_  | ~\new_[1034]_  | ~\new_[857]_  | ~\new_[1181]_ ;
  assign \new_[607]_  = ~\new_[5190]_  | (~\new_[774]_  & ~\new_[916]_ );
  assign \new_[608]_  = ~\new_[1061]_  | ~\new_[827]_  | ~\new_[1079]_  | ~\new_[1253]_ ;
  assign \new_[609]_  = ~\new_[699]_  | ~\new_[4417]_ ;
  assign \new_[610]_  = ~\new_[860]_  | (~\new_[809]_  & ~\new_[4961]_ );
  assign \new_[611]_  = ~\new_[719]_  | ~\new_[698]_ ;
  assign \new_[612]_  = ~\new_[1036]_  & (~\new_[795]_  | ~\new_[1172]_ );
  assign \new_[613]_  = ~\new_[1014]_  & ~\new_[708]_ ;
  assign \new_[614]_  = ~\new_[4961]_  & (~\new_[790]_  | ~\new_[1127]_ );
  assign \new_[615]_  = ~\new_[1179]_  | ~\new_[755]_  | ~\new_[4417]_ ;
  assign \new_[616]_  = ~\new_[1020]_  & ~\new_[673]_ ;
  assign \new_[617]_  = ~\new_[733]_  | ~\new_[5000]_ ;
  assign \new_[618]_  = ~\new_[4894]_  | (~\new_[742]_  & ~\new_[963]_ );
  assign \new_[619]_  = ~\new_[728]_  | ~\new_[5046]_ ;
  assign \new_[620]_  = ~\new_[727]_  | ~\new_[4999]_ ;
  assign \new_[621]_  = ~\new_[850]_  & ~\new_[718]_ ;
  assign \new_[622]_  = ~\new_[5046]_  | (~\new_[779]_  & ~\new_[5292]_ );
  assign \new_[623]_  = ~\new_[714]_  | ~\new_[4390]_ ;
  assign \new_[624]_  = ~\new_[725]_  | ~\new_[1172]_ ;
  assign \new_[625]_  = ~\new_[680]_  & (~\new_[968]_  | ~\new_[1508]_ );
  assign \new_[626]_  = ~\new_[1520]_  & (~\new_[789]_  | ~\new_[1149]_ );
  assign \new_[627]_  = ~\new_[681]_  & ~\new_[928]_ ;
  assign \new_[628]_  = ~\new_[682]_  | ~\new_[1521]_ ;
  assign \new_[629]_  = ~\new_[678]_  | ~\new_[5082]_ ;
  assign \new_[630]_  = ~\new_[760]_  | ~\new_[1176]_ ;
  assign \new_[631]_  = ~\new_[771]_  | ~\new_[5046]_ ;
  assign \new_[632]_  = ~\new_[996]_  | ~\new_[763]_ ;
  assign \new_[633]_  = ~\new_[1043]_  | ~\new_[748]_ ;
  assign \new_[634]_  = ~\new_[1018]_  & ~\new_[782]_ ;
  assign \new_[635]_  = ~\new_[1405]_  | (~\new_[912]_  & ~\new_[1333]_ );
  assign \new_[636]_  = ~\new_[4389]_  | (~\new_[918]_  & ~\new_[1366]_ );
  assign \new_[637]_  = ~\new_[1404]_  | (~\new_[815]_  & ~\new_[945]_ );
  assign \new_[638]_  = ~\new_[5191]_  | (~\new_[913]_  & ~\new_[923]_ );
  assign \new_[639]_  = ~\new_[1023]_  & (~\new_[813]_  | ~\new_[1039]_ );
  assign \new_[640]_  = ~\new_[784]_  | ~\new_[1077]_ ;
  assign \new_[641]_  = ~\new_[739]_  & ~\new_[781]_ ;
  assign \new_[642]_  = ~\new_[1033]_  | (~\new_[819]_  & ~\new_[1405]_ );
  assign \new_[643]_  = ~\new_[780]_  | (~\new_[1422]_  & ~\new_[1259]_ );
  assign \new_[644]_  = ~\new_[791]_  | ~\new_[1013]_ ;
  assign \new_[645]_  = ~\new_[749]_  | ~\new_[1013]_ ;
  assign \new_[646]_  = ~\new_[1520]_  | (~\new_[826]_  & ~\new_[1295]_ );
  assign \new_[647]_  = ~\new_[1029]_  & (~\new_[829]_  | ~\new_[914]_ );
  assign \new_[648]_  = ~\new_[818]_  & ~\new_[807]_ ;
  assign \new_[649]_  = ~\new_[806]_  | ~\new_[1404]_ ;
  assign \new_[650]_  = ~\new_[808]_  & ~\new_[940]_ ;
  assign \new_[651]_  = ~\new_[810]_  | ~\new_[4975]_ ;
  assign \new_[652]_  = ~\new_[5046]_  | (~\new_[955]_  & ~\new_[874]_ );
  assign \new_[653]_  = ~\new_[4388]_  | (~\new_[843]_  & ~\new_[1462]_ );
  assign \new_[654]_  = ~\new_[4390]_  | (~\new_[969]_  & ~\new_[838]_ );
  assign \new_[655]_  = ~\new_[1179]_  | (~\new_[877]_  & ~\new_[983]_ );
  assign \new_[656]_  = ~\new_[1427]_  | (~\new_[875]_  & ~\new_[1002]_ );
  assign \new_[657]_  = ~\new_[796]_  & ~\new_[930]_ ;
  assign \new_[658]_  = ~\new_[4391]_  | (~\new_[867]_  & ~\new_[1449]_ );
  assign \new_[659]_  = ~\new_[5189]_  | (~\new_[872]_  & ~\new_[1452]_ );
  assign \new_[660]_  = ~\new_[998]_  & (~\new_[863]_  | ~\new_[5284]_ );
  assign \new_[661]_  = ~\new_[1417]_  | (~\new_[873]_  & ~\new_[1063]_ );
  assign \new_[662]_  = ~\new_[994]_  | (~\new_[866]_  & ~\new_[5000]_ );
  assign \new_[663]_  = (~\new_[878]_  | ~\new_[5286]_ ) & (~\new_[1522]_  | ~\new_[1445]_ );
  assign \new_[664]_  = ~\new_[1198]_  | ~\new_[1021]_  | ~\new_[898]_ ;
  assign \new_[665]_  = ~\new_[964]_  | ~\new_[783]_ ;
  assign \new_[666]_  = ~\new_[724]_ ;
  assign \new_[667]_  = ~\new_[1521]_  & (~\new_[880]_  | ~\new_[1075]_ );
  assign \new_[668]_  = ~\new_[777]_  | ~\new_[4388]_ ;
  assign \new_[669]_  = ~\new_[847]_  | ~\new_[763]_ ;
  assign \new_[670]_  = ~\new_[744]_  | ~\new_[1404]_ ;
  assign \new_[671]_  = ~\new_[765]_  | ~\new_[1518]_ ;
  assign \new_[672]_  = ~\new_[842]_  | ~\new_[836]_ ;
  assign \new_[673]_  = ~\new_[973]_  | (~\new_[4565]_  & ~\new_[5082]_ );
  assign \new_[674]_  = ~\new_[1071]_  & ~\new_[816]_ ;
  assign \new_[675]_  = ~\new_[1292]_  | ~\new_[897]_ ;
  assign \new_[676]_  = ~\new_[902]_  | ~\new_[1438]_ ;
  assign \new_[677]_  = ~\new_[901]_  | ~\new_[5083]_ ;
  assign \new_[678]_  = ~\new_[891]_  | ~\new_[1152]_ ;
  assign \new_[679]_  = ~\new_[1417]_  | ~\new_[1093]_ ;
  assign \new_[680]_  = ~\new_[1571]_  & ~\new_[881]_ ;
  assign \new_[681]_  = ~\new_[1017]_  & ~\new_[1572]_  & ~\new_[1176]_ ;
  assign \new_[682]_  = ~\new_[906]_  | ~\new_[1234]_ ;
  assign \new_[683]_  = ~\new_[896]_  | ~\new_[1515]_ ;
  assign \new_[684]_  = ~\new_[924]_  & ~\new_[889]_ ;
  assign \new_[685]_  = ~\new_[915]_  | ~\new_[5115]_ ;
  assign \new_[686]_  = ~\new_[758]_ ;
  assign \new_[687]_  = ~\new_[899]_  | ~\new_[5083]_ ;
  assign \new_[688]_  = \new_[887]_  & \new_[1202]_ ;
  assign \new_[689]_  = ~\new_[1274]_  | ~\new_[5191]_  | ~\new_[1022]_ ;
  assign \new_[690]_  = ~\new_[903]_  & ~\new_[1158]_ ;
  assign \new_[691]_  = ~\new_[879]_  | ~\new_[4461]_ ;
  assign \new_[692]_  = ~\new_[776]_ ;
  assign \new_[693]_  = ~\new_[978]_  & ~\new_[888]_ ;
  assign \new_[694]_  = ~\new_[886]_  & (~\new_[1428]_  | ~\new_[1269]_ );
  assign \new_[695]_  = ~\new_[1508]_  | (~\new_[931]_  & ~\new_[1136]_ );
  assign \new_[696]_  = ~\new_[1055]_  | ~\new_[1122]_  | ~\new_[991]_ ;
  assign \new_[697]_  = ~\new_[1098]_  & (~\new_[947]_  | ~\new_[4391]_ );
  assign \new_[698]_  = ~\new_[956]_  & (~\new_[942]_  | ~\new_[5046]_ );
  assign \new_[699]_  = ~\new_[1124]_  | ~\new_[934]_  | ~\new_[935]_ ;
  assign \new_[700]_  = ~\new_[4390]_  | (~\new_[957]_  & ~\new_[1453]_ );
  assign \new_[701]_  = ~\new_[937]_  & ~\new_[907]_ ;
  assign \new_[702]_  = ~\new_[910]_  | ~\new_[1306]_ ;
  assign \new_[703]_  = ~\new_[1171]_  | (~\new_[962]_  & ~\new_[1068]_ );
  assign \new_[704]_  = ~\new_[783]_ ;
  assign \new_[705]_  = ~\new_[1044]_  | ~\new_[941]_  | ~\new_[4583]_ ;
  assign \new_[706]_  = ~\new_[1310]_  | (~\new_[929]_  & ~\new_[1150]_ );
  assign \new_[707]_  = ~\new_[5191]_  | (~\new_[944]_  & ~\new_[1120]_ );
  assign \new_[708]_  = ~\new_[5083]_  & (~\new_[967]_  | ~\new_[1364]_ );
  assign \new_[709]_  = ~\new_[917]_  | ~\new_[4757]_ ;
  assign \new_[710]_  = ~\new_[909]_  | ~\new_[1172]_ ;
  assign \new_[711]_  = ~\new_[1073]_  & ~\new_[908]_ ;
  assign \new_[712]_  = ~\new_[862]_  | ~\new_[1417]_ ;
  assign \new_[713]_  = ~\new_[983]_  & (~\new_[988]_  | ~\new_[1521]_ );
  assign \new_[714]_  = ~\new_[869]_  | ~\new_[1369]_ ;
  assign \new_[715]_  = ~\new_[868]_  | ~\new_[5154]_ ;
  assign \new_[716]_  = ~\new_[868]_  | ~\new_[4388]_ ;
  assign \new_[717]_  = ~\new_[870]_  | ~\new_[4388]_ ;
  assign \new_[718]_  = ~\new_[1189]_  | ~\new_[1066]_  | ~\new_[1182]_  | ~\new_[1065]_ ;
  assign \new_[719]_  = ~\new_[950]_  & ~\new_[5197]_ ;
  assign \new_[720]_  = ~\new_[858]_  & ~\new_[927]_ ;
  assign \new_[721]_  = ~\new_[4999]_  & ~\new_[846]_ ;
  assign \new_[722]_  = ~\new_[828]_  | ~\new_[1167]_ ;
  assign \new_[723]_  = ~\new_[873]_  & ~\new_[853]_ ;
  assign \new_[724]_  = ~\new_[825]_  | ~\new_[1051]_ ;
  assign \new_[725]_  = ~\new_[933]_  | ~\new_[4806]_ ;
  assign \new_[726]_  = ~\new_[794]_ ;
  assign \new_[727]_  = ~\new_[871]_  | ~\new_[1215]_ ;
  assign \new_[728]_  = ~\new_[1328]_  | ~\new_[876]_  | ~\new_[1373]_ ;
  assign \new_[729]_  = ~\new_[1041]_  & (~\new_[989]_  | ~\new_[1083]_ );
  assign \new_[730]_  = ~\new_[837]_  | ~\new_[1217]_ ;
  assign \new_[731]_  = ~\new_[861]_  & ~\new_[919]_ ;
  assign \new_[732]_  = ~\new_[1047]_  | ~\new_[1048]_ ;
  assign \new_[733]_  = ~\new_[852]_  | ~\new_[1049]_ ;
  assign \new_[734]_  = ~\new_[824]_  | ~\new_[5083]_ ;
  assign \new_[735]_  = ~\new_[1041]_  | (~\new_[987]_  & ~\new_[1251]_ );
  assign \new_[736]_  = ~\new_[1080]_  & (~\new_[1010]_  | ~\new_[1041]_ );
  assign \new_[737]_  = ~\new_[814]_ ;
  assign \new_[738]_  = ~\new_[1147]_  | (~\new_[1131]_  & ~\new_[1520]_ );
  assign \new_[739]_  = ~\new_[1232]_  & ~\new_[4999]_ ;
  assign \new_[740]_  = ~\new_[1003]_  | ~\new_[1423]_ ;
  assign \new_[741]_  = ~\new_[1008]_  | ~\new_[1423]_ ;
  assign \new_[742]_  = ~\new_[1435]_  | ~\new_[1201]_ ;
  assign \new_[743]_  = ~\new_[922]_  & ~\new_[990]_ ;
  assign \new_[744]_  = ~\new_[1007]_  | ~\new_[1204]_ ;
  assign \new_[745]_  = \new_[972]_  | \new_[4398]_ ;
  assign \new_[746]_  = ~\new_[1201]_  | ~\new_[1186]_ ;
  assign \new_[747]_  = ~\new_[1006]_  | ~\new_[1040]_ ;
  assign \new_[748]_  = ~\new_[1005]_  | ~\new_[1412]_ ;
  assign \new_[749]_  = ~\new_[1016]_  | ~\new_[1109]_ ;
  assign \new_[750]_  = ~\new_[1134]_  | ~\new_[1510]_  | ~\new_[1171]_ ;
  assign \new_[751]_  = ~\new_[1004]_  | ~\new_[1506]_ ;
  assign \new_[752]_  = ~\new_[1254]_  & ~\new_[980]_ ;
  assign \new_[753]_  = ~\new_[1418]_  | ~\new_[979]_ ;
  assign \new_[754]_  = \new_[1077]_  & \new_[1012]_ ;
  assign \new_[755]_  = ~\new_[1149]_  | ~\new_[1059]_  | ~\new_[1257]_ ;
  assign \new_[756]_  = ~\new_[1286]_  & ~\new_[4975]_  & ~\new_[1137]_ ;
  assign \new_[757]_  = ~\new_[1321]_  & ~\new_[1350]_  & ~\new_[5284]_ ;
  assign \new_[758]_  = ~\new_[986]_  & ~\new_[1172]_ ;
  assign \new_[759]_  = ~\new_[1021]_  | ~\new_[4603]_ ;
  assign \new_[760]_  = ~\new_[1185]_  | ~\new_[1094]_ ;
  assign \new_[761]_  = \new_[1187]_  & \new_[1201]_ ;
  assign \new_[762]_  = ~\new_[1076]_  & ~\new_[981]_ ;
  assign \new_[763]_  = ~\new_[1410]_  | ~\new_[4398]_  | ~\new_[1175]_  | ~\new_[1415]_ ;
  assign \new_[764]_  = ~\new_[831]_ ;
  assign \new_[765]_  = ~\new_[1025]_  | ~\new_[1326]_ ;
  assign \new_[766]_  = ~\new_[1009]_  | ~\new_[5286]_ ;
  assign \new_[767]_  = ~\new_[1287]_  & ~\new_[5053]_  & ~\new_[1039]_ ;
  assign \new_[768]_  = ~\new_[1022]_  | ~\new_[1121]_ ;
  assign \new_[769]_  = ~\new_[844]_ ;
  assign \new_[770]_  = ~\new_[1011]_  | ~\new_[5286]_ ;
  assign \new_[771]_  = ~\new_[1229]_  | ~\new_[1000]_ ;
  assign \new_[772]_  = ~\new_[853]_ ;
  assign \new_[773]_  = ~\new_[985]_  | ~\new_[1179]_ ;
  assign \new_[774]_  = ~\new_[1040]_  & ~\new_[1225]_ ;
  assign \new_[775]_  = ~\new_[984]_  & ~\new_[1062]_ ;
  assign \new_[776]_  = ~\new_[1145]_  | (~\new_[1143]_  & ~\new_[1616]_ );
  assign \new_[777]_  = ~\new_[1001]_  | ~\new_[1111]_ ;
  assign \new_[778]_  = ~\new_[861]_ ;
  assign \new_[779]_  = ~\new_[1025]_  | ~\new_[1104]_ ;
  assign \new_[780]_  = ~\new_[1515]_  | ~\new_[1015]_ ;
  assign \new_[781]_  = ~\new_[1050]_  | ~\new_[1048]_  | ~\new_[1074]_ ;
  assign \new_[782]_  = ~\new_[887]_ ;
  assign \new_[783]_  = ~\new_[1015]_  | ~\new_[1520]_ ;
  assign \new_[784]_  = ~\new_[1569]_  | ~\new_[1015]_ ;
  assign \new_[785]_  = ~\new_[1264]_  | ~\new_[5041]_ ;
  assign \new_[786]_  = (~\new_[1056]_  | ~\new_[1310]_ ) & (~\new_[1237]_  | ~\new_[1611]_ );
  assign \new_[787]_  = ~\new_[5189]_  & (~\new_[1326]_  | ~\new_[1044]_ );
  assign \new_[788]_  = ~\new_[1035]_  | ~\new_[925]_  | ~\new_[1167]_ ;
  assign \new_[789]_  = ~\new_[896]_ ;
  assign \new_[790]_  = ~\new_[4721]_  & (~\new_[1086]_  | ~\new_[5041]_ );
  assign \new_[791]_  = ~\new_[1329]_  | ~\new_[1316]_  | ~\new_[1306]_ ;
  assign \new_[792]_  = ~\new_[4999]_  | ~\new_[946]_ ;
  assign \new_[793]_  = ~\new_[926]_  & ~\new_[1036]_ ;
  assign \new_[794]_  = ~\new_[4583]_  | ~\new_[5196]_ ;
  assign \new_[795]_  = ~\new_[1324]_  | ~\new_[966]_  | ~\new_[1125]_ ;
  assign \new_[796]_  = ~\new_[921]_  | ~\new_[1031]_ ;
  assign \new_[797]_  = ~\new_[1205]_  & ~\new_[953]_ ;
  assign \new_[798]_  = ~\new_[945]_  | ~\new_[1412]_ ;
  assign \new_[799]_  = ~\new_[949]_  & ~\new_[954]_ ;
  assign \new_[800]_  = ~\new_[4583]_  | ~\new_[1054]_ ;
  assign \new_[801]_  = ~\new_[943]_  & ~\new_[995]_ ;
  assign \new_[802]_  = ~\new_[1119]_  | ~\new_[1039]_  | ~\new_[5046]_ ;
  assign \new_[803]_  = ~\new_[1506]_  | (~\new_[1126]_  & ~\new_[1242]_ );
  assign \new_[804]_  = ~\new_[1119]_  | ~\new_[1040]_  | ~\new_[1311]_ ;
  assign \new_[805]_  = ~\new_[916]_ ;
  assign \new_[806]_  = ~\new_[961]_  | ~\new_[1055]_ ;
  assign \new_[807]_  = ~\new_[1310]_  & (~\new_[1200]_  | ~\new_[1072]_ );
  assign \new_[808]_  = ~\new_[939]_  | ~\new_[938]_ ;
  assign \new_[809]_  = ~\new_[981]_  & (~\new_[1130]_  | ~\new_[5286]_ );
  assign \new_[810]_  = ~\new_[974]_  | ~\new_[1038]_ ;
  assign \new_[811]_  = ~\new_[992]_  & (~\new_[1128]_  | ~\new_[5161]_ );
  assign \new_[812]_  = ~\new_[920]_ ;
  assign \new_[813]_  = ~\new_[1045]_  | ~\new_[1046]_ ;
  assign \new_[814]_  = ~\new_[5161]_  & (~\new_[1209]_  | ~\new_[1290]_ );
  assign \new_[815]_  = ~\new_[1100]_  | (~\new_[1313]_  & ~\new_[1204]_ );
  assign \new_[816]_  = ~\new_[1508]_  & (~\new_[1248]_  | ~\new_[1243]_ );
  assign \new_[817]_  = ~\new_[1091]_  | ~\new_[1323]_ ;
  assign \new_[818]_  = ~\new_[1510]_  & ~\new_[1088]_ ;
  assign \new_[819]_  = ~\new_[1123]_  & ~\new_[1224]_ ;
  assign \new_[820]_  = ~\new_[927]_ ;
  assign \new_[821]_  = ~\new_[1129]_  & ~\new_[1428]_ ;
  assign \new_[822]_  = ~\new_[1281]_  | ~\new_[1175]_  | ~\new_[4999]_ ;
  assign \new_[823]_  = ~\new_[883]_  & ~\new_[1063]_ ;
  assign \new_[824]_  = ~\new_[1271]_  | ~\new_[1260]_  | ~\new_[1438]_ ;
  assign \new_[825]_  = ~\new_[1241]_  | ~\new_[1594]_  | ~\new_[1309]_ ;
  assign \new_[826]_  = ~\new_[1077]_  | ~\new_[1394]_ ;
  assign \new_[827]_  = ~\new_[1520]_  | (~\new_[1235]_  & ~\new_[1478]_ );
  assign \new_[828]_  = ~\new_[1431]_  | ~\new_[1309]_  | ~\new_[4802]_ ;
  assign \new_[829]_  = ~\new_[1090]_  & ~\new_[1153]_ ;
  assign \new_[830]_  = ~\new_[1171]_  & ~\new_[1088]_ ;
  assign \new_[831]_  = ~\new_[1216]_  | ~\new_[1103]_ ;
  assign \new_[832]_  = ~\new_[1493]_  | ~\new_[1492]_  | ~\new_[1039]_  | ~\new_[5053]_ ;
  assign \new_[833]_  = ~\new_[5153]_  | ~\new_[1430]_  | ~\new_[4391]_ ;
  assign \new_[834]_  = ~\new_[4390]_  | ~\new_[1108]_ ;
  assign \new_[835]_  = ~\new_[1039]_  | ~\new_[1206]_ ;
  assign \new_[836]_  = ~\new_[5116]_  | ~\new_[1097]_ ;
  assign \new_[837]_  = ~\new_[946]_ ;
  assign \new_[838]_  = ~\new_[1456]_  | ~\new_[1112]_ ;
  assign \new_[839]_  = ~\new_[5161]_  | ~\new_[1110]_ ;
  assign \new_[840]_  = ~\new_[1465]_  | ~\new_[4388]_  | ~\new_[1312]_ ;
  assign \new_[841]_  = ~\new_[1314]_  | ~\new_[1101]_ ;
  assign \new_[842]_  = ~\new_[5116]_  | ~\new_[1114]_ ;
  assign \new_[843]_  = ~\new_[1096]_  | ~\new_[1216]_ ;
  assign \new_[844]_  = ~\new_[1105]_  | ~\new_[1227]_ ;
  assign \new_[845]_  = ~\new_[951]_ ;
  assign \new_[846]_  = ~\new_[953]_ ;
  assign \new_[847]_  = ~\new_[1281]_  | ~\new_[1316]_  | ~\new_[5000]_ ;
  assign \new_[848]_  = ~\new_[1111]_  | ~\new_[1112]_ ;
  assign \new_[849]_  = ~\new_[4391]_  | ~\new_[1113]_ ;
  assign \new_[850]_  = ~\new_[1563]_  & (~\new_[1240]_  | ~\new_[1398]_ );
  assign \new_[851]_  = ~\new_[1322]_  | ~\new_[1089]_ ;
  assign \new_[852]_  = ~\new_[1224]_  & ~\new_[1101]_ ;
  assign \new_[853]_  = ~\new_[1249]_  & ~\new_[1606]_  & ~\new_[1508]_ ;
  assign \new_[854]_  = ~\new_[1286]_  & ~\new_[1171]_  & ~\new_[1524]_ ;
  assign \new_[855]_  = ~\new_[1256]_  | ~\new_[1106]_  | ~\new_[1358]_ ;
  assign \new_[856]_  = ~\new_[5116]_  | ~\new_[1121]_ ;
  assign \new_[857]_  = ~\new_[1057]_  | ~\new_[1508]_ ;
  assign \new_[858]_  = ~\new_[1414]_  & ~\new_[1284]_  & ~\new_[1490]_ ;
  assign \new_[859]_  = ~\new_[1269]_  | ~\new_[1322]_  | ~\new_[5082]_ ;
  assign \new_[860]_  = ~\new_[1060]_  | ~\new_[1522]_ ;
  assign \new_[861]_  = ~\new_[1032]_  & ~\new_[5115]_ ;
  assign \new_[862]_  = ~\new_[1094]_  | (~\new_[1571]_  & ~\new_[1539]_ );
  assign \new_[863]_  = ~\new_[1084]_  | ~\new_[1350]_ ;
  assign \new_[864]_  = ~\new_[1140]_  | ~\new_[4603]_ ;
  assign \new_[865]_  = ~\new_[1070]_  | ~\new_[1199]_ ;
  assign \new_[866]_  = ~\new_[1205]_  & ~\new_[1154]_ ;
  assign \new_[867]_  = ~\new_[1099]_  | ~\new_[1456]_ ;
  assign \new_[868]_  = ~\new_[1367]_  | ~\new_[1095]_ ;
  assign \new_[869]_  = ~\new_[1375]_  & (~\new_[1622]_  | ~\new_[5153]_ );
  assign \new_[870]_  = ~\new_[1448]_  | ~\new_[1103]_ ;
  assign \new_[871]_  = ~\new_[1107]_  | ~\new_[1501]_ ;
  assign \new_[872]_  = ~\new_[1156]_  | ~\new_[1326]_ ;
  assign \new_[873]_  = ~\new_[1082]_  | ~\new_[1187]_ ;
  assign \new_[874]_  = ~\new_[1116]_  | ~\new_[1208]_ ;
  assign \new_[875]_  = ~\new_[1081]_  | ~\new_[1360]_ ;
  assign \new_[876]_  = ~\new_[1160]_  & (~\new_[5111]_  | ~\new_[1452]_ );
  assign \new_[877]_  = ~\new_[1058]_  | ~\new_[1288]_ ;
  assign \new_[878]_  = ~\new_[1381]_  | ~\new_[1085]_ ;
  assign \new_[879]_  = ~\new_[1422]_  | ~\new_[1352]_ ;
  assign \new_[880]_  = ~\new_[1421]_  | ~\new_[1146]_ ;
  assign \new_[881]_  = ~\new_[1343]_  | ~\new_[1508]_ ;
  assign \new_[882]_  = ~\new_[1150]_  | ~\new_[1310]_ ;
  assign \new_[883]_  = ~\new_[1185]_ ;
  assign \new_[884]_  = ~\new_[1607]_  | ~\new_[1138]_ ;
  assign \new_[885]_  = ~\new_[5079]_ ;
  assign \new_[886]_  = ~\new_[1516]_  & ~\new_[1139]_ ;
  assign \new_[887]_  = ~\new_[1571]_  | ~\new_[1138]_ ;
  assign \new_[888]_  = ~\new_[5291]_  | ~\new_[1132]_ ;
  assign \new_[889]_  = ~\new_[985]_ ;
  assign \new_[890]_  = ~\new_[1390]_  | ~\new_[1582]_  | ~\new_[1168]_ ;
  assign \new_[891]_  = ~\new_[990]_ ;
  assign \new_[892]_  = ~\new_[1584]_  | ~\new_[1159]_ ;
  assign \new_[893]_  = ~\new_[1526]_  | ~\new_[1159]_ ;
  assign \new_[894]_  = \new_[5116]_  | \new_[1287]_ ;
  assign \new_[895]_  = \new_[4956]_  & \new_[4725]_ ;
  assign \new_[896]_  = ~\new_[1566]_  & (~\new_[1300]_  | ~\new_[1166]_ );
  assign \new_[897]_  = ~\new_[1299]_  | ~\new_[1142]_ ;
  assign \new_[898]_  = ~\new_[1135]_  | ~\new_[5084]_ ;
  assign \new_[899]_  = ~\new_[1162]_  | ~\new_[1362]_ ;
  assign \new_[900]_  = ~\new_[1176]_  | ~\new_[4782]_  | ~\new_[1193]_ ;
  assign \new_[901]_  = ~\new_[1141]_  | ~\new_[1364]_ ;
  assign \new_[902]_  = ~\new_[1467]_  & (~\new_[1180]_  | ~\new_[1482]_ );
  assign \new_[903]_  = ~\new_[1247]_  | ~\new_[4642]_ ;
  assign \new_[904]_  = ~\new_[1353]_  | ~\new_[1148]_ ;
  assign \new_[905]_  = ~\new_[1012]_ ;
  assign \new_[906]_  = ~\new_[1015]_ ;
  assign \new_[907]_  = ~\new_[1167]_  | ~\new_[1035]_ ;
  assign \new_[908]_  = ~\new_[1176]_  & (~\new_[1191]_  | ~\new_[1250]_ );
  assign \new_[909]_  = ~\new_[1031]_  | ~\new_[4755]_ ;
  assign \new_[910]_  = ~\new_[1042]_  | ~\new_[1204]_ ;
  assign \new_[911]_  = ~\new_[1183]_  | ~\new_[1051]_ ;
  assign \new_[912]_  = ~\new_[1047]_  | ~\new_[1217]_ ;
  assign \new_[913]_  = ~\new_[1052]_  | ~\new_[1225]_ ;
  assign \new_[914]_  = ~\new_[1020]_ ;
  assign \new_[915]_  = ~\new_[1030]_  | ~\new_[1493]_ ;
  assign \new_[916]_  = ~\new_[1053]_  | ~\new_[1054]_ ;
  assign \new_[917]_  = ~\new_[1173]_  | ~\new_[1088]_ ;
  assign \new_[918]_  = ~\new_[1203]_  | (~\new_[1220]_  & ~\new_[1409]_ );
  assign \new_[919]_  = ~\new_[1025]_ ;
  assign \new_[920]_  = ~\new_[1203]_  | (~\new_[1430]_  & ~\new_[1223]_ );
  assign \new_[921]_  = ~\new_[4807]_  | ~\new_[1408]_  | ~\new_[1638]_ ;
  assign \new_[922]_  = ~\new_[4880]_ ;
  assign \new_[923]_  = ~\new_[1226]_  | (~\new_[5115]_  & ~\new_[1320]_ );
  assign \new_[924]_  = \new_[5201]_  | \new_[1179]_ ;
  assign \new_[925]_  = ~\new_[1418]_  | ~\new_[1190]_ ;
  assign \new_[926]_  = ~\new_[1031]_ ;
  assign \new_[927]_  = ~\new_[1490]_  & ~\new_[1218]_ ;
  assign \new_[928]_  = ~\new_[1034]_ ;
  assign \new_[929]_  = ~\new_[1200]_  | ~\new_[1323]_ ;
  assign \new_[930]_  = ~\new_[1035]_ ;
  assign \new_[931]_  = ~\new_[1201]_  | ~\new_[1243]_ ;
  assign \new_[932]_  = ~\new_[4757]_  | ~\new_[1325]_ ;
  assign \new_[933]_  = ~\new_[1036]_ ;
  assign \new_[934]_  = ~\new_[1391]_  | ~\new_[1616]_  | ~\new_[1570]_  | ~\new_[1521]_ ;
  assign \new_[935]_  = ~\new_[1566]_  | ~\new_[1400]_  | ~\new_[1570]_  | ~\new_[1521]_ ;
  assign \new_[936]_  = ~\new_[1510]_  | ~\new_[1195]_ ;
  assign \new_[937]_  = ~\new_[1037]_ ;
  assign \new_[938]_  = ~\new_[1437]_  | ~\new_[4803]_  | ~\new_[1310]_ ;
  assign \new_[939]_  = ~\new_[1431]_  | ~\new_[1418]_  | ~\new_[1310]_ ;
  assign \new_[940]_  = ~\new_[1038]_ ;
  assign \new_[941]_  = ~\new_[1206]_  | ~\new_[5116]_ ;
  assign \new_[942]_  = ~\new_[1208]_  | ~\new_[1207]_ ;
  assign \new_[943]_  = ~\new_[4389]_  & ~\new_[1586]_  & ~\new_[1372]_ ;
  assign \new_[944]_  = ~\new_[1228]_  | ~\new_[1326]_ ;
  assign \new_[945]_  = ~\new_[1221]_  | ~\new_[1210]_ ;
  assign \new_[946]_  = ~\new_[1230]_  | ~\new_[1215]_ ;
  assign \new_[947]_  = ~\new_[1278]_  | ~\new_[1213]_ ;
  assign \new_[948]_  = ~\new_[1219]_  & ~\new_[1315]_ ;
  assign \new_[949]_  = ~\new_[1315]_  & ~\new_[1217]_ ;
  assign \new_[950]_  = ~\new_[1046]_ ;
  assign \new_[951]_  = ~\new_[1213]_  | ~\new_[1216]_ ;
  assign \new_[952]_  = ~\new_[5046]_  | ~\new_[1214]_ ;
  assign \new_[953]_  = ~\new_[1411]_  & ~\new_[1218]_ ;
  assign \new_[954]_  = ~\new_[1047]_ ;
  assign \new_[955]_  = ~\new_[1229]_  | ~\new_[1225]_ ;
  assign \new_[956]_  = ~\new_[1052]_ ;
  assign \new_[957]_  = ~\new_[1285]_  | ~\new_[1222]_ ;
  assign \new_[958]_  = ~\new_[1357]_  | ~\new_[5285]_  | ~\new_[1396]_ ;
  assign \new_[959]_  = ~\new_[1233]_  | ~\new_[1197]_ ;
  assign \new_[960]_  = ~\new_[1053]_ ;
  assign \new_[961]_  = ~\new_[1335]_  & ~\new_[1231]_ ;
  assign \new_[962]_  = ~\new_[1236]_  | (~\new_[4802]_  & ~\new_[1439]_ );
  assign \new_[963]_  = ~\new_[1192]_  | ~\new_[1186]_ ;
  assign \new_[964]_  = ~\new_[1254]_  & (~\new_[5201]_  | ~\new_[1379]_ );
  assign \new_[965]_  = ~\new_[1357]_  | ~\new_[1612]_  | ~\new_[1619]_ ;
  assign \new_[966]_  = ~\new_[1196]_  | ~\new_[4802]_ ;
  assign \new_[967]_  = ~\new_[1245]_  & (~\new_[4604]_  | ~\new_[1363]_ );
  assign \new_[968]_  = ~\new_[1261]_  | ~\new_[1202]_ ;
  assign \new_[969]_  = ~\new_[1212]_  | ~\new_[1223]_ ;
  assign \new_[970]_  = ~\new_[1552]_  | ~\new_[1252]_ ;
  assign \new_[971]_  = ~\new_[4802]_  | ~\new_[1277]_ ;
  assign \new_[972]_  = ~\new_[1415]_  | ~\new_[1239]_ ;
  assign \new_[973]_  = ~\new_[1525]_  | ~\new_[1269]_ ;
  assign \new_[974]_  = ~\new_[1431]_  | ~\new_[1241]_ ;
  assign \new_[975]_  = ~\new_[1072]_ ;
  assign \new_[976]_  = ~\new_[5081]_  | ~\new_[1532]_ ;
  assign \new_[977]_  = ~\new_[1571]_  | ~\new_[1238]_ ;
  assign \new_[978]_  = ~\new_[1258]_  | ~\new_[1253]_ ;
  assign \new_[979]_  = ~\new_[1408]_  & ~\new_[1439]_ ;
  assign \new_[980]_  = ~\new_[1075]_ ;
  assign \new_[981]_  = ~\new_[5042]_  & ~\new_[1256]_ ;
  assign \new_[982]_  = ~\new_[1076]_ ;
  assign \new_[983]_  = ~\new_[1569]_  & ~\new_[1253]_ ;
  assign \new_[984]_  = ~\new_[1291]_  & ~\new_[1608]_  & ~\new_[1507]_ ;
  assign \new_[985]_  = ~\new_[1470]_  | ~\new_[1259]_ ;
  assign \new_[986]_  = ~\new_[1252]_  | ~\new_[1531]_ ;
  assign \new_[987]_  = ~\new_[1360]_  | ~\new_[4612]_ ;
  assign \new_[988]_  = ~\new_[1258]_  | ~\new_[5291]_ ;
  assign \new_[989]_  = ~\new_[1582]_  | ~\new_[1441]_ ;
  assign \new_[990]_  = ~\new_[4604]_  & ~\new_[1270]_ ;
  assign \new_[991]_  = ~\new_[1313]_  | ~\new_[1281]_ ;
  assign \new_[992]_  = ~\new_[1096]_ ;
  assign \new_[993]_  = ~\new_[5041]_  & ~\new_[1273]_ ;
  assign \new_[994]_  = ~\new_[1415]_  | ~\new_[4397]_  | ~\new_[1314]_ ;
  assign \new_[995]_  = ~\new_[1103]_ ;
  assign \new_[996]_  = ~\new_[1412]_  | ~\new_[1281]_ ;
  assign \new_[997]_  = ~\new_[1105]_ ;
  assign \new_[998]_  = ~\new_[1106]_ ;
  assign \new_[999]_  = ~\new_[1584]_  & ~\new_[1290]_ ;
  assign \new_[1000]_  = ~\new_[1120]_ ;
  assign \new_[1001]_  = ~\new_[1526]_  | ~\new_[1527]_  | ~\new_[1312]_ ;
  assign \new_[1002]_  = ~\new_[4612]_  | ~\new_[1263]_ ;
  assign \new_[1003]_  = ~\new_[1272]_  | ~\new_[1279]_ ;
  assign \new_[1004]_  = ~\new_[1246]_  | ~\new_[1249]_ ;
  assign \new_[1005]_  = ~\new_[1275]_  | ~\new_[1537]_ ;
  assign \new_[1006]_  = ~\new_[1283]_  | ~\new_[1373]_ ;
  assign \new_[1007]_  = ~\new_[1276]_  & ~\new_[1458]_ ;
  assign \new_[1008]_  = ~\new_[1129]_ ;
  assign \new_[1009]_  = ~\new_[1255]_  | ~\new_[1350]_ ;
  assign \new_[1010]_  = ~\new_[1262]_  | ~\new_[1354]_ ;
  assign \new_[1011]_  = ~\new_[1266]_  | ~\new_[1358]_ ;
  assign \new_[1012]_  = ~\new_[1302]_  | ~\new_[1383]_  | ~\new_[1521]_ ;
  assign \new_[1013]_  = ~\new_[1415]_  | ~\new_[1457]_  | ~\new_[1306]_  | ~\new_[1316]_ ;
  assign \new_[1014]_  = ~\new_[1420]_  & ~\new_[1164]_ ;
  assign \new_[1015]_  = ~\new_[1132]_ ;
  assign \new_[1016]_  = ~\new_[1412]_  & ~\new_[5000]_ ;
  assign \new_[1017]_  = ~\new_[1138]_ ;
  assign \new_[1018]_  = ~\new_[1142]_ ;
  assign \new_[1019]_  = ~\new_[5041]_  & ~\new_[1480]_ ;
  assign \new_[1020]_  = ~\new_[1403]_  & ~\new_[1481]_ ;
  assign \new_[1021]_  = ~\new_[4840]_  | ~\new_[1170]_ ;
  assign \new_[1022]_  = ~\new_[1155]_ ;
  assign \new_[1023]_  = ~\new_[4584]_  & ~\new_[1328]_  & ~\new_[5190]_ ;
  assign \new_[1024]_  = ~\new_[1169]_  | ~\new_[1553]_ ;
  assign \new_[1025]_  = ~\new_[1169]_  | ~\new_[1493]_ ;
  assign \new_[1026]_  = ~\new_[1174]_  & ~\new_[1551]_ ;
  assign \new_[1027]_  = \new_[5285]_  & \new_[4962]_ ;
  assign \new_[1028]_  = ~\new_[1164]_ ;
  assign \new_[1029]_  = ~\new_[1165]_ ;
  assign \new_[1030]_  = ~\new_[5110]_  & ~\new_[1425]_ ;
  assign \new_[1031]_  = ~\new_[1552]_  | ~\new_[1611]_  | ~\new_[1511]_  | ~\new_[1406]_ ;
  assign \new_[1032]_  = ~\new_[5110]_  | ~\new_[5192]_ ;
  assign \new_[1033]_  = ~\new_[1457]_  | ~\new_[1491]_  | ~\new_[1498]_ ;
  assign \new_[1034]_  = ~\new_[1609]_  | ~\new_[1466]_  | ~\new_[1571]_  | ~\new_[1506]_ ;
  assign \new_[1035]_  = ~\new_[1419]_  | ~\new_[1325]_ ;
  assign \new_[1036]_  = ~\new_[1323]_  & ~\new_[1418]_ ;
  assign \new_[1037]_  = ~\new_[1509]_  | ~\new_[4760]_ ;
  assign \new_[1038]_  = ~\new_[1310]_  | ~\new_[4857]_ ;
  assign \new_[1039]_  = ~\new_[5116]_ ;
  assign \new_[1040]_  = ~\new_[4584]_ ;
  assign \new_[1041]_  = ~\new_[5041]_ ;
  assign \new_[1042]_  = ~\new_[1412]_  | ~\new_[1331]_ ;
  assign \new_[1043]_  = ~\new_[1413]_  | ~\new_[1335]_ ;
  assign \new_[1044]_  = ~\new_[5110]_  | ~\new_[1327]_ ;
  assign \new_[1045]_  = ~\new_[1518]_  | ~\new_[1327]_ ;
  assign \new_[1046]_  = ~\new_[5191]_  | ~\new_[1334]_ ;
  assign \new_[1047]_  = ~\new_[1497]_  | ~\new_[1505]_  | ~\new_[1502]_  | ~\new_[4397]_ ;
  assign \new_[1048]_  = ~\new_[1411]_  | ~\new_[1329]_ ;
  assign \new_[1049]_  = ~\new_[1332]_  | ~\new_[1413]_ ;
  assign \new_[1050]_  = ~\new_[1411]_  | ~\new_[1335]_ ;
  assign \new_[1051]_  = ~\new_[1431]_  | ~\new_[1309]_  | ~\new_[1509]_ ;
  assign \new_[1052]_  = ~\new_[4795]_  | ~\new_[1553]_  | ~\new_[5110]_  | ~\new_[5049]_ ;
  assign \new_[1053]_  = ~\new_[1320]_  | ~\new_[4744]_ ;
  assign \new_[1054]_  = ~\new_[1320]_  | ~\new_[1327]_ ;
  assign \new_[1055]_  = ~\new_[1501]_  | ~\new_[1330]_ ;
  assign \new_[1056]_  = ~\new_[1337]_  | (~\new_[1419]_  & ~\new_[5282]_ );
  assign \new_[1057]_  = ~\new_[1435]_  | ~\new_[1344]_ ;
  assign \new_[1058]_  = ~\new_[1515]_  | ~\new_[1349]_ ;
  assign \new_[1059]_  = ~\new_[1351]_  | ~\new_[1570]_ ;
  assign \new_[1060]_  = ~\new_[4962]_  & ~\new_[1355]_ ;
  assign \new_[1061]_  = ~\new_[5211]_  | ~\new_[1379]_ ;
  assign \new_[1062]_  = ~\new_[1507]_  & ~\new_[1342]_ ;
  assign \new_[1063]_  = ~\new_[1188]_ ;
  assign \new_[1064]_  = ~\new_[1189]_ ;
  assign \new_[1065]_  = ~\new_[1563]_  | ~\new_[1345]_ ;
  assign \new_[1066]_  = ~\new_[1607]_  | ~\new_[1347]_ ;
  assign \new_[1067]_  = ~\new_[1497]_  & ~\new_[1339]_ ;
  assign \new_[1068]_  = ~\new_[1337]_  & ~\new_[1509]_ ;
  assign \new_[1069]_  = ~\new_[1362]_  | ~\new_[1472]_ ;
  assign \new_[1070]_  = ~\new_[1525]_  | ~\new_[1346]_ ;
  assign \new_[1071]_  = ~\new_[1571]_  & ~\new_[1338]_ ;
  assign \new_[1072]_  = ~\new_[1509]_  | ~\new_[1377]_ ;
  assign \new_[1073]_  = ~\new_[1572]_  & ~\new_[1341]_ ;
  assign \new_[1074]_  = ~\new_[1490]_  | ~\new_[1458]_ ;
  assign \new_[1075]_  = ~\new_[1569]_  | ~\new_[5200]_ ;
  assign \new_[1076]_  = ~\new_[1618]_  & ~\new_[1348]_ ;
  assign \new_[1077]_  = ~\new_[1395]_  | ~\new_[1514]_  | ~\new_[5211]_ ;
  assign \new_[1078]_  = ~\new_[1520]_  | ~\new_[1352]_ ;
  assign \new_[1079]_  = ~\new_[1351]_  | ~\new_[5211]_ ;
  assign \new_[1080]_  = ~\new_[1427]_  & ~\new_[1350]_ ;
  assign \new_[1081]_  = ~\new_[5041]_  | ~\new_[1442]_ ;
  assign \new_[1082]_  = ~\new_[1512]_  | ~\new_[1637]_  | ~\new_[1608]_  | ~\new_[1609]_ ;
  assign \new_[1083]_  = ~\new_[4613]_  | ~\new_[4624]_  | ~\new_[1612]_  | ~\new_[1643]_ ;
  assign \new_[1084]_  = ~\new_[1579]_  | ~\new_[1356]_ ;
  assign \new_[1085]_  = ~\new_[1612]_  | ~\new_[1356]_ ;
  assign \new_[1086]_  = ~\new_[1359]_  | ~\new_[1354]_ ;
  assign \new_[1087]_  = ~\new_[1294]_  | ~\new_[1355]_ ;
  assign \new_[1088]_  = ~\new_[1195]_ ;
  assign \new_[1089]_  = ~\new_[1362]_  | ~\new_[1361]_ ;
  assign \new_[1090]_  = ~\new_[1198]_ ;
  assign \new_[1091]_  = ~\new_[1564]_  | ~\new_[1594]_  | ~\new_[1406]_ ;
  assign \new_[1092]_  = ~\new_[1419]_  & ~\new_[1374]_ ;
  assign \new_[1093]_  = ~\new_[1201]_ ;
  assign \new_[1094]_  = ~\new_[1608]_  | ~\new_[1343]_ ;
  assign \new_[1095]_  = ~\new_[1585]_  | ~\new_[1366]_ ;
  assign \new_[1096]_  = ~\new_[1645]_  | ~\new_[5249]_  | ~\new_[1622]_  | ~\new_[1409]_ ;
  assign \new_[1097]_  = ~\new_[1207]_ ;
  assign \new_[1098]_  = ~\new_[1209]_ ;
  assign \new_[1099]_  = ~\new_[1584]_  | ~\new_[1375]_ ;
  assign \new_[1100]_  = ~\new_[1370]_  | ~\new_[1504]_ ;
  assign \new_[1101]_  = ~\new_[1210]_ ;
  assign \new_[1102]_  = ~\new_[1316]_  | ~\new_[1455]_ ;
  assign \new_[1103]_  = ~\new_[1626]_  | ~\new_[5245]_  | ~\new_[1622]_  | ~\new_[1409]_ ;
  assign \new_[1104]_  = ~\new_[1320]_  | ~\new_[1533]_ ;
  assign \new_[1105]_  = ~\new_[1583]_  | ~\new_[1380]_ ;
  assign \new_[1106]_  = ~\new_[4724]_  | ~\new_[1357]_ ;
  assign \new_[1107]_  = ~\new_[1535]_  | ~\new_[1536]_ ;
  assign \new_[1108]_  = ~\new_[1216]_ ;
  assign \new_[1109]_  = ~\new_[1219]_ ;
  assign \new_[1110]_  = ~\new_[1220]_ ;
  assign \new_[1111]_  = ~\new_[1583]_  | ~\new_[1371]_ ;
  assign \new_[1112]_  = ~\new_[1624]_  | ~\new_[1376]_ ;
  assign \new_[1113]_  = ~\new_[1222]_ ;
  assign \new_[1114]_  = ~\new_[1225]_ ;
  assign \new_[1115]_  = ~\new_[4615]_  | ~\new_[1357]_ ;
  assign \new_[1116]_  = ~\new_[1320]_  | ~\new_[5047]_ ;
  assign \new_[1117]_  = ~\new_[5154]_  | ~\new_[1376]_ ;
  assign \new_[1118]_  = ~\new_[1489]_  | ~\new_[1430]_  | ~\new_[4390]_ ;
  assign \new_[1119]_  = ~\new_[1228]_ ;
  assign \new_[1120]_  = ~\new_[1320]_  & ~\new_[5055]_ ;
  assign \new_[1121]_  = ~\new_[1518]_  & ~\new_[1382]_ ;
  assign \new_[1122]_  = ~\new_[1231]_ ;
  assign \new_[1123]_  = ~\new_[1232]_ ;
  assign \new_[1124]_  = ~\new_[1395]_  | ~\new_[5210]_  | ~\new_[1521]_ ;
  assign \new_[1125]_  = ~\new_[1510]_  | ~\new_[1552]_  | ~\new_[1408]_ ;
  assign \new_[1126]_  = ~\new_[1378]_  | ~\new_[1344]_ ;
  assign \new_[1127]_  = ~\new_[1336]_  & ~\new_[1368]_ ;
  assign \new_[1128]_  = ~\new_[1365]_  | ~\new_[1459]_ ;
  assign \new_[1129]_  = ~\new_[1549]_  & ~\new_[1346]_ ;
  assign \new_[1130]_  = ~\new_[1402]_  | ~\new_[1358]_ ;
  assign \new_[1131]_  = ~\new_[1293]_  & (~\new_[1515]_  | ~\new_[1395]_ );
  assign \new_[1132]_  = ~\new_[1568]_  | ~\new_[1301]_ ;
  assign \new_[1133]_  = \new_[4999]_  & \new_[1318]_ ;
  assign \new_[1134]_  = ~\new_[1236]_ ;
  assign \new_[1135]_  = ~\new_[1305]_  | ~\new_[1386]_ ;
  assign \new_[1136]_  = ~\new_[1240]_ ;
  assign \new_[1137]_  = ~\new_[1241]_ ;
  assign \new_[1138]_  = ~\new_[1576]_  & ~\new_[1474]_ ;
  assign \new_[1139]_  = ~\new_[1245]_ ;
  assign \new_[1140]_  = ~\new_[1420]_  | ~\new_[1304]_ ;
  assign \new_[1141]_  = ~\new_[1525]_  | ~\new_[4842]_ ;
  assign \new_[1142]_  = ~\new_[1512]_  | ~\new_[1399]_ ;
  assign \new_[1143]_  = ~\new_[1179]_  | ~\new_[1296]_ ;
  assign \new_[1144]_  = ~\new_[4612]_ ;
  assign \new_[1145]_  = ~\new_[5201]_  | ~\new_[1303]_ ;
  assign \new_[1146]_  = ~\new_[1253]_ ;
  assign \new_[1147]_  = ~\new_[1581]_  | ~\new_[1296]_ ;
  assign \new_[1148]_  = ~\new_[1566]_  | ~\new_[1303]_ ;
  assign \new_[1149]_  = ~\new_[1569]_  | ~\new_[1302]_ ;
  assign \new_[1150]_  = ~\new_[1267]_ ;
  assign \new_[1151]_  = ~\new_[4645]_  | ~\new_[1304]_ ;
  assign \new_[1152]_  = ~\new_[1428]_  | ~\new_[4840]_ ;
  assign \new_[1153]_  = ~\new_[1270]_ ;
  assign \new_[1154]_  = ~\new_[1497]_  & ~\new_[1411]_ ;
  assign \new_[1155]_  = ~\new_[5110]_  | ~\new_[4874]_ ;
  assign \new_[1156]_  = ~\new_[1553]_  | ~\new_[1320]_ ;
  assign \new_[1157]_  = ~\new_[1278]_ ;
  assign \new_[1158]_  = ~\new_[1279]_ ;
  assign \new_[1159]_  = ~\new_[1285]_ ;
  assign \new_[1160]_  = ~\new_[1298]_  & ~\new_[1554]_ ;
  assign \new_[1161]_  = \new_[1526]_  & \new_[4390]_ ;
  assign \new_[1162]_  = ~\new_[4607]_  | ~\new_[1304]_ ;
  assign \new_[1163]_  = ~\new_[1296]_ ;
  assign \new_[1164]_  = ~\new_[1429]_  | ~\new_[5084]_ ;
  assign \new_[1165]_  = ~\new_[5082]_  & ~\new_[5121]_ ;
  assign \new_[1166]_  = ~\new_[1302]_ ;
  assign \new_[1167]_  = ~\new_[1510]_  | ~\new_[4857]_ ;
  assign \new_[1168]_  = \new_[1579]_  & \new_[5287]_ ;
  assign \new_[1169]_  = ~\new_[4794]_  & ~\new_[5111]_ ;
  assign \new_[1170]_  = ~\new_[1305]_ ;
  assign \new_[1171]_  = ~\new_[1310]_ ;
  assign \new_[1172]_  = ~\new_[1310]_ ;
  assign \new_[1173]_  = ~\new_[1419]_  | ~\new_[4857]_ ;
  assign \new_[1174]_  = ~\new_[1312]_ ;
  assign \new_[1175]_  = ~\new_[1314]_ ;
  assign \new_[1176]_  = ~\new_[1506]_ ;
  assign \new_[1177]_  = ~\new_[1318]_ ;
  assign \new_[1178]_  = ~\new_[1319]_ ;
  assign \new_[1179]_  = ~\new_[1520]_ ;
  assign \new_[1180]_  = ~\new_[1322]_ ;
  assign \new_[1181]_  = ~\new_[1507]_  | ~\new_[1434]_ ;
  assign \new_[1182]_  = ~\new_[1562]_  | ~\new_[1433]_ ;
  assign \new_[1183]_  = ~\new_[1418]_  | ~\new_[1531]_ ;
  assign \new_[1184]_  = ~\new_[1417]_  | ~\new_[1436]_ ;
  assign \new_[1185]_  = ~\new_[1607]_  | ~\new_[1433]_ ;
  assign \new_[1186]_  = ~\new_[1565]_  | ~\new_[1662]_  | ~\new_[1563]_  | ~\new_[1517]_ ;
  assign \new_[1187]_  = ~\new_[1565]_  | ~\new_[1637]_  | ~\new_[1605]_  | ~\new_[1517]_ ;
  assign \new_[1188]_  = ~\new_[1605]_  | ~\new_[1436]_ ;
  assign \new_[1189]_  = ~\new_[1471]_  | ~\new_[1517]_  | ~\new_[1512]_ ;
  assign \new_[1190]_  = ~\new_[1323]_ ;
  assign \new_[1191]_  = ~\new_[1607]_  | ~\new_[1434]_ ;
  assign \new_[1192]_  = ~\new_[1542]_  | ~\new_[1574]_  | ~\new_[1471]_ ;
  assign \new_[1193]_  = ~\new_[1435]_  | ~\new_[1398]_ ;
  assign \new_[1194]_  = ~\new_[1325]_ ;
  assign \new_[1195]_  = ~\new_[1407]_  & ~\new_[1530]_ ;
  assign \new_[1196]_  = ~\new_[1530]_  | ~\new_[1460]_ ;
  assign \new_[1197]_  = ~\new_[1442]_  & ~\new_[1441]_ ;
  assign \new_[1198]_  = ~\new_[1429]_  | ~\new_[1446]_ ;
  assign \new_[1199]_  = ~\new_[4604]_  | ~\new_[1532]_ ;
  assign \new_[1200]_  = ~\new_[1408]_  | ~\new_[1531]_ ;
  assign \new_[1201]_  = ~\new_[1634]_  | ~\new_[1432]_ ;
  assign \new_[1202]_  = ~\new_[1607]_  | ~\new_[1436]_ ;
  assign \new_[1203]_  = ~\new_[1667]_  | ~\new_[5250]_  | ~\new_[1621]_  | ~\new_[1496]_ ;
  assign \new_[1204]_  = ~\new_[1455]_  | ~\new_[1416]_ ;
  assign \new_[1205]_  = ~\new_[1504]_  & ~\new_[1450]_ ;
  assign \new_[1206]_  = ~\new_[1326]_ ;
  assign \new_[1207]_  = ~\new_[5049]_  | ~\new_[1452]_ ;
  assign \new_[1208]_  = ~\new_[4585]_  | ~\new_[1533]_ ;
  assign \new_[1209]_  = ~\new_[1583]_  | ~\new_[1447]_ ;
  assign \new_[1210]_  = ~\new_[1416]_  | ~\new_[1454]_ ;
  assign \new_[1211]_  = ~\new_[1622]_  | ~\new_[1462]_ ;
  assign \new_[1212]_  = ~\new_[1645]_  | ~\new_[1451]_ ;
  assign \new_[1213]_  = ~\new_[1585]_  | ~\new_[1449]_ ;
  assign \new_[1214]_  = ~\new_[1328]_ ;
  assign \new_[1215]_  = ~\new_[1329]_ ;
  assign \new_[1216]_  = ~\new_[1645]_  | ~\new_[5250]_  | ~\new_[1622]_  | ~\new_[1495]_ ;
  assign \new_[1217]_  = ~\new_[1330]_ ;
  assign \new_[1218]_  = ~\new_[1331]_ ;
  assign \new_[1219]_  = ~\new_[4397]_  | ~\new_[1458]_ ;
  assign \new_[1220]_  = ~\new_[1465]_  | ~\new_[1585]_ ;
  assign \new_[1221]_  = ~\new_[1332]_ ;
  assign \new_[1222]_  = ~\new_[1623]_  | ~\new_[5246]_  | ~\new_[1644]_  | ~\new_[1494]_ ;
  assign \new_[1223]_  = ~\new_[1409]_  | ~\new_[1465]_ ;
  assign \new_[1224]_  = ~\new_[1499]_  & ~\new_[1464]_ ;
  assign \new_[1225]_  = ~\new_[1519]_  | ~\new_[5047]_ ;
  assign \new_[1226]_  = ~\new_[1463]_  | ~\new_[5111]_ ;
  assign \new_[1227]_  = ~\new_[1583]_  | ~\new_[1462]_ ;
  assign \new_[1228]_  = ~\new_[1334]_ ;
  assign \new_[1229]_  = ~\new_[4744]_ ;
  assign \new_[1230]_  = ~\new_[1335]_ ;
  assign \new_[1231]_  = ~\new_[1503]_  & ~\new_[1464]_ ;
  assign \new_[1232]_  = ~\new_[1559]_  | ~\new_[1497]_  | ~\new_[1500]_ ;
  assign \new_[1233]_  = ~\new_[1443]_  & ~\new_[1444]_ ;
  assign \new_[1234]_  = ~\new_[1478]_  & (~\new_[1581]_  | ~\new_[1477]_ );
  assign \new_[1235]_  = ~\new_[5211]_  & ~\new_[4699]_ ;
  assign \new_[1236]_  = ~\new_[1552]_  | ~\new_[4720]_ ;
  assign \new_[1237]_  = ~\new_[1511]_  & ~\new_[4758]_ ;
  assign \new_[1238]_  = ~\new_[1338]_ ;
  assign \new_[1239]_  = ~\new_[1339]_ ;
  assign \new_[1240]_  = ~\new_[1605]_  | ~\new_[1389]_ ;
  assign \new_[1241]_  = ~\new_[1340]_ ;
  assign \new_[1242]_  = ~\new_[1341]_ ;
  assign \new_[1243]_  = ~\new_[1343]_ ;
  assign \new_[1244]_  = ~\new_[4888]_  & ~\new_[1472]_ ;
  assign \new_[1245]_  = ~\new_[4885]_  & ~\new_[4841]_ ;
  assign \new_[1246]_  = ~\new_[1573]_  | ~\new_[1389]_ ;
  assign \new_[1247]_  = ~\new_[4644]_  | ~\new_[1397]_ ;
  assign \new_[1248]_  = ~\new_[1565]_  | ~\new_[1399]_ ;
  assign \new_[1249]_  = ~\new_[1347]_ ;
  assign \new_[1250]_  = ~\new_[1605]_  | ~\new_[1385]_ ;
  assign \new_[1251]_  = ~\new_[1348]_ ;
  assign \new_[1252]_  = ~\new_[4803]_  & ~\new_[1407]_ ;
  assign \new_[1253]_  = ~\new_[1400]_  | ~\new_[1567]_ ;
  assign \new_[1254]_  = ~\new_[1581]_  & ~\new_[1393]_ ;
  assign \new_[1255]_  = ~\new_[1619]_  | ~\new_[1387]_ ;
  assign \new_[1256]_  = ~\new_[4615]_  | ~\new_[4723]_ ;
  assign \new_[1257]_  = ~\new_[1384]_  | ~\new_[1580]_ ;
  assign \new_[1258]_  = ~\new_[1351]_ ;
  assign \new_[1259]_  = ~\new_[1352]_ ;
  assign \new_[1260]_  = ~\new_[1428]_  | ~\new_[1467]_ ;
  assign \new_[1261]_  = ~\new_[1385]_  | ~\new_[1488]_ ;
  assign \new_[1262]_  = ~\new_[1613]_  | ~\new_[4392]_ ;
  assign \new_[1263]_  = ~\new_[1619]_  | ~\new_[4723]_ ;
  assign \new_[1264]_  = \new_[1550]_  & \new_[1387]_ ;
  assign \new_[1265]_  = ~\new_[1565]_  | ~\new_[1488]_ ;
  assign \new_[1266]_  = ~\new_[1388]_  | ~\new_[4615]_ ;
  assign \new_[1267]_  = ~\new_[1564]_  | ~\new_[1406]_  | ~\new_[1638]_ ;
  assign \new_[1268]_  = ~\new_[1361]_ ;
  assign \new_[1269]_  = ~\new_[1362]_ ;
  assign \new_[1270]_  = ~\new_[1363]_ ;
  assign \new_[1271]_  = ~\new_[4888]_  | ~\new_[1482]_ ;
  assign \new_[1272]_  = ~\new_[4604]_  | ~\new_[1544]_ ;
  assign \new_[1273]_  = ~\new_[1368]_ ;
  assign \new_[1274]_  = ~\new_[1373]_ ;
  assign \new_[1275]_  = ~\new_[1410]_  | ~\new_[1504]_ ;
  assign \new_[1276]_  = ~\new_[1410]_  & ~\new_[1498]_ ;
  assign \new_[1277]_  = ~\new_[1374]_ ;
  assign \new_[1278]_  = ~\new_[1625]_  | ~\new_[1409]_ ;
  assign \new_[1279]_  = ~\new_[4607]_  | ~\new_[1397]_ ;
  assign \new_[1280]_  = ~\new_[5190]_  & ~\new_[4873]_ ;
  assign \new_[1281]_  = ~\new_[1535]_ ;
  assign \new_[1282]_  = ~\new_[1375]_ ;
  assign \new_[1283]_  = ~\new_[1553]_  | ~\new_[5048]_ ;
  assign \new_[1284]_  = ~\new_[1458]_ ;
  assign \new_[1285]_  = ~\new_[1409]_  | ~\new_[1548]_ ;
  assign \new_[1286]_  = ~\new_[1377]_ ;
  assign \new_[1287]_  = ~\new_[4795]_  | ~\new_[1518]_ ;
  assign \new_[1288]_  = ~\new_[1384]_  | ~\new_[1581]_ ;
  assign \new_[1289]_  = ~\new_[4624]_  & ~\new_[1401]_ ;
  assign \new_[1290]_  = ~\new_[1380]_ ;
  assign \new_[1291]_  = ~\new_[1385]_ ;
  assign \new_[1292]_  = \new_[1508]_  & \new_[4894]_ ;
  assign \new_[1293]_  = ~\new_[1580]_  & ~\new_[1513]_ ;
  assign \new_[1294]_  = ~\new_[1388]_ ;
  assign \new_[1295]_  = ~\new_[1616]_  & ~\new_[1513]_ ;
  assign \new_[1296]_  = ~\new_[1392]_ ;
  assign \new_[1297]_  = ~\new_[1527]_  | ~\new_[1526]_ ;
  assign \new_[1298]_  = ~\new_[5054]_  | ~\new_[5112]_ ;
  assign \new_[1299]_  = ~\new_[1662]_  | ~\new_[1609]_ ;
  assign \new_[1300]_  = ~\new_[1395]_ ;
  assign \new_[1301]_  = ~\new_[4699]_ ;
  assign \new_[1302]_  = ~\new_[4699]_ ;
  assign \new_[1303]_  = ~\new_[1580]_  & ~\new_[1521]_ ;
  assign \new_[1304]_  = ~\new_[1403]_ ;
  assign \new_[1305]_  = ~\new_[1525]_  | ~\new_[1642]_ ;
  assign \new_[1306]_  = ~\new_[1405]_ ;
  assign \new_[1307]_  = ~\new_[4535]_ ;
  assign \new_[1308]_  = ~\new_[4535]_ ;
  assign \new_[1309]_  = ~\new_[1408]_ ;
  assign \new_[1310]_  = ~\new_[4758]_ ;
  assign \new_[1311]_  = ~\new_[4873]_ ;
  assign \new_[1312]_  = ~\new_[1409]_ ;
  assign \new_[1313]_  = ~\new_[1412]_ ;
  assign \new_[1314]_  = ~\new_[1413]_ ;
  assign \new_[1315]_  = ~\new_[1414]_ ;
  assign \new_[1316]_  = \new_[1414]_ ;
  assign \new_[1317]_  = ~\new_[4417]_ ;
  assign \new_[1318]_  = ~\new_[1424]_ ;
  assign \new_[1319]_  = ~\new_[4782]_ ;
  assign \new_[1320]_  = ~\new_[4585]_ ;
  assign \new_[1321]_  = ~\new_[1427]_ ;
  assign \new_[1322]_  = ~\new_[1429]_ ;
  assign \new_[1323]_  = ~\new_[1638]_  | ~\new_[5243]_  | ~\new_[1594]_ ;
  assign \new_[1324]_  = ~\new_[4857]_ ;
  assign \new_[1325]_  = ~\new_[5282]_  & ~\new_[5243]_ ;
  assign \new_[1326]_  = ~\new_[1519]_  | ~\new_[1533]_ ;
  assign \new_[1327]_  = ~\new_[5050]_  & ~\new_[1534]_ ;
  assign \new_[1328]_  = ~\new_[1554]_  | ~\new_[1577]_  | ~\new_[4795]_ ;
  assign \new_[1329]_  = ~\new_[1559]_  & ~\new_[1536]_ ;
  assign \new_[1330]_  = ~\new_[1505]_  & ~\new_[1537]_ ;
  assign \new_[1331]_  = ~\new_[1559]_  & ~\new_[1538]_ ;
  assign \new_[1332]_  = ~\new_[1559]_  & ~\new_[1537]_ ;
  assign \new_[1333]_  = ~\new_[1501]_  & ~\new_[1538]_ ;
  assign \new_[1334]_  = ~\new_[5054]_  & ~\new_[5127]_ ;
  assign \new_[1335]_  = ~\new_[1538]_  & ~\new_[1505]_ ;
  assign \new_[1336]_  = ~\new_[4613]_  & ~\new_[1485]_ ;
  assign \new_[1337]_  = ~\new_[1594]_  | ~\new_[4719]_ ;
  assign \new_[1338]_  = ~\new_[1563]_  | ~\new_[1473]_ ;
  assign \new_[1339]_  = ~\new_[1498]_  | ~\new_[5001]_ ;
  assign \new_[1340]_  = ~\new_[4803]_  | ~\new_[4759]_ ;
  assign \new_[1341]_  = ~\new_[1432]_ ;
  assign \new_[1342]_  = ~\new_[1433]_ ;
  assign \new_[1343]_  = ~\new_[1474]_  & ~\new_[1575]_ ;
  assign \new_[1344]_  = ~\new_[1512]_  | ~\new_[1488]_ ;
  assign \new_[1345]_  = ~\new_[1609]_  & ~\new_[4568]_ ;
  assign \new_[1346]_  = ~\new_[1438]_ ;
  assign \new_[1347]_  = ~\new_[1575]_  & ~\new_[4568]_ ;
  assign \new_[1348]_  = ~\new_[1613]_  | ~\new_[1469]_ ;
  assign \new_[1349]_  = ~\new_[1484]_  & ~\new_[4838]_ ;
  assign \new_[1350]_  = ~\new_[1440]_ ;
  assign \new_[1351]_  = ~\new_[1470]_  & ~\new_[1580]_ ;
  assign \new_[1352]_  = ~\new_[4838]_  & ~\new_[1486]_ ;
  assign \new_[1353]_  = ~\new_[1514]_  | ~\new_[1479]_ ;
  assign \new_[1354]_  = ~\new_[1441]_ ;
  assign \new_[1355]_  = ~\new_[1442]_ ;
  assign \new_[1356]_  = ~\new_[1468]_  | ~\new_[1480]_ ;
  assign \new_[1357]_  = ~\new_[1468]_  | ~\new_[1540]_ ;
  assign \new_[1358]_  = ~\new_[1475]_  | ~\new_[1612]_ ;
  assign \new_[1359]_  = ~\new_[1444]_ ;
  assign \new_[1360]_  = ~\new_[1445]_ ;
  assign \new_[1361]_  = ~\new_[4893]_  | ~\new_[4884]_  | ~\new_[4644]_ ;
  assign \new_[1362]_  = ~\new_[4885]_  | ~\new_[4842]_ ;
  assign \new_[1363]_  = ~\new_[4885]_  & ~\new_[1472]_ ;
  assign \new_[1364]_  = ~\new_[1446]_ ;
  assign \new_[1365]_  = ~\new_[1447]_ ;
  assign \new_[1366]_  = ~\new_[1590]_  & ~\new_[1494]_ ;
  assign \new_[1367]_  = ~\new_[1585]_  | ~\new_[1483]_ ;
  assign \new_[1368]_  = ~\new_[1578]_  & ~\new_[1485]_ ;
  assign \new_[1369]_  = ~\new_[1449]_ ;
  assign \new_[1370]_  = ~\new_[1450]_ ;
  assign \new_[1371]_  = ~\new_[1495]_  & ~\new_[1547]_ ;
  assign \new_[1372]_  = ~\new_[1451]_ ;
  assign \new_[1373]_  = ~\new_[1519]_  | ~\new_[1493]_ ;
  assign \new_[1374]_  = ~\new_[1663]_  | ~\new_[5243]_ ;
  assign \new_[1375]_  = ~\new_[5246]_  & ~\new_[1495]_ ;
  assign \new_[1376]_  = ~\new_[1667]_  & ~\new_[1496]_ ;
  assign \new_[1377]_  = ~\new_[1460]_ ;
  assign \new_[1378]_  = ~\new_[1637]_  | ~\new_[1488]_ ;
  assign \new_[1379]_  = ~\new_[4831]_  & ~\new_[1486]_ ;
  assign \new_[1380]_  = ~\new_[1494]_  & ~\new_[1551]_ ;
  assign \new_[1381]_  = ~\new_[4624]_  | ~\new_[1487]_ ;
  assign \new_[1382]_  = ~\new_[1463]_ ;
  assign \new_[1383]_  = ~\new_[1568]_  & ~\new_[5211]_ ;
  assign \new_[1384]_  = ~\new_[1567]_  & ~\new_[1570]_ ;
  assign \new_[1385]_  = ~\new_[4568]_ ;
  assign \new_[1386]_  = ~\new_[1467]_ ;
  assign \new_[1387]_  = ~\new_[1468]_ ;
  assign \new_[1388]_  = ~\new_[1640]_  & ~\new_[4377]_ ;
  assign \new_[1389]_  = ~\new_[1474]_ ;
  assign \new_[1390]_  = ~\new_[1475]_ ;
  assign \new_[1391]_  = ~\new_[1476]_ ;
  assign \new_[1392]_  = ~\new_[1567]_  | ~\new_[5211]_ ;
  assign \new_[1393]_  = ~\new_[1477]_ ;
  assign \new_[1394]_  = ~\new_[1479]_ ;
  assign \new_[1395]_  = ~\new_[1484]_ ;
  assign \new_[1396]_  = ~\new_[4724]_ ;
  assign \new_[1397]_  = ~\new_[4888]_  & ~\new_[1642]_ ;
  assign \new_[1398]_  = ~\new_[1637]_  | ~\new_[1576]_ ;
  assign \new_[1399]_  = ~\new_[1634]_  & ~\new_[1574]_ ;
  assign \new_[1400]_  = ~\new_[1486]_ ;
  assign \new_[1401]_  = ~\new_[1487]_ ;
  assign \new_[1402]_  = ~\new_[1619]_  | ~\new_[1578]_ ;
  assign \new_[1403]_  = ~\new_[4888]_  | ~\new_[4885]_ ;
  assign \new_[1404]_  = ~\new_[1490]_ ;
  assign \new_[1405]_  = ~\new_[1491]_ ;
  assign \new_[1406]_  = ~\new_[4719]_ ;
  assign \new_[1407]_  = ~\new_[4719]_ ;
  assign \new_[1408]_  = \new_[4719]_ ;
  assign \new_[1409]_  = ~\new_[1494]_ ;
  assign \new_[1410]_  = ~\new_[1497]_ ;
  assign \new_[1411]_  = ~\new_[1498]_ ;
  assign \new_[1412]_  = ~\new_[1499]_ ;
  assign \new_[1413]_  = ~\new_[1501]_ ;
  assign \new_[1414]_  = ~\new_[1502]_ ;
  assign \new_[1415]_  = ~\new_[1504]_ ;
  assign \new_[1416]_  = ~\new_[1505]_ ;
  assign \new_[1417]_  = ~\new_[1508]_ ;
  assign \new_[1418]_  = ~\new_[1510]_ ;
  assign \new_[1419]_  = ~\new_[1511]_ ;
  assign \new_[1420]_  = ~\new_[4645]_ ;
  assign \new_[1421]_  = ~\new_[1515]_ ;
  assign \new_[1422]_  = ~\new_[5209]_ ;
  assign \new_[1423]_  = ~\new_[1516]_ ;
  assign \new_[1424]_  = ~\new_[1587]_  & (~\new_[1652]_  | ~\new_[2601]_ );
  assign \new_[1425]_  = ~\new_[5049]_ ;
  assign \new_[1426]_  = ~\new_[1521]_ ;
  assign \new_[1427]_  = ~\new_[1522]_ ;
  assign \new_[1428]_  = ~\new_[1525]_ ;
  assign \new_[1429]_  = \new_[1525]_ ;
  assign \new_[1430]_  = ~\new_[1526]_ ;
  assign \new_[1431]_  = ~\new_[1530]_ ;
  assign \new_[1432]_  = ~\new_[1610]_  & ~\new_[1542]_ ;
  assign \new_[1433]_  = ~\new_[1539]_  & ~\new_[1575]_ ;
  assign \new_[1434]_  = ~\new_[1574]_  & ~\new_[1542]_ ;
  assign \new_[1435]_  = ~\new_[1609]_  | ~\new_[1565]_  | ~\new_[1634]_ ;
  assign \new_[1436]_  = ~\new_[1609]_  & ~\new_[1539]_ ;
  assign \new_[1437]_  = ~\new_[4761]_ ;
  assign \new_[1438]_  = ~\new_[4885]_  | ~\new_[1544]_ ;
  assign \new_[1439]_  = ~\new_[1531]_ ;
  assign \new_[1440]_  = ~\new_[1543]_  & ~\new_[1620]_ ;
  assign \new_[1441]_  = ~\new_[1540]_  & ~\new_[1640]_ ;
  assign \new_[1442]_  = ~\new_[4628]_  & ~\new_[1540]_ ;
  assign \new_[1443]_  = ~\new_[4377]_  & ~\new_[1592]_ ;
  assign \new_[1444]_  = ~\new_[1614]_  & ~\new_[1543]_ ;
  assign \new_[1445]_  = ~\new_[4617]_  & ~\new_[1543]_ ;
  assign \new_[1446]_  = ~\new_[1642]_  & ~\new_[1545]_ ;
  assign \new_[1447]_  = ~\new_[1555]_  & ~\new_[1547]_ ;
  assign \new_[1448]_  = ~\new_[1622]_  | ~\new_[1546]_ ;
  assign \new_[1449]_  = ~\new_[1555]_  & ~\new_[1590]_ ;
  assign \new_[1450]_  = ~\new_[1558]_  | ~\new_[4398]_ ;
  assign \new_[1451]_  = ~\new_[1555]_  & ~\new_[1623]_ ;
  assign \new_[1452]_  = ~\new_[1534]_ ;
  assign \new_[1453]_  = ~\new_[1585]_  & ~\new_[1547]_ ;
  assign \new_[1454]_  = ~\new_[1535]_ ;
  assign \new_[1455]_  = ~\new_[1536]_ ;
  assign \new_[1456]_  = ~\new_[1621]_  | ~\new_[1548]_ ;
  assign \new_[1457]_  = ~\new_[1537]_ ;
  assign \new_[1458]_  = ~\new_[1556]_  & ~\new_[1559]_ ;
  assign \new_[1459]_  = ~\new_[1585]_  | ~\new_[1548]_ ;
  assign \new_[1460]_  = ~\new_[5244]_  | ~\new_[1663]_ ;
  assign \new_[1461]_  = ~\new_[1578]_  | ~\new_[1550]_ ;
  assign \new_[1462]_  = ~\new_[1555]_  & ~\new_[1591]_ ;
  assign \new_[1463]_  = ~\new_[4745]_ ;
  assign \new_[1464]_  = ~\new_[1556]_  | ~\new_[1559]_ ;
  assign \new_[1465]_  = ~\new_[1591]_  | ~\new_[1551]_ ;
  assign \new_[1466]_  = ~\new_[1539]_ ;
  assign \new_[1467]_  = ~\new_[4608]_  & ~\new_[4885]_ ;
  assign \new_[1468]_  = ~\new_[4378]_  | ~\new_[4625]_ ;
  assign \new_[1469]_  = ~\new_[1540]_ ;
  assign \new_[1470]_  = ~\new_[1617]_  | ~\new_[5069]_ ;
  assign \new_[1471]_  = ~\new_[1634]_  & ~\new_[1602]_ ;
  assign \new_[1472]_  = ~\new_[4608]_  | ~\new_[4891]_ ;
  assign \new_[1473]_  = ~\new_[1542]_ ;
  assign \new_[1474]_  = ~\new_[4572]_  | ~\new_[4574]_ ;
  assign \new_[1475]_  = ~\new_[1543]_ ;
  assign \new_[1476]_  = ~\new_[1617]_  | ~\new_[1604]_ ;
  assign \new_[1477]_  = ~\new_[4838]_  & ~\new_[5211]_ ;
  assign \new_[1478]_  = ~\new_[1617]_  & ~\new_[1604]_ ;
  assign \new_[1479]_  = ~\new_[1616]_  & ~\new_[5211]_ ;
  assign \new_[1480]_  = ~\new_[4378]_  | ~\new_[4618]_ ;
  assign \new_[1481]_  = ~\new_[1544]_ ;
  assign \new_[1482]_  = ~\new_[1545]_ ;
  assign \new_[1483]_  = ~\new_[1547]_ ;
  assign \new_[1484]_  = ~\new_[1615]_  | ~\new_[4611]_ ;
  assign \new_[1485]_  = ~\new_[1614]_  | ~\new_[1643]_ ;
  assign \new_[1486]_  = ~\new_[4700]_  | ~\new_[4611]_ ;
  assign \new_[1487]_  = ~\new_[1614]_  & ~\new_[4616]_ ;
  assign \new_[1488]_  = ~\new_[1660]_  & ~\new_[1610]_ ;
  assign \new_[1489]_  = ~\new_[1551]_ ;
  assign \new_[1490]_  = ~\new_[5001]_ ;
  assign \new_[1491]_  = ~\new_[5001]_ ;
  assign \new_[1492]_  = ~\new_[1553]_ ;
  assign \new_[1493]_  = ~\new_[4795]_ ;
  assign \new_[1494]_  = ~\new_[1555]_ ;
  assign \new_[1495]_  = ~\new_[1555]_ ;
  assign \new_[1496]_  = ~\new_[1555]_ ;
  assign \new_[1497]_  = ~\new_[1556]_ ;
  assign \new_[1498]_  = ~\new_[1557]_ ;
  assign \new_[1499]_  = ~\new_[1557]_ ;
  assign \new_[1500]_  = ~\new_[1557]_ ;
  assign \new_[1501]_  = ~\new_[1558]_ ;
  assign \new_[1502]_  = ~\new_[1558]_ ;
  assign \new_[1503]_  = ~\new_[1558]_ ;
  assign \new_[1504]_  = ~\new_[1559]_ ;
  assign \new_[1505]_  = ~\new_[1559]_ ;
  assign \new_[1506]_  = ~\new_[1562]_ ;
  assign \new_[1507]_  = \new_[1562]_ ;
  assign \new_[1508]_  = ~\new_[1563]_ ;
  assign \new_[1509]_  = ~\new_[1564]_ ;
  assign \new_[1510]_  = ~\new_[1564]_ ;
  assign \new_[1511]_  = ~\new_[1564]_ ;
  assign \new_[1512]_  = ~\new_[1565]_ ;
  assign \new_[1513]_  = ~\new_[1566]_ ;
  assign \new_[1514]_  = ~\new_[1566]_ ;
  assign \new_[1515]_  = ~\new_[5211]_ ;
  assign \new_[1516]_  = ~\new_[5084]_ ;
  assign \new_[1517]_  = ~\new_[1576]_ ;
  assign \new_[1518]_  = ~\new_[5192]_ ;
  assign \new_[1519]_  = ~\new_[1577]_ ;
  assign \new_[1520]_  = ~\new_[4831]_ ;
  assign \new_[1521]_  = ~\new_[4832]_ ;
  assign \new_[1522]_  = ~\new_[1579]_ ;
  assign \new_[1523]_  = \new_[4975]_ ;
  assign \new_[1524]_  = ~\new_[4975]_ ;
  assign \new_[1525]_  = ~\new_[4888]_ ;
  assign \new_[1526]_  = ~\new_[1585]_ ;
  assign \new_[1527]_  = ~\new_[1586]_ ;
  assign \new_[1528]_  = ~\new_[1628]_  | ~\new_[3147]_ ;
  assign \new_[1529]_  = \new_[1628]_  | \new_[3147]_ ;
  assign \new_[1530]_  = ~\new_[1593]_  | ~\new_[1663]_ ;
  assign \new_[1531]_  = ~\new_[1588]_ ;
  assign \new_[1532]_  = ~\new_[4885]_  & ~\new_[1589]_ ;
  assign \new_[1533]_  = ~\new_[5133]_  & ~\new_[4747]_ ;
  assign \new_[1534]_  = ~\new_[4747]_  | ~\new_[5133]_ ;
  assign \new_[1535]_  = ~\new_[1597]_  | ~\new_[4399]_ ;
  assign \new_[1536]_  = ~\new_[1596]_  | ~\new_[4400]_ ;
  assign \new_[1537]_  = ~\new_[1597]_  | ~\new_[4400]_ ;
  assign \new_[1538]_  = ~\new_[1596]_  | ~\new_[4399]_ ;
  assign \new_[1539]_  = ~\new_[4573]_  | ~\new_[4574]_ ;
  assign \new_[1540]_  = ~\new_[4672]_  | ~\new_[4626]_ ;
  assign \new_[1541]_  = ~\new_[1633]_  | ~\new_[4892]_ ;
  assign \new_[1542]_  = ~\new_[4573]_  | ~\new_[4569]_ ;
  assign \new_[1543]_  = ~\new_[1639]_  | ~\new_[4672]_ ;
  assign \new_[1544]_  = ~\new_[1589]_ ;
  assign \new_[1545]_  = ~\new_[4646]_  | ~\new_[1665]_ ;
  assign \new_[1546]_  = ~\new_[1590]_ ;
  assign \new_[1547]_  = ~\new_[1667]_  | ~\new_[5247]_ ;
  assign \new_[1548]_  = ~\new_[1591]_ ;
  assign \new_[1549]_  = ~\new_[4890]_  & ~\new_[4884]_ ;
  assign \new_[1550]_  = ~\new_[1592]_ ;
  assign \new_[1551]_  = ~\new_[1680]_  | ~\new_[5250]_ ;
  assign \new_[1552]_  = ~\new_[1594]_ ;
  assign \new_[1553]_  = ~\new_[4796]_ ;
  assign \new_[1554]_  = ~\new_[4796]_ ;
  assign \new_[1555]_  = ~\new_[1595]_ ;
  assign \new_[1556]_  = ~\new_[1597]_ ;
  assign \new_[1557]_  = ~\new_[1598]_ ;
  assign \new_[1558]_  = \new_[1598]_ ;
  assign \new_[1559]_  = ~\new_[1599]_ ;
  assign \new_[1560]_  = ~\new_[1651]_  | ~\new_[4464]_ ;
  assign \new_[1561]_  = \new_[1651]_  | \new_[4464]_ ;
  assign \new_[1562]_  = ~\new_[1602]_ ;
  assign \new_[1563]_  = ~\new_[1602]_ ;
  assign \new_[1564]_  = ~\new_[1603]_ ;
  assign \new_[1565]_  = \new_[4572]_ ;
  assign \new_[1566]_  = \new_[1604]_ ;
  assign \new_[1567]_  = ~\new_[1604]_ ;
  assign \new_[1568]_  = ~\new_[4838]_ ;
  assign \new_[1569]_  = \new_[5211]_ ;
  assign \new_[1570]_  = ~\new_[5211]_ ;
  assign \new_[1571]_  = ~\new_[1607]_ ;
  assign \new_[1572]_  = ~\new_[1606]_ ;
  assign \new_[1573]_  = ~\new_[1606]_ ;
  assign \new_[1574]_  = ~\new_[1609]_ ;
  assign \new_[1575]_  = ~\new_[1610]_ ;
  assign \new_[1576]_  = \new_[1610]_ ;
  assign \new_[1577]_  = ~\new_[4794]_ ;
  assign \new_[1578]_  = ~\new_[4624]_ ;
  assign \new_[1579]_  = ~\new_[1614]_ ;
  assign \new_[1580]_  = ~\new_[1616]_ ;
  assign \new_[1581]_  = \new_[1617]_ ;
  assign \new_[1582]_  = ~\new_[1618]_ ;
  assign \new_[1583]_  = ~\new_[1621]_ ;
  assign \new_[1584]_  = ~\new_[1622]_ ;
  assign \new_[1585]_  = ~\new_[1624]_ ;
  assign \new_[1586]_  = ~\new_[1625]_ ;
  assign \new_[1587]_  = ~\new_[1652]_  & ~\new_[2601]_ ;
  assign \new_[1588]_  = ~\new_[4862]_  | ~\new_[4861]_ ;
  assign \new_[1589]_  = ~\new_[4648]_  | ~\new_[4892]_ ;
  assign \new_[1590]_  = ~\new_[1680]_  | ~\new_[5248]_ ;
  assign \new_[1591]_  = ~\new_[1666]_  | ~\new_[5248]_ ;
  assign \new_[1592]_  = ~\new_[1664]_  | ~\new_[4628]_ ;
  assign \new_[1593]_  = ~\new_[4862]_ ;
  assign \new_[1594]_  = ~\new_[4862]_ ;
  assign \new_[1595]_  = ~\new_[1675]_  | ~\new_[1657]_ ;
  assign \new_[1596]_  = \new_[1629]_ ;
  assign \new_[1597]_  = ~\new_[1629]_ ;
  assign \new_[1598]_  = ~\new_[1677]_  | ~\new_[1658]_ ;
  assign \new_[1599]_  = ~\new_[1678]_  | ~\new_[1659]_ ;
  assign \new_[1600]_  = ~\new_[1670]_  | ~n1035;
  assign \new_[1601]_  = ~\new_[1671]_  | ~n1190;
  assign \new_[1602]_  = ~\new_[1682]_  | ~\new_[1669]_ ;
  assign \new_[1603]_  = ~\new_[4804]_ ;
  assign \new_[1604]_  = ~\new_[5069]_ ;
  assign \new_[1605]_  = ~\new_[1634]_ ;
  assign \new_[1606]_  = \new_[1635]_ ;
  assign \new_[1607]_  = ~\new_[1635]_ ;
  assign \new_[1608]_  = \new_[1635]_ ;
  assign \new_[1609]_  = ~\new_[1636]_ ;
  assign \new_[1610]_  = ~\new_[1636]_ ;
  assign \new_[1611]_  = ~\new_[1638]_ ;
  assign \new_[1612]_  = ~\new_[1640]_ ;
  assign \new_[1613]_  = \new_[1640]_ ;
  assign \new_[1614]_  = ~\new_[1641]_ ;
  assign \new_[1615]_  = ~\new_[4700]_ ;
  assign \new_[1616]_  = ~\new_[4700]_ ;
  assign \new_[1617]_  = \new_[4708]_ ;
  assign \new_[1618]_  = \new_[1643]_ ;
  assign \new_[1619]_  = ~\new_[1643]_ ;
  assign \new_[1620]_  = ~\new_[4617]_ ;
  assign \new_[1621]_  = ~\new_[4710]_ ;
  assign \new_[1622]_  = ~\new_[4710]_ ;
  assign \new_[1623]_  = ~\new_[4710]_ ;
  assign \new_[1624]_  = ~\new_[4710]_ ;
  assign \new_[1625]_  = ~\new_[1645]_ ;
  assign \new_[1626]_  = ~\new_[1645]_ ;
  assign \new_[1627]_  = ~\new_[1672]_  | ~n1025;
  assign \new_[1628]_  = ~\new_[1711]_  | ~\new_[2117]_  | ~\new_[2366]_  | ~\new_[1978]_ ;
  assign \new_[1629]_  = ~\new_[1676]_  | (~\new_[1716]_  & ~\new_[3284]_ );
  assign \new_[1630]_  = ~\new_[1685]_  | ~\new_[2595]_ ;
  assign \new_[1631]_  = ~\new_[1686]_  | ~\new_[3284]_ ;
  assign \new_[1632]_  = ~\new_[1687]_  | ~n1020;
  assign \new_[1633]_  = ~\new_[4648]_ ;
  assign \new_[1634]_  = ~\new_[1660]_ ;
  assign \new_[1635]_  = \new_[1660]_ ;
  assign \new_[1636]_  = ~\new_[1661]_ ;
  assign \new_[1637]_  = ~\new_[1662]_ ;
  assign \new_[1638]_  = ~\new_[1663]_ ;
  assign \new_[1639]_  = ~\new_[4626]_ ;
  assign \new_[1640]_  = ~\new_[1664]_ ;
  assign \new_[1641]_  = ~\new_[1664]_ ;
  assign \new_[1642]_  = ~\new_[4885]_ ;
  assign \new_[1643]_  = ~\new_[4618]_ ;
  assign \new_[1644]_  = ~\new_[1667]_ ;
  assign \new_[1645]_  = ~\new_[1667]_ ;
  assign \new_[1646]_  = ~\new_[1700]_  | ~\new_[1681]_ ;
  assign \new_[1647]_  = ~\new_[1690]_  | ~\new_[4704]_ ;
  assign \new_[1648]_  = ~\new_[1689]_  | ~\new_[2226]_ ;
  assign \new_[1649]_  = ~\new_[4735]_  | ~\new_[2442]_ ;
  assign \new_[1650]_  = \new_[1690]_  | \new_[4704]_ ;
  assign \new_[1651]_  = ~\new_[1730]_  | ~\new_[2629]_  | ~\new_[1833]_  | ~\new_[1835]_ ;
  assign \new_[1652]_  = ~\new_[1731]_  | ~\new_[1914]_  | ~\new_[1841]_  | ~\new_[2086]_ ;
  assign \new_[1653]_  = ~\new_[1881]_  & ~\new_[1691]_ ;
  assign \new_[1654]_  = ~\new_[1729]_  | ~\new_[2012]_  | ~\new_[2145]_  | ~\new_[2011]_ ;
  assign \new_[1655]_  = ~\new_[4839]_  | ~n1240;
  assign \new_[1656]_  = ~\new_[5134]_  | ~\new_[2580]_ ;
  assign \new_[1657]_  = ~\new_[1703]_  | ~n1140;
  assign \new_[1658]_  = ~\new_[1705]_  | ~n1110;
  assign \new_[1659]_  = ~\new_[1704]_  | ~n1115;
  assign \new_[1660]_  = n1225 ? \new_[1719]_  : \new_[2692]_ ;
  assign \new_[1661]_  = n1135 ? \new_[5060]_  : \new_[2669]_ ;
  assign \new_[1662]_  = ~\new_[4569]_ ;
  assign \new_[1663]_  = \new_[4833]_ ;
  assign \new_[1664]_  = ~\new_[1679]_ ;
  assign \new_[1665]_  = ~\new_[4892]_ ;
  assign \new_[1666]_  = ~\new_[1680]_ ;
  assign \new_[1667]_  = ~\new_[1680]_ ;
  assign \new_[1668]_  = ~\new_[1706]_  | ~n990;
  assign \new_[1669]_  = ~\new_[1707]_  | ~n1010;
  assign \new_[1670]_  = ~\new_[1685]_ ;
  assign \new_[1671]_  = ~\new_[1686]_ ;
  assign \new_[1672]_  = ~\new_[4735]_ ;
  assign \new_[1673]_  = ~\new_[1692]_ ;
  assign \new_[1674]_  = ~\new_[1695]_ ;
  assign \new_[1675]_  = ~\new_[4691]_  | ~\new_[2732]_ ;
  assign \new_[1676]_  = ~\new_[1716]_  | ~\new_[3284]_ ;
  assign \new_[1677]_  = ~\new_[1718]_  | ~\new_[2854]_ ;
  assign \new_[1678]_  = ~\new_[1717]_  | ~\new_[2853]_ ;
  assign \new_[1679]_  = \new_[2992]_  ? \new_[1736]_  : \new_[2851]_ ;
  assign \new_[1680]_  = ~\new_[1699]_ ;
  assign \new_[1681]_  = ~\new_[1725]_  | ~n1140;
  assign \new_[1682]_  = ~\new_[4591]_  | ~\new_[2597]_ ;
  assign \new_[1683]_  = ~\new_[1720]_  | ~\new_[3256]_ ;
  assign \new_[1684]_  = ~\new_[1721]_  | ~n1005;
  assign \new_[1685]_  = ~\new_[1756]_  | ~\new_[2165]_  | ~\new_[1803]_  | ~\new_[1972]_ ;
  assign \new_[1686]_  = ~\new_[1804]_  | ~\new_[2028]_  | ~\new_[1757]_  | ~\new_[1979]_ ;
  assign \new_[1687]_  = ~\new_[5134]_ ;
  assign \new_[1688]_  = ~\new_[1854]_  | ~\new_[1853]_  | ~\new_[1758]_  | ~\new_[1861]_ ;
  assign \new_[1689]_  = ~\new_[1706]_ ;
  assign \new_[1690]_  = ~\new_[1980]_  | ~\new_[1760]_  | ~\new_[1847]_  | ~\new_[1974]_ ;
  assign \new_[1691]_  = ~\new_[2166]_  | ~\new_[1740]_  | ~\new_[1898]_ ;
  assign \new_[1692]_  = (~\new_[1743]_  & ~\new_[3713]_ ) | (~\new_[2872]_  & ~\new_[4311]_ );
  assign \new_[1693]_  = (~\new_[1751]_  | ~\new_[3739]_ ) & (~\new_[3713]_  | ~\desIn[22] );
  assign \new_[1694]_  = ~\new_[4987]_ ;
  assign \new_[1695]_  = (~\new_[1748]_  & ~\new_[3713]_ ) | (~\new_[2872]_  & ~\new_[4361]_ );
  assign \new_[1696]_  = ~\new_[1710]_ ;
  assign \new_[1697]_  = ~\new_[1712]_ ;
  assign \new_[1698]_  = ~\new_[1713]_ ;
  assign \new_[1699]_  = n995 ? \new_[4599]_  : \new_[2602]_ ;
  assign \new_[1700]_  = ~\new_[4814]_  | ~\new_[2732]_ ;
  assign \new_[1701]_  = ~\new_[1733]_  | ~\new_[3149]_ ;
  assign \new_[1702]_  = ~\new_[4728]_  | ~\new_[2599]_ ;
  assign \new_[1703]_  = ~\new_[4691]_ ;
  assign \new_[1704]_  = ~\new_[1717]_ ;
  assign \new_[1705]_  = ~\new_[1718]_ ;
  assign \new_[1706]_  = ~\new_[1844]_  & ~\new_[5212]_ ;
  assign \new_[1707]_  = ~\new_[4591]_ ;
  assign \new_[1708]_  = ~\new_[1724]_ ;
  assign \new_[1709]_  = ~\new_[1728]_ ;
  assign \new_[1710]_  = (~\new_[1769]_  & ~\new_[3713]_ ) | (~\new_[3739]_  & ~\new_[4358]_ );
  assign \new_[1711]_  = ~\new_[2115]_  & ~\new_[1742]_ ;
  assign \new_[1712]_  = (~\new_[1771]_  & ~\new_[3713]_ ) | (~\new_[3739]_  & ~\new_[4357]_ );
  assign \new_[1713]_  = (~\new_[1772]_  & ~\new_[3713]_ ) | (~\new_[2872]_  & ~\new_[4363]_ );
  assign \new_[1714]_  = (~\new_[1754]_  | ~\new_[3739]_ ) & (~\new_[3713]_  | ~\desIn[54] );
  assign \new_[1715]_  = ~\new_[4942]_  | ~\new_[2853]_ ;
  assign \new_[1716]_  = ~\new_[2353]_  | ~\new_[1957]_  | ~\new_[1790]_  | ~\new_[2354]_ ;
  assign \new_[1717]_  = ~\new_[2132]_  | ~\new_[1789]_  | ~\new_[1888]_  | ~\new_[1994]_ ;
  assign \new_[1718]_  = ~\new_[2357]_  | ~\new_[1792]_  | ~\new_[1775]_  | ~\new_[1992]_ ;
  assign \new_[1719]_  = ~\new_[1836]_  & ~\new_[4473]_ ;
  assign \new_[1720]_  = ~\new_[1733]_ ;
  assign \new_[1721]_  = ~\new_[4728]_ ;
  assign \new_[1722]_  = ~\new_[1735]_ ;
  assign \new_[1723]_  = ~\new_[1737]_ ;
  assign \new_[1724]_  = ~\new_[2338]_  | ~\new_[1805]_  | ~\new_[1797]_  | ~\new_[2342]_ ;
  assign \new_[1725]_  = ~\new_[4814]_ ;
  assign \new_[1726]_  = ~\new_[1886]_  | ~\new_[1800]_  | ~\new_[2100]_  | ~\new_[2330]_ ;
  assign \new_[1727]_  = ~\new_[1806]_  | ~\new_[1807]_  | ~\new_[1988]_  | ~\new_[1911]_ ;
  assign \new_[1728]_  = (~\new_[1777]_  & ~\new_[3713]_ ) | (~\new_[2872]_  & ~\new_[4297]_ );
  assign \new_[1729]_  = ~\new_[1902]_  & ~\new_[1759]_ ;
  assign \new_[1730]_  = ~\new_[1738]_ ;
  assign \new_[1731]_  = ~\new_[1739]_ ;
  assign \new_[1732]_  = \new_[4930]_  | \new_[4939]_  | \new_[3290]_  | \new_[4938]_ ;
  assign \new_[1733]_  = ~\new_[1935]_  & ~\new_[4664]_ ;
  assign \new_[1734]_  = ~\new_[2101]_  | ~\new_[1875]_  | ~\new_[1827]_  | ~\new_[1970]_ ;
  assign \new_[1735]_  = ~\new_[2317]_  | ~\new_[1826]_  | ~\new_[2319]_  | ~\new_[1874]_ ;
  assign \new_[1736]_  = ~\new_[2104]_  | ~\new_[1830]_  | ~\new_[1845]_  | ~\new_[2107]_ ;
  assign \new_[1737]_  = ~\new_[2109]_  | ~\new_[2110]_  | ~\new_[1831]_  | ~\new_[1877]_ ;
  assign \new_[1738]_  = ~\new_[1890]_  | ~\new_[1834]_  | ~\new_[1862]_  | ~\new_[1858]_ ;
  assign \new_[1739]_  = ~\new_[1960]_  | ~\new_[1857]_  | ~\new_[1998]_  | ~\new_[2299]_ ;
  assign \new_[1740]_  = ~\new_[4853]_ ;
  assign \new_[1741]_  = ~\new_[1761]_ ;
  assign \new_[1742]_  = ~\new_[1779]_  | ~\new_[1780]_ ;
  assign \new_[1743]_  = (~\new_[1809]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[454]_ );
  assign \new_[1744]_  = (~\new_[1810]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[436]_ );
  assign \new_[1745]_  = \new_[474]_  ? \new_[3489]_  : \new_[1811]_ ;
  assign \new_[1746]_  = \new_[473]_  ? \new_[3489]_  : \new_[1812]_ ;
  assign \new_[1747]_  = (~\new_[1784]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[4346]_ );
  assign \new_[1748]_  = (~\new_[1781]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[442]_ );
  assign \new_[1749]_  = (~\new_[1782]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[492]_ );
  assign \new_[1750]_  = (~\new_[1785]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[4370]_ );
  assign \new_[1751]_  = \new_[438]_  ? \new_[3489]_  : \new_[1783]_ ;
  assign \new_[1752]_  = \new_[463]_  ? \new_[3489]_  : \new_[1786]_ ;
  assign \new_[1753]_  = (~\new_[1787]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[503]_ );
  assign \new_[1754]_  = \new_[440]_  ? \new_[3712]_  : \new_[1828]_ ;
  assign \new_[1755]_  = \new_[494]_  ? \new_[3489]_  : \new_[1829]_ ;
  assign \new_[1756]_  = ~\new_[1793]_  & ~\new_[1840]_ ;
  assign \new_[1757]_  = ~\new_[1848]_  & ~\new_[1794]_ ;
  assign \new_[1758]_  = ~\new_[1795]_  & ~\new_[1855]_ ;
  assign \new_[1759]_  = ~\new_[1808]_  | ~\new_[1852]_ ;
  assign \new_[1760]_  = ~\new_[1843]_  & ~\new_[1802]_ ;
  assign \new_[1761]_  = ~\new_[2164]_  | ~\new_[1801]_  | ~\new_[1968]_ ;
  assign \new_[1762]_  = \new_[490]_  ? \new_[3489]_  : \new_[1815]_ ;
  assign \new_[1763]_  = (~\new_[1813]_  & ~\new_[3754]_ ) | (~\new_[3712]_  & ~\new_[485]_ );
  assign \new_[1764]_  = \new_[472]_  ? \new_[3489]_  : \new_[1814]_ ;
  assign \new_[1765]_  = \new_[434]_  ? \new_[3489]_  : \new_[1816]_ ;
  assign \new_[1766]_  = \new_[477]_  ? \new_[3489]_  : \new_[1817]_ ;
  assign \new_[1767]_  = (~\new_[1818]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[452]_ );
  assign \new_[1768]_  = \new_[465]_  ? \new_[3489]_  : \new_[1819]_ ;
  assign \new_[1769]_  = (~\new_[1820]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[459]_ );
  assign \new_[1770]_  = \new_[476]_  ? \new_[3489]_  : \new_[1821]_ ;
  assign \new_[1771]_  = (~\new_[1822]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[505]_ );
  assign \new_[1772]_  = (~\new_[1823]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[448]_ );
  assign \new_[1773]_  = (~\new_[1865]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[456]_ );
  assign \new_[1774]_  = \new_[470]_  ? \new_[3489]_  : \new_[1872]_ ;
  assign \new_[1775]_  = ~\new_[1856]_  & ~\new_[1991]_ ;
  assign \new_[1776]_  = (~\new_[1912]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[466]_ );
  assign \new_[1777]_  = (~\new_[1863]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[475]_ );
  assign \new_[1778]_  = \new_[455]_  ? \new_[3489]_  : \new_[1864]_ ;
  assign \new_[1779]_  = ~\new_[1907]_  & ~\new_[1859]_ ;
  assign \new_[1780]_  = ~\new_[1860]_  & ~\new_[2167]_ ;
  assign \new_[1781]_  = \new_[1922]_  ? \new_[5307]_  : \new_[442]_ ;
  assign \new_[1782]_  = \new_[1923]_  ? \new_[5307]_  : \new_[492]_ ;
  assign \new_[1783]_  = \new_[1930]_  ? \new_[5307]_  : \new_[438]_ ;
  assign \new_[1784]_  = \new_[1929]_  ? \new_[5307]_  : \new_[4346]_ ;
  assign \new_[1785]_  = \new_[1924]_  ? \new_[5307]_  : \new_[4370]_ ;
  assign \new_[1786]_  = \new_[1932]_  ? \new_[5307]_  : \new_[463]_ ;
  assign \new_[1787]_  = \new_[1931]_  ? \new_[5307]_  : \new_[503]_ ;
  assign \new_[1788]_  = ~\new_[2081]_  | ~\new_[2084]_  | ~\new_[2168]_  | ~\new_[2082]_ ;
  assign \new_[1789]_  = ~\new_[1959]_  & ~\new_[1871]_ ;
  assign \new_[1790]_  = ~\new_[2079]_  & ~\new_[1867]_ ;
  assign \new_[1791]_  = ~\new_[2294]_  & ~\new_[1869]_ ;
  assign \new_[1792]_  = ~\new_[1868]_  & ~\new_[1958]_ ;
  assign \new_[1793]_  = ~\new_[1884]_  | ~\new_[2362]_ ;
  assign \new_[1794]_  = ~\new_[1882]_  | ~\new_[1883]_ ;
  assign \new_[1795]_  = ~\new_[1889]_  | ~\new_[1996]_ ;
  assign \new_[1796]_  = ~\new_[1949]_  & ~\new_[1876]_ ;
  assign \new_[1797]_  = ~\new_[1953]_  & ~\new_[1885]_ ;
  assign \new_[1798]_  = (~\new_[2030]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[446]_ );
  assign \new_[1799]_  = (~\new_[1913]_  | ~\new_[3489]_ ) & (~\new_[3754]_  | ~\new_[483]_ );
  assign \new_[1800]_  = ~\new_[2133]_  & ~\new_[1896]_ ;
  assign \new_[1801]_  = ~\new_[1906]_  & ~\new_[1967]_ ;
  assign \new_[1802]_  = ~\new_[2102]_  | ~\new_[1897]_ ;
  assign \new_[1803]_  = ~\new_[2003]_  & ~\new_[1895]_ ;
  assign \new_[1804]_  = \new_[2142]_  & \new_[1899]_ ;
  assign \new_[1805]_  = ~\new_[1908]_  & ~\new_[2118]_ ;
  assign \new_[1806]_  = ~\new_[1909]_  & ~\new_[1900]_ ;
  assign \new_[1807]_  = ~\new_[1986]_  & ~\new_[1901]_ ;
  assign \new_[1808]_  = ~\new_[1910]_  & ~\new_[1903]_ ;
  assign \new_[1809]_  = \new_[1928]_  ? \new_[5307]_  : \new_[454]_ ;
  assign \new_[1810]_  = \new_[1926]_  ? \new_[5307]_  : \new_[436]_ ;
  assign \new_[1811]_  = \new_[1925]_  ? \new_[5307]_  : \new_[474]_ ;
  assign \new_[1812]_  = \new_[1927]_  ? \new_[5307]_  : \new_[473]_ ;
  assign \new_[1813]_  = ~\new_[1915]_  & (~\new_[4313]_  | ~\new_[5307]_ );
  assign \new_[1814]_  = \new_[2065]_  ? \new_[5307]_  : \new_[472]_ ;
  assign \new_[1815]_  = \new_[2066]_  ? \new_[5307]_  : \new_[490]_ ;
  assign \new_[1816]_  = \new_[2067]_  ? \new_[5307]_  : \new_[434]_ ;
  assign \new_[1817]_  = \new_[2069]_  ? \new_[5307]_  : \new_[477]_ ;
  assign \new_[1818]_  = \new_[2070]_  ? \new_[5307]_  : \new_[452]_ ;
  assign \new_[1819]_  = \new_[2064]_  ? \new_[5307]_  : \new_[465]_ ;
  assign \new_[1820]_  = \new_[2068]_  ? \new_[5307]_  : \new_[459]_ ;
  assign \new_[1821]_  = \new_[2071]_  ? \new_[5307]_  : \new_[476]_ ;
  assign \new_[1822]_  = \new_[2073]_  ? \new_[5307]_  : \new_[505]_ ;
  assign \new_[1823]_  = \new_[2074]_  ? \new_[5307]_  : \new_[448]_ ;
  assign \new_[1824]_  = ~\new_[1933]_  & ~\new_[1936]_ ;
  assign \new_[1825]_  = ~\new_[1942]_  & ~\new_[1939]_ ;
  assign \new_[1826]_  = ~\new_[1943]_  & ~\new_[1944]_ ;
  assign \new_[1827]_  = ~\new_[1952]_  & ~\new_[1951]_ ;
  assign \new_[1828]_  = \new_[2077]_  ? \new_[5307]_  : \new_[440]_ ;
  assign \new_[1829]_  = \new_[2076]_  ? \new_[5307]_  : \new_[494]_ ;
  assign \new_[1830]_  = ~\new_[1947]_  & ~\new_[1948]_ ;
  assign \new_[1831]_  = ~\new_[2287]_  & ~\new_[1950]_ ;
  assign \new_[1832]_  = ~\new_[1954]_  & ~\new_[1955]_ ;
  assign \new_[1833]_  = \new_[1999]_  & \new_[1961]_ ;
  assign \new_[1834]_  = \new_[2035]_  & \new_[2015]_ ;
  assign \new_[1835]_  = ~\new_[2000]_  & (~\new_[2550]_  | ~\new_[4226]_ );
  assign \new_[1836]_  = ~\new_[2043]_  | ~\new_[2088]_  | ~\new_[2380]_ ;
  assign \new_[1837]_  = ~\new_[2002]_  | ~\new_[1965]_ ;
  assign \new_[1838]_  = \new_[2005]_  & \new_[1966]_ ;
  assign \new_[1839]_  = ~\new_[2127]_  & ~\new_[1969]_ ;
  assign \new_[1840]_  = ~\new_[1971]_  | ~\new_[2099]_ ;
  assign \new_[1841]_  = \new_[2004]_  & \new_[2298]_ ;
  assign \new_[1842]_  = ~\new_[2119]_  | ~\new_[2234]_  | ~\new_[2032]_ ;
  assign \new_[1843]_  = ~\new_[1981]_  | ~\new_[2315]_ ;
  assign \new_[1844]_  = ~\new_[2136]_  | ~\new_[1975]_ ;
  assign \new_[1845]_  = ~\new_[2006]_  & ~\new_[1976]_ ;
  assign \new_[1846]_  = ~\new_[2007]_  & ~\new_[1977]_ ;
  assign \new_[1847]_  = \new_[2096]_  & \new_[1973]_ ;
  assign \new_[1848]_  = ~\new_[2008]_  | ~\new_[2116]_ ;
  assign \new_[1849]_  = ~\new_[2413]_  | ~\new_[1984]_  | ~\new_[2917]_ ;
  assign \new_[1850]_  = ~\new_[2010]_  & ~\new_[2147]_ ;
  assign \new_[1851]_  = ~\new_[2144]_  | ~\new_[1985]_ ;
  assign \new_[1852]_  = ~\new_[1989]_  & ~\new_[1990]_ ;
  assign \new_[1853]_  = ~\new_[2013]_  & ~\new_[1995]_ ;
  assign \new_[1854]_  = \new_[2014]_  & \new_[2249]_ ;
  assign \new_[1855]_  = ~\new_[2420]_  | ~\new_[1997]_  | ~\new_[2654]_ ;
  assign \new_[1856]_  = ~\new_[2378]_  | ~\new_[2017]_ ;
  assign \new_[1857]_  = ~\new_[1917]_  & (~\new_[2771]_  | ~\new_[4102]_ );
  assign \new_[1858]_  = \new_[1918]_  & \new_[2213]_ ;
  assign \new_[1859]_  = ~\new_[2244]_  | ~\new_[1919]_ ;
  assign \new_[1860]_  = ~\new_[2205]_  | ~\new_[1920]_ ;
  assign \new_[1861]_  = \new_[1921]_  & \new_[2268]_ ;
  assign \new_[1862]_  = \new_[2887]_  & \new_[1916]_ ;
  assign \new_[1863]_  = \new_[2269]_  ? \new_[5307]_  : \new_[475]_ ;
  assign \new_[1864]_  = \new_[2271]_  ? \new_[5307]_  : \new_[455]_ ;
  assign \new_[1865]_  = \new_[2295]_  ? \new_[5307]_  : \new_[456]_ ;
  assign \new_[1866]_  = ~\new_[2616]_  | ~\new_[2078]_ ;
  assign \new_[1867]_  = ~\new_[2982]_  | ~\new_[2600]_  | ~\new_[2214]_ ;
  assign \new_[1868]_  = ~\new_[2085]_  | ~\new_[2374]_ ;
  assign \new_[1869]_  = ~\new_[2301]_  | ~\new_[2877]_  | ~\new_[2858]_ ;
  assign \new_[1870]_  = ~\new_[2717]_  | ~\new_[2080]_  | ~\new_[2418]_ ;
  assign \new_[1871]_  = ~\new_[2296]_  | ~\new_[2083]_ ;
  assign \new_[1872]_  = \new_[2169]_  ? \new_[5307]_  : \new_[470]_ ;
  assign \new_[1873]_  = ~\new_[2406]_  | ~\new_[2091]_  | ~\new_[2645]_ ;
  assign \new_[1874]_  = ~\new_[2097]_  & ~\new_[2120]_ ;
  assign \new_[1875]_  = ~\new_[2093]_  & ~\new_[2092]_ ;
  assign \new_[1876]_  = ~\new_[2398]_  | ~\new_[2328]_  | ~\new_[2174]_ ;
  assign \new_[1877]_  = ~\new_[2139]_  & ~\new_[2108]_ ;
  assign \new_[1878]_  = ~\new_[2140]_  & ~\new_[2114]_ ;
  assign \new_[1879]_  = ~\new_[2331]_  | ~\new_[2111]_ ;
  assign \new_[1880]_  = ~\new_[2333]_  | ~\new_[2112]_ ;
  assign \new_[1881]_  = ~\new_[2141]_  | ~\new_[2113]_ ;
  assign \new_[1882]_  = ~\new_[2151]_  & (~\new_[2782]_  | ~\new_[4074]_ );
  assign \new_[1883]_  = ~\new_[2152]_  & (~\new_[2281]_  | ~\new_[4065]_ );
  assign \new_[1884]_  = ~\new_[2150]_  & (~\new_[2181]_  | ~\new_[4214]_ );
  assign \new_[1885]_  = ~\new_[2388]_  | ~\new_[2341]_  | ~\new_[2177]_ ;
  assign \new_[1886]_  = ~\new_[2143]_  & ~\new_[2361]_ ;
  assign \new_[1887]_  = ~\new_[2371]_  & ~\new_[2123]_ ;
  assign \new_[1888]_  = ~\new_[2130]_  & ~\new_[2131]_ ;
  assign \new_[1889]_  = ~\new_[2033]_  & (~\new_[5271]_  | ~\new_[4098]_ );
  assign \new_[1890]_  = \new_[2264]_  & \new_[2042]_ ;
  assign \new_[1891]_  = ~\new_[2193]_  & (~\new_[2275]_  | ~\new_[4214]_ );
  assign \new_[1892]_  = ~\new_[2037]_  & (~\new_[2793]_  | ~\new_[4116]_ );
  assign \new_[1893]_  = ~\new_[2046]_  | ~\new_[2055]_ ;
  assign \new_[1894]_  = ~\new_[2191]_  | ~\new_[2036]_ ;
  assign \new_[1895]_  = ~\new_[2223]_  | ~\new_[2044]_ ;
  assign \new_[1896]_  = ~\new_[2038]_  | ~\new_[2492]_ ;
  assign \new_[1897]_  = ~\new_[2215]_  & (~\new_[2277]_  | ~\new_[5068]_ );
  assign \new_[1898]_  = ~\new_[2516]_  & (~\new_[2278]_  | ~\new_[4121]_ );
  assign \new_[1899]_  = ~\new_[2052]_  & (~\new_[2820]_  | ~\new_[4226]_ );
  assign \new_[1900]_  = ~\new_[2259]_  | ~\new_[2059]_ ;
  assign \new_[1901]_  = ~\new_[2060]_  | ~\new_[2260]_ ;
  assign \new_[1902]_  = \new_[2061]_  | \new_[2589]_ ;
  assign \new_[1903]_  = \new_[2534]_  | \new_[2063]_ ;
  assign \new_[1904]_  = ~\new_[2045]_  & (~\new_[3366]_  | ~\new_[4069]_ );
  assign \new_[1905]_  = ~\new_[2637]_  | ~\new_[2054]_ ;
  assign \new_[1906]_  = ~\new_[2893]_  | ~\new_[2047]_ ;
  assign \new_[1907]_  = ~\new_[2175]_  | ~\new_[2051]_ ;
  assign \new_[1908]_  = ~\new_[2041]_  | ~\new_[2409]_ ;
  assign \new_[1909]_  = ~\new_[2415]_  | ~\new_[2058]_ ;
  assign \new_[1910]_  = ~\new_[2650]_  | ~\new_[2062]_ ;
  assign \new_[1911]_  = ~\new_[2029]_ ;
  assign \new_[1912]_  = \new_[2270]_  ? \new_[5307]_  : \new_[466]_ ;
  assign \new_[1913]_  = \new_[2547]_  ? \new_[5307]_  : \new_[483]_ ;
  assign \new_[1914]_  = (~\new_[2827]_  | ~\new_[4069]_ ) & (~\new_[2581]_  | ~\new_[4222]_ );
  assign \new_[1915]_  = ~\new_[2272]_  & ~\new_[5307]_ ;
  assign \new_[1916]_  = ~\new_[2034]_ ;
  assign \new_[1917]_  = ~\new_[4197]_  & (~\new_[2961]_  | ~\new_[3433]_ );
  assign \new_[1918]_  = ~\new_[2273]_  | ~\new_[4214]_ ;
  assign \new_[1919]_  = ~\new_[2283]_  | ~\new_[4240]_ ;
  assign \new_[1920]_  = ~\new_[2280]_  | ~\new_[4121]_ ;
  assign \new_[1921]_  = ~\new_[2279]_  | ~\new_[4047]_ ;
  assign \new_[1922]_  = \\L_reg[15] ;
  assign \new_[1923]_  = \\L_reg[23] ;
  assign \new_[1924]_  = \\L_reg[30] ;
  assign \new_[1925]_  = \\L_reg[19] ;
  assign \new_[1926]_  = \\L_reg[11] ;
  assign \new_[1927]_  = \\L_reg[27] ;
  assign \new_[1928]_  = \\L_reg[28] ;
  assign \new_[1929]_  = \\L_reg[17] ;
  assign \new_[1930]_  = \\L_reg[3] ;
  assign \new_[1931]_  = \\L_reg[24] ;
  assign \new_[1932]_  = \\L_reg[31] ;
  assign \new_[1933]_  = ~\new_[2621]_  | ~\new_[2303]_ ;
  assign \new_[1934]_  = ~\new_[2360]_  | ~\new_[2607]_ ;
  assign \new_[1935]_  = ~\new_[2659]_  | ~\new_[2304]_  | ~\new_[2901]_ ;
  assign \new_[1936]_  = ~\new_[2340]_  | ~\new_[2318]_ ;
  assign \new_[1937]_  = ~\new_[2524]_  | ~\new_[2335]_  | ~\new_[2383]_ ;
  assign \new_[1938]_  = ~\new_[2894]_  | ~\new_[2306]_  | ~\new_[2636]_ ;
  assign \new_[1939]_  = ~\new_[2605]_  | ~\new_[2312]_ ;
  assign \new_[1940]_  = ~\new_[2363]_  | ~\new_[2862]_ ;
  assign \new_[1941]_  = ~\new_[2900]_  | ~\new_[2311]_  | ~\new_[2395]_ ;
  assign \new_[1942]_  = ~\new_[2337]_  | ~\new_[2313]_ ;
  assign \new_[1943]_  = ~\new_[2336]_  | ~\new_[2609]_ ;
  assign \new_[1944]_  = ~\new_[2320]_  | ~\new_[2863]_ ;
  assign \new_[1945]_  = ~\new_[2364]_  | ~\new_[2321]_ ;
  assign \new_[1946]_  = ~\new_[2322]_  | ~\new_[2323]_ ;
  assign \new_[1947]_  = ~\new_[2504]_  | ~\new_[2326]_  | ~\new_[2396]_ ;
  assign \new_[1948]_  = ~\new_[2400]_  | ~\new_[2327]_  | ~\new_[2399]_ ;
  assign \new_[1949]_  = ~\new_[2365]_  | ~\new_[2325]_ ;
  assign \new_[1950]_  = ~\new_[2909]_  | ~\new_[2402]_  | ~\new_[2329]_ ;
  assign \new_[1951]_  = ~\new_[2316]_  | ~\new_[2300]_ ;
  assign \new_[1952]_  = ~\new_[2314]_  | ~\new_[2611]_ ;
  assign \new_[1953]_  = ~\new_[2368]_  | ~\new_[2339]_ ;
  assign \new_[1954]_  = ~\new_[2372]_  | ~\new_[2349]_ ;
  assign \new_[1955]_  = ~\new_[2920]_  | ~\new_[2350]_  | ~\new_[2919]_ ;
  assign \new_[1956]_  = ~\new_[2615]_  | ~\new_[2351]_ ;
  assign \new_[1957]_  = ~\new_[2624]_  & ~\new_[2352]_ ;
  assign \new_[1958]_  = ~\new_[2375]_  | ~\new_[2358]_ ;
  assign \new_[1959]_  = ~\new_[2606]_  | ~\new_[2359]_ ;
  assign \new_[1960]_  = ~\new_[2656]_  & (~\new_[2583]_  | ~\new_[4116]_ );
  assign \new_[1961]_  = ~\new_[2212]_  & (~\new_[2773]_  | ~\new_[4122]_ );
  assign \new_[1962]_  = ~\new_[2225]_  & (~\new_[2838]_  | ~\new_[4170]_ );
  assign \new_[1963]_  = ~\new_[2944]_  & (~\new_[2582]_  | ~\new_[4256]_ );
  assign \new_[1964]_  = ~\new_[2186]_  | ~\new_[2466]_ ;
  assign \new_[1965]_  = ~\new_[2540]_  & (~\new_[2591]_  | ~\new_[5097]_ );
  assign \new_[1966]_  = ~\new_[2219]_  & (~\new_[2800]_  | ~\new_[4102]_ );
  assign \new_[1967]_  = \new_[2476]_  | \new_[2220]_ ;
  assign \new_[1968]_  = \new_[2221]_  & \new_[2189]_ ;
  assign \new_[1969]_  = ~\new_[2222]_  | ~\new_[2482]_ ;
  assign \new_[1970]_  = ~\new_[2187]_  & (~\new_[3053]_  | ~\new_[4166]_ );
  assign \new_[1971]_  = ~\new_[2248]_  & (~\new_[2558]_  | ~\new_[4074]_ );
  assign \new_[1972]_  = \new_[2252]_  & \new_[2243]_ ;
  assign \new_[1973]_  = ~\new_[2227]_  & (~\new_[2556]_  | ~\new_[4069]_ );
  assign \new_[1974]_  = \new_[2254]_  & \new_[2437]_ ;
  assign \new_[1975]_  = ~\new_[2722]_  & (~\new_[2579]_  | ~\new_[4122]_ );
  assign \new_[1976]_  = ~\new_[2196]_  | ~\new_[2233]_ ;
  assign \new_[1977]_  = ~\new_[2199]_  | ~\new_[2235]_ ;
  assign \new_[1978]_  = ~\new_[2204]_  & (~\new_[2575]_  | ~\new_[4074]_ );
  assign \new_[1979]_  = \new_[2206]_  & \new_[2250]_ ;
  assign \new_[1980]_  = \new_[2224]_  & \new_[2195]_ ;
  assign \new_[1981]_  = ~\new_[2185]_  & (~\new_[2567]_  | ~\new_[4108]_ );
  assign \new_[1982]_  = ~\new_[2255]_  | ~\new_[2490]_ ;
  assign \new_[1983]_  = ~\new_[2544]_  & (~\new_[2584]_  | ~\new_[4245]_ );
  assign \new_[1984]_  = ~\new_[2530]_  & (~\new_[2586]_  | ~\new_[5097]_ );
  assign \new_[1985]_  = ~\new_[2258]_  & (~\new_[2814]_  | ~\new_[4023]_ );
  assign \new_[1986]_  = ~\new_[2436]_  | ~\new_[2208]_ ;
  assign \new_[1987]_  = ~\new_[2754]_  & (~\new_[2588]_  | ~\new_[4125]_ );
  assign \new_[1988]_  = ~\new_[2266]_  & (~\new_[2845]_  | ~\new_[4226]_ );
  assign \new_[1989]_  = \new_[2535]_  | \new_[2262]_ ;
  assign \new_[1990]_  = \new_[2682]_  | \new_[2209]_ ;
  assign \new_[1991]_  = ~\new_[2687]_  | ~\new_[2232]_ ;
  assign \new_[1992]_  = ~\new_[2766]_  & (~\new_[2592]_  | ~\new_[4116]_ );
  assign \new_[1993]_  = ~\new_[2183]_  & (~\new_[2555]_  | ~\new_[4245]_ );
  assign \new_[1994]_  = ~\new_[2767]_  & (~\new_[2622]_  | ~\new_[4222]_ );
  assign \new_[1995]_  = \new_[2210]_  | \new_[2545]_ ;
  assign \new_[1996]_  = ~\new_[2768]_  & (~\new_[2570]_  | ~\new_[4240]_ );
  assign \new_[1997]_  = ~\new_[2267]_  & (~\new_[3145]_  | ~\new_[5097]_ );
  assign \new_[1998]_  = ~\new_[2216]_  & (~\new_[2705]_  | ~\new_[4220]_ );
  assign \new_[1999]_  = ~\new_[2211]_  & (~\new_[3345]_  | ~\new_[4222]_ );
  assign \new_[2000]_  = ~\new_[4143]_  & (~\new_[3165]_  | ~\new_[2772]_ );
  assign \new_[2001]_  = ~\new_[2171]_  | ~\new_[2253]_ ;
  assign \new_[2002]_  = ~\new_[2251]_  & (~\new_[3334]_  | ~\new_[4021]_ );
  assign \new_[2003]_  = ~\new_[2394]_  | ~\new_[2192]_ ;
  assign \new_[2004]_  = ~\new_[2464]_  & (~\new_[2578]_  | ~\new_[4098]_ );
  assign \new_[2005]_  = ~\new_[2228]_  & (~\new_[3012]_  | ~\new_[4220]_ );
  assign \new_[2006]_  = ~\new_[2173]_  | ~\new_[2231]_ ;
  assign \new_[2007]_  = ~\new_[2397]_  | ~\new_[2198]_ ;
  assign \new_[2008]_  = ~\new_[2245]_  & (~\new_[2578]_  | ~\new_[4220]_ );
  assign \new_[2009]_  = ~\new_[2178]_  | ~\new_[2527]_ ;
  assign \new_[2010]_  = ~\new_[2414]_  | ~\new_[2261]_ ;
  assign \new_[2011]_  = ~\new_[2218]_  & (~\new_[3248]_  | ~\new_[4098]_ );
  assign \new_[2012]_  = ~\new_[2263]_  & (~\new_[3476]_  | ~\new_[4069]_ );
  assign \new_[2013]_  = ~\new_[2632]_  | ~\new_[2265]_ ;
  assign \new_[2014]_  = ~\new_[2148]_ ;
  assign \new_[2015]_  = ~\new_[2170]_  | ~\new_[4065]_ ;
  assign \new_[2016]_  = \\FP_R_reg[49] ;
  assign \new_[2017]_  = ~\new_[2182]_  | ~\new_[5068]_ ;
  assign \new_[2018]_  = \\FP_R_reg[35] ;
  assign \new_[2019]_  = \\FP_R_reg[56] ;
  assign \new_[2020]_  = \\FP_R_reg[55] ;
  assign \new_[2021]_  = \\FP_R_reg[62] ;
  assign \new_[2022]_  = \\FP_R_reg[47] ;
  assign \new_[2023]_  = \\FP_R_reg[60] ;
  assign \new_[2024]_  = \\FP_R_reg[59] ;
  assign \new_[2025]_  = \\FP_R_reg[43] ;
  assign \new_[2026]_  = \\FP_R_reg[51] ;
  assign \new_[2027]_  = \\FP_R_reg[63] ;
  assign \new_[2028]_  = ~\new_[2176]_  & (~\new_[2581]_  | ~\new_[4069]_ );
  assign \new_[2029]_  = ~\new_[2179]_  | ~\new_[2180]_ ;
  assign \new_[2030]_  = \new_[2546]_  ? \new_[5307]_  : \new_[446]_ ;
  assign \new_[2031]_  = \\FP_R_reg[64] ;
  assign \new_[2032]_  = ~\new_[5270]_  | ~\new_[4220]_ ;
  assign \new_[2033]_  = ~\new_[4104]_  & (~\new_[3255]_  | ~\new_[2772]_ );
  assign \new_[2034]_  = ~\new_[4203]_  & (~\new_[3277]_  | ~\new_[3564]_ );
  assign \new_[2035]_  = ~\new_[2184]_ ;
  assign \new_[2036]_  = ~\new_[2561]_  | ~\new_[4158]_ ;
  assign \new_[2037]_  = ~\new_[5174]_  & (~\new_[3186]_  | ~\new_[3488]_ );
  assign \new_[2038]_  = ~\new_[2563]_  | ~\new_[4212]_ ;
  assign \new_[2039]_  = ~\new_[2553]_  | ~\new_[4208]_ ;
  assign \new_[2040]_  = ~\new_[2203]_ ;
  assign \new_[2041]_  = ~\new_[2554]_  | ~\new_[4174]_ ;
  assign \new_[2042]_  = ~\new_[2549]_  | ~\new_[4047]_ ;
  assign \new_[2043]_  = ~\new_[2552]_  | ~\new_[4226]_ ;
  assign \new_[2044]_  = ~\new_[2566]_  | ~\new_[4240]_ ;
  assign \new_[2045]_  = ~\new_[4189]_  & (~\new_[3402]_  | ~\new_[5178]_ );
  assign \new_[2046]_  = ~\new_[2557]_  | ~\new_[4108]_ ;
  assign \new_[2047]_  = ~\new_[2564]_  | ~\new_[4121]_ ;
  assign \new_[2048]_  = ~\new_[2571]_  | ~\new_[4176]_ ;
  assign \new_[2049]_  = ~\new_[2585]_  | ~\new_[4226]_ ;
  assign \new_[2050]_  = ~\new_[2574]_  | ~\new_[5068]_ ;
  assign \new_[2051]_  = ~\new_[2577]_  | ~\new_[4023]_ ;
  assign \new_[2052]_  = ~\new_[4184]_  & (~\new_[3277]_  | ~\new_[3314]_ );
  assign \new_[2053]_  = ~\new_[4085]_  & (~\new_[3186]_  | ~\new_[3264]_ );
  assign \new_[2054]_  = ~\new_[2569]_  | ~\new_[4200]_ ;
  assign \new_[2055]_  = ~\new_[2560]_  | ~\new_[5068]_ ;
  assign \new_[2056]_  = ~\new_[2551]_  | ~\new_[4214]_ ;
  assign \new_[2057]_  = ~\new_[2593]_  | ~\new_[4170]_ ;
  assign \new_[2058]_  = ~\new_[2587]_  | ~\new_[4256]_ ;
  assign \new_[2059]_  = ~\new_[2576]_  | ~\new_[5068]_ ;
  assign \new_[2060]_  = ~\new_[2559]_  | ~\new_[4125]_ ;
  assign \new_[2061]_  = ~\new_[4189]_  & (~\new_[3309]_  | ~\new_[2880]_ );
  assign \new_[2062]_  = ~\new_[2610]_  | ~\new_[4214]_ ;
  assign \new_[2063]_  = \new_[2590]_  & \new_[4065]_ ;
  assign \new_[2064]_  = \\L_reg[8] ;
  assign \new_[2065]_  = \\L_reg[26] ;
  assign \new_[2066]_  = \\L_reg[32] ;
  assign \new_[2067]_  = \\L_reg[25] ;
  assign \new_[2068]_  = \\L_reg[13] ;
  assign \new_[2069]_  = \\L_reg[6] ;
  assign \new_[2070]_  = \\L_reg[5] ;
  assign \new_[2071]_  = \\L_reg[21] ;
  assign \new_[2072]_  = ~\new_[2734]_  | ~\new_[2866]_  | ~\new_[2865]_ ;
  assign \new_[2073]_  = \\L_reg[16] ;
  assign \new_[2074]_  = \\L_reg[22] ;
  assign \new_[2075]_  = ~\new_[2433]_  | ~\new_[2884]_ ;
  assign \new_[2076]_  = \\L_reg[1] ;
  assign \new_[2077]_  = \\L_reg[7] ;
  assign \new_[2078]_  = ~\new_[3190]_  & (~\new_[2651]_  | ~\new_[5099]_ );
  assign \new_[2079]_  = ~\new_[3179]_  | ~\new_[2874]_  | ~\new_[2761]_ ;
  assign \new_[2080]_  = ~\new_[2627]_  & (~\new_[2959]_  | ~\new_[4793]_ );
  assign \new_[2081]_  = ~\new_[2625]_  & ~\new_[2618]_ ;
  assign \new_[2082]_  = ~\new_[2619]_  & ~\new_[2620]_ ;
  assign \new_[2083]_  = ~\new_[2928]_  & ~\new_[2630]_ ;
  assign \new_[2084]_  = ~\new_[2628]_  & (~\new_[3392]_  | ~\new_[5097]_ );
  assign \new_[2085]_  = ~\new_[2626]_  & (~\new_[3037]_  | ~\new_[4131]_ );
  assign \new_[2086]_  = ~\new_[2421]_  & (~\new_[2824]_  | ~\new_[4121]_ );
  assign \new_[2087]_  = ~\new_[2493]_  & (~\new_[2825]_  | ~\new_[4170]_ );
  assign \new_[2088]_  = ~\new_[2658]_  & ~\new_[2467]_ ;
  assign \new_[2089]_  = ~\new_[2675]_  | ~\new_[2471]_ ;
  assign \new_[2090]_  = ~\new_[2472]_  | ~\new_[2423]_ ;
  assign \new_[2091]_  = ~\new_[2424]_  & ~\new_[2698]_ ;
  assign \new_[2092]_  = ~\new_[2488]_  | ~\new_[2519]_ ;
  assign \new_[2093]_  = ~\new_[2434]_  | ~\new_[2541]_ ;
  assign \new_[2094]_  = ~\new_[2712]_  | ~\new_[2430]_ ;
  assign \new_[2095]_  = ~\new_[2713]_  | ~\new_[2483]_ ;
  assign \new_[2096]_  = ~\new_[2487]_  & (~\new_[2826]_  | ~\new_[4023]_ );
  assign \new_[2097]_  = ~\new_[2665]_  | ~\new_[2525]_ ;
  assign \new_[2098]_  = ~\new_[2696]_  | ~\new_[2470]_ ;
  assign \new_[2099]_  = ~\new_[2885]_  & (~\new_[2819]_  | ~\new_[4250]_ );
  assign \new_[2100]_  = ~\new_[2491]_  & (~\new_[3068]_  | ~\new_[4166]_ );
  assign \new_[2101]_  = ~\new_[2431]_  & (~\new_[2993]_  | ~\new_[4232]_ );
  assign \new_[2102]_  = ~\new_[2748]_  & ~\new_[2522]_ ;
  assign \new_[2103]_  = ~\new_[2440]_  | ~\new_[2439]_ ;
  assign \new_[2104]_  = ~\new_[2444]_  & (~\new_[2834]_  | ~\new_[4108]_ );
  assign \new_[2105]_  = ~\new_[2503]_  | ~\new_[2509]_ ;
  assign \new_[2106]_  = ~\new_[2958]_  & (~\new_[2794]_  | ~\new_[4232]_ );
  assign \new_[2107]_  = ~\new_[2506]_  & (~\new_[3082]_  | ~\new_[5068]_ );
  assign \new_[2108]_  = ~\new_[2445]_  | ~\new_[2507]_ ;
  assign \new_[2109]_  = ~\new_[2508]_  & (~\new_[2812]_  | ~\new_[4209]_ );
  assign \new_[2110]_  = ~\new_[2510]_  & (~\new_[2813]_  | ~\new_[4233]_ );
  assign \new_[2111]_  = ~\new_[2673]_  & (~\new_[2816]_  | ~\new_[5068]_ );
  assign \new_[2112]_  = ~\new_[2447]_  & (~\new_[3122]_  | ~\new_[4237]_ );
  assign \new_[2113]_  = ~\new_[2448]_  & (~\new_[3133]_  | ~\new_[4226]_ );
  assign \new_[2114]_  = ~\new_[2933]_  | ~\new_[2523]_ ;
  assign \new_[2115]_  = \new_[2520]_  | \new_[2521]_ ;
  assign \new_[2116]_  = ~\new_[2450]_  & (~\new_[2832]_  | ~\new_[5068]_ );
  assign \new_[2117]_  = ~\new_[2644]_  & (~\new_[2796]_  | ~\new_[5068]_ );
  assign \new_[2118]_  = ~\new_[2454]_  | ~\new_[2526]_ ;
  assign \new_[2119]_  = ~\new_[2975]_  & (~\new_[2777]_  | ~\new_[4109]_ );
  assign \new_[2120]_  = ~\new_[2486]_  | ~\new_[2484]_ ;
  assign \new_[2121]_  = ~\new_[2529]_  & (~\new_[3169]_  | ~\new_[4239]_ );
  assign \new_[2122]_  = ~\new_[2532]_  | ~\new_[2463]_ ;
  assign \new_[2123]_  = ~\new_[2458]_  | ~\new_[2459]_ ;
  assign \new_[2124]_  = ~\new_[2757]_  & (~\new_[2804]_  | ~\new_[4214]_ );
  assign \new_[2125]_  = ~\new_[2536]_  | ~\new_[2537]_ ;
  assign \new_[2126]_  = ~\new_[2538]_  | ~\new_[2937]_ ;
  assign \new_[2127]_  = ~\new_[2461]_  | ~\new_[2662]_ ;
  assign \new_[2128]_  = ~\new_[2485]_  | ~\new_[2432]_ ;
  assign \new_[2129]_  = ~\new_[2462]_  | ~\new_[2542]_ ;
  assign \new_[2130]_  = ~\new_[2452]_  | ~\new_[2743]_ ;
  assign \new_[2131]_  = ~\new_[2543]_  | ~\new_[2438]_ ;
  assign \new_[2132]_  = ~\new_[2477]_  & (~\new_[2997]_  | ~\new_[4122]_ );
  assign \new_[2133]_  = ~\new_[2389]_  | ~\new_[2480]_ ;
  assign \new_[2134]_  = ~\new_[2390]_  | ~\new_[2962]_ ;
  assign \new_[2135]_  = ~\new_[2635]_  | ~\new_[2518]_ ;
  assign \new_[2136]_  = ~\new_[2441]_  & (~\new_[3233]_  | ~\new_[4222]_ );
  assign \new_[2137]_  = ~\new_[2641]_  | ~\new_[2495]_ ;
  assign \new_[2138]_  = ~\new_[2906]_  | ~\new_[2502]_ ;
  assign \new_[2139]_  = ~\new_[2401]_  | ~\new_[2716]_ ;
  assign \new_[2140]_  = ~\new_[2403]_  | ~\new_[2449]_ ;
  assign \new_[2141]_  = ~\new_[2515]_  & (~\new_[3137]_  | ~\new_[4069]_ );
  assign \new_[2142]_  = ~\new_[2740]_  & (~\new_[2827]_  | ~\new_[4222]_ );
  assign \new_[2143]_  = ~\new_[2646]_  | ~\new_[2494]_ ;
  assign \new_[2144]_  = ~\new_[2457]_  & (~\new_[3006]_  | ~\new_[4222]_ );
  assign \new_[2145]_  = ~\new_[2460]_  & (~\new_[3126]_  | ~\new_[4222]_ );
  assign \new_[2146]_  = ~\new_[2896]_  | ~\new_[2429]_ ;
  assign \new_[2147]_  = ~\new_[2416]_  | ~\new_[2505]_ ;
  assign \new_[2148]_  = ~\new_[4203]_  & (~\new_[2779]_  | ~\new_[3151]_ );
  assign \new_[2149]_  = ~\new_[4177]_  & (~\new_[3646]_  | ~\new_[2779]_ );
  assign \new_[2150]_  = ~\new_[4169]_  & (~\new_[3316]_  | ~\new_[2779]_ );
  assign \new_[2151]_  = ~\new_[4169]_  & (~\new_[2772]_  | ~\new_[3270]_ );
  assign \new_[2152]_  = ~\new_[4197]_  & (~\new_[2779]_  | ~\new_[3404]_ );
  assign \new_[2153]_  = \\FP_R_reg[58] ;
  assign \new_[2154]_  = \\FP_R_reg[54] ;
  assign \new_[2155]_  = \\FP_R_reg[53] ;
  assign \new_[2156]_  = \\FP_R_reg[40] ;
  assign \new_[2157]_  = \\FP_R_reg[38] ;
  assign \new_[2158]_  = \\FP_R_reg[37] ;
  assign \new_[2159]_  = \\FP_R_reg[45] ;
  assign \new_[2160]_  = \\FP_R_reg[57] ;
  assign \new_[2161]_  = \\FP_R_reg[48] ;
  assign \new_[2162]_  = \\FP_R_reg[33] ;
  assign \new_[2163]_  = \\FP_R_reg[39] ;
  assign \new_[2164]_  = \new_[2895]_  & \new_[2385]_ ;
  assign \new_[2165]_  = \new_[2914]_  & \new_[2386]_ ;
  assign \new_[2166]_  = (~\new_[3095]_  | ~\new_[4098]_ ) & (~\new_[2821]_  | ~\new_[4222]_ );
  assign \new_[2167]_  = ~\new_[2407]_  | ~\new_[2408]_ ;
  assign \new_[2168]_  = ~\new_[2377]_ ;
  assign \new_[2169]_  = \\L_reg[12] ;
  assign \new_[2170]_  = ~\new_[2779]_  | ~\new_[3278]_ ;
  assign \new_[2171]_  = ~\new_[2783]_  | ~\new_[4220]_ ;
  assign \new_[2172]_  = ~\new_[2778]_  | ~\new_[4222]_ ;
  assign \new_[2173]_  = ~\new_[2776]_  | ~\new_[4220]_ ;
  assign \new_[2174]_  = ~\new_[2811]_  | ~\new_[4242]_ ;
  assign \new_[2175]_  = ~\new_[2776]_  | ~\new_[4098]_ ;
  assign \new_[2176]_  = \new_[2705]_  & \new_[4098]_ ;
  assign \new_[2177]_  = ~\new_[2821]_  | ~\new_[4176]_ ;
  assign \new_[2178]_  = ~\new_[2811]_  | ~\new_[4698]_ ;
  assign \new_[2179]_  = ~\new_[2783]_  | ~\new_[4098]_ ;
  assign \new_[2180]_  = ~\new_[2778]_  | ~\new_[4069]_ ;
  assign \new_[2181]_  = ~\new_[3277]_  | ~\new_[3216]_ ;
  assign \new_[2182]_  = ~\new_[3498]_  | ~\new_[2779]_ ;
  assign \new_[2183]_  = ~\new_[5098]_  & (~\new_[3488]_  | ~\new_[3273]_ );
  assign \new_[2184]_  = ~\new_[5174]_  & (~\new_[3587]_  | ~\new_[3314]_ );
  assign \new_[2185]_  = ~\new_[5174]_  & (~\new_[3316]_  | ~\new_[3433]_ );
  assign \new_[2186]_  = ~\new_[2810]_  | ~\new_[4074]_ ;
  assign \new_[2187]_  = ~\new_[4163]_  & (~\new_[3281]_  | ~\new_[2978]_ );
  assign \new_[2188]_  = ~\new_[2799]_  | ~\new_[4158]_ ;
  assign \new_[2189]_  = ~\new_[2427]_ ;
  assign \new_[2190]_  = ~\new_[4269]_  & (~\new_[3152]_  | ~\new_[3479]_ );
  assign \new_[2191]_  = ~\new_[2787]_  | ~\new_[4250]_ ;
  assign \new_[2192]_  = ~\new_[2784]_  | ~\new_[5097]_ ;
  assign \new_[2193]_  = ~\new_[4203]_  & (~\new_[3310]_  | ~\new_[3309]_ );
  assign \new_[2194]_  = \\FP_R_reg[52] ;
  assign \new_[2195]_  = ~\new_[2435]_ ;
  assign \new_[2196]_  = ~\new_[2803]_  | ~\new_[4158]_ ;
  assign \new_[2197]_  = ~\new_[4269]_  & (~\new_[3421]_  | ~\new_[3426]_ );
  assign \new_[2198]_  = ~\new_[2806]_  | ~\new_[4241]_ ;
  assign \new_[2199]_  = ~\new_[2808]_  | ~\new_[4199]_ ;
  assign \new_[2200]_  = ~\new_[2830]_  | ~\new_[5097]_ ;
  assign \new_[2201]_  = ~\new_[2446]_ ;
  assign \new_[2202]_  = ~\new_[5098]_  & (~\new_[3155]_  | ~\new_[5241]_ );
  assign \new_[2203]_  = ~\new_[4192]_  & (~\new_[4380]_  | ~\new_[4385]_ );
  assign \new_[2204]_  = ~\new_[4203]_  & (~\new_[4790]_  | ~\new_[3170]_ );
  assign \new_[2205]_  = ~\new_[2829]_  | ~\new_[5097]_ ;
  assign \new_[2206]_  = ~\new_[2453]_ ;
  assign \new_[2207]_  = \\FP_R_reg[36] ;
  assign \new_[2208]_  = ~\new_[2844]_  | ~\new_[4199]_ ;
  assign \new_[2209]_  = ~\new_[5174]_  & (~\new_[4402]_  | ~\new_[2978]_ );
  assign \new_[2210]_  = ~\new_[5174]_  & (~\new_[3265]_  | ~\new_[3414]_ );
  assign \new_[2211]_  = ~\new_[3958]_  & (~\new_[3316]_  | ~\new_[3425]_ );
  assign \new_[2212]_  = ~\new_[4792]_  & (~\new_[3265]_  | ~\new_[3404]_ );
  assign \new_[2213]_  = ~\new_[2795]_  | ~\new_[5068]_ ;
  assign \new_[2214]_  = ~\new_[2652]_  | ~\new_[4239]_ ;
  assign \new_[2215]_  = ~\new_[4169]_  & (~\new_[3154]_  | ~\new_[3485]_ );
  assign \new_[2216]_  = ~\new_[4115]_  & (~\new_[3154]_  | ~\new_[3550]_ );
  assign \new_[2217]_  = \\FP_R_reg[42] ;
  assign \new_[2218]_  = ~\new_[4792]_  & (~\new_[3331]_  | ~\new_[5241]_ );
  assign \new_[2219]_  = ~\new_[5063]_  & (~\new_[3293]_  | ~\new_[2978]_ );
  assign \new_[2220]_  = ~\new_[4184]_  & (~\new_[4790]_  | ~\new_[3155]_ );
  assign \new_[2221]_  = ~\new_[2786]_  | ~\new_[4226]_ ;
  assign \new_[2222]_  = ~\new_[2797]_  | ~\new_[4176]_ ;
  assign \new_[2223]_  = ~\new_[2723]_  | ~\new_[4226]_ ;
  assign \new_[2224]_  = ~\new_[2775]_  | ~\new_[4121]_ ;
  assign \new_[2225]_  = ~\new_[4184]_  & (~\new_[5240]_  | ~\new_[3280]_ );
  assign \new_[2226]_  = ~n990;
  assign \new_[2227]_  = ~\new_[4168]_  & (~\new_[3153]_  | ~\new_[3199]_ );
  assign \new_[2228]_  = ~\new_[4115]_  & (~\new_[3275]_  | ~\new_[5241]_ );
  assign \new_[2229]_  = ~\new_[2846]_  | ~\new_[4133]_ ;
  assign \new_[2230]_  = ~\new_[2801]_  | ~\new_[4109]_ ;
  assign \new_[2231]_  = ~\new_[2802]_  | ~\new_[4228]_ ;
  assign \new_[2232]_  = ~\new_[2823]_  | ~\new_[4228]_ ;
  assign \new_[2233]_  = ~\new_[2839]_  | ~\new_[4214]_ ;
  assign \new_[2234]_  = ~\new_[2805]_  | ~\new_[5068]_ ;
  assign \new_[2235]_  = ~\new_[2809]_  | ~\new_[4237]_ ;
  assign \new_[2236]_  = ~\new_[4169]_  & (~\new_[3309]_  | ~\new_[3273]_ );
  assign \new_[2237]_  = ~\new_[4168]_  & (~\new_[3443]_  | ~\new_[3263]_ );
  assign n1030 = ~\new_[5194]_ ;
  assign \new_[2239]_  = ~\new_[2842]_  | ~\new_[4116]_ ;
  assign \new_[2240]_  = ~\new_[2788]_  | ~\new_[3985]_ ;
  assign \new_[2241]_  = ~\new_[2683]_  | ~\new_[4214]_ ;
  assign \new_[2242]_  = ~\new_[2833]_  | ~\new_[4170]_ ;
  assign \new_[2243]_  = ~\new_[2791]_  | ~\new_[4121]_ ;
  assign \new_[2244]_  = ~\new_[2836]_  | ~\new_[4226]_ ;
  assign \new_[2245]_  = ~\new_[4164]_  & (~\new_[3153]_  | ~\new_[3255]_ );
  assign \new_[2246]_  = ~\new_[4104]_  & (~\new_[3157]_  | ~\new_[3199]_ );
  assign \new_[2247]_  = \\FP_R_reg[34] ;
  assign \new_[2248]_  = ~\new_[4247]_  & (~\new_[3153]_  | ~\new_[3165]_ );
  assign \new_[2249]_  = ~\new_[2719]_  | ~\new_[4065]_ ;
  assign \new_[2250]_  = ~\new_[2835]_  | ~\new_[4121]_ ;
  assign \new_[2251]_  = ~\new_[4189]_  & (~\new_[3503]_  | ~\new_[3151]_ );
  assign \new_[2252]_  = ~\new_[2828]_  | ~\new_[4023]_ ;
  assign \new_[2253]_  = ~\new_[2837]_  | ~\new_[4108]_ ;
  assign \new_[2254]_  = ~\new_[2840]_  | ~\new_[4226]_ ;
  assign \new_[2255]_  = ~\new_[2770]_  | ~\new_[4232]_ ;
  assign \new_[2256]_  = ~\new_[4179]_  & (~\new_[3268]_  | ~\new_[3151]_ );
  assign \new_[2257]_  = ~\new_[2843]_  | ~\new_[5068]_ ;
  assign \new_[2258]_  = ~\new_[4792]_  & (~\new_[4405]_  | ~\new_[3443]_ );
  assign \new_[2259]_  = ~\new_[2785]_  | ~\new_[4108]_ ;
  assign \new_[2260]_  = ~\new_[2789]_  | ~\new_[4228]_ ;
  assign \new_[2261]_  = ~\new_[2781]_  | ~\new_[4160]_ ;
  assign \new_[2262]_  = ~\new_[5063]_  & (~\new_[5183]_  | ~\new_[3488]_ );
  assign \new_[2263]_  = ~\new_[3958]_  & (~\new_[3531]_  | ~\new_[3155]_ );
  assign \new_[2264]_  = ~\new_[2774]_  | ~\new_[3985]_ ;
  assign \new_[2265]_  = ~\new_[2847]_  | ~\new_[3985]_ ;
  assign \new_[2266]_  = ~\new_[4184]_  & (~\new_[3517]_  | ~\new_[2978]_ );
  assign \new_[2267]_  = ~\new_[4792]_  & (~\new_[3165]_  | ~\new_[3314]_ );
  assign \new_[2268]_  = ~\new_[2831]_  | ~\new_[4214]_ ;
  assign \new_[2269]_  = \\L_reg[10] ;
  assign \new_[2270]_  = \\L_reg[20] ;
  assign \new_[2271]_  = \\L_reg[14] ;
  assign \new_[2272]_  = ~\\L_reg[18] ;
  assign \new_[2273]_  = ~\new_[3261]_  | ~\new_[3460]_ ;
  assign \new_[2274]_  = \\FP_R_reg[50] ;
  assign \new_[2275]_  = ~\new_[3189]_  | ~\new_[2848]_ ;
  assign \new_[2276]_  = ~\new_[3186]_  | ~\new_[3336]_ ;
  assign \new_[2277]_  = \new_[3413]_  | \new_[3260]_ ;
  assign \new_[2278]_  = ~\new_[3300]_  | ~\new_[3279]_ ;
  assign \new_[2279]_  = ~\new_[3460]_  | ~\new_[3703]_ ;
  assign \new_[2280]_  = ~\new_[3310]_  | ~\new_[2848]_ ;
  assign \new_[2281]_  = \new_[3267]_  | \new_[3164]_ ;
  assign \new_[2282]_  = ~\new_[2848]_  | ~\new_[3271]_ ;
  assign \new_[2283]_  = ~\new_[3186]_  | ~\new_[3156]_ ;
  assign \new_[2284]_  = \new_[444]_  ? \new_[3489]_  : \new_[3303]_ ;
  assign \new_[2285]_  = ~\new_[2878]_  | ~\new_[2859]_ ;
  assign \new_[2286]_  = ~\new_[2911]_  | ~\new_[2860]_  | ~\new_[2892]_ ;
  assign \new_[2287]_  = ~\new_[2879]_  | ~\new_[2864]_ ;
  assign n1005 = ~\new_[2599]_ ;
  assign n1000 = ~\new_[2596]_ ;
  assign n1020 = ~\new_[2580]_ ;
  assign \new_[2291]_  = ~\new_[2867]_  | ~\new_[2868]_ ;
  assign n1010 = ~\new_[2597]_ ;
  assign n1025 = ~\new_[2442]_ ;
  assign \new_[2294]_  = ~\new_[2881]_  | ~\new_[2876]_ ;
  assign \new_[2295]_  = \\L_reg[2] ;
  assign \new_[2296]_  = ~\new_[2883]_  & (~\new_[3298]_  | ~\new_[4190]_ );
  assign n1035 = ~\new_[2595]_ ;
  assign \new_[2298]_  = ~\new_[2690]_  & (~\new_[3032]_  | ~\new_[4023]_ );
  assign \new_[2299]_  = ~\new_[2655]_  & (~\new_[3021]_  | ~\new_[5068]_ );
  assign \new_[2300]_  = ~\new_[3205]_  & (~\new_[3101]_  | ~\new_[4206]_ );
  assign \new_[2301]_  = ~\new_[4176]_  | ~\new_[2633]_ ;
  assign \new_[2302]_  = ~\new_[2943]_  & (~\new_[2972]_  | ~\new_[4252]_ );
  assign \new_[2303]_  = ~\new_[2695]_  & (~\new_[3018]_  | ~\new_[4186]_ );
  assign \new_[2304]_  = ~\new_[2946]_  & (~\new_[3150]_  | ~\new_[4240]_ );
  assign \new_[2305]_  = ~\new_[2661]_  | ~\new_[2949]_ ;
  assign \new_[2306]_  = ~\new_[2707]_  & (~\new_[3052]_  | ~\new_[4252]_ );
  assign \new_[2307]_  = ~\new_[2708]_  & (~\new_[3246]_  | ~\new_[4232]_ );
  assign \new_[2308]_  = ~\new_[2709]_  | ~\new_[2710]_ ;
  assign \new_[2309]_  = ~\new_[2631]_  | ~\new_[4242]_ ;
  assign \new_[2310]_  = ~\new_[2715]_  & (~\new_[3057]_  | ~\new_[4121]_ );
  assign \new_[2311]_  = ~\new_[2741]_  & (~\new_[3100]_  | ~\new_[4121]_ );
  assign \new_[2312]_  = ~\new_[3195]_  & (~\new_[3051]_  | ~\new_[5068]_ );
  assign \new_[2313]_  = ~\new_[2935]_  & (~\new_[3107]_  | ~\new_[4235]_ );
  assign \new_[2314]_  = ~\new_[2666]_  & (~\new_[3002]_  | ~\new_[4242]_ );
  assign \new_[2315]_  = ~\new_[2678]_  & (~\new_[3039]_  | ~\new_[4233]_ );
  assign \new_[2316]_  = ~\new_[2744]_  & (~\new_[3250]_  | ~\new_[4222]_ );
  assign \new_[2317]_  = ~\new_[2759]_  & (~\new_[2994]_  | ~\new_[4170]_ );
  assign \new_[2318]_  = ~\new_[2689]_  & (~\new_[3019]_  | ~\new_[4198]_ );
  assign \new_[2319]_  = ~\new_[2670]_  & (~\new_[3049]_  | ~\new_[4176]_ );
  assign \new_[2320]_  = ~\new_[2668]_  & (~\new_[3071]_  | ~\new_[5068]_ );
  assign \new_[2321]_  = ~\new_[2724]_  & (~\new_[3125]_  | ~\new_[5068]_ );
  assign \new_[2322]_  = ~\new_[2725]_  & (~\new_[3118]_  | ~\new_[4108]_ );
  assign \new_[2323]_  = ~\new_[2726]_  & (~\new_[3069]_  | ~\new_[4233]_ );
  assign \new_[2324]_  = ~\new_[2727]_  & (~\new_[2995]_  | ~\new_[4109]_ );
  assign \new_[2325]_  = ~\new_[2729]_  & (~\new_[3238]_  | ~\new_[5099]_ );
  assign \new_[2326]_  = ~\new_[2728]_  & (~\new_[3076]_  | ~\new_[4212]_ );
  assign \new_[2327]_  = ~\new_[2731]_  & ~\new_[2957]_ ;
  assign \new_[2328]_  = ~\new_[2730]_  & (~\new_[3243]_  | ~\new_[4239]_ );
  assign \new_[2329]_  = ~\new_[3202]_  & ~\new_[2733]_ ;
  assign \new_[2330]_  = ~\new_[2672]_  & ~\new_[3167]_ ;
  assign \new_[2331]_  = ~\new_[2735]_  & (~\new_[3085]_  | ~\new_[4152]_ );
  assign \new_[2332]_  = ~\new_[3713]_  | ~\desIn[32] ;
  assign \new_[2333]_  = ~\new_[2674]_  & (~\new_[3086]_  | ~\new_[4232]_ );
  assign \new_[2334]_  = ~\new_[3713]_  | ~\desIn[20] ;
  assign \new_[2335]_  = ~\new_[2737]_  & ~\new_[3183]_ ;
  assign \new_[2336]_  = ~\new_[2693]_  & (~\new_[3011]_  | ~\new_[4262]_ );
  assign \new_[2337]_  = ~\new_[2927]_  & (~\new_[3054]_  | ~\new_[4270]_ );
  assign \new_[2338]_  = ~\new_[2869]_  & ~\new_[2745]_ ;
  assign \new_[2339]_  = ~\new_[2677]_  & (~\new_[3113]_  | ~\new_[4793]_ );
  assign \new_[2340]_  = ~\new_[2703]_  & (~\new_[3105]_  | ~\new_[5068]_ );
  assign \new_[2341]_  = ~\new_[2965]_  & (~\new_[3123]_  | ~\new_[4239]_ );
  assign \new_[2342]_  = ~\new_[2747]_  & (~\new_[3028]_  | ~\new_[4102]_ );
  assign \new_[2343]_  = ~\new_[2721]_  & (~\new_[3143]_  | ~\new_[4116]_ );
  assign \new_[2344]_  = ~\new_[2694]_  & (~\new_[3124]_  | ~\new_[4239]_ );
  assign \new_[2345]_  = ~\new_[2749]_  & (~\new_[3383]_  | ~\new_[5097]_ );
  assign \new_[2346]_  = \\FP_R_reg[44] ;
  assign \new_[2347]_  = ~\new_[3208]_  & (~\new_[3043]_  | ~\new_[4170]_ );
  assign \new_[2348]_  = \\L_reg[4] ;
  assign \new_[2349]_  = ~\new_[2755]_  & (~\new_[3129]_  | ~\new_[4206]_ );
  assign \new_[2350]_  = ~\new_[2756]_  & (~\new_[3132]_  | ~\new_[4252]_ );
  assign \new_[2351]_  = ~\new_[2760]_  & (~\new_[3393]_  | ~\new_[4239]_ );
  assign \new_[2352]_  = ~\new_[2684]_  | ~\new_[2981]_ ;
  assign \new_[2353]_  = ~\new_[2685]_  & (~\new_[3139]_  | ~\new_[4237]_ );
  assign \new_[2354]_  = ~\new_[2762]_  & (~\new_[3096]_  | ~\new_[4109]_ );
  assign \new_[2355]_  = ~\new_[3287]_  & (~\new_[3140]_  | ~\new_[4228]_ );
  assign \new_[2356]_  = ~\new_[2763]_  & (~\new_[3365]_  | ~\new_[5097]_ );
  assign \new_[2357]_  = ~\new_[2688]_  & (~\new_[3131]_  | ~\new_[4214]_ );
  assign \new_[2358]_  = ~\new_[2676]_  & (~\new_[3142]_  | ~\new_[4206]_ );
  assign \new_[2359]_  = ~\new_[2739]_  & (~\new_[3491]_  | ~\new_[4216]_ );
  assign \new_[2360]_  = ~\new_[2691]_  & (~\new_[3476]_  | ~\new_[4222]_ );
  assign \new_[2361]_  = ~\new_[2634]_  | ~\new_[2951]_ ;
  assign \new_[2362]_  = ~\new_[2720]_  & (~\new_[3232]_  | ~\new_[4220]_ );
  assign \new_[2363]_  = ~\new_[2664]_  & (~\new_[4176]_  | ~\new_[3109]_ );
  assign \new_[2364]_  = ~\new_[2671]_  & (~\new_[3526]_  | ~\new_[4698]_ );
  assign \new_[2365]_  = ~\new_[2956]_  & (~\new_[3075]_  | ~\new_[4222]_ );
  assign \new_[2366]_  = ~\new_[2738]_  & (~\new_[3080]_  | ~\new_[4220]_ );
  assign \new_[2367]_  = ~\new_[2657]_  & (~\new_[3006]_  | ~\new_[4176]_ );
  assign \new_[2368]_  = ~\new_[2746]_  & (~\new_[3092]_  | ~\new_[4242]_ );
  assign \new_[2369]_  = ~\new_[3197]_  & (~\new_[3075]_  | ~\new_[4176]_ );
  assign \new_[2370]_  = ~\new_[2648]_  | ~\new_[2750]_ ;
  assign \new_[2371]_  = ~\new_[2649]_  | ~\new_[2753]_ ;
  assign \new_[2372]_  = ~\new_[2681]_  & (~\new_[3046]_  | ~\new_[4131]_ );
  assign \new_[2373]_  = ~\new_[2653]_  | ~\new_[2939]_ ;
  assign \new_[2374]_  = ~\new_[2960]_  & (~\new_[2999]_  | ~\new_[4242]_ );
  assign \new_[2375]_  = ~\new_[2765]_  & (~\new_[3334]_  | ~\new_[4113]_ );
  assign \new_[2376]_  = \\FP_R_reg[46] ;
  assign \new_[2377]_  = ~\new_[2912]_  | ~\new_[2640]_ ;
  assign \new_[2378]_  = ~\new_[3017]_  | ~\new_[4196]_ ;
  assign \new_[2379]_  = ~\new_[3130]_  | ~\new_[4208]_ ;
  assign \new_[2380]_  = ~\new_[3048]_  | ~\new_[4222]_ ;
  assign \new_[2381]_  = ~\new_[3012]_  | ~\new_[4242]_ ;
  assign \new_[2382]_  = ~\new_[3117]_  | ~\new_[4196]_ ;
  assign \new_[2383]_  = ~\new_[3116]_  | ~\new_[4113]_ ;
  assign \new_[2384]_  = ~\new_[2999]_  | ~\new_[4220]_ ;
  assign \new_[2385]_  = ~\new_[3048]_  | ~\new_[4069]_ ;
  assign \new_[2386]_  = ~\new_[3116]_  | ~\new_[4021]_ ;
  assign \new_[2387]_  = ~\new_[2952]_  | ~\new_[4196]_ ;
  assign \new_[2388]_  = ~\new_[3137]_  | ~\new_[4113]_ ;
  assign \new_[2389]_  = ~\new_[2915]_  | ~\new_[4222]_ ;
  assign \new_[2390]_  = ~\new_[3135]_  | ~\new_[4698]_ ;
  assign \new_[2391]_  = ~\new_[3017]_  | ~\new_[4208]_ ;
  assign \new_[2392]_  = ~\new_[3037]_  | ~\new_[4222]_ ;
  assign \new_[2393]_  = \new_[3109]_  & \new_[4222]_ ;
  assign \new_[2394]_  = ~\new_[3117]_  | ~\new_[4098]_ ;
  assign \new_[2395]_  = ~\new_[3135]_  | ~\new_[4242]_ ;
  assign \new_[2396]_  = ~\new_[3000]_  | ~\new_[4176]_ ;
  assign \new_[2397]_  = ~\new_[3073]_  | ~\new_[4161]_ ;
  assign \new_[2398]_  = ~\new_[3077]_  | ~\new_[4176]_ ;
  assign \new_[2399]_  = ~\new_[3078]_  | ~\new_[4222]_ ;
  assign \new_[2400]_  = ~\new_[3080]_  | ~\new_[4208]_ ;
  assign \new_[2401]_  = ~\new_[3136]_  | ~\new_[4188]_ ;
  assign \new_[2402]_  = ~\new_[3127]_  | ~\new_[4176]_ ;
  assign \new_[2403]_  = ~\new_[4161]_  | ~\new_[3087]_ ;
  assign \new_[2404]_  = ~\new_[3092]_  | ~\new_[4220]_ ;
  assign \new_[2405]_  = \new_[3087]_  & \new_[4242]_ ;
  assign \new_[2406]_  = ~\new_[3126]_  | ~\new_[4176]_ ;
  assign \new_[2407]_  = ~\new_[3078]_  | ~\new_[4021]_ ;
  assign \new_[2408]_  = ~\new_[3000]_  | ~\new_[4222]_ ;
  assign \new_[2409]_  = ~\new_[3095]_  | ~\new_[4698]_ ;
  assign \new_[2410]_  = ~\new_[3077]_  | ~\new_[4222]_ ;
  assign \new_[2411]_  = ~\new_[3073]_  | ~\new_[4242]_ ;
  assign \new_[2412]_  = \\FP_R_reg[61] ;
  assign \new_[2413]_  = ~\new_[2952]_  | ~\new_[4098]_ ;
  assign \new_[2414]_  = ~\new_[3127]_  | ~\new_[4222]_ ;
  assign \new_[2415]_  = ~\new_[3130]_  | ~\new_[4196]_ ;
  assign \new_[2416]_  = ~\new_[3136]_  | ~\new_[4208]_ ;
  assign \new_[2417]_  = \\FP_R_reg[41] ;
  assign \new_[2418]_  = ~\new_[3046]_  | ~\new_[4222]_ ;
  assign n985 = ~\new_[4570]_ ;
  assign \new_[2420]_  = ~\new_[2915]_  | ~\new_[4069]_ ;
  assign \new_[2421]_  = ~\new_[4143]_  & (~\new_[3503]_  | ~\new_[3292]_ );
  assign \new_[2422]_  = ~\new_[4203]_  & (~\new_[5288]_  | ~\new_[3543]_ );
  assign \new_[2423]_  = ~\new_[3015]_  | ~\new_[4185]_ ;
  assign \new_[2424]_  = ~\new_[5098]_  & (~\new_[5182]_  | ~\new_[3187]_ );
  assign \new_[2425]_  = ~\new_[3161]_  | ~\new_[4241]_ ;
  assign \new_[2426]_  = ~\new_[4269]_  & (~\new_[3533]_  | ~\new_[3599]_ );
  assign \new_[2427]_  = ~\new_[4143]_  & (~\new_[3336]_  | ~\new_[3263]_ );
  assign \new_[2428]_  = ~\new_[3027]_  | ~\new_[4173]_ ;
  assign \new_[2429]_  = ~\new_[3168]_  | ~\new_[5097]_ ;
  assign \new_[2430]_  = ~\new_[3029]_  | ~\new_[4173]_ ;
  assign \new_[2431]_  = ~\new_[4244]_  & (~\new_[3280]_  | ~\new_[3537]_ );
  assign \new_[2432]_  = ~\new_[3041]_  | ~\new_[4198]_ ;
  assign \new_[2433]_  = ~\new_[3093]_  | ~\new_[4216]_ ;
  assign \new_[2434]_  = ~\new_[3050]_  | ~\new_[4233]_ ;
  assign \new_[2435]_  = ~\new_[4178]_  & (~\new_[3261]_  | ~\new_[3524]_ );
  assign \new_[2436]_  = ~\new_[3001]_  | ~\new_[4174]_ ;
  assign \new_[2437]_  = ~\new_[2667]_ ;
  assign \new_[2438]_  = ~\new_[3091]_  | ~\new_[4208]_ ;
  assign \new_[2439]_  = ~\new_[3060]_  | ~\new_[4199]_ ;
  assign \new_[2440]_  = ~\new_[3059]_  | ~\new_[4174]_ ;
  assign \new_[2441]_  = ~\new_[5098]_  & (~\new_[5289]_  | ~\new_[3421]_ );
  assign \new_[2442]_  = (~\new_[3291]_  | ~\new_[3739]_ ) & (~\new_[3759]_  | ~\desIn[21] );
  assign \new_[2443]_  = ~\new_[2886]_  | ~\new_[5097]_ ;
  assign \new_[2444]_  = ~\new_[4269]_  & (~\new_[4393]_  | ~\new_[3299]_ );
  assign \new_[2445]_  = ~\new_[3079]_  | ~\new_[4185]_ ;
  assign \new_[2446]_  = ~\new_[4163]_  & (~\new_[3517]_  | ~\new_[3189]_ );
  assign \new_[2447]_  = ~\new_[4269]_  & (~\new_[3186]_  | ~\new_[3402]_ );
  assign \new_[2448]_  = ~\new_[4143]_  & (~\new_[3281]_  | ~\new_[3305]_ );
  assign \new_[2449]_  = ~\new_[3097]_  | ~\new_[4250]_ ;
  assign \new_[2450]_  = ~\new_[4203]_  & (~\new_[3265]_  | ~\new_[3646]_ );
  assign \new_[2451]_  = ~\new_[2998]_  | ~\new_[4173]_ ;
  assign \new_[2452]_  = ~\new_[2934]_  | ~\new_[5097]_ ;
  assign \new_[2453]_  = ~\new_[4143]_  & (~\new_[3468]_  | ~\new_[3278]_ );
  assign \new_[2454]_  = ~\new_[3010]_  | ~\new_[4158]_ ;
  assign \new_[2455]_  = ~\new_[4244]_  & (~\new_[3276]_  | ~\new_[4790]_ );
  assign \new_[2456]_  = ~\new_[4192]_  & (~\new_[3270]_  | ~\new_[3550]_ );
  assign \new_[2457]_  = ~\new_[4143]_  & (~\new_[3257]_  | ~\new_[3276]_ );
  assign \new_[2458]_  = ~\new_[3084]_  | ~\new_[4174]_ ;
  assign \new_[2459]_  = ~\new_[3128]_  | ~\new_[4199]_ ;
  assign \new_[2460]_  = ~\new_[4143]_  & (~\new_[3271]_  | ~\new_[4387]_ );
  assign \new_[2461]_  = ~\new_[3106]_  | ~\new_[5097]_ ;
  assign \new_[2462]_  = ~\new_[3065]_  | ~\new_[4241]_ ;
  assign \new_[2463]_  = ~\new_[2926]_  | ~\new_[5175]_ ;
  assign \new_[2464]_  = ~\new_[4189]_  & (~\new_[3332]_  | ~\new_[3254]_ );
  assign \new_[2465]_  = ~\new_[3044]_  | ~\new_[4109]_ ;
  assign \new_[2466]_  = ~\new_[3112]_  | ~\new_[4102]_ ;
  assign \new_[2467]_  = ~\new_[4184]_  & (~\new_[3300]_  | ~\new_[3299]_ );
  assign \new_[2468]_  = ~\new_[3034]_  | ~\new_[4276]_ ;
  assign \new_[2469]_  = ~\new_[3024]_  | ~\new_[4108]_ ;
  assign \new_[2470]_  = ~\new_[3023]_  | ~\new_[4228]_ ;
  assign \new_[2471]_  = ~\new_[3104]_  | ~\new_[5068]_ ;
  assign \new_[2472]_  = ~\new_[3089]_  | ~\new_[4116]_ ;
  assign \new_[2473]_  = ~\new_[4253]_  & (~\new_[3269]_  | ~\new_[3705]_ );
  assign \new_[2474]_  = ~\new_[3058]_  | ~\new_[3985]_ ;
  assign \new_[2475]_  = ~\new_[3003]_  | ~\new_[4214]_ ;
  assign \new_[2476]_  = ~\new_[4104]_  & (~\new_[5289]_  | ~\new_[3405]_ );
  assign \new_[2477]_  = ~\new_[4189]_  & (~\new_[3261]_  | ~\new_[3485]_ );
  assign \new_[2478]_  = ~\new_[3025]_  | ~\new_[4228]_ ;
  assign \new_[2479]_  = ~\new_[3026]_  | ~\new_[5068]_ ;
  assign \new_[2480]_  = ~\new_[3030]_  | ~\new_[4206]_ ;
  assign \new_[2481]_  = ~\new_[3115]_  | ~\new_[4160]_ ;
  assign \new_[2482]_  = ~\new_[3040]_  | ~\new_[4226]_ ;
  assign \new_[2483]_  = ~\new_[3045]_  | ~\new_[4270]_ ;
  assign \new_[2484]_  = ~\new_[3103]_  | ~\new_[4252]_ ;
  assign \new_[2485]_  = ~\new_[3056]_  | ~\new_[4133]_ ;
  assign \new_[2486]_  = ~\new_[3042]_  | ~\new_[4226]_ ;
  assign \new_[2487]_  = ~\new_[4271]_  & (~\new_[3265]_  | ~\new_[3456]_ );
  assign \new_[2488]_  = ~\new_[3108]_  | ~\new_[4133]_ ;
  assign n990 = ~\new_[3589]_  | (~\new_[3295]_  & ~\new_[3759]_ );
  assign \new_[2490]_  = ~\new_[3090]_  | ~\new_[5068]_ ;
  assign \new_[2491]_  = ~\new_[4255]_  & (~\new_[3266]_  | ~\new_[3485]_ );
  assign \new_[2492]_  = ~\new_[3061]_  | ~\new_[4245]_ ;
  assign \new_[2493]_  = ~\new_[4792]_  & (~\new_[3269]_  | ~\new_[4382]_ );
  assign \new_[2494]_  = ~\new_[3063]_  | ~\new_[4240]_ ;
  assign \new_[2495]_  = ~\new_[3005]_  | ~\new_[4232]_ ;
  assign \new_[2496]_  = ~\new_[3062]_  | ~\new_[5068]_ ;
  assign \new_[2497]_  = ~\new_[3144]_  | ~\new_[4256]_ ;
  assign \new_[2498]_  = ~\new_[4104]_  & (~\new_[5181]_  | ~\new_[3263]_ );
  assign \new_[2499]_  = ~\new_[3066]_  | ~\new_[4160]_ ;
  assign \new_[2500]_  = ~\new_[3067]_  | ~\new_[4121]_ ;
  assign \new_[2501]_  = ~\new_[4189]_  & (~\new_[3336]_  | ~\new_[3271]_ );
  assign \new_[2502]_  = ~\new_[3072]_  | ~\new_[4793]_ ;
  assign \new_[2503]_  = ~\new_[3074]_  | ~\new_[4226]_ ;
  assign \new_[2504]_  = ~\new_[3064]_  | ~\new_[4126]_ ;
  assign \new_[2505]_  = ~\new_[3020]_  | ~\new_[4240]_ ;
  assign \new_[2506]_  = ~\new_[4085]_  & (~\new_[3418]_  | ~\new_[3517]_ );
  assign \new_[2507]_  = ~\new_[3081]_  | ~\new_[4186]_ ;
  assign \new_[2508]_  = ~\new_[4181]_  & (~\new_[3592]_  | ~\new_[3558]_ );
  assign \new_[2509]_  = ~\new_[3083]_  | ~\new_[4239]_ ;
  assign \new_[2510]_  = ~\new_[4264]_  & (~\new_[5182]_  | ~\new_[4383]_ );
  assign \new_[2511]_  = ~\new_[4164]_  & (~\new_[5183]_  | ~\new_[3336]_ );
  assign \new_[2512]_  = ~\new_[4197]_  & (~\new_[3405]_  | ~\new_[3276]_ );
  assign \new_[2513]_  = ~\new_[4189]_  & (~\new_[3299]_  | ~\new_[4784]_ );
  assign \new_[2514]_  = ~\new_[4271]_  & (~\new_[3531]_  | ~\new_[4384]_ );
  assign \new_[2515]_  = ~\new_[3958]_  & (~\new_[3450]_  | ~\new_[3262]_ );
  assign \new_[2516]_  = ~\new_[4168]_  & (~\new_[3419]_  | ~\new_[3531]_ );
  assign \new_[2517]_  = ~\new_[3008]_  | ~\new_[5068]_ ;
  assign \new_[2518]_  = ~\new_[3014]_  | ~\new_[4140]_ ;
  assign \new_[2519]_  = ~\new_[3110]_  | ~\new_[4152]_ ;
  assign \new_[2520]_  = ~\new_[4169]_  & (~\new_[3293]_  | ~\new_[3263]_ );
  assign \new_[2521]_  = ~\new_[4179]_  & (~\new_[3189]_  | ~\new_[3336]_ );
  assign \new_[2522]_  = \new_[3171]_  & \new_[4214]_ ;
  assign \new_[2523]_  = ~\new_[2963]_  | ~\new_[4200]_ ;
  assign \new_[2524]_  = ~\new_[3114]_  | ~\new_[4245]_ ;
  assign \new_[2525]_  = ~\new_[3038]_  | ~\new_[4113]_ ;
  assign \new_[2526]_  = ~\new_[3119]_  | ~\new_[4256]_ ;
  assign \new_[2527]_  = ~\new_[3121]_  | ~\new_[4152]_ ;
  assign \new_[2528]_  = ~\new_[3070]_  | ~\new_[4047]_ ;
  assign \new_[2529]_  = ~\new_[4268]_  & (~\new_[3186]_  | ~\new_[4401]_ );
  assign \new_[2530]_  = ~\new_[4189]_  & (~\new_[3460]_  | ~\new_[3400]_ );
  assign \new_[2531]_  = ~\new_[2930]_  | ~\new_[4121]_ ;
  assign \new_[2532]_  = ~\new_[3141]_  | ~\new_[4133]_ ;
  assign \new_[2533]_  = ~\new_[4264]_  & (~\new_[3299]_  | ~\new_[3545]_ );
  assign \new_[2534]_  = ~\new_[4164]_  & (~\new_[3279]_  | ~\new_[5263]_ );
  assign \new_[2535]_  = ~\new_[4085]_  & (~\new_[3276]_  | ~\new_[3299]_ );
  assign \new_[2536]_  = ~\new_[3013]_  | ~\new_[4133]_ ;
  assign \new_[2537]_  = ~\new_[3031]_  | ~\new_[4209]_ ;
  assign \new_[2538]_  = ~\new_[2996]_  | ~\new_[4152]_ ;
  assign \new_[2539]_  = ~\new_[5063]_  & (~\new_[3199]_  | ~\new_[3550]_ );
  assign \new_[2540]_  = ~\new_[4184]_  & (~\new_[3533]_  | ~\new_[3255]_ );
  assign \new_[2541]_  = ~\new_[3055]_  | ~\new_[4204]_ ;
  assign \new_[2542]_  = ~\new_[3007]_  | ~\new_[4140]_ ;
  assign \new_[2543]_  = ~\new_[3102]_  | ~\new_[4170]_ ;
  assign \new_[2544]_  = ~\new_[4184]_  & (~\new_[3254]_  | ~\new_[3468]_ );
  assign \new_[2545]_  = ~\new_[5063]_  & (~\new_[3268]_  | ~\new_[3278]_ );
  assign \new_[2546]_  = \\L_reg[29] ;
  assign \new_[2547]_  = \\L_reg[9] ;
  assign \new_[2548]_  = ~\new_[4405]_  | ~\new_[3488]_ ;
  assign \new_[2549]_  = ~\new_[3454]_  | ~\new_[3468]_ ;
  assign \new_[2550]_  = ~\new_[3153]_  | ~\new_[3703]_ ;
  assign \new_[2551]_  = ~\new_[3157]_  | ~\new_[3703]_ ;
  assign \new_[2552]_  = ~\new_[4382]_  | ~\new_[3443]_ ;
  assign \new_[2553]_  = ~\new_[3300]_  | ~\new_[5241]_ ;
  assign \new_[2554]_  = ~\new_[3501]_  | ~\new_[3488]_ ;
  assign \new_[2555]_  = ~\new_[4385]_  | ~\new_[3405]_ ;
  assign \new_[2556]_  = ~\new_[3454]_  | ~\new_[3645]_ ;
  assign \new_[2557]_  = ~\new_[3266]_  | ~\new_[3314]_ ;
  assign \new_[2558]_  = ~\new_[3154]_  | ~\new_[3564]_ ;
  assign \new_[2559]_  = ~\new_[3488]_  | ~\new_[3271]_ ;
  assign \new_[2560]_  = ~\new_[3414]_  | ~\new_[3433]_ ;
  assign \new_[2561]_  = ~\new_[2961]_  | ~\new_[3407]_ ;
  assign \new_[2562]_  = ~\new_[3254]_  | ~\new_[3433]_ ;
  assign \new_[2563]_  = ~\new_[3409]_  | ~\new_[3306]_ ;
  assign \new_[2564]_  = ~\new_[3170]_  | ~\new_[3421]_ ;
  assign \new_[2565]_  = \new_[4791]_  | \new_[3477]_ ;
  assign \new_[2566]_  = ~\new_[3174]_  | ~\new_[3404]_ ;
  assign \new_[2567]_  = \new_[3166]_  | \new_[3509]_ ;
  assign \new_[2568]_  = ~\new_[3406]_  | ~\new_[4385]_ ;
  assign \new_[2569]_  = ~\new_[2961]_  | ~\new_[3757]_ ;
  assign \new_[2570]_  = ~\new_[3261]_  | ~\new_[2902]_ ;
  assign \new_[2571]_  = ~\new_[4382]_  | ~\new_[3488]_ ;
  assign \new_[2572]_  = ~\new_[2978]_  | ~\new_[4387]_ ;
  assign \new_[2573]_  = \new_[3158]_  | \new_[3677]_ ;
  assign \new_[2574]_  = ~\new_[3170]_  | ~\new_[3257]_ ;
  assign \new_[2575]_  = ~\new_[3435]_  | ~\new_[3155]_ ;
  assign \new_[2576]_  = ~\new_[3299]_  | ~\new_[3426]_ ;
  assign \new_[2577]_  = ~\new_[3269]_  | ~\new_[2978]_ ;
  assign \new_[2578]_  = ~\new_[3587]_  | ~\new_[3157]_ ;
  assign \new_[2579]_  = \new_[3548]_  | \new_[3148]_ ;
  assign \new_[2580]_  = (~\new_[3294]_  | ~\new_[3739]_ ) & (~\new_[3759]_  | ~\desIn[17] );
  assign \new_[2581]_  = ~\new_[3174]_  | ~\new_[3414]_ ;
  assign \new_[2582]_  = ~\new_[3407]_  | ~\new_[3414]_ ;
  assign \new_[2583]_  = ~\new_[3266]_  | ~\new_[5273]_ ;
  assign \new_[2584]_  = ~\new_[3425]_  | ~\new_[3414]_ ;
  assign \new_[2585]_  = ~\new_[5181]_  | ~\new_[2978]_ ;
  assign \new_[2586]_  = ~\new_[3314]_  | ~\new_[3255]_ ;
  assign \new_[2587]_  = ~\new_[4385]_  | ~\new_[5240]_ ;
  assign \new_[2588]_  = ~\new_[2902]_  | ~\new_[3400]_ ;
  assign \new_[2589]_  = ~\new_[4168]_  & (~\new_[3405]_  | ~\new_[3262]_ );
  assign \new_[2590]_  = ~\new_[4385]_  | ~\new_[3257]_ ;
  assign \new_[2591]_  = \new_[3146]_  | \new_[3598]_ ;
  assign \new_[2592]_  = ~\new_[3261]_  | ~\new_[3153]_ ;
  assign \new_[2593]_  = ~\new_[3535]_  | ~\new_[3404]_ ;
  assign n1105 = \new_[4713]_ ;
  assign \new_[2595]_  = ~\new_[3159]_  & (~\new_[3713]_  | ~\desIn[49] );
  assign \new_[2596]_  = (~\new_[3272]_  | ~\new_[3809]_ ) & (~\new_[3759]_  | ~\desIn[51] );
  assign \new_[2597]_  = (~\new_[3274]_  | ~\new_[3739]_ ) & (~\new_[3837]_  | ~\desIn[53] );
  assign n1125 = ~\new_[2700]_ ;
  assign \new_[2599]_  = (~\new_[3289]_  | ~\new_[3809]_ ) & (~\new_[3914]_  | ~\desIn[41] );
  assign \new_[2600]_  = ~\new_[3214]_  & (~\new_[3180]_  | ~\new_[4118]_ );
  assign \new_[2601]_  = ~n995;
  assign \new_[2602]_  = ~n995;
  assign n1110 = ~\new_[2854]_ ;
  assign n1155 = ~\new_[4882]_ ;
  assign \new_[2605]_  = ~\new_[3184]_  & (~\new_[3297]_  | ~\new_[4262]_ );
  assign \new_[2606]_  = ~\new_[2989]_  & (~\new_[3381]_  | ~\new_[4262]_ );
  assign \new_[2607]_  = ~\new_[2945]_  & (~\new_[3222]_  | ~\new_[4118]_ );
  assign \new_[2608]_  = ~\new_[2925]_  | ~\new_[2950]_ ;
  assign \new_[2609]_  = ~\new_[2938]_  & (~\new_[3586]_  | ~\new_[4215]_ );
  assign \new_[2610]_  = ~\new_[3273]_  | ~\new_[3443]_ ;
  assign \new_[2611]_  = ~\new_[2967]_  & (~\new_[3223]_  | ~\new_[4176]_ );
  assign \new_[2612]_  = ~\new_[2976]_  | ~\new_[2964]_ ;
  assign \new_[2613]_  = ~\new_[2968]_  | ~\new_[2969]_ ;
  assign \new_[2614]_  = ~\new_[2970]_  | ~\new_[3160]_ ;
  assign \new_[2615]_  = ~\new_[3193]_  & (~\new_[3285]_  | ~\new_[4121]_ );
  assign \new_[2616]_  = ~\new_[3211]_  & (~\new_[3251]_  | ~\new_[4222]_ );
  assign \new_[2617]_  = ~\new_[2985]_  | ~\new_[2940]_ ;
  assign \new_[2618]_  = ~\new_[2987]_  | ~\new_[2988]_ ;
  assign \new_[2619]_  = ~\new_[2990]_  | ~\new_[2991]_ ;
  assign \new_[2620]_  = ~\new_[2942]_  | ~\new_[2941]_ ;
  assign \new_[2621]_  = ~\new_[2979]_  & (~\new_[3348]_  | ~\new_[4161]_ );
  assign \new_[2622]_  = ~\new_[3533]_  | ~\new_[3458]_ ;
  assign \new_[2623]_  = ~\new_[3317]_  & (~\new_[3233]_  | ~\new_[4176]_ );
  assign \new_[2624]_  = ~\new_[2921]_  | ~\new_[2980]_ ;
  assign \new_[2625]_  = ~\new_[2924]_  | ~\new_[2986]_ ;
  assign \new_[2626]_  = ~\new_[4180]_  & (~\new_[3587]_  | ~\new_[3216]_ );
  assign \new_[2627]_  = ~\new_[4272]_  & (~\new_[3700]_  | ~\new_[3217]_ );
  assign \new_[2628]_  = ~\new_[4268]_  & (~\new_[3664]_  | ~\new_[3221]_ );
  assign \new_[2629]_  = (~\new_[3347]_  | ~\new_[4069]_ ) & (~\new_[3219]_  | ~\new_[4098]_ );
  assign \new_[2630]_  = ~\new_[4162]_  & (~\new_[3409]_  | ~\new_[3221]_ );
  assign \new_[2631]_  = ~\new_[3221]_  | ~\new_[3676]_ ;
  assign \new_[2632]_  = ~\new_[3229]_  | ~\new_[4220]_ ;
  assign \new_[2633]_  = ~\new_[3675]_  | ~\new_[3221]_ ;
  assign \new_[2634]_  = ~\new_[3237]_  | ~\new_[4176]_ ;
  assign \new_[2635]_  = ~\new_[3248]_  | ~\new_[4161]_ ;
  assign \new_[2636]_  = ~\new_[3232]_  | ~\new_[4242]_ ;
  assign \new_[2637]_  = ~\new_[3234]_  | ~\new_[4698]_ ;
  assign \new_[2638]_  = ~\new_[3224]_  | ~\new_[4242]_ ;
  assign \new_[2639]_  = ~\new_[2898]_ ;
  assign \new_[2640]_  = ~\new_[3177]_  | ~\new_[4242]_ ;
  assign \new_[2641]_  = ~\new_[3224]_  | ~\new_[4698]_ ;
  assign \new_[2642]_  = ~\new_[3230]_  | ~\new_[4208]_ ;
  assign \new_[2643]_  = ~\new_[3242]_  | ~\new_[4222]_ ;
  assign \new_[2644]_  = ~\new_[4197]_  & (~\new_[4784]_  | ~\new_[3421]_ );
  assign \new_[2645]_  = ~\new_[3283]_  | ~\new_[4242]_ ;
  assign \new_[2646]_  = ~\new_[3229]_  | ~\new_[4242]_ ;
  assign \new_[2647]_  = ~\new_[3242]_  | ~\new_[4131]_ ;
  assign \new_[2648]_  = ~\new_[3230]_  | ~\new_[4188]_ ;
  assign \new_[2649]_  = ~\new_[3177]_  | ~\new_[4196]_ ;
  assign \new_[2650]_  = ~\new_[3283]_  | ~\new_[4220]_ ;
  assign \new_[2651]_  = ~\new_[3694]_  | ~\new_[3221]_ ;
  assign \new_[2652]_  = ~\new_[3655]_  | ~\new_[3221]_ ;
  assign \new_[2653]_  = ~\new_[3219]_  | ~\new_[4188]_ ;
  assign \new_[2654]_  = ~\new_[3237]_  | ~\new_[4222]_ ;
  assign \new_[2655]_  = ~\new_[5174]_  & (~\new_[3412]_  | ~\new_[3535]_ );
  assign \new_[2656]_  = ~\new_[4203]_  & (~\new_[3387]_  | ~\new_[3645]_ );
  assign \new_[2657]_  = ~\new_[4143]_  & (~\new_[3558]_  | ~\new_[3419]_ );
  assign \new_[2658]_  = ~\new_[4143]_  & (~\new_[3418]_  | ~\new_[4403]_ );
  assign \new_[2659]_  = ~\new_[3236]_  | ~\new_[4212]_ ;
  assign \new_[2660]_  = ~\new_[4269]_  & (~\new_[3408]_  | ~\new_[3528]_ );
  assign \new_[2661]_  = ~\new_[3226]_  | ~\new_[5175]_ ;
  assign \new_[2662]_  = ~\new_[3253]_  | ~\new_[4242]_ ;
  assign \new_[2663]_  = ~\new_[4192]_  & (~\new_[3534]_  | ~\new_[3313]_ );
  assign \new_[2664]_  = ~\new_[5098]_  & (~\new_[3479]_  | ~\new_[3533]_ );
  assign \new_[2665]_  = ~\new_[3220]_  | ~\new_[5097]_ ;
  assign \new_[2666]_  = ~\new_[5098]_  & (~\new_[4657]_  | ~\new_[3707]_ );
  assign \new_[2667]_  = ~\new_[4143]_  & (~\new_[3332]_  | ~\new_[3387]_ );
  assign \new_[2668]_  = ~\new_[4238]_  & (~\new_[3409]_  | ~\new_[3663]_ );
  assign \new_[2669]_  = ~n1135;
  assign \new_[2670]_  = ~\new_[4178]_  & (~\new_[3315]_  | ~\new_[3408]_ );
  assign \new_[2671]_  = ~\new_[4211]_  & (~\new_[3501]_  | ~\new_[3635]_ );
  assign \new_[2672]_  = ~\new_[4203]_  & (~\new_[3544]_  | ~\new_[3433]_ );
  assign \new_[2673]_  = ~\new_[4238]_  & (~\new_[3450]_  | ~\new_[3426]_ );
  assign \new_[2674]_  = ~\new_[4244]_  & (~\new_[3472]_  | ~\new_[3309]_ );
  assign \new_[2675]_  = ~\new_[3258]_  | ~\new_[4250]_ ;
  assign \new_[2676]_  = ~\new_[5098]_  & (~\new_[3482]_  | ~\new_[3581]_ );
  assign \new_[2677]_  = ~\new_[5098]_  & (~\new_[3402]_  | ~\new_[3319]_ );
  assign \new_[2678]_  = ~\new_[4163]_  & (~\new_[3588]_  | ~\new_[3313]_ );
  assign \new_[2679]_  = ~\new_[3239]_  | ~\new_[4212]_ ;
  assign \new_[2680]_  = ~\new_[4244]_  & (~\new_[3621]_  | ~\new_[3484]_ );
  assign \new_[2681]_  = ~\new_[5098]_  & (~\new_[3414]_  | ~\new_[3753]_ );
  assign \new_[2682]_  = ~\new_[4192]_  & (~\new_[3517]_  | ~\new_[4405]_ );
  assign \new_[2683]_  = ~\new_[3418]_  | ~\new_[3492]_ ;
  assign \new_[2684]_  = ~\new_[3252]_  | ~\new_[4185]_ ;
  assign \new_[2685]_  = ~\new_[4269]_  & (~\new_[3458]_  | ~\new_[3432]_ );
  assign \new_[2686]_  = ~\new_[4211]_  & (~\new_[3420]_  | ~\new_[3614]_ );
  assign \new_[2687]_  = ~\new_[3244]_  | ~\new_[4174]_ ;
  assign \new_[2688]_  = ~\new_[5174]_  & (~\new_[3332]_  | ~\new_[3408]_ );
  assign \new_[2689]_  = ~\new_[4269]_  & (~\new_[3443]_  | ~\new_[3319]_ );
  assign \new_[2690]_  = ~\new_[4168]_  & (~\new_[3534]_  | ~\new_[3400]_ );
  assign \new_[2691]_  = ~\new_[4272]_  & (~\new_[3725]_  | ~\new_[3640]_ );
  assign \new_[2692]_  = ~n1225;
  assign \new_[2693]_  = ~\new_[4167]_  & (~\new_[3655]_  | ~\new_[3760]_ );
  assign \new_[2694]_  = ~\new_[4268]_  & (~\new_[5288]_  | ~\new_[5240]_ );
  assign \new_[2695]_  = ~\new_[4181]_  & (~\new_[3636]_  | ~\new_[3426]_ );
  assign \new_[2696]_  = ~\new_[3218]_  | ~\new_[4190]_ ;
  assign \new_[2697]_  = ~\new_[4792]_  & (~\new_[4393]_  | ~\new_[3531]_ );
  assign \new_[2698]_  = ~\new_[4792]_  & (~\new_[3341]_  | ~\new_[3662]_ );
  assign \new_[2699]_  = ~\new_[4135]_  & (~\new_[3503]_  | ~\new_[3676]_ );
  assign \new_[2700]_  = (~\new_[3462]_  | ~\new_[3809]_ ) & (~\new_[3914]_  | ~\desIn[47] );
  assign \new_[2701]_  = ~\new_[3247]_  | ~\new_[4215]_ ;
  assign \new_[2702]_  = ~\new_[4180]_  & (~\new_[3418]_  | ~\new_[3717]_ );
  assign \new_[2703]_  = ~\new_[4253]_  & (~\new_[3649]_  | ~\new_[4386]_ );
  assign \new_[2704]_  = ~\new_[4264]_  & (~\new_[4379]_  | ~\new_[3426]_ );
  assign \new_[2705]_  = ~\new_[3444]_  | ~\new_[3599]_ ;
  assign \new_[2706]_  = ~\new_[4181]_  & (~\new_[3649]_  | ~\new_[3402]_ );
  assign \new_[2707]_  = ~\new_[4104]_  & (~\new_[3503]_  | ~\new_[3414]_ );
  assign \new_[2708]_  = ~\new_[4164]_  & (~\new_[3482]_  | ~\new_[3457]_ );
  assign \new_[2709]_  = ~\new_[3228]_  | ~\new_[4118]_ ;
  assign \new_[2710]_  = ~\new_[3235]_  | ~\new_[4239]_ ;
  assign \new_[2711]_  = ~\new_[4259]_  & (~\new_[3454]_  | ~\new_[3407]_ );
  assign \new_[2712]_  = ~\new_[3225]_  | ~\new_[4108]_ ;
  assign \new_[2713]_  = ~\new_[3215]_  | ~\new_[4190]_ ;
  assign \new_[2714]_  = ~\new_[4189]_  & (~\new_[3588]_  | ~\new_[3401]_ );
  assign \new_[2715]_  = ~\new_[4271]_  & (~\new_[3305]_  | ~\new_[3309]_ );
  assign \new_[2716]_  = ~\new_[3206]_  | ~\new_[4108]_ ;
  assign \new_[2717]_  = ~\new_[3249]_  | ~\new_[4126]_ ;
  assign \new_[2718]_  = ~\new_[4169]_  & (~\new_[3315]_  | ~\new_[3457]_ );
  assign \new_[2719]_  = ~\new_[3564]_  | ~\new_[3270]_ ;
  assign \new_[2720]_  = ~\new_[4255]_  & (~\new_[3454]_  | ~\new_[3482]_ );
  assign \new_[2721]_  = ~\new_[4164]_  & (~\new_[3313]_  | ~\new_[3446]_ );
  assign \new_[2722]_  = ~\new_[4189]_  & (~\new_[3419]_  | ~\new_[4380]_ );
  assign \new_[2723]_  = ~\new_[3444]_  | ~\new_[3270]_ ;
  assign \new_[2724]_  = ~\new_[4169]_  & (~\new_[3631]_  | ~\new_[5240]_ );
  assign \new_[2725]_  = ~\new_[4264]_  & (~\new_[3488]_  | ~\new_[3319]_ );
  assign \new_[2726]_  = ~\new_[4255]_  & (~\new_[3537]_  | ~\new_[3426]_ );
  assign \new_[2727]_  = ~\new_[4164]_  & (~\new_[3443]_  | ~\new_[3472]_ );
  assign \new_[2728]_  = ~\new_[4272]_  & (~\new_[3492]_  | ~\new_[3429]_ );
  assign \new_[2729]_  = ~\new_[4792]_  & (~\new_[3492]_  | ~\new_[3484]_ );
  assign \new_[2730]_  = ~\new_[4189]_  & (~\new_[3341]_  | ~\new_[3629]_ );
  assign \new_[2731]_  = ~\new_[4189]_  & (~\new_[3725]_  | ~\new_[4657]_ );
  assign \new_[2732]_  = ~n1140;
  assign \new_[2733]_  = ~\new_[4792]_  & (~\new_[3490]_  | ~\new_[3725]_ );
  assign \new_[2734]_  = ~\new_[3245]_  | ~\new_[4215]_ ;
  assign \new_[2735]_  = ~\new_[4164]_  & (~\new_[3419]_  | ~\new_[3537]_ );
  assign \new_[2736]_  = ~\new_[4168]_  & (~\new_[3435]_  | ~\new_[5263]_ );
  assign \new_[2737]_  = ~\new_[4268]_  & (~\new_[3480]_  | ~\new_[3624]_ );
  assign \new_[2738]_  = ~\new_[4115]_  & (~\new_[5181]_  | ~\new_[4405]_ );
  assign \new_[2739]_  = ~\new_[4264]_  & (~\new_[3423]_  | ~\new_[3420]_ );
  assign \new_[2740]_  = ~\new_[3958]_  & (~\new_[3588]_  | ~\new_[3703]_ );
  assign \new_[2741]_  = ~\new_[4189]_  & (~\new_[3423]_  | ~\new_[5278]_ );
  assign \new_[2742]_  = ~\new_[4135]_  & (~\new_[5269]_  | ~\new_[3387]_ );
  assign \new_[2743]_  = ~\new_[3240]_  | ~\new_[4121]_ ;
  assign \new_[2744]_  = ~\new_[4189]_  & (~\new_[3471]_  | ~\new_[3426]_ );
  assign \new_[2745]_  = ~\new_[4169]_  & (~\new_[3405]_  | ~\new_[4785]_ );
  assign \new_[2746]_  = ~\new_[4139]_  & (~\new_[5240]_  | ~\new_[3640]_ );
  assign \new_[2747]_  = ~\new_[5063]_  & (~\new_[3336]_  | ~\new_[4405]_ );
  assign \new_[2748]_  = ~\new_[4179]_  & (~\new_[3534]_  | ~\new_[3442]_ );
  assign \new_[2749]_  = ~\new_[4792]_  & (~\new_[3501]_  | ~\new_[3312]_ );
  assign \new_[2750]_  = ~\new_[3231]_  | ~\new_[4228]_ ;
  assign \new_[2751]_  = ~\new_[4181]_  & (~\new_[3438]_  | ~\new_[3443]_ );
  assign \new_[2752]_  = ~\new_[4169]_  & (~\new_[5280]_  | ~\new_[3333]_ );
  assign \new_[2753]_  = ~\new_[3241]_  | ~\new_[4232]_ ;
  assign \new_[2754]_  = ~\new_[4164]_  & (~\new_[3329]_  | ~\new_[3564]_ );
  assign \new_[2755]_  = ~\new_[4180]_  & (~\new_[3478]_  | ~\new_[5279]_ );
  assign \new_[2756]_  = ~\new_[4189]_  & (~\new_[3758]_  | ~\new_[3433]_ );
  assign \new_[2757]_  = ~\new_[4247]_  & (~\new_[3645]_  | ~\new_[3417]_ );
  assign \new_[2758]_  = ~\new_[4247]_  & (~\new_[3422]_  | ~\new_[3533]_ );
  assign \new_[2759]_  = ~\new_[4792]_  & (~\new_[3676]_  | ~\new_[3608]_ );
  assign \new_[2760]_  = ~\new_[4259]_  & (~\new_[3420]_  | ~\new_[3625]_ );
  assign \new_[2761]_  = ~\new_[3181]_  | ~\new_[4176]_ ;
  assign \new_[2762]_  = ~\new_[5063]_  & (~\new_[3446]_  | ~\new_[3401]_ );
  assign \new_[2763]_  = ~\new_[4792]_  & (~\new_[3333]_  | ~\new_[3760]_ );
  assign \new_[2764]_  = ~\new_[4264]_  & (~\new_[3638]_  | ~\new_[3480]_ );
  assign \new_[2765]_  = ~\new_[4168]_  & (~\new_[3422]_  | ~\new_[3460]_ );
  assign \new_[2766]_  = ~\new_[4115]_  & (~\new_[3534]_  | ~\new_[3327]_ );
  assign \new_[2767]_  = ~\new_[4080]_  & (~\new_[3446]_  | ~\new_[3329]_ );
  assign \new_[2768]_  = ~\new_[4189]_  & (~\new_[3454]_  | ~\new_[3560]_ );
  assign \new_[2769]_  = ~\new_[3576]_  | ~\new_[3465]_ ;
  assign \new_[2770]_  = ~\new_[3402]_  | ~\new_[3415]_ ;
  assign \new_[2771]_  = ~\new_[3533]_  | ~\new_[3199]_ ;
  assign \new_[2772]_  = ~\new_[3344]_ ;
  assign \new_[2773]_  = ~\new_[3528]_  | ~\new_[3646]_ ;
  assign \new_[2774]_  = ~\new_[3498]_  | ~\new_[3268]_ ;
  assign \new_[2775]_  = ~\new_[3444]_  | ~\new_[3266]_ ;
  assign \new_[2776]_  = ~\new_[3264]_  | ~\new_[3273]_ ;
  assign \new_[2777]_  = ~\new_[3533]_  | ~\new_[3442]_ ;
  assign \new_[2778]_  = ~\new_[3576]_  | ~\new_[3406]_ ;
  assign \new_[2779]_  = ~\new_[3004]_ ;
  assign \new_[2780]_  = ~\new_[3275]_  | ~\new_[3450]_ ;
  assign \new_[2781]_  = ~\new_[5263]_  | ~\new_[3299]_ ;
  assign \new_[2782]_  = \new_[3307]_  | \new_[3302]_ ;
  assign \new_[2783]_  = ~\new_[3418]_  | ~\new_[3643]_ ;
  assign \new_[2784]_  = ~\new_[3261]_  | ~\new_[3588]_ ;
  assign \new_[2785]_  = ~\new_[3402]_  | ~\new_[3438]_ ;
  assign \new_[2786]_  = ~\new_[3269]_  | ~\new_[4405]_ ;
  assign \new_[2787]_  = ~\new_[3292]_  | ~\new_[3560]_ ;
  assign \new_[2788]_  = ~\new_[3435]_  | ~\new_[3331]_ ;
  assign \new_[2789]_  = ~\new_[3273]_  | ~\new_[4386]_ ;
  assign \new_[2790]_  = \new_[3509]_  | \new_[3487]_ ;
  assign \new_[2791]_  = ~\new_[3528]_  | ~\new_[3278]_ ;
  assign \new_[2792]_  = ~n1130;
  assign \new_[2793]_  = ~\new_[4380]_  | ~\new_[4384]_ ;
  assign \new_[2794]_  = ~\new_[3281]_  | ~\new_[3418]_ ;
  assign \new_[2795]_  = ~\new_[3588]_  | ~\new_[3270]_ ;
  assign \new_[2796]_  = ~\new_[5289]_  | ~\new_[4380]_ ;
  assign \new_[2797]_  = ~\new_[3492]_  | ~\new_[3319]_ ;
  assign \new_[2798]_  = ~\new_[3485]_  | ~\new_[3329]_ ;
  assign \new_[2799]_  = ~\new_[3485]_  | ~\new_[3401]_ ;
  assign \new_[2800]_  = ~\new_[3406]_  | ~\new_[4784]_ ;
  assign \new_[2801]_  = ~\new_[3269]_  | ~\new_[3501]_ ;
  assign \new_[2802]_  = ~\new_[4402]_  | ~\new_[3438]_ ;
  assign \new_[2803]_  = ~\new_[3300]_  | ~\new_[3403]_ ;
  assign \new_[2804]_  = ~\new_[3254]_  | ~\new_[3560]_ ;
  assign \new_[2805]_  = ~\new_[3332]_  | ~\new_[3292]_ ;
  assign \new_[2806]_  = ~\new_[3592]_  | ~\new_[3530]_ ;
  assign \new_[2807]_  = ~\new_[4383]_  | ~\new_[4402]_ ;
  assign \new_[2808]_  = ~\new_[3419]_  | ~\new_[3707]_ ;
  assign \new_[2809]_  = ~\new_[4395]_  | ~\new_[3279]_ ;
  assign \new_[2810]_  = ~\new_[3511]_  | ~\new_[4384]_ ;
  assign \new_[2811]_  = ~\new_[3186]_  | ~\new_[4386]_ ;
  assign \new_[2812]_  = ~\new_[3186]_  | ~\new_[3492]_ ;
  assign \new_[2813]_  = ~\new_[3269]_  | ~\new_[3305]_ ;
  assign \new_[2814]_  = \new_[5177]_  | \new_[3178]_ ;
  assign \new_[2815]_  = ~\new_[3275]_  | ~\new_[4380]_ ;
  assign \new_[2816]_  = ~\new_[3269]_  | ~\new_[3719]_ ;
  assign \new_[2817]_  = ~\new_[3264]_  | ~\new_[4405]_ ;
  assign \new_[2818]_  = ~\new_[3262]_  | ~\new_[3421]_ ;
  assign \new_[2819]_  = ~\new_[3587]_  | ~\new_[3460]_ ;
  assign \new_[2820]_  = ~\new_[3316]_  | ~\new_[3268]_ ;
  assign \new_[2821]_  = ~\new_[3186]_  | ~\new_[3635]_ ;
  assign \new_[2822]_  = ~\new_[3277]_  | ~\new_[3485]_ ;
  assign \new_[2823]_  = ~\new_[3588]_  | ~\new_[3277]_ ;
  assign \new_[2824]_  = ~\new_[3485]_  | ~\new_[3313]_ ;
  assign \new_[2825]_  = ~\new_[3616]_  | ~\new_[3492]_ ;
  assign \new_[2826]_  = ~\new_[3587]_  | ~\new_[3533]_ ;
  assign \new_[2827]_  = ~\new_[3498]_  | ~\new_[3560]_ ;
  assign \new_[2828]_  = ~\new_[3498]_  | ~\new_[3468]_ ;
  assign \new_[2829]_  = ~\new_[3406]_  | ~\new_[4384]_ ;
  assign \new_[2830]_  = ~\new_[3501]_  | ~\new_[3735]_ ;
  assign \new_[2831]_  = ~\new_[3468]_  | ~\new_[3646]_ ;
  assign \new_[2832]_  = \new_[3582]_  | \new_[3519]_ ;
  assign \new_[2833]_  = ~\new_[3558]_  | ~\new_[3576]_ ;
  assign \new_[2834]_  = ~\new_[4383]_  | ~\new_[4386]_ ;
  assign \new_[2835]_  = ~\new_[3261]_  | ~\new_[3564]_ ;
  assign \new_[2836]_  = ~\new_[3275]_  | ~\new_[3405]_ ;
  assign \new_[2837]_  = ~\new_[3281]_  | ~\new_[3189]_ ;
  assign \new_[2838]_  = ~\new_[3279]_  | ~\new_[3437]_ ;
  assign \new_[2839]_  = ~\new_[3280]_  | ~\new_[3531]_ ;
  assign \new_[2840]_  = ~\new_[3528]_  | ~\new_[3292]_ ;
  assign \new_[2841]_  = ~\new_[3269]_  | ~\new_[3273]_ ;
  assign \new_[2842]_  = ~\new_[3280]_  | ~\new_[3543]_ ;
  assign \new_[2843]_  = ~\new_[3599]_  | ~\new_[3564]_ ;
  assign \new_[2844]_  = ~\new_[4379]_  | ~\new_[3653]_ ;
  assign \new_[2845]_  = \new_[3301]_  | \new_[3483]_ ;
  assign \new_[2846]_  = ~\new_[3717]_  | ~\new_[3319]_ ;
  assign \new_[2847]_  = ~\new_[3588]_  | ~\new_[3599]_ ;
  assign \new_[2848]_  = ~\new_[3148]_ ;
  assign n1120 = ~\new_[4674]_ ;
  assign n1185 = \new_[2992]_ ;
  assign \new_[2851]_  = ~\new_[2992]_ ;
  assign \new_[2852]_  = ~n1145;
  assign \new_[2853]_  = ~n1115;
  assign \new_[2854]_  = (~\new_[3464]_  | ~\new_[3739]_ ) & (~\new_[3713]_  | ~\desIn[43] );
  assign n995 = ~\new_[3756]_  | ~\new_[3288]_ ;
  assign \new_[2856]_  = ~n1150;
  assign n1215 = ~\new_[3147]_ ;
  assign \new_[2858]_  = ~\new_[3172]_  | ~\new_[4242]_ ;
  assign \new_[2859]_  = ~\new_[3194]_  & (~\new_[3379]_  | ~\new_[4207]_ );
  assign \new_[2860]_  = ~\new_[3196]_  & (~\new_[3440]_  | ~\new_[4231]_ );
  assign \new_[2861]_  = ~\new_[3175]_  | ~\new_[4176]_ ;
  assign \new_[2862]_  = ~\new_[3198]_  & (~\new_[3372]_  | ~\new_[4160]_ );
  assign \new_[2863]_  = ~\new_[3185]_  & (~\new_[3376]_  | ~\new_[4276]_ );
  assign \new_[2864]_  = ~\new_[3201]_  & (~\new_[3371]_  | ~\new_[5097]_ );
  assign \new_[2865]_  = ~\new_[4698]_  | ~\new_[3172]_ ;
  assign \new_[2866]_  = ~\new_[3188]_  & (~\new_[3373]_  | ~\new_[4262]_ );
  assign \new_[2867]_  = ~\new_[3203]_  & (~\new_[3375]_  | ~\new_[5175]_ );
  assign \new_[2868]_  = ~\new_[3204]_  & (~\new_[3324]_  | ~\new_[5068]_ );
  assign \new_[2869]_  = ~\new_[4164]_  & (~\new_[5288]_  | ~\new_[3403]_ );
  assign \new_[2870]_  = ~\new_[3175]_  | ~\new_[4222]_ ;
  assign \new_[2871]_  = ~\new_[3713]_ ;
  assign \new_[2872]_  = ~\new_[3713]_ ;
  assign \new_[2873]_  = ~\new_[3207]_  & (~\new_[3363]_  | ~\new_[4231]_ );
  assign \new_[2874]_  = ~\new_[3191]_  & (~\new_[3398]_  | ~\new_[4249]_ );
  assign \new_[2875]_  = ~\new_[3213]_  & (~\new_[3427]_  | ~\new_[4207]_ );
  assign \new_[2876]_  = ~\new_[3337]_  & (~\new_[3339]_  | ~\new_[4231]_ );
  assign \new_[2877]_  = ~\new_[3192]_  & (~\new_[3384]_  | ~\new_[5097]_ );
  assign \new_[2878]_  = ~\new_[3182]_  & (~\new_[3351]_  | ~\new_[4176]_ );
  assign \new_[2879]_  = ~\new_[3200]_  & (~\new_[3366]_  | ~\new_[4222]_ );
  assign \new_[2880]_  = ~\new_[3158]_ ;
  assign \new_[2881]_  = ~\new_[3210]_  & (~\new_[4222]_  | ~\new_[3449]_ );
  assign \new_[2882]_  = ~\new_[3212]_  & (~\new_[3347]_  | ~\new_[4222]_ );
  assign \new_[2883]_  = ~\new_[4211]_  & (~\new_[3479]_  | ~\new_[3529]_ );
  assign \new_[2884]_  = ~\new_[3173]_  | ~\new_[5068]_ ;
  assign \new_[2885]_  = ~\new_[4115]_  & (~\new_[3412]_  | ~\new_[3425]_ );
  assign \new_[2886]_  = ~\new_[3649]_  | ~\new_[3309]_ ;
  assign \new_[2887]_  = ~\new_[3346]_  | ~\new_[4220]_ ;
  assign \new_[2888]_  = ~\new_[3386]_  | ~\new_[4176]_ ;
  assign \new_[2889]_  = ~\new_[3385]_  | ~\new_[4698]_ ;
  assign \new_[2890]_  = ~\new_[3351]_  | ~\new_[4249]_ ;
  assign \new_[2891]_  = ~\new_[3355]_  | ~\new_[4242]_ ;
  assign \new_[2892]_  = ~\new_[3385]_  | ~\new_[4242]_ ;
  assign \new_[2893]_  = ~\new_[3361]_  | ~\new_[4098]_ ;
  assign \new_[2894]_  = ~\new_[3391]_  | ~\new_[4176]_ ;
  assign \new_[2895]_  = ~\new_[3386]_  | ~\new_[4222]_ ;
  assign \new_[2896]_  = ~\new_[3389]_  | ~\new_[4222]_ ;
  assign \new_[2897]_  = ~\new_[3359]_  | ~\new_[4176]_ ;
  assign \new_[2898]_  = ~\new_[3713]_ ;
  assign \new_[2899]_  = ~\new_[3361]_  | ~\new_[4220]_ ;
  assign \new_[2900]_  = ~\new_[3359]_  | ~\new_[4222]_ ;
  assign \new_[2901]_  = ~\new_[3352]_  | ~\new_[4176]_ ;
  assign \new_[2902]_  = ~\new_[3495]_ ;
  assign \new_[2903]_  = ~\new_[3350]_  | ~\new_[4176]_ ;
  assign \new_[2904]_  = ~\new_[3368]_  | ~\new_[4176]_ ;
  assign \new_[2905]_  = ~\new_[3369]_  | ~\new_[4208]_ ;
  assign \new_[2906]_  = ~\new_[4176]_  | ~\new_[3449]_ ;
  assign \new_[2907]_  = ~\new_[3428]_  | ~\new_[3735]_ ;
  assign \new_[2908]_  = \new_[3713]_ ;
  assign \new_[2909]_  = ~\new_[3348]_  | ~\new_[4242]_ ;
  assign \new_[2910]_  = ~\new_[3394]_  | ~\new_[4242]_ ;
  assign \new_[2911]_  = ~\new_[3352]_  | ~\new_[4222]_ ;
  assign \new_[2912]_  = ~\new_[3390]_  | ~\new_[4176]_ ;
  assign \new_[2913]_  = ~\new_[3355]_  | ~\new_[4220]_ ;
  assign \new_[2914]_  = ~\new_[3391]_  | ~\new_[4222]_ ;
  assign \new_[2915]_  = ~\new_[3607]_  | ~\new_[3330]_ ;
  assign \new_[2916]_  = ~\new_[3368]_  | ~\new_[4222]_ ;
  assign \new_[2917]_  = ~\new_[3389]_  | ~\new_[4021]_ ;
  assign \new_[2918]_  = ~\new_[3350]_  | ~\new_[4222]_ ;
  assign \new_[2919]_  = ~\new_[3390]_  | ~\new_[4222]_ ;
  assign \new_[2920]_  = ~\new_[3340]_  | ~\new_[4242]_ ;
  assign \new_[2921]_  = ~\new_[3394]_  | ~\new_[4188]_ ;
  assign \new_[2922]_  = ~\new_[3346]_  | ~\new_[4242]_ ;
  assign \new_[2923]_  = ~\new_[3345]_  | ~\new_[4176]_ ;
  assign \new_[2924]_  = ~\new_[3340]_  | ~\new_[4698]_ ;
  assign \new_[2925]_  = ~\new_[3360]_  | ~\new_[4248]_ ;
  assign \new_[2926]_  = ~\new_[4395]_  | ~\new_[5240]_ ;
  assign \new_[2927]_  = ~\new_[4238]_  & (~\new_[4394]_  | ~\new_[3537]_ );
  assign \new_[2928]_  = ~\new_[4238]_  & (~\new_[3757]_  | ~\new_[3670]_ );
  assign n1135 = ~\new_[3748]_  | ~\new_[3451]_ ;
  assign \new_[2930]_  = ~\new_[3511]_  | ~\new_[3419]_ ;
  assign n1190 = ~\new_[3284]_ ;
  assign \new_[2932]_  = ~\new_[5098]_  & (~\new_[3544]_  | ~\new_[5268]_ );
  assign \new_[2933]_  = ~\new_[3380]_  | ~\new_[4198]_ ;
  assign \new_[2934]_  = ~\new_[3587]_  | ~\new_[3444]_ ;
  assign \new_[2935]_  = ~\new_[4269]_  & (~\new_[4403]_  | ~\new_[3660]_ );
  assign \new_[2936]_  = ~\new_[3588]_  | ~\new_[3329]_ ;
  assign \new_[2937]_  = ~\new_[3473]_  | ~\new_[4198]_ ;
  assign \new_[2938]_  = ~\new_[5174]_  & (~\new_[3532]_  | ~\new_[3738]_ );
  assign \new_[2939]_  = ~\new_[3378]_  | ~\new_[4173]_ ;
  assign \new_[2940]_  = ~\new_[3436]_  | ~\new_[4212]_ ;
  assign \new_[2941]_  = ~\new_[3434]_  | ~\new_[5175]_ ;
  assign \new_[2942]_  = ~\new_[3320]_  | ~\new_[4241]_ ;
  assign \new_[2943]_  = ~\new_[4189]_  & (~\new_[4395]_  | ~\new_[3727]_ );
  assign \new_[2944]_  = ~\new_[5063]_  & (~\new_[3646]_  | ~\new_[3535]_ );
  assign \new_[2945]_  = ~\new_[4259]_  & (~\new_[3592]_  | ~\new_[3727]_ );
  assign \new_[2946]_  = ~\new_[4189]_  & (~\new_[3718]_  | ~\new_[3653]_ );
  assign \new_[2947]_  = ~\new_[3353]_  | ~\new_[4262]_ ;
  assign \new_[2948]_  = ~\new_[3367]_  | ~\new_[4235]_ ;
  assign \new_[2949]_  = ~\new_[3362]_  | ~\new_[4276]_ ;
  assign \new_[2950]_  = ~\new_[3357]_  | ~\new_[5068]_ ;
  assign \new_[2951]_  = ~\new_[3354]_  | ~\new_[4226]_ ;
  assign \new_[2952]_  = ~\new_[3454]_  | ~\new_[3433]_ ;
  assign \new_[2953]_  = ~\new_[3358]_  | ~\new_[4121]_ ;
  assign \new_[2954]_  = ~\new_[3444]_  | ~\new_[3700]_ ;
  assign \new_[2955]_  = ~\new_[4259]_  & (~\new_[4401]_  | ~\new_[3705]_ );
  assign \new_[2956]_  = ~\new_[4259]_  & (~\new_[3726]_  | ~\new_[3610]_ );
  assign \new_[2957]_  = ~\new_[4180]_  & (~\new_[3604]_  | ~\new_[5178]_ );
  assign \new_[2958]_  = ~\new_[5063]_  & (~\new_[3543]_  | ~\new_[3545]_ );
  assign \new_[2959]_  = ~\new_[3628]_  | ~\new_[3422]_ ;
  assign \new_[2960]_  = ~\new_[4189]_  & (~\new_[3544]_  | ~\new_[3658]_ );
  assign \new_[2961]_  = ~\new_[3260]_ ;
  assign \new_[2962]_  = ~\new_[3377]_  | ~\new_[4262]_ ;
  assign \new_[2963]_  = ~\new_[3478]_  | ~\new_[3432]_ ;
  assign \new_[2964]_  = ~\new_[3395]_  | ~\new_[4121]_ ;
  assign \new_[2965]_  = ~\new_[4189]_  & (~\new_[3660]_  | ~\new_[3735]_ );
  assign \new_[2966]_  = ~\new_[3388]_  | ~\new_[4207]_ ;
  assign \new_[2967]_  = ~\new_[4272]_  & (~\new_[4403]_  | ~\new_[3649]_ );
  assign \new_[2968]_  = ~\new_[3322]_  | ~\new_[4215]_ ;
  assign \new_[2969]_  = ~\new_[3382]_  | ~\new_[5068]_ ;
  assign \new_[2970]_  = ~\new_[3356]_  | ~\new_[4235]_ ;
  assign \new_[2971]_  = ~\new_[5182]_  | ~\new_[3684]_ ;
  assign \new_[2972]_  = ~\new_[3305]_  | ~\new_[3735]_ ;
  assign n1140 = ~\new_[3755]_  | ~\new_[3475]_ ;
  assign \new_[2974]_  = ~\new_[4255]_  & (~\new_[3592]_  | ~\new_[3725]_ );
  assign \new_[2975]_  = ~\new_[4164]_  & (~\new_[3587]_  | ~\new_[3524]_ );
  assign \new_[2976]_  = ~\new_[3311]_  | ~\new_[4231]_ ;
  assign n1130 = ~\new_[3751]_  | ~\new_[3452]_ ;
  assign \new_[2978]_  = ~\new_[3259]_ ;
  assign \new_[2979]_  = ~\new_[4115]_  & (~\new_[3530]_  | ~\new_[4785]_ );
  assign \new_[2980]_  = ~\new_[3343]_  | ~\new_[4140]_ ;
  assign \new_[2981]_  = ~\new_[3318]_  | ~\new_[4186]_ ;
  assign \new_[2982]_  = ~\new_[3396]_  | ~\new_[4121]_ ;
  assign \new_[2983]_  = ~\new_[4264]_  & (~\new_[3533]_  | ~\new_[3614]_ );
  assign \new_[2984]_  = ~\new_[3335]_  | ~\new_[4176]_ ;
  assign \new_[2985]_  = ~\new_[3455]_  | ~\new_[4226]_ ;
  assign \new_[2986]_  = ~\new_[3374]_  | ~\new_[4215]_ ;
  assign \new_[2987]_  = ~\new_[3349]_  | ~\new_[4235]_ ;
  assign \new_[2988]_  = ~\new_[3370]_  | ~\new_[4276]_ ;
  assign \new_[2989]_  = ~\new_[4247]_  & (~\new_[3591]_  | ~\new_[3638]_ );
  assign \new_[2990]_  = ~\new_[3397]_  | ~\new_[4262]_ ;
  assign \new_[2991]_  = ~\new_[3342]_  | ~\new_[5068]_ ;
  assign \new_[2992]_  = ~\new_[3698]_  | (~\new_[3568]_  & ~\new_[3837]_ );
  assign \new_[2993]_  = ~\new_[3428]_  | ~\new_[3443]_ ;
  assign \new_[2994]_  = ~\new_[3433]_  | ~\new_[3417]_ ;
  assign \new_[2995]_  = ~\new_[4403]_  | ~\new_[3305]_ ;
  assign \new_[2996]_  = ~\new_[3628]_  | ~\new_[3458]_ ;
  assign \new_[2997]_  = ~\new_[3454]_  | ~\new_[3315]_ ;
  assign \new_[2998]_  = ~\new_[4657]_  | ~\new_[3727]_ ;
  assign \new_[2999]_  = ~\new_[3714]_  | ~\new_[3738]_ ;
  assign \new_[3000]_  = ~\new_[3419]_  | ~\new_[5240]_ ;
  assign \new_[3001]_  = ~\new_[3331]_  | ~\new_[3405]_ ;
  assign \new_[3002]_  = ~\new_[3305]_  | ~\new_[3402]_ ;
  assign \new_[3003]_  = ~\new_[5273]_  | ~\new_[3527]_ ;
  assign \new_[3004]_  = ~\new_[3221]_ ;
  assign \new_[3005]_  = ~\new_[3310]_  | ~\new_[3735]_ ;
  assign \new_[3006]_  = ~\new_[3471]_  | ~\new_[4785]_ ;
  assign \new_[3007]_  = ~\new_[3515]_  | ~\new_[3414]_ ;
  assign \new_[3008]_  = ~\new_[4785]_  | ~\new_[5240]_ ;
  assign \new_[3009]_  = ~\new_[3406]_  | ~\new_[5263]_ ;
  assign \new_[3010]_  = ~\new_[3310]_  | ~\new_[4386]_ ;
  assign \new_[3011]_  = ~\new_[3399]_  | ~\new_[3753]_ ;
  assign \new_[3012]_  = ~\new_[3718]_  | ~\new_[3481]_ ;
  assign \new_[3013]_  = ~\new_[3444]_  | ~\new_[3738]_ ;
  assign \new_[3014]_  = ~\new_[4395]_  | ~\new_[3416]_ ;
  assign \new_[3015]_  = ~\new_[3305]_  | ~\new_[3643]_ ;
  assign \new_[3016]_  = ~\new_[3558]_  | ~\new_[3490]_ ;
  assign \new_[3017]_  = ~\new_[3442]_  | ~\new_[3673]_ ;
  assign \new_[3018]_  = ~\new_[3437]_  | ~\new_[5240]_ ;
  assign \new_[3019]_  = ~\new_[3517]_  | ~\new_[3719]_ ;
  assign \new_[3020]_  = ~\new_[3331]_  | ~\new_[4379]_ ;
  assign \new_[3021]_  = ~\new_[3315]_  | ~\new_[3456]_ ;
  assign \new_[3022]_  = ~\new_[3482]_  | ~\new_[3670]_ ;
  assign \new_[3023]_  = ~\new_[3576]_  | ~\new_[3471]_ ;
  assign \new_[3024]_  = ~\new_[3341]_  | ~\new_[4657]_ ;
  assign \new_[3025]_  = ~\new_[3400]_  | ~\new_[3524]_ ;
  assign \new_[3026]_  = ~\new_[3587]_  | ~\new_[3485]_ ;
  assign \new_[3027]_  = ~\new_[3717]_  | ~\new_[3429]_ ;
  assign \new_[3028]_  = ~\new_[4380]_  | ~\new_[5263]_ ;
  assign \new_[3029]_  = ~\new_[3591]_  | ~\new_[3624]_ ;
  assign \new_[3030]_  = ~\new_[3422]_  | ~\new_[5272]_ ;
  assign \new_[3031]_  = ~\new_[3581]_  | ~\new_[3658]_ ;
  assign \new_[3032]_  = ~\new_[3442]_  | ~\new_[3524]_ ;
  assign \new_[3033]_  = ~\new_[3312]_  | ~\new_[3319]_ ;
  assign \new_[3034]_  = ~\new_[3604]_  | ~\new_[3438]_ ;
  assign \new_[3035]_  = ~\new_[3456]_  | ~\new_[3645]_ ;
  assign \new_[3036]_  = ~\new_[3456]_  | ~\new_[3535]_ ;
  assign \new_[3037]_  = ~\new_[3674]_  | ~\new_[3758]_ ;
  assign \new_[3038]_  = ~\new_[3479]_  | ~\new_[3673]_ ;
  assign \new_[3039]_  = \new_[3431]_  | \new_[3721]_ ;
  assign \new_[3040]_  = ~\new_[3418]_  | ~\new_[3488]_ ;
  assign \new_[3041]_  = ~\new_[3444]_  | ~\new_[3527]_ ;
  assign \new_[3042]_  = ~\new_[3314]_  | ~\new_[3326]_ ;
  assign \new_[3043]_  = ~\new_[3469]_  | ~\new_[3615]_ ;
  assign \new_[3044]_  = ~\new_[3313]_  | ~\new_[3723]_ ;
  assign \new_[3045]_  = ~\new_[3683]_  | ~\new_[3673]_ ;
  assign \new_[3046]_  = ~\new_[3333]_  | ~\new_[3658]_ ;
  assign \new_[3047]_  = ~\new_[3482]_  | ~\new_[3720]_ ;
  assign \new_[3048]_  = ~\new_[3472]_  | ~\new_[4387]_ ;
  assign \new_[3049]_  = ~\new_[3485]_  | ~\new_[3327]_ ;
  assign \new_[3050]_  = ~\new_[3545]_  | ~\new_[5240]_ ;
  assign \new_[3051]_  = ~\new_[3438]_  | ~\new_[3615]_ ;
  assign \new_[3052]_  = ~\new_[3333]_  | ~\new_[3608]_ ;
  assign \new_[3053]_  = ~\new_[3629]_  | ~\new_[3403]_ ;
  assign \new_[3054]_  = ~\new_[3610]_  | ~\new_[3429]_ ;
  assign \new_[3055]_  = ~\new_[3437]_  | ~\new_[3530]_ ;
  assign \new_[3056]_  = ~\new_[5269]_  | ~\new_[3330]_ ;
  assign \new_[3057]_  = ~\new_[3465]_  | ~\new_[3545]_ ;
  assign \new_[3058]_  = ~\new_[3315]_  | ~\new_[3417]_ ;
  assign \new_[3059]_  = ~\new_[3718]_  | ~\new_[4785]_ ;
  assign \new_[3060]_  = ~\new_[3450]_  | ~\new_[3631]_ ;
  assign \new_[3061]_  = ~\new_[3638]_  | ~\new_[3650]_ ;
  assign \new_[3062]_  = ~\new_[3490]_  | ~\new_[3406]_ ;
  assign \new_[3063]_  = ~\new_[3611]_  | ~\new_[3614]_ ;
  assign \new_[3064]_  = ~\new_[3305]_  | ~\new_[3443]_ ;
  assign \new_[3065]_  = ~\new_[3485]_  | ~\new_[3527]_ ;
  assign \new_[3066]_  = ~\new_[3403]_  | ~\new_[4785]_ ;
  assign \new_[3067]_  = ~\new_[4380]_  | ~\new_[3437]_ ;
  assign \new_[3068]_  = ~\new_[3503]_  | ~\new_[3387]_ ;
  assign \new_[3069]_  = ~\new_[3719]_  | ~\new_[4386]_ ;
  assign \new_[3070]_  = ~\new_[3646]_  | ~\new_[3560]_ ;
  assign \new_[3071]_  = ~\new_[3614]_  | ~\new_[3624]_ ;
  assign \new_[3072]_  = ~\new_[3420]_  | ~\new_[3700]_ ;
  assign \new_[3073]_  = ~\new_[3321]_  | ~\new_[5182]_ ;
  assign \new_[3074]_  = ~\new_[5260]_  | ~\new_[3333]_ ;
  assign \new_[3075]_  = ~\new_[4657]_  | ~\new_[3718]_ ;
  assign \new_[3076]_  = ~\new_[3471]_  | ~\new_[3653]_ ;
  assign \new_[3077]_  = ~\new_[3490]_  | ~\new_[3636]_ ;
  assign \new_[3078]_  = ~\new_[3450]_  | ~\new_[3437]_ ;
  assign \new_[3079]_  = ~\new_[3418]_  | ~\new_[3735]_ ;
  assign \new_[3080]_  = ~\new_[3705]_  | ~\new_[3488]_ ;
  assign \new_[3081]_  = ~\new_[3709]_  | ~\new_[3341]_ ;
  assign \new_[3082]_  = ~\new_[3511]_  | ~\new_[3331]_ ;
  assign \new_[3083]_  = ~\new_[3628]_  | ~\new_[3480]_ ;
  assign \new_[3084]_  = ~\new_[3456]_  | ~\new_[3407]_ ;
  assign \new_[3085]_  = ~\new_[3406]_  | ~\new_[5289]_ ;
  assign \new_[3086]_  = ~\new_[3640]_  | ~\new_[3727]_ ;
  assign \new_[3087]_  = ~\new_[3683]_  | ~\new_[5272]_ ;
  assign \new_[3088]_  = ~\new_[3442]_  | ~\new_[5273]_ ;
  assign \new_[3089]_  = ~\new_[4863]_  | ~\new_[3419]_ ;
  assign \new_[3090]_  = ~\new_[3537]_  | ~\new_[4384]_ ;
  assign \new_[3091]_  = ~\new_[3468]_  | ~\new_[3447]_ ;
  assign \new_[3092]_  = ~\new_[3490]_  | ~\new_[3707]_ ;
  assign \new_[3093]_  = ~\new_[3622]_  | ~\new_[3430]_ ;
  assign \new_[3094]_  = ~\new_[3511]_  | ~\new_[4393]_ ;
  assign \new_[3095]_  = ~\new_[4863]_  | ~\new_[4657]_ ;
  assign \new_[3096]_  = ~\new_[3407]_  | ~\new_[3404]_ ;
  assign \new_[3097]_  = ~\new_[3663]_  | ~\new_[3330]_ ;
  assign \new_[3098]_  = \new_[3467]_  | \new_[3598]_ ;
  assign \new_[3099]_  = ~\new_[3725]_  | ~\new_[3629]_ ;
  assign \new_[3100]_  = ~\new_[3664]_  | ~\new_[3603]_ ;
  assign \new_[3101]_  = ~\new_[3488]_  | ~\new_[3438]_ ;
  assign \new_[3102]_  = ~\new_[3482]_  | ~\new_[3387]_ ;
  assign \new_[3103]_  = ~\new_[3644]_  | ~\new_[3447]_ ;
  assign \new_[3104]_  = ~\new_[3305]_  | ~\new_[3610]_ ;
  assign \new_[3105]_  = ~\new_[3312]_  | ~\new_[3428]_ ;
  assign \new_[3106]_  = ~\new_[5178]_  | ~\new_[3443]_ ;
  assign \new_[3107]_  = ~\new_[4657]_  | ~\new_[3730]_ ;
  assign \new_[3108]_  = ~\new_[3418]_  | ~\new_[3309]_ ;
  assign \new_[3109]_  = ~\new_[3693]_  | ~\new_[3667]_ ;
  assign \new_[3110]_  = ~\new_[5178]_  | ~\new_[4387]_ ;
  assign \new_[3111]_  = ~\new_[3457]_  | ~\new_[3433]_ ;
  assign \new_[3112]_  = ~\new_[5181]_  | ~\new_[3472]_ ;
  assign \new_[3113]_  = ~\new_[3426]_  | ~\new_[3416]_ ;
  assign \new_[3114]_  = ~\new_[3753]_  | ~\new_[3675]_ ;
  assign \new_[3115]_  = ~\new_[3607]_  | ~\new_[3409]_ ;
  assign \new_[3116]_  = ~\new_[3700]_  | ~\new_[3430]_ ;
  assign \new_[3117]_  = ~\new_[3387]_  | ~\new_[3407]_ ;
  assign \new_[3118]_  = ~\new_[3640]_  | ~\new_[3707]_ ;
  assign \new_[3119]_  = ~\new_[3309]_  | ~\new_[3415]_ ;
  assign \new_[3120]_  = ~\new_[3471]_  | ~\new_[4385]_ ;
  assign \new_[3121]_  = ~\new_[3643]_  | ~\new_[3319]_ ;
  assign \new_[3122]_  = ~\new_[3616]_  | ~\new_[3643]_ ;
  assign \new_[3123]_  = ~\new_[3481]_  | ~\new_[3727]_ ;
  assign \new_[3124]_  = ~\new_[3616]_  | ~\new_[3488]_ ;
  assign \new_[3125]_  = ~\new_[3660]_  | ~\new_[3402]_ ;
  assign \new_[3126]_  = ~\new_[3684]_  | ~\new_[3716]_ ;
  assign \new_[3127]_  = ~\new_[3484]_  | ~\new_[3643]_ ;
  assign \new_[3128]_  = ~\new_[3663]_  | ~\new_[3457]_ ;
  assign \new_[3129]_  = ~\new_[3614]_  | ~\new_[3430]_ ;
  assign \new_[3130]_  = ~\new_[4402]_  | ~\new_[3415]_ ;
  assign \new_[3131]_  = ~\new_[3694]_  | ~\new_[3528]_ ;
  assign \new_[3132]_  = ~\new_[5273]_  | ~\new_[3738]_ ;
  assign \new_[3133]_  = ~\new_[3472]_  | ~\new_[3517]_ ;
  assign \new_[3134]_  = ~\new_[3479]_  | ~\new_[5279]_ ;
  assign \new_[3135]_  = ~\new_[3607]_  | ~\new_[3308]_ ;
  assign \new_[3136]_  = ~\new_[3470]_  | ~\new_[3640]_ ;
  assign \new_[3137]_  = ~\new_[3621]_  | ~\new_[3429]_ ;
  assign \new_[3138]_  = ~\new_[3444]_  | ~\new_[3326]_ ;
  assign \new_[3139]_  = ~\new_[3314]_  | ~\new_[3625]_ ;
  assign \new_[3140]_  = ~\new_[3306]_  | ~\new_[3664]_ ;
  assign \new_[3141]_  = ~\new_[3305]_  | ~\new_[3488]_ ;
  assign \new_[3142]_  = ~\new_[3444]_  | ~\new_[3458]_ ;
  assign \new_[3143]_  = ~\new_[3314]_  | ~\new_[3667]_ ;
  assign \new_[3144]_  = ~\new_[4790]_  | ~\new_[4384]_ ;
  assign \new_[3145]_  = ~\new_[3425]_  | ~\new_[3408]_ ;
  assign \new_[3146]_  = ~\new_[3254]_ ;
  assign \new_[3147]_  = \new_[3256]_ ;
  assign \new_[3148]_  = ~\new_[3402]_ ;
  assign \new_[3149]_  = ~\new_[3256]_ ;
  assign \new_[3150]_  = ~\new_[5182]_  | ~\new_[3438]_ ;
  assign \new_[3151]_  = ~\new_[3302]_ ;
  assign \new_[3152]_  = ~\new_[3296]_ ;
  assign \new_[3153]_  = ~\new_[3296]_ ;
  assign \new_[3154]_  = ~\new_[3286]_ ;
  assign \new_[3155]_  = ~\new_[3500]_ ;
  assign \new_[3156]_  = ~\new_[3178]_ ;
  assign \new_[3157]_  = ~\new_[3495]_ ;
  assign \new_[3158]_  = ~\new_[3438]_ ;
  assign \new_[3159]_  = ~\new_[3713]_  & (~\new_[3686]_  | ~\new_[3577]_ );
  assign \new_[3160]_  = ~\new_[3364]_  | ~\new_[4276]_ ;
  assign \new_[3161]_  = ~\new_[3416]_  | ~\new_[3481]_ ;
  assign n1225 = ~\new_[3627]_  | (~\new_[3551]_  & ~\new_[3713]_ );
  assign n1220 = ~\new_[3290]_ ;
  assign \new_[3164]_  = ~\new_[3460]_ ;
  assign \new_[3165]_  = ~\new_[3267]_ ;
  assign \new_[3166]_  = ~\new_[3277]_ ;
  assign \new_[3167]_  = ~\new_[4244]_  & (~\new_[3498]_  | ~\new_[3645]_ );
  assign \new_[3168]_  = ~\new_[3638]_  | ~\new_[3453]_ ;
  assign \new_[3169]_  = ~\new_[3490]_  | ~\new_[3470]_ ;
  assign \new_[3170]_  = ~\new_[3301]_ ;
  assign \new_[3171]_  = ~\new_[3412]_  | ~\new_[3315]_ ;
  assign \new_[3172]_  = ~\new_[3529]_  | ~\new_[3650]_ ;
  assign \new_[3173]_  = ~\new_[3529]_  | ~\new_[3738]_ ;
  assign \new_[3174]_  = ~\new_[3413]_ ;
  assign \new_[3175]_  = ~\new_[3614]_  | ~\new_[3529]_ ;
  assign \new_[3176]_  = ~\new_[3526]_  | ~\new_[4242]_ ;
  assign \new_[3177]_  = ~\new_[3521]_  | ~\new_[3625]_ ;
  assign \new_[3178]_  = ~\new_[3309]_ ;
  assign \new_[3179]_  = ~\new_[3536]_  | ~\new_[4242]_ ;
  assign \new_[3180]_  = ~\new_[3667]_  | ~\new_[3529]_ ;
  assign \new_[3181]_  = ~\new_[3591]_  | ~\new_[5278]_ ;
  assign \new_[3182]_  = ~\new_[5098]_  & (~\new_[3631]_  | ~\new_[3637]_ );
  assign \new_[3183]_  = ~\new_[5098]_  & (~\new_[3614]_  | ~\new_[5279]_ );
  assign \new_[3184]_  = ~\new_[5174]_  & (~\new_[3604]_  | ~\new_[3649]_ );
  assign \new_[3185]_  = ~\new_[4269]_  & (~\new_[5272]_  | ~\new_[3706]_ );
  assign \new_[3186]_  = ~\new_[3411]_ ;
  assign \new_[3187]_  = ~\new_[3411]_ ;
  assign \new_[3188]_  = ~\new_[4269]_  & (~\new_[3674]_  | ~\new_[3733]_ );
  assign \new_[3189]_  = ~\new_[3410]_ ;
  assign \new_[3190]_  = ~\new_[4178]_  & (~\new_[3638]_  | ~\new_[3706]_ );
  assign \new_[3191]_  = ~\new_[5098]_  & (~\new_[3673]_  | ~\new_[3738]_ );
  assign \new_[3192]_  = ~\new_[4259]_  & (~\new_[3673]_  | ~\new_[3612]_ );
  assign \new_[3193]_  = ~\new_[4150]_  & (~\new_[5280]_  | ~\new_[3720]_ );
  assign \new_[3194]_  = ~\new_[4792]_  & (~\new_[5100]_  | ~\new_[3719]_ );
  assign \new_[3195]_  = ~\new_[4164]_  & (~\new_[5276]_  | ~\new_[3619]_ );
  assign \new_[3196]_  = ~\new_[4189]_  & (~\new_[3636]_  | ~\new_[3640]_ );
  assign \new_[3197]_  = ~\new_[4259]_  & (~\new_[3649]_  | ~\new_[3735]_ );
  assign \new_[3198]_  = ~\new_[4272]_  & (~\new_[5257]_  | ~\new_[3760]_ );
  assign \new_[3199]_  = \new_[3326]_ ;
  assign \new_[3200]_  = ~\new_[4272]_  & (~\new_[3662]_  | ~\new_[5276]_ );
  assign \new_[3201]_  = ~\new_[4268]_  & (~\new_[3616]_  | ~\new_[3604]_ );
  assign \new_[3202]_  = ~\new_[4259]_  & (~\new_[4863]_  | ~\new_[4762]_ );
  assign \new_[3203]_  = ~\new_[4264]_  & (~\new_[3665]_  | ~\new_[5280]_ );
  assign \new_[3204]_  = ~\new_[4167]_  & (~\new_[3638]_  | ~\new_[3701]_ );
  assign \new_[3205]_  = ~\new_[4792]_  & (~\new_[3610]_  | ~\new_[3660]_ );
  assign \new_[3206]_  = ~\new_[3576]_  | ~\new_[3727]_ ;
  assign \new_[3207]_  = ~\new_[4268]_  & (~\new_[5276]_  | ~\new_[3715]_ );
  assign \new_[3208]_  = ~\new_[4792]_  & (~\new_[4403]_  | ~\new_[3620]_ );
  assign \new_[3209]_  = ~\new_[3512]_  | ~\new_[4222]_ ;
  assign \new_[3210]_  = ~\new_[4189]_  & (~\new_[3760]_  | ~\new_[3648]_ );
  assign \new_[3211]_  = ~\new_[4189]_  & (~\new_[3665]_  | ~\new_[3663]_ );
  assign \new_[3212]_  = ~\new_[4268]_  & (~\new_[3700]_  | ~\new_[3723]_ );
  assign \new_[3213]_  = ~\new_[4272]_  & (~\new_[3664]_  | ~\new_[3753]_ );
  assign \new_[3214]_  = ~\new_[4259]_  & (~\new_[3670]_  | ~\new_[3608]_ );
  assign \new_[3215]_  = ~\new_[3663]_  | ~\new_[3670]_ ;
  assign \new_[3216]_  = ~\new_[3344]_ ;
  assign \new_[3217]_  = ~\new_[3344]_ ;
  assign \new_[3218]_  = ~\new_[3511]_  | ~\new_[3653]_ ;
  assign \new_[3219]_  = ~\new_[3544]_  | ~\new_[3608]_ ;
  assign \new_[3220]_  = ~\new_[3527]_  | ~\new_[3723]_ ;
  assign \new_[3221]_  = ~\new_[3304]_ ;
  assign \new_[3222]_  = ~\new_[3492]_  | ~\new_[3652]_ ;
  assign \new_[3223]_  = ~\new_[4396]_  | ~\new_[4380]_ ;
  assign \new_[3224]_  = ~\new_[3726]_  | ~\new_[3618]_ ;
  assign \new_[3225]_  = ~\new_[3542]_  | ~\new_[3608]_ ;
  assign \new_[3226]_  = ~\new_[3601]_  | ~\new_[3730]_ ;
  assign \new_[3227]_  = ~\new_[3642]_  | (~\new_[3641]_  & ~\new_[3818]_ );
  assign \new_[3228]_  = ~\new_[3591]_  | ~\new_[3533]_ ;
  assign \new_[3229]_  = ~\new_[3591]_  | ~\new_[3723]_ ;
  assign \new_[3230]_  = ~\new_[3492]_  | ~\new_[3649]_ ;
  assign \new_[3231]_  = ~\new_[3496]_  | ~\new_[3541]_ ;
  assign \new_[3232]_  = ~\new_[3515]_  | ~\new_[3758]_ ;
  assign \new_[3233]_  = ~\new_[3734]_  | ~\new_[3637]_ ;
  assign \new_[3234]_  = ~\new_[3665]_  | ~\new_[3753]_ ;
  assign \new_[3235]_  = ~\new_[3542]_  | ~\new_[3757]_ ;
  assign \new_[3236]_  = ~\new_[4396]_  | ~\new_[3725]_ ;
  assign \new_[3237]_  = ~\new_[3542]_  | ~\new_[3753]_ ;
  assign \new_[3238]_  = ~\new_[5276]_  | ~\new_[3576]_ ;
  assign \new_[3239]_  = ~\new_[4382]_  | ~\new_[3492]_ ;
  assign \new_[3240]_  = ~\new_[3515]_  | ~\new_[3581]_ ;
  assign \new_[3241]_  = ~\new_[3599]_  | ~\new_[3723]_ ;
  assign \new_[3242]_  = ~\new_[3541]_  | ~\new_[3735]_ ;
  assign \new_[3243]_  = ~\new_[3717]_  | ~\new_[3508]_ ;
  assign \new_[3244]_  = ~\new_[5269]_  | ~\new_[3670]_ ;
  assign \new_[3245]_  = ~\new_[3622]_  | ~\new_[3521]_ ;
  assign \new_[3246]_  = ~\new_[3544]_  | ~\new_[3515]_ ;
  assign \new_[3247]_  = ~\new_[3504]_  | ~\new_[3729]_ ;
  assign \new_[3248]_  = ~\new_[3511]_  | ~\new_[4785]_ ;
  assign \new_[3249]_  = ~\new_[3622]_  | ~\new_[3638]_ ;
  assign \new_[3250]_  = ~\new_[5277]_  | ~\new_[3631]_ ;
  assign \new_[3251]_  = ~\new_[3544]_  | ~\new_[3644]_ ;
  assign \new_[3252]_  = ~\new_[3622]_  | ~\new_[3723]_ ;
  assign \new_[3253]_  = ~\new_[3725]_  | ~\new_[5263]_ ;
  assign \new_[3254]_  = \new_[3330]_ ;
  assign \new_[3255]_  = \new_[3401]_ ;
  assign \new_[3256]_  = ~\new_[3575]_  & (~\new_[3747]_  | ~\new_[3831]_ );
  assign \new_[3257]_  = \new_[3465]_ ;
  assign \new_[3258]_  = ~\new_[3492]_  | ~\new_[3541]_ ;
  assign \new_[3259]_  = ~\new_[3319]_ ;
  assign \new_[3260]_  = ~\new_[3409]_ ;
  assign \new_[3261]_  = ~\new_[3323]_ ;
  assign \new_[3262]_  = ~\new_[3338]_ ;
  assign \new_[3263]_  = \new_[3415]_ ;
  assign \new_[3264]_  = ~\new_[3486]_ ;
  assign \new_[3265]_  = \new_[3482]_ ;
  assign \new_[3266]_  = \new_[3479]_ ;
  assign \new_[3267]_  = ~\new_[3458]_ ;
  assign \new_[3268]_  = \new_[3407]_ ;
  assign \new_[3269]_  = ~\new_[3325]_ ;
  assign \new_[3270]_  = \new_[3327]_ ;
  assign \new_[3271]_  = \new_[3428]_ ;
  assign \new_[3272]_  = ~\new_[3744]_  | ~\new_[3579]_  | ~\new_[3697]_ ;
  assign \new_[3273]_  = ~\new_[3424]_ ;
  assign \new_[3274]_  = ~\new_[3689]_  | ~\new_[3687]_  | ~\new_[3806]_ ;
  assign \new_[3275]_  = \new_[3490]_ ;
  assign \new_[3276]_  = \new_[3481]_ ;
  assign \new_[3277]_  = ~\new_[3439]_ ;
  assign \new_[3278]_  = ~\new_[3467]_ ;
  assign \new_[3279]_  = \new_[3470]_ ;
  assign \new_[3280]_  = ~\new_[3445]_ ;
  assign \new_[3281]_  = ~\new_[3448]_ ;
  assign n1240 = ~\new_[4905]_ ;
  assign \new_[3283]_  = ~\new_[3576]_  | ~\new_[3639]_ ;
  assign \new_[3284]_  = ~\new_[3795]_  & ~\new_[3572]_ ;
  assign \new_[3285]_  = ~\new_[3591]_  | ~\new_[3678]_ ;
  assign \new_[3286]_  = ~\new_[3423]_ ;
  assign \new_[3287]_  = ~\new_[4115]_  & (~\new_[3607]_  | ~\new_[3676]_ );
  assign \new_[3288]_  = ~\new_[3506]_  | ~\new_[3809]_ ;
  assign \new_[3289]_  = ~\new_[3609]_  | ~\new_[3688]_  | ~\new_[3803]_ ;
  assign \new_[3290]_  = (~\new_[3606]_  | ~\new_[3987]_ ) & (~\new_[3914]_  | ~\desIn[31] );
  assign \new_[3291]_  = \new_[2025]_  ? \new_[3712]_  : \new_[3695]_ ;
  assign \new_[3292]_  = \new_[3447]_ ;
  assign \new_[3293]_  = ~\new_[3677]_ ;
  assign \new_[3294]_  = \new_[2024]_  ? \new_[3712]_  : \new_[3647]_ ;
  assign \new_[3295]_  = (~\new_[3696]_  | ~\new_[3818]_ ) & (~\new_[3754]_  | ~\new_[2018]_ );
  assign \new_[3296]_  = ~\new_[3420]_ ;
  assign \new_[3297]_  = ~\new_[3629]_  | ~\new_[3707]_ ;
  assign \new_[3298]_  = ~\new_[3544]_  | ~\new_[3607]_ ;
  assign \new_[3299]_  = ~\new_[3441]_ ;
  assign \new_[3300]_  = ~\new_[3477]_ ;
  assign \new_[3301]_  = ~\new_[5263]_ ;
  assign \new_[3302]_  = ~\new_[3417]_ ;
  assign \new_[3303]_  = \new_[2348]_  ? \new_[5307]_  : \new_[444]_ ;
  assign \new_[3304]_  = ~\new_[3523]_ ;
  assign \new_[3305]_  = ~\new_[3493]_ ;
  assign \new_[3306]_  = ~\new_[3567]_ ;
  assign \new_[3307]_  = ~\new_[3528]_ ;
  assign \new_[3308]_  = ~\new_[3494]_ ;
  assign \new_[3309]_  = ~\new_[3513]_ ;
  assign \new_[3310]_  = ~\new_[3555]_ ;
  assign \new_[3311]_  = ~\new_[3665]_  | ~\new_[3603]_ ;
  assign \new_[3312]_  = ~\new_[3513]_ ;
  assign \new_[3313]_  = ~\new_[3556]_ ;
  assign \new_[3314]_  = ~\new_[3554]_ ;
  assign \new_[3315]_  = ~\new_[3567]_ ;
  assign \new_[3316]_  = \new_[3581]_ ;
  assign \new_[3317]_  = ~\new_[5098]_  & (~\new_[3736]_  | ~\new_[3730]_ );
  assign \new_[3318]_  = ~\new_[3663]_  | ~\new_[3758]_ ;
  assign \new_[3319]_  = ~\new_[3539]_ ;
  assign \new_[3320]_  = ~\new_[3694]_  | ~\new_[5281]_ ;
  assign \new_[3321]_  = ~\new_[3507]_ ;
  assign \new_[3322]_  = ~\new_[4863]_  | ~\new_[3653]_ ;
  assign \new_[3323]_  = ~\new_[3622]_ ;
  assign \new_[3324]_  = ~\new_[3607]_  | ~\new_[3664]_ ;
  assign \new_[3325]_  = ~\new_[3621]_ ;
  assign \new_[3326]_  = ~\new_[3593]_ ;
  assign \new_[3327]_  = ~\new_[3553]_ ;
  assign \new_[3328]_  = ~\new_[3685]_  | ~\new_[3809]_ ;
  assign \new_[3329]_  = ~\new_[3593]_ ;
  assign \new_[3330]_  = ~\new_[3499]_ ;
  assign \new_[3331]_  = ~\new_[3552]_ ;
  assign \new_[3332]_  = \new_[3515]_ ;
  assign \new_[3333]_  = ~\new_[3510]_ ;
  assign \new_[3334]_  = ~\new_[3664]_  | ~\new_[3663]_ ;
  assign \new_[3335]_  = ~\new_[3628]_  | ~\new_[3612]_ ;
  assign \new_[3336]_  = ~\new_[3497]_ ;
  assign \new_[3337]_  = ~\new_[4792]_  & (~\new_[3738]_  | ~\new_[3723]_ );
  assign \new_[3338]_  = ~\new_[3653]_ ;
  assign \new_[3339]_  = ~\new_[5278]_  | ~\new_[3625]_ ;
  assign \new_[3340]_  = ~\new_[3657]_  | ~\new_[3678]_ ;
  assign \new_[3341]_  = ~\new_[3540]_ ;
  assign \new_[3342]_  = ~\new_[5259]_  | ~\new_[5257]_ ;
  assign \new_[3343]_  = ~\new_[3694]_  | ~\new_[3753]_ ;
  assign \new_[3344]_  = ~\new_[3529]_ ;
  assign \new_[3345]_  = ~\new_[3611]_  | ~\new_[3706]_ ;
  assign \new_[3346]_  = ~\new_[5268]_  | ~\new_[3720]_ ;
  assign \new_[3347]_  = ~\new_[3626]_  | ~\new_[3624]_ ;
  assign \new_[3348]_  = ~\new_[3654]_  | ~\new_[3653]_ ;
  assign \new_[3349]_  = ~\new_[5255]_  | ~\new_[3611]_ ;
  assign \new_[3350]_  = ~\new_[3725]_  | ~\new_[3619]_ ;
  assign \new_[3351]_  = ~\new_[4863]_  | ~\new_[3736]_ ;
  assign \new_[3352]_  = ~\new_[3662]_  | ~\new_[3707]_ ;
  assign \new_[3353]_  = ~\new_[3724]_  | ~\new_[3656]_ ;
  assign \new_[3354]_  = ~\new_[5268]_  | ~\new_[3676]_ ;
  assign \new_[3355]_  = ~\new_[3616]_  | ~\new_[3635]_ ;
  assign \new_[3356]_  = ~\new_[4762]_  | ~\new_[3623]_ ;
  assign \new_[3357]_  = ~\new_[3605]_  | ~\new_[3623]_ ;
  assign \new_[3358]_  = ~\new_[3665]_  | ~\new_[3674]_ ;
  assign \new_[3359]_  = ~\new_[3701]_  | ~\new_[3723]_ ;
  assign \new_[3360]_  = ~\new_[3671]_  | ~\new_[3709]_ ;
  assign \new_[3361]_  = ~\new_[3709]_  | ~\new_[3636]_ ;
  assign \new_[3362]_  = ~\new_[5277]_  | ~\new_[3734]_ ;
  assign \new_[3363]_  = ~\new_[3604]_  | ~\new_[3660]_ ;
  assign \new_[3364]_  = ~\new_[3717]_  | ~\new_[3656]_ ;
  assign \new_[3365]_  = ~\new_[5272]_  | ~\new_[3650]_ ;
  assign \new_[3366]_  = ~\new_[3613]_  | ~\new_[3652]_ ;
  assign \new_[3367]_  = ~\new_[3726]_  | ~\new_[3604]_ ;
  assign \new_[3368]_  = ~\new_[3616]_  | ~\new_[3729]_ ;
  assign \new_[3369]_  = ~\new_[3662]_  | ~\new_[3730]_ ;
  assign \new_[3370]_  = ~\new_[5268]_  | ~\new_[3733]_ ;
  assign \new_[3371]_  = ~\new_[3717]_  | ~\new_[3705]_ ;
  assign \new_[3372]_  = ~\new_[5281]_  | ~\new_[3676]_ ;
  assign \new_[3373]_  = ~\new_[3626]_  | ~\new_[3611]_ ;
  assign \new_[3374]_  = ~\new_[3714]_  | ~\new_[3683]_ ;
  assign \new_[3375]_  = ~\new_[3694]_  | ~\new_[3757]_ ;
  assign \new_[3376]_  = ~\new_[3667]_  | ~\new_[5278]_ ;
  assign \new_[3377]_  = ~\new_[3658]_  | ~\new_[3648]_ ;
  assign \new_[3378]_  = ~\new_[3638]_  | ~\new_[3667]_ ;
  assign \new_[3379]_  = ~\new_[3643]_  | ~\new_[3660]_ ;
  assign \new_[3380]_  = ~\new_[3658]_  | ~\new_[3676]_ ;
  assign \new_[3381]_  = ~\new_[3665]_  | ~\new_[5269]_ ;
  assign \new_[3382]_  = ~\new_[3604]_  | ~\new_[3705]_ ;
  assign \new_[3383]_  = ~\new_[4380]_  | ~\new_[4785]_ ;
  assign \new_[3384]_  = ~\new_[3720]_  | ~\new_[3608]_ ;
  assign \new_[3385]_  = ~\new_[3621]_  | ~\new_[5180]_ ;
  assign \new_[3386]_  = ~\new_[5182]_  | ~\new_[3660]_ ;
  assign \new_[3387]_  = ~\new_[3520]_ ;
  assign \new_[3388]_  = ~\new_[5269]_  | ~\new_[3675]_ ;
  assign \new_[3389]_  = ~\new_[3622]_  | ~\new_[5273]_ ;
  assign \new_[3390]_  = ~\new_[3757]_  | ~\new_[3648]_ ;
  assign \new_[3391]_  = ~\new_[3638]_  | ~\new_[3738]_ ;
  assign \new_[3392]_  = ~\new_[3665]_  | ~\new_[3607]_ ;
  assign \new_[3393]_  = ~\new_[3701]_  | ~\new_[3673]_ ;
  assign \new_[3394]_  = ~\new_[5259]_  | ~\new_[5261]_ ;
  assign \new_[3395]_  = ~\new_[5257]_  | ~\new_[3757]_ ;
  assign \new_[3396]_  = ~\new_[3658]_  | ~\new_[3720]_ ;
  assign \new_[3397]_  = ~\new_[3701]_  | ~\new_[3693]_ ;
  assign \new_[3398]_  = ~\new_[3628]_  | ~\new_[3612]_ ;
  assign \new_[3399]_  = ~\new_[3499]_ ;
  assign \new_[3400]_  = \new_[3527]_ ;
  assign \new_[3401]_  = ~\new_[3583]_ ;
  assign \new_[3402]_  = ~\new_[3522]_ ;
  assign \new_[3403]_  = ~\new_[3570]_ ;
  assign \new_[3404]_  = ~\new_[3525]_ ;
  assign \new_[3405]_  = \new_[3537]_ ;
  assign \new_[3406]_  = ~\new_[3546]_ ;
  assign \new_[3407]_  = ~\new_[3563]_ ;
  assign \new_[3408]_  = ~\new_[3525]_ ;
  assign \new_[3409]_  = ~\new_[3510]_ ;
  assign \new_[3410]_  = ~\new_[3501]_ ;
  assign \new_[3411]_  = ~\new_[3504]_ ;
  assign \new_[3412]_  = \new_[3544]_ ;
  assign \new_[3413]_  = ~\new_[5269]_ ;
  assign \new_[3414]_  = ~\new_[3494]_ ;
  assign \new_[3415]_  = ~\new_[3596]_ ;
  assign \new_[3416]_  = ~\new_[3546]_ ;
  assign \new_[3417]_  = ~\new_[3600]_ ;
  assign \new_[3418]_  = ~\new_[3569]_ ;
  assign \new_[3419]_  = ~\new_[3547]_ ;
  assign \new_[3420]_  = ~\new_[3580]_ ;
  assign \new_[3421]_  = ~\new_[3549]_ ;
  assign \new_[3422]_  = ~\new_[3565]_ ;
  assign \new_[3423]_  = ~\new_[3565]_ ;
  assign \new_[3424]_  = ~\new_[3660]_ ;
  assign \new_[3425]_  = ~\new_[3519]_ ;
  assign \new_[3426]_  = ~\new_[3500]_ ;
  assign \new_[3427]_  = ~\new_[3674]_  | ~\new_[5261]_ ;
  assign \new_[3428]_  = ~\new_[3507]_ ;
  assign \new_[3429]_  = ~\new_[3507]_ ;
  assign \new_[3430]_  = ~\new_[3554]_ ;
  assign \new_[3431]_  = ~\new_[3498]_ ;
  assign \new_[3432]_  = ~\new_[3495]_ ;
  assign \new_[3433]_  = ~\new_[3557]_ ;
  assign \new_[3434]_  = ~\new_[3674]_  | ~\new_[3670]_ ;
  assign \new_[3435]_  = ~\new_[3597]_ ;
  assign \new_[3436]_  = ~\new_[3714]_  | ~\new_[3700]_ ;
  assign \new_[3437]_  = ~\new_[3502]_ ;
  assign \new_[3438]_  = ~\new_[3595]_ ;
  assign \new_[3439]_  = ~\new_[3591]_ ;
  assign \new_[3440]_  = ~\new_[3652]_  | ~\new_[3615]_ ;
  assign \new_[3441]_  = ~\new_[3707]_ ;
  assign \new_[3442]_  = ~\new_[3559]_ ;
  assign \new_[3443]_  = ~\new_[3538]_ ;
  assign \new_[3444]_  = ~\new_[3584]_ ;
  assign \new_[3445]_  = ~\new_[3576]_ ;
  assign \new_[3446]_  = ~\new_[3561]_ ;
  assign \new_[3447]_  = ~\new_[3562]_ ;
  assign \new_[3448]_  = ~\new_[3604]_ ;
  assign \new_[3449]_  = ~\new_[3670]_  | ~\new_[3603]_ ;
  assign \new_[3450]_  = ~\new_[3540]_ ;
  assign \new_[3451]_  = ~\new_[3679]_  | ~\new_[3987]_ ;
  assign \new_[3452]_  = ~\new_[3680]_  | ~\new_[3987]_ ;
  assign \new_[3453]_  = ~\new_[3565]_ ;
  assign \new_[3454]_  = ~\new_[3582]_ ;
  assign \new_[3455]_  = ~\new_[3701]_  | ~\new_[5273]_ ;
  assign \new_[3456]_  = ~\new_[3571]_ ;
  assign \new_[3457]_  = ~\new_[3562]_ ;
  assign \new_[3458]_  = ~\new_[3518]_ ;
  assign \new_[3459]_  = \new_[3764]_  ? \new_[3754]_  : \new_[2026]_ ;
  assign \new_[3460]_  = ~\new_[3561]_ ;
  assign \new_[3461]_  = (~\new_[3793]_  | ~\new_[3818]_ ) & (~\new_[3918]_  | ~\new_[2153]_ );
  assign \new_[3462]_  = \new_[2157]_  ? \new_[3883]_  : \new_[3761]_ ;
  assign \new_[3463]_  = ~\new_[3750]_  | (~\new_[3732]_  & ~\new_[3883]_ );
  assign \new_[3464]_  = \new_[3710]_  | \new_[3737]_ ;
  assign \new_[3465]_  = ~\new_[3570]_ ;
  assign \new_[3466]_  = ~\new_[3681]_  | ~\new_[3987]_ ;
  assign \new_[3467]_  = ~\new_[3670]_ ;
  assign \new_[3468]_  = ~\new_[3585]_ ;
  assign \new_[3469]_  = ~\new_[3569]_ ;
  assign \new_[3470]_  = ~\new_[3590]_ ;
  assign \new_[3471]_  = ~\new_[3590]_ ;
  assign \new_[3472]_  = ~\new_[3548]_ ;
  assign \new_[3473]_  = ~\new_[5269]_  | ~\new_[3758]_ ;
  assign \new_[3474]_  = ~\new_[3704]_  | ~\new_[3987]_ ;
  assign \new_[3475]_  = ~\new_[3682]_  | ~\new_[3987]_ ;
  assign \new_[3476]_  = ~\new_[3604]_  | ~\new_[3719]_ ;
  assign \new_[3477]_  = ~\new_[3592]_ ;
  assign \new_[3478]_  = ~\new_[3583]_ ;
  assign \new_[3479]_  = ~\new_[3514]_ ;
  assign \new_[3480]_  = ~\new_[3514]_ ;
  assign \new_[3481]_  = ~\new_[3502]_ ;
  assign \new_[3482]_  = ~\new_[3594]_ ;
  assign \new_[3483]_  = ~\new_[3531]_ ;
  assign \new_[3484]_  = ~\new_[3595]_ ;
  assign \new_[3485]_  = ~\new_[3516]_ ;
  assign \new_[3486]_  = ~\new_[3717]_ ;
  assign \new_[3487]_  = ~\new_[3599]_ ;
  assign \new_[3488]_  = ~\new_[3602]_ ;
  assign \new_[3489]_  = ~\new_[3754]_ ;
  assign \new_[3490]_  = \new_[3601]_ ;
  assign \new_[3491]_  = ~\new_[3628]_  | ~\new_[3700]_ ;
  assign \new_[3492]_  = ~\new_[3634]_ ;
  assign \new_[3493]_  = ~\new_[3656]_ ;
  assign \new_[3494]_  = ~\new_[3655]_ ;
  assign \new_[3495]_  = ~\new_[3624]_ ;
  assign \new_[3496]_  = ~\new_[3666]_ ;
  assign \new_[3497]_  = ~\new_[3643]_ ;
  assign \new_[3498]_  = \new_[3665]_ ;
  assign \new_[3499]_  = ~\new_[5262]_ ;
  assign \new_[3500]_  = ~\new_[3619]_ ;
  assign \new_[3501]_  = \new_[3652]_ ;
  assign \new_[3502]_  = ~\new_[3715]_ ;
  assign \new_[3503]_  = ~\new_[3721]_ ;
  assign \new_[3504]_  = ~\new_[3749]_  | ~\new_[3961]_ ;
  assign \new_[3505]_  = (~\new_[3813]_  | ~\new_[3952]_ ) & (~\new_[3884]_  | ~\new_[2274]_ );
  assign \new_[3506]_  = ~\new_[3790]_  | ~\new_[3728]_ ;
  assign \new_[3507]_  = ~\new_[3620]_ ;
  assign \new_[3508]_  = ~\new_[5179]_ ;
  assign \new_[3509]_  = ~\new_[5273]_ ;
  assign \new_[3510]_  = ~\new_[3630]_ ;
  assign \new_[3511]_  = \new_[5277]_ ;
  assign \new_[3512]_  = ~\new_[5255]_  | ~\new_[5279]_ ;
  assign \new_[3513]_  = ~\new_[3618]_ ;
  assign \new_[3514]_  = ~\new_[3657]_ ;
  assign \new_[3515]_  = \new_[5281]_ ;
  assign \new_[3516]_  = ~\new_[3714]_ ;
  assign \new_[3517]_  = ~\new_[3666]_ ;
  assign \new_[3518]_  = ~\new_[3683]_ ;
  assign \new_[3519]_  = ~\new_[3663]_ ;
  assign \new_[3520]_  = ~\new_[3664]_ ;
  assign \new_[3521]_  = ~\new_[3708]_ ;
  assign \new_[3522]_  = ~\new_[3716]_ ;
  assign \new_[3523]_  = ~\new_[3722]_  | ~\new_[3969]_ ;
  assign \new_[3524]_  = \new_[5279]_ ;
  assign \new_[3525]_  = ~\new_[3648]_ ;
  assign \new_[3526]_  = ~\new_[3736]_  | ~\new_[3727]_ ;
  assign \new_[3527]_  = \new_[3612]_ ;
  assign \new_[3528]_  = \new_[3607]_ ;
  assign \new_[3529]_  = ~\new_[3722]_  | ~\new_[3966]_ ;
  assign \new_[3530]_  = ~\new_[3633]_ ;
  assign \new_[3531]_  = ~\new_[3633]_ ;
  assign \new_[3532]_  = ~\new_[3708]_ ;
  assign \new_[3533]_  = ~\new_[3708]_ ;
  assign \new_[3534]_  = \new_[3638]_ ;
  assign \new_[3535]_  = ~\new_[3702]_ ;
  assign \new_[3536]_  = ~\new_[3733]_  | ~\new_[3760]_ ;
  assign \new_[3537]_  = \new_[3637]_ ;
  assign \new_[3538]_  = ~\new_[3635]_ ;
  assign \new_[3539]_  = ~\new_[4808]_ ;
  assign \new_[3540]_  = ~\new_[3623]_ ;
  assign \new_[3541]_  = ~\new_[5179]_ ;
  assign \new_[3542]_  = ~\new_[3651]_ ;
  assign \new_[3543]_  = ~\new_[3632]_ ;
  assign \new_[3544]_  = \new_[5258]_ ;
  assign \new_[3545]_  = \new_[3653]_ ;
  assign \new_[3546]_  = ~\new_[3654]_ ;
  assign \new_[3547]_  = ~\new_[3709]_ ;
  assign \new_[3548]_  = ~\new_[3705]_ ;
  assign \new_[3549]_  = ~\new_[3727]_ ;
  assign \new_[3550]_  = ~\new_[3661]_ ;
  assign \new_[3551]_  = ~\new_[3742]_  & (~\new_[3884]_  | ~\new_[2376]_ );
  assign \new_[3552]_  = ~\new_[3629]_ ;
  assign \new_[3553]_  = ~\new_[3625]_ ;
  assign \new_[3554]_  = ~\new_[3617]_ ;
  assign \new_[3555]_  = ~\new_[3616]_ ;
  assign \new_[3556]_  = ~\new_[3614]_ ;
  assign \new_[3557]_  = ~\new_[3603]_ ;
  assign \new_[3558]_  = \new_[3718]_ ;
  assign \new_[3559]_  = ~\new_[3700]_ ;
  assign \new_[3560]_  = \new_[3608]_ ;
  assign \new_[3561]_  = ~\new_[3678]_ ;
  assign \new_[3562]_  = ~\new_[3675]_ ;
  assign \new_[3563]_  = ~\new_[3644]_ ;
  assign \new_[3564]_  = \new_[3673]_ ;
  assign \new_[3565]_  = ~\new_[3626]_ ;
  assign \new_[3566]_  = \new_[3746]_  | \new_[3743]_ ;
  assign \new_[3567]_  = ~\new_[3674]_ ;
  assign \new_[3568]_  = (~\new_[3802]_  | ~\new_[3952]_ ) & (~\new_[3884]_  | ~\new_[2217]_ );
  assign \new_[3569]_  = ~\new_[3684]_ ;
  assign \new_[3570]_  = ~\new_[3636]_ ;
  assign \new_[3571]_  = ~\new_[3676]_ ;
  assign \new_[3572]_  = \new_[3741]_  & \new_[3987]_ ;
  assign \new_[3573]_  = \new_[3794]_  ? \new_[3918]_  : \new_[2023]_ ;
  assign \new_[3574]_  = ~\new_[3810]_  | (~\new_[3797]_  & ~\new_[3818]_ );
  assign \new_[3575]_  = ~\new_[3821]_  | (~\new_[3768]_  & ~\new_[3986]_ );
  assign \new_[3576]_  = \new_[3605]_ ;
  assign \new_[3577]_  = ~\new_[467]_  | ~\new_[3830]_ ;
  assign \new_[3578]_  = ~\new_[3759]_  | ~\desIn[9] ;
  assign \new_[3579]_  = ~\new_[5306]_  | ~\new_[3818]_  | ~\new_[2020]_ ;
  assign \new_[3580]_  = ~\new_[3693]_ ;
  assign \new_[3581]_  = ~\new_[3651]_ ;
  assign \new_[3582]_  = ~\new_[3694]_ ;
  assign \new_[3583]_  = ~\new_[3706]_ ;
  assign \new_[3584]_  = ~\new_[3611]_ ;
  assign \new_[3585]_  = ~\new_[3658]_ ;
  assign \new_[3586]_  = ~\new_[3757]_  | ~\new_[3758]_ ;
  assign \new_[3587]_  = \new_[3701]_ ;
  assign \new_[3588]_  = \new_[3628]_ ;
  assign \new_[3589]_  = ~\new_[3759]_  | ~\desIn[23] ;
  assign \new_[3590]_  = ~\new_[3671]_ ;
  assign \new_[3591]_  = ~\new_[3669]_ ;
  assign \new_[3592]_  = ~\new_[3711]_ ;
  assign \new_[3593]_  = ~\new_[3650]_ ;
  assign \new_[3594]_  = ~\new_[5260]_ ;
  assign \new_[3595]_  = ~\new_[3668]_ ;
  assign \new_[3596]_  = ~\new_[3719]_ ;
  assign \new_[3597]_  = ~\new_[3718]_ ;
  assign \new_[3598]_  = ~\new_[3645]_ ;
  assign \new_[3599]_  = \new_[3667]_ ;
  assign \new_[3600]_  = ~\new_[3720]_ ;
  assign \new_[3601]_  = ~\new_[3749]_  | ~\new_[4830]_ ;
  assign \new_[3602]_  = ~\new_[5100]_ ;
  assign \new_[3603]_  = ~\new_[3783]_  | ~\new_[3949]_ ;
  assign \new_[3604]_  = ~\new_[3792]_  | ~\new_[3981]_ ;
  assign \new_[3605]_  = ~\new_[4768]_  | ~\new_[3771]_ ;
  assign \new_[3606]_  = ~\new_[3823]_  | ~\new_[3791]_  | ~\new_[3839]_ ;
  assign \new_[3607]_  = ~\new_[5267]_  | ~\new_[3960]_ ;
  assign \new_[3608]_  = ~\new_[5295]_  | ~\new_[3782]_ ;
  assign \new_[3609]_  = ~\new_[5309]_  | ~\new_[3883]_  | ~\new_[496]_ ;
  assign \new_[3610]_  = \new_[3729]_ ;
  assign \new_[3611]_  = ~\new_[3769]_  | ~\new_[3855]_ ;
  assign \new_[3612]_  = ~\new_[3949]_  | ~\new_[3777]_ ;
  assign \new_[3613]_  = ~\new_[3774]_  | ~\new_[5296]_ ;
  assign \new_[3614]_  = ~\new_[3763]_  | ~\new_[5101]_ ;
  assign \new_[3615]_  = ~\new_[3805]_  | ~\new_[3948]_ ;
  assign \new_[3616]_  = ~\new_[3781]_  | ~\new_[3893]_ ;
  assign \new_[3617]_  = ~\new_[3804]_  | ~\new_[3906]_ ;
  assign \new_[3618]_  = ~\new_[3807]_  | ~\new_[3905]_ ;
  assign \new_[3619]_  = ~\new_[3765]_  | ~\new_[3949]_ ;
  assign \new_[3620]_  = ~\new_[4658]_  | ~\new_[4810]_ ;
  assign \new_[3621]_  = ~\new_[5295]_  | ~\new_[4866]_ ;
  assign \new_[3622]_  = ~\new_[3801]_  | ~\new_[5101]_ ;
  assign \new_[3623]_  = ~\new_[4788]_  | ~\new_[3784]_ ;
  assign \new_[3624]_  = ~\new_[3782]_  | ~\new_[3893]_ ;
  assign \new_[3625]_  = ~\new_[3785]_  | ~\new_[3947]_ ;
  assign \new_[3626]_  = ~\new_[3965]_  | ~\new_[3800]_ ;
  assign \new_[3627]_  = ~\new_[3713]_  | ~\desIn[45] ;
  assign \new_[3628]_  = ~\new_[3775]_  | ~\new_[3906]_ ;
  assign \new_[3629]_  = \new_[3736]_ ;
  assign \new_[3630]_  = ~\new_[3788]_  | ~\new_[4661]_ ;
  assign \new_[3631]_  = ~\new_[4809]_  | ~\new_[3949]_ ;
  assign \new_[3632]_  = ~\new_[3725]_ ;
  assign \new_[3633]_  = ~\new_[3730]_ ;
  assign \new_[3634]_  = ~\new_[3724]_ ;
  assign \new_[3635]_  = ~\new_[3786]_  | ~\new_[3917]_ ;
  assign \new_[3636]_  = ~\new_[3972]_  | ~\new_[3805]_ ;
  assign \new_[3637]_  = ~\new_[3855]_  | ~\new_[3807]_ ;
  assign \new_[3638]_  = ~\new_[3776]_  | ~\new_[3966]_ ;
  assign \new_[3639]_  = ~\new_[3796]_  | ~\new_[3885]_ ;
  assign \new_[3640]_  = ~\new_[3773]_  | ~\new_[3949]_ ;
  assign \new_[3641]_  = ~\new_[3809]_  | ~\new_[2163]_ ;
  assign \new_[3642]_  = ~\new_[3837]_  | ~\desIn[55] ;
  assign \new_[3643]_  = ~\new_[3767]_  | ~\new_[3905]_ ;
  assign \new_[3644]_  = ~\new_[3804]_  | ~\new_[4787]_ ;
  assign \new_[3645]_  = \new_[3760]_ ;
  assign \new_[3646]_  = \new_[3758]_ ;
  assign \new_[3647]_  = \new_[481]_  ? \new_[5306]_  : \new_[2024]_ ;
  assign \new_[3648]_  = ~\new_[3920]_  | ~\new_[3785]_ ;
  assign \new_[3649]_  = ~\new_[3972]_  | ~\new_[3765]_ ;
  assign \new_[3650]_  = ~\new_[3762]_  | ~\new_[3905]_ ;
  assign \new_[3651]_  = ~\new_[3733]_ ;
  assign \new_[3652]_  = ~\new_[3773]_  | ~\new_[3893]_ ;
  assign \new_[3653]_  = ~\new_[3770]_  | ~\new_[3980]_ ;
  assign \new_[3654]_  = ~\new_[3885]_  | ~\new_[3767]_ ;
  assign \new_[3655]_  = ~\new_[3772]_  | ~\new_[3966]_ ;
  assign \new_[3656]_  = ~\new_[4763]_  | ~\new_[3975]_ ;
  assign \new_[3657]_  = ~\new_[3788]_  | ~\new_[3948]_ ;
  assign \new_[3658]_  = ~\new_[3808]_  | ~\new_[3905]_ ;
  assign \new_[3659]_  = ~\new_[3906]_  | ~\new_[5106]_ ;
  assign \new_[3660]_  = ~\new_[3811]_  | ~\new_[3961]_ ;
  assign \new_[3661]_  = ~\new_[3723]_ ;
  assign \new_[3662]_  = ~\new_[3781]_  | ~\new_[5295]_ ;
  assign \new_[3663]_  = ~\new_[3780]_  | ~\new_[4787]_ ;
  assign \new_[3664]_  = ~\new_[5086]_  | ~\new_[4014]_ ;
  assign \new_[3665]_  = ~\new_[3799]_  | ~\new_[3855]_ ;
  assign \new_[3666]_  = ~\new_[3729]_ ;
  assign \new_[3667]_  = ~\new_[3772]_  | ~\new_[3947]_ ;
  assign \new_[3668]_  = ~\new_[3770]_  | ~\new_[3961]_ ;
  assign \new_[3669]_  = ~\new_[5256]_ ;
  assign \new_[3670]_  = ~\new_[3778]_  | ~\new_[4014]_ ;
  assign \new_[3671]_  = ~\new_[3774]_  | ~\new_[4718]_ ;
  assign \new_[3672]_  = \new_[3834]_  ? \new_[3918]_  : \new_[2031]_ ;
  assign \new_[3673]_  = ~\new_[3780]_  | ~\new_[3957]_ ;
  assign \new_[3674]_  = ~\new_[3789]_  | ~\new_[5296]_ ;
  assign \new_[3675]_  = ~\new_[3762]_  | ~\new_[3957]_ ;
  assign \new_[3676]_  = ~\new_[3885]_  | ~\new_[3763]_ ;
  assign \new_[3677]_  = ~\new_[3735]_ ;
  assign \new_[3678]_  = ~\new_[3808]_  | ~\new_[3855]_ ;
  assign \new_[3679]_  = (~\new_[3827]_  & ~\new_[3951]_ ) | (~\new_[3952]_  & ~\new_[4320]_ );
  assign \new_[3680]_  = (~\new_[3815]_  & ~\new_[3951]_ ) | (~\new_[3952]_  & ~\new_[4355]_ );
  assign \new_[3681]_  = (~\new_[3828]_  & ~\new_[3951]_ ) | (~\new_[3952]_  & ~\new_[4336]_ );
  assign \new_[3682]_  = (~\new_[3826]_  & ~\new_[3951]_ ) | (~\new_[3952]_  & ~\new_[4376]_ );
  assign \new_[3683]_  = ~\new_[3778]_  | ~\new_[3917]_ ;
  assign \new_[3684]_  = ~\new_[3771]_  | ~\new_[3966]_ ;
  assign \new_[3685]_  = (~\new_[4319]_  & ~\new_[3879]_ ) | (~\new_[3830]_  & ~\new_[4343]_ );
  assign \new_[3686]_  = ~\new_[2027]_  | ~\new_[3879]_ ;
  assign \new_[3687]_  = ~\new_[5300]_  | ~\new_[3883]_  | ~\new_[2022]_ ;
  assign \new_[3688]_  = ~\new_[5300]_  | ~\new_[3883]_  | ~\new_[2021]_ ;
  assign \new_[3689]_  = ~\new_[5299]_  | ~\new_[3883]_  | ~\new_[443]_ ;
  assign \new_[3690]_  = \new_[439]_  ? \new_[5300]_  : \new_[2163]_ ;
  assign \new_[3691]_  = \new_[451]_  ? \new_[5310]_  : \new_[2247]_ ;
  assign \new_[3692]_  = ~\new_[3713]_  | ~\desIn[61] ;
  assign \new_[3693]_  = ~\new_[5266]_  | ~\new_[3906]_ ;
  assign \new_[3694]_  = ~\new_[3801]_  | ~\new_[4810]_ ;
  assign \new_[3695]_  = \new_[437]_  ? \new_[5300]_  : \new_[2025]_ ;
  assign \new_[3696]_  = \new_[441]_  ? \new_[5306]_  : \new_[2018]_ ;
  assign \new_[3697]_  = ~\new_[3918]_  | ~\new_[2020]_ ;
  assign \new_[3698]_  = ~\new_[3837]_  | ~\desIn[13] ;
  assign \new_[3699]_  = ~\new_[3837]_  | ~\desIn[11] ;
  assign \new_[3700]_  = ~\new_[5086]_  | ~\new_[3965]_ ;
  assign \new_[3701]_  = ~\new_[3799]_  | ~\new_[4768]_ ;
  assign \new_[3702]_  = ~\new_[3753]_ ;
  assign \new_[3703]_  = \new_[3738]_ ;
  assign \new_[3704]_  = ~\new_[3829]_  | (~\new_[3816]_  & ~\new_[3951]_ );
  assign \new_[3705]_  = ~\new_[3779]_  | ~\new_[4718]_ ;
  assign \new_[3706]_  = ~\new_[3798]_  | ~\new_[3905]_ ;
  assign \new_[3707]_  = ~\new_[3786]_  | ~\new_[3961]_ ;
  assign \new_[3708]_  = ~\new_[3731]_ ;
  assign \new_[3709]_  = ~\new_[3779]_  | ~\new_[3917]_ ;
  assign \new_[3710]_  = \new_[2154]_  & \new_[3879]_ ;
  assign \new_[3711]_  = ~\new_[3734]_ ;
  assign \new_[3712]_  = ~\new_[3754]_ ;
  assign \new_[3713]_  = ~\new_[3739]_ ;
  assign \new_[3714]_  = ~\new_[3789]_  | ~\new_[4810]_ ;
  assign \new_[3715]_  = ~\new_[3811]_  | ~\new_[3917]_ ;
  assign \new_[3716]_  = ~\new_[3796]_  | ~\new_[3965]_ ;
  assign \new_[3717]_  = ~\new_[3784]_  | ~\new_[3949]_ ;
  assign \new_[3718]_  = ~\new_[3787]_  | ~\new_[3920]_ ;
  assign \new_[3719]_  = ~\new_[4786]_  | ~\new_[3972]_ ;
  assign \new_[3720]_  = ~\new_[3798]_  | ~\new_[4810]_ ;
  assign \new_[3721]_  = ~\new_[3757]_ ;
  assign \new_[3722]_  = ~\new_[4134]_  | ~\new_[3916]_  | ~\new_[3946]_  | ~\new_[4067]_ ;
  assign \new_[3723]_  = ~\new_[3819]_  | ~\new_[4810]_ ;
  assign \new_[3724]_  = ~\new_[3822]_  | ~\new_[5296]_ ;
  assign \new_[3725]_  = ~\new_[3822]_  | ~\new_[3975]_ ;
  assign \new_[3726]_  = ~\new_[3824]_  | ~\new_[3906]_ ;
  assign \new_[3727]_  = ~\new_[3832]_  | ~\new_[3975]_ ;
  assign \new_[3728]_  = ~\new_[504]_  | ~\new_[3830]_ ;
  assign \new_[3729]_  = ~\new_[3820]_  | ~\new_[5296]_ ;
  assign \new_[3730]_  = ~\new_[3820]_  | ~\new_[4014]_ ;
  assign \new_[3731]_  = ~\new_[3836]_  | ~\new_[4051]_ ;
  assign \new_[3732]_  = ~\new_[3739]_  | ~\new_[2247]_ ;
  assign \new_[3733]_  = ~\new_[4014]_  | ~\new_[3825]_ ;
  assign \new_[3734]_  = ~\new_[3824]_  | ~\new_[5296]_ ;
  assign \new_[3735]_  = ~\new_[3832]_  | ~\new_[3947]_ ;
  assign \new_[3736]_  = ~\new_[3838]_  | ~\new_[3965]_ ;
  assign \new_[3737]_  = \new_[449]_  & \new_[3830]_ ;
  assign \new_[3738]_  = ~\new_[3835]_  | ~\new_[5296]_ ;
  assign \new_[3739]_  = ~\new_[3837]_ ;
  assign \new_[3740]_  = ~\new_[3833]_  | ~\new_[3817]_ ;
  assign \new_[3741]_  = \new_[2194]_  ? \new_[3883]_  : \new_[3888]_ ;
  assign \new_[3742]_  = ~\new_[3884]_  & (~\new_[3921]_  | ~\new_[3880]_ );
  assign \new_[3743]_  = \new_[2156]_  ? \new_[3853]_  : \new_[3909]_ ;
  assign \new_[3744]_  = ~\new_[5299]_  | ~\new_[3952]_  | ~\new_[493]_ ;
  assign \new_[3745]_  = ~\new_[3837]_  | ~\desIn[35] ;
  assign \new_[3746]_  = ~\new_[3814]_ ;
  assign \new_[3747]_  = \new_[471]_  ? \new_[5303]_  : \new_[2346]_ ;
  assign \new_[3748]_  = ~\new_[3837]_  | ~\desIn[37] ;
  assign \new_[3749]_  = ~\new_[4136]_  | ~\new_[4045]_  | ~\new_[3925]_  | ~\new_[3990]_ ;
  assign \new_[3750]_  = ~\new_[3837]_  | ~\desIn[15] ;
  assign \new_[3751]_  = ~\new_[3914]_  | ~\desIn[39] ;
  assign \new_[3752]_  = ~\new_[3914]_  | ~\desIn[3] ;
  assign \new_[3753]_  = ~\new_[5295]_  | ~\new_[3819]_ ;
  assign \new_[3754]_  = ~\new_[3883]_ ;
  assign \new_[3755]_  = ~\new_[3914]_  | ~\desIn[1] ;
  assign \new_[3756]_  = ~\new_[3837]_  | ~\desIn[59] ;
  assign \new_[3757]_  = ~\new_[3836]_  | ~\new_[3960]_ ;
  assign \new_[3758]_  = ~\new_[3835]_  | ~\new_[3957]_ ;
  assign \new_[3759]_  = ~\new_[3809]_ ;
  assign \new_[3760]_  = ~\new_[4715]_  | ~\new_[5295]_ ;
  assign \new_[3761]_  = \new_[482]_  ? \new_[5310]_  : \new_[2157]_ ;
  assign \new_[3762]_  = ~\new_[3841]_  | ~\new_[3874]_ ;
  assign \new_[3763]_  = ~\new_[3931]_  | ~\new_[3871]_ ;
  assign \new_[3764]_  = \new_[479]_  ? \new_[5303]_  : \new_[2026]_ ;
  assign \new_[3765]_  = ~\new_[3845]_  | ~\new_[3945]_ ;
  assign \new_[3766]_  = \new_[3894]_  ? \new_[3951]_  : \new_[2417]_ ;
  assign \new_[3767]_  = ~\new_[3882]_  | ~\new_[3860]_ ;
  assign \new_[3768]_  = ~\new_[3809]_  | ~\new_[2346]_ ;
  assign \new_[3769]_  = ~\new_[3868]_  | ~\new_[3935]_ ;
  assign \new_[3770]_  = ~\new_[3857]_  | ~\new_[3910]_ ;
  assign \new_[3771]_  = ~\new_[4119]_  | ~\new_[3967]_  | ~\new_[3974]_  | ~\new_[3959]_ ;
  assign \new_[3772]_  = ~\new_[3908]_  | ~\new_[3858]_ ;
  assign \new_[3773]_  = ~\new_[3911]_  | ~\new_[3852]_ ;
  assign \new_[3774]_  = ~\new_[3863]_  | ~\new_[3901]_ ;
  assign \new_[3775]_  = ~\new_[3872]_  | ~\new_[3913]_ ;
  assign \new_[3776]_  = ~\new_[3861]_  | ~\new_[3956]_ ;
  assign \new_[3777]_  = ~\new_[3859]_  | ~\new_[3919]_ ;
  assign \new_[3778]_  = ~\new_[3940]_  | ~\new_[3864]_ ;
  assign \new_[3779]_  = ~\new_[3955]_  | ~\new_[3854]_ ;
  assign \new_[3780]_  = ~\new_[3979]_  | ~\new_[3842]_  | ~\new_[3962]_ ;
  assign \new_[3781]_  = ~\new_[3928]_  | ~\new_[5221]_ ;
  assign \new_[3782]_  = ~\new_[3846]_  | ~\new_[3896]_ ;
  assign \new_[3783]_  = ~\new_[3944]_  | ~\new_[3840]_ ;
  assign \new_[3784]_  = ~\new_[3847]_  | ~\new_[3953]_ ;
  assign \new_[3785]_  = ~\new_[3907]_  | ~\new_[3856]_ ;
  assign \new_[3786]_  = ~\new_[3886]_  | ~\new_[3922]_ ;
  assign \new_[3787]_  = ~\new_[3877]_  | ~\new_[3881]_ ;
  assign \new_[3788]_  = ~\new_[3851]_  | ~\new_[3937]_ ;
  assign \new_[3789]_  = ~\new_[3870]_  | ~\new_[3939]_ ;
  assign \new_[3790]_  = ~\new_[2019]_  | ~\new_[3879]_ ;
  assign \new_[3791]_  = ~\new_[5310]_  | ~\new_[3853]_  | ~\new_[2207]_ ;
  assign \new_[3792]_  = ~\new_[3850]_  | ~\new_[3933]_ ;
  assign \new_[3793]_  = \new_[464]_  ? \new_[5310]_  : \new_[2153]_ ;
  assign \new_[3794]_  = ~\new_[3950]_  | ~\new_[3878]_ ;
  assign \new_[3795]_  = \new_[3837]_  & \desIn[27] ;
  assign \new_[3796]_  = ~\new_[3867]_  | ~\new_[3915]_ ;
  assign \new_[3797]_  = ~\new_[3987]_  | ~\new_[2162]_ ;
  assign \new_[3798]_  = ~\new_[3941]_  | ~\new_[3862]_ ;
  assign \new_[3799]_  = ~\new_[3843]_  | ~\new_[3890]_ ;
  assign \new_[3800]_  = ~\new_[3873]_  | ~\new_[3899]_ ;
  assign \new_[3801]_  = ~\new_[3866]_  | ~\new_[3904]_ ;
  assign \new_[3802]_  = \new_[478]_  ? \new_[5303]_  : \new_[2217]_ ;
  assign \new_[3803]_  = ~\new_[3884]_  | ~\new_[2021]_ ;
  assign \new_[3804]_  = ~\new_[3943]_  | ~\new_[3849]_ ;
  assign \new_[3805]_  = ~\new_[3895]_  | ~\new_[3844]_ ;
  assign \new_[3806]_  = ~\new_[3884]_  | ~\new_[2022]_ ;
  assign \new_[3807]_  = ~\new_[3942]_  | ~\new_[3875]_ ;
  assign \new_[3808]_  = ~\new_[3869]_  | ~\new_[3936]_ ;
  assign \new_[3809]_  = ~\new_[3914]_ ;
  assign \new_[3810]_  = ~\new_[3837]_  | ~\desIn[7] ;
  assign \new_[3811]_  = ~\new_[3865]_  | ~\new_[3900]_ ;
  assign \new_[3812]_  = \new_[495]_  ? \new_[5310]_  : \new_[2162]_ ;
  assign \new_[3813]_  = \new_[486]_  ? \new_[5306]_  : \new_[2274]_ ;
  assign \new_[3814]_  = ~\new_[2156]_  | ~\new_[3883]_  | ~\new_[5300]_ ;
  assign \new_[3815]_  = \new_[4324]_  ? \new_[5310]_  : \new_[4355]_ ;
  assign \new_[3816]_  = \new_[4303]_  ? \new_[5306]_  : \new_[4373]_ ;
  assign \new_[3817]_  = ~\new_[3889]_  | ~\new_[3952]_ ;
  assign \new_[3818]_  = ~\new_[3918]_ ;
  assign \new_[3819]_  = ~\new_[3927]_  | ~\new_[3897]_ ;
  assign \new_[3820]_  = ~\new_[3903]_  | ~\new_[3929]_ ;
  assign \new_[3821]_  = ~\new_[3914]_  | ~\desIn[29] ;
  assign \new_[3822]_  = ~\new_[3938]_  | ~\new_[3924]_ ;
  assign \new_[3823]_  = ~\new_[5302]_  | ~\new_[3952]_  | ~\new_[445]_ ;
  assign \new_[3824]_  = ~\new_[3934]_  | ~\new_[3988]_ ;
  assign \new_[3825]_  = ~\new_[3887]_  | ~\new_[3902]_ ;
  assign \new_[3826]_  = \new_[4304]_  ? \new_[5303]_  : \new_[4376]_ ;
  assign \new_[3827]_  = \new_[4333]_  ? \new_[5312]_  : \new_[4320]_ ;
  assign \new_[3828]_  = \new_[4371]_  ? \new_[5304]_  : \new_[4336]_ ;
  assign \new_[3829]_  = \new_[3952]_  | \new_[4373]_ ;
  assign \new_[3830]_  = ~\new_[3879]_ ;
  assign \new_[3831]_  = ~\new_[3951]_  & ~\new_[3914]_ ;
  assign \new_[3832]_  = ~\new_[3930]_  | ~\new_[3892]_ ;
  assign \new_[3833]_  = ~\new_[3951]_  | ~\new_[2412]_ ;
  assign \new_[3834]_  = \new_[491]_  ? \new_[5310]_  : \new_[2031]_ ;
  assign \new_[3835]_  = ~\new_[3926]_  | ~\new_[3973]_ ;
  assign \new_[3836]_  = ~\new_[3932]_  | ~\new_[3978]_ ;
  assign \new_[3837]_  = ~\new_[3987]_ ;
  assign \new_[3838]_  = ~\new_[3898]_  | ~\new_[3954]_ ;
  assign \new_[3839]_  = \new_[3986]_  | \new_[4299]_ ;
  assign \new_[3840]_  = ~\new_[4058]_  & ~\new_[3964]_ ;
  assign \new_[3841]_  = ~\new_[3982]_  & (~\new_[4094]_  | ~\key1[29] );
  assign \new_[3842]_  = ~\new_[4073]_  & (~\new_[4005]_  | ~\key2[8] );
  assign \new_[3843]_  = (~\new_[4034]_  | ~\key2[28] ) & (~\new_[4227]_  | ~\key3[28] );
  assign \new_[3844]_  = ~\new_[4157]_  & ~\new_[3989]_ ;
  assign \new_[3845]_  = (~\new_[4010]_  | ~\key2[3] ) & (~\new_[4172]_  | ~\key3[3] );
  assign \new_[3846]_  = ~\new_[4151]_  & (~\new_[4036]_  | ~\key2[35] );
  assign \new_[3847]_  = (~\new_[4001]_  | ~\key2[10] ) & (~\new_[4246]_  | ~\key3[10] );
  assign \new_[3848]_  = (~\new_[4039]_  | ~\key2[46] ) & (~\new_[4172]_  | ~\key3[46] );
  assign \new_[3849]_  = (~\new_[3995]_  | ~\key2[49] ) & (~\new_[4172]_  | ~\key3[49] );
  assign \new_[3850]_  = ~\new_[3976]_  & (~\new_[4227]_  | ~\key3[39] );
  assign \new_[3851]_  = ~\new_[4147]_  & (~\new_[4007]_  | ~\key2[15] );
  assign \new_[3852]_  = ~\new_[4114]_  & (~\new_[4031]_  | ~\key2[18] );
  assign \new_[3853]_  = ~\new_[3918]_ ;
  assign \new_[3854]_  = ~\new_[3977]_  & (~\new_[4260]_  | ~\key3[33] );
  assign \new_[3855]_  = ~\new_[4864]_ ;
  assign \new_[3856]_  = (~\new_[4006]_  | ~\key2[31] ) & (~\new_[4260]_  | ~\key3[31] );
  assign \new_[3857]_  = ~\new_[4061]_  & (~\new_[4019]_  | ~\key2[34] );
  assign \new_[3858]_  = ~\new_[4092]_  & (~\new_[3997]_  | ~\key2[16] );
  assign \new_[3859]_  = ~\new_[4146]_  & (~\new_[4025]_  | ~\key2[2] );
  assign \new_[3860]_  = ~\new_[4132]_  & (~\new_[3998]_  | ~\key2[41] );
  assign \new_[3861]_  = ~\new_[4107]_  & (~\new_[3996]_  | ~\key2[37] );
  assign \new_[3862]_  = ~\new_[4129]_  & (~\new_[4026]_  | ~\key2[30] );
  assign \new_[3863]_  = ~\new_[4060]_  & (~\new_[4038]_  | ~\key2[25] );
  assign \new_[3864]_  = ~\new_[4091]_  & (~\new_[3992]_  | ~\key2[45] );
  assign \new_[3865]_  = (~\new_[4037]_  | ~\key2[17] ) & (~\new_[4217]_  | ~\key3[17] );
  assign \new_[3866]_  = (~\new_[4008]_  | ~\key2[0] ) & (~\new_[4260]_  | ~\key3[0] );
  assign \new_[3867]_  = (~\new_[4040]_  | ~\key2[55] ) & (~\new_[4227]_  | ~\key3[55] );
  assign \new_[3868]_  = (~\new_[4009]_  | ~\key2[23] ) & (~\new_[4217]_  | ~\key3[23] );
  assign \new_[3869]_  = (~\new_[3995]_  | ~\key2[22] ) & (~\new_[4246]_  | ~\key3[22] );
  assign \new_[3870]_  = (~\new_[4040]_  | ~\key2[51] ) & (~\new_[4227]_  | ~\key3[51] );
  assign \new_[3871]_  = (~\new_[4037]_  | ~\key2[43] ) & (~\new_[4260]_  | ~\key3[43] );
  assign \new_[3872]_  = (~\new_[4008]_  | ~\key2[50] ) & (~\new_[4172]_  | ~\key3[50] );
  assign \new_[3873]_  = (~\new_[4039]_  | ~\key2[42] ) & (~\new_[4217]_  | ~\key3[42] );
  assign \new_[3874]_  = (~\new_[4001]_  | ~\key2[29] ) & (~\new_[4172]_  | ~\key3[29] );
  assign \new_[3875]_  = (~\new_[4009]_  | ~\key2[12] ) & (~\new_[4246]_  | ~\key3[12] );
  assign \new_[3876]_  = ~\new_[3983]_  & (~\new_[4095]_  | ~\key1[32] );
  assign \new_[3877]_  = ~\new_[3963]_  & (~\new_[4097]_  | ~\key1[24] );
  assign \new_[3878]_  = \new_[4339]_  | \new_[5310]_ ;
  assign \new_[3879]_  = ~\new_[3986]_  | ~\new_[5311]_ ;
  assign \new_[3880]_  = \new_[4338]_  | \new_[5301]_ ;
  assign \new_[3881]_  = ~\new_[3970]_  & (~\new_[4260]_  | ~\key3[24] );
  assign \new_[3882]_  = ~\new_[3984]_  & (~\new_[4057]_  | ~\key1[41] );
  assign \new_[3883]_  = ~\new_[3918]_ ;
  assign \new_[3884]_  = ~\new_[3952]_ ;
  assign \new_[3885]_  = ~\new_[3948]_ ;
  assign \new_[3886]_  = (~\new_[4006]_  | ~\key2[54] ) & (~\new_[4227]_  | ~\key3[54] );
  assign \new_[3887]_  = (~\new_[4070]_  | ~\key2[14] ) & (~\new_[4217]_  | ~\key3[14] );
  assign \new_[3888]_  = \new_[468]_  ? \new_[5310]_  : \new_[2194]_ ;
  assign \new_[3889]_  = \new_[447]_  ? \new_[5310]_  : \new_[2412]_ ;
  assign \new_[3890]_  = (~\new_[4095]_  | ~\key1[28] ) & (~\key3[28]  | ~\new_[4144]_ );
  assign \new_[3891]_  = ~\new_[4032]_  & (~\new_[4056]_  | ~\key1[46] );
  assign \new_[3892]_  = (~\new_[4087]_  | ~\key2[27] ) & (~\new_[4227]_  | ~\key3[27] );
  assign \new_[3893]_  = ~\new_[4829]_ ;
  assign \new_[3894]_  = \new_[484]_  ? \new_[5305]_  : \new_[2417]_ ;
  assign \new_[3895]_  = ~\new_[3993]_  & (~\new_[4055]_  | ~\key1[40] );
  assign \new_[3896]_  = (~\new_[4081]_  | ~\key1[35] ) & (~\key3[35]  | ~\new_[4144]_ );
  assign \new_[3897]_  = (~\new_[4053]_  | ~\key2[21] ) & (~\new_[4172]_  | ~\key3[21] );
  assign \new_[3898]_  = ~\new_[4003]_  & (~\new_[4096]_  | ~\key1[20] );
  assign \new_[3899]_  = (~\new_[4071]_  | ~\key1[42] ) & (~\key3[42]  | ~\new_[4165]_ );
  assign \new_[3900]_  = ~\new_[4000]_  & (~\new_[4963]_  | ~\key1[17] );
  assign \new_[3901]_  = (~\new_[4075]_  | ~\key1[25] ) & (~\key3[25]  | ~\new_[4120]_ );
  assign \new_[3902]_  = (~\new_[4078]_  | ~\key1[14] ) & (~\key3[14]  | ~\new_[4182]_ );
  assign \new_[3903]_  = (~\new_[4053]_  | ~\key2[11] ) & (~\new_[4246]_  | ~\key3[11] );
  assign \new_[3904]_  = (~\new_[4078]_  | ~\key1[0] ) & (~\key3[0]  | ~\new_[4144]_ );
  assign \new_[3905]_  = \new_[4813]_ ;
  assign \new_[3906]_  = ~\new_[4829]_ ;
  assign \new_[3907]_  = (~\new_[4089]_  | ~\key1[31] ) & (~\new_[4088]_  | ~\key3[31] );
  assign \new_[3908]_  = (~\new_[4076]_  | ~\key1[16] ) & (~\key3[16]  | ~\new_[4165]_ );
  assign \new_[3909]_  = \new_[469]_  & \new_[5311]_ ;
  assign \new_[3910]_  = ~\new_[4041]_  & (~\new_[4054]_  | ~\key1[34] );
  assign \new_[3911]_  = (~\new_[4077]_  | ~\key1[18] ) & (~\key3[18]  | ~\new_[4144]_ );
  assign \new_[3912]_  = (~\new_[4077]_  | ~\key1[9] ) & (~\key3[9]  | ~\new_[4120]_ );
  assign \new_[3913]_  = ~\new_[3999]_  & (~\new_[4963]_  | ~\key1[50] );
  assign \new_[3914]_  = ~\new_[3987]_ ;
  assign \new_[3915]_  = ~\new_[4033]_  & (~\new_[4094]_  | ~\key1[55] );
  assign \new_[3916]_  = ~\new_[4052]_  | ~\key2[36] ;
  assign \new_[3917]_  = ~\new_[3968]_ ;
  assign \new_[3918]_  = ~\new_[3986]_ ;
  assign \new_[3919]_  = ~\new_[4013]_  & (~\new_[4081]_  | ~\key1[2] );
  assign \new_[3920]_  = ~\new_[3980]_ ;
  assign \new_[3921]_  = \new_[4356]_  | \new_[5313]_ ;
  assign \new_[3922]_  = ~\new_[4018]_  & (~\new_[4089]_  | ~\key1[54] );
  assign \new_[3923]_  = (~\new_[4070]_  | ~\key2[32] ) & (~\new_[4260]_  | ~\key3[32] );
  assign \new_[3924]_  = (~\new_[4059]_  | ~\key2[53] ) & (~\new_[4246]_  | ~\key3[53] );
  assign \new_[3925]_  = ~\new_[4049]_  | ~\key2[47] ;
  assign \new_[3926]_  = (~\new_[4093]_  | ~\key1[44] ) & (~\key3[44]  | ~\new_[4165]_ );
  assign \new_[3927]_  = ~\new_[3991]_  & (~\new_[4062]_  | ~\key1[21] );
  assign \new_[3928]_  = (~\new_[4063]_  | ~\key1[4] ) & (~\key3[4]  | ~\new_[4144]_ );
  assign \new_[3929]_  = ~\new_[4012]_  & (~\new_[4062]_  | ~\key1[11] );
  assign \new_[3930]_  = ~\new_[4046]_  & (~\new_[4096]_  | ~\key1[27] );
  assign \new_[3931]_  = ~\new_[4042]_  & (~\new_[4963]_  | ~\key1[43] );
  assign \new_[3932]_  = (~\new_[4064]_  | ~\key1[38] ) & (~\key3[38]  | ~\new_[4194]_ );
  assign \new_[3933]_  = ~\new_[4043]_  & (~\new_[4075]_  | ~\key1[39] );
  assign \new_[3934]_  = (~\new_[4100]_  | ~\key1[19] ) & (~\key3[19]  | ~\new_[4182]_ );
  assign \new_[3935]_  = ~\new_[4024]_  & (~\new_[4056]_  | ~\key1[23] );
  assign \new_[3936]_  = (~\new_[4086]_  | ~\key1[22] ) & (~\key3[22]  | ~\new_[4120]_ );
  assign \new_[3937]_  = (~\new_[4063]_  | ~\key1[15] ) & (~\key3[15]  | ~\new_[4165]_ );
  assign \new_[3938]_  = (~\new_[4082]_  | ~\key1[53] ) & (~\key3[53]  | ~\new_[4182]_ );
  assign \new_[3939]_  = ~\new_[4020]_  & (~\new_[4100]_  | ~\key1[51] );
  assign \new_[3940]_  = ~\new_[4015]_  & (~\new_[4057]_  | ~\key1[45] );
  assign \new_[3941]_  = (~\new_[4055]_  | ~\key1[30] ) & (~\new_[4083]_  | ~\key3[30] );
  assign \new_[3942]_  = (~\new_[4064]_  | ~\key1[12] ) & (~\key3[12]  | ~\new_[4144]_ );
  assign \new_[3943]_  = ~\new_[4016]_  & (~\new_[4086]_  | ~\key1[49] );
  assign \new_[3944]_  = ~\new_[4022]_  & (~\new_[4076]_  | ~\key1[52] );
  assign \new_[3945]_  = (~\new_[4084]_  | ~\key1[3] ) & (~\key3[3]  | ~\new_[4156]_ );
  assign \new_[3946]_  = ~\new_[4044]_  & ~\new_[4111]_ ;
  assign \new_[3947]_  = ~\new_[3961]_ ;
  assign \new_[3948]_  = ~\new_[4769]_ ;
  assign \new_[3949]_  = ~\new_[5102]_ ;
  assign \new_[3950]_  = \new_[4372]_  | \new_[5313]_ ;
  assign \new_[3951]_  = \new_[3971]_ ;
  assign \new_[3952]_  = ~\new_[3971]_ ;
  assign \new_[3953]_  = ~\new_[4050]_  & (~\new_[4072]_  | ~\key1[10] );
  assign \new_[3954]_  = (~\new_[4087]_  | ~\key2[20] ) & (~\new_[4217]_  | ~\key3[20] );
  assign \new_[3955]_  = ~\new_[4011]_  & (~\new_[4090]_  | ~\key1[33] );
  assign \new_[3956]_  = ~\new_[4027]_  & (~\new_[4097]_  | ~\key1[37] );
  assign \new_[3957]_  = ~\new_[4830]_ ;
  assign \new_[3958]_  = ~\new_[4023]_ ;
  assign \new_[3959]_  = ~\new_[4066]_  | ~\key1[48] ;
  assign \new_[3960]_  = ~\new_[4051]_ ;
  assign \new_[3961]_  = ~\new_[4030]_ ;
  assign \new_[3962]_  = ~\key3[8]  | ~\new_[4088]_ ;
  assign \new_[3963]_  = ~\new_[4295]_  & ~\new_[4079]_ ;
  assign \new_[3964]_  = ~\new_[4312]_  & (~\new_[5227]_  | ~\new_[5223]_ );
  assign \new_[3965]_  = ~\new_[4051]_ ;
  assign \new_[3966]_  = ~\new_[4048]_ ;
  assign \new_[3967]_  = ~\new_[4099]_  | ~\key2[48] ;
  assign \new_[3968]_  = ~\new_[4048]_ ;
  assign \new_[3969]_  = ~\new_[4051]_ ;
  assign \new_[3970]_  = ~\new_[4322]_  & (~\new_[4234]_  | ~\new_[4155]_ );
  assign \new_[3971]_  = \new_[4002]_ ;
  assign \new_[3972]_  = \new_[4051]_ ;
  assign \new_[3973]_  = ~\new_[4068]_  & (~\new_[4193]_  | ~\key2[44] );
  assign \new_[3974]_  = ~\key3[48]  | ~\new_[4088]_ ;
  assign \new_[3975]_  = ~\new_[4030]_ ;
  assign \new_[3976]_  = ~\new_[4323]_  & (~\new_[4110]_  | ~\new_[4236]_ );
  assign \new_[3977]_  = ~\new_[4301]_  & (~\new_[5223]_  | ~\new_[4234]_ );
  assign \new_[3978]_  = (~\new_[4141]_  | ~\key2[38] ) & (~\new_[4219]_  | ~\key3[38] );
  assign \new_[3979]_  = ~\new_[4090]_  | ~\key1[8] ;
  assign \new_[3980]_  = ~\new_[4051]_ ;
  assign \new_[3981]_  = ~\new_[4051]_ ;
  assign \new_[3982]_  = ~\new_[4306]_  & ~\new_[4079]_ ;
  assign \new_[3983]_  = ~\new_[4354]_  & ~\new_[4079]_ ;
  assign \new_[3984]_  = ~\new_[4317]_  & ~\new_[4079]_ ;
  assign \new_[3985]_  = ~\new_[4115]_ ;
  assign \new_[3986]_  = ~\new_[4002]_ ;
  assign \new_[3987]_  = ~\new_[4029]_ ;
  assign \new_[3988]_  = (~\new_[4141]_  | ~\key2[19] ) & (~\new_[4246]_  | ~\key3[19] );
  assign \new_[3989]_  = ~\new_[4292]_  & (~\new_[5227]_  | ~\new_[4912]_ );
  assign \new_[3990]_  = ~\new_[4093]_  | ~\key1[47] ;
  assign \new_[3991]_  = ~\new_[4148]_  & ~\new_[4332]_ ;
  assign \new_[3992]_  = ~\new_[4229]_  | ~\new_[4105]_ ;
  assign \new_[3993]_  = ~\new_[4345]_  & ~\new_[4128]_ ;
  assign \new_[3994]_  = ~\new_[4367]_  & ~\new_[4149]_ ;
  assign \new_[3995]_  = ~\new_[4229]_  | ~\new_[4110]_ ;
  assign \new_[3996]_  = ~\new_[4251]_  | ~\new_[4110]_ ;
  assign \new_[3997]_  = ~\new_[4913]_  | ~\new_[4105]_ ;
  assign \new_[3998]_  = ~\new_[4234]_  | ~\new_[4155]_ ;
  assign \new_[3999]_  = ~\new_[4348]_  & ~\new_[4154]_ ;
  assign \new_[4000]_  = ~\new_[4302]_  & ~\new_[4101]_ ;
  assign \new_[4001]_  = ~\new_[4110]_  | ~\new_[4236]_ ;
  assign \new_[4002]_  = ~\new_[4257]_  & ~\new_[4106]_ ;
  assign \new_[4003]_  = ~\new_[4326]_  & ~\new_[4128]_ ;
  assign \new_[4004]_  = ~\new_[4234]_  | ~\new_[5223]_ ;
  assign \new_[4005]_  = ~\new_[5227]_  | ~\new_[4912]_ ;
  assign \new_[4006]_  = ~\new_[4110]_  | ~\new_[4236]_ ;
  assign \new_[4007]_  = ~\new_[4229]_  | ~\new_[4110]_ ;
  assign \new_[4008]_  = ~\new_[4912]_  | ~\new_[4913]_ ;
  assign \new_[4009]_  = ~\new_[4112]_  | ~\new_[4225]_ ;
  assign \new_[4010]_  = ~\new_[4110]_  | ~\new_[4229]_ ;
  assign \new_[4011]_  = ~\new_[4308]_  & ~\new_[4153]_ ;
  assign \new_[4012]_  = ~\new_[4337]_  & ~\new_[4128]_ ;
  assign \new_[4013]_  = ~\new_[4374]_  & ~\new_[4130]_ ;
  assign \new_[4014]_  = \new_[4789]_ ;
  assign \new_[4015]_  = ~\new_[4340]_  & ~\new_[4148]_ ;
  assign \new_[4016]_  = ~\new_[4291]_  & ~\new_[4154]_ ;
  assign \new_[4017]_  = ~\new_[4341]_  & ~\new_[4101]_ ;
  assign \new_[4018]_  = ~\new_[4309]_  & ~\new_[4117]_ ;
  assign \new_[4019]_  = ~\new_[4103]_  | ~\new_[4913]_ ;
  assign \new_[4020]_  = ~\new_[4369]_  & ~\new_[4148]_ ;
  assign \new_[4021]_  = ~\new_[4080]_ ;
  assign \new_[4022]_  = ~\new_[4342]_  & ~\new_[4148]_ ;
  assign \new_[4023]_  = \new_[4170]_ ;
  assign \new_[4024]_  = ~\new_[4300]_  & ~\new_[4101]_ ;
  assign \new_[4025]_  = ~\new_[5227]_  | ~\new_[5223]_ ;
  assign \new_[4026]_  = ~\new_[4234]_  | ~\new_[4155]_ ;
  assign \new_[4027]_  = ~\new_[4344]_  & ~\new_[4101]_ ;
  assign \new_[4028]_  = ~\new_[4365]_  & ~\new_[4128]_ ;
  assign \new_[4029]_  = ~\new_[4223]_  & ~\new_[4106]_ ;
  assign \new_[4030]_  = ~\new_[4789]_ ;
  assign \new_[4031]_  = ~\new_[4234]_  | ~\new_[4155]_ ;
  assign \new_[4032]_  = ~\new_[4293]_  & ~\new_[4154]_ ;
  assign \new_[4033]_  = ~\new_[4352]_  & ~\new_[4117]_ ;
  assign \new_[4034]_  = ~\new_[4110]_  | ~\new_[4229]_ ;
  assign \new_[4035]_  = ~\new_[4912]_  | ~\new_[5227]_ ;
  assign \new_[4036]_  = ~\new_[4234]_  | ~\new_[5223]_ ;
  assign \new_[4037]_  = ~\new_[4124]_  | ~\new_[4251]_ ;
  assign \new_[4038]_  = ~\new_[4912]_  | ~\new_[4913]_ ;
  assign \new_[4039]_  = ~\new_[4124]_  | ~\new_[4225]_ ;
  assign \new_[4040]_  = ~\new_[4110]_  | ~\new_[4236]_ ;
  assign \new_[4041]_  = ~\new_[4298]_  & ~\new_[4123]_ ;
  assign \new_[4042]_  = ~\new_[4347]_  & ~\new_[4154]_ ;
  assign \new_[4043]_  = ~\new_[4318]_  & ~\new_[4138]_ ;
  assign \new_[4044]_  = ~\new_[4325]_  & ~\new_[4137]_ ;
  assign \new_[4045]_  = ~\key3[47]  | ~\new_[4156]_ ;
  assign \new_[4046]_  = ~\new_[4327]_  & ~\new_[4153]_ ;
  assign \new_[4047]_  = ~\new_[4085]_ ;
  assign \new_[4048]_  = ~\new_[4789]_ ;
  assign \new_[4049]_  = ~\new_[4225]_  | ~\new_[4112]_ ;
  assign \new_[4050]_  = ~\new_[4315]_  & ~\new_[4117]_ ;
  assign \new_[4051]_  = \new_[4663]_ ;
  assign \new_[4052]_  = ~\new_[4124]_  | ~\new_[4225]_ ;
  assign \new_[4053]_  = ~\new_[4251]_  | ~\new_[4187]_ ;
  assign \new_[4054]_  = ~\new_[4230]_  | ~\new_[4159]_ ;
  assign \new_[4055]_  = ~\new_[4243]_  | ~\new_[4202]_ ;
  assign \new_[4056]_  = ~\new_[4205]_  | ~\new_[4243]_ ;
  assign \new_[4057]_  = ~\new_[4230]_  | ~\new_[4159]_ ;
  assign \new_[4058]_  = ~\new_[4171]_  & ~\new_[4342]_ ;
  assign \new_[4059]_  = ~\new_[4187]_  | ~\new_[4251]_ ;
  assign \new_[4060]_  = ~\new_[4171]_  & ~\new_[4328]_ ;
  assign \new_[4061]_  = ~\new_[4171]_  & ~\new_[4298]_ ;
  assign \new_[4062]_  = ~\new_[4243]_  | ~\new_[4202]_ ;
  assign \new_[4063]_  = ~\new_[4243]_  | ~\new_[4205]_ ;
  assign \new_[4064]_  = ~\new_[4213]_  | ~\new_[4964]_ ;
  assign \new_[4065]_  = ~\new_[4255]_ ;
  assign \new_[4066]_  = ~\new_[4205]_  | ~\new_[4243]_ ;
  assign \new_[4067]_  = ~\new_[4172]_  | ~\key3[36] ;
  assign \new_[4068]_  = ~\new_[4171]_  & ~\new_[4331]_ ;
  assign \new_[4069]_  = \new_[4131]_ ;
  assign \new_[4070]_  = ~\new_[4251]_  | ~\new_[4187]_ ;
  assign \new_[4071]_  = ~\new_[4243]_  | ~\new_[4202]_ ;
  assign \new_[4072]_  = ~\new_[4243]_  | ~\new_[4202]_ ;
  assign \new_[4073]_  = ~\new_[4171]_  & ~\new_[4360]_ ;
  assign \new_[4074]_  = ~\new_[5174]_ ;
  assign \new_[4075]_  = ~\new_[4213]_  | ~\new_[4964]_ ;
  assign \new_[4076]_  = ~\new_[4243]_  | ~\new_[4202]_ ;
  assign \new_[4077]_  = ~\new_[4213]_  | ~\new_[4202]_ ;
  assign \new_[4078]_  = ~\new_[4230]_  | ~\new_[4159]_ ;
  assign \new_[4079]_  = ~\new_[4156]_ ;
  assign \new_[4080]_  = ~\new_[4131]_ ;
  assign \new_[4081]_  = ~\new_[4213]_  | ~\new_[4202]_ ;
  assign \new_[4082]_  = ~\new_[4243]_  | ~\new_[4205]_ ;
  assign \new_[4083]_  = ~\new_[4138]_ ;
  assign \new_[4084]_  = ~\new_[4213]_  | ~\new_[4202]_ ;
  assign \new_[4085]_  = ~\new_[4125]_ ;
  assign \new_[4086]_  = ~\new_[4213]_  | ~\new_[4202]_ ;
  assign \new_[4087]_  = ~\new_[4187]_  | ~\new_[4225]_ ;
  assign \new_[4088]_  = ~\new_[4138]_ ;
  assign \new_[4089]_  = ~\new_[4230]_  | ~\new_[4159]_ ;
  assign \new_[4090]_  = ~\new_[4213]_  | ~\new_[4202]_ ;
  assign \new_[4091]_  = ~\new_[4171]_  & ~\new_[4340]_ ;
  assign \new_[4092]_  = ~\new_[4171]_  & ~\new_[4330]_ ;
  assign \new_[4093]_  = ~\new_[4969]_  | ~\new_[4201]_ ;
  assign \new_[4094]_  = ~\new_[4230]_  | ~\new_[4159]_ ;
  assign \new_[4095]_  = ~\new_[4213]_  | ~\new_[4202]_ ;
  assign \new_[4096]_  = ~\new_[4243]_  | ~\new_[4202]_ ;
  assign \new_[4097]_  = ~\new_[4243]_  | ~\new_[4205]_ ;
  assign \new_[4098]_  = ~\new_[4178]_ ;
  assign \new_[4099]_  = ~\new_[4187]_  | ~\new_[4225]_ ;
  assign \new_[4100]_  = ~\new_[4230]_  | ~\new_[4159]_ ;
  assign \new_[4101]_  = ~\new_[4194]_ ;
  assign \new_[4102]_  = ~\new_[4179]_ ;
  assign \new_[4103]_  = ~\new_[4191]_ ;
  assign \new_[4104]_  = ~\new_[4170]_ ;
  assign \new_[4105]_  = ~\new_[4191]_ ;
  assign \new_[4106]_  = ~\new_[4349]_  | ~\new_[4261]_  | ~\new_[4329]_ ;
  assign \new_[4107]_  = ~\new_[4258]_  & ~\new_[4344]_ ;
  assign \new_[4108]_  = ~\new_[4164]_ ;
  assign \new_[4109]_  = ~\new_[4167]_ ;
  assign \new_[4110]_  = ~\new_[4175]_ ;
  assign \new_[4111]_  = ~\new_[4243]_  & ~\new_[4334]_ ;
  assign \new_[4112]_  = ~\new_[4175]_ ;
  assign \new_[4113]_  = ~\new_[4271]_ ;
  assign \new_[4114]_  = ~\new_[4254]_  & ~\new_[4307]_ ;
  assign \new_[4115]_  = ~\new_[4215]_ ;
  assign \new_[4116]_  = ~\new_[4169]_ ;
  assign \new_[4117]_  = ~\new_[4165]_ ;
  assign \new_[4118]_  = ~\new_[4189]_ ;
  assign \new_[4119]_  = ~\new_[4246]_  | ~\key3[48] ;
  assign \new_[4120]_  = ~\new_[4195]_ ;
  assign \new_[4121]_  = ~\new_[4792]_ ;
  assign \new_[4122]_  = ~\new_[4168]_ ;
  assign \new_[4123]_  = ~\new_[4165]_ ;
  assign \new_[4124]_  = ~\new_[4175]_ ;
  assign \new_[4125]_  = \new_[4190]_ ;
  assign \new_[4126]_  = ~\new_[4259]_ ;
  assign \new_[4127]_  = ~\new_[4254]_  & ~\new_[4350]_ ;
  assign \new_[4128]_  = ~\new_[4183]_ ;
  assign \new_[4129]_  = ~\new_[4254]_  & ~\new_[4368]_ ;
  assign \new_[4130]_  = ~\new_[4182]_ ;
  assign \new_[4131]_  = \new_[4176]_ ;
  assign \new_[4132]_  = ~\new_[4254]_  & ~\new_[4317]_ ;
  assign \new_[4133]_  = ~\new_[4162]_ ;
  assign \new_[4134]_  = ~\new_[4274]_  | ~\new_[4285]_  | ~\key1[36]  | ~\new_[4286]_ ;
  assign \new_[4135]_  = ~\new_[4190]_ ;
  assign \new_[4136]_  = ~\new_[4217]_  | ~\key3[47] ;
  assign \new_[4137]_  = ~\new_[4194]_ ;
  assign \new_[4138]_  = ~\new_[4194]_ ;
  assign \new_[4139]_  = ~\new_[4160]_ ;
  assign \new_[4140]_  = ~\new_[4162]_ ;
  assign \new_[4141]_  = ~\new_[4225]_  | ~\new_[5225]_ ;
  assign \new_[4142]_  = ~\new_[4287]_  | ~\new_[4224]_  | ~\new_[4288]_ ;
  assign \new_[4143]_  = ~\new_[5097]_ ;
  assign \new_[4144]_  = ~\new_[4195]_ ;
  assign \new_[4145]_  = ~\new_[4254]_  & ~\new_[4367]_ ;
  assign \new_[4146]_  = ~\new_[4254]_  & ~\new_[4374]_ ;
  assign \new_[4147]_  = ~\new_[4258]_  & ~\new_[4364]_ ;
  assign \new_[4148]_  = ~\new_[4183]_ ;
  assign \new_[4149]_  = ~\new_[4182]_ ;
  assign \new_[4150]_  = ~\new_[4176]_ ;
  assign \new_[4151]_  = ~\new_[4254]_  & ~\new_[4366]_ ;
  assign \new_[4152]_  = ~\new_[4167]_ ;
  assign \new_[4153]_  = ~\new_[4182]_ ;
  assign \new_[4154]_  = ~\new_[4165]_ ;
  assign \new_[4155]_  = ~\new_[4191]_ ;
  assign \new_[4156]_  = ~\new_[4195]_ ;
  assign \new_[4157]_  = ~\new_[4258]_  & ~\new_[4345]_ ;
  assign \new_[4158]_  = \new_[5175]_ ;
  assign \new_[4159]_  = ~\new_[4965]_ ;
  assign \new_[4160]_  = ~\new_[4259]_ ;
  assign \new_[4161]_  = ~\new_[4238]_ ;
  assign \new_[4162]_  = ~\new_[4215]_ ;
  assign \new_[4163]_  = ~\new_[4220]_ ;
  assign \new_[4164]_  = ~\new_[4215]_ ;
  assign \new_[4165]_  = ~\new_[4221]_ ;
  assign \new_[4166]_  = ~\new_[4253]_ ;
  assign \new_[4167]_  = ~\new_[4235]_ ;
  assign \new_[4168]_  = ~\new_[4239]_ ;
  assign \new_[4169]_  = ~\new_[4235]_ ;
  assign \new_[4170]_  = ~\new_[4259]_ ;
  assign \new_[4171]_  = ~\new_[4219]_ ;
  assign \new_[4172]_  = ~\new_[4258]_ ;
  assign \new_[4173]_  = ~\new_[4244]_ ;
  assign \new_[4174]_  = \new_[4216]_ ;
  assign \new_[4175]_  = ~\new_[5225]_ ;
  assign \new_[4176]_  = ~\new_[4210]_ ;
  assign \new_[4177]_  = ~\new_[4245]_ ;
  assign \new_[4178]_  = ~\new_[4242]_ ;
  assign \new_[4179]_  = ~\new_[4228]_ ;
  assign \new_[4180]_  = ~\new_[4121]_ ;
  assign \new_[4181]_  = ~\new_[4235]_ ;
  assign \new_[4182]_  = ~\new_[4221]_ ;
  assign \new_[4183]_  = ~\new_[4221]_ ;
  assign \new_[4184]_  = ~\new_[4240]_ ;
  assign \new_[4185]_  = ~\new_[4211]_ ;
  assign \new_[4186]_  = ~\new_[4255]_ ;
  assign \new_[4187]_  = \new_[5225]_ ;
  assign \new_[4188]_  = ~\new_[4238]_ ;
  assign \new_[4189]_  = ~\new_[4226]_ ;
  assign \new_[4190]_  = \new_[4235]_ ;
  assign \new_[4191]_  = ~\new_[5225]_ ;
  assign \new_[4192]_  = ~\new_[4250]_ ;
  assign \new_[4193]_  = ~\new_[4414]_  & (~\new_[4286]_  | ~\new_[4282]_ );
  assign \new_[4194]_  = \new_[4218]_ ;
  assign \new_[4195]_  = ~\new_[4218]_ ;
  assign \new_[4196]_  = ~\new_[4238]_ ;
  assign \new_[4197]_  = ~\new_[4214]_ ;
  assign \new_[4198]_  = ~\new_[4211]_ ;
  assign \new_[4199]_  = ~\new_[4211]_ ;
  assign \new_[4200]_  = ~\new_[4255]_ ;
  assign \new_[4201]_  = ~\new_[4965]_ ;
  assign \new_[4202]_  = ~\new_[4965]_ ;
  assign \new_[4203]_  = ~\new_[4233]_ ;
  assign \new_[4204]_  = ~\new_[4247]_ ;
  assign \new_[4205]_  = ~\new_[4965]_ ;
  assign \new_[4206]_  = ~\new_[4259]_ ;
  assign \new_[4207]_  = ~\new_[4259]_ ;
  assign \new_[4208]_  = \new_[4242]_ ;
  assign \new_[4209]_  = ~\new_[4247]_ ;
  assign \new_[4210]_  = ~\new_[4290]_  | ~\new_[4275]_ ;
  assign \new_[4211]_  = ~\new_[5175]_ ;
  assign \new_[4212]_  = ~\new_[5098]_ ;
  assign \new_[4213]_  = ~\new_[4968]_ ;
  assign \new_[4214]_  = ~\new_[4264]_ ;
  assign \new_[4215]_  = \new_[4275]_  & \new_[4280]_ ;
  assign \new_[4216]_  = ~\new_[4269]_ ;
  assign \new_[4217]_  = \new_[4266]_ ;
  assign \new_[4218]_  = ~\new_[4406]_ ;
  assign \new_[4219]_  = ~\new_[4265]_ ;
  assign \new_[4220]_  = \new_[4698]_ ;
  assign \new_[4221]_  = \new_[4406]_ ;
  assign \new_[4222]_  = ~\new_[4271]_ ;
  assign \new_[4223]_  = \new_[4281]_  | \new_[4277]_ ;
  assign \new_[4224]_  = \new_[4274]_  & \new_[4285]_ ;
  assign \new_[4225]_  = ~\new_[4273]_ ;
  assign \new_[4226]_  = ~\new_[4268]_ ;
  assign \new_[4227]_  = \new_[4266]_ ;
  assign \new_[4228]_  = \new_[4262]_ ;
  assign \new_[4229]_  = ~\new_[5228]_ ;
  assign \new_[4230]_  = ~\new_[4968]_ ;
  assign \new_[4231]_  = ~\new_[4272]_ ;
  assign \new_[4232]_  = \new_[4262]_ ;
  assign \new_[4233]_  = ~\new_[4269]_ ;
  assign \new_[4234]_  = ~\new_[4267]_ ;
  assign \new_[4235]_  = \new_[4275]_  & \new_[4288]_ ;
  assign \new_[4236]_  = ~\new_[5228]_ ;
  assign \new_[4237]_  = ~\new_[4264]_ ;
  assign \new_[4238]_  = ~\new_[4698]_ ;
  assign \new_[4239]_  = ~\new_[4272]_ ;
  assign \new_[4240]_  = ~\new_[4272]_ ;
  assign \new_[4241]_  = ~\new_[4269]_ ;
  assign \new_[4242]_  = ~\new_[4263]_ ;
  assign \new_[4243]_  = ~\new_[4968]_ ;
  assign \new_[4244]_  = ~\new_[5175]_ ;
  assign \new_[4245]_  = ~\new_[4792]_ ;
  assign \new_[4246]_  = ~\new_[4265]_ ;
  assign \new_[4247]_  = ~\new_[5068]_ ;
  assign \new_[4248]_  = ~\new_[4269]_ ;
  assign \new_[4249]_  = ~\new_[4271]_ ;
  assign \new_[4250]_  = ~\new_[4269]_ ;
  assign \new_[4251]_  = ~\new_[4267]_ ;
  assign \new_[4252]_  = ~\new_[4272]_ ;
  assign \new_[4253]_  = ~\new_[4270]_ ;
  assign \new_[4254]_  = \new_[4265]_ ;
  assign \new_[4255]_  = ~\new_[4262]_ ;
  assign \new_[4256]_  = ~\new_[4264]_ ;
  assign \new_[4257]_  = ~\new_[4287]_  | ~\new_[4277]_ ;
  assign \new_[4258]_  = ~\new_[4266]_ ;
  assign \new_[4259]_  = ~\new_[4275]_  | ~\new_[4283]_ ;
  assign \new_[4260]_  = \new_[4266]_ ;
  assign \new_[4261]_  = ~\new_[4274]_ ;
  assign \new_[4262]_  = \new_[4290]_  & \new_[4284]_ ;
  assign \new_[4263]_  = ~\new_[4288]_  | ~\new_[4287]_ ;
  assign \new_[4264]_  = ~\new_[4276]_ ;
  assign \new_[4265]_  = \new_[4843]_ ;
  assign \new_[4266]_  = ~\new_[4843]_ ;
  assign \new_[4267]_  = ~\new_[5229]_ ;
  assign \new_[4268]_  = ~\new_[4279]_  | ~\new_[4280]_ ;
  assign \new_[4269]_  = ~\new_[4280]_  | ~\new_[4287]_ ;
  assign \new_[4270]_  = \new_[4276]_ ;
  assign \new_[4271]_  = ~\new_[4290]_  | ~\new_[4279]_ ;
  assign \new_[4272]_  = ~\new_[4283]_  | ~\new_[4284]_ ;
  assign \new_[4273]_  = ~\new_[5229]_ ;
  assign \new_[4274]_  = ~\new_[4278]_ ;
  assign \new_[4275]_  = \roundSel[2]  & \roundSel[3] ;
  assign \new_[4276]_  = \new_[4290]_  & \new_[4287]_ ;
  assign \new_[4277]_  = ~\new_[4285]_ ;
  assign \new_[4278]_  = ~\new_[4635]_ ;
  assign \new_[4279]_  = ~\new_[4314]_  & ~\roundSel[3] ;
  assign \new_[4280]_  = ~\roundSel[0]  & ~\new_[4349]_ ;
  assign \new_[4281]_  = ~\new_[4287]_ ;
  assign \new_[4282]_  = ~\new_[4286]_ ;
  assign \new_[4283]_  = ~\roundSel[1]  & ~\new_[4329]_ ;
  assign \new_[4284]_  = \new_[4314]_  & \roundSel[3] ;
  assign \new_[4285]_  = ~\new_[4289]_ ;
  assign \new_[4286]_  = ~\new_[4321]_ ;
  assign \new_[4287]_  = ~\roundSel[2]  & ~\roundSel[3] ;
  assign \new_[4288]_  = ~\roundSel[0]  & ~\roundSel[1] ;
  assign \new_[4289]_  = ~\new_[4967]_ ;
  assign \new_[4290]_  = \roundSel[0]  & \roundSel[1] ;
  assign \new_[4291]_  = ~\key3[49] ;
  assign \new_[4292]_  = ~\key2[40] ;
  assign \new_[4293]_  = ~\key3[46] ;
  assign \new_[4294]_  = ~\key2[1] ;
  assign \new_[4295]_  = ~\key3[24] ;
  assign \new_[4296]_  = ~\desIn[26] ;
  assign \new_[4297]_  = ~\desIn[12] ;
  assign \new_[4298]_  = ~\key3[34] ;
  assign \new_[4299]_  = ~\new_[2207]_ ;
  assign \new_[4300]_  = ~\key3[23] ;
  assign \new_[4301]_  = ~\key2[33] ;
  assign \new_[4302]_  = ~\key3[17] ;
  assign \new_[4303]_  = ~\new_[502]_ ;
  assign \new_[4304]_  = ~\new_[435]_ ;
  assign \new_[4305]_  = ~\key3[4] ;
  assign \new_[4306]_  = ~\key3[29] ;
  assign \new_[4307]_  = ~\key3[18] ;
  assign \new_[4308]_  = ~\key3[33] ;
  assign \new_[4309]_  = ~\key3[54] ;
  assign \new_[4310]_  = ~\desIn[4] ;
  assign \new_[4311]_  = ~\desIn[24] ;
  assign \new_[4312]_  = ~\key2[52] ;
  assign \new_[4313]_  = ~\new_[485]_ ;
  assign \new_[4314]_  = ~\roundSel[2] ;
  assign \new_[4315]_  = ~\key3[10] ;
  assign \new_[4316]_  = ~\desIn[58] ;
  assign \new_[4317]_  = ~\key3[41] ;
  assign \new_[4318]_  = ~\key3[39] ;
  assign \new_[4319]_  = ~\new_[506]_ ;
  assign \new_[4320]_  = ~\new_[2159]_ ;
  assign \new_[4321]_  = ~decrypt;
  assign \new_[4322]_  = ~\key2[24] ;
  assign \new_[4323]_  = ~\key2[39] ;
  assign \new_[4324]_  = ~\new_[453]_ ;
  assign \new_[4325]_  = ~\key3[36] ;
  assign \new_[4326]_  = ~\key3[20] ;
  assign \new_[4327]_  = ~\key3[27] ;
  assign \new_[4328]_  = ~\key3[25] ;
  assign \new_[4329]_  = ~\roundSel[0] ;
  assign \new_[4330]_  = ~\key3[16] ;
  assign \new_[4331]_  = ~\key3[44] ;
  assign \new_[4332]_  = ~\key3[21] ;
  assign \new_[4333]_  = ~\new_[457]_ ;
  assign \new_[4334]_  = ~\key1[36] ;
  assign \new_[4335]_  = ~\desIn[40] ;
  assign \new_[4336]_  = ~\new_[2155]_ ;
  assign \new_[4337]_  = ~\key3[11] ;
  assign \new_[4338]_  = ~\new_[450]_ ;
  assign \new_[4339]_  = ~\new_[458]_ ;
  assign \new_[4340]_  = ~\key3[45] ;
  assign \new_[4341]_  = ~\key3[1] ;
  assign \new_[4342]_  = ~\key3[52] ;
  assign \new_[4343]_  = ~\new_[2161]_ ;
  assign \new_[4344]_  = ~\key3[37] ;
  assign \new_[4345]_  = ~\key3[40] ;
  assign \new_[4346]_  = ~\new_[501]_ ;
  assign \new_[4347]_  = ~\key3[43] ;
  assign \new_[4348]_  = ~\key3[50] ;
  assign \new_[4349]_  = ~\roundSel[1] ;
  assign \new_[4350]_  = ~\key3[5] ;
  assign \new_[4351]_  = ~\key3[9] ;
  assign \new_[4352]_  = ~\key3[55] ;
  assign \new_[4353]_  = ~\desIn[38] ;
  assign \new_[4354]_  = ~\key3[32] ;
  assign \new_[4355]_  = ~\new_[2158]_ ;
  assign \new_[4356]_  = ~\new_[2376]_ ;
  assign \new_[4357]_  = ~\desIn[60] ;
  assign \new_[4358]_  = ~\desIn[36] ;
  assign \new_[4359]_  = ~\desIn[2] ;
  assign \new_[4360]_  = ~\key3[8] ;
  assign \new_[4361]_  = ~\desIn[52] ;
  assign \new_[4362]_  = ~\desIn[50] ;
  assign \new_[4363]_  = ~\desIn[42] ;
  assign \new_[4364]_  = ~\key3[15] ;
  assign \new_[4365]_  = ~\key3[7] ;
  assign \new_[4366]_  = ~\key3[35] ;
  assign \new_[4367]_  = ~\key3[6] ;
  assign \new_[4368]_  = ~\key3[30] ;
  assign \new_[4369]_  = ~\key3[51] ;
  assign \new_[4370]_  = ~\new_[489]_ ;
  assign \new_[4371]_  = ~\new_[480]_ ;
  assign \new_[4372]_  = ~\new_[2023]_ ;
  assign \new_[4373]_  = ~\new_[2016]_ ;
  assign \new_[4374]_  = ~\key3[2] ;
  assign \new_[4375]_  = ~\desIn[14] ;
  assign \new_[4376]_  = ~\new_[2160]_ ;
  assign \new_[4377]_  = ~\new_[4378]_ ;
  assign \new_[4378]_  = ~\new_[4672]_ ;
  assign \new_[4379]_  = ~\new_[4381]_ ;
  assign \new_[4380]_  = ~\new_[4381]_ ;
  assign \new_[4381]_  = ~\new_[3639]_ ;
  assign \new_[4382]_  = \new_[3726]_ ;
  assign \new_[4383]_  = \new_[3726]_ ;
  assign \new_[4384]_  = \new_[3640]_ ;
  assign \new_[4385]_  = \new_[4657]_ ;
  assign \new_[4386]_  = \new_[3615]_ ;
  assign \new_[4387]_  = \new_[3615]_ ;
  assign \new_[4388]_  = ~\new_[4389]_ ;
  assign \new_[4389]_  = \new_[5155]_ ;
  assign \new_[4390]_  = ~\new_[5161]_ ;
  assign \new_[4391]_  = ~\new_[5154]_ ;
  assign \new_[4392]_  = \new_[4723]_ ;
  assign \new_[4393]_  = \new_[4394]_ ;
  assign \new_[4394]_  = \new_[4762]_ ;
  assign \new_[4395]_  = \new_[4762]_ ;
  assign \new_[4396]_  = \new_[4762]_ ;
  assign \new_[4397]_  = ~\new_[4398]_ ;
  assign \new_[4398]_  = ~\new_[4399]_ ;
  assign \new_[4399]_  = ~\new_[1646]_ ;
  assign \new_[4400]_  = \new_[1646]_ ;
  assign \new_[4401]_  = \new_[3613]_ ;
  assign \new_[4402]_  = \new_[4403]_ ;
  assign \new_[4403]_  = ~\new_[4404]_ ;
  assign \new_[4404]_  = ~\new_[3613]_ ;
  assign \new_[4405]_  = \new_[3649]_ ;
  assign \new_[4406]_  = ~\new_[4407]_  | ~\new_[4408]_ ;
  assign \new_[4407]_  = ~\new_[4970]_ ;
  assign \new_[4408]_  = ~decrypt & ~\roundSel[4] ;
  assign n665 = \new_[4410]_  ? \new_[4993]_  : \new_[4411]_ ;
  assign \new_[4410]_  = ~\new_[4411]_ ;
  assign \new_[4411]_  = (~\desIn[30]  | ~\new_[2908]_ ) & (~\new_[2284]_  | ~\new_[2898]_ );
  assign \new_[4412]_  = ~\new_[4413]_  | ~\roundSel[4] ;
  assign \new_[4413]_  = ~\roundSel[5] ;
  assign \new_[4414]_  = ~\new_[4413]_  | ~\roundSel[4] ;
  assign \new_[4415]_  = ~\new_[770]_  | ~\new_[895]_ ;
  assign \new_[4416]_  = ~\new_[890]_  | ~\new_[958]_ ;
  assign \new_[4417]_  = ~\new_[4462]_ ;
  assign \new_[4418]_  = ~\new_[1253]_  | ~\new_[906]_  | ~\new_[1059]_ ;
  assign \new_[4419]_  = \new_[1179]_  & \new_[4462]_ ;
  assign \new_[4420]_  = ~\new_[934]_  | ~\new_[754]_  | ~\new_[1078]_ ;
  assign n615 = \new_[4422]_  ? \new_[4424]_  : \new_[4423]_ ;
  assign \new_[4422]_  = (~\desIn[0]  | ~\new_[2639]_ ) & (~\new_[1765]_  | ~\new_[2898]_ );
  assign \new_[4423]_  = ~\new_[4422]_ ;
  assign \new_[4424]_  = ~\new_[4425]_  & ~\new_[529]_ ;
  assign \new_[4425]_  = ~\new_[4428]_  | ~\new_[4426]_  | ~\new_[4427]_ ;
  assign \new_[4426]_  = ~\new_[569]_ ;
  assign \new_[4427]_  = ~\new_[767]_ ;
  assign \new_[4428]_  = ~\new_[956]_ ;
  assign n785 = \new_[4430]_  ? \new_[4432]_  : \new_[4431]_ ;
  assign \new_[4430]_  = ~\new_[4431]_ ;
  assign \new_[4431]_  = (~\desIn[8]  | ~\new_[2908]_ ) & (~\new_[1764]_  | ~\new_[2871]_ );
  assign \new_[4432]_  = ~\new_[531]_  | ~\new_[772]_ ;
  assign n760 = \new_[4434]_  ? \new_[4436]_  : \new_[4435]_ ;
  assign \new_[4434]_  = ~\new_[4435]_ ;
  assign \new_[4435]_  = (~\desIn[48]  | ~\new_[2908]_ ) & (~\new_[1752]_  | ~\new_[2898]_ );
  assign \new_[4436]_  = \new_[544]_  | \new_[4437]_ ;
  assign \new_[4437]_  = ~\new_[560]_  | ~\new_[4438]_ ;
  assign \new_[4438]_  = ~\new_[4490]_  & ~\new_[905]_ ;
  assign \new_[4439]_  = \new_[4440]_  & \new_[2517]_ ;
  assign \new_[4440]_  = ~\new_[2706]_  & ~\new_[4441]_ ;
  assign \new_[4441]_  = ~\new_[2913]_ ;
  assign \new_[4442]_  = ~\new_[2286]_  & (~\new_[3033]_  | ~\new_[4228]_ );
  assign \new_[4443]_  = ~\new_[4444]_  & (~\new_[2907]_  | ~\new_[4140]_ );
  assign \new_[4444]_  = ~\new_[2425]_  | ~\new_[2451]_ ;
  assign \new_[4445]_  = ~\new_[2704]_  & ~\new_[2285]_ ;
  assign n890 = \new_[4447]_  ? \new_[4449]_  : \new_[4448]_ ;
  assign \new_[4447]_  = ~\new_[4448]_ ;
  assign \new_[4448]_  = (~\desIn[6]  | ~\new_[3713]_ ) & (~\new_[1755]_  | ~\new_[2898]_ );
  assign \new_[4449]_  = ~\new_[556]_  | ~\new_[547]_  | ~\new_[543]_ ;
  assign \new_[4450]_  = ~\new_[4451]_  | ~\new_[4452]_ ;
  assign \new_[4451]_  = ~\new_[855]_  | ~\new_[1027]_ ;
  assign \new_[4452]_  = ~\new_[4721]_ ;
  assign \new_[4453]_  = ~\new_[4962]_ ;
  assign \new_[4454]_  = ~\new_[4455]_  | ~\new_[4456]_ ;
  assign \new_[4455]_  = ~\new_[959]_  | ~\new_[5286]_ ;
  assign \new_[4456]_  = ~\new_[4392]_  | ~\new_[1550]_ ;
  assign \new_[4457]_  = ~\new_[1317]_  | (~\new_[597]_  & ~\new_[684]_ );
  assign \new_[4458]_  = ~\new_[4417]_  | (~\new_[4459]_  & ~\new_[4460]_ );
  assign \new_[4459]_  = ~\new_[628]_  | ~\new_[773]_ ;
  assign \new_[4460]_  = ~\new_[683]_  | ~\new_[4461]_ ;
  assign \new_[4461]_  = ~\new_[5290]_  | ~\new_[5209]_ ;
  assign \new_[4462]_  = n1220 ? \new_[1653]_  : \new_[3290]_ ;
  assign \new_[4463]_  = ~\new_[1179]_  | ~\new_[691]_ ;
  assign \new_[4464]_  = ~n1015;
  assign n1015 = \new_[3573]_  ? \new_[3914]_  : \desIn[25] ;
  assign \new_[4466]_  = ~\new_[4472]_  | ~\new_[4471]_  | ~\new_[4470]_  | ~\new_[4467]_ ;
  assign \new_[4467]_  = \new_[4468]_  & \new_[4469]_ ;
  assign \new_[4468]_  = ~\new_[2798]_  | ~\new_[4166]_ ;
  assign \new_[4469]_  = ~\new_[3088]_  | ~\new_[5068]_ ;
  assign \new_[4470]_  = ~\new_[2128]_  & ~\new_[1905]_ ;
  assign \new_[4471]_  = ~\new_[1940]_  & ~\new_[1941]_ ;
  assign \new_[4472]_  = ~\new_[2718]_  & ~\new_[2663]_ ;
  assign \new_[4473]_  = ~\new_[4478]_  | ~\new_[4474]_  | ~\new_[4477]_ ;
  assign \new_[4474]_  = ~\new_[4475]_  & ~\new_[4476]_ ;
  assign \new_[4475]_  = ~\new_[2899]_  | ~\new_[2381]_  | ~\new_[2888]_ ;
  assign \new_[4476]_  = ~\new_[2469]_  | ~\new_[2468]_  | ~\new_[2428]_ ;
  assign \new_[4477]_  = ~\new_[2089]_  & (~\new_[3099]_  | ~\new_[4160]_ );
  assign \new_[4478]_  = ~\new_[2098]_  & ~\new_[2697]_ ;
  assign n705 = \new_[4480]_  ? \new_[4483]_  : \new_[4481]_ ;
  assign \new_[4480]_  = ~\new_[4481]_ ;
  assign \new_[4481]_  = ~\new_[4482]_  | (~\new_[1767]_  & ~\new_[3713]_ );
  assign \new_[4482]_  = \new_[4353]_  | \new_[3739]_ ;
  assign \new_[4483]_  = ~\new_[686]_  | ~\new_[536]_  | ~\new_[537]_ ;
  assign \new_[4484]_  = ~\new_[4485]_  & (~\new_[4420]_  | ~\new_[4462]_ );
  assign \new_[4485]_  = \new_[704]_  & \new_[5209]_ ;
  assign \new_[4486]_  = ~\new_[4417]_  | (~\new_[665]_  & ~\new_[738]_ );
  assign \new_[4487]_  = ~\new_[4488]_  & (~\new_[4419]_  | ~\new_[4418]_ );
  assign \new_[4488]_  = ~\new_[5291]_  & ~\new_[1421]_  & ~\new_[1521]_ ;
  assign \new_[4489]_  = ~\new_[4490]_  & ~\new_[667]_ ;
  assign \new_[4490]_  = ~\new_[1163]_  & ~\new_[1426]_  & ~\new_[1580]_ ;
  assign \new_[4491]_  = ~\new_[4497]_  | ~\new_[4496]_  | ~\new_[4492]_  | ~\new_[4494]_ ;
  assign \new_[4492]_  = ~\new_[4493]_ ;
  assign \new_[4493]_  = ~\new_[1516]_  & (~\new_[1151]_  | ~\new_[1152]_ );
  assign \new_[4494]_  = ~\new_[4495]_  & (~\new_[5082]_  | ~\new_[1089]_ );
  assign \new_[4495]_  = ~\new_[4604]_  & ~\new_[1481]_  & ~\new_[5083]_ ;
  assign \new_[4496]_  = ~\new_[1180]_  | ~\new_[1532]_ ;
  assign \new_[4497]_  = ~\new_[1482]_  | ~\new_[1028]_  | ~\new_[4649]_ ;
  assign \new_[4498]_  = ~\new_[4499]_ ;
  assign \new_[4499]_  = ~\new_[2334]_  | (~\new_[1744]_  & ~\new_[3713]_ );
  assign \new_[4500]_  = ~\new_[594]_  | ~\new_[585]_  | ~\new_[533]_  | ~\new_[532]_ ;
  assign \new_[4501]_  = ~\new_[4511]_  | ~\new_[4509]_  | ~\new_[4502]_  | ~\new_[4507]_ ;
  assign \new_[4502]_  = ~\new_[4503]_ ;
  assign \new_[4503]_  = ~\new_[4504]_  | ~\new_[4505]_ ;
  assign \new_[4504]_  = ~\new_[3009]_  | ~\new_[4214]_ ;
  assign \new_[4505]_  = ~\new_[4506]_  & ~\new_[2455]_ ;
  assign \new_[4506]_  = ~\new_[2411]_  | ~\new_[2410]_ ;
  assign \new_[4507]_  = ~\new_[4508]_  & ~\new_[1982]_ ;
  assign \new_[4508]_  = ~\new_[2344]_  | ~\new_[2369]_ ;
  assign \new_[4509]_  = ~\new_[2197]_  & ~\new_[4510]_ ;
  assign \new_[4510]_  = ~\new_[2345]_ ;
  assign \new_[4511]_  = ~\new_[2009]_  & (~\new_[2841]_  | ~\new_[3985]_ );
  assign n675 = \new_[4513]_  ? \new_[4515]_  : \new_[4514]_ ;
  assign \new_[4513]_  = ~\new_[4514]_ ;
  assign \new_[4514]_  = ~\new_[2332]_  | (~\new_[1798]_  & ~\new_[3713]_ );
  assign \new_[4515]_  = ~\new_[4516]_  | ~\new_[527]_  | ~\new_[545]_ ;
  assign \new_[4516]_  = \new_[745]_  & \new_[1049]_ ;
  assign \new_[4517]_  = ~\new_[4518]_ ;
  assign \new_[4518]_  = ~\new_[5174]_  & (~\new_[3331]_  | ~\new_[3406]_ );
  assign \new_[4519]_  = ~\new_[2511]_ ;
  assign \new_[4520]_  = ~\new_[2050]_  | ~\new_[4521]_ ;
  assign \new_[4521]_  = ~\new_[2512]_  & (~\new_[2818]_  | ~\new_[4021]_ );
  assign \new_[4522]_  = ~\new_[2282]_  | ~\new_[4170]_ ;
  assign \new_[4523]_  = ~\new_[2202]_ ;
  assign \new_[4524]_  = ~\new_[4530]_  | ~\new_[4525]_  | ~\new_[4529]_ ;
  assign \new_[4525]_  = ~\new_[4528]_  | (~\new_[4526]_  & ~\new_[4527]_ );
  assign \new_[4526]_  = ~\new_[1021]_  | ~\new_[4603]_  | ~\new_[743]_  | ~\new_[687]_ ;
  assign \new_[4527]_  = ~\new_[1199]_  | ~\new_[740]_ ;
  assign \new_[4528]_  = ~\new_[5126]_ ;
  assign \new_[4529]_  = ~\new_[4491]_  | ~\new_[5126]_ ;
  assign \new_[4530]_  = ~\new_[647]_  & (~\new_[759]_  | ~\new_[5081]_ );
  assign \new_[4531]_  = ~\new_[4538]_  | ~\new_[4536]_  | ~\new_[4532]_  | ~\new_[4533]_ ;
  assign \new_[4532]_  = ~\new_[572]_  | ~\new_[1307]_ ;
  assign \new_[4533]_  = ~\new_[4534]_  | ~\new_[4535]_ ;
  assign \new_[4534]_  = ~\new_[1118]_  | ~\new_[769]_  | ~\new_[801]_  | ~\new_[700]_ ;
  assign \new_[4535]_  = ~\new_[1561]_  | ~\new_[1560]_ ;
  assign \new_[4536]_  = ~\new_[4537]_  | ~\new_[1430]_ ;
  assign \new_[4537]_  = ~\new_[1117]_ ;
  assign \new_[4538]_  = ~\new_[587]_  & (~\new_[1161]_  | ~\new_[1157]_ );
  assign \new_[4539]_  = ~\new_[4540]_ ;
  assign \new_[4540]_  = (~\desIn[16]  | ~\new_[2639]_ ) & (~\new_[1746]_  | ~\new_[2898]_ );
  assign \new_[4541]_  = ~\new_[4542]_  & ~\new_[2501]_ ;
  assign \new_[4542]_  = ~\new_[2499]_  | ~\new_[2643]_ ;
  assign \new_[4543]_  = ~\new_[4544]_  & ~\new_[1945]_ ;
  assign \new_[4544]_  = ~\new_[2443]_  | ~\new_[2904]_ ;
  assign \new_[4545]_  = ~\new_[4546]_  & ~\new_[1946]_ ;
  assign \new_[4546]_  = ~\new_[2500]_  | ~\new_[2905]_ ;
  assign \new_[4547]_  = ~\new_[2568]_  | ~\new_[4240]_ ;
  assign \new_[4548]_  = ~\new_[4783]_ ;
  assign \new_[4549]_  = ~\new_[4550]_  | ~\new_[4551]_ ;
  assign \new_[4550]_  = ~\new_[2736]_ ;
  assign \new_[4551]_  = ~\new_[2817]_  | ~\new_[4222]_ ;
  assign \new_[4552]_  = ~\new_[2200]_  | ~\new_[4553]_ ;
  assign \new_[4553]_  = ~\new_[2815]_  | ~\new_[4160]_ ;
  assign \new_[4554]_  = ~\new_[2190]_  & (~\new_[2954]_  | ~\new_[4237]_ );
  assign \new_[4555]_  = ~\new_[4556]_  & (~\new_[2936]_  | ~\new_[4199]_ );
  assign \new_[4556]_  = ~\new_[2309]_  | ~\new_[2481]_ ;
  assign \new_[4557]_  = ~\new_[4558]_  & ~\new_[2308]_ ;
  assign \new_[4558]_  = ~\new_[2861]_  | ~\new_[2953]_ ;
  assign \new_[4559]_  = ~\new_[2146]_  & ~\new_[2742]_ ;
  assign \new_[4560]_  = ~\new_[4567]_  | ~\new_[4561]_  | ~\new_[4563]_ ;
  assign \new_[4561]_  = ~\new_[4562]_  & (~\new_[676]_  | ~\new_[1165]_ );
  assign \new_[4562]_  = ~\new_[4528]_  & (~\new_[851]_  | ~\new_[4603]_ );
  assign \new_[4563]_  = ~\new_[4564]_  & (~\new_[864]_  | ~\new_[5081]_ );
  assign \new_[4564]_  = ~\new_[4565]_  & ~\new_[4566]_ ;
  assign \new_[4565]_  = ~\new_[1532]_  & ~\new_[1244]_ ;
  assign \new_[4566]_  = ~\new_[1423]_  | ~\new_[5126]_ ;
  assign \new_[4567]_  = ~\new_[563]_  | ~\new_[4528]_ ;
  assign \new_[4568]_  = ~\new_[4569]_  | ~\new_[4572]_ ;
  assign \new_[4569]_  = \new_[4570]_  ? \new_[4571]_  : n985;
  assign \new_[4570]_  = \new_[3474]_  & \new_[3752]_ ;
  assign \new_[4571]_  = ~\new_[4445]_  | ~\new_[4443]_  | ~\new_[4439]_  | ~\new_[4442]_ ;
  assign \new_[4572]_  = ~\new_[4573]_ ;
  assign \new_[4573]_  = ~\new_[1683]_  | ~\new_[1701]_ ;
  assign \new_[4574]_  = n985 ? \new_[4571]_  : \new_[4570]_ ;
  assign \new_[4575]_  = ~\new_[4576]_  | ~\new_[4579]_ ;
  assign \new_[4576]_  = \new_[4577]_  & \new_[4578]_ ;
  assign \new_[4577]_  = ~\new_[580]_  | ~\new_[4874]_ ;
  assign \new_[4578]_  = ~\new_[611]_  | ~\new_[4873]_ ;
  assign \new_[4579]_  = ~\new_[4580]_  & ~\new_[589]_ ;
  assign \new_[4580]_  = ~\new_[778]_  | ~\new_[5045]_ ;
  assign \new_[4581]_  = ~\new_[705]_  | ~\new_[5189]_ ;
  assign \new_[4582]_  = ~\new_[4577]_  | ~\new_[4578]_ ;
  assign \new_[4583]_  = ~\new_[4744]_  | ~\new_[4584]_ ;
  assign \new_[4584]_  = ~\new_[1320]_ ;
  assign \new_[4585]_  = \new_[5112]_ ;
  assign n720 = \new_[4587]_  ? \new_[4589]_  : \new_[4588]_ ;
  assign \new_[4587]_  = ~\new_[4588]_ ;
  assign \new_[4588]_  = (~\new_[3739]_  & ~\new_[4375]_ ) | (~\new_[1773]_  & ~\new_[3713]_ );
  assign \new_[4589]_  = ~\new_[4590]_  & ~\new_[5117]_ ;
  assign \new_[4590]_  = ~\new_[4528]_  & (~\new_[554]_  | ~\new_[1199]_ );
  assign \new_[4591]_  = ~\new_[4597]_  | ~\new_[4592]_  | ~\new_[4595]_ ;
  assign \new_[4592]_  = ~\new_[4593]_  & ~\new_[2001]_ ;
  assign \new_[4593]_  = ~\new_[4594]_  | ~\new_[2367]_  | ~\new_[2172]_  | ~\new_[2302]_ ;
  assign \new_[4594]_  = ~\new_[2780]_  | ~\new_[4214]_ ;
  assign \new_[4595]_  = ~\new_[1964]_  & ~\new_[4596]_ ;
  assign \new_[4596]_  = \new_[2053]_  | \new_[2422]_ ;
  assign \new_[4597]_  = ~\new_[4598]_  & (~\new_[2565]_  | ~\new_[5068]_ );
  assign \new_[4598]_  = ~\new_[2087]_  | ~\new_[2379]_ ;
  assign \new_[4599]_  = ~\new_[4600]_  & ~\new_[4650]_ ;
  assign \new_[4600]_  = ~\new_[4602]_  | ~\new_[2355]_  | ~\new_[4601]_ ;
  assign \new_[4601]_  = ~\new_[2752]_  & (~\new_[3536]_  | ~\new_[4161]_ );
  assign \new_[4602]_  = ~\new_[2686]_ ;
  assign \new_[4603]_  = ~\new_[4607]_  | ~\new_[4646]_  | ~\new_[4649]_  | ~\new_[4604]_ ;
  assign \new_[4604]_  = ~\new_[4887]_ ;
  assign \new_[4605]_  = ~\new_[1708]_  | ~n1125;
  assign \new_[4606]_  = ~\new_[2700]_  | ~\new_[1724]_ ;
  assign \new_[4607]_  = ~\new_[4890]_ ;
  assign \new_[4608]_  = ~\new_[4646]_ ;
  assign \new_[4609]_  = ~\new_[1723]_  | ~n1130;
  assign \new_[4610]_  = ~\new_[2792]_  | ~\new_[1737]_ ;
  assign \new_[4611]_  = ~\new_[4708]_ ;
  assign \new_[4612]_  = ~\new_[4623]_  | ~\new_[4615]_  | ~\new_[4613]_ ;
  assign \new_[4613]_  = \new_[4614]_ ;
  assign \new_[4614]_  = ~\new_[4672]_ ;
  assign \new_[4615]_  = ~\new_[4616]_ ;
  assign \new_[4616]_  = ~\new_[4617]_ ;
  assign \new_[4617]_  = ~\new_[4618]_ ;
  assign \new_[4618]_  = ~\new_[4619]_ ;
  assign \new_[4619]_  = \new_[4620]_  ? \new_[4622]_  : n1245;
  assign \new_[4620]_  = ~n1245;
  assign n1245 = \new_[3766]_  ? \new_[3837]_  : \desIn[5] ;
  assign \new_[4622]_  = ~\new_[1993]_  | ~\new_[1824]_  | ~\new_[1850]_  | ~\new_[1904]_ ;
  assign \new_[4623]_  = ~\new_[4624]_ ;
  assign \new_[4624]_  = ~\new_[4625]_ ;
  assign \new_[4625]_  = ~\new_[4626]_ ;
  assign \new_[4626]_  = ~\new_[4627]_ ;
  assign \new_[4627]_  = \new_[2669]_  ? \new_[1734]_  : n1135;
  assign \new_[4628]_  = \new_[4618]_ ;
  assign \new_[4629]_  = ~\new_[4630]_ ;
  assign \new_[4630]_  = (~\desIn[62]  | ~\new_[2639]_ ) & (~\new_[1768]_  | ~\new_[2898]_ );
  assign \new_[4631]_  = ~\new_[2257]_  | ~\new_[4632]_ ;
  assign \new_[4632]_  = (~\new_[4108]_  | ~\new_[3098]_ ) & (~\new_[2631]_  | ~\new_[4220]_ );
  assign \new_[4633]_  = ~\new_[2256]_ ;
  assign \new_[4634]_  = ~\new_[2528]_ ;
  assign \new_[4635]_  = ~\new_[4970]_ ;
  assign \new_[4636]_  = ~\new_[4638]_  | ~\new_[4637]_  | ~\new_[2201]_ ;
  assign \new_[4637]_  = ~\new_[2513]_  & ~\new_[2237]_ ;
  assign \new_[4638]_  = ~\new_[2572]_  | ~\new_[4245]_ ;
  assign \new_[4639]_  = ~\new_[2573]_  | ~\new_[4098]_ ;
  assign \new_[4640]_  = n1240 ? \new_[4641]_  : \new_[4905]_ ;
  assign \new_[4641]_  = ~\new_[1870]_  & ~\new_[1788]_ ;
  assign \new_[4642]_  = ~\new_[4644]_  | ~\new_[4649]_  | ~\new_[5083]_  | ~\new_[4604]_ ;
  assign \new_[4643]_  = \new_[4885]_ ;
  assign \new_[4644]_  = ~\new_[4645]_ ;
  assign \new_[4645]_  = \new_[4646]_ ;
  assign \new_[4646]_  = ~\new_[4647]_ ;
  assign \new_[4647]_  = ~\new_[4836]_  | ~\new_[1732]_ ;
  assign \new_[4648]_  = ~\new_[4837]_  | ~\new_[1732]_ ;
  assign \new_[4649]_  = ~\new_[4643]_ ;
  assign \new_[4650]_  = ~\new_[4655]_  | ~\new_[4654]_  | ~\new_[4651]_  | ~\new_[4653]_ ;
  assign \new_[4651]_  = ~\new_[4652]_  & ~\new_[2612]_ ;
  assign \new_[4652]_  = ~\new_[2984]_  | ~\new_[3209]_ ;
  assign \new_[4653]_  = ~\new_[3138]_  | ~\new_[4233]_ ;
  assign \new_[4654]_  = ~\new_[2617]_  & ~\new_[2764]_ ;
  assign \new_[4655]_  = ~\new_[4656]_  & ~\new_[2758]_ ;
  assign \new_[4656]_  = ~\new_[2910]_  | ~\new_[2966]_ ;
  assign \new_[4657]_  = ~\new_[5295]_  | ~\new_[4658]_ ;
  assign \new_[4658]_  = ~\new_[4659]_  | ~\new_[4660]_ ;
  assign \new_[4659]_  = ~\new_[3994]_  & (~\new_[4004]_  | ~\key2[6] );
  assign \new_[4660]_  = ~\new_[4145]_  & (~\new_[4054]_  | ~\key1[6] );
  assign \new_[4661]_  = ~\new_[4662]_ ;
  assign \new_[4662]_  = ~\new_[4663]_ ;
  assign \new_[4663]_  = ~\new_[5105]_ ;
  assign \new_[4664]_  = ~\new_[4671]_  | ~\new_[4668]_  | ~\new_[4666]_  | ~\new_[4665]_ ;
  assign \new_[4665]_  = ~\new_[2955]_  & ~\new_[2702]_ ;
  assign \new_[4666]_  = ~\new_[4667]_ ;
  assign \new_[4667]_  = ~\new_[2889]_  | ~\new_[2891]_  | ~\new_[2890]_ ;
  assign \new_[4668]_  = ~\new_[4669]_  & ~\new_[4670]_ ;
  assign \new_[4669]_  = ~\new_[2701]_  | ~\new_[2947]_ ;
  assign \new_[4670]_  = ~\new_[2948]_ ;
  assign \new_[4671]_  = ~\new_[2608]_  & ~\new_[2305]_ ;
  assign \new_[4672]_  = ~\new_[4673]_ ;
  assign \new_[4673]_  = \new_[4674]_  ? \new_[4678]_  : \new_[4677]_ ;
  assign \new_[4674]_  = \new_[4675]_  & \new_[4676]_ ;
  assign \new_[4675]_  = ~\new_[3566]_  | ~\new_[3987]_ ;
  assign \new_[4676]_  = ~\new_[3914]_  | ~\desIn[63] ;
  assign \new_[4677]_  = ~\new_[4674]_ ;
  assign \new_[4678]_  = ~\new_[2310]_  | ~\new_[1962]_  | ~\new_[1839]_  | ~\new_[1825]_ ;
  assign n765 = \new_[4680]_  ? \new_[4682]_  : \new_[4681]_ ;
  assign \new_[4680]_  = (~\new_[3739]_  & ~\new_[4296]_ ) | (~\new_[1776]_  & ~\new_[3713]_ );
  assign \new_[4681]_  = ~\new_[4680]_ ;
  assign \new_[4682]_  = ~\new_[4683]_  | ~\new_[4686]_ ;
  assign \new_[4683]_  = ~\new_[4684]_  & ~\new_[4685]_ ;
  assign \new_[4684]_  = ~\new_[4782]_  & (~\new_[621]_  | ~\new_[823]_ );
  assign \new_[4685]_  = ~\new_[4894]_  & ~\new_[571]_ ;
  assign \new_[4686]_  = ~\new_[4687]_  & ~\new_[4688]_ ;
  assign \new_[4687]_  = ~\new_[1176]_  & ~\new_[1201]_ ;
  assign \new_[4688]_  = ~\new_[630]_  | ~\new_[4689]_ ;
  assign \new_[4689]_  = ~\new_[4690]_ ;
  assign \new_[4690]_  = ~\new_[1186]_  & ~\new_[1571]_ ;
  assign \new_[4691]_  = ~\new_[4696]_  | ~\new_[4695]_  | ~\new_[4692]_  | ~\new_[4693]_ ;
  assign \new_[4692]_  = ~\new_[1956]_  & ~\new_[1866]_ ;
  assign \new_[4693]_  = ~\new_[4694]_  & ~\new_[2660]_ ;
  assign \new_[4694]_  = ~\new_[4179]_  & (~\new_[3261]_  | ~\new_[3216]_ );
  assign \new_[4695]_  = ~\new_[2126]_  & ~\new_[2125]_ ;
  assign \new_[4696]_  = ~\new_[4697]_  & (~\new_[3022]_  | ~\new_[4256]_ );
  assign \new_[4697]_  = ~\new_[4238]_  & (~\new_[3423]_  | ~\new_[3314]_ );
  assign \new_[4698]_  = \new_[4284]_  & \new_[4288]_ ;
  assign \new_[4699]_  = ~\new_[4700]_  | ~\new_[4708]_ ;
  assign \new_[4700]_  = ~\new_[4701]_  | ~\new_[4706]_ ;
  assign \new_[4701]_  = ~\new_[4702]_  | ~\new_[4704]_ ;
  assign \new_[4702]_  = ~\new_[1796]_  | ~\new_[4707]_  | ~\new_[1846]_ ;
  assign \new_[4703]_  = ~\new_[2106]_  | ~\new_[2324]_ ;
  assign \new_[4704]_  = ~n1055;
  assign n1055 = \new_[3672]_  ? \new_[3914]_  : \desIn[57] ;
  assign \new_[4706]_  = ~n1055 | ~\new_[1796]_  | ~\new_[4707]_  | ~\new_[1846]_ ;
  assign \new_[4707]_  = ~\new_[4703]_ ;
  assign \new_[4708]_  = ~\new_[4610]_  | ~\new_[4609]_ ;
  assign \new_[4709]_  = \new_[4217]_  & \key3[7] ;
  assign \new_[4710]_  = ~\new_[4711]_ ;
  assign \new_[4711]_  = \new_[4712]_  ? \new_[4714]_  : \new_[4713]_ ;
  assign \new_[4712]_  = ~\new_[4713]_ ;
  assign \new_[4713]_  = ~\new_[3578]_  | (~\new_[3461]_  & ~\new_[3837]_ );
  assign \new_[4714]_  = ~\new_[2124]_  | ~\new_[1987]_  | ~\new_[1887]_  | ~\new_[1832]_ ;
  assign \new_[4715]_  = ~\new_[4717]_  | ~\new_[4716]_ ;
  assign \new_[4716]_  = ~\new_[4709]_  & (~\new_[4072]_  | ~\key1[7] );
  assign \new_[4717]_  = ~\new_[4028]_  & (~\new_[4059]_  | ~\key2[7] );
  assign \new_[4718]_  = ~\new_[4813]_ ;
  assign \new_[4719]_  = ~\new_[4720]_ ;
  assign \new_[4720]_  = ~\new_[1655]_  | ~\new_[4901]_ ;
  assign \new_[4721]_  = ~\new_[5042]_  & ~\new_[4722]_ ;
  assign \new_[4722]_  = ~\new_[4723]_  | ~\new_[4724]_ ;
  assign \new_[4723]_  = \new_[4614]_  & \new_[4626]_ ;
  assign \new_[4724]_  = \new_[1641]_  & \new_[4618]_ ;
  assign \new_[4725]_  = ~\new_[4723]_  | ~\new_[4724]_ ;
  assign \new_[4726]_  = ~\new_[1774]_  | ~\new_[3739]_ ;
  assign \new_[4727]_  = ~\new_[3713]_  | ~\desIn[28] ;
  assign \new_[4728]_  = ~\new_[4734]_  | ~\new_[4731]_  | ~\new_[4733]_  | ~\new_[4729]_ ;
  assign \new_[4729]_  = ~\new_[4730]_  & (~\new_[2562]_  | ~\new_[4116]_ );
  assign \new_[4730]_  = ~\new_[2382]_  | ~\new_[2474]_ ;
  assign \new_[4731]_  = ~\new_[4732]_  & (~\new_[3035]_  | ~\new_[4228]_ );
  assign \new_[4732]_  = ~\new_[2188]_  | ~\new_[2475]_ ;
  assign \new_[4733]_  = ~\new_[1937]_  & ~\new_[1938]_ ;
  assign \new_[4734]_  = ~\new_[2426]_  & ~\new_[2539]_ ;
  assign \new_[4735]_  = ~\new_[4742]_  | ~\new_[4736]_  | ~\new_[4739]_ ;
  assign \new_[4736]_  = ~\new_[4737]_  & ~\new_[4520]_ ;
  assign \new_[4737]_  = ~\new_[4738]_  | ~\new_[4517]_ ;
  assign \new_[4738]_  = ~\new_[2514]_  & (~\new_[2548]_  | ~\new_[4102]_ );
  assign \new_[4739]_  = ~\new_[4740]_ ;
  assign \new_[4740]_  = ~\new_[4519]_  | ~\new_[4522]_  | ~\new_[4741]_  | ~\new_[4523]_ ;
  assign \new_[4741]_  = ~\new_[2236]_ ;
  assign \new_[4742]_  = ~\new_[4743]_  & ~\new_[4636]_ ;
  assign \new_[4743]_  = ~\new_[2040]_  | ~\new_[4639]_ ;
  assign \new_[4744]_  = ~\new_[5133]_  & ~\new_[4745]_ ;
  assign \new_[4745]_  = ~\new_[4746]_  | ~\new_[4747]_ ;
  assign \new_[4746]_  = ~\new_[5294]_ ;
  assign \new_[4747]_  = \new_[5129]_ ;
  assign n895 = \new_[4749]_  ? \new_[4752]_  : \new_[4750]_ ;
  assign \new_[4749]_  = ~\new_[4750]_ ;
  assign \new_[4750]_  = ~\new_[4751]_  | (~\new_[1750]_  & ~\new_[3713]_ );
  assign \new_[4751]_  = \new_[4335]_  | \new_[3739]_ ;
  assign \new_[4752]_  = ~\new_[785]_  | ~\new_[548]_  | ~\new_[565]_ ;
  assign \new_[4753]_  = ~\new_[4754]_  | ~\new_[4757]_ ;
  assign \new_[4754]_  = ~\new_[4755]_  | ~\new_[970]_  | ~\new_[1374]_ ;
  assign \new_[4755]_  = ~\new_[5244]_  | ~\new_[1594]_  | ~\new_[4756]_ ;
  assign \new_[4756]_  = \new_[4860]_ ;
  assign \new_[4757]_  = \new_[4758]_ ;
  assign \new_[4758]_  = ~\new_[4759]_ ;
  assign \new_[4759]_  = ~\new_[1600]_  | ~\new_[1630]_ ;
  assign \new_[4760]_  = ~\new_[4755]_ ;
  assign \new_[4761]_  = ~\new_[1594]_  | ~\new_[4756]_ ;
  assign \new_[4762]_  = ~\new_[4763]_  | ~\new_[4768]_ ;
  assign \new_[4763]_  = ~\new_[4764]_  | ~\new_[4765]_ ;
  assign \new_[4764]_  = ~\new_[4127]_  & (~\new_[4035]_  | ~\key2[5] );
  assign \new_[4765]_  = \new_[4766]_  & \new_[4767]_ ;
  assign \new_[4766]_  = ~\new_[4066]_  | ~\key1[5] ;
  assign \new_[4767]_  = ~\new_[4120]_  | ~\key3[5] ;
  assign \new_[4768]_  = ~\new_[4769]_ ;
  assign \new_[4769]_  = ~\new_[5103]_ ;
  assign n715 = \new_[4771]_  ? \new_[4773]_  : \new_[4772]_ ;
  assign \new_[4771]_  = ~\new_[4772]_ ;
  assign \new_[4772]_  = (~\desIn[44]  | ~\new_[2908]_ ) & (~\new_[1778]_  | ~\new_[2871]_ );
  assign \new_[4773]_  = ~\new_[530]_  | ~\new_[534]_ ;
  assign \new_[4774]_  = ~\new_[4779]_  | ~\new_[4775]_  | ~\new_[4776]_ ;
  assign \new_[4775]_  = ~\new_[582]_  | ~\new_[1178]_ ;
  assign \new_[4776]_  = \new_[4777]_  & \new_[4778]_ ;
  assign \new_[4777]_  = ~\new_[1506]_  | (~\new_[883]_  & ~\new_[873]_ );
  assign \new_[4778]_  = ~\new_[1064]_  & ~\new_[4690]_ ;
  assign \new_[4779]_  = ~\new_[1319]_  | ~\new_[4780]_ ;
  assign \new_[4780]_  = ~\new_[4781]_  | ~\new_[1185]_  | ~\new_[674]_  | ~\new_[775]_ ;
  assign \new_[4781]_  = \new_[1265]_  & \new_[1188]_ ;
  assign \new_[4782]_  = ~\new_[4894]_ ;
  assign \new_[4783]_  = ~\new_[4792]_  & (~\new_[4784]_  | ~\new_[4790]_ );
  assign \new_[4784]_  = \new_[4785]_ ;
  assign \new_[4785]_  = ~\new_[4786]_  | ~\new_[4787]_ ;
  assign \new_[4786]_  = ~\new_[3876]_  | ~\new_[3923]_ ;
  assign \new_[4787]_  = ~\new_[4788]_ ;
  assign \new_[4788]_  = ~\new_[4030]_ ;
  assign \new_[4789]_  = ~\new_[5105]_ ;
  assign \new_[4790]_  = ~\new_[4791]_ ;
  assign \new_[4791]_  = ~\new_[4863]_ ;
  assign \new_[4792]_  = ~\new_[4284]_  | ~\new_[4280]_ ;
  assign \new_[4793]_  = ~\new_[4792]_ ;
  assign \new_[4794]_  = \new_[5294]_ ;
  assign \new_[4795]_  = ~\new_[5133]_ ;
  assign \new_[4796]_  = ~\new_[5128]_ ;
  assign \new_[4797]_  = ~\new_[4800]_  | ~\new_[4798]_  | ~\new_[4799]_ ;
  assign \new_[4798]_  = ~\new_[1171]_  | (~\new_[1092]_  & ~\new_[817]_ );
  assign \new_[4799]_  = ~\new_[911]_  | ~\new_[1310]_ ;
  assign \new_[4800]_  = ~\new_[4801]_  & ~\new_[4805]_ ;
  assign \new_[4801]_  = \new_[4760]_  & \new_[4802]_ ;
  assign \new_[4802]_  = ~\new_[4803]_ ;
  assign \new_[4803]_  = ~\new_[4804]_ ;
  assign \new_[4804]_  = ~\new_[1684]_  | ~\new_[1702]_ ;
  assign \new_[4805]_  = ~\new_[4802]_  & (~\new_[1194]_  | ~\new_[1200]_ );
  assign \new_[4806]_  = ~\new_[4801]_ ;
  assign \new_[4807]_  = ~\new_[4802]_ ;
  assign \new_[4808]_  = ~\new_[4809]_  | ~\new_[4810]_ ;
  assign \new_[4809]_  = ~\new_[3891]_  | ~\new_[3848]_ ;
  assign \new_[4810]_  = \new_[4865]_ ;
  assign \new_[4811]_  = ~\new_[4414]_  | ~\new_[4286]_ ;
  assign \new_[4812]_  = ~\new_[4321]_  | ~\new_[4278]_  | ~\new_[4289]_ ;
  assign \new_[4813]_  = ~\new_[5104]_ ;
  assign \new_[4814]_  = ~\new_[4821]_  | ~\new_[4819]_  | ~\new_[4815]_  | ~\new_[4818]_ ;
  assign \new_[4815]_  = ~\new_[4816]_  & (~\new_[3111]_  | ~\new_[4232]_ );
  assign \new_[4816]_  = ~\new_[2356]_  | ~\new_[4817]_ ;
  assign \new_[4817]_  = ~\new_[2983]_ ;
  assign \new_[4818]_  = ~\new_[2373]_  & ~\new_[2129]_ ;
  assign \new_[4819]_  = ~\new_[4820]_  & (~\new_[3134]_  | ~\new_[4209]_ );
  assign \new_[4820]_  = ~\new_[2882]_  | ~\new_[2875]_ ;
  assign \new_[4821]_  = ~\new_[4822]_  & ~\new_[2699]_ ;
  assign \new_[4822]_  = ~\new_[2923]_  | ~\new_[2922]_ ;
  assign \new_[4823]_  = ~\new_[4824]_  & ~\new_[5091]_ ;
  assign \new_[4824]_  = ~\new_[4827]_  | ~\new_[4826]_  | ~\new_[4825]_ ;
  assign \new_[4825]_  = ~\new_[2149]_ ;
  assign \new_[4826]_  = ~\new_[2094]_  & (~\new_[3234]_  | ~\new_[4208]_ );
  assign \new_[4827]_  = ~\new_[4828]_  & ~\new_[2134]_ ;
  assign \new_[4828]_  = ~\new_[2897]_ ;
  assign \new_[4829]_  = \new_[4662]_ ;
  assign \new_[4830]_  = \new_[4662]_ ;
  assign \new_[4831]_  = ~\new_[1648]_  | ~\new_[1668]_ ;
  assign \new_[4832]_  = ~\new_[1648]_  | ~\new_[1668]_ ;
  assign \new_[4833]_  = \new_[4464]_  ? \new_[4466]_  : n1015;
  assign n790 = \new_[4539]_  ? \new_[4972]_  : \new_[4540]_ ;
  assign n830 = \new_[4539]_  ? \new_[4972]_  : \new_[4540]_ ;
  assign \new_[4836]_  = ~\new_[4928]_  | ~\new_[3290]_ ;
  assign \new_[4837]_  = ~\new_[4928]_  | ~\new_[3290]_ ;
  assign \new_[4838]_  = ~\new_[5076]_  | ~\new_[5072]_ ;
  assign \new_[4839]_  = ~\new_[4906]_  & ~\new_[4907]_ ;
  assign \new_[4840]_  = ~\new_[4841]_ ;
  assign \new_[4841]_  = ~\new_[4842]_ ;
  assign \new_[4842]_  = ~\new_[1541]_ ;
  assign \new_[4843]_  = ~decrypt | ~\new_[4970]_  | ~\new_[4844]_ ;
  assign \new_[4844]_  = ~\roundSel[4] ;
  assign \new_[4845]_  = ~\new_[4850]_  | ~\new_[4847]_  | ~\new_[4846]_ ;
  assign \new_[4846]_  = ~\new_[729]_  & (~\new_[1019]_  | ~\new_[1321]_ );
  assign \new_[4847]_  = ~\new_[4848]_  | ~\new_[4849]_ ;
  assign \new_[4848]_  = ~\new_[736]_  | ~\new_[656]_ ;
  assign \new_[4849]_  = ~\new_[4961]_ ;
  assign \new_[4850]_  = ~\new_[4961]_  | ~\new_[586]_ ;
  assign \new_[4851]_  = ~\new_[4849]_  | ~\new_[4848]_ ;
  assign \new_[4852]_  = ~\new_[4961]_  | ~\new_[586]_ ;
  assign \new_[4853]_  = \new_[4854]_  | \new_[5169]_ ;
  assign \new_[4854]_  = ~\new_[2404]_  | ~\new_[2239]_  | ~\new_[2240]_  | ~\new_[2241]_ ;
  assign \new_[4855]_  = ~\new_[2039]_  | ~\new_[4548]_ ;
  assign \new_[4856]_  = ~\new_[2049]_  | ~\new_[2048]_ ;
  assign \new_[4857]_  = ~\new_[5244]_  & ~\new_[5283]_ ;
  assign \new_[4858]_  = ~\new_[1655]_  | ~\new_[4901]_ ;
  assign \new_[4859]_  = n1150 ? \new_[4823]_  : \new_[5075]_ ;
  assign \new_[4860]_  = n1015 ? \new_[4466]_  : \new_[4464]_ ;
  assign \new_[4861]_  = ~\new_[4860]_ ;
  assign \new_[4862]_  = ~\new_[4859]_ ;
  assign \new_[4863]_  = ~\new_[3855]_  | ~\new_[4866]_ ;
  assign \new_[4864]_  = ~\new_[4865]_ ;
  assign \new_[4865]_  = \new_[5104]_ ;
  assign \new_[4866]_  = ~\new_[4869]_  | ~\new_[4867]_  | ~\new_[4868]_ ;
  assign \new_[4867]_  = (~\key3[13]  | ~\new_[4144]_ ) & (~\new_[4227]_  | ~\key3[13] );
  assign \new_[4868]_  = ~\new_[4010]_  | ~\key2[13] ;
  assign \new_[4869]_  = ~\new_[4084]_  | ~\key1[13] ;
  assign \new_[4870]_  = ~\new_[5045]_  | ~\new_[5188]_  | ~\new_[4871]_  | ~\new_[4875]_ ;
  assign \new_[4871]_  = ~\new_[4872]_  | ~\new_[4873]_ ;
  assign \new_[4872]_  = ~\new_[604]_  | ~\new_[894]_ ;
  assign \new_[4873]_  = ~\new_[4874]_ ;
  assign \new_[4874]_  = ~\new_[1601]_  | ~\new_[1631]_ ;
  assign \new_[4875]_  = ~\new_[4874]_  | ~\new_[579]_ ;
  assign n780 = \new_[4877]_  ? \new_[4879]_  : \new_[4878]_ ;
  assign \new_[4877]_  = ~\new_[4726]_  | ~\new_[4727]_ ;
  assign \new_[4878]_  = ~\new_[4877]_ ;
  assign \new_[4879]_  = ~\new_[535]_  | ~\new_[541]_ ;
  assign \new_[4880]_  = ~\new_[4890]_  | ~\new_[4887]_  | ~\new_[4881]_  | ~\new_[4884]_ ;
  assign \new_[4881]_  = ~\new_[5084]_ ;
  assign \new_[4882]_  = ~\new_[3227]_  & (~\new_[3690]_  | ~\new_[3831]_ );
  assign \new_[4883]_  = ~\new_[1851]_  & ~\new_[1727]_ ;
  assign \new_[4884]_  = \new_[4885]_ ;
  assign \new_[4885]_  = ~\new_[4886]_ ;
  assign \new_[4886]_  = \new_[2792]_  ? \new_[4501]_  : n1130;
  assign \new_[4887]_  = ~\new_[4888]_ ;
  assign \new_[4888]_  = ~\new_[4889]_ ;
  assign \new_[4889]_  = ~\new_[4605]_  | ~\new_[4606]_ ;
  assign \new_[4890]_  = ~\new_[4891]_ ;
  assign \new_[4891]_  = ~\new_[4892]_ ;
  assign \new_[4892]_  = \new_[4620]_  ? \new_[5011]_  : n1245;
  assign \new_[4893]_  = ~\new_[4890]_ ;
  assign \new_[4894]_  = n1145 ^ \new_[4895]_ ;
  assign \new_[4895]_  = ~\new_[1838]_  | ~\new_[1741]_  | ~\new_[4896]_ ;
  assign \new_[4896]_  = \new_[1892]_  & \new_[1891]_ ;
  assign \new_[4897]_  = ~\new_[1963]_  | ~\new_[4899]_  | ~\new_[1791]_ ;
  assign \new_[4898]_  = ~\new_[1878]_  | ~\new_[2343]_ ;
  assign \new_[4899]_  = ~\new_[4898]_ ;
  assign n1145 = ~\new_[3328]_  | ~\new_[3692]_ ;
  assign \new_[4901]_  = ~\new_[4905]_  | (~\new_[4902]_  & ~\new_[4903]_ );
  assign \new_[4902]_  = ~\new_[4559]_  | ~\new_[4557]_  | ~\new_[4555]_  | ~\new_[2307]_ ;
  assign \new_[4903]_  = ~\new_[4904]_  | ~\new_[4554]_ ;
  assign \new_[4904]_  = \new_[2387]_  & \new_[2479]_ ;
  assign \new_[4905]_  = (~\new_[3809]_  | ~\new_[3740]_ ) & (~\new_[3837]_  | ~\desIn[33] );
  assign \new_[4906]_  = ~\new_[2479]_  | ~\new_[2307]_  | ~\new_[2387]_ ;
  assign \new_[4907]_  = ~\new_[4559]_  | ~\new_[4557]_  | ~\new_[4555]_  | ~\new_[4554]_ ;
  assign \new_[4908]_  = ~\new_[2478]_ ;
  assign \new_[4909]_  = ~\new_[2465]_  | ~\new_[2392]_ ;
  assign \new_[4910]_  = ~\new_[4914]_  & (~\new_[4911]_  | ~\key2[9] );
  assign \new_[4911]_  = ~\new_[4912]_  | ~\new_[4913]_ ;
  assign \new_[4912]_  = ~\new_[5224]_ ;
  assign \new_[4913]_  = ~\new_[5228]_ ;
  assign \new_[4914]_  = ~\new_[4351]_  & ~\new_[4171]_ ;
  assign n825 = \new_[4916]_  ? \new_[4918]_  : \new_[4917]_ ;
  assign \new_[4916]_  = ~\new_[4917]_ ;
  assign \new_[4917]_  = (~\new_[2898]_  | ~\new_[1770]_ ) & (~\new_[2639]_  | ~\desIn[34] );
  assign \new_[4918]_  = ~\new_[4921]_  | ~\new_[4920]_  | ~\new_[4919]_ ;
  assign \new_[4919]_  = ~\new_[4797]_  | ~\new_[1524]_ ;
  assign \new_[4920]_  = ~\new_[567]_  | ~\new_[1523]_ ;
  assign \new_[4921]_  = ~\new_[4922]_  & (~\new_[1150]_  | ~\new_[1172]_ );
  assign \new_[4922]_  = \new_[830]_  & \new_[1418]_ ;
  assign n835 = \new_[4924]_  ? \new_[4926]_  : \new_[4925]_ ;
  assign \new_[4924]_  = ~\new_[4925]_ ;
  assign \new_[4925]_  = (~\new_[2871]_  | ~\new_[1766]_ ) & (~\new_[2908]_  | ~\desIn[46] );
  assign \new_[4926]_  = ~\new_[4927]_  | ~\new_[4951]_  | ~\new_[5037]_ ;
  assign \new_[4927]_  = ~\new_[610]_ ;
  assign \new_[4928]_  = ~\new_[4929]_  | ~\new_[4936]_ ;
  assign \new_[4929]_  = ~\new_[4930]_ ;
  assign \new_[4930]_  = ~\new_[4935]_  | ~\new_[4933]_  | ~\new_[4931]_  | ~\new_[4932]_ ;
  assign \new_[4931]_  = ~\new_[2613]_  & ~\new_[2614]_ ;
  assign \new_[4932]_  = \new_[3176]_  & \new_[2916]_ ;
  assign \new_[4933]_  = ~\new_[4934]_  & (~\new_[2971]_  | ~\new_[4248]_ );
  assign \new_[4934]_  = \new_[4698]_  & \new_[3369]_ ;
  assign \new_[4935]_  = ~\new_[2974]_  & ~\new_[2680]_ ;
  assign \new_[4936]_  = ~\new_[4937]_  & ~\new_[4938]_ ;
  assign \new_[4937]_  = ~\new_[2242]_  | ~\new_[2531]_ ;
  assign \new_[4938]_  = ~\new_[2679]_  | ~\new_[2121]_  | ~\new_[2647]_ ;
  assign \new_[4939]_  = ~\new_[2531]_  | ~\new_[2242]_ ;
  assign \new_[4940]_  = \new_[2853]_  | \new_[4942]_ ;
  assign n1115 = ~\new_[3466]_  | ~\new_[3745]_ ;
  assign \new_[4942]_  = ~\new_[4949]_  | ~\new_[4948]_  | ~\new_[4944]_  | ~\new_[4943]_ ;
  assign \new_[4943]_  = ~\new_[2291]_  & ~\new_[2105]_ ;
  assign \new_[4944]_  = ~\new_[2138]_  & ~\new_[4945]_ ;
  assign \new_[4945]_  = ~\new_[4946]_  | ~\new_[4947]_ ;
  assign \new_[4946]_  = ~\new_[2932]_ ;
  assign \new_[4947]_  = ~\new_[2633]_  | ~\new_[4222]_ ;
  assign \new_[4948]_  = ~\new_[2822]_  | ~\new_[4126]_ ;
  assign \new_[4949]_  = ~\new_[2405]_  & ~\new_[2072]_ ;
  assign \new_[4950]_  = \new_[4310]_  | \new_[2872]_ ;
  assign \new_[4951]_  = ~\new_[4952]_  | ~\new_[4961]_ ;
  assign \new_[4952]_  = ~\new_[4960]_  | ~\new_[4953]_  | ~\new_[4958]_ ;
  assign \new_[4953]_  = ~\new_[4954]_  & ~\new_[4957]_ ;
  assign \new_[4954]_  = ~\new_[4955]_  | ~\new_[4956]_ ;
  assign \new_[4955]_  = ~\new_[1475]_  | ~\new_[5285]_  | ~\new_[1618]_  | ~\new_[1522]_ ;
  assign \new_[4956]_  = ~\new_[1445]_  | ~\new_[1613]_  | ~\new_[5042]_ ;
  assign \new_[4957]_  = ~\new_[965]_  | ~\new_[1083]_  | ~\new_[4725]_ ;
  assign \new_[4958]_  = ~\new_[4959]_  | ~\new_[1168]_  | ~\new_[1618]_ ;
  assign \new_[4959]_  = ~\new_[4613]_ ;
  assign \new_[4960]_  = \new_[1612]_  | \new_[1115]_ ;
  assign \new_[4961]_  = \new_[4962]_ ;
  assign \new_[4962]_  = ~\new_[1529]_  | ~\new_[1528]_ ;
  assign \new_[4963]_  = ~\new_[4964]_  | ~\new_[4213]_ ;
  assign \new_[4964]_  = ~\new_[4965]_ ;
  assign \new_[4965]_  = ~\new_[4966]_ ;
  assign \new_[4966]_  = ~decrypt | ~\new_[4635]_  | ~\new_[4967]_ ;
  assign \new_[4967]_  = ~\roundSel[4] ;
  assign \new_[4968]_  = ~\new_[4969]_ ;
  assign \new_[4969]_  = ~\new_[4971]_  | ~\new_[4970]_  | ~\new_[4967]_ ;
  assign \new_[4970]_  = ~\roundSel[5] ;
  assign \new_[4971]_  = ~decrypt;
  assign \new_[4972]_  = ~\new_[566]_  | ~\new_[4978]_  | ~\new_[4973]_  | ~\new_[4976]_ ;
  assign \new_[4973]_  = ~\new_[4974]_  | ~\new_[1524]_ ;
  assign \new_[4974]_  = ~\new_[1091]_  | ~\new_[793]_  | ~\new_[706]_  | ~\new_[709]_ ;
  assign \new_[4975]_  = ~\new_[1650]_  | ~\new_[1647]_ ;
  assign \new_[4976]_  = ~\new_[4977]_  & ~\new_[758]_ ;
  assign \new_[4977]_  = ~\new_[750]_  | ~\new_[651]_ ;
  assign \new_[4978]_  = ~\new_[722]_  | ~\new_[1310]_ ;
  assign n905 = \new_[4980]_  ? \new_[4982]_  : \new_[4981]_ ;
  assign \new_[4980]_  = (~\new_[1747]_  & ~\new_[3713]_ ) | (~\new_[3739]_  & ~\new_[4359]_ );
  assign \new_[4981]_  = ~\new_[4980]_ ;
  assign \new_[4982]_  = ~\new_[4985]_  | ~\new_[4983]_  | ~\new_[4984]_ ;
  assign \new_[4983]_  = ~\new_[1317]_  | ~\new_[564]_ ;
  assign \new_[4984]_  = ~\new_[588]_  & (~\new_[643]_  | ~\new_[1520]_ );
  assign \new_[4985]_  = ~\new_[626]_  | ~\new_[4417]_ ;
  assign \new_[4986]_  = ~\new_[4987]_  | ~\new_[4988]_ ;
  assign \new_[4987]_  = (~\desIn[10]  | ~\new_[2908]_ ) & (~\new_[1763]_  | ~\new_[2871]_ );
  assign \new_[4988]_  = ~\new_[976]_  | ~\new_[557]_  | ~\new_[555]_  | ~\new_[629]_ ;
  assign \new_[4989]_  = ~\new_[4988]_ ;
  assign \new_[4990]_  = ~n1205;
  assign n1205 = ~\new_[3699]_  | (~\new_[3505]_  & ~\new_[3837]_ );
  assign \new_[4992]_  = ~\new_[1842]_  & ~\new_[1726]_ ;
  assign \new_[4993]_  = ~\new_[5005]_  | ~\new_[4994]_  | ~\new_[4995]_ ;
  assign \new_[4994]_  = ~\new_[559]_  | ~\new_[1318]_ ;
  assign \new_[4995]_  = ~\new_[4996]_ ;
  assign \new_[4996]_  = ~\new_[4997]_  | ~\new_[5003]_ ;
  assign \new_[4997]_  = ~\new_[4998]_  | ~\new_[4999]_ ;
  assign \new_[4998]_  = ~\new_[798]_  | ~\new_[1102]_ ;
  assign \new_[4999]_  = ~\new_[5000]_ ;
  assign \new_[5000]_  = \new_[5001]_ ;
  assign \new_[5001]_  = ~\new_[5002]_ ;
  assign \new_[5002]_  = n1000 ? \new_[1688]_  : \new_[2596]_ ;
  assign \new_[5003]_  = ~\new_[5004]_  | ~\new_[730]_  | ~\new_[1412]_ ;
  assign \new_[5004]_  = ~\new_[4999]_ ;
  assign \new_[5005]_  = ~\new_[1424]_  | (~\new_[669]_  & ~\new_[662]_ );
  assign n880 = \new_[5007]_  ? \new_[5010]_  : \new_[5008]_ ;
  assign \new_[5007]_  = ~\new_[5008]_ ;
  assign \new_[5008]_  = ~\new_[5009]_  | (~\new_[1749]_  & ~\new_[2639]_ );
  assign \new_[5009]_  = \new_[4362]_  | \new_[3739]_ ;
  assign \new_[5010]_  = ~\new_[4489]_  | ~\new_[4487]_  | ~\new_[4484]_  | ~\new_[4486]_ ;
  assign \new_[5011]_  = ~\new_[5018]_  | ~\new_[5016]_  | ~\new_[5012]_  | ~\new_[5015]_ ;
  assign \new_[5012]_  = ~\new_[2533]_  & ~\new_[5013]_ ;
  assign \new_[5013]_  = ~\new_[5014]_  | ~\new_[2347]_ ;
  assign \new_[5014]_  = ~\new_[2751]_ ;
  assign \new_[5015]_  = ~\new_[2370]_  & ~\new_[2122]_ ;
  assign \new_[5016]_  = ~\new_[5017]_  & (~\new_[3120]_  | ~\new_[4209]_ );
  assign \new_[5017]_  = ~\new_[2623]_  | ~\new_[2873]_ ;
  assign \new_[5018]_  = ~\new_[5019]_  & (~\new_[2769]_  | ~\new_[4233]_ );
  assign \new_[5019]_  = ~\new_[2918]_  | ~\new_[2638]_ ;
  assign \new_[5020]_  = ~\new_[5026]_  | ~\new_[5024]_  | ~\new_[5021]_  | ~\new_[5023]_ ;
  assign \new_[5021]_  = ~\new_[5022]_ ;
  assign \new_[5022]_  = ~\new_[849]_  | (~\new_[812]_  & ~\new_[4391]_ );
  assign \new_[5023]_  = ~\new_[1307]_  | (~\new_[591]_  & ~\new_[920]_ );
  assign \new_[5024]_  = ~\new_[5025]_ ;
  assign \new_[5025]_  = ~\new_[1308]_  & (~\new_[715]_  | ~\new_[1222]_ );
  assign \new_[5026]_  = ~\new_[592]_  | ~\new_[4535]_ ;
  assign \new_[5027]_  = ~\new_[5023]_  | ~\new_[5026]_ ;
  assign \new_[5028]_  = ~\new_[1308]_  & (~\new_[1222]_  | ~\new_[715]_ );
  assign n870 = \new_[5030]_  ? \new_[5032]_  : \new_[5031]_ ;
  assign \new_[5030]_  = ~\new_[5031]_ ;
  assign \new_[5031]_  = (~\new_[2871]_  | ~\new_[1762]_ ) & (~\new_[2908]_  | ~\desIn[56] );
  assign \new_[5032]_  = ~\new_[5035]_  | ~\new_[5033]_  | ~\new_[5034]_ ;
  assign \new_[5033]_  = ~\new_[1308]_  | ~\new_[574]_ ;
  assign \new_[5034]_  = ~\new_[4535]_  | ~\new_[581]_ ;
  assign \new_[5035]_  = ~\new_[5036]_  & (~\new_[5161]_  | ~\new_[1108]_ );
  assign \new_[5036]_  = \new_[4390]_  & \new_[848]_ ;
  assign \new_[5037]_  = ~\new_[5040]_  & (~\new_[5038]_  | ~\new_[5039]_ );
  assign \new_[5038]_  = \new_[1289]_  | \new_[1002]_ ;
  assign \new_[5039]_  = ~\new_[5286]_  & ~\new_[4962]_ ;
  assign \new_[5040]_  = ~\new_[5042]_  & (~\new_[982]_  | ~\new_[1461]_ );
  assign \new_[5041]_  = ~\new_[5042]_ ;
  assign \new_[5042]_  = \new_[5043]_ ;
  assign \new_[5043]_  = ~\new_[1627]_  | ~\new_[1649]_ ;
  assign \new_[5044]_  = ~\new_[1627]_  | ~\new_[1649]_ ;
  assign \new_[5045]_  = ~\new_[5048]_  | ~\new_[5116]_  | ~\new_[5046]_  | ~\new_[5047]_ ;
  assign \new_[5046]_  = ~\new_[1518]_ ;
  assign \new_[5047]_  = ~\new_[5127]_ ;
  assign \new_[5048]_  = ~\new_[5049]_ ;
  assign \new_[5049]_  = \new_[5050]_ ;
  assign \new_[5050]_  = ~\new_[5293]_ ;
  assign \new_[5051]_  = ~\new_[1722]_  | ~n985;
  assign \new_[5052]_  = ~\new_[4570]_  | ~\new_[1735]_ ;
  assign \new_[5053]_  = ~\new_[5048]_ ;
  assign \new_[5054]_  = ~\new_[5050]_ ;
  assign \new_[5055]_  = ~\new_[5047]_ ;
  assign \new_[5056]_  = ~\new_[3691]_  | ~\new_[3831]_ ;
  assign \new_[5057]_  = ~\new_[3463]_ ;
  assign \new_[5058]_  = ~\new_[1880]_  & ~\new_[4856]_ ;
  assign \new_[5059]_  = ~\new_[4552]_  & ~\new_[1879]_ ;
  assign \new_[5060]_  = ~\new_[5066]_  | ~\new_[5061]_  | ~\new_[5064]_  | ~\new_[5065]_ ;
  assign \new_[5061]_  = ~\new_[5062]_  & (~\new_[3016]_  | ~\new_[4232]_ );
  assign \new_[5062]_  = ~\new_[5063]_  & (~\new_[3717]_  | ~\new_[3310]_ );
  assign \new_[5063]_  = ~\new_[4279]_  | ~\new_[4283]_ ;
  assign \new_[5064]_  = ~\new_[1934]_  & ~\new_[1873]_ ;
  assign \new_[5065]_  = ~\new_[2135]_  & ~\new_[2090]_ ;
  assign \new_[5066]_  = ~\new_[5067]_  & ~\new_[2473]_ ;
  assign \new_[5067]_  = ~\new_[4192]_  & (~\new_[3735]_  | ~\new_[4382]_ );
  assign \new_[5068]_  = ~\new_[5063]_ ;
  assign \new_[5069]_  = ~\new_[5070]_  | ~\new_[5072]_ ;
  assign \new_[5070]_  = ~\new_[2856]_  | ~\new_[5071]_ ;
  assign \new_[5071]_  = ~\new_[4547]_  | ~\new_[4543]_  | ~\new_[4541]_  | ~\new_[4545]_ ;
  assign \new_[5072]_  = ~n1150 | ~\new_[4543]_  | ~\new_[5073]_  | ~\new_[4541]_ ;
  assign \new_[5073]_  = \new_[4547]_  & \new_[4545]_ ;
  assign n1150 = ~\new_[5075]_ ;
  assign \new_[5075]_  = ~\new_[3574]_  & (~\new_[3812]_  | ~\new_[3831]_ );
  assign \new_[5076]_  = ~\new_[2856]_  | ~\new_[5071]_ ;
  assign \new_[5077]_  = ~\new_[5133]_ ;
  assign \new_[5078]_  = \new_[5293]_  & \new_[5129]_ ;
  assign \new_[5079]_  = ~\new_[4607]_  | ~\new_[1322]_  | ~\new_[4643]_  | ~\new_[1420]_ ;
  assign \new_[5080]_  = ~\new_[1180]_  | ~\new_[1467]_ ;
  assign \new_[5081]_  = ~\new_[5082]_ ;
  assign \new_[5082]_  = ~\new_[5083]_ ;
  assign \new_[5083]_  = ~\new_[5084]_ ;
  assign \new_[5084]_  = ~\new_[5085]_ ;
  assign \new_[5085]_  = \new_[4882]_  ? \new_[4883]_  : n1155;
  assign \new_[5086]_  = ~\new_[5087]_  | ~\new_[5089]_ ;
  assign \new_[5087]_  = ~\new_[5088]_  & (~\new_[4082]_  | ~\key1[1] );
  assign \new_[5088]_  = ~\new_[4294]_  & (~\new_[4103]_  | ~\new_[4234]_ );
  assign \new_[5089]_  = ~\new_[5090]_  & ~\new_[4017]_ ;
  assign \new_[5090]_  = ~\new_[4258]_  & ~\new_[4341]_ ;
  assign \new_[5091]_  = ~\new_[5095]_  | ~\new_[5094]_  | ~\new_[5092]_  | ~\new_[5093]_ ;
  assign \new_[5092]_  = ~\new_[2714]_  & ~\new_[2095]_ ;
  assign \new_[5093]_  = ~\new_[2711]_  & (~\new_[3047]_  | ~\new_[4122]_ );
  assign \new_[5094]_  = ~\new_[2393]_  & ~\new_[2075]_ ;
  assign \new_[5095]_  = ~\new_[5096]_  | ~\new_[5097]_ ;
  assign \new_[5096]_  = ~\new_[3327]_  | ~\new_[3446]_ ;
  assign \new_[5097]_  = ~\new_[5098]_ ;
  assign \new_[5098]_  = ~\new_[4279]_  | ~\new_[4288]_ ;
  assign \new_[5099]_  = ~\new_[5098]_ ;
  assign \new_[5100]_  = ~\new_[5101]_  | ~\new_[5106]_ ;
  assign \new_[5101]_  = ~\new_[5102]_ ;
  assign \new_[5102]_  = ~\new_[5103]_ ;
  assign \new_[5103]_  = ~\new_[5104]_ ;
  assign \new_[5104]_  = ~\new_[5105]_ ;
  assign \new_[5105]_  = ~\new_[4811]_  | ~\new_[4812]_ ;
  assign \new_[5106]_  = ~\new_[5109]_  | ~\new_[5107]_  | ~\new_[5108]_ ;
  assign \new_[5107]_  = (~\key3[26]  | ~\new_[4144]_ ) & (~\new_[4260]_  | ~\key3[26] );
  assign \new_[5108]_  = ~\new_[4034]_  | ~\key2[26] ;
  assign \new_[5109]_  = ~\new_[4071]_  | ~\key1[26] ;
  assign \new_[5110]_  = ~\new_[5111]_ ;
  assign \new_[5111]_  = ~\new_[5112]_ ;
  assign \new_[5112]_  = ~\new_[5114]_  | ~\new_[5113]_ ;
  assign \new_[5113]_  = ~\new_[4992]_  | ~n1205;
  assign \new_[5114]_  = ~\new_[4990]_  | (~\new_[1726]_  & ~\new_[1842]_ );
  assign \new_[5115]_  = ~\new_[5078]_  | ~\new_[5077]_ ;
  assign \new_[5116]_  = ~\new_[5110]_ ;
  assign \new_[5117]_  = ~\new_[5125]_  | ~\new_[5124]_  | ~\new_[5118]_  | ~\new_[5122]_ ;
  assign \new_[5118]_  = ~\new_[5121]_  | ~\new_[5119]_  | ~\new_[5083]_ ;
  assign \new_[5119]_  = ~\new_[5120]_ ;
  assign \new_[5120]_  = ~\new_[1268]_  & (~\new_[1428]_  | ~\new_[1069]_ );
  assign \new_[5121]_  = \new_[4674]_  ? \new_[1654]_  : \new_[4677]_ ;
  assign \new_[5122]_  = ~\new_[5123]_  | ~\new_[5082]_ ;
  assign \new_[5123]_  = ~\new_[5080]_  | ~\new_[5079]_ ;
  assign \new_[5124]_  = ~\new_[865]_  | ~\new_[5081]_ ;
  assign \new_[5125]_  = ~\new_[664]_  | ~\new_[5121]_ ;
  assign \new_[5126]_  = ~\new_[5121]_ ;
  assign \new_[5127]_  = ~\new_[5128]_  | ~\new_[5130]_ ;
  assign \new_[5128]_  = ~\new_[5129]_ ;
  assign \new_[5129]_  = ~\new_[4940]_  | ~\new_[1715]_ ;
  assign \new_[5130]_  = ~\new_[5131]_  | ~\new_[5132]_ ;
  assign \new_[5131]_  = ~n1145 | ~\new_[1963]_  | ~\new_[4899]_  | ~\new_[1791]_ ;
  assign \new_[5132]_  = ~\new_[4897]_  | ~\new_[2852]_ ;
  assign \new_[5133]_  = ~\new_[5132]_  | ~\new_[5131]_ ;
  assign \new_[5134]_  = ~\new_[5141]_  | ~\new_[5135]_  | ~\new_[5139]_ ;
  assign \new_[5135]_  = ~\new_[5136]_  & ~\new_[1849]_ ;
  assign \new_[5136]_  = ~\new_[4633]_  | ~\new_[5137]_ ;
  assign \new_[5137]_  = ~\new_[5138]_  | ~\new_[4074]_ ;
  assign \new_[5138]_  = ~\new_[3165]_  | ~\new_[3524]_ ;
  assign \new_[5139]_  = ~\new_[4631]_  & ~\new_[5140]_ ;
  assign \new_[5140]_  = \new_[2456]_  | \new_[4634]_ ;
  assign \new_[5141]_  = ~\new_[5142]_ ;
  assign \new_[5142]_  = ~\new_[2870]_  | ~\new_[2057]_  | ~\new_[1983]_  | ~\new_[2056]_ ;
  assign \new_[5143]_  = ~\new_[5148]_  | ~\new_[5146]_  | ~\new_[5144]_  | ~\new_[5145]_ ;
  assign \new_[5144]_  = ~\new_[1893]_  & ~\new_[1894]_ ;
  assign \new_[5145]_  = ~\new_[4908]_  & (~\new_[2790]_  | ~\new_[4121]_ );
  assign \new_[5146]_  = ~\new_[5147]_  & ~\new_[2246]_ ;
  assign \new_[5147]_  = ~\new_[2391]_  | ~\new_[2384]_ ;
  assign \new_[5148]_  = ~\new_[4909]_  & (~\new_[3036]_  | ~\new_[4166]_ );
  assign \new_[5149]_  = ~\new_[5160]_  | ~\new_[5150]_  | ~\new_[5156]_ ;
  assign \new_[5150]_  = ~\new_[5151]_  | ~\new_[5154]_ ;
  assign \new_[5151]_  = ~\new_[5152]_  | ~\new_[1297]_  | ~\new_[1282]_ ;
  assign \new_[5152]_  = ~\new_[5153]_ ;
  assign \new_[5153]_  = \new_[5249]_  & \new_[1494]_ ;
  assign \new_[5154]_  = \new_[5155]_ ;
  assign \new_[5155]_  = ~\new_[1632]_  | ~\new_[1656]_ ;
  assign \new_[5156]_  = ~\new_[5157]_ ;
  assign \new_[5157]_  = ~\new_[1095]_  | ~\new_[5158]_  | ~\new_[1227]_ ;
  assign \new_[5158]_  = ~\new_[5159]_  & ~\new_[999]_ ;
  assign \new_[5159]_  = ~\new_[1203]_  | ~\new_[1222]_ ;
  assign \new_[5160]_  = ~\new_[4388]_  | ~\new_[1026]_ ;
  assign \new_[5161]_  = ~\new_[5155]_ ;
  assign n820 = \new_[5163]_  ? \new_[5165]_  : \new_[5164]_ ;
  assign \new_[5163]_  = ~\new_[5164]_ ;
  assign \new_[5164]_  = (~\desIn[18]  | ~\new_[2908]_ ) & (~\new_[1745]_  | ~\new_[2898]_ );
  assign \new_[5165]_  = ~\new_[5168]_  | ~\new_[5166]_  | ~\new_[5167]_ ;
  assign \new_[5166]_  = ~\new_[1177]_  | ~\new_[576]_ ;
  assign \new_[5167]_  = ~\new_[721]_  & ~\new_[645]_ ;
  assign \new_[5168]_  = ~\new_[584]_  | ~\new_[1318]_ ;
  assign \new_[5169]_  = ~\new_[5170]_  | ~\new_[5172]_ ;
  assign \new_[5170]_  = ~\new_[5171]_  & (~\new_[2807]_  | ~\new_[5068]_ );
  assign \new_[5171]_  = ~\new_[4192]_  & (~\new_[2880]_  | ~\new_[3264]_ );
  assign \new_[5172]_  = ~\new_[5173]_  & (~\new_[3094]_  | ~\new_[4065]_ );
  assign \new_[5173]_  = ~\new_[5174]_  & ~\new_[5176]_ ;
  assign \new_[5174]_  = ~\new_[5175]_ ;
  assign \new_[5175]_  = \new_[4287]_  & \new_[4283]_ ;
  assign \new_[5176]_  = \new_[5178]_  & \new_[5181]_ ;
  assign \new_[5177]_  = ~\new_[5178]_ ;
  assign \new_[5178]_  = ~\new_[5179]_ ;
  assign \new_[5179]_  = ~\new_[5180]_ ;
  assign \new_[5180]_  = ~\new_[3838]_  | ~\new_[3855]_ ;
  assign \new_[5181]_  = \new_[5182]_ ;
  assign \new_[5182]_  = ~\new_[3787]_  | ~\new_[3917]_ ;
  assign \new_[5183]_  = ~\new_[5177]_ ;
  assign n845 = \new_[5185]_  ? \new_[5187]_  : \new_[5186]_ ;
  assign \new_[5185]_  = ~\new_[4950]_  | (~\new_[1799]_  & ~\new_[3713]_ );
  assign \new_[5186]_  = ~\new_[5185]_ ;
  assign \new_[5187]_  = ~\new_[4463]_  | ~\new_[4458]_  | ~\new_[4457]_ ;
  assign \new_[5188]_  = ~\new_[5198]_  & (~\new_[5189]_  | ~\new_[5197]_ );
  assign \new_[5189]_  = ~\new_[5190]_ ;
  assign \new_[5190]_  = ~\new_[5191]_ ;
  assign \new_[5191]_  = ~\new_[5192]_ ;
  assign \new_[5192]_  = ~\new_[5193]_ ;
  assign \new_[5193]_  = \new_[5194]_  ? \new_[5195]_  : n1030;
  assign \new_[5194]_  = (~\new_[3459]_  & ~\new_[3914]_ ) | (~\new_[3809]_  & ~\desIn[19] );
  assign \new_[5195]_  = ~\new_[1837]_  & ~\new_[5143]_ ;
  assign \new_[5196]_  = ~\new_[5197]_ ;
  assign \new_[5197]_  = ~\new_[5115]_  & ~\new_[5110]_ ;
  assign \new_[5198]_  = ~\new_[802]_  | ~\new_[856]_ ;
  assign \new_[5199]_  = ~\new_[5200]_  | ~\new_[5201]_ ;
  assign \new_[5200]_  = ~\new_[1580]_  & ~\new_[1476]_ ;
  assign \new_[5201]_  = \new_[5202]_ ;
  assign \new_[5202]_  = ~\new_[5203]_  | ~\new_[5207]_ ;
  assign \new_[5203]_  = ~n1210 | (~\new_[5204]_  & ~\new_[5205]_ );
  assign \new_[5204]_  = ~\new_[5059]_  | ~\new_[5297]_ ;
  assign \new_[5205]_  = ~\new_[5058]_ ;
  assign n1210 = ~\new_[5056]_  | ~\new_[5057]_ ;
  assign \new_[5207]_  = ~\new_[5208]_  | ~\new_[5059]_  | ~\new_[5058]_  | ~\new_[5298]_ ;
  assign \new_[5208]_  = ~n1210;
  assign \new_[5209]_  = ~\new_[5201]_ ;
  assign \new_[5210]_  = ~\new_[5201]_ ;
  assign \new_[5211]_  = ~\new_[5202]_ ;
  assign \new_[5212]_  = ~\new_[5218]_  | ~\new_[5216]_  | ~\new_[5213]_  | ~\new_[5214]_ ;
  assign \new_[5213]_  = ~\new_[2498]_  & ~\new_[2103]_ ;
  assign \new_[5214]_  = ~\new_[2137]_  & ~\new_[5215]_ ;
  assign \new_[5215]_  = ~\new_[2230]_ ;
  assign \new_[5216]_  = ~\new_[5217]_  & (~\new_[2276]_  | ~\new_[4245]_ );
  assign \new_[5217]_  = ~\new_[2229]_  | ~\new_[2496]_ ;
  assign \new_[5218]_  = ~\new_[5219]_  & ~\new_[5220]_ ;
  assign \new_[5219]_  = ~\new_[2642]_  | ~\new_[2903]_ ;
  assign \new_[5220]_  = ~\new_[2497]_ ;
  assign \new_[5221]_  = ~\new_[5230]_  & (~\new_[5222]_  | ~\key2[4] );
  assign \new_[5222]_  = ~\new_[5223]_  | ~\new_[5227]_ ;
  assign \new_[5223]_  = ~\new_[5224]_ ;
  assign \new_[5224]_  = ~\new_[5225]_ ;
  assign \new_[5225]_  = ~\new_[5226]_ ;
  assign \new_[5226]_  = ~\new_[4971]_  & ~\new_[4412]_ ;
  assign \new_[5227]_  = ~\new_[5228]_ ;
  assign \new_[5228]_  = ~\new_[5229]_ ;
  assign \new_[5229]_  = ~\roundSel[4]  | ~\new_[4321]_  | ~\new_[4970]_ ;
  assign \new_[5230]_  = ~\new_[4305]_  & ~\new_[4254]_ ;
  assign \new_[5231]_  = (~\new_[3739]_  & ~\new_[4316]_ ) | (~\new_[1753]_  & ~\new_[3713]_ );
  assign \new_[5232]_  = ~\new_[5231]_ ;
  assign \new_[5233]_  = ~\new_[5237]_  | ~\new_[5236]_  | ~\new_[5235]_  | ~\new_[5234]_ ;
  assign \new_[5234]_  = ~\new_[4450]_  & ~\new_[757]_ ;
  assign \new_[5235]_  = ~\new_[4454]_  | ~\new_[4962]_ ;
  assign \new_[5236]_  = ~\new_[4453]_  | (~\new_[4415]_  & ~\new_[4416]_ );
  assign \new_[5237]_  = ~\new_[1144]_  | ~\new_[1041]_  | ~\new_[1321]_ ;
  assign n725 = ~\new_[511]_  | ~\new_[508]_ ;
  assign n735 = ~\new_[511]_  | ~\new_[508]_ ;
  assign \new_[5240]_  = ~\new_[5242]_ ;
  assign \new_[5241]_  = \new_[5240]_ ;
  assign \new_[5242]_  = ~\new_[3659]_ ;
  assign \new_[5243]_  = ~\new_[5244]_ ;
  assign \new_[5244]_  = \new_[4858]_ ;
  assign \new_[5245]_  = ~\new_[5246]_ ;
  assign \new_[5246]_  = \new_[5248]_ ;
  assign \new_[5247]_  = ~\new_[5248]_ ;
  assign \new_[5248]_  = ~\new_[4640]_ ;
  assign \new_[5249]_  = ~\new_[5250]_ ;
  assign \new_[5250]_  = \new_[4640]_ ;
  assign n750 = \new_[4629]_  ? \new_[4870]_  : \new_[4630]_ ;
  assign n770 = \new_[4629]_  ? \new_[4870]_  : \new_[4630]_ ;
  assign n620 = \new_[4498]_  ? \new_[4500]_  : \new_[4499]_ ;
  assign n625 = \new_[4498]_  ? \new_[4500]_  : \new_[4499]_ ;
  assign \new_[5255]_  = ~\new_[3825]_  | ~\new_[3965]_ ;
  assign \new_[5256]_  = ~\new_[3825]_  | ~\new_[3965]_ ;
  assign \new_[5257]_  = ~\new_[3800]_  | ~\new_[4014]_ ;
  assign \new_[5258]_  = ~\new_[3800]_  | ~\new_[4014]_ ;
  assign \new_[5259]_  = ~\new_[3775]_  | ~\new_[3917]_ ;
  assign \new_[5260]_  = ~\new_[3775]_  | ~\new_[3917]_ ;
  assign \new_[5261]_  = ~\new_[3777]_  | ~\new_[3906]_ ;
  assign \new_[5262]_  = ~\new_[3777]_  | ~\new_[3906]_ ;
  assign \new_[5263]_  = \new_[3631]_ ;
  assign n850 = ~\new_[4986]_  | ~\new_[523]_ ;
  assign n855 = ~\new_[4986]_  | ~\new_[523]_ ;
  assign \new_[5266]_  = ~\new_[4910]_  | ~\new_[3912]_ ;
  assign \new_[5267]_  = ~\new_[4910]_  | ~\new_[3912]_ ;
  assign \new_[5268]_  = ~\new_[3769]_  | ~\new_[3969]_ ;
  assign \new_[5269]_  = ~\new_[3769]_  | ~\new_[3969]_ ;
  assign \new_[5270]_  = ~\new_[3153]_  | ~\new_[3527]_ ;
  assign \new_[5271]_  = ~\new_[3153]_  | ~\new_[3527]_ ;
  assign \new_[5272]_  = ~\new_[3783]_  | ~\new_[4014]_ ;
  assign \new_[5273]_  = ~\new_[3783]_  | ~\new_[4014]_ ;
  assign n910 = \new_[5231]_  ? \new_[5233]_  : \new_[5232]_ ;
  assign n915 = \new_[5231]_  ? \new_[5233]_  : \new_[5232]_ ;
  assign \new_[5276]_  = ~\new_[3792]_  | ~\new_[5102]_ ;
  assign \new_[5277]_  = ~\new_[3792]_  | ~\new_[5102]_ ;
  assign \new_[5278]_  = ~\new_[4715]_  | ~\new_[4718]_ ;
  assign \new_[5279]_  = ~\new_[4715]_  | ~\new_[4718]_ ;
  assign \new_[5280]_  = ~\new_[3776]_  | ~\new_[3960]_ ;
  assign \new_[5281]_  = ~\new_[3776]_  | ~\new_[3960]_ ;
  assign \new_[5282]_  = ~\new_[4862]_  | ~\new_[4860]_ ;
  assign \new_[5283]_  = ~\new_[4862]_  | ~\new_[4860]_ ;
  assign \new_[5284]_  = ~\new_[5286]_ ;
  assign \new_[5285]_  = ~\new_[5287]_ ;
  assign \new_[5286]_  = \new_[5287]_ ;
  assign \new_[5287]_  = ~\new_[5044]_ ;
  assign \new_[5288]_  = \new_[3662]_ ;
  assign \new_[5289]_  = \new_[3662]_ ;
  assign \new_[5290]_  = ~\new_[5291]_ ;
  assign \new_[5291]_  = ~\new_[1349]_ ;
  assign \new_[5292]_  = \new_[1327]_ ;
  assign \new_[5293]_  = ~\new_[5051]_  | ~\new_[5052]_ ;
  assign \new_[5294]_  = ~\new_[5051]_  | ~\new_[5052]_ ;
  assign \new_[5295]_  = ~\new_[4661]_ ;
  assign \new_[5296]_  = ~\new_[4661]_ ;
  assign \new_[5297]_  = ~\new_[4855]_  & ~\new_[4549]_ ;
  assign \new_[5298]_  = ~\new_[4855]_  & ~\new_[4549]_ ;
  assign \new_[5299]_  = ~\new_[5300]_ ;
  assign \new_[5300]_  = ~\new_[5302]_ ;
  assign \new_[5301]_  = ~\new_[5302]_ ;
  assign \new_[5302]_  = ~\new_[5304]_ ;
  assign \new_[5303]_  = \new_[5304]_ ;
  assign \new_[5304]_  = ~\new_[5311]_ ;
  assign \new_[5305]_  = ~\new_[5311]_ ;
  assign \new_[5306]_  = ~\new_[5308]_ ;
  assign \new_[5307]_  = ~\new_[5308]_ ;
  assign \new_[5308]_  = \new_[5311]_ ;
  assign \new_[5309]_  = ~\new_[5310]_ ;
  assign \new_[5310]_  = ~\new_[5311]_ ;
  assign \new_[5311]_  = ~\new_[5314]_ ;
  assign \new_[5312]_  = ~\new_[5313]_ ;
  assign \new_[5313]_  = \new_[5311]_ ;
  assign \new_[5314]_  = ~\new_[4142]_ ;
  assign \desOut[0]  = n615;
  assign \desOut[1]  = n1140;
  assign \desOut[2]  = n905;
  assign \desOut[3]  = n985;
  assign \desOut[4]  = n845;
  assign \desOut[5]  = n1245;
  assign \desOut[6]  = n890;
  assign \desOut[7]  = n1150;
  assign \desOut[8]  = n785;
  assign \desOut[9]  = n1105;
  assign \desOut[10]  = n850;
  assign \desOut[11]  = n1205;
  assign \desOut[12]  = n815;
  assign \desOut[13]  = n1185;
  assign \desOut[14]  = n720;
  assign \desOut[15]  = n1210;
  assign \desOut[16]  = n790;
  assign \desOut[17]  = n1020;
  assign \desOut[18]  = n820;
  assign \desOut[19]  = n1030;
  assign \desOut[20]  = n620;
  assign \desOut[21]  = n1025;
  assign \desOut[22]  = n645;
  assign \desOut[23]  = n990;
  assign \desOut[24]  = n730;
  assign \desOut[25]  = n1015;
  assign \desOut[26]  = n765;
  assign \desOut[27]  = n1190;
  assign \desOut[28]  = n780;
  assign \desOut[29]  = n1215;
  assign \desOut[30]  = n665;
  assign \desOut[31]  = n1220;
  assign \desOut[32]  = n675;
  assign \desOut[33]  = n1240;
  assign \desOut[34]  = n825;
  assign \desOut[35]  = n1115;
  assign \desOut[36]  = n725;
  assign \desOut[37]  = n1135;
  assign \desOut[38]  = n705;
  assign \desOut[39]  = n1130;
  assign \desOut[40]  = n895;
  assign \desOut[41]  = n1005;
  assign \desOut[42]  = n685;
  assign \desOut[43]  = n1110;
  assign \desOut[44]  = n715;
  assign \desOut[45]  = n1225;
  assign \desOut[46]  = n835;
  assign \desOut[47]  = n1125;
  assign \desOut[48]  = n760;
  assign \desOut[49]  = n1035;
  assign \desOut[50]  = n880;
  assign \desOut[51]  = n1000;
  assign \desOut[52]  = n655;
  assign \desOut[53]  = n1010;
  assign \desOut[54]  = n640;
  assign \desOut[55]  = n1155;
  assign \desOut[56]  = n870;
  assign \desOut[57]  = n1055;
  assign \desOut[58]  = n910;
  assign \desOut[59]  = n995;
  assign \desOut[60]  = n925;
  assign \desOut[61]  = n1145;
  assign \desOut[62]  = n750;
  assign \desOut[63]  = n1120;
  assign n610 = n615;
  assign n630 = n645;
  assign n635 = n640;
  assign n650 = n655;
  assign n660 = n665;
  assign n670 = n675;
  assign n680 = n685;
  assign n690 = n715;
  assign n695 = n720;
  assign n700 = n705;
  assign n710 = n730;
  assign n740 = n760;
  assign n745 = n785;
  assign n755 = n765;
  assign n775 = n780;
  assign n795 = n820;
  assign n800 = n815;
  assign n805 = n825;
  assign n810 = n835;
  assign n840 = n845;
  assign n860 = n895;
  assign n865 = n870;
  assign n875 = n880;
  assign n885 = n890;
  assign n900 = n905;
  assign n920 = n925;
  assign n930 = n1010;
  assign n935 = n1000;
  assign n940 = n1005;
  assign n945 = n1030;
  assign n950 = n1025;
  assign n955 = n1020;
  assign n960 = n1015;
  assign n965 = n985;
  assign n970 = n990;
  assign n975 = n995;
  assign n980 = n1035;
  assign n1040 = n1055;
  assign n1045 = n1120;
  assign n1050 = n1105;
  assign n1060 = n1140;
  assign n1065 = n1135;
  assign n1070 = n1125;
  assign n1075 = n1130;
  assign n1080 = n1115;
  assign n1085 = n1145;
  assign n1090 = n1110;
  assign n1095 = n1150;
  assign n1100 = n1155;
  assign n1160 = n1215;
  assign n1165 = n1190;
  assign n1170 = n1220;
  assign n1175 = n1185;
  assign n1180 = n1210;
  assign n1195 = n1225;
  assign n1200 = n1205;
  assign n1230 = n1240;
  assign n1235 = n1245;
  always @ (posedge clock) begin
    \\FP_R_reg[25]  <= n610;
    \\R_reg[25]  <= n615;
    \\FP_R_reg[11]  <= n620;
    \\R_reg[11]  <= n625;
    \\FP_R_reg[3]  <= n630;
    \\R_reg[7]  <= n635;
    \\FP_R_reg[7]  <= n640;
    \\R_reg[3]  <= n645;
    \\FP_R_reg[15]  <= n650;
    \\R_reg[15]  <= n655;
    \\FP_R_reg[4]  <= n660;
    \\R_reg[4]  <= n665;
    \\FP_R_reg[29]  <= n670;
    \\R_reg[29]  <= n675;
    \\FP_R_reg[22]  <= n680;
    \\R_reg[22]  <= n685;
    \\R_reg[14]  <= n690;
    \\R_reg[2]  <= n695;
    \\FP_R_reg[5]  <= n700;
    \\R_reg[5]  <= n705;
    \\FP_R_reg[28]  <= n710;
    \\FP_R_reg[14]  <= n715;
    \\FP_R_reg[2]  <= n720;
    \\R_reg[13]  <= n725;
    \\R_reg[28]  <= n730;
    \\FP_R_reg[13]  <= n735;
    \\FP_R_reg[31]  <= n740;
    \\R_reg[26]  <= n745;
    \\FP_R_reg[8]  <= n750;
    \\FP_R_reg[20]  <= n755;
    \\R_reg[31]  <= n760;
    \\R_reg[20]  <= n765;
    \\R_reg[8]  <= n770;
    \\FP_R_reg[12]  <= n775;
    \\R_reg[12]  <= n780;
    \\FP_R_reg[26]  <= n785;
    \\FP_R_reg[27]  <= n790;
    \\FP_R_reg[19]  <= n795;
    \\FP_R_reg[10]  <= n800;
    \\FP_R_reg[21]  <= n805;
    \\FP_R_reg[6]  <= n810;
    \\R_reg[10]  <= n815;
    \\R_reg[19]  <= n820;
    \\R_reg[21]  <= n825;
    \\R_reg[27]  <= n830;
    \\R_reg[6]  <= n835;
    \\FP_R_reg[9]  <= n840;
    \\R_reg[9]  <= n845;
    \\FP_R_reg[18]  <= n850;
    \\R_reg[18]  <= n855;
    \\FP_R_reg[30]  <= n860;
    \\FP_R_reg[32]  <= n865;
    \\R_reg[32]  <= n870;
    \\FP_R_reg[23]  <= n875;
    \\R_reg[23]  <= n880;
    \\FP_R_reg[1]  <= n885;
    \\R_reg[1]  <= n890;
    \\R_reg[30]  <= n895;
    \\FP_R_reg[17]  <= n900;
    \\R_reg[17]  <= n905;
    \\FP_R_reg[24]  <= n910;
    \\R_reg[24]  <= n915;
    \\FP_R_reg[16]  <= n920;
    \\R_reg[16]  <= n925;
    \\L_reg[15]  <= n930;
    \\L_reg[23]  <= n935;
    \\L_reg[30]  <= n940;
    \\L_reg[19]  <= n945;
    \\L_reg[11]  <= n950;
    \\L_reg[27]  <= n955;
    \\L_reg[28]  <= n960;
    \\L_reg[17]  <= n965;
    \\L_reg[3]  <= n970;
    \\L_reg[24]  <= n975;
    \\L_reg[31]  <= n980;
    \\FP_R_reg[49]  <= n985;
    \\FP_R_reg[35]  <= n990;
    \\FP_R_reg[56]  <= n995;
    \\FP_R_reg[55]  <= n1000;
    \\FP_R_reg[62]  <= n1005;
    \\FP_R_reg[47]  <= n1010;
    \\FP_R_reg[60]  <= n1015;
    \\FP_R_reg[59]  <= n1020;
    \\FP_R_reg[43]  <= n1025;
    \\FP_R_reg[51]  <= n1030;
    \\FP_R_reg[63]  <= n1035;
    \\FP_R_reg[64]  <= n1040;
    \\L_reg[8]  <= n1045;
    \\L_reg[26]  <= n1050;
    \\L_reg[32]  <= n1055;
    \\L_reg[25]  <= n1060;
    \\L_reg[13]  <= n1065;
    \\L_reg[6]  <= n1070;
    \\L_reg[5]  <= n1075;
    \\L_reg[21]  <= n1080;
    \\L_reg[16]  <= n1085;
    \\L_reg[22]  <= n1090;
    \\L_reg[1]  <= n1095;
    \\L_reg[7]  <= n1100;
    \\FP_R_reg[58]  <= n1105;
    \\FP_R_reg[54]  <= n1110;
    \\FP_R_reg[53]  <= n1115;
    \\FP_R_reg[40]  <= n1120;
    \\FP_R_reg[38]  <= n1125;
    \\FP_R_reg[37]  <= n1130;
    \\FP_R_reg[45]  <= n1135;
    \\FP_R_reg[57]  <= n1140;
    \\FP_R_reg[48]  <= n1145;
    \\FP_R_reg[33]  <= n1150;
    \\FP_R_reg[39]  <= n1155;
    \\L_reg[12]  <= n1160;
    \\FP_R_reg[52]  <= n1165;
    \\FP_R_reg[36]  <= n1170;
    \\FP_R_reg[42]  <= n1175;
    \\FP_R_reg[34]  <= n1180;
    \\L_reg[10]  <= n1185;
    \\L_reg[20]  <= n1190;
    \\L_reg[14]  <= n1195;
    \\L_reg[18]  <= n1200;
    \\FP_R_reg[50]  <= n1205;
    \\L_reg[2]  <= n1210;
    \\FP_R_reg[44]  <= n1215;
    \\L_reg[4]  <= n1220;
    \\FP_R_reg[46]  <= n1225;
    \\FP_R_reg[61]  <= n1230;
    \\FP_R_reg[41]  <= n1235;
    \\L_reg[29]  <= n1240;
    \\L_reg[9]  <= n1245;
  end
endmodule


