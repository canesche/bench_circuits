module top ( 
    pa, pb, pc, pd, pe, pf, pg, ph, pi, pj,
    pp, pk, pl, pm, pn, po  );
  input  pa, pb, pc, pd, pe, pf, pg, ph, pi, pj;
  output pp, pk, pl, pm, pn, po;
  wire new_n17_, new_n19_, new_n21_, new_n22_, new_n23_, new_n25_, new_n26_,
    new_n27_, new_n28_, new_n29_, new_n30_, new_n31_, new_n32_, new_n33_,
    new_n34_, new_n35_, new_n36_, new_n37_, new_n38_, new_n39_, new_n40_,
    new_n41_, new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n47_,
    new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_,
    new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_,
    new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_,
    new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_;
  assign new_n17_ = ~pa & ~pc;
  assign pn = pb & pd;
  assign new_n19_ = ~pb & ~pd;
  assign pm = pn | new_n19_;
  assign new_n21_ = new_n17_ & pm;
  assign new_n22_ = pa & pc;
  assign new_n23_ = pm & new_n22_;
  assign pp = new_n21_ | new_n23_;
  assign new_n25_ = pa & pg;
  assign new_n26_ = ph & new_n25_;
  assign new_n27_ = ~pj & new_n26_;
  assign new_n28_ = ~pg & ~ph;
  assign new_n29_ = ~pj & new_n28_;
  assign new_n30_ = ~pf & ~pg;
  assign new_n31_ = ~pj & new_n30_;
  assign new_n32_ = ~new_n29_ & ~new_n31_;
  assign new_n33_ = ~pa & ~new_n32_;
  assign new_n34_ = ~pe & new_n33_;
  assign new_n35_ = ~pa & pc;
  assign new_n36_ = pg & ~ph;
  assign new_n37_ = pf & pj;
  assign new_n38_ = new_n35_ & new_n36_;
  assign new_n39_ = new_n37_ & new_n38_;
  assign new_n40_ = ~pe & new_n39_;
  assign new_n41_ = ~ph & ~pj;
  assign new_n42_ = ~pg & new_n41_;
  assign new_n43_ = pg & pj;
  assign new_n44_ = ~new_n42_ & ~new_n43_;
  assign new_n45_ = pe & ~pf;
  assign new_n46_ = ~new_n44_ & new_n45_;
  assign new_n47_ = ~new_n17_ & new_n46_;
  assign new_n48_ = pa & ~pc;
  assign new_n49_ = new_n37_ & new_n48_;
  assign new_n50_ = ~pe & new_n49_;
  assign new_n51_ = ~new_n36_ & new_n37_;
  assign new_n52_ = ~pe & new_n51_;
  assign new_n53_ = ~pf & pg;
  assign new_n54_ = ph & ~pj;
  assign new_n55_ = new_n53_ & new_n54_;
  assign new_n56_ = pe & new_n55_;
  assign new_n57_ = pe & pf;
  assign new_n58_ = new_n36_ & new_n57_;
  assign new_n59_ = ~new_n52_ & ~new_n56_;
  assign new_n60_ = ~new_n58_ & new_n59_;
  assign new_n61_ = ~pc & ~new_n60_;
  assign new_n62_ = ~pe & ~pf;
  assign new_n63_ = ph & new_n62_;
  assign new_n64_ = pj & new_n63_;
  assign new_n65_ = ~pg & new_n64_;
  assign new_n66_ = new_n22_ & new_n65_;
  assign new_n67_ = new_n36_ & new_n62_;
  assign new_n68_ = new_n22_ & new_n67_;
  assign new_n69_ = ph & new_n57_;
  assign new_n70_ = pj & new_n69_;
  assign new_n71_ = ~pg & new_n70_;
  assign new_n72_ = new_n22_ & new_n71_;
  assign new_n73_ = ~new_n34_ & ~new_n40_;
  assign new_n74_ = ~new_n47_ & ~new_n50_;
  assign new_n75_ = new_n73_ & new_n74_;
  assign new_n76_ = ~new_n68_ & ~new_n72_;
  assign new_n77_ = ~new_n61_ & ~new_n66_;
  assign new_n78_ = new_n76_ & new_n77_;
  assign new_n79_ = new_n75_ & new_n78_;
  assign new_n80_ = ~pg & ~new_n79_;
  assign new_n81_ = ~pe & new_n80_;
  assign new_n82_ = pc & new_n81_;
  assign new_n83_ = ~pj & new_n82_;
  assign new_n84_ = new_n57_ & new_n79_;
  assign new_n85_ = ~pg & new_n84_;
  assign new_n86_ = ph & new_n85_;
  assign new_n87_ = pj & new_n86_;
  assign new_n88_ = ~new_n57_ & new_n79_;
  assign new_n89_ = ph & new_n88_;
  assign new_n90_ = new_n25_ & new_n89_;
  assign new_n91_ = pj & new_n90_;
  assign new_n92_ = pg & new_n79_;
  assign new_n93_ = ~new_n80_ & ~new_n92_;
  assign new_n94_ = ~pe & pf;
  assign new_n95_ = ~ph & ~new_n93_;
  assign new_n96_ = new_n94_ & new_n95_;
  assign new_n97_ = pj & new_n96_;
  assign new_n98_ = pj & new_n36_;
  assign new_n99_ = new_n22_ & new_n45_;
  assign new_n100_ = new_n98_ & new_n99_;
  assign new_n101_ = new_n62_ & new_n79_;
  assign new_n102_ = new_n98_ & new_n101_;
  assign new_n103_ = ~pe & ph;
  assign new_n104_ = new_n37_ & new_n103_;
  assign new_n105_ = pa & new_n104_;
  assign new_n106_ = pa & ~new_n79_;
  assign new_n107_ = new_n57_ & new_n106_;
  assign new_n108_ = new_n98_ & new_n107_;
  assign new_n109_ = ~new_n79_ & new_n104_;
  assign new_n110_ = ~new_n108_ & ~new_n109_;
  assign new_n111_ = ~new_n100_ & ~new_n102_;
  assign new_n112_ = ~new_n105_ & new_n111_;
  assign new_n113_ = new_n110_ & new_n112_;
  assign new_n114_ = pg & new_n57_;
  assign new_n115_ = ~ph & new_n113_;
  assign new_n116_ = new_n114_ & new_n115_;
  assign new_n117_ = pj & new_n116_;
  assign new_n118_ = ph & new_n114_;
  assign new_n119_ = ~pa & new_n118_;
  assign new_n120_ = pj & new_n119_;
  assign new_n121_ = ~pg & new_n22_;
  assign new_n122_ = new_n104_ & new_n121_;
  assign new_n123_ = new_n45_ & new_n98_;
  assign new_n124_ = new_n113_ & new_n123_;
  assign new_n125_ = ~new_n122_ & ~new_n124_;
  assign new_n126_ = pe & new_n53_;
  assign new_n127_ = ~ph & new_n126_;
  assign new_n128_ = ~new_n79_ & new_n127_;
  assign new_n129_ = pj & new_n128_;
  assign new_n130_ = new_n125_ & new_n129_;
  assign new_n131_ = new_n53_ & ~new_n113_;
  assign new_n132_ = ~ph & new_n131_;
  assign new_n133_ = ~pa & new_n132_;
  assign new_n134_ = pj & new_n133_;
  assign new_n135_ = ~pe & new_n134_;
  assign new_n136_ = new_n94_ & new_n113_;
  assign new_n137_ = ~pg & new_n136_;
  assign new_n138_ = ph & new_n137_;
  assign new_n139_ = pj & new_n138_;
  assign new_n140_ = ~new_n125_ & new_n139_;
  assign new_n141_ = new_n79_ & new_n127_;
  assign new_n142_ = pj & new_n141_;
  assign new_n143_ = ~new_n125_ & new_n142_;
  assign new_n144_ = new_n94_ & ~new_n113_;
  assign new_n145_ = ~pg & new_n144_;
  assign new_n146_ = ph & new_n145_;
  assign new_n147_ = pj & new_n146_;
  assign new_n148_ = new_n125_ & new_n147_;
  assign new_n149_ = pe & new_n35_;
  assign new_n150_ = ~pf & new_n149_;
  assign new_n151_ = ~pg & new_n150_;
  assign new_n152_ = pj & new_n151_;
  assign new_n153_ = ~pa & new_n62_;
  assign new_n154_ = ph & new_n153_;
  assign new_n155_ = ~new_n79_ & new_n154_;
  assign new_n156_ = pj & new_n155_;
  assign new_n157_ = pe & new_n48_;
  assign new_n158_ = ~pf & new_n157_;
  assign new_n159_ = ~pg & new_n158_;
  assign new_n160_ = pj & new_n159_;
  assign new_n161_ = pa & ~pe;
  assign new_n162_ = new_n79_ & new_n161_;
  assign new_n163_ = ~pf & new_n162_;
  assign new_n164_ = ~pg & new_n163_;
  assign new_n165_ = pj & new_n164_;
  assign new_n166_ = new_n113_ & new_n161_;
  assign new_n167_ = ~pf & new_n166_;
  assign new_n168_ = ~ph & new_n167_;
  assign new_n169_ = pj & new_n168_;
  assign new_n170_ = pa & ~new_n57_;
  assign new_n171_ = ~pg & new_n170_;
  assign new_n172_ = ~ph & new_n171_;
  assign new_n173_ = pj & new_n172_;
  assign new_n174_ = ~pa & ~new_n79_;
  assign new_n175_ = pg & new_n174_;
  assign new_n176_ = ph & new_n175_;
  assign new_n177_ = pj & new_n176_;
  assign new_n178_ = ~new_n140_ & ~new_n143_;
  assign new_n179_ = ~new_n130_ & ~new_n135_;
  assign new_n180_ = new_n178_ & new_n179_;
  assign new_n181_ = ~new_n117_ & ~new_n120_;
  assign new_n182_ = ~new_n87_ & ~new_n91_;
  assign new_n183_ = ~new_n97_ & new_n182_;
  assign new_n184_ = new_n181_ & new_n183_;
  assign new_n185_ = new_n180_ & new_n184_;
  assign new_n186_ = ~new_n173_ & ~new_n177_;
  assign new_n187_ = ~new_n165_ & ~new_n169_;
  assign new_n188_ = new_n186_ & new_n187_;
  assign new_n189_ = ~new_n148_ & ~new_n152_;
  assign new_n190_ = ~new_n156_ & ~new_n160_;
  assign new_n191_ = new_n189_ & new_n190_;
  assign new_n192_ = new_n188_ & new_n191_;
  assign new_n193_ = new_n185_ & new_n192_;
  assign new_n194_ = ~pi & new_n193_;
  assign new_n195_ = pj & new_n194_;
  assign new_n196_ = ~pg & new_n57_;
  assign new_n197_ = ~ph & new_n196_;
  assign new_n198_ = pj & new_n197_;
  assign new_n199_ = pi & ~new_n193_;
  assign new_n200_ = pj & new_n199_;
  assign new_n201_ = ~ph & new_n45_;
  assign new_n202_ = ~pc & new_n201_;
  assign new_n203_ = ~pj & new_n202_;
  assign new_n204_ = pg & new_n203_;
  assign new_n205_ = ~pf & new_n79_;
  assign new_n206_ = ~ph & new_n205_;
  assign new_n207_ = pe & new_n206_;
  assign new_n208_ = ~pj & new_n207_;
  assign new_n209_ = ~pg & new_n208_;
  assign new_n210_ = pg & ~new_n79_;
  assign new_n211_ = ph & new_n210_;
  assign new_n212_ = ~pf & new_n211_;
  assign new_n213_ = ~pj & new_n212_;
  assign new_n214_ = pe & ~pg;
  assign new_n215_ = new_n35_ & new_n214_;
  assign new_n216_ = ph & new_n215_;
  assign new_n217_ = ~pf & new_n216_;
  assign new_n218_ = ~pj & new_n217_;
  assign new_n219_ = new_n17_ & new_n36_;
  assign new_n220_ = ~pe & new_n219_;
  assign new_n221_ = pf & new_n220_;
  assign new_n222_ = ~pj & new_n221_;
  assign new_n223_ = pg & new_n106_;
  assign new_n224_ = pe & new_n223_;
  assign new_n225_ = pf & new_n224_;
  assign new_n226_ = ~pj & new_n225_;
  assign new_n227_ = ph & new_n22_;
  assign new_n228_ = pf & new_n227_;
  assign new_n229_ = ~pj & new_n228_;
  assign new_n230_ = ~pe & pg;
  assign new_n231_ = pf & new_n22_;
  assign new_n232_ = new_n230_ & new_n231_;
  assign new_n233_ = ~pj & new_n232_;
  assign new_n234_ = pc & new_n103_;
  assign new_n235_ = pf & new_n234_;
  assign new_n236_ = ~pj & new_n235_;
  assign new_n237_ = ph & new_n230_;
  assign new_n238_ = ~pf & new_n237_;
  assign new_n239_ = ~pj & new_n238_;
  assign new_n240_ = ph & new_n161_;
  assign new_n241_ = ~pf & new_n240_;
  assign new_n242_ = ~pj & new_n241_;
  assign new_n243_ = ~pe & ~new_n93_;
  assign new_n244_ = ~pf & new_n243_;
  assign new_n245_ = ~pj & new_n244_;
  assign new_n246_ = ph & new_n48_;
  assign new_n247_ = ~pf & new_n246_;
  assign new_n248_ = ~pj & new_n247_;
  assign new_n249_ = ~new_n245_ & ~new_n248_;
  assign new_n250_ = ~new_n239_ & ~new_n242_;
  assign new_n251_ = new_n249_ & new_n250_;
  assign new_n252_ = ~new_n233_ & ~new_n236_;
  assign new_n253_ = ~new_n222_ & ~new_n226_;
  assign new_n254_ = ~new_n229_ & new_n253_;
  assign new_n255_ = new_n252_ & new_n254_;
  assign new_n256_ = new_n251_ & new_n255_;
  assign new_n257_ = ~new_n213_ & ~new_n218_;
  assign new_n258_ = ~new_n204_ & ~new_n209_;
  assign new_n259_ = new_n257_ & new_n258_;
  assign new_n260_ = ~new_n198_ & ~new_n200_;
  assign new_n261_ = ~new_n27_ & ~new_n83_;
  assign new_n262_ = ~new_n195_ & new_n261_;
  assign new_n263_ = new_n260_ & new_n262_;
  assign new_n264_ = new_n259_ & new_n263_;
  assign pk = ~new_n256_ | ~new_n264_;
  assign new_n266_ = ~new_n19_ & new_n45_;
  assign new_n267_ = ~new_n44_ & new_n266_;
  assign new_n268_ = ~pb & ~new_n32_;
  assign new_n269_ = ~pe & new_n268_;
  assign new_n270_ = ~pf & new_n36_;
  assign new_n271_ = pn & new_n270_;
  assign new_n272_ = pj & new_n271_;
  assign new_n273_ = ~pe & new_n271_;
  assign new_n274_ = ~pd & ~new_n60_;
  assign new_n275_ = pb & ~pd;
  assign new_n276_ = pf & new_n275_;
  assign new_n277_ = ~pe & new_n276_;
  assign new_n278_ = ~new_n35_ & new_n277_;
  assign new_n279_ = pj & new_n278_;
  assign new_n280_ = ~pb & pd;
  assign new_n281_ = pf & ~new_n35_;
  assign new_n282_ = ~pe & new_n281_;
  assign new_n283_ = new_n36_ & new_n282_;
  assign new_n284_ = pj & new_n283_;
  assign new_n285_ = new_n280_ & new_n284_;
  assign new_n286_ = ~pf & new_n25_;
  assign new_n287_ = ~pe & new_n286_;
  assign new_n288_ = ph & new_n287_;
  assign new_n289_ = pj & new_n288_;
  assign new_n290_ = pf & new_n35_;
  assign new_n291_ = pj & new_n290_;
  assign new_n292_ = ~pe & new_n291_;
  assign new_n293_ = new_n19_ & new_n292_;
  assign new_n294_ = ~pg & pn;
  assign new_n295_ = ~pf & ph;
  assign new_n296_ = pj & new_n295_;
  assign new_n297_ = ~pe & new_n296_;
  assign new_n298_ = new_n294_ & new_n297_;
  assign new_n299_ = ph & new_n37_;
  assign new_n300_ = pe & new_n299_;
  assign new_n301_ = new_n294_ & new_n300_;
  assign new_n302_ = pn & new_n35_;
  assign new_n303_ = ~pe & new_n302_;
  assign new_n304_ = new_n36_ & new_n303_;
  assign new_n305_ = pj & new_n304_;
  assign new_n306_ = ~new_n298_ & ~new_n301_;
  assign new_n307_ = ~new_n305_ & new_n306_;
  assign new_n308_ = ~new_n285_ & ~new_n289_;
  assign new_n309_ = ~new_n293_ & new_n308_;
  assign new_n310_ = new_n307_ & new_n309_;
  assign new_n311_ = ~new_n267_ & ~new_n269_;
  assign new_n312_ = ~new_n272_ & new_n311_;
  assign new_n313_ = ~new_n273_ & ~new_n274_;
  assign new_n314_ = ~new_n279_ & new_n313_;
  assign new_n315_ = new_n312_ & new_n314_;
  assign new_n316_ = new_n310_ & new_n315_;
  assign new_n317_ = ~pg & ~new_n316_;
  assign new_n318_ = ~pe & new_n317_;
  assign new_n319_ = pd & new_n318_;
  assign new_n320_ = ~pj & new_n319_;
  assign new_n321_ = ~pf & new_n318_;
  assign new_n322_ = ~pj & new_n321_;
  assign new_n323_ = ~pf & new_n214_;
  assign new_n324_ = new_n22_ & new_n323_;
  assign new_n325_ = new_n19_ & new_n324_;
  assign new_n326_ = ph & new_n325_;
  assign new_n327_ = pj & new_n326_;
  assign new_n328_ = new_n280_ & new_n323_;
  assign new_n329_ = ~new_n22_ & new_n328_;
  assign new_n330_ = pj & new_n329_;
  assign new_n331_ = pd & new_n323_;
  assign new_n332_ = ~ph & new_n331_;
  assign new_n333_ = pj & new_n332_;
  assign new_n334_ = new_n62_ & new_n316_;
  assign new_n335_ = new_n98_ & new_n334_;
  assign new_n336_ = pn & new_n45_;
  assign new_n337_ = new_n98_ & new_n336_;
  assign new_n338_ = pb & new_n104_;
  assign new_n339_ = pb & ~new_n316_;
  assign new_n340_ = new_n57_ & new_n339_;
  assign new_n341_ = new_n98_ & new_n340_;
  assign new_n342_ = new_n104_ & ~new_n316_;
  assign new_n343_ = ~new_n341_ & ~new_n342_;
  assign new_n344_ = ~new_n335_ & ~new_n337_;
  assign new_n345_ = ~new_n338_ & new_n344_;
  assign new_n346_ = new_n343_ & new_n345_;
  assign new_n347_ = new_n57_ & new_n113_;
  assign new_n348_ = new_n346_ & new_n347_;
  assign new_n349_ = pg & new_n348_;
  assign new_n350_ = ~ph & new_n349_;
  assign new_n351_ = pj & new_n350_;
  assign new_n352_ = pn & new_n324_;
  assign new_n353_ = pj & new_n352_;
  assign new_n354_ = new_n123_ & new_n346_;
  assign new_n355_ = new_n104_ & new_n294_;
  assign new_n356_ = ~new_n354_ & ~new_n355_;
  assign new_n357_ = ~new_n113_ & ~new_n125_;
  assign new_n358_ = new_n94_ & ~new_n346_;
  assign new_n359_ = ~pg & new_n358_;
  assign new_n360_ = ph & new_n359_;
  assign new_n361_ = pj & new_n360_;
  assign new_n362_ = new_n356_ & new_n361_;
  assign new_n363_ = ~new_n357_ & new_n362_;
  assign new_n364_ = pb & new_n25_;
  assign new_n365_ = ph & new_n364_;
  assign new_n366_ = new_n57_ & new_n365_;
  assign new_n367_ = pj & new_n366_;
  assign new_n368_ = new_n94_ & new_n346_;
  assign new_n369_ = ~pg & new_n368_;
  assign new_n370_ = ph & new_n369_;
  assign new_n371_ = pj & new_n370_;
  assign new_n372_ = ~new_n356_ & new_n371_;
  assign new_n373_ = ~new_n357_ & new_n372_;
  assign new_n374_ = pa & ~new_n113_;
  assign new_n375_ = ~new_n346_ & ~new_n374_;
  assign new_n376_ = new_n346_ & new_n374_;
  assign new_n377_ = ~new_n375_ & ~new_n376_;
  assign new_n378_ = ~pb & ~new_n377_;
  assign new_n379_ = pg & new_n378_;
  assign new_n380_ = ~ph & new_n379_;
  assign new_n381_ = pj & new_n380_;
  assign new_n382_ = new_n62_ & new_n381_;
  assign new_n383_ = new_n57_ & ~new_n113_;
  assign new_n384_ = pg & new_n383_;
  assign new_n385_ = ~ph & new_n384_;
  assign new_n386_ = pj & new_n385_;
  assign new_n387_ = ~new_n346_ & new_n386_;
  assign new_n388_ = ~pb & new_n57_;
  assign new_n389_ = pg & new_n388_;
  assign new_n390_ = ph & new_n389_;
  assign new_n391_ = pj & new_n390_;
  assign new_n392_ = ~pa & new_n391_;
  assign new_n393_ = ~new_n79_ & ~new_n125_;
  assign new_n394_ = new_n45_ & ~new_n316_;
  assign new_n395_ = pg & new_n394_;
  assign new_n396_ = ~ph & new_n395_;
  assign new_n397_ = pj & new_n396_;
  assign new_n398_ = new_n356_ & new_n397_;
  assign new_n399_ = ~new_n393_ & new_n398_;
  assign new_n400_ = ~new_n79_ & ~new_n316_;
  assign new_n401_ = ~ph & new_n400_;
  assign new_n402_ = new_n94_ & new_n401_;
  assign new_n403_ = pj & new_n402_;
  assign new_n404_ = new_n45_ & new_n316_;
  assign new_n405_ = pg & new_n404_;
  assign new_n406_ = ~ph & new_n405_;
  assign new_n407_ = pj & new_n406_;
  assign new_n408_ = ~new_n356_ & new_n407_;
  assign new_n409_ = ~new_n393_ & new_n408_;
  assign new_n410_ = ~new_n62_ & ~new_n230_;
  assign new_n411_ = ~new_n53_ & new_n410_;
  assign new_n412_ = ~new_n106_ & new_n316_;
  assign new_n413_ = new_n106_ & ~new_n316_;
  assign new_n414_ = ~new_n412_ & ~new_n413_;
  assign new_n415_ = pb & ~new_n411_;
  assign new_n416_ = ~new_n414_ & new_n415_;
  assign new_n417_ = ph & new_n416_;
  assign new_n418_ = pj & new_n417_;
  assign new_n419_ = new_n356_ & new_n371_;
  assign new_n420_ = new_n357_ & new_n419_;
  assign new_n421_ = ~pb & ~new_n411_;
  assign new_n422_ = new_n414_ & new_n421_;
  assign new_n423_ = ph & new_n422_;
  assign new_n424_ = pj & new_n423_;
  assign new_n425_ = ~new_n356_ & new_n361_;
  assign new_n426_ = new_n357_ & new_n425_;
  assign new_n427_ = new_n80_ & ~new_n316_;
  assign new_n428_ = ph & new_n427_;
  assign new_n429_ = new_n57_ & new_n428_;
  assign new_n430_ = pj & new_n429_;
  assign new_n431_ = new_n356_ & new_n407_;
  assign new_n432_ = new_n393_ & new_n431_;
  assign new_n433_ = new_n79_ & new_n316_;
  assign new_n434_ = new_n94_ & new_n433_;
  assign new_n435_ = pg & new_n434_;
  assign new_n436_ = ~ph & new_n435_;
  assign new_n437_ = pj & new_n436_;
  assign new_n438_ = ~new_n356_ & new_n397_;
  assign new_n439_ = new_n393_ & new_n438_;
  assign new_n440_ = new_n57_ & new_n433_;
  assign new_n441_ = ~pg & new_n440_;
  assign new_n442_ = ph & new_n441_;
  assign new_n443_ = pj & new_n442_;
  assign new_n444_ = pb & ~new_n57_;
  assign new_n445_ = ~pg & new_n444_;
  assign new_n446_ = ~ph & new_n445_;
  assign new_n447_ = pj & new_n446_;
  assign new_n448_ = pb & ~pe;
  assign new_n449_ = ~ph & new_n377_;
  assign new_n450_ = new_n448_ & new_n449_;
  assign new_n451_ = ~pf & new_n450_;
  assign new_n452_ = pj & new_n451_;
  assign new_n453_ = new_n94_ & ~new_n316_;
  assign new_n454_ = ~pg & new_n453_;
  assign new_n455_ = ~ph & new_n454_;
  assign new_n456_ = pj & new_n455_;
  assign new_n457_ = new_n275_ & new_n323_;
  assign new_n458_ = ~new_n22_ & new_n457_;
  assign new_n459_ = pj & new_n458_;
  assign new_n460_ = new_n30_ & ~new_n414_;
  assign new_n461_ = new_n448_ & new_n460_;
  assign new_n462_ = pj & new_n461_;
  assign new_n463_ = ~new_n456_ & ~new_n459_;
  assign new_n464_ = ~new_n462_ & new_n463_;
  assign new_n465_ = ~new_n447_ & ~new_n452_;
  assign new_n466_ = ~new_n439_ & ~new_n443_;
  assign new_n467_ = new_n465_ & new_n466_;
  assign new_n468_ = new_n464_ & new_n467_;
  assign new_n469_ = ~new_n424_ & ~new_n426_;
  assign new_n470_ = ~new_n418_ & ~new_n420_;
  assign new_n471_ = new_n469_ & new_n470_;
  assign new_n472_ = ~new_n430_ & ~new_n432_;
  assign new_n473_ = ~new_n437_ & new_n472_;
  assign new_n474_ = new_n471_ & new_n473_;
  assign new_n475_ = new_n468_ & new_n474_;
  assign new_n476_ = ~new_n399_ & ~new_n403_;
  assign new_n477_ = ~new_n409_ & new_n476_;
  assign new_n478_ = ~new_n387_ & ~new_n392_;
  assign new_n479_ = ~new_n373_ & ~new_n382_;
  assign new_n480_ = new_n478_ & new_n479_;
  assign new_n481_ = new_n477_ & new_n480_;
  assign new_n482_ = ~new_n353_ & ~new_n363_;
  assign new_n483_ = ~new_n367_ & new_n482_;
  assign new_n484_ = ~new_n327_ & ~new_n330_;
  assign new_n485_ = ~new_n333_ & ~new_n351_;
  assign new_n486_ = new_n484_ & new_n485_;
  assign new_n487_ = new_n483_ & new_n486_;
  assign new_n488_ = new_n481_ & new_n487_;
  assign new_n489_ = new_n475_ & new_n488_;
  assign new_n490_ = pi & ~new_n489_;
  assign new_n491_ = pj & new_n490_;
  assign new_n492_ = new_n193_ & ~new_n489_;
  assign new_n493_ = pj & new_n492_;
  assign new_n494_ = pe & new_n339_;
  assign new_n495_ = pf & new_n494_;
  assign new_n496_ = pg & new_n495_;
  assign new_n497_ = ~pj & new_n496_;
  assign new_n498_ = new_n19_ & new_n36_;
  assign new_n499_ = pf & new_n498_;
  assign new_n500_ = ~pe & new_n499_;
  assign new_n501_ = ~pj & new_n500_;
  assign new_n502_ = ~ph & new_n53_;
  assign new_n503_ = ~pd & new_n502_;
  assign new_n504_ = ~pj & new_n503_;
  assign new_n505_ = pe & new_n504_;
  assign new_n506_ = ~pg & new_n316_;
  assign new_n507_ = ~ph & new_n506_;
  assign new_n508_ = ~pf & new_n507_;
  assign new_n509_ = ~pj & new_n508_;
  assign new_n510_ = pe & new_n509_;
  assign new_n511_ = ph & pn;
  assign new_n512_ = pf & new_n511_;
  assign new_n513_ = ~pj & new_n512_;
  assign new_n514_ = pf & pn;
  assign new_n515_ = new_n230_ & new_n514_;
  assign new_n516_ = ~pj & new_n515_;
  assign new_n517_ = pg & ~new_n316_;
  assign new_n518_ = ph & new_n517_;
  assign new_n519_ = ~pf & new_n518_;
  assign new_n520_ = ~pj & new_n519_;
  assign new_n521_ = new_n214_ & new_n280_;
  assign new_n522_ = ph & new_n521_;
  assign new_n523_ = ~pf & new_n522_;
  assign new_n524_ = ~pj & new_n523_;
  assign new_n525_ = ph & new_n448_;
  assign new_n526_ = ~pf & new_n525_;
  assign new_n527_ = ~pj & new_n526_;
  assign new_n528_ = pd & new_n103_;
  assign new_n529_ = pf & new_n528_;
  assign new_n530_ = ~pj & new_n529_;
  assign new_n531_ = ph & new_n275_;
  assign new_n532_ = ~pf & new_n531_;
  assign new_n533_ = ~pj & new_n532_;
  assign new_n534_ = ~pf & new_n316_;
  assign new_n535_ = new_n230_ & new_n534_;
  assign new_n536_ = ~pj & new_n535_;
  assign new_n537_ = ~pi & new_n489_;
  assign new_n538_ = ~new_n193_ & new_n537_;
  assign new_n539_ = pj & new_n538_;
  assign new_n540_ = pg & ph;
  assign new_n541_ = pb & new_n540_;
  assign new_n542_ = ~pj & new_n541_;
  assign new_n543_ = ~new_n539_ & ~new_n542_;
  assign new_n544_ = ~new_n239_ & ~new_n533_;
  assign new_n545_ = ~new_n536_ & new_n544_;
  assign new_n546_ = new_n543_ & new_n545_;
  assign new_n547_ = ~new_n527_ & ~new_n530_;
  assign new_n548_ = ~new_n516_ & ~new_n520_;
  assign new_n549_ = ~new_n524_ & new_n548_;
  assign new_n550_ = new_n547_ & new_n549_;
  assign new_n551_ = new_n546_ & new_n550_;
  assign new_n552_ = ~new_n198_ & ~new_n493_;
  assign new_n553_ = ~new_n320_ & ~new_n322_;
  assign new_n554_ = ~new_n491_ & new_n553_;
  assign new_n555_ = new_n552_ & new_n554_;
  assign new_n556_ = ~new_n510_ & ~new_n513_;
  assign new_n557_ = ~new_n497_ & ~new_n501_;
  assign new_n558_ = ~new_n505_ & new_n557_;
  assign new_n559_ = new_n556_ & new_n558_;
  assign new_n560_ = new_n555_ & new_n559_;
  assign pl = ~new_n551_ | ~new_n560_;
  assign new_n562_ = ~pi & ~new_n489_;
  assign new_n563_ = ~new_n193_ & new_n562_;
  assign new_n564_ = pj & new_n563_;
  assign new_n565_ = ph & ~new_n19_;
  assign new_n566_ = new_n324_ & new_n565_;
  assign new_n567_ = pj & new_n566_;
  assign new_n568_ = ~ph & new_n348_;
  assign new_n569_ = pj & new_n568_;
  assign new_n570_ = new_n196_ & new_n433_;
  assign new_n571_ = pj & new_n570_;
  assign new_n572_ = ~pg & ~new_n356_;
  assign new_n573_ = ph & new_n572_;
  assign new_n574_ = new_n94_ & new_n573_;
  assign new_n575_ = pj & new_n574_;
  assign new_n576_ = new_n357_ & new_n575_;
  assign new_n577_ = pe & ~new_n356_;
  assign new_n578_ = ~ph & new_n577_;
  assign new_n579_ = new_n53_ & new_n578_;
  assign new_n580_ = pj & new_n579_;
  assign new_n581_ = ~new_n316_ & new_n580_;
  assign new_n582_ = new_n393_ & new_n580_;
  assign new_n583_ = pe & ~new_n316_;
  assign new_n584_ = ~ph & new_n583_;
  assign new_n585_ = new_n53_ & new_n584_;
  assign new_n586_ = pj & new_n585_;
  assign new_n587_ = new_n393_ & new_n586_;
  assign new_n588_ = ~new_n346_ & new_n374_;
  assign new_n589_ = ~ph & new_n588_;
  assign new_n590_ = new_n53_ & new_n589_;
  assign new_n591_ = pj & new_n590_;
  assign new_n592_ = ~pe & new_n591_;
  assign new_n593_ = ~pe & ~new_n346_;
  assign new_n594_ = ~ph & new_n593_;
  assign new_n595_ = new_n53_ & new_n594_;
  assign new_n596_ = pj & new_n595_;
  assign new_n597_ = pb & new_n596_;
  assign new_n598_ = ~pg & new_n94_;
  assign new_n599_ = ph & new_n598_;
  assign new_n600_ = ~new_n346_ & new_n599_;
  assign new_n601_ = pj & new_n600_;
  assign new_n602_ = ~new_n356_ & new_n601_;
  assign new_n603_ = new_n357_ & new_n601_;
  assign new_n604_ = pb & new_n106_;
  assign new_n605_ = ph & new_n604_;
  assign new_n606_ = ~new_n411_ & new_n605_;
  assign new_n607_ = pj & new_n606_;
  assign new_n608_ = ph & new_n413_;
  assign new_n609_ = ~new_n411_ & new_n608_;
  assign new_n610_ = pj & new_n609_;
  assign new_n611_ = ~pa & ~pb;
  assign new_n612_ = ph & new_n611_;
  assign new_n613_ = new_n114_ & new_n612_;
  assign new_n614_ = pj & new_n613_;
  assign new_n615_ = pf & new_n230_;
  assign new_n616_ = new_n433_ & new_n615_;
  assign new_n617_ = ~ph & new_n616_;
  assign new_n618_ = pj & new_n617_;
  assign new_n619_ = new_n374_ & new_n448_;
  assign new_n620_ = ~ph & new_n619_;
  assign new_n621_ = new_n53_ & new_n620_;
  assign new_n622_ = pj & new_n621_;
  assign new_n623_ = new_n323_ & new_n511_;
  assign new_n624_ = pj & new_n623_;
  assign new_n625_ = ph & new_n339_;
  assign new_n626_ = ~new_n411_ & new_n625_;
  assign new_n627_ = pj & new_n626_;
  assign new_n628_ = ~new_n624_ & ~new_n627_;
  assign new_n629_ = ~new_n614_ & ~new_n618_;
  assign new_n630_ = ~new_n622_ & new_n629_;
  assign new_n631_ = new_n628_ & new_n630_;
  assign new_n632_ = ~new_n607_ & ~new_n610_;
  assign new_n633_ = ~new_n597_ & ~new_n602_;
  assign new_n634_ = ~new_n603_ & new_n633_;
  assign new_n635_ = new_n632_ & new_n634_;
  assign new_n636_ = new_n631_ & new_n635_;
  assign new_n637_ = ~new_n569_ & ~new_n571_;
  assign new_n638_ = ~new_n564_ & ~new_n567_;
  assign new_n639_ = ~new_n198_ & new_n638_;
  assign new_n640_ = new_n637_ & new_n639_;
  assign new_n641_ = ~new_n587_ & ~new_n592_;
  assign new_n642_ = ~new_n576_ & ~new_n581_;
  assign new_n643_ = ~new_n582_ & new_n642_;
  assign new_n644_ = new_n641_ & new_n643_;
  assign new_n645_ = new_n640_ & new_n644_;
  assign po = ~new_n636_ | ~new_n645_;
endmodule

