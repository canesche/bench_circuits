module top ( 
    pp, pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0, pw, px,
    py, pz, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn, po,
    ph0, pi0, pj0, pk0, pl0, pm0, pn0, po0, pp0, pq0, pr0, ps0, pt0, pu0,
    pv0, pw0, px0  );
  input  pp, pa0, pq, pb0, pr, pc0, ps, pd0, pt, pe0, pu, pf0, pv, pg0,
    pw, px, py, pz, pa, pb, pc, pd, pe, pf, pg, ph, pi, pj, pk, pl, pm, pn,
    po;
  output ph0, pi0, pj0, pk0, pl0, pm0, pn0, po0, pp0, pq0, pr0, ps0, pt0, pu0,
    pv0, pw0, px0;
  wire new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_,
    new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_,
    new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n117_,
    new_n118_, new_n119_, new_n120_, new_n121_, new_n122_, new_n123_,
    new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_,
    new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n287_, new_n288_, new_n289_;
  assign new_n51_ = ~pp & ~pg0;
  assign new_n52_ = ~pf0 & ~pg0;
  assign new_n53_ = ~pp & ~pf0;
  assign new_n54_ = ~new_n51_ & ~new_n52_;
  assign new_n55_ = ~new_n53_ & new_n54_;
  assign new_n56_ = ~po & ~new_n55_;
  assign new_n57_ = ~pe0 & ~new_n55_;
  assign new_n58_ = ~pe0 & ~po;
  assign new_n59_ = ~new_n56_ & ~new_n57_;
  assign new_n60_ = ~new_n58_ & new_n59_;
  assign new_n61_ = ~pn & ~new_n60_;
  assign new_n62_ = ~pd0 & ~new_n60_;
  assign new_n63_ = ~pd0 & ~pn;
  assign new_n64_ = ~new_n61_ & ~new_n62_;
  assign new_n65_ = ~new_n63_ & new_n64_;
  assign new_n66_ = ~pm & ~new_n65_;
  assign new_n67_ = ~pc0 & ~new_n65_;
  assign new_n68_ = ~pc0 & ~pm;
  assign new_n69_ = ~new_n66_ & ~new_n67_;
  assign new_n70_ = ~new_n68_ & new_n69_;
  assign new_n71_ = ~pl & ~new_n70_;
  assign new_n72_ = ~pb0 & ~new_n70_;
  assign new_n73_ = ~pb0 & ~pl;
  assign new_n74_ = ~new_n71_ & ~new_n72_;
  assign new_n75_ = ~new_n73_ & new_n74_;
  assign new_n76_ = ~pk & ~new_n75_;
  assign new_n77_ = ~pa0 & ~new_n75_;
  assign new_n78_ = ~pa0 & ~pk;
  assign new_n79_ = ~new_n76_ & ~new_n77_;
  assign new_n80_ = ~new_n78_ & new_n79_;
  assign new_n81_ = ~pj & ~new_n80_;
  assign new_n82_ = ~pz & ~new_n80_;
  assign new_n83_ = ~pz & ~pj;
  assign new_n84_ = ~new_n81_ & ~new_n82_;
  assign new_n85_ = ~new_n83_ & new_n84_;
  assign new_n86_ = ~pi & ~new_n85_;
  assign new_n87_ = ~py & ~new_n85_;
  assign new_n88_ = ~py & ~pi;
  assign new_n89_ = ~new_n86_ & ~new_n87_;
  assign new_n90_ = ~new_n88_ & new_n89_;
  assign new_n91_ = ~ph & ~new_n90_;
  assign new_n92_ = ~px & ~new_n90_;
  assign new_n93_ = ~px & ~ph;
  assign new_n94_ = ~new_n91_ & ~new_n92_;
  assign new_n95_ = ~new_n93_ & new_n94_;
  assign new_n96_ = ~pg & ~new_n95_;
  assign new_n97_ = ~pw & ~new_n95_;
  assign new_n98_ = ~pw & ~pg;
  assign new_n99_ = ~new_n96_ & ~new_n97_;
  assign new_n100_ = ~new_n98_ & new_n99_;
  assign new_n101_ = ~pf & ~new_n100_;
  assign new_n102_ = ~pv & ~new_n100_;
  assign new_n103_ = ~pv & ~pf;
  assign new_n104_ = ~new_n101_ & ~new_n102_;
  assign new_n105_ = ~new_n103_ & new_n104_;
  assign new_n106_ = ~pe & ~new_n105_;
  assign new_n107_ = ~pu & ~new_n105_;
  assign new_n108_ = ~pu & ~pe;
  assign new_n109_ = ~new_n106_ & ~new_n107_;
  assign new_n110_ = ~new_n108_ & new_n109_;
  assign new_n111_ = ~pd & ~new_n110_;
  assign new_n112_ = ~pt & ~new_n110_;
  assign new_n113_ = ~pt & ~pd;
  assign new_n114_ = ~new_n111_ & ~new_n112_;
  assign new_n115_ = ~new_n113_ & new_n114_;
  assign new_n116_ = ~pc & ~new_n115_;
  assign new_n117_ = ~ps & ~new_n115_;
  assign new_n118_ = ~ps & ~pc;
  assign new_n119_ = ~new_n116_ & ~new_n117_;
  assign new_n120_ = ~new_n118_ & new_n119_;
  assign new_n121_ = ~pb & ~new_n120_;
  assign new_n122_ = ~pr & ~new_n120_;
  assign new_n123_ = ~pr & ~pb;
  assign new_n124_ = ~new_n121_ & ~new_n122_;
  assign new_n125_ = ~new_n123_ & new_n124_;
  assign new_n126_ = ~pq & new_n125_;
  assign new_n127_ = pa & new_n126_;
  assign new_n128_ = ~pq & ~new_n125_;
  assign new_n129_ = ~pa & new_n128_;
  assign new_n130_ = pq & new_n125_;
  assign new_n131_ = ~pa & new_n130_;
  assign new_n132_ = pq & ~new_n125_;
  assign new_n133_ = pa & new_n132_;
  assign new_n134_ = ~new_n131_ & ~new_n133_;
  assign new_n135_ = ~new_n127_ & ~new_n129_;
  assign ph0 = new_n134_ & new_n135_;
  assign new_n137_ = ~pr & new_n120_;
  assign new_n138_ = pb & new_n137_;
  assign new_n139_ = ~pb & new_n122_;
  assign new_n140_ = pr & new_n120_;
  assign new_n141_ = ~pb & new_n140_;
  assign new_n142_ = pr & ~new_n120_;
  assign new_n143_ = pb & new_n142_;
  assign new_n144_ = ~new_n141_ & ~new_n143_;
  assign new_n145_ = ~new_n138_ & ~new_n139_;
  assign pi0 = new_n144_ & new_n145_;
  assign new_n147_ = ~ps & new_n115_;
  assign new_n148_ = pc & new_n147_;
  assign new_n149_ = ~pc & new_n117_;
  assign new_n150_ = ps & new_n115_;
  assign new_n151_ = ~pc & new_n150_;
  assign new_n152_ = ps & ~new_n115_;
  assign new_n153_ = pc & new_n152_;
  assign new_n154_ = ~new_n151_ & ~new_n153_;
  assign new_n155_ = ~new_n148_ & ~new_n149_;
  assign pj0 = new_n154_ & new_n155_;
  assign new_n157_ = ~pt & new_n110_;
  assign new_n158_ = pd & new_n157_;
  assign new_n159_ = ~pd & new_n112_;
  assign new_n160_ = pt & new_n110_;
  assign new_n161_ = ~pd & new_n160_;
  assign new_n162_ = pt & ~new_n110_;
  assign new_n163_ = pd & new_n162_;
  assign new_n164_ = ~new_n161_ & ~new_n163_;
  assign new_n165_ = ~new_n158_ & ~new_n159_;
  assign pk0 = new_n164_ & new_n165_;
  assign new_n167_ = ~pu & new_n105_;
  assign new_n168_ = pe & new_n167_;
  assign new_n169_ = ~pe & new_n107_;
  assign new_n170_ = pu & new_n105_;
  assign new_n171_ = ~pe & new_n170_;
  assign new_n172_ = pu & ~new_n105_;
  assign new_n173_ = pe & new_n172_;
  assign new_n174_ = ~new_n171_ & ~new_n173_;
  assign new_n175_ = ~new_n168_ & ~new_n169_;
  assign pl0 = new_n174_ & new_n175_;
  assign new_n177_ = ~pv & new_n100_;
  assign new_n178_ = pf & new_n177_;
  assign new_n179_ = ~pf & new_n102_;
  assign new_n180_ = pv & new_n100_;
  assign new_n181_ = ~pf & new_n180_;
  assign new_n182_ = pv & ~new_n100_;
  assign new_n183_ = pf & new_n182_;
  assign new_n184_ = ~new_n181_ & ~new_n183_;
  assign new_n185_ = ~new_n178_ & ~new_n179_;
  assign pm0 = new_n184_ & new_n185_;
  assign new_n187_ = ~pw & new_n95_;
  assign new_n188_ = pg & new_n187_;
  assign new_n189_ = ~pg & new_n97_;
  assign new_n190_ = pw & new_n95_;
  assign new_n191_ = ~pg & new_n190_;
  assign new_n192_ = pw & ~new_n95_;
  assign new_n193_ = pg & new_n192_;
  assign new_n194_ = ~new_n191_ & ~new_n193_;
  assign new_n195_ = ~new_n188_ & ~new_n189_;
  assign pn0 = new_n194_ & new_n195_;
  assign new_n197_ = ~px & new_n90_;
  assign new_n198_ = ph & new_n197_;
  assign new_n199_ = ~ph & new_n92_;
  assign new_n200_ = px & new_n90_;
  assign new_n201_ = ~ph & new_n200_;
  assign new_n202_ = px & ~new_n90_;
  assign new_n203_ = ph & new_n202_;
  assign new_n204_ = ~new_n201_ & ~new_n203_;
  assign new_n205_ = ~new_n198_ & ~new_n199_;
  assign po0 = new_n204_ & new_n205_;
  assign new_n207_ = ~py & new_n85_;
  assign new_n208_ = pi & new_n207_;
  assign new_n209_ = ~pi & new_n87_;
  assign new_n210_ = py & new_n85_;
  assign new_n211_ = ~pi & new_n210_;
  assign new_n212_ = py & ~new_n85_;
  assign new_n213_ = pi & new_n212_;
  assign new_n214_ = ~new_n211_ & ~new_n213_;
  assign new_n215_ = ~new_n208_ & ~new_n209_;
  assign pp0 = new_n214_ & new_n215_;
  assign new_n217_ = ~pz & new_n80_;
  assign new_n218_ = pj & new_n217_;
  assign new_n219_ = ~pj & new_n82_;
  assign new_n220_ = pz & new_n80_;
  assign new_n221_ = ~pj & new_n220_;
  assign new_n222_ = pz & ~new_n80_;
  assign new_n223_ = pj & new_n222_;
  assign new_n224_ = ~new_n221_ & ~new_n223_;
  assign new_n225_ = ~new_n218_ & ~new_n219_;
  assign pq0 = new_n224_ & new_n225_;
  assign new_n227_ = ~pa0 & new_n75_;
  assign new_n228_ = pk & new_n227_;
  assign new_n229_ = ~pk & new_n77_;
  assign new_n230_ = pa0 & new_n75_;
  assign new_n231_ = ~pk & new_n230_;
  assign new_n232_ = pa0 & ~new_n75_;
  assign new_n233_ = pk & new_n232_;
  assign new_n234_ = ~new_n231_ & ~new_n233_;
  assign new_n235_ = ~new_n228_ & ~new_n229_;
  assign pr0 = new_n234_ & new_n235_;
  assign new_n237_ = ~pb0 & new_n70_;
  assign new_n238_ = pl & new_n237_;
  assign new_n239_ = ~pl & new_n72_;
  assign new_n240_ = pb0 & new_n70_;
  assign new_n241_ = ~pl & new_n240_;
  assign new_n242_ = pb0 & ~new_n70_;
  assign new_n243_ = pl & new_n242_;
  assign new_n244_ = ~new_n241_ & ~new_n243_;
  assign new_n245_ = ~new_n238_ & ~new_n239_;
  assign ps0 = new_n244_ & new_n245_;
  assign new_n247_ = ~pc0 & new_n65_;
  assign new_n248_ = pm & new_n247_;
  assign new_n249_ = ~pm & new_n67_;
  assign new_n250_ = pc0 & new_n65_;
  assign new_n251_ = ~pm & new_n250_;
  assign new_n252_ = pc0 & ~new_n65_;
  assign new_n253_ = pm & new_n252_;
  assign new_n254_ = ~new_n251_ & ~new_n253_;
  assign new_n255_ = ~new_n248_ & ~new_n249_;
  assign pt0 = new_n254_ & new_n255_;
  assign new_n257_ = ~pd0 & new_n60_;
  assign new_n258_ = pn & new_n257_;
  assign new_n259_ = ~pn & new_n62_;
  assign new_n260_ = pd0 & new_n60_;
  assign new_n261_ = ~pn & new_n260_;
  assign new_n262_ = pd0 & ~new_n60_;
  assign new_n263_ = pn & new_n262_;
  assign new_n264_ = ~new_n261_ & ~new_n263_;
  assign new_n265_ = ~new_n258_ & ~new_n259_;
  assign pu0 = new_n264_ & new_n265_;
  assign new_n267_ = ~pe0 & new_n55_;
  assign new_n268_ = po & new_n267_;
  assign new_n269_ = ~po & new_n57_;
  assign new_n270_ = pe0 & new_n55_;
  assign new_n271_ = ~po & new_n270_;
  assign new_n272_ = pe0 & ~new_n55_;
  assign new_n273_ = po & new_n272_;
  assign new_n274_ = ~new_n271_ & ~new_n273_;
  assign new_n275_ = ~new_n268_ & ~new_n269_;
  assign pv0 = new_n274_ & new_n275_;
  assign new_n277_ = ~pp & new_n52_;
  assign new_n278_ = ~pf0 & pg0;
  assign new_n279_ = pp & new_n278_;
  assign new_n280_ = pf0 & ~pg0;
  assign new_n281_ = pp & new_n280_;
  assign new_n282_ = pf0 & pg0;
  assign new_n283_ = ~pp & new_n282_;
  assign new_n284_ = ~new_n281_ & ~new_n283_;
  assign new_n285_ = ~new_n277_ & ~new_n279_;
  assign pw0 = new_n284_ & new_n285_;
  assign new_n287_ = ~pa & ~new_n125_;
  assign new_n288_ = ~pq & ~pa;
  assign new_n289_ = ~new_n128_ & ~new_n287_;
  assign px0 = ~new_n288_ & new_n289_;
endmodule

